

module b17_C_SARLock_k_128_10 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, U355, U356, U357, U358, U359, U360, U361, 
        U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, 
        U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, U376, U247, 
        U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, 
        U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223, 
        U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254, U255, 
        U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, 
        U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, 
        U280, U281, U282, U212, U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, 
        P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, 
        P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, 
        P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, 
        P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, 
        P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, 
        P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, 
        P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, 
        P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, 
        P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, 
        P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, 
        P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, 
        P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, 
        P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, 
        P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, 
        P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, 
        P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, 
        P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, 
        P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, 
        P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, 
        P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, 
        P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, 
        P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, 
        P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, 
        P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, 
        P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, 
        P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, 
        P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, 
        P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, 
        P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, 
        P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, 
        P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, 
        P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, 
        P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, 
        P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, 
        P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, 
        P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, 
        P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, 
        P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, 
        P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, 
        P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, 
        P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, 
        P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, 
        P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, 
        P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, 
        P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, 
        P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, 
        P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, 
        P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, 
        P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, 
        P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, 
        P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, 
        P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, 
        P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, 
        P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, 
        P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, 
        P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, 
        P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, 
        P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, 
        P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, 
        P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, 
        P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, 
        P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, 
        P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, 
        P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, 
        P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, 
        P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, 
        P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, 
        P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, 
        P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, 
        P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, 
        P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, 
        P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, 
        P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, 
        P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, 
        P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, 
        P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, 
        P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, 
        P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, 
        P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, 
        P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, 
        P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, 
        P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, 
        P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, 
        P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, 
        P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, 
        P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, 
        P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, 
        P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, 
        P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, 
        P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, 
        P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, 
        P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, 
        P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, 
        P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, 
        P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, 
        P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, 
        P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, 
        P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, 
        P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, 
        P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, 
        P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, 
        P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, 
        P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, 
        P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, 
        P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, 
        P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, 
        P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, 
        P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, 
        P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, 
        P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, 
        P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, 
        P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, 
        P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, 
        P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, 
        P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, 
        P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, 
        P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, 
        P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, 
        P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, 
        P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, 
        P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, 
        P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, 
        P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, 
        P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, 
        P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, 
        P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, 
        P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, 
        P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, 
        P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, 
        P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, 
        P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, 
        P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, 
        P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, 
        P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, 
        P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, 
        P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, 
        P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, 
        P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, 
        P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, 
        P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, 
        P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, 
        P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, 
        P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, 
        P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, 
        P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, 
        P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, 
        P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, 
        P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, 
        P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, 
        P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, 
        P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, 
        P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, 
        P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, 
        P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, 
        P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, 
        P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, 
        P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, 
        P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, 
        P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, 
        P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, 
        P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, 
        P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, 
        P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, 
        P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, 
        P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, 
        P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, 
        P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, 
        P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, 
        P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, 
        P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, 
        P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, 
        P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, 
        P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, 
        P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, 
        P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, 
        P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, 
        P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, 
        P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801
 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9720, n9721, n9722, n9723, n9724, n9725, n9727, n9728, n9729, n9730,
         n9731, n9734, n9735, n9736, n9737, n9738, n9740, n9741, n9743, n9744,
         n9745, n9746, n9747, n9748, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
         n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
         n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
         n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654,
         n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662,
         n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
         n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
         n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702,
         n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
         n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718,
         n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
         n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
         n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
         n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750,
         n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
         n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766,
         n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
         n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782,
         n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
         n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798,
         n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806,
         n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
         n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822,
         n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
         n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838,
         n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
         n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
         n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
         n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870,
         n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
         n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
         n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894,
         n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
         n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910,
         n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918,
         n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926,
         n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
         n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942,
         n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
         n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
         n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966,
         n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
         n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982,
         n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990,
         n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998,
         n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
         n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014,
         n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
         n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030,
         n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038,
         n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046,
         n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054,
         n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062,
         n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070,
         n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078,
         n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086,
         n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094,
         n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102,
         n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110,
         n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
         n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126,
         n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134,
         n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142,
         n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150,
         n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158,
         n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
         n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
         n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182,
         n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
         n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198,
         n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206,
         n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214,
         n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222,
         n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230,
         n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
         n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246,
         n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254,
         n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262,
         n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270,
         n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278,
         n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286,
         n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294,
         n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302,
         n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
         n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
         n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326,
         n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
         n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342,
         n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358,
         n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
         n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
         n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
         n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
         n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
         n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
         n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
         n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
         n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
         n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
         n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
         n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
         n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462,
         n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
         n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
         n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486,
         n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494,
         n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502,
         n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510,
         n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518,
         n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526,
         n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
         n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542,
         n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550,
         n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558,
         n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566,
         n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
         n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598,
         n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
         n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614,
         n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622,
         n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630,
         n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638,
         n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646,
         n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654,
         n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662,
         n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670,
         n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
         n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686,
         n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694,
         n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702,
         n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710,
         n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
         n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726,
         n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734,
         n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742,
         n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750,
         n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758,
         n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
         n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774,
         n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
         n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
         n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798,
         n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806,
         n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814,
         n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822,
         n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830,
         n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838,
         n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846,
         n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854,
         n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
         n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870,
         n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878,
         n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886,
         n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
         n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
         n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
         n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
         n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926,
         n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934,
         n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942,
         n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950,
         n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
         n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
         n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974,
         n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
         n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
         n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998,
         n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006,
         n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014,
         n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022,
         n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030,
         n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
         n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046,
         n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054,
         n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
         n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070,
         n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078,
         n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086,
         n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094,
         n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102,
         n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110,
         n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118,
         n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126,
         n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134,
         n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142,
         n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150,
         n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158,
         n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166,
         n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
         n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182,
         n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190,
         n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
         n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206,
         n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214,
         n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222,
         n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230,
         n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238,
         n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246,
         n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
         n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262,
         n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
         n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278,
         n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286,
         n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294,
         n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302,
         n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310,
         n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326,
         n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334,
         n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350,
         n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358,
         n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
         n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
         n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
         n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390,
         n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
         n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
         n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422,
         n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
         n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
         n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454,
         n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462,
         n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470,
         n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478,
         n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
         n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
         n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502,
         n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510,
         n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
         n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
         n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534,
         n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
         n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
         n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
         n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566,
         n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
         n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
         n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638,
         n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646,
         n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
         n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
         n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
         n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
         n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
         n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
         n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
         n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
         n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
         n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286,
         n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
         n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
         n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
         n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358,
         n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366,
         n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374,
         n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
         n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
         n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398,
         n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
         n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414,
         n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422,
         n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430,
         n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438,
         n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446,
         n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
         n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462,
         n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470,
         n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
         n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
         n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
         n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
         n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510,
         n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518,
         n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
         n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
         n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542,
         n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
         n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
         n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
         n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574,
         n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582,
         n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
         n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
         n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
         n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614,
         n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
         n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630,
         n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
         n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
         n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654,
         n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662,
         n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
         n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678,
         n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686,
         n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
         n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702,
         n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
         n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718,
         n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726,
         n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734,
         n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
         n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750,
         n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758,
         n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
         n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774,
         n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782,
         n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
         n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798,
         n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806,
         n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814,
         n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822,
         n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830,
         n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
         n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846,
         n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870,
         n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878,
         n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
         n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894,
         n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902,
         n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
         n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918,
         n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926,
         n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934,
         n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942,
         n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950,
         n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
         n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966,
         n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974,
         n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
         n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990,
         n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
         n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006,
         n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014,
         n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022,
         n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030,
         n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038,
         n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046,
         n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
         n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062,
         n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
         n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078,
         n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086,
         n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094,
         n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
         n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110,
         n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118,
         n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
         n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134,
         n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
         n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150,
         n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158,
         n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166,
         n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
         n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182,
         n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190,
         n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
         n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
         n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214,
         n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222,
         n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230,
         n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238,
         n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
         n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254,
         n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262,
         n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
         n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278,
         n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286,
         n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294,
         n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302,
         n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310,
         n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
         n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326,
         n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334,
         n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342,
         n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350,
         n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358,
         n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366,
         n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374,
         n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382,
         n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
         n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398,
         n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406,
         n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
         n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422,
         n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430,
         n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438,
         n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446,
         n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454,
         n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
         n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470,
         n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478,
         n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486,
         n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494,
         n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502,
         n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510,
         n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518,
         n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526,
         n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
         n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542,
         n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550,
         n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
         n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566,
         n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574,
         n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582,
         n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
         n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
         n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
         n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614,
         n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
         n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
         n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
         n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
         n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
         n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
         n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
         n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
         n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
         n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758,
         n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
         n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
         n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
         n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
         n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
         n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806,
         n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
         n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
         n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830,
         n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838,
         n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
         n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
         n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
         n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
         n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
         n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
         n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926,
         n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
         n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
         n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
         n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
         n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
         n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
         n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
         n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
         n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
         n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
         n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
         n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
         n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
         n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
         n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
         n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
         n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
         n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
         n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
         n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
         n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
         n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
         n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
         n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
         n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790,
         n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
         n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806,
         n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814,
         n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
         n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
         n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838,
         n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846,
         n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
         n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862,
         n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
         n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878,
         n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886,
         n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
         n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
         n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910,
         n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918,
         n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
         n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934,
         n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942,
         n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950,
         n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958,
         n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
         n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
         n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982,
         n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990,
         n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998,
         n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006,
         n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014,
         n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022,
         n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030,
         n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038,
         n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
         n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054,
         n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062,
         n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070,
         n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078,
         n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086,
         n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094,
         n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102,
         n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110,
         n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118,
         n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126,
         n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134,
         n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142,
         n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150,
         n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158,
         n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166,
         n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174,
         n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182,
         n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190,
         n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198,
         n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206,
         n21207;

  AOI21_X1 U11165 ( .B1(n13913), .B2(n9787), .A(n13912), .ZN(n14296) );
  OAI21_X1 U11166 ( .B1(n13952), .B2(n13953), .A(n13939), .ZN(n14326) );
  INV_X1 U11167 ( .A(n20027), .ZN(n20016) );
  NAND2_X1 U11168 ( .A1(n14323), .A2(n14333), .ZN(n14322) );
  NOR2_X1 U11169 ( .A1(n17436), .A2(n17253), .ZN(n17248) );
  AND2_X1 U11170 ( .A1(n14828), .A2(n12369), .ZN(n14815) );
  NAND2_X1 U11171 ( .A1(n9908), .A2(n18835), .ZN(n18658) );
  NAND2_X1 U11172 ( .A1(n10116), .A2(n9764), .ZN(n14444) );
  NAND2_X1 U11173 ( .A1(n10126), .A2(n12512), .ZN(n10125) );
  BUF_X1 U11174 ( .A(n12089), .Z(n19002) );
  INV_X1 U11175 ( .A(n16815), .ZN(n16852) );
  NAND2_X1 U11176 ( .A1(n20114), .A2(n20113), .ZN(n20112) );
  NOR4_X2 U11177 ( .A1(n15560), .A2(n15586), .A3(n15564), .A4(n18183), .ZN(
        n17416) );
  NAND2_X1 U11178 ( .A1(n12474), .A2(n12425), .ZN(n12502) );
  CLKBUF_X2 U11179 ( .A(n10736), .Z(n10762) );
  CLKBUF_X2 U11180 ( .A(n10733), .Z(n10847) );
  CLKBUF_X2 U11181 ( .A(n10765), .Z(n10848) );
  INV_X1 U11182 ( .A(n18835), .ZN(n16523) );
  NOR2_X1 U11183 ( .A1(n10484), .A2(n10491), .ZN(n19442) );
  XNOR2_X1 U11184 ( .A(n11343), .B(n11312), .ZN(n12426) );
  NAND2_X1 U11185 ( .A1(n11215), .A2(n11214), .ZN(n11312) );
  INV_X1 U11186 ( .A(n12253), .ZN(n12260) );
  OR2_X1 U11187 ( .A1(n11218), .A2(n11217), .ZN(n11247) );
  INV_X2 U11188 ( .A(n11016), .ZN(n10102) );
  CLKBUF_X3 U11189 ( .A(n15647), .Z(n17166) );
  BUF_X2 U11190 ( .A(n9727), .Z(n17146) );
  BUF_X2 U11191 ( .A(n15491), .Z(n17049) );
  CLKBUF_X2 U11193 ( .A(n15401), .Z(n9727) );
  INV_X2 U11194 ( .A(n15694), .ZN(n17118) );
  INV_X1 U11195 ( .A(n15669), .ZN(n17153) );
  INV_X1 U11196 ( .A(n9776), .ZN(n17170) );
  CLKBUF_X2 U11197 ( .A(n11176), .Z(n11460) );
  AND2_X1 U11198 ( .A1(n10518), .A2(n12956), .ZN(n10580) );
  AND2_X1 U11199 ( .A1(n13884), .A2(n12956), .ZN(n10581) );
  AND2_X1 U11200 ( .A1(n10518), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10607) );
  AND2_X1 U11201 ( .A1(n10510), .A2(n10511), .ZN(n10546) );
  NAND2_X1 U11202 ( .A1(n18803), .A2(n18793), .ZN(n15388) );
  NOR2_X1 U11203 ( .A1(n12623), .A2(n11131), .ZN(n11132) );
  BUF_X2 U11204 ( .A(n10512), .Z(n13886) );
  CLKBUF_X1 U11205 ( .A(n10399), .Z(n19243) );
  BUF_X1 U11207 ( .A(n10409), .Z(n16300) );
  AND2_X4 U11208 ( .A1(n11044), .A2(n11045), .ZN(n11168) );
  CLKBUF_X1 U11209 ( .A(n10385), .Z(n19223) );
  AND2_X1 U11210 ( .A1(n12780), .A2(n11035), .ZN(n11547) );
  AND2_X1 U11211 ( .A1(n11046), .A2(n13150), .ZN(n9745) );
  INV_X1 U11212 ( .A(n11827), .ZN(n11789) );
  INV_X1 U11213 ( .A(n9779), .ZN(n11820) );
  INV_X1 U11214 ( .A(n12773), .ZN(n14646) );
  NAND2_X1 U11215 ( .A1(n13151), .A2(n10031), .ZN(n11815) );
  NAND2_X1 U11216 ( .A1(n12780), .A2(n11044), .ZN(n11827) );
  NAND2_X1 U11217 ( .A1(n13151), .A2(n11028), .ZN(n11700) );
  NAND4_X1 U11218 ( .A1(n11027), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A4(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11787) );
  AND3_X1 U11219 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13147) );
  NOR2_X2 U11220 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12777) );
  NAND2_X1 U11221 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12773) );
  NOR2_X2 U11222 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13151) );
  OAI21_X1 U11223 ( .B1(n14376), .B2(n12518), .A(n15923), .ZN(n9720) );
  INV_X1 U11224 ( .A(n14361), .ZN(n9721) );
  OAI21_X1 U11225 ( .B1(n14376), .B2(n12518), .A(n15923), .ZN(n14371) );
  NAND2_X1 U11226 ( .A1(n9858), .A2(n14370), .ZN(n14308) );
  XNOR2_X2 U11228 ( .A(n14304), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14482) );
  NAND2_X2 U11229 ( .A1(n11226), .A2(n11225), .ZN(n11252) );
  CLKBUF_X1 U11230 ( .A(n18690), .Z(n9722) );
  NOR2_X1 U11231 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18787), .ZN(n18690) );
  NOR2_X1 U11232 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10279) );
  INV_X1 U11233 ( .A(n11813), .ZN(n11790) );
  CLKBUF_X2 U11234 ( .A(n13621), .Z(n9728) );
  AND2_X1 U11235 ( .A1(n13885), .A2(n12956), .ZN(n12959) );
  INV_X1 U11236 ( .A(n15672), .ZN(n15682) );
  INV_X1 U11237 ( .A(n14409), .ZN(n10122) );
  AND2_X1 U11238 ( .A1(n11052), .A2(n11051), .ZN(n11139) );
  NAND2_X1 U11239 ( .A1(n20112), .A2(n12462), .ZN(n15954) );
  NAND2_X1 U11240 ( .A1(n11100), .A2(n10272), .ZN(n20184) );
  INV_X1 U11241 ( .A(n11139), .ZN(n11204) );
  INV_X1 U11242 ( .A(n9783), .ZN(n17037) );
  NOR2_X1 U11243 ( .A1(n17375), .A2(n17855), .ZN(n15710) );
  NAND2_X1 U11244 ( .A1(n18818), .A2(n18811), .ZN(n16884) );
  INV_X1 U11245 ( .A(n15458), .ZN(n17107) );
  AND4_X1 U11246 ( .A1(n11061), .A2(n11060), .A3(n11059), .A4(n11058), .ZN(
        n9784) );
  OAI21_X1 U11247 ( .B1(n20162), .B2(n10179), .A(n11354), .ZN(n13199) );
  OAI21_X1 U11248 ( .B1(n10122), .B2(n10040), .A(n10120), .ZN(n14376) );
  NAND2_X1 U11251 ( .A1(n11346), .A2(n11356), .ZN(n20162) );
  NAND2_X1 U11252 ( .A1(n11320), .A2(n11319), .ZN(n20247) );
  OR2_X1 U11253 ( .A1(n16065), .A2(n16064), .ZN(n9998) );
  AND2_X1 U11254 ( .A1(n9731), .A2(n12626), .ZN(n13357) );
  NAND2_X2 U11255 ( .A1(n9784), .A2(n9848), .ZN(n20209) );
  NOR2_X2 U11256 ( .A1(n12064), .A2(n14960), .ZN(n12063) );
  NOR2_X1 U11257 ( .A1(n12074), .A2(n15041), .ZN(n12075) );
  INV_X1 U11258 ( .A(n17579), .ZN(n17766) );
  INV_X1 U11259 ( .A(n19980), .ZN(n19996) );
  AOI211_X1 U11260 ( .C1(n15932), .C2(n14329), .A(n14328), .B(n14327), .ZN(
        n14330) );
  INV_X1 U11261 ( .A(n9724), .ZN(n17375) );
  NOR2_X1 U11262 ( .A1(n20184), .A2(n20189), .ZN(n13180) );
  INV_X1 U11263 ( .A(n20184), .ZN(n12974) );
  NOR2_X4 U11264 ( .A1(n14738), .A2(n14737), .ZN(n14740) );
  AND2_X1 U11265 ( .A1(n14646), .A2(n12777), .ZN(n9723) );
  AND2_X2 U11266 ( .A1(n10418), .A2(n10417), .ZN(n12364) );
  NAND2_X1 U11267 ( .A1(n14733), .A2(n14736), .ZN(n14735) );
  XNOR2_X1 U11268 ( .A(n13760), .B(n13761), .ZN(n14733) );
  NAND2_X2 U11269 ( .A1(n13322), .A2(n9961), .ZN(n9960) );
  INV_X1 U11270 ( .A(n11929), .ZN(n13179) );
  NOR2_X2 U11271 ( .A1(n11929), .A2(n13909), .ZN(n12004) );
  AOI21_X2 U11274 ( .B1(n15018), .B2(n15015), .A(n14945), .ZN(n15009) );
  XNOR2_X2 U11275 ( .A(n10940), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15008) );
  NOR2_X2 U11276 ( .A1(n17976), .A2(n17755), .ZN(n17661) );
  NOR3_X2 U11278 ( .A1(n16796), .A2(n17188), .A3(n17187), .ZN(n17186) );
  NOR2_X2 U11279 ( .A1(n15407), .A2(n15406), .ZN(n18183) );
  NOR2_X1 U11280 ( .A1(n15386), .A2(n15385), .ZN(n15401) );
  AND2_X4 U11281 ( .A1(n13832), .A2(n19576), .ZN(n12253) );
  INV_X4 U11282 ( .A(n16316), .ZN(n13832) );
  AND2_X1 U11283 ( .A1(n13878), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13621) );
  AOI21_X2 U11284 ( .B1(n15009), .B2(n15008), .A(n14947), .ZN(n14999) );
  OAI21_X1 U11285 ( .B1(n14735), .B2(n10247), .A(n10245), .ZN(n10243) );
  NAND2_X1 U11286 ( .A1(n14322), .A2(n10052), .ZN(n10054) );
  AOI21_X1 U11287 ( .B1(n14935), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n14933), .ZN(n9922) );
  NAND2_X1 U11288 ( .A1(n10990), .A2(n10989), .ZN(n14935) );
  NAND2_X1 U11289 ( .A1(n9926), .A2(n10915), .ZN(n15293) );
  CLKBUF_X1 U11290 ( .A(n14376), .Z(n14601) );
  CLKBUF_X1 U11291 ( .A(n14409), .Z(n15936) );
  NOR2_X1 U11292 ( .A1(n9778), .A2(n14766), .ZN(n14767) );
  OAI21_X1 U11293 ( .B1(n10659), .B2(n9924), .A(n18998), .ZN(n10886) );
  NAND2_X1 U11295 ( .A1(n9920), .A2(n9919), .ZN(n10658) );
  AND2_X1 U11296 ( .A1(n15203), .A2(n9832), .ZN(n15156) );
  NOR2_X1 U11297 ( .A1(n10644), .A2(n12132), .ZN(n9920) );
  OAI21_X1 U11298 ( .B1(n10973), .B2(n9977), .A(n10972), .ZN(n9976) );
  NAND2_X1 U11299 ( .A1(n10138), .A2(n10573), .ZN(n10644) );
  NOR2_X1 U11300 ( .A1(n17976), .A2(n17974), .ZN(n17577) );
  AOI22_X1 U11301 ( .A1(n18027), .A2(n17848), .B1(n17766), .B2(n18029), .ZN(
        n17755) );
  OR2_X1 U11302 ( .A1(n10485), .A2(n10492), .ZN(n19544) );
  AND2_X1 U11303 ( .A1(n12847), .A2(n12898), .ZN(n12897) );
  INV_X1 U11304 ( .A(n12838), .ZN(n13322) );
  NOR2_X1 U11305 ( .A1(n13019), .A2(n12125), .ZN(n13078) );
  NAND2_X1 U11306 ( .A1(n14710), .A2(n10916), .ZN(n10926) );
  NOR2_X1 U11307 ( .A1(n9736), .A2(n18154), .ZN(n18149) );
  INV_X1 U11308 ( .A(n18057), .ZN(n18641) );
  CLKBUF_X2 U11309 ( .A(n12693), .Z(n12879) );
  NAND2_X1 U11310 ( .A1(n10403), .A2(n16319), .ZN(n13859) );
  AND2_X2 U11311 ( .A1(n12269), .A2(n13757), .ZN(n10765) );
  AND2_X1 U11312 ( .A1(n12848), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10733) );
  NOR2_X2 U11313 ( .A1(n12066), .A2(n15019), .ZN(n12067) );
  NAND2_X1 U11314 ( .A1(n12096), .A2(n16316), .ZN(n12241) );
  CLKBUF_X3 U11315 ( .A(n11152), .Z(n9729) );
  BUF_X2 U11316 ( .A(n10414), .Z(n19250) );
  AND2_X1 U11317 ( .A1(n10293), .A2(n10292), .ZN(n10413) );
  NAND2_X1 U11318 ( .A1(n10357), .A2(n10356), .ZN(n10399) );
  NAND2_X2 U11319 ( .A1(n11080), .A2(n10273), .ZN(n11155) );
  CLKBUF_X3 U11320 ( .A(n15648), .Z(n9734) );
  CLKBUF_X2 U11321 ( .A(n11057), .Z(n11800) );
  NOR2_X2 U11322 ( .A1(n15384), .A2(n16884), .ZN(n15533) );
  INV_X1 U11324 ( .A(n11232), .ZN(n11767) );
  INV_X2 U11325 ( .A(n11700), .ZN(n11729) );
  CLKBUF_X2 U11326 ( .A(n10509), .Z(n13880) );
  NOR2_X2 U11327 ( .A1(n16885), .A2(n15389), .ZN(n15645) );
  INV_X2 U11328 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11027) );
  INV_X2 U11329 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11038) );
  INV_X4 U11330 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12956) );
  AND2_X2 U11331 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10510) );
  AOI21_X1 U11332 ( .B1(n14726), .B2(n10249), .A(n14721), .ZN(n13838) );
  AND2_X1 U11333 ( .A1(n12385), .A2(n12384), .ZN(n12386) );
  NAND2_X1 U11334 ( .A1(n10244), .A2(n13788), .ZN(n10249) );
  NOR2_X1 U11335 ( .A1(n14291), .A2(n9852), .ZN(n14481) );
  NOR2_X1 U11336 ( .A1(n9853), .A2(n14475), .ZN(n9852) );
  AND2_X1 U11337 ( .A1(n9853), .A2(n14475), .ZN(n14291) );
  NAND2_X1 U11338 ( .A1(n12522), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9879) );
  OAI21_X1 U11339 ( .B1(n13763), .B2(n10247), .A(n14727), .ZN(n10246) );
  NAND2_X1 U11340 ( .A1(n10049), .A2(n10054), .ZN(n9853) );
  OR2_X1 U11341 ( .A1(n15302), .A2(n15310), .ZN(n15303) );
  NAND2_X1 U11342 ( .A1(n15320), .A2(n12372), .ZN(n15159) );
  NAND2_X1 U11343 ( .A1(n15293), .A2(n15290), .ZN(n15275) );
  NAND2_X1 U11344 ( .A1(n16203), .A2(n10692), .ZN(n15320) );
  NAND2_X1 U11345 ( .A1(n12520), .A2(n14411), .ZN(n14370) );
  NAND2_X1 U11346 ( .A1(n9917), .A2(n9822), .ZN(n9916) );
  OR2_X1 U11347 ( .A1(n14405), .A2(n9847), .ZN(n12520) );
  XNOR2_X1 U11348 ( .A(n10689), .B(n10687), .ZN(n15040) );
  INV_X1 U11349 ( .A(n9998), .ZN(n16063) );
  AND2_X1 U11350 ( .A1(n10041), .A2(n12501), .ZN(n9891) );
  NAND2_X1 U11351 ( .A1(n15052), .A2(n10211), .ZN(n15067) );
  AOI21_X1 U11352 ( .B1(n10123), .B2(n10125), .A(n10121), .ZN(n10120) );
  AND2_X1 U11353 ( .A1(n10664), .A2(n10643), .ZN(n10889) );
  NAND2_X1 U11354 ( .A1(n13503), .A2(n12499), .ZN(n10116) );
  NAND2_X1 U11355 ( .A1(n12494), .A2(n15947), .ZN(n13503) );
  NAND3_X1 U11356 ( .A1(n10141), .A2(n13438), .A3(n10139), .ZN(n13443) );
  XNOR2_X1 U11357 ( .A(n10886), .B(n13449), .ZN(n13437) );
  NOR2_X1 U11358 ( .A1(n12516), .A2(n15920), .ZN(n15909) );
  OAI22_X1 U11359 ( .A1(n14676), .A2(n9988), .B1(n19002), .B2(n16092), .ZN(
        n16090) );
  AND2_X1 U11360 ( .A1(n10118), .A2(n12484), .ZN(n10117) );
  INV_X1 U11361 ( .A(n9976), .ZN(n9975) );
  NOR2_X1 U11362 ( .A1(n10032), .A2(n14423), .ZN(n12513) );
  INV_X1 U11363 ( .A(n14404), .ZN(n10121) );
  NAND2_X1 U11364 ( .A1(n10644), .A2(n10645), .ZN(n9971) );
  NAND2_X1 U11365 ( .A1(n13195), .A2(n12454), .ZN(n20114) );
  AND2_X1 U11366 ( .A1(n10615), .A2(n10614), .ZN(n10657) );
  AND2_X1 U11367 ( .A1(n11384), .A2(n10155), .ZN(n10154) );
  NAND2_X1 U11368 ( .A1(n10137), .A2(n10526), .ZN(n10645) );
  AND2_X1 U11369 ( .A1(n12480), .A2(n12479), .ZN(n13422) );
  OR2_X1 U11370 ( .A1(n12486), .A2(n11311), .ZN(n10153) );
  INV_X2 U11371 ( .A(n12502), .ZN(n14411) );
  INV_X1 U11372 ( .A(n12502), .ZN(n14342) );
  OR2_X1 U11373 ( .A1(n10602), .A2(n10601), .ZN(n10615) );
  XNOR2_X1 U11374 ( .A(n12474), .B(n11306), .ZN(n12486) );
  OR2_X1 U11375 ( .A1(n11374), .A2(n11373), .ZN(n12474) );
  AND2_X1 U11376 ( .A1(n10496), .A2(n10497), .ZN(n19477) );
  AND2_X1 U11377 ( .A1(n10496), .A2(n10495), .ZN(n19510) );
  INV_X1 U11378 ( .A(n19544), .ZN(n9730) );
  OR2_X1 U11379 ( .A1(n10485), .A2(n10491), .ZN(n19568) );
  OR2_X1 U11380 ( .A1(n14704), .A2(n10981), .ZN(n10957) );
  OR2_X1 U11381 ( .A1(n18882), .A2(n18881), .ZN(n18884) );
  NAND2_X2 U11382 ( .A1(n20040), .A2(n20209), .ZN(n14194) );
  CLKBUF_X3 U11383 ( .A(n12087), .Z(n9753) );
  INV_X1 U11384 ( .A(n10498), .ZN(n10492) );
  NOR2_X1 U11385 ( .A1(n14190), .A2(n14107), .ZN(n14109) );
  NAND2_X1 U11386 ( .A1(n12684), .A2(n12683), .ZN(n12836) );
  OR2_X1 U11387 ( .A1(n15893), .A2(n14188), .ZN(n14190) );
  AND2_X1 U11388 ( .A1(n10467), .A2(n10743), .ZN(n10745) );
  NAND2_X1 U11389 ( .A1(n19155), .A2(n12888), .ZN(n12684) );
  AND2_X2 U11390 ( .A1(n10480), .A2(n10478), .ZN(n19155) );
  XNOR2_X1 U11391 ( .A(n10856), .B(n10855), .ZN(n12051) );
  NAND2_X1 U11392 ( .A1(n11326), .A2(n10135), .ZN(n12437) );
  NAND2_X1 U11394 ( .A1(n10128), .A2(n11327), .ZN(n11326) );
  OR2_X1 U11395 ( .A1(n11245), .A2(n11246), .ZN(n11225) );
  NAND2_X1 U11396 ( .A1(n11231), .A2(n11230), .ZN(n20322) );
  AND2_X1 U11397 ( .A1(n10433), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10457) );
  OAI22_X1 U11398 ( .A1(n10433), .A2(n10432), .B1(n10733), .B2(n10431), .ZN(
        n10437) );
  AND3_X1 U11399 ( .A1(n10440), .A2(n10439), .A3(n10438), .ZN(n10470) );
  AND2_X1 U11400 ( .A1(n10073), .A2(n11935), .ZN(n10072) );
  NOR2_X1 U11401 ( .A1(n12867), .A2(n12115), .ZN(n12120) );
  AOI22_X1 U11402 ( .A1(n13859), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n12588), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10404) );
  INV_X2 U11403 ( .A(n19073), .ZN(n12748) );
  NOR2_X1 U11404 ( .A1(n12865), .A2(n12866), .ZN(n12867) );
  AOI22_X1 U11405 ( .A1(n11144), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n11210), 
        .B2(n11154), .ZN(n11145) );
  NOR2_X2 U11406 ( .A1(n10883), .A2(n10866), .ZN(n10891) );
  AND2_X1 U11407 ( .A1(n10423), .A2(n10422), .ZN(n10425) );
  NAND2_X1 U11408 ( .A1(n10885), .A2(n10884), .ZN(n10883) );
  INV_X1 U11409 ( .A(n12269), .ZN(n16319) );
  NOR2_X2 U11410 ( .A1(n17342), .A2(n15748), .ZN(n17761) );
  AND2_X1 U11411 ( .A1(n12688), .A2(n10188), .ZN(n12114) );
  AND2_X1 U11412 ( .A1(n10874), .A2(n10869), .ZN(n10885) );
  INV_X1 U11413 ( .A(n10406), .ZN(n12269) );
  AND2_X1 U11414 ( .A1(n12892), .A2(n12891), .ZN(n12893) );
  OR2_X2 U11415 ( .A1(n17414), .A2(n18678), .ZN(n17482) );
  NAND2_X1 U11416 ( .A1(n13357), .A2(n10045), .ZN(n10047) );
  NOR2_X1 U11417 ( .A1(n10430), .A2(n10394), .ZN(n12848) );
  NAND2_X1 U11418 ( .A1(n12364), .A2(n12344), .ZN(n12377) );
  NOR2_X1 U11419 ( .A1(n10875), .A2(n10876), .ZN(n10874) );
  INV_X1 U11420 ( .A(n11152), .ZN(n12626) );
  NAND2_X2 U11421 ( .A1(n10400), .A2(n16300), .ZN(n16302) );
  AND2_X1 U11422 ( .A1(n10046), .A2(n13180), .ZN(n10045) );
  AND2_X1 U11423 ( .A1(n10410), .A2(n12340), .ZN(n10418) );
  CLKBUF_X1 U11424 ( .A(n12340), .Z(n12661) );
  AND2_X1 U11425 ( .A1(n12295), .A2(n19250), .ZN(n10393) );
  AND3_X2 U11426 ( .A1(n12686), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13832), 
        .ZN(n13757) );
  AND3_X1 U11427 ( .A1(n10269), .A2(n10386), .A3(n19234), .ZN(n10400) );
  NAND4_X1 U11428 ( .A1(n10035), .A2(n11130), .A3(n10033), .A4(n9785), .ZN(
        n11152) );
  INV_X1 U11429 ( .A(n10385), .ZN(n12294) );
  AND3_X1 U11430 ( .A1(n16316), .A2(n10860), .A3(n19250), .ZN(n12094) );
  NOR2_X1 U11431 ( .A1(n10413), .A2(n10385), .ZN(n10333) );
  NAND2_X1 U11432 ( .A1(n11155), .A2(n20209), .ZN(n12970) );
  INV_X1 U11433 ( .A(n16316), .ZN(n9740) );
  INV_X2 U11434 ( .A(n16454), .ZN(n16451) );
  NOR2_X1 U11435 ( .A1(n11155), .A2(n11307), .ZN(n11500) );
  INV_X2 U11436 ( .A(n20166), .ZN(n9731) );
  OR2_X1 U11437 ( .A1(n10571), .A2(n10572), .ZN(n10723) );
  INV_X1 U11438 ( .A(n19212), .ZN(n10409) );
  NOR2_X2 U11439 ( .A1(n15395), .A2(n15394), .ZN(n18835) );
  INV_X1 U11440 ( .A(n10399), .ZN(n12686) );
  NAND2_X1 U11441 ( .A1(n10307), .A2(n10306), .ZN(n10385) );
  INV_X2 U11442 ( .A(U212), .ZN(n16449) );
  NAND2_X2 U11443 ( .A1(n9948), .A2(n9946), .ZN(n19212) );
  NAND2_X1 U11444 ( .A1(n10345), .A2(n10344), .ZN(n10865) );
  NAND2_X1 U11445 ( .A1(n10332), .A2(n10331), .ZN(n10414) );
  NAND2_X1 U11446 ( .A1(n9944), .A2(n9942), .ZN(n10411) );
  AND4_X1 U11447 ( .A1(n11079), .A2(n11078), .A3(n11077), .A4(n11076), .ZN(
        n11080) );
  AND4_X1 U11448 ( .A1(n11095), .A2(n11094), .A3(n11093), .A4(n11092), .ZN(
        n11100) );
  AND2_X1 U11449 ( .A1(n10295), .A2(n10294), .ZN(n10299) );
  NAND2_X2 U11450 ( .A1(n18779), .A2(n18714), .ZN(n18760) );
  AND2_X2 U11451 ( .A1(n13879), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10574) );
  BUF_X2 U11452 ( .A(n11799), .Z(n9752) );
  AND2_X1 U11453 ( .A1(n11037), .A2(n11036), .ZN(n11042) );
  AND2_X1 U11455 ( .A1(n10314), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10318) );
  AND3_X1 U11456 ( .A1(n10309), .A2(n10308), .A3(n12956), .ZN(n10313) );
  INV_X1 U11457 ( .A(n11703), .ZN(n11176) );
  INV_X2 U11458 ( .A(n13660), .ZN(n13879) );
  AND2_X2 U11459 ( .A1(n13878), .A2(n12956), .ZN(n13652) );
  INV_X2 U11460 ( .A(n16487), .ZN(U215) );
  AND2_X2 U11461 ( .A1(n10506), .A2(n12956), .ZN(n12162) );
  BUF_X2 U11462 ( .A(n15533), .Z(n17171) );
  NAND2_X2 U11463 ( .A1(n19944), .A2(n19842), .ZN(n19889) );
  NAND2_X1 U11465 ( .A1(n11044), .A2(n11039), .ZN(n9779) );
  BUF_X4 U11466 ( .A(n15396), .Z(n9735) );
  OR2_X2 U11467 ( .A1(n12416), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n19990) );
  BUF_X2 U11468 ( .A(n10513), .Z(n13878) );
  CLKBUF_X1 U11469 ( .A(n10508), .Z(n13660) );
  INV_X4 U11470 ( .A(n18169), .ZN(n9736) );
  AND2_X2 U11471 ( .A1(n10278), .A2(n10444), .ZN(n10506) );
  INV_X2 U11472 ( .A(n10508), .ZN(n10507) );
  NAND2_X1 U11473 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18803), .ZN(
        n15386) );
  NAND3_X1 U11474 ( .A1(n10114), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10508) );
  NOR2_X1 U11475 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11040) );
  INV_X4 U11476 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10444) );
  AND2_X1 U11477 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11028) );
  NAND2_X1 U11478 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16885) );
  INV_X1 U11479 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18818) );
  INV_X2 U11480 ( .A(n13225), .ZN(n9911) );
  AOI21_X2 U11481 ( .B1(n12833), .B2(n12888), .A(n12832), .ZN(n12863) );
  AND2_X1 U11482 ( .A1(n12104), .A2(n16316), .ZN(n12343) );
  OAI21_X1 U11483 ( .B1(n9725), .B2(n15846), .A(n18830), .ZN(n17368) );
  NAND2_X2 U11484 ( .A1(n14780), .A2(n14781), .ZN(n14776) );
  NOR2_X4 U11485 ( .A1(n13575), .A2(n10251), .ZN(n14780) );
  NAND2_X2 U11486 ( .A1(n11218), .A2(n11145), .ZN(n11219) );
  OR2_X1 U11487 ( .A1(n13735), .A2(n13734), .ZN(n13736) );
  OAI21_X1 U11488 ( .B1(n12436), .B2(n11317), .A(n11318), .ZN(n11215) );
  NOR2_X2 U11489 ( .A1(n15845), .A2(n9863), .ZN(n17212) );
  AND2_X1 U11490 ( .A1(n10278), .A2(n10444), .ZN(n9737) );
  AND2_X2 U11491 ( .A1(n10278), .A2(n10444), .ZN(n9738) );
  OR2_X1 U11492 ( .A1(n12833), .A2(n19155), .ZN(n10494) );
  AOI21_X2 U11493 ( .B1(n14999), .B2(n15000), .A(n14951), .ZN(n14991) );
  NOR2_X2 U11494 ( .A1(n14077), .A2(n10171), .ZN(n14047) );
  NAND2_X2 U11495 ( .A1(n10043), .A2(n11143), .ZN(n12388) );
  NOR2_X2 U11496 ( .A1(n12070), .A2(n16174), .ZN(n12071) );
  OR2_X2 U11497 ( .A1(n11114), .A2(n11113), .ZN(n20166) );
  OAI22_X2 U11498 ( .A1(n12051), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n16324), 
        .B2(n10698), .ZN(n12089) );
  INV_X4 U11499 ( .A(n11232), .ZN(n11120) );
  NAND2_X1 U11500 ( .A1(n13147), .A2(n12774), .ZN(n11232) );
  AOI21_X2 U11501 ( .B1(n12864), .B2(n12863), .A(n12837), .ZN(n12896) );
  NOR2_X2 U11502 ( .A1(n13214), .A2(n13213), .ZN(n13212) );
  NAND2_X1 U11503 ( .A1(n20219), .A2(n11250), .ZN(n13170) );
  NOR2_X2 U11504 ( .A1(n12055), .A2(n9999), .ZN(n12053) );
  NOR2_X2 U11505 ( .A1(n13475), .A2(n11415), .ZN(n13510) );
  OAI21_X1 U11506 ( .B1(n15778), .B2(n9993), .A(n9992), .ZN(n12551) );
  XNOR2_X2 U11507 ( .A(n12446), .B(n20156), .ZN(n13126) );
  NAND2_X2 U11508 ( .A1(n13057), .A2(n12445), .ZN(n12446) );
  NOR2_X2 U11509 ( .A1(n14030), .A2(n10163), .ZN(n13976) );
  INV_X1 U11510 ( .A(n11138), .ZN(n9743) );
  INV_X1 U11511 ( .A(n9743), .ZN(n9744) );
  AND2_X1 U11512 ( .A1(n11046), .A2(n13150), .ZN(n9746) );
  AND2_X1 U11513 ( .A1(n11046), .A2(n13150), .ZN(n11638) );
  NOR2_X4 U11514 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11044) );
  AND2_X1 U11515 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11045) );
  NAND2_X1 U11516 ( .A1(n20285), .A2(n11163), .ZN(n11250) );
  NAND2_X2 U11517 ( .A1(n13952), .A2(n13953), .ZN(n13939) );
  NOR2_X4 U11518 ( .A1(n13966), .A2(n13967), .ZN(n13952) );
  INV_X2 U11519 ( .A(n11827), .ZN(n9747) );
  INV_X1 U11520 ( .A(n11813), .ZN(n9748) );
  NAND2_X1 U11523 ( .A1(n13150), .A2(n11040), .ZN(n11813) );
  INV_X1 U11524 ( .A(n9779), .ZN(n11799) );
  INV_X1 U11525 ( .A(n12089), .ZN(n12087) );
  AND2_X4 U11526 ( .A1(n12780), .A2(n14646), .ZN(n11194) );
  INV_X1 U11527 ( .A(n10645), .ZN(n9919) );
  INV_X1 U11528 ( .A(n10660), .ZN(n10640) );
  AND2_X1 U11529 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10511) );
  AND2_X1 U11530 ( .A1(n11251), .A2(n9888), .ZN(n9884) );
  NOR2_X1 U11531 ( .A1(n9890), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9888) );
  INV_X1 U11532 ( .A(n11266), .ZN(n9890) );
  AND2_X1 U11533 ( .A1(n12774), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10031) );
  NAND2_X1 U11534 ( .A1(n13000), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11263) );
  NOR2_X1 U11535 ( .A1(n20209), .A2(n11307), .ZN(n11333) );
  INV_X1 U11536 ( .A(n11728), .ZN(n11189) );
  NAND2_X1 U11537 ( .A1(n11138), .A2(n20189), .ZN(n11103) );
  NAND2_X1 U11538 ( .A1(n11265), .A2(n11263), .ZN(n11895) );
  AND3_X1 U11539 ( .A1(n20166), .A2(n11204), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11898) );
  NOR2_X1 U11540 ( .A1(n10185), .A2(n10184), .ZN(n10183) );
  INV_X1 U11541 ( .A(n14091), .ZN(n10184) );
  NAND2_X1 U11542 ( .A1(n10156), .A2(n10179), .ZN(n10155) );
  INV_X1 U11543 ( .A(n11338), .ZN(n11845) );
  NOR3_X1 U11544 ( .A1(n14411), .A2(n14476), .A3(n10053), .ZN(n10052) );
  NAND2_X1 U11545 ( .A1(n10891), .A2(n10105), .ZN(n10913) );
  AND2_X1 U11546 ( .A1(n9786), .A2(n10906), .ZN(n10105) );
  INV_X1 U11547 ( .A(n13757), .ZN(n13786) );
  NAND2_X1 U11548 ( .A1(n13736), .A2(n14745), .ZN(n13760) );
  NOR2_X1 U11549 ( .A1(n10406), .A2(n9740), .ZN(n10408) );
  NOR2_X1 U11550 ( .A1(n13347), .A2(n13346), .ZN(n10082) );
  AOI21_X1 U11551 ( .B1(n10690), .B2(n16245), .A(n10148), .ZN(n10147) );
  INV_X1 U11552 ( .A(n16204), .ZN(n10148) );
  INV_X1 U11553 ( .A(n10657), .ZN(n9938) );
  AND2_X1 U11554 ( .A1(n10160), .A2(n16181), .ZN(n10159) );
  OR2_X1 U11555 ( .A1(n10636), .A2(n10635), .ZN(n12134) );
  NAND2_X1 U11556 ( .A1(n15345), .A2(n10663), .ZN(n10689) );
  OAI21_X1 U11557 ( .B1(n13257), .B2(n13256), .A(n9758), .ZN(n10145) );
  INV_X1 U11558 ( .A(n10145), .ZN(n10143) );
  AND2_X1 U11559 ( .A1(n10573), .A2(n10526), .ZN(n10136) );
  INV_X1 U11560 ( .A(n10723), .ZN(n12118) );
  NAND2_X1 U11561 ( .A1(n17376), .A2(n15582), .ZN(n15598) );
  INV_X2 U11562 ( .A(n11689), .ZN(n11847) );
  AND2_X1 U11563 ( .A1(n11307), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11846) );
  OR2_X1 U11564 ( .A1(n12979), .A2(n19949), .ZN(n12805) );
  AOI21_X1 U11565 ( .B1(n14308), .B2(n14411), .A(n10050), .ZN(n10048) );
  INV_X1 U11566 ( .A(n10051), .ZN(n10050) );
  AOI21_X1 U11567 ( .B1(n14411), .B2(n14309), .A(n10055), .ZN(n10051) );
  NAND2_X1 U11568 ( .A1(n12983), .A2(n12982), .ZN(n13005) );
  NAND2_X1 U11569 ( .A1(n16096), .A2(n16081), .ZN(n16080) );
  INV_X1 U11570 ( .A(n14813), .ZN(n12268) );
  NAND2_X1 U11571 ( .A1(n12268), .A2(n12267), .ZN(n15052) );
  AND2_X1 U11572 ( .A1(n12664), .A2(n12663), .ZN(n12679) );
  NAND2_X1 U11573 ( .A1(n9962), .A2(n11010), .ZN(n14899) );
  AND2_X1 U11574 ( .A1(n12337), .A2(n19815), .ZN(n12382) );
  OR2_X1 U11575 ( .A1(n16815), .A2(n17537), .ZN(n10004) );
  AND2_X1 U11576 ( .A1(n14416), .A2(n12420), .ZN(n15932) );
  INV_X2 U11577 ( .A(n14416), .ZN(n20111) );
  NAND2_X1 U11578 ( .A1(n12291), .A2(n10732), .ZN(n12587) );
  OR2_X1 U11579 ( .A1(n19053), .A2(n19250), .ZN(n16132) );
  NAND2_X1 U11580 ( .A1(n10396), .A2(n10395), .ZN(n10423) );
  NAND2_X1 U11581 ( .A1(n10394), .A2(n10384), .ZN(n10395) );
  AND2_X1 U11582 ( .A1(n11886), .A2(n11885), .ZN(n11888) );
  NAND2_X1 U11583 ( .A1(n9731), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11265) );
  NOR2_X1 U11584 ( .A1(n10058), .A2(n11293), .ZN(n10057) );
  INV_X1 U11585 ( .A(n11355), .ZN(n10058) );
  AND2_X1 U11586 ( .A1(n11188), .A2(n11187), .ZN(n11209) );
  NAND2_X1 U11587 ( .A1(n9886), .A2(n9889), .ZN(n9885) );
  AOI21_X1 U11588 ( .B1(n9884), .B2(n11252), .A(n9883), .ZN(n9882) );
  NAND2_X1 U11589 ( .A1(n9881), .A2(n9889), .ZN(n9880) );
  INV_X1 U11590 ( .A(n13357), .ZN(n12763) );
  AND2_X1 U11591 ( .A1(n12625), .A2(n12624), .ZN(n12756) );
  INV_X1 U11592 ( .A(n10692), .ZN(n9955) );
  AND4_X1 U11593 ( .A1(n10490), .A2(n10489), .A3(n10488), .A4(n10487), .ZN(
        n10505) );
  NAND2_X1 U11594 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10275) );
  NAND2_X1 U11595 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18793), .ZN(
        n15384) );
  NAND2_X1 U11596 ( .A1(n18818), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15387) );
  NOR2_X1 U11597 ( .A1(n17350), .A2(n15733), .ZN(n15731) );
  INV_X1 U11598 ( .A(n15426), .ZN(n9907) );
  INV_X1 U11599 ( .A(n15434), .ZN(n9862) );
  NAND2_X1 U11600 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n9861) );
  NOR2_X1 U11601 ( .A1(n14086), .A2(n10064), .ZN(n10063) );
  INV_X1 U11602 ( .A(n14094), .ZN(n10064) );
  NAND2_X1 U11603 ( .A1(n10167), .A2(n10166), .ZN(n10165) );
  INV_X1 U11604 ( .A(n14006), .ZN(n10166) );
  INV_X1 U11605 ( .A(n10168), .ZN(n10167) );
  NAND2_X1 U11606 ( .A1(n14016), .A2(n10169), .ZN(n10168) );
  INV_X1 U11607 ( .A(n14032), .ZN(n10169) );
  NAND2_X1 U11608 ( .A1(n10173), .A2(n10172), .ZN(n10171) );
  INV_X1 U11609 ( .A(n14049), .ZN(n10172) );
  CLKBUF_X1 U11610 ( .A(n11338), .Z(n11914) );
  NAND2_X1 U11611 ( .A1(n14003), .A2(n14019), .ZN(n10068) );
  NAND2_X1 U11612 ( .A1(n12512), .A2(n10127), .ZN(n10124) );
  INV_X1 U11613 ( .A(n14410), .ZN(n10126) );
  NOR2_X1 U11614 ( .A1(n10079), .A2(n10078), .ZN(n10077) );
  INV_X1 U11615 ( .A(n13536), .ZN(n10078) );
  INV_X1 U11616 ( .A(n13499), .ZN(n10076) );
  NAND2_X1 U11617 ( .A1(n10080), .A2(n13517), .ZN(n10079) );
  INV_X1 U11618 ( .A(n13500), .ZN(n10080) );
  AND2_X1 U11619 ( .A1(n15953), .A2(n12482), .ZN(n9865) );
  NAND2_X1 U11620 ( .A1(n12482), .A2(n10119), .ZN(n10118) );
  INV_X1 U11621 ( .A(n12472), .ZN(n10119) );
  INV_X1 U11622 ( .A(n13234), .ZN(n10073) );
  INV_X1 U11623 ( .A(n13126), .ZN(n9855) );
  INV_X1 U11624 ( .A(n12447), .ZN(n9871) );
  OR2_X1 U11625 ( .A1(n11242), .A2(n11241), .ZN(n12465) );
  NOR2_X1 U11626 ( .A1(n10134), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10133) );
  INV_X1 U11627 ( .A(n11150), .ZN(n10134) );
  NAND2_X1 U11628 ( .A1(n11268), .A2(n11312), .ZN(n11356) );
  AND2_X1 U11629 ( .A1(n12756), .A2(n12978), .ZN(n12786) );
  AND2_X1 U11630 ( .A1(n11115), .A2(n12626), .ZN(n10043) );
  INV_X1 U11631 ( .A(n20250), .ZN(n20287) );
  AND2_X1 U11632 ( .A1(n11228), .A2(n20707), .ZN(n20443) );
  INV_X1 U11633 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11122) );
  NOR2_X1 U11634 ( .A1(n11128), .A2(n10036), .ZN(n10035) );
  NAND2_X1 U11635 ( .A1(n20773), .A2(n20165), .ZN(n20327) );
  OR2_X1 U11636 ( .A1(n10986), .A2(n10985), .ZN(n10994) );
  INV_X1 U11637 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n10099) );
  AOI21_X1 U11638 ( .B1(n12885), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12884), .ZN(n12891) );
  NAND2_X1 U11639 ( .A1(n9822), .A2(n14750), .ZN(n9915) );
  NAND2_X1 U11640 ( .A1(n10093), .A2(n14693), .ZN(n10092) );
  INV_X1 U11641 ( .A(n14797), .ZN(n10093) );
  NOR2_X1 U11642 ( .A1(n9987), .A2(n9986), .ZN(n9985) );
  NAND2_X1 U11643 ( .A1(n10685), .A2(n9924), .ZN(n10691) );
  INV_X1 U11644 ( .A(n10664), .ZN(n10685) );
  AND2_X1 U11645 ( .A1(n10097), .A2(n13047), .ZN(n10096) );
  NOR2_X1 U11646 ( .A1(n10098), .A2(n13032), .ZN(n10097) );
  INV_X1 U11647 ( .A(n13043), .ZN(n10098) );
  AND4_X1 U11648 ( .A1(n10668), .A2(n10667), .A3(n10666), .A4(n10665), .ZN(
        n10684) );
  INV_X1 U11649 ( .A(n12043), .ZN(n10088) );
  INV_X1 U11650 ( .A(n14836), .ZN(n10221) );
  OR2_X1 U11651 ( .A1(n13037), .A2(n10218), .ZN(n10217) );
  INV_X1 U11652 ( .A(n13061), .ZN(n10218) );
  OR2_X1 U11653 ( .A1(n10147), .A2(n9955), .ZN(n9953) );
  NAND2_X1 U11654 ( .A1(n9952), .A2(n10690), .ZN(n9954) );
  NOR2_X1 U11655 ( .A1(n15040), .A2(n9955), .ZN(n9952) );
  NAND2_X1 U11656 ( .A1(n10639), .A2(n10638), .ZN(n10660) );
  OR2_X1 U11657 ( .A1(n10626), .A2(n10625), .ZN(n10639) );
  NOR2_X1 U11658 ( .A1(n10552), .A2(n10551), .ZN(n16267) );
  NAND2_X1 U11659 ( .A1(n10190), .A2(n10189), .ZN(n12124) );
  NAND3_X1 U11660 ( .A1(n10388), .A2(n16300), .A3(n10387), .ZN(n12347) );
  AND2_X1 U11661 ( .A1(n12833), .A2(n19035), .ZN(n10498) );
  INV_X1 U11662 ( .A(n17487), .ZN(n10008) );
  OR2_X1 U11663 ( .A1(n15386), .A2(n15387), .ZN(n15669) );
  OR2_X1 U11664 ( .A1(n16884), .A2(n15388), .ZN(n9776) );
  NAND2_X1 U11665 ( .A1(n18811), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15385) );
  NAND2_X1 U11666 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17567), .ZN(
        n17532) );
  NOR2_X1 U11667 ( .A1(n17618), .A2(n10014), .ZN(n10013) );
  INV_X1 U11668 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10014) );
  NOR2_X1 U11669 ( .A1(n15827), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16341) );
  OR2_X1 U11670 ( .A1(n16388), .A2(n15828), .ZN(n16343) );
  INV_X1 U11671 ( .A(n17651), .ZN(n15768) );
  NAND2_X1 U11672 ( .A1(n15731), .A2(n17345), .ZN(n15748) );
  NOR2_X1 U11673 ( .A1(n10238), .A2(n10237), .ZN(n10235) );
  NAND2_X1 U11674 ( .A1(n10239), .A2(n21143), .ZN(n10237) );
  AND2_X1 U11675 ( .A1(n15574), .A2(n17263), .ZN(n15601) );
  NAND2_X1 U11676 ( .A1(n9931), .A2(n15742), .ZN(n15745) );
  NAND2_X1 U11677 ( .A1(n11931), .A2(n11930), .ZN(n13187) );
  NAND2_X1 U11678 ( .A1(n13357), .A2(n10044), .ZN(n12766) );
  AND2_X1 U11679 ( .A1(n13180), .A2(n13181), .ZN(n10044) );
  OR2_X1 U11680 ( .A1(n11695), .A2(n11694), .ZN(n13991) );
  OR2_X1 U11681 ( .A1(n11631), .A2(n11630), .ZN(n11636) );
  INV_X1 U11682 ( .A(n13511), .ZN(n11415) );
  INV_X1 U11683 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11379) );
  NAND2_X1 U11684 ( .A1(n14308), .A2(n12521), .ZN(n9857) );
  OAI21_X1 U11685 ( .B1(n14308), .B2(n14309), .A(n14411), .ZN(n14333) );
  AND2_X1 U11686 ( .A1(n14614), .A2(n14457), .ZN(n14604) );
  OR2_X1 U11687 ( .A1(n20142), .A2(n14618), .ZN(n16017) );
  NAND2_X1 U11688 ( .A1(n11252), .A2(n11251), .ZN(n13145) );
  INV_X1 U11689 ( .A(n19949), .ZN(n12982) );
  INV_X1 U11690 ( .A(n20535), .ZN(n20419) );
  AND2_X1 U11691 ( .A1(n20563), .A2(n20213), .ZN(n20497) );
  INV_X1 U11692 ( .A(n20536), .ZN(n20488) );
  OR2_X1 U11693 ( .A1(n20639), .A2(n20610), .ZN(n20650) );
  NAND2_X1 U11694 ( .A1(n13405), .A2(n11344), .ZN(n20639) );
  AND2_X1 U11695 ( .A1(n11907), .A2(n11906), .ZN(n12979) );
  NAND2_X1 U11696 ( .A1(n10104), .A2(n10103), .ZN(n10862) );
  NAND2_X1 U11697 ( .A1(n12338), .A2(n12317), .ZN(n10103) );
  OR2_X1 U11698 ( .A1(n10723), .A2(n12338), .ZN(n10104) );
  XNOR2_X1 U11699 ( .A(n11012), .B(n11011), .ZN(n16066) );
  NOR2_X1 U11700 ( .A1(n16080), .A2(n11001), .ZN(n11012) );
  INV_X1 U11701 ( .A(n14930), .ZN(n9989) );
  NAND2_X1 U11702 ( .A1(n10999), .A2(n11018), .ZN(n16096) );
  NOR2_X1 U11703 ( .A1(n16112), .A2(n9753), .ZN(n14676) );
  NAND2_X1 U11704 ( .A1(n9990), .A2(n9989), .ZN(n9991) );
  INV_X1 U11705 ( .A(n14676), .ZN(n9990) );
  NOR2_X1 U11706 ( .A1(n12551), .A2(n9753), .ZN(n16113) );
  OR2_X1 U11707 ( .A1(n15778), .A2(n15779), .ZN(n9994) );
  NOR2_X1 U11708 ( .A1(n9753), .A2(n12563), .ZN(n15778) );
  NOR2_X1 U11709 ( .A1(n16291), .A2(n16333), .ZN(n12578) );
  NAND2_X1 U11710 ( .A1(n13351), .A2(n9820), .ZN(n10257) );
  INV_X1 U11711 ( .A(n10257), .ZN(n10256) );
  NOR2_X1 U11712 ( .A1(n13224), .A2(n9913), .ZN(n9912) );
  INV_X1 U11713 ( .A(n13227), .ZN(n13224) );
  NOR2_X1 U11714 ( .A1(n13030), .A2(n13039), .ZN(n13031) );
  AND2_X1 U11715 ( .A1(n12901), .A2(n12900), .ZN(n12902) );
  NAND2_X1 U11716 ( .A1(n16296), .A2(n16293), .ZN(n12849) );
  NAND2_X1 U11717 ( .A1(n10252), .A2(n13606), .ZN(n10251) );
  INV_X1 U11718 ( .A(n10253), .ZN(n10252) );
  NAND2_X1 U11719 ( .A1(n13446), .A2(n10204), .ZN(n10203) );
  INV_X1 U11720 ( .A(n13137), .ZN(n10204) );
  NAND2_X1 U11721 ( .A1(n10000), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9999) );
  NOR2_X1 U11722 ( .A1(n14668), .A2(n10002), .ZN(n10000) );
  CLKBUF_X1 U11723 ( .A(n12055), .Z(n12056) );
  CLKBUF_X1 U11724 ( .A(n12060), .Z(n12061) );
  AND2_X1 U11725 ( .A1(n10810), .A2(n10809), .ZN(n12567) );
  AND2_X1 U11726 ( .A1(n10777), .A2(n10776), .ZN(n13346) );
  INV_X1 U11727 ( .A(n10082), .ZN(n13391) );
  AND2_X1 U11728 ( .A1(n10764), .A2(n10763), .ZN(n13116) );
  OAI21_X1 U11729 ( .B1(n10149), .B2(n15040), .A(n10147), .ZN(n16203) );
  NAND2_X1 U11730 ( .A1(n10140), .A2(n13445), .ZN(n10139) );
  INV_X1 U11731 ( .A(n10659), .ZN(n10859) );
  OR3_X1 U11732 ( .A1(n14689), .A2(n10981), .A3(n21137), .ZN(n14923) );
  NAND2_X1 U11733 ( .A1(n10993), .A2(n15124), .ZN(n9923) );
  INV_X1 U11734 ( .A(n9922), .ZN(n9921) );
  AOI21_X1 U11735 ( .B1(n9975), .B2(n9781), .A(n9974), .ZN(n9973) );
  NAND2_X1 U11736 ( .A1(n13207), .A2(n13220), .ZN(n13219) );
  NAND2_X1 U11737 ( .A1(n15275), .A2(n10924), .ZN(n14943) );
  OR2_X1 U11738 ( .A1(n10217), .A2(n13088), .ZN(n10216) );
  OR2_X1 U11739 ( .A1(n12940), .A2(n10217), .ZN(n13087) );
  NAND2_X1 U11740 ( .A1(n10910), .A2(n16177), .ZN(n16181) );
  AND2_X1 U11741 ( .A1(n10904), .A2(n10161), .ZN(n10160) );
  INV_X1 U11742 ( .A(n15322), .ZN(n10161) );
  AND2_X1 U11743 ( .A1(n19186), .A2(n19192), .ZN(n15307) );
  NAND2_X1 U11744 ( .A1(n12134), .A2(n12225), .ZN(n10207) );
  NAND2_X1 U11745 ( .A1(n10192), .A2(n10196), .ZN(n12923) );
  AOI21_X1 U11746 ( .B1(n10198), .B2(n10205), .A(n10197), .ZN(n10196) );
  AOI21_X1 U11747 ( .B1(n10203), .B2(n10207), .A(n12692), .ZN(n10200) );
  NAND2_X1 U11748 ( .A1(n16302), .A2(n16319), .ZN(n16292) );
  INV_X1 U11749 ( .A(n12954), .ZN(n16295) );
  NAND2_X1 U11750 ( .A1(n19266), .A2(n19928), .ZN(n19413) );
  NAND2_X1 U11751 ( .A1(n19266), .A2(n19265), .ZN(n19450) );
  NAND2_X1 U11752 ( .A1(n19902), .A2(n19265), .ZN(n19633) );
  NAND2_X1 U11753 ( .A1(n16815), .A2(n10011), .ZN(n10010) );
  NAND2_X1 U11754 ( .A1(n16852), .A2(n17507), .ZN(n10011) );
  AND2_X1 U11755 ( .A1(n10003), .A2(n9837), .ZN(n16586) );
  AOI211_X1 U11756 ( .C1(n15582), .C2(n16515), .A(n18707), .B(n18654), .ZN(
        n15847) );
  NOR2_X1 U11757 ( .A1(n17849), .A2(n17498), .ZN(n16528) );
  OR2_X1 U11758 ( .A1(n17598), .A2(n17505), .ZN(n15828) );
  NAND2_X1 U11759 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17518), .ZN(
        n17498) );
  NOR2_X1 U11760 ( .A1(n17787), .A2(n10023), .ZN(n10021) );
  NAND2_X1 U11761 ( .A1(n10024), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10023) );
  INV_X1 U11762 ( .A(n17703), .ZN(n10024) );
  AOI21_X1 U11763 ( .B1(n17563), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n18566), .ZN(n17702) );
  NOR2_X1 U11764 ( .A1(n16348), .A2(n10228), .ZN(n10227) );
  NAND2_X1 U11765 ( .A1(n16344), .A2(n10229), .ZN(n10228) );
  OR2_X1 U11766 ( .A1(n17761), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10229) );
  NAND2_X1 U11767 ( .A1(n16343), .A2(n10230), .ZN(n15829) );
  NAND2_X1 U11768 ( .A1(n16341), .A2(n17598), .ZN(n10230) );
  NAND2_X1 U11769 ( .A1(n15829), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16342) );
  AND2_X1 U11770 ( .A1(n10232), .A2(n10231), .ZN(n17646) );
  NAND2_X1 U11771 ( .A1(n17651), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10231) );
  NOR2_X1 U11772 ( .A1(n10234), .A2(n17650), .ZN(n10232) );
  AND2_X1 U11773 ( .A1(n17761), .A2(n17992), .ZN(n10234) );
  NOR2_X1 U11774 ( .A1(n17722), .A2(n21143), .ZN(n18029) );
  NAND2_X1 U11775 ( .A1(n15727), .A2(n17762), .ZN(n18027) );
  INV_X1 U11776 ( .A(n18027), .ZN(n17974) );
  INV_X1 U11777 ( .A(n18029), .ZN(n17973) );
  INV_X1 U11778 ( .A(n15751), .ZN(n10238) );
  NOR2_X1 U11779 ( .A1(n9936), .A2(n21143), .ZN(n17759) );
  INV_X1 U11780 ( .A(n15761), .ZN(n9936) );
  XNOR2_X1 U11781 ( .A(n15749), .B(n9935), .ZN(n17773) );
  INV_X1 U11782 ( .A(n15750), .ZN(n9935) );
  AOI21_X1 U11783 ( .B1(n15562), .B2(n18835), .A(n15598), .ZN(n15604) );
  NOR3_X1 U11784 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18719), .A3(n18698), 
        .ZN(n16518) );
  OR2_X1 U11785 ( .A1(n15820), .A2(n20773), .ZN(n19949) );
  XNOR2_X1 U11786 ( .A(n10061), .B(n13910), .ZN(n14477) );
  INV_X1 U11787 ( .A(n13911), .ZN(n10061) );
  AND2_X1 U11788 ( .A1(n15908), .A2(n13068), .ZN(n14273) );
  INV_X1 U11789 ( .A(n15908), .ZN(n14289) );
  XNOR2_X1 U11790 ( .A(n11920), .B(n11919), .ZN(n13364) );
  XNOR2_X1 U11791 ( .A(n13912), .B(n11848), .ZN(n12423) );
  NAND2_X1 U11792 ( .A1(n19955), .A2(n12417), .ZN(n14416) );
  OAI211_X1 U11793 ( .C1(n14291), .C2(n9877), .A(n9873), .B(n9872), .ZN(n14451) );
  NAND2_X1 U11794 ( .A1(n9879), .A2(n10115), .ZN(n9877) );
  NAND2_X1 U11795 ( .A1(n9875), .A2(n9874), .ZN(n9873) );
  NAND2_X1 U11796 ( .A1(n14291), .A2(n9808), .ZN(n9872) );
  INV_X1 U11797 ( .A(n14477), .ZN(n10060) );
  INV_X1 U11798 ( .A(n16017), .ZN(n15969) );
  NAND2_X1 U11799 ( .A1(n20420), .A2(n20419), .ZN(n20442) );
  NOR2_X1 U11800 ( .A1(n10721), .A2(n10729), .ZN(n19937) );
  OR2_X1 U11801 ( .A1(n12237), .A2(n12236), .ZN(n13463) );
  NAND2_X1 U11802 ( .A1(n10209), .A2(n9824), .ZN(n10208) );
  NAND2_X1 U11803 ( .A1(n14883), .A2(n13903), .ZN(n10209) );
  OR2_X1 U11804 ( .A1(n12268), .A2(n12267), .ZN(n10211) );
  NAND2_X1 U11805 ( .A1(n12680), .A2(n19815), .ZN(n19053) );
  OR2_X1 U11806 ( .A1(n19053), .A2(n12104), .ZN(n16133) );
  INV_X1 U11807 ( .A(n10858), .ZN(n10085) );
  XNOR2_X1 U11808 ( .A(n12281), .B(n10851), .ZN(n16057) );
  NOR2_X1 U11809 ( .A1(n9957), .A2(n15218), .ZN(n9956) );
  INV_X1 U11810 ( .A(n9958), .ZN(n9957) );
  OR2_X1 U11811 ( .A1(n12587), .A2(n9740), .ZN(n19159) );
  AND2_X1 U11812 ( .A1(n16225), .A2(n19916), .ZN(n19156) );
  AND2_X1 U11813 ( .A1(n11023), .A2(n13832), .ZN(n19162) );
  NAND2_X1 U11814 ( .A1(n10146), .A2(n9846), .ZN(n10699) );
  XNOR2_X1 U11815 ( .A(n11022), .B(n11021), .ZN(n15047) );
  NAND2_X1 U11816 ( .A1(n12382), .A2(n12379), .ZN(n16266) );
  AND2_X1 U11817 ( .A1(n12382), .A2(n19938), .ZN(n19182) );
  INV_X1 U11818 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19908) );
  NAND2_X1 U11819 ( .A1(n16551), .A2(n16907), .ZN(n10030) );
  AND2_X1 U11820 ( .A1(n10005), .A2(n16815), .ZN(n16598) );
  NOR2_X2 U11821 ( .A1(n18679), .A2(n16525), .ZN(n16876) );
  INV_X1 U11822 ( .A(n17263), .ZN(n18222) );
  NOR2_X1 U11823 ( .A1(n17115), .A2(n17131), .ZN(n17101) );
  AND2_X1 U11824 ( .A1(n17101), .A2(P3_EBX_REG_13__SCAN_IN), .ZN(n17074) );
  NAND2_X1 U11825 ( .A1(n17145), .A2(P3_EBX_REG_11__SCAN_IN), .ZN(n17131) );
  AND2_X1 U11826 ( .A1(n17183), .A2(P3_EBX_REG_9__SCAN_IN), .ZN(n17133) );
  AND2_X1 U11827 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17186), .ZN(n17183) );
  INV_X1 U11828 ( .A(n17212), .ZN(n17215) );
  NOR2_X2 U11829 ( .A1(n17215), .A2(n18222), .ZN(n17216) );
  INV_X1 U11830 ( .A(n16403), .ZN(n17342) );
  NAND2_X1 U11831 ( .A1(n17692), .A2(n17658), .ZN(n9901) );
  NOR2_X1 U11832 ( .A1(n9896), .A2(n9895), .ZN(n9894) );
  NOR2_X1 U11833 ( .A1(n17764), .A2(n17997), .ZN(n9895) );
  AND2_X1 U11834 ( .A1(n9898), .A2(n17995), .ZN(n9897) );
  INV_X1 U11835 ( .A(n11252), .ZN(n9881) );
  INV_X1 U11836 ( .A(n9887), .ZN(n9883) );
  AOI21_X1 U11837 ( .B1(n9889), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n9759), .ZN(
        n9887) );
  INV_X1 U11838 ( .A(n11251), .ZN(n9886) );
  NOR2_X1 U11839 ( .A1(n11266), .A2(n9782), .ZN(n9889) );
  NAND2_X1 U11840 ( .A1(n11121), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11037) );
  AND2_X1 U11841 ( .A1(n10595), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10537) );
  NAND2_X1 U11842 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10287) );
  NAND2_X1 U11843 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10309) );
  OR2_X1 U11844 ( .A1(n11857), .A2(n11863), .ZN(n11859) );
  AND2_X1 U11845 ( .A1(n11859), .A2(n11850), .ZN(n11876) );
  NAND2_X1 U11846 ( .A1(n11877), .A2(n11854), .ZN(n11886) );
  NAND2_X1 U11847 ( .A1(n11204), .A2(n20209), .ZN(n11091) );
  NAND2_X1 U11848 ( .A1(n9851), .A2(n20209), .ZN(n12411) );
  NAND2_X1 U11849 ( .A1(n13181), .A2(n11155), .ZN(n9851) );
  OR2_X1 U11850 ( .A1(n11278), .A2(n11277), .ZN(n12464) );
  NOR2_X1 U11851 ( .A1(n11262), .A2(n11261), .ZN(n12449) );
  NOR2_X1 U11852 ( .A1(n11205), .A2(n20773), .ZN(n11208) );
  OR2_X1 U11853 ( .A1(n11174), .A2(n11173), .ZN(n12431) );
  INV_X1 U11854 ( .A(n11208), .ZN(n12424) );
  INV_X1 U11855 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11025) );
  INV_X1 U11856 ( .A(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11026) );
  NOR2_X1 U11857 ( .A1(n11027), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11035) );
  NOR2_X1 U11858 ( .A1(n12774), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11046) );
  OR2_X1 U11859 ( .A1(n11895), .A2(n11856), .ZN(n11896) );
  AND2_X1 U11860 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19924), .ZN(
        n10700) );
  INV_X1 U11861 ( .A(n13680), .ZN(n9917) );
  OR2_X1 U11862 ( .A1(n10588), .A2(n10587), .ZN(n12129) );
  NAND2_X1 U11863 ( .A1(n10398), .A2(n10397), .ZN(n10433) );
  NAND2_X1 U11864 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10294) );
  AOI22_X1 U11865 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10509), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10329) );
  NOR2_X1 U11866 ( .A1(n17358), .A2(n15739), .ZN(n15734) );
  NAND2_X1 U11867 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15389) );
  NAND2_X1 U11868 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n11855), .ZN(
        n11911) );
  AND2_X1 U11869 ( .A1(n11332), .A2(n11330), .ZN(n11163) );
  XNOR2_X1 U11870 ( .A(n11149), .B(n11218), .ZN(n20285) );
  NAND2_X1 U11871 ( .A1(n10181), .A2(n13924), .ZN(n10180) );
  INV_X1 U11872 ( .A(n13940), .ZN(n10181) );
  NOR2_X1 U11873 ( .A1(n10175), .A2(n10174), .ZN(n10173) );
  INV_X1 U11874 ( .A(n14173), .ZN(n10174) );
  INV_X1 U11875 ( .A(n11842), .ZN(n11806) );
  NAND2_X1 U11876 ( .A1(n14066), .A2(n10176), .ZN(n10175) );
  INV_X1 U11877 ( .A(n14271), .ZN(n10176) );
  NAND2_X1 U11878 ( .A1(n9829), .A2(n9769), .ZN(n10185) );
  NAND2_X1 U11879 ( .A1(n10186), .A2(n11446), .ZN(n14104) );
  OR2_X1 U11880 ( .A1(n11186), .A2(n11185), .ZN(n12496) );
  AND2_X1 U11881 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11308), .ZN(
        n11347) );
  NAND2_X1 U11882 ( .A1(n10056), .A2(n14314), .ZN(n10055) );
  NAND2_X1 U11883 ( .A1(n10039), .A2(n10038), .ZN(n10037) );
  NAND2_X1 U11884 ( .A1(n14444), .A2(n12501), .ZN(n14409) );
  NAND2_X1 U11885 ( .A1(n11922), .A2(n20166), .ZN(n12005) );
  OR2_X1 U11886 ( .A1(n11200), .A2(n11199), .ZN(n12439) );
  INV_X1 U11887 ( .A(n10130), .ZN(n10129) );
  OAI21_X1 U11888 ( .B1(n11203), .B2(n10131), .A(n12485), .ZN(n10130) );
  NOR2_X1 U11889 ( .A1(n12970), .A2(n20198), .ZN(n10046) );
  INV_X1 U11890 ( .A(n11143), .ZN(n11154) );
  AND2_X1 U11891 ( .A1(n15820), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11246) );
  NAND2_X1 U11892 ( .A1(n12762), .A2(n9866), .ZN(n12993) );
  INV_X1 U11893 ( .A(n9867), .ZN(n9866) );
  OAI21_X1 U11894 ( .B1(n11143), .B2(n12763), .A(n12789), .ZN(n9867) );
  INV_X1 U11895 ( .A(n11053), .ZN(n9850) );
  NAND3_X1 U11896 ( .A1(n11054), .A2(n11055), .A3(n11056), .ZN(n9849) );
  NAND2_X1 U11897 ( .A1(n12753), .A2(n20773), .ZN(n11244) );
  INV_X1 U11898 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20566) );
  INV_X1 U11899 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20492) );
  NAND2_X1 U11900 ( .A1(n11898), .A2(n12485), .ZN(n11904) );
  INV_X1 U11901 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n10109) );
  NOR2_X1 U11902 ( .A1(n10929), .A2(n10113), .ZN(n10112) );
  NAND2_X1 U11903 ( .A1(n10935), .A2(n10930), .ZN(n10113) );
  INV_X1 U11904 ( .A(n10897), .ZN(n10106) );
  NOR2_X1 U11905 ( .A1(n10900), .A2(n10108), .ZN(n10107) );
  INV_X1 U11906 ( .A(n10890), .ZN(n10108) );
  NAND2_X1 U11907 ( .A1(n10101), .A2(n10100), .ZN(n10876) );
  NAND2_X1 U11908 ( .A1(n11016), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10100) );
  NAND2_X1 U11909 ( .A1(n10862), .A2(n10102), .ZN(n10101) );
  NOR2_X1 U11910 ( .A1(n10214), .A2(n10213), .ZN(n10212) );
  INV_X1 U11911 ( .A(n14873), .ZN(n10214) );
  INV_X1 U11912 ( .A(n14696), .ZN(n10213) );
  NAND2_X1 U11913 ( .A1(n10254), .A2(n10267), .ZN(n10253) );
  INV_X1 U11914 ( .A(n14795), .ZN(n10254) );
  NOR2_X1 U11915 ( .A1(n10613), .A2(n10612), .ZN(n12097) );
  NAND2_X1 U11916 ( .A1(n10338), .A2(n12956), .ZN(n10345) );
  NOR2_X1 U11917 ( .A1(n9983), .A2(n9981), .ZN(n9980) );
  INV_X1 U11918 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n9981) );
  NAND2_X1 U11919 ( .A1(n10443), .A2(n10442), .ZN(n10469) );
  OAI21_X1 U11920 ( .B1(n10441), .B2(n10473), .A(n10470), .ZN(n10443) );
  NAND2_X1 U11921 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12079) );
  INV_X1 U11922 ( .A(n13571), .ZN(n10087) );
  AND2_X1 U11923 ( .A1(n11003), .A2(n9964), .ZN(n9963) );
  NOR2_X1 U11924 ( .A1(n14915), .A2(n9965), .ZN(n9964) );
  INV_X1 U11925 ( .A(n14924), .ZN(n9965) );
  INV_X1 U11926 ( .A(n14851), .ZN(n10222) );
  NAND2_X1 U11927 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n9941) );
  NAND2_X1 U11928 ( .A1(n9929), .A2(n10915), .ZN(n9927) );
  INV_X1 U11929 ( .A(n15149), .ZN(n9974) );
  INV_X1 U11930 ( .A(n15290), .ZN(n9978) );
  AND2_X1 U11931 ( .A1(n12248), .A2(n12247), .ZN(n15201) );
  AND2_X1 U11932 ( .A1(n10769), .A2(n10768), .ZN(n13228) );
  NOR2_X1 U11933 ( .A1(n16177), .A2(n15328), .ZN(n9951) );
  OR2_X1 U11934 ( .A1(n10691), .A2(n16246), .ZN(n10692) );
  NOR2_X1 U11935 ( .A1(n10206), .A2(n10194), .ZN(n10193) );
  INV_X1 U11936 ( .A(n10207), .ZN(n10194) );
  INV_X1 U11937 ( .A(n10200), .ZN(n10198) );
  INV_X1 U11938 ( .A(n12751), .ZN(n10197) );
  NAND2_X1 U11939 ( .A1(n10157), .A2(n18985), .ZN(n10893) );
  NAND2_X1 U11940 ( .A1(n10466), .A2(n10465), .ZN(n10743) );
  NOR2_X1 U11941 ( .A1(n10562), .A2(n10561), .ZN(n12109) );
  OR2_X1 U11942 ( .A1(n10524), .A2(n10523), .ZN(n12126) );
  NAND2_X1 U11943 ( .A1(n10401), .A2(n16302), .ZN(n10407) );
  OR2_X1 U11944 ( .A1(n12358), .A2(n12357), .ZN(n12954) );
  NAND2_X1 U11945 ( .A1(n10479), .A2(n19155), .ZN(n10491) );
  NAND3_X1 U11946 ( .A1(n12882), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19753), 
        .ZN(n19204) );
  INV_X1 U11947 ( .A(n12327), .ZN(n12330) );
  OR2_X1 U11948 ( .A1(n16885), .A2(n15388), .ZN(n9783) );
  NOR2_X1 U11949 ( .A1(n15388), .A2(n15387), .ZN(n15396) );
  NOR2_X1 U11950 ( .A1(n16885), .A2(n15384), .ZN(n15671) );
  NOR2_X1 U11951 ( .A1(n15385), .A2(n15384), .ZN(n15647) );
  INV_X1 U11952 ( .A(n15378), .ZN(n17169) );
  NAND2_X1 U11953 ( .A1(n15601), .A2(n18197), .ZN(n15586) );
  OR2_X1 U11954 ( .A1(n10240), .A2(n17515), .ZN(n9934) );
  NAND2_X1 U11955 ( .A1(n9793), .A2(n10241), .ZN(n10240) );
  NAND2_X1 U11956 ( .A1(n17761), .A2(n17866), .ZN(n10241) );
  NOR2_X1 U11957 ( .A1(n17777), .A2(n18094), .ZN(n15722) );
  INV_X1 U11958 ( .A(n15598), .ZN(n16514) );
  NOR2_X1 U11959 ( .A1(n17761), .A2(n15761), .ZN(n17722) );
  NAND2_X1 U11960 ( .A1(n17772), .A2(n15751), .ZN(n15761) );
  NAND2_X1 U11961 ( .A1(n17784), .A2(n15747), .ZN(n15749) );
  INV_X1 U11962 ( .A(n18210), .ZN(n15560) );
  NAND2_X1 U11963 ( .A1(n15425), .A2(n9905), .ZN(n15574) );
  NOR2_X1 U11964 ( .A1(n9907), .A2(n9906), .ZN(n9905) );
  INV_X1 U11965 ( .A(n15427), .ZN(n9906) );
  OR2_X1 U11966 ( .A1(n9860), .A2(n15433), .ZN(n15608) );
  NAND2_X1 U11967 ( .A1(n9904), .A2(n9903), .ZN(n17376) );
  INV_X1 U11968 ( .A(n18847), .ZN(n9903) );
  INV_X1 U11969 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15881) );
  OR3_X1 U11970 ( .A1(n20854), .A2(n15817), .A3(n11916), .ZN(n19982) );
  OR2_X1 U11971 ( .A1(n20005), .A2(n20003), .ZN(n14112) );
  AND2_X1 U11972 ( .A1(n14109), .A2(n9815), .ZN(n14176) );
  NAND2_X1 U11973 ( .A1(n14109), .A2(n10063), .ZN(n15872) );
  OR2_X1 U11974 ( .A1(n13187), .A2(n13186), .ZN(n13235) );
  INV_X1 U11975 ( .A(n14078), .ZN(n11507) );
  INV_X1 U11976 ( .A(n20159), .ZN(n20160) );
  OR2_X1 U11977 ( .A1(n11811), .A2(n14298), .ZN(n11918) );
  NOR2_X1 U11978 ( .A1(n11760), .A2(n14325), .ZN(n11761) );
  NAND2_X1 U11979 ( .A1(n11761), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11811) );
  NAND2_X1 U11980 ( .A1(n11723), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11724) );
  OR2_X1 U11981 ( .A1(n11724), .A2(n13968), .ZN(n11760) );
  INV_X1 U11982 ( .A(n11720), .ZN(n11723) );
  NAND2_X1 U11983 ( .A1(n11696), .A2(n10164), .ZN(n10163) );
  INV_X1 U11984 ( .A(n10165), .ZN(n10164) );
  NAND2_X1 U11985 ( .A1(n11635), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11692) );
  INV_X1 U11986 ( .A(n11636), .ZN(n11635) );
  AND2_X1 U11987 ( .A1(n11634), .A2(n11633), .ZN(n14016) );
  OR2_X1 U11988 ( .A1(n14368), .A2(n11845), .ZN(n11633) );
  CLKBUF_X1 U11989 ( .A(n14030), .Z(n14031) );
  CLKBUF_X1 U11990 ( .A(n14047), .Z(n14048) );
  AND2_X1 U11991 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n11559), .ZN(
        n11560) );
  INV_X1 U11992 ( .A(n11558), .ZN(n11559) );
  NOR2_X1 U11993 ( .A1(n11523), .A2(n14083), .ZN(n11524) );
  NAND2_X1 U11994 ( .A1(n11524), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11558) );
  NAND2_X1 U11995 ( .A1(n11491), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11523) );
  NOR2_X1 U11996 ( .A1(n11476), .A2(n14111), .ZN(n11491) );
  OR2_X1 U11997 ( .A1(n11471), .A2(n15881), .ZN(n11476) );
  AND2_X1 U11998 ( .A1(n11441), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11442) );
  NOR2_X1 U11999 ( .A1(n11426), .A2(n13521), .ZN(n11441) );
  NAND2_X1 U12000 ( .A1(n11376), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11401) );
  NOR2_X1 U12001 ( .A1(n11375), .A2(n11379), .ZN(n11376) );
  AOI21_X1 U12002 ( .B1(n12473), .B2(n11500), .A(n11383), .ZN(n13411) );
  NAND2_X1 U12003 ( .A1(n11369), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11375) );
  INV_X1 U12004 ( .A(n13265), .ZN(n11372) );
  AND2_X1 U12005 ( .A1(n11347), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11369) );
  AOI21_X1 U12006 ( .B1(n11316), .B2(n10179), .A(n10178), .ZN(n10177) );
  INV_X1 U12007 ( .A(n11342), .ZN(n10178) );
  NAND2_X1 U12008 ( .A1(n12005), .A2(n13909), .ZN(n13006) );
  NAND2_X1 U12009 ( .A1(n9879), .A2(n9876), .ZN(n9875) );
  NAND2_X1 U12010 ( .A1(n15937), .A2(n10115), .ZN(n9876) );
  NAND2_X1 U12011 ( .A1(n12522), .A2(n9774), .ZN(n9874) );
  NAND2_X1 U12012 ( .A1(n14301), .A2(n9811), .ZN(n10049) );
  NOR2_X1 U12013 ( .A1(n13938), .A2(n13926), .ZN(n13925) );
  OR2_X1 U12014 ( .A1(n13951), .A2(n13936), .ZN(n13938) );
  OR2_X1 U12015 ( .A1(n13965), .A2(n13949), .ZN(n13951) );
  NAND2_X1 U12016 ( .A1(n10067), .A2(n10066), .ZN(n10065) );
  NOR2_X1 U12017 ( .A1(n10068), .A2(n13998), .ZN(n10067) );
  INV_X1 U12018 ( .A(n11988), .ZN(n10066) );
  INV_X1 U12019 ( .A(n14308), .ZN(n14361) );
  NOR3_X1 U12020 ( .A1(n14170), .A2(n11988), .A3(n10069), .ZN(n14017) );
  NOR2_X1 U12021 ( .A1(n14170), .A2(n11988), .ZN(n14035) );
  NAND2_X1 U12022 ( .A1(n9892), .A2(n10123), .ZN(n14405) );
  NAND2_X1 U12023 ( .A1(n14444), .A2(n9891), .ZN(n9892) );
  INV_X1 U12024 ( .A(n10125), .ZN(n10041) );
  NOR2_X1 U12025 ( .A1(n15923), .A2(n21157), .ZN(n10032) );
  NAND2_X1 U12026 ( .A1(n14109), .A2(n14094), .ZN(n14096) );
  NOR2_X1 U12027 ( .A1(n10075), .A2(n15890), .ZN(n10074) );
  INV_X1 U12028 ( .A(n10077), .ZN(n10075) );
  NAND2_X1 U12029 ( .A1(n10076), .A2(n10077), .ZN(n15891) );
  NOR2_X1 U12030 ( .A1(n13499), .A2(n10079), .ZN(n13537) );
  NOR2_X1 U12031 ( .A1(n13499), .A2(n13500), .ZN(n13518) );
  OR2_X1 U12032 ( .A1(n13469), .A2(n13468), .ZN(n13499) );
  NAND2_X1 U12033 ( .A1(n15954), .A2(n9865), .ZN(n9859) );
  INV_X1 U12034 ( .A(n20858), .ZN(n13002) );
  NOR2_X1 U12035 ( .A1(n13187), .A2(n10071), .ZN(n16036) );
  NAND2_X1 U12036 ( .A1(n15954), .A2(n15953), .ZN(n15952) );
  OR2_X1 U12037 ( .A1(n13187), .A2(n10070), .ZN(n16032) );
  INV_X1 U12038 ( .A(n10072), .ZN(n10070) );
  NAND2_X1 U12039 ( .A1(n9871), .A2(n12448), .ZN(n9870) );
  NAND2_X1 U12040 ( .A1(n9855), .A2(n9789), .ZN(n9854) );
  NAND2_X1 U12041 ( .A1(n13197), .A2(n13196), .ZN(n13195) );
  INV_X1 U12042 ( .A(n20142), .ZN(n14616) );
  AND2_X1 U12043 ( .A1(n12996), .A2(n12995), .ZN(n14614) );
  NAND2_X1 U12044 ( .A1(n12934), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12933) );
  NAND2_X1 U12045 ( .A1(n10132), .A2(n9792), .ZN(n10135) );
  INV_X1 U12047 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20565) );
  NOR2_X1 U12048 ( .A1(n11129), .A2(n10034), .ZN(n10033) );
  AND3_X1 U12049 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20773), .A3(n20165), 
        .ZN(n20210) );
  NAND2_X1 U12050 ( .A1(n20247), .A2(n20164), .ZN(n20535) );
  NOR2_X2 U12051 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20717) );
  AOI21_X1 U12052 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20602), .A(n20327), 
        .ZN(n20716) );
  AND2_X1 U12053 ( .A1(n12364), .A2(n12365), .ZN(n16293) );
  CLKBUF_X1 U12054 ( .A(n10720), .Z(n10721) );
  NAND2_X1 U12055 ( .A1(n14815), .A2(n14814), .ZN(n14813) );
  NOR2_X1 U12056 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n16097), .ZN(n16082) );
  NOR2_X1 U12057 ( .A1(n10994), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10995) );
  AND2_X1 U12058 ( .A1(n10994), .A2(n10987), .ZN(n12552) );
  AND2_X1 U12059 ( .A1(n15203), .A2(n9826), .ZN(n15153) );
  NOR2_X1 U12060 ( .A1(n10929), .A2(n10111), .ZN(n10110) );
  INV_X1 U12061 ( .A(n10935), .ZN(n10111) );
  NAND2_X1 U12062 ( .A1(n10943), .A2(n9766), .ZN(n10937) );
  NAND2_X1 U12063 ( .A1(n10943), .A2(n10941), .ZN(n10945) );
  AND2_X1 U12064 ( .A1(n10891), .A2(n9786), .ZN(n10907) );
  NAND2_X1 U12065 ( .A1(n10891), .A2(n10890), .ZN(n10902) );
  AND2_X1 U12066 ( .A1(n10826), .A2(n10825), .ZN(n14678) );
  AND2_X1 U12067 ( .A1(n10785), .A2(n10784), .ZN(n12542) );
  INV_X1 U12068 ( .A(n10246), .ZN(n10245) );
  NAND2_X1 U12069 ( .A1(n14735), .A2(n13763), .ZN(n10244) );
  CLKBUF_X1 U12070 ( .A(n14769), .Z(n14770) );
  NOR2_X1 U12071 ( .A1(n15202), .A2(n15201), .ZN(n15203) );
  AND2_X1 U12072 ( .A1(n15203), .A2(n14873), .ZN(n14871) );
  INV_X1 U12073 ( .A(n15234), .ZN(n12246) );
  NAND2_X1 U12074 ( .A1(n12246), .A2(n14880), .ZN(n15202) );
  CLKBUF_X1 U12075 ( .A(n13575), .Z(n13496) );
  NAND2_X1 U12076 ( .A1(n12108), .A2(n12107), .ZN(n10188) );
  OR2_X1 U12077 ( .A1(n16267), .A2(n12241), .ZN(n12108) );
  NOR3_X1 U12078 ( .A1(n12055), .A2(n16078), .A3(n14668), .ZN(n12052) );
  INV_X1 U12079 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14668) );
  AND2_X1 U12080 ( .A1(n10814), .A2(n10813), .ZN(n14766) );
  NAND2_X1 U12081 ( .A1(n10091), .A2(n10090), .ZN(n10089) );
  NOR2_X1 U12082 ( .A1(n10094), .A2(n12567), .ZN(n10090) );
  INV_X1 U12083 ( .A(n10092), .ZN(n10091) );
  INV_X1 U12084 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14960) );
  CLKBUF_X1 U12085 ( .A(n12064), .Z(n12090) );
  INV_X1 U12086 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14984) );
  CLKBUF_X1 U12087 ( .A(n12088), .Z(n12091) );
  NOR2_X1 U12088 ( .A1(n14805), .A2(n14797), .ZN(n14799) );
  NOR3_X1 U12089 ( .A1(n14805), .A2(n10094), .A3(n14797), .ZN(n14790) );
  AND2_X1 U12090 ( .A1(n9985), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9984) );
  NOR2_X1 U12091 ( .A1(n15252), .A2(n15260), .ZN(n9958) );
  CLKBUF_X1 U12092 ( .A(n12066), .Z(n12085) );
  AND2_X1 U12093 ( .A1(n10781), .A2(n10780), .ZN(n13390) );
  NAND2_X1 U12094 ( .A1(n10082), .A2(n10081), .ZN(n13393) );
  INV_X1 U12095 ( .A(n13390), .ZN(n10081) );
  CLKBUF_X1 U12096 ( .A(n12068), .Z(n12084) );
  CLKBUF_X1 U12097 ( .A(n12070), .Z(n12083) );
  AND2_X1 U12098 ( .A1(n13042), .A2(n9801), .ZN(n13240) );
  INV_X1 U12099 ( .A(n13116), .ZN(n10095) );
  CLKBUF_X1 U12100 ( .A(n12072), .Z(n12082) );
  NAND2_X1 U12101 ( .A1(n13042), .A2(n10096), .ZN(n13115) );
  AND2_X1 U12102 ( .A1(n10742), .A2(n10741), .ZN(n13032) );
  AND2_X1 U12103 ( .A1(n13042), .A2(n10097), .ZN(n13046) );
  CLKBUF_X1 U12104 ( .A(n12074), .Z(n12081) );
  NAND2_X1 U12105 ( .A1(n13042), .A2(n13043), .ZN(n13041) );
  AND2_X1 U12106 ( .A1(n10753), .A2(n10752), .ZN(n12904) );
  CLKBUF_X1 U12107 ( .A(n12076), .Z(n12080) );
  INV_X1 U12108 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n21074) );
  NOR2_X1 U12109 ( .A1(n15103), .A2(n9941), .ZN(n9940) );
  XNOR2_X1 U12110 ( .A(n15052), .B(n15051), .ZN(n16056) );
  AND4_X1 U12111 ( .A1(n10672), .A2(n10671), .A3(n10670), .A4(n10669), .ZN(
        n10683) );
  AND4_X1 U12112 ( .A1(n10676), .A2(n10675), .A3(n10674), .A4(n10673), .ZN(
        n10682) );
  AND2_X1 U12113 ( .A1(n14852), .A2(n9836), .ZN(n14828) );
  INV_X1 U12114 ( .A(n14829), .ZN(n10220) );
  NAND2_X1 U12115 ( .A1(n14852), .A2(n9823), .ZN(n14839) );
  AND2_X1 U12116 ( .A1(n15110), .A2(n12373), .ZN(n15089) );
  OR2_X1 U12117 ( .A1(n14756), .A2(n14678), .ZN(n14738) );
  AND2_X1 U12118 ( .A1(n10830), .A2(n10829), .ZN(n14737) );
  NAND2_X1 U12119 ( .A1(n14852), .A2(n9821), .ZN(n14837) );
  INV_X1 U12120 ( .A(n9941), .ZN(n9939) );
  NAND2_X1 U12121 ( .A1(n14852), .A2(n14851), .ZN(n14854) );
  OR2_X1 U12122 ( .A1(n14754), .A2(n14753), .ZN(n14756) );
  NAND2_X1 U12123 ( .A1(n10146), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14936) );
  INV_X1 U12124 ( .A(n10924), .ZN(n9979) );
  OR2_X1 U12125 ( .A1(n15781), .A2(n10982), .ZN(n15148) );
  NOR2_X1 U12126 ( .A1(n14993), .A2(n15195), .ZN(n14983) );
  OR2_X1 U12127 ( .A1(n15002), .A2(n20943), .ZN(n14993) );
  NOR2_X1 U12128 ( .A1(n13393), .A2(n12542), .ZN(n13484) );
  NAND2_X1 U12129 ( .A1(n13484), .A2(n13483), .ZN(n14806) );
  NOR2_X1 U12130 ( .A1(n13219), .A2(n12544), .ZN(n15232) );
  NAND2_X1 U12131 ( .A1(n15273), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15025) );
  OR2_X1 U12132 ( .A1(n10216), .A2(n10219), .ZN(n10215) );
  INV_X1 U12133 ( .A(n13209), .ZN(n10219) );
  NAND2_X1 U12134 ( .A1(n9930), .A2(n9928), .ZN(n9926) );
  NAND2_X1 U12135 ( .A1(n9796), .A2(n9954), .ZN(n16176) );
  OAI211_X1 U12136 ( .C1(n10889), .C2(n13443), .A(n10661), .B(n9950), .ZN(
        n15346) );
  NAND2_X1 U12137 ( .A1(n15346), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15345) );
  NAND2_X1 U12138 ( .A1(n10888), .A2(n10887), .ZN(n15348) );
  CLKBUF_X1 U12139 ( .A(n12377), .Z(n12950) );
  CLKBUF_X1 U12140 ( .A(n12889), .Z(n12947) );
  NOR2_X1 U12141 ( .A1(n9924), .A2(n21153), .ZN(n9970) );
  NAND2_X1 U12142 ( .A1(n12124), .A2(n10191), .ZN(n13018) );
  NAND2_X1 U12143 ( .A1(n12681), .A2(n19576), .ZN(n12885) );
  AND2_X1 U12144 ( .A1(n16324), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12888) );
  INV_X1 U12145 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n21098) );
  NAND2_X1 U12146 ( .A1(n19909), .A2(n19910), .ZN(n19506) );
  AOI21_X2 U12147 ( .B1(n16324), .B2(n16327), .A(n15842), .ZN(n19682) );
  AND2_X1 U12148 ( .A1(n16330), .A2(n15841), .ZN(n15842) );
  OR2_X1 U12149 ( .A1(n19909), .A2(n19920), .ZN(n19640) );
  NAND2_X1 U12150 ( .A1(n9943), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9942) );
  NAND2_X1 U12151 ( .A1(n9945), .A2(n12956), .ZN(n9944) );
  INV_X1 U12152 ( .A(n19233), .ZN(n19249) );
  NAND2_X1 U12153 ( .A1(n19902), .A2(n19928), .ZN(n19678) );
  INV_X1 U12154 ( .A(n19247), .ZN(n19255) );
  OR2_X1 U12155 ( .A1(n19909), .A2(n19910), .ZN(n19899) );
  NOR2_X2 U12156 ( .A1(n19205), .A2(n19204), .ZN(n19246) );
  NOR2_X2 U12157 ( .A1(n13897), .A2(n19204), .ZN(n19247) );
  OR2_X1 U12158 ( .A1(n17416), .A2(n15587), .ZN(n9904) );
  OAI22_X1 U12159 ( .A1(n16340), .A2(n18658), .B1(n18655), .B2(n16339), .ZN(
        n18666) );
  NAND2_X1 U12160 ( .A1(n16528), .A2(n9765), .ZN(n16371) );
  NAND2_X1 U12161 ( .A1(n10010), .A2(n10008), .ZN(n10006) );
  OR2_X1 U12162 ( .A1(n16610), .A2(n9830), .ZN(n10003) );
  OR2_X1 U12163 ( .A1(n16610), .A2(n17550), .ZN(n10005) );
  NAND2_X1 U12164 ( .A1(n17088), .A2(P3_EBX_REG_15__SCAN_IN), .ZN(n17046) );
  INV_X1 U12165 ( .A(n16981), .ZN(n17080) );
  AOI211_X1 U12166 ( .C1(n9727), .C2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n15654), .B(n15653), .ZN(n15655) );
  AOI21_X1 U12167 ( .B1(n15602), .B2(n18660), .A(n15479), .ZN(n15845) );
  NOR3_X1 U12168 ( .A1(n17376), .A2(n18833), .A3(n17414), .ZN(n17394) );
  NOR2_X1 U12169 ( .A1(n18685), .A2(n18654), .ZN(n17415) );
  NOR2_X1 U12170 ( .A1(n17532), .A2(n17533), .ZN(n17518) );
  AND2_X1 U12171 ( .A1(n17639), .A2(n9816), .ZN(n17567) );
  INV_X1 U12172 ( .A(n17584), .ZN(n10012) );
  INV_X1 U12173 ( .A(n16658), .ZN(n17580) );
  NAND2_X1 U12174 ( .A1(n17639), .A2(n9760), .ZN(n17583) );
  NAND2_X1 U12175 ( .A1(n17639), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17617) );
  NOR2_X1 U12176 ( .A1(n16537), .A2(n17656), .ZN(n17639) );
  OR2_X1 U12177 ( .A1(n17663), .A2(n17659), .ZN(n9898) );
  NAND2_X1 U12178 ( .A1(n17661), .A2(n17992), .ZN(n9900) );
  NAND2_X1 U12179 ( .A1(n17660), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9899) );
  AND2_X1 U12180 ( .A1(n9757), .A2(n10022), .ZN(n17678) );
  NOR2_X1 U12181 ( .A1(n17787), .A2(n17703), .ZN(n10022) );
  NAND2_X1 U12182 ( .A1(n9757), .A2(n10025), .ZN(n17701) );
  INV_X1 U12183 ( .A(n17787), .ZN(n10025) );
  INV_X1 U12184 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17735) );
  NOR2_X1 U12185 ( .A1(n17787), .A2(n17788), .ZN(n17757) );
  AOI21_X1 U12186 ( .B1(n18136), .B2(n17822), .A(n15740), .ZN(n17814) );
  NOR2_X1 U12187 ( .A1(n17810), .A2(n17843), .ZN(n17790) );
  NOR2_X1 U12188 ( .A1(n18835), .A2(n16498), .ZN(n16353) );
  INV_X1 U12189 ( .A(n15828), .ZN(n16401) );
  NAND2_X1 U12190 ( .A1(n15770), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17505) );
  INV_X1 U12191 ( .A(n9934), .ZN(n15770) );
  OAI211_X1 U12192 ( .C1(n17896), .C2(n17529), .A(n17528), .B(n9813), .ZN(
        n17516) );
  NOR2_X1 U12193 ( .A1(n17516), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17515) );
  NOR3_X1 U12194 ( .A1(n17543), .A2(n17558), .A3(n17901), .ZN(n17529) );
  OR2_X1 U12195 ( .A1(n17761), .A2(n17543), .ZN(n17528) );
  NAND2_X1 U12196 ( .A1(n17605), .A2(n15767), .ZN(n17544) );
  NAND2_X1 U12197 ( .A1(n15768), .A2(n15764), .ZN(n15766) );
  NOR2_X1 U12198 ( .A1(n17544), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17543) );
  NAND2_X1 U12199 ( .A1(n17645), .A2(n17598), .ZN(n17605) );
  NAND2_X1 U12200 ( .A1(n17646), .A2(n17970), .ZN(n17645) );
  NAND2_X1 U12201 ( .A1(n17694), .A2(n10233), .ZN(n17650) );
  OR2_X1 U12202 ( .A1(n17761), .A2(n15763), .ZN(n10233) );
  NAND2_X1 U12203 ( .A1(n15761), .A2(n9937), .ZN(n17651) );
  AND2_X1 U12204 ( .A1(n15760), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9937) );
  NAND2_X1 U12205 ( .A1(n17662), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17976) );
  INV_X1 U12206 ( .A(n17577), .ZN(n18000) );
  NOR2_X1 U12207 ( .A1(n18014), .A2(n17699), .ZN(n18015) );
  NOR2_X1 U12208 ( .A1(n17779), .A2(n17778), .ZN(n17777) );
  NAND2_X1 U12209 ( .A1(n17801), .A2(n15746), .ZN(n17785) );
  NAND2_X1 U12210 ( .A1(n17785), .A2(n17786), .ZN(n17784) );
  XNOR2_X1 U12211 ( .A(n15745), .B(n15744), .ZN(n17802) );
  NAND2_X1 U12212 ( .A1(n17802), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17801) );
  INV_X1 U12213 ( .A(n18658), .ZN(n18001) );
  XNOR2_X1 U12214 ( .A(n15737), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17838) );
  NAND2_X1 U12215 ( .A1(n15560), .A2(n18197), .ZN(n15611) );
  INV_X1 U12216 ( .A(n16885), .ZN(n18634) );
  INV_X1 U12217 ( .A(n18628), .ZN(n18643) );
  NAND2_X1 U12218 ( .A1(n15602), .A2(n18847), .ZN(n18659) );
  NAND2_X1 U12219 ( .A1(n15604), .A2(n15576), .ZN(n16515) );
  INV_X1 U12220 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18646) );
  INV_X1 U12221 ( .A(n15574), .ZN(n18200) );
  INV_X1 U12222 ( .A(n15608), .ZN(n18197) );
  INV_X1 U12223 ( .A(n15561), .ZN(n18206) );
  INV_X1 U12224 ( .A(n17222), .ZN(n18215) );
  INV_X1 U12225 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n16516) );
  OR2_X1 U12226 ( .A1(n12618), .A2(n19949), .ZN(n12605) );
  AND2_X1 U12227 ( .A1(n12023), .A2(n12021), .ZN(n20005) );
  INV_X1 U12228 ( .A(n20024), .ZN(n20006) );
  AND2_X1 U12229 ( .A1(n19982), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20024) );
  NOR2_X1 U12230 ( .A1(n11252), .A2(n20562), .ZN(n12858) );
  INV_X1 U12231 ( .A(n20005), .ZN(n19994) );
  AND2_X1 U12232 ( .A1(n12023), .A2(n12015), .ZN(n20025) );
  AND2_X1 U12233 ( .A1(n12023), .A2(n12022), .ZN(n20021) );
  OR2_X1 U12234 ( .A1(n13177), .A2(n19949), .ZN(n13184) );
  NAND2_X1 U12235 ( .A1(n20040), .A2(n13185), .ZN(n14196) );
  INV_X1 U12236 ( .A(n14197), .ZN(n14278) );
  INV_X1 U12237 ( .A(n14285), .ZN(n15905) );
  NAND2_X1 U12238 ( .A1(n12392), .A2(n13091), .ZN(n15908) );
  AOI21_X1 U12239 ( .B1(n12797), .B2(n12982), .A(n12391), .ZN(n12392) );
  NOR2_X1 U12240 ( .A1(n13069), .A2(n14273), .ZN(n14285) );
  NAND2_X1 U12241 ( .A1(n20077), .A2(n20050), .ZN(n20047) );
  INV_X2 U12242 ( .A(n20047), .ZN(n20074) );
  INV_X1 U12243 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14325) );
  INV_X1 U12244 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14399) );
  CLKBUF_X1 U12245 ( .A(n13529), .Z(n13530) );
  INV_X1 U12246 ( .A(n20161), .ZN(n20117) );
  OR2_X1 U12247 ( .A1(n16045), .A2(n20711), .ZN(n20161) );
  NAND2_X1 U12248 ( .A1(n14322), .A2(n14468), .ZN(n14303) );
  AND2_X1 U12249 ( .A1(n14533), .A2(n14463), .ZN(n14522) );
  INV_X1 U12250 ( .A(n20139), .ZN(n20127) );
  NOR2_X1 U12251 ( .A1(n14616), .A2(n14631), .ZN(n20140) );
  OR2_X1 U12252 ( .A1(n14555), .A2(n14557), .ZN(n20142) );
  INV_X1 U12253 ( .A(n14614), .ZN(n20141) );
  OR2_X1 U12254 ( .A1(n13005), .A2(n12988), .ZN(n20147) );
  NOR2_X1 U12255 ( .A1(n13005), .A2(n12987), .ZN(n14555) );
  INV_X1 U12256 ( .A(n20717), .ZN(n20711) );
  INV_X1 U12257 ( .A(n12987), .ZN(n15787) );
  INV_X1 U12258 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13568) );
  NOR2_X1 U12259 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n14657) );
  OAI211_X1 U12260 ( .C1(n20175), .C2(n11307), .A(n20497), .B(n20171), .ZN(
        n20216) );
  OAI21_X1 U12261 ( .B1(n20345), .B2(n20328), .A(n20655), .ZN(n20347) );
  INV_X1 U12262 ( .A(n20329), .ZN(n20346) );
  OAI211_X1 U12263 ( .C1(n20464), .C2(n20573), .A(n20497), .B(n20448), .ZN(
        n20466) );
  INV_X1 U12264 ( .A(n20442), .ZN(n20465) );
  OAI211_X1 U12265 ( .C1(n20500), .C2(n20499), .A(n20498), .B(n20497), .ZN(
        n20524) );
  OAI211_X1 U12266 ( .C1(n20657), .C2(n20656), .A(n20655), .B(n20654), .ZN(
        n20703) );
  INV_X1 U12267 ( .A(n20646), .ZN(n21195) );
  INV_X1 U12268 ( .A(n20665), .ZN(n20729) );
  INV_X1 U12269 ( .A(n20672), .ZN(n20735) );
  INV_X1 U12270 ( .A(n20684), .ZN(n20747) );
  OR2_X1 U12271 ( .A1(n20639), .A2(n20535), .ZN(n20759) );
  INV_X1 U12272 ( .A(n20691), .ZN(n20753) );
  INV_X1 U12273 ( .A(n20697), .ZN(n20762) );
  NOR2_X1 U12274 ( .A1(n20573), .A2(n12979), .ZN(n15823) );
  NOR2_X1 U12275 ( .A1(n11307), .A2(n20772), .ZN(n16047) );
  INV_X1 U12276 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20772) );
  INV_X1 U12277 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20573) );
  NAND2_X1 U12278 ( .A1(n9998), .A2(n19002), .ZN(n9997) );
  NOR2_X1 U12279 ( .A1(n11012), .A2(n11002), .ZN(n14672) );
  NOR2_X1 U12280 ( .A1(n12283), .A2(n12093), .ZN(n19032) );
  NAND2_X1 U12281 ( .A1(n14917), .A2(n9989), .ZN(n9988) );
  AND2_X1 U12282 ( .A1(n9991), .A2(n19002), .ZN(n16091) );
  INV_X1 U12283 ( .A(n9991), .ZN(n14675) );
  NAND2_X1 U12284 ( .A1(n9995), .A2(n16153), .ZN(n9993) );
  NAND2_X1 U12285 ( .A1(n9753), .A2(n9995), .ZN(n9992) );
  INV_X1 U12286 ( .A(n16138), .ZN(n9995) );
  INV_X1 U12287 ( .A(n9994), .ZN(n15777) );
  INV_X1 U12288 ( .A(n19037), .ZN(n18996) );
  AND2_X1 U12289 ( .A1(n12276), .A2(n12275), .ZN(n19026) );
  NOR2_X1 U12290 ( .A1(n19073), .A2(n12275), .ZN(n19015) );
  INV_X1 U12291 ( .A(n19820), .ZN(n19021) );
  INV_X1 U12292 ( .A(n19034), .ZN(n19020) );
  NOR2_X1 U12293 ( .A1(n10255), .A2(n9910), .ZN(n9909) );
  NAND2_X1 U12294 ( .A1(n10256), .A2(n13463), .ZN(n10255) );
  INV_X1 U12295 ( .A(n9912), .ZN(n9910) );
  OR2_X1 U12296 ( .A1(n12184), .A2(n12183), .ZN(n13227) );
  NOR2_X1 U12297 ( .A1(n12172), .A2(n12171), .ZN(n13243) );
  OR2_X1 U12298 ( .A1(n12158), .A2(n12157), .ZN(n13113) );
  CLKBUF_X1 U12299 ( .A(n13223), .Z(n13112) );
  OR2_X1 U12300 ( .A1(n12144), .A2(n12143), .ZN(n13050) );
  AND2_X1 U12301 ( .A1(n9767), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10250) );
  INV_X1 U12302 ( .A(n14811), .ZN(n14783) );
  OR2_X1 U12303 ( .A1(n12944), .A2(n12945), .ZN(n12946) );
  OR2_X1 U12304 ( .A1(n14804), .A2(n12851), .ZN(n14811) );
  CLKBUF_X1 U12305 ( .A(n14733), .Z(n14734) );
  CLKBUF_X1 U12306 ( .A(n14743), .Z(n14744) );
  CLKBUF_X1 U12307 ( .A(n14760), .Z(n14761) );
  INV_X1 U12308 ( .A(n19059), .ZN(n19044) );
  NOR2_X1 U12309 ( .A1(n12940), .A2(n13037), .ZN(n13060) );
  OR2_X1 U12310 ( .A1(n13136), .A2(n10203), .ZN(n10199) );
  NOR2_X1 U12311 ( .A1(n19064), .A2(n19055), .ZN(n19070) );
  INV_X1 U12312 ( .A(n16133), .ZN(n19064) );
  NOR2_X1 U12313 ( .A1(n12836), .A2(n12687), .ZN(n19265) );
  AND4_X1 U12314 ( .A1(n12686), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n12685), 
        .A4(n19576), .ZN(n12687) );
  AND2_X1 U12315 ( .A1(n19075), .A2(n19828), .ZN(n19131) );
  INV_X1 U12316 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14927) );
  INV_X1 U12317 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15019) );
  INV_X1 U12318 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16159) );
  AND2_X1 U12319 ( .A1(n13391), .A2(n13348), .ZN(n18933) );
  INV_X1 U12320 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16174) );
  NAND2_X1 U12321 ( .A1(n15335), .A2(n10690), .ZN(n16205) );
  INV_X1 U12322 ( .A(n19159), .ZN(n16186) );
  AND2_X1 U12323 ( .A1(n13274), .A2(n10144), .ZN(n13441) );
  INV_X1 U12324 ( .A(n16217), .ZN(n19152) );
  INV_X1 U12325 ( .A(n19156), .ZN(n16211) );
  INV_X1 U12326 ( .A(n19162), .ZN(n16219) );
  INV_X1 U12327 ( .A(n16225), .ZN(n19154) );
  NAND2_X1 U12328 ( .A1(n14899), .A2(n14896), .ZN(n10152) );
  OR2_X1 U12329 ( .A1(n13574), .A2(n13573), .ZN(n16070) );
  NAND2_X1 U12330 ( .A1(n14925), .A2(n14924), .ZN(n14913) );
  AND2_X1 U12331 ( .A1(n15337), .A2(n12371), .ZN(n15329) );
  NAND2_X1 U12332 ( .A1(n19202), .A2(n19175), .ZN(n9959) );
  AND2_X1 U12333 ( .A1(n10158), .A2(n10160), .ZN(n16179) );
  OR2_X1 U12334 ( .A1(n13279), .A2(n12360), .ZN(n15330) );
  NAND2_X1 U12335 ( .A1(n10158), .A2(n10904), .ZN(n15324) );
  INV_X1 U12336 ( .A(n10195), .ZN(n12752) );
  AOI21_X1 U12337 ( .B1(n10201), .B2(n10200), .A(n10206), .ZN(n10195) );
  NAND2_X1 U12338 ( .A1(n13136), .A2(n10207), .ZN(n10201) );
  NAND2_X1 U12339 ( .A1(n12382), .A2(n12367), .ZN(n16251) );
  NAND2_X1 U12340 ( .A1(n15040), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15335) );
  CLKBUF_X1 U12341 ( .A(n12947), .Z(n16255) );
  INV_X1 U12342 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19185) );
  AND2_X1 U12343 ( .A1(n12355), .A2(n16262), .ZN(n19186) );
  INV_X1 U12344 ( .A(n16266), .ZN(n19199) );
  AND2_X1 U12345 ( .A1(n19175), .A2(n15226), .ZN(n19192) );
  INV_X1 U12346 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19933) );
  INV_X1 U12347 ( .A(n19265), .ZN(n19928) );
  INV_X1 U12348 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19924) );
  XNOR2_X1 U12349 ( .A(n12863), .B(n12864), .ZN(n19920) );
  INV_X1 U12350 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19915) );
  INV_X1 U12351 ( .A(n19920), .ZN(n19910) );
  XNOR2_X1 U12352 ( .A(n12896), .B(n12897), .ZN(n19909) );
  INV_X1 U12353 ( .A(n19266), .ZN(n19902) );
  AOI21_X1 U12354 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n16324), .A(n12669), 
        .ZN(n15376) );
  NOR2_X1 U12355 ( .A1(n19899), .A2(n19413), .ZN(n19459) );
  NOR2_X1 U12356 ( .A1(n19899), .A2(n19450), .ZN(n19471) );
  INV_X1 U12357 ( .A(n19773), .ZN(n19614) );
  INV_X1 U12358 ( .A(n19787), .ZN(n19620) );
  INV_X1 U12359 ( .A(n19602), .ZN(n19632) );
  OAI22_X1 U12360 ( .A1(n19207), .A2(n19255), .B1(n19206), .B2(n19253), .ZN(
        n19688) );
  INV_X1 U12361 ( .A(n19772), .ZN(n19704) );
  AND2_X1 U12362 ( .A1(n19223), .A2(n19249), .ZN(n19703) );
  OAI21_X1 U12363 ( .B1(n19693), .B2(n19692), .A(n19691), .ZN(n19734) );
  INV_X1 U12364 ( .A(n19705), .ZN(n19736) );
  AND2_X1 U12365 ( .A1(n19250), .A2(n19249), .ZN(n19733) );
  INV_X1 U12366 ( .A(n19648), .ZN(n19755) );
  INV_X1 U12367 ( .A(n19688), .ZN(n19758) );
  INV_X1 U12368 ( .A(n19653), .ZN(n19762) );
  INV_X1 U12369 ( .A(n19726), .ZN(n19790) );
  INV_X1 U12370 ( .A(n19813), .ZN(n19798) );
  INV_X1 U12371 ( .A(n19809), .ZN(n19801) );
  NOR2_X1 U12372 ( .A1(n19899), .A2(n19633), .ZN(n19809) );
  OR2_X1 U12373 ( .A1(n12270), .A2(n19441), .ZN(n16333) );
  INV_X1 U12374 ( .A(n16333), .ZN(n19815) );
  INV_X2 U12375 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n16324) );
  INV_X1 U12376 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19576) );
  XNOR2_X1 U12377 ( .A(n16523), .B(n17377), .ZN(n18847) );
  INV_X1 U12378 ( .A(n9904), .ZN(n16497) );
  NOR2_X1 U12379 ( .A1(n16575), .A2(n16576), .ZN(n16574) );
  NOR2_X1 U12380 ( .A1(n16585), .A2(n16852), .ZN(n16575) );
  NOR2_X1 U12381 ( .A1(n18756), .A2(n16620), .ZN(n16618) );
  NOR2_X1 U12382 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16643), .ZN(n16629) );
  INV_X1 U12383 ( .A(n16862), .ZN(n16892) );
  NOR2_X1 U12384 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16705), .ZN(n16691) );
  NOR2_X1 U12385 ( .A1(n20974), .A2(n18695), .ZN(n16853) );
  NOR2_X1 U12386 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16763), .ZN(n16762) );
  NOR2_X1 U12387 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16798), .ZN(n16785) );
  INV_X1 U12388 ( .A(n16520), .ZN(n16893) );
  NOR2_X2 U12389 ( .A1(n18787), .A2(n16768), .ZN(n16880) );
  NAND4_X1 U12390 ( .A1(n18169), .A2(n18846), .A3(n18693), .A4(n18683), .ZN(
        n16897) );
  NAND2_X1 U12391 ( .A1(n16944), .A2(n9842), .ZN(n16938) );
  NAND2_X1 U12392 ( .A1(n16946), .A2(n17197), .ZN(n16944) );
  NAND2_X1 U12393 ( .A1(n16955), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n16946) );
  NOR2_X1 U12394 ( .A1(n16952), .A2(n16901), .ZN(n16955) );
  AND3_X1 U12395 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(P3_EBX_REG_19__SCAN_IN), 
        .A3(n16993), .ZN(n16991) );
  NOR2_X1 U12396 ( .A1(n17263), .A2(n17046), .ZN(n17059) );
  AND2_X1 U12397 ( .A1(n17074), .A2(P3_EBX_REG_14__SCAN_IN), .ZN(n17088) );
  AND2_X1 U12398 ( .A1(n17133), .A2(P3_EBX_REG_10__SCAN_IN), .ZN(n17145) );
  INV_X1 U12399 ( .A(n17195), .ZN(n17193) );
  NOR2_X1 U12400 ( .A1(n17215), .A2(n17202), .ZN(n17196) );
  NAND2_X1 U12401 ( .A1(n17196), .A2(P3_EBX_REG_4__SCAN_IN), .ZN(n17195) );
  NAND2_X1 U12402 ( .A1(n16523), .A2(n9864), .ZN(n9863) );
  NOR2_X1 U12403 ( .A1(n18183), .A2(n18685), .ZN(n9864) );
  INV_X1 U12404 ( .A(n17301), .ZN(n17290) );
  INV_X1 U12405 ( .A(n17271), .ZN(n17297) );
  NOR2_X1 U12406 ( .A1(n17368), .A2(n18222), .ZN(n17325) );
  NOR2_X1 U12407 ( .A1(n15634), .A2(n15633), .ZN(n17350) );
  INV_X1 U12408 ( .A(n17369), .ZN(n17367) );
  INV_X1 U12409 ( .A(n17335), .ZN(n17374) );
  NOR2_X1 U12410 ( .A1(n18642), .A2(n17362), .ZN(n17369) );
  OAI211_X1 U12411 ( .C1(n18835), .C2(n18836), .A(n17416), .B(n17415), .ZN(
        n17469) );
  NOR2_X1 U12412 ( .A1(n18835), .A2(n17479), .ZN(n17476) );
  BUF_X1 U12413 ( .A(n17469), .Z(n17479) );
  NAND2_X1 U12415 ( .A1(n10019), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10017) );
  OR2_X1 U12416 ( .A1(n16528), .A2(n16544), .ZN(n10016) );
  INV_X1 U12417 ( .A(n17702), .ZN(n17654) );
  NOR2_X1 U12418 ( .A1(n17973), .A2(n17976), .ZN(n17578) );
  NOR2_X1 U12419 ( .A1(n17843), .A2(n17856), .ZN(n17563) );
  NAND2_X1 U12420 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17790), .ZN(n17709) );
  INV_X1 U12421 ( .A(n17578), .ZN(n17998) );
  AND2_X1 U12422 ( .A1(n10027), .A2(n10026), .ZN(n17726) );
  NOR2_X1 U12423 ( .A1(n16349), .A2(n17735), .ZN(n10026) );
  NOR2_X1 U12424 ( .A1(n17767), .A2(n16774), .ZN(n10027) );
  INV_X1 U12425 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16349) );
  NOR2_X1 U12426 ( .A1(n17809), .A2(n17821), .ZN(n17806) );
  INV_X1 U12427 ( .A(n17850), .ZN(n17840) );
  INV_X1 U12428 ( .A(n18219), .ZN(n18566) );
  INV_X1 U12429 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17849) );
  INV_X1 U12430 ( .A(n17848), .ZN(n17861) );
  NAND2_X1 U12431 ( .A1(n16347), .A2(n10226), .ZN(n16397) );
  NAND2_X1 U12432 ( .A1(n16342), .A2(n10227), .ZN(n10226) );
  AND2_X1 U12433 ( .A1(n18154), .A2(n17939), .ZN(n17991) );
  OAI21_X1 U12434 ( .B1(n18002), .B2(n17975), .A(n18154), .ZN(n18076) );
  AND2_X1 U12435 ( .A1(n17772), .A2(n10236), .ZN(n17760) );
  NOR2_X1 U12436 ( .A1(n10238), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10236) );
  NAND2_X1 U12437 ( .A1(n10223), .A2(n17822), .ZN(n17824) );
  INV_X1 U12438 ( .A(n18659), .ZN(n18639) );
  INV_X1 U12439 ( .A(n18170), .ZN(n18154) );
  NAND2_X1 U12440 ( .A1(n15604), .A2(n15603), .ZN(n18628) );
  INV_X1 U12441 ( .A(n18130), .ZN(n18166) );
  INV_X1 U12442 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18477) );
  INV_X1 U12443 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21113) );
  INV_X1 U12444 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18665) );
  NAND2_X1 U12445 ( .A1(n16517), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18685) );
  INV_X1 U12446 ( .A(n14221), .ZN(n20159) );
  OAI21_X1 U12448 ( .B1(n14451), .B2(n19955), .A(n12523), .ZN(P1_U2968) );
  AND2_X1 U12449 ( .A1(n14473), .A2(n14474), .ZN(n9878) );
  OAI211_X1 U12450 ( .C1(n14481), .C2(n15986), .A(n10062), .B(n10059), .ZN(
        P1_U3001) );
  AOI21_X1 U12451 ( .B1(n14479), .B2(n14480), .A(n14478), .ZN(n10062) );
  NAND2_X1 U12452 ( .A1(n10060), .A2(n20133), .ZN(n10059) );
  AND2_X1 U12453 ( .A1(n10210), .A2(n9833), .ZN(n13904) );
  OR2_X1 U12454 ( .A1(n16132), .A2(n15067), .ZN(n10210) );
  AOI21_X1 U12455 ( .B1(n15047), .B2(n19162), .A(n10084), .ZN(n10083) );
  OAI21_X1 U12456 ( .B1(n15062), .B2(n19159), .A(n10085), .ZN(n10084) );
  OAI211_X1 U12457 ( .C1(n15058), .C2(n16266), .A(n10268), .B(n15057), .ZN(
        n15059) );
  OAI21_X1 U12458 ( .B1(n16546), .B2(n9843), .A(n10028), .ZN(P3_U2640) );
  NOR2_X1 U12459 ( .A1(n16542), .A2(n10029), .ZN(n10028) );
  INV_X1 U12460 ( .A(n17074), .ZN(n17100) );
  INV_X1 U12461 ( .A(n17133), .ZN(n17163) );
  NAND2_X1 U12462 ( .A1(n9902), .A2(n9893), .ZN(P3_U2814) );
  NAND2_X1 U12463 ( .A1(n17657), .A2(n17656), .ZN(n9902) );
  AND2_X1 U12464 ( .A1(n9901), .A2(n9894), .ZN(n9893) );
  INV_X1 U12465 ( .A(n10540), .ZN(n13627) );
  INV_X1 U12466 ( .A(n17008), .ZN(n15491) );
  BUF_X1 U12467 ( .A(n15491), .Z(n17167) );
  AND2_X1 U12468 ( .A1(n12067), .A2(n9985), .ZN(n9754) );
  AND2_X1 U12469 ( .A1(n9765), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9755) );
  NAND2_X1 U12470 ( .A1(n12094), .A2(n19576), .ZN(n12121) );
  INV_X1 U12471 ( .A(n10546), .ZN(n13625) );
  INV_X1 U12472 ( .A(n15671), .ZN(n15458) );
  NAND2_X1 U12473 ( .A1(n12063), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12062) );
  OR2_X1 U12474 ( .A1(n14030), .A2(n10168), .ZN(n9756) );
  NAND2_X1 U12475 ( .A1(n12067), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12065) );
  INV_X1 U12476 ( .A(n11327), .ZN(n10131) );
  AND2_X1 U12477 ( .A1(n17726), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9757) );
  INV_X1 U12478 ( .A(n11121), .ZN(n11711) );
  OR2_X1 U12479 ( .A1(n10655), .A2(n21153), .ZN(n9758) );
  NAND2_X1 U12480 ( .A1(n11131), .A2(n11328), .ZN(n11137) );
  AND2_X1 U12481 ( .A1(n11266), .A2(n9782), .ZN(n9759) );
  INV_X1 U12482 ( .A(n14887), .ZN(n10151) );
  AND2_X1 U12483 ( .A1(n10013), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9760) );
  OR2_X1 U12484 ( .A1(n17702), .A2(n16537), .ZN(n9761) );
  NAND2_X1 U12485 ( .A1(n12899), .A2(n12898), .ZN(n12944) );
  NOR2_X1 U12486 ( .A1(n14760), .A2(n13680), .ZN(n14749) );
  NAND2_X1 U12487 ( .A1(n10242), .A2(n10248), .ZN(n14726) );
  AND2_X1 U12488 ( .A1(n9994), .A2(n19002), .ZN(n9762) );
  AND2_X1 U12489 ( .A1(n10894), .A2(n9804), .ZN(n9763) );
  AND2_X1 U12490 ( .A1(n9797), .A2(n12500), .ZN(n9764) );
  NAND2_X1 U12491 ( .A1(n17947), .A2(n18643), .ZN(n17867) );
  INV_X1 U12492 ( .A(n17867), .ZN(n9908) );
  OR2_X1 U12493 ( .A1(n12209), .A2(n12208), .ZN(n13351) );
  NAND2_X1 U12494 ( .A1(n13352), .A2(n13351), .ZN(n13413) );
  NAND2_X1 U12495 ( .A1(n9911), .A2(n9909), .ZN(n9914) );
  AND2_X1 U12496 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n9765) );
  AND2_X1 U12497 ( .A1(n10941), .A2(n9825), .ZN(n9766) );
  AND2_X1 U12498 ( .A1(n12914), .A2(n13031), .ZN(n9767) );
  OR2_X1 U12499 ( .A1(n13575), .A2(n10253), .ZN(n9768) );
  OR2_X1 U12500 ( .A1(n10187), .A2(n11446), .ZN(n9769) );
  OR2_X2 U12501 ( .A1(n9914), .A2(n9845), .ZN(n13575) );
  NAND3_X1 U12502 ( .A1(n10016), .A2(n10015), .A3(n10017), .ZN(n16815) );
  INV_X1 U12503 ( .A(n19202), .ZN(n16231) );
  NAND2_X1 U12504 ( .A1(n12382), .A2(n19937), .ZN(n19202) );
  AND2_X1 U12505 ( .A1(n9827), .A2(n10087), .ZN(n9770) );
  AND2_X1 U12506 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n9771) );
  AND2_X1 U12507 ( .A1(n9771), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9772) );
  AND2_X1 U12508 ( .A1(n9772), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9773) );
  AND2_X1 U12509 ( .A1(n10115), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9774) );
  OR2_X1 U12510 ( .A1(n19250), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n9775) );
  NOR2_X1 U12511 ( .A1(n15385), .A2(n15389), .ZN(n15379) );
  NAND2_X1 U12512 ( .A1(n11035), .A2(n12777), .ZN(n11703) );
  OR2_X1 U12513 ( .A1(n14170), .A2(n10065), .ZN(n9777) );
  OR2_X1 U12514 ( .A1(n14805), .A2(n10089), .ZN(n9778) );
  AND2_X1 U12515 ( .A1(n14919), .A2(n9772), .ZN(n9780) );
  NOR2_X1 U12516 ( .A1(n14030), .A2(n10165), .ZN(n13990) );
  NOR2_X1 U12517 ( .A1(n14030), .A2(n14032), .ZN(n14015) );
  OR2_X1 U12518 ( .A1(n10973), .A2(n9979), .ZN(n9781) );
  NOR2_X1 U12519 ( .A1(n12449), .A2(n11263), .ZN(n9782) );
  BUF_X1 U12520 ( .A(n10381), .Z(n19227) );
  INV_X1 U12521 ( .A(n10206), .ZN(n10205) );
  NOR2_X1 U12522 ( .A1(n10981), .A2(n12241), .ZN(n10206) );
  NOR2_X1 U12523 ( .A1(n14077), .A2(n10175), .ZN(n14064) );
  NAND2_X1 U12524 ( .A1(n10170), .A2(n10173), .ZN(n14046) );
  NOR2_X1 U12525 ( .A1(n14077), .A2(n14271), .ZN(n14063) );
  AND2_X1 U12526 ( .A1(n9923), .A2(n9921), .ZN(n14925) );
  OAI21_X1 U12527 ( .B1(n15293), .B2(n9781), .A(n9975), .ZN(n15147) );
  NAND2_X1 U12528 ( .A1(n9930), .A2(n10912), .ZN(n15304) );
  INV_X1 U12529 ( .A(n10249), .ZN(n14719) );
  AND2_X1 U12530 ( .A1(n11119), .A2(n11117), .ZN(n9785) );
  AND2_X1 U12531 ( .A1(n10107), .A2(n10106), .ZN(n9786) );
  AND2_X1 U12532 ( .A1(n12901), .A2(n12895), .ZN(n12945) );
  NAND3_X1 U12533 ( .A1(n9885), .A2(n9882), .A3(n9880), .ZN(n11343) );
  OR2_X1 U12534 ( .A1(n13939), .A2(n10180), .ZN(n9787) );
  AND2_X1 U12535 ( .A1(n10146), .A2(n9939), .ZN(n9788) );
  AND2_X1 U12536 ( .A1(n12447), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9789) );
  NOR2_X1 U12537 ( .A1(n14749), .A2(n14750), .ZN(n9790) );
  NAND2_X1 U12538 ( .A1(n10865), .A2(n10399), .ZN(n10390) );
  AND2_X1 U12539 ( .A1(n16034), .A2(n16033), .ZN(n9791) );
  INV_X1 U12540 ( .A(n10690), .ZN(n10149) );
  AND2_X1 U12541 ( .A1(n11203), .A2(n10131), .ZN(n9792) );
  INV_X1 U12542 ( .A(n13529), .ZN(n10186) );
  INV_X1 U12543 ( .A(n14077), .ZN(n10170) );
  OR2_X1 U12544 ( .A1(n17529), .A2(n17598), .ZN(n9793) );
  AND2_X1 U12545 ( .A1(n10224), .A2(n15738), .ZN(n9794) );
  INV_X1 U12546 ( .A(n9933), .ZN(n17504) );
  NAND2_X1 U12547 ( .A1(n9934), .A2(n17871), .ZN(n9933) );
  AND2_X1 U12548 ( .A1(n9729), .A2(n20198), .ZN(n12485) );
  INV_X1 U12549 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12774) );
  INV_X1 U12550 ( .A(n11131), .ZN(n13181) );
  BUF_X1 U12551 ( .A(n11131), .Z(n20198) );
  AND2_X1 U12552 ( .A1(n9966), .A2(n13851), .ZN(n9795) );
  INV_X1 U12553 ( .A(n10040), .ZN(n10123) );
  NAND2_X1 U12554 ( .A1(n15909), .A2(n10124), .ZN(n10040) );
  AND2_X1 U12555 ( .A1(n9953), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9796) );
  OR2_X1 U12556 ( .A1(n15923), .A2(n13542), .ZN(n9797) );
  AND2_X1 U12557 ( .A1(n13763), .A2(n10247), .ZN(n9798) );
  AND2_X1 U12558 ( .A1(n10249), .A2(n10248), .ZN(n9799) );
  OAI21_X1 U12559 ( .B1(n16066), .B2(n10981), .A(n15076), .ZN(n14896) );
  AND2_X1 U12560 ( .A1(n9975), .A2(n9927), .ZN(n9800) );
  AND2_X1 U12561 ( .A1(n10096), .A2(n10095), .ZN(n9801) );
  NOR2_X1 U12562 ( .A1(n13529), .A2(n10185), .ZN(n14090) );
  NAND2_X1 U12563 ( .A1(n14803), .A2(n10267), .ZN(n14794) );
  NOR2_X1 U12564 ( .A1(n12076), .A2(n16224), .ZN(n12077) );
  NOR2_X1 U12565 ( .A1(n12072), .A2(n16195), .ZN(n12073) );
  NOR2_X1 U12566 ( .A1(n12068), .A2(n16159), .ZN(n12069) );
  AND3_X1 U12567 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12078) );
  AND2_X1 U12568 ( .A1(n17639), .A2(n10013), .ZN(n9802) );
  AND2_X1 U12569 ( .A1(n12063), .A2(n9980), .ZN(n9803) );
  NAND2_X1 U12570 ( .A1(n11244), .A2(n11243), .ZN(n11344) );
  NOR2_X1 U12571 ( .A1(n16198), .A2(n16196), .ZN(n9804) );
  AND2_X1 U12572 ( .A1(n15203), .A2(n10212), .ZN(n12569) );
  AND3_X1 U12573 ( .A1(n10153), .A2(n10154), .A3(n11385), .ZN(n13459) );
  NOR2_X1 U12574 ( .A1(n14806), .A2(n14807), .ZN(n10794) );
  AND2_X1 U12575 ( .A1(n11143), .A2(n11115), .ZN(n9805) );
  NAND2_X1 U12576 ( .A1(n9859), .A2(n10117), .ZN(n15946) );
  NAND2_X1 U12577 ( .A1(n10116), .A2(n12500), .ZN(n13541) );
  NAND2_X1 U12578 ( .A1(n15952), .A2(n12472), .ZN(n13421) );
  INV_X1 U12579 ( .A(n14342), .ZN(n15937) );
  NOR2_X1 U12580 ( .A1(n12940), .A2(n10215), .ZN(n13207) );
  NAND2_X1 U12581 ( .A1(n17773), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17772) );
  XNOR2_X1 U12582 ( .A(n12836), .B(n12834), .ZN(n12864) );
  OR3_X1 U12583 ( .A1(n14170), .A2(n11988), .A3(n10068), .ZN(n9806) );
  OR3_X1 U12584 ( .A1(n14805), .A2(n10092), .A3(n10094), .ZN(n9807) );
  AND2_X1 U12585 ( .A1(n14411), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9808) );
  INV_X1 U12586 ( .A(n10981), .ZN(n9924) );
  NAND2_X1 U12587 ( .A1(n12944), .A2(n12945), .ZN(n12943) );
  AND2_X1 U12588 ( .A1(n14068), .A2(n15871), .ZN(n9809) );
  OR2_X1 U12589 ( .A1(n12197), .A2(n12196), .ZN(n13249) );
  INV_X1 U12590 ( .A(n13249), .ZN(n9913) );
  NAND2_X1 U12591 ( .A1(n15305), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9810) );
  NOR2_X1 U12592 ( .A1(n15923), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9811) );
  OR2_X1 U12593 ( .A1(n16868), .A2(n16544), .ZN(n9812) );
  INV_X1 U12594 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17788) );
  OR2_X1 U12595 ( .A1(n17598), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9813) );
  INV_X1 U12596 ( .A(n9929), .ZN(n9928) );
  NAND2_X1 U12597 ( .A1(n10912), .A2(n9810), .ZN(n9929) );
  NOR2_X1 U12598 ( .A1(n14424), .A2(n10032), .ZN(n9814) );
  AND2_X1 U12599 ( .A1(n10063), .A2(n9809), .ZN(n9815) );
  AND2_X1 U12600 ( .A1(n9760), .A2(n10012), .ZN(n9816) );
  AND2_X1 U12601 ( .A1(n9766), .A2(n10099), .ZN(n9817) );
  AND2_X1 U12602 ( .A1(n10159), .A2(n10915), .ZN(n9818) );
  INV_X1 U12603 ( .A(n14804), .ZN(n14808) );
  INV_X1 U12604 ( .A(n13100), .ZN(n20083) );
  INV_X1 U12605 ( .A(n13788), .ZN(n10247) );
  INV_X1 U12606 ( .A(n14808), .ZN(n14791) );
  INV_X1 U12607 ( .A(n11500), .ZN(n10179) );
  NAND2_X1 U12608 ( .A1(n12915), .A2(n12914), .ZN(n13029) );
  NOR2_X1 U12609 ( .A1(n16037), .A2(n16036), .ZN(n9819) );
  INV_X1 U12610 ( .A(n20149), .ZN(n20133) );
  NAND2_X1 U12611 ( .A1(n12915), .A2(n9767), .ZN(n13048) );
  NOR2_X1 U12612 ( .A1(n13225), .A2(n13224), .ZN(n13248) );
  NOR2_X1 U12613 ( .A1(n13349), .A2(n10257), .ZN(n13462) );
  NAND2_X1 U12614 ( .A1(n18884), .A2(n19002), .ZN(n14690) );
  INV_X1 U12615 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20773) );
  OR2_X1 U12616 ( .A1(n12224), .A2(n12223), .ZN(n9820) );
  NOR2_X1 U12617 ( .A1(n14680), .A2(n10222), .ZN(n9821) );
  OR3_X1 U12618 ( .A1(n13707), .A2(n13706), .A3(n14752), .ZN(n9822) );
  AND2_X1 U12619 ( .A1(n9821), .A2(n10221), .ZN(n9823) );
  NOR2_X1 U12620 ( .A1(n13239), .A2(n13228), .ZN(n13229) );
  NOR2_X1 U12621 ( .A1(n12060), .A2(n14927), .ZN(n12058) );
  OR2_X1 U12622 ( .A1(n19060), .A2(n13896), .ZN(n9824) );
  OR2_X1 U12623 ( .A1(n10102), .A2(n10927), .ZN(n9825) );
  AND2_X1 U12624 ( .A1(n10212), .A2(n12570), .ZN(n9826) );
  AND2_X1 U12625 ( .A1(n10088), .A2(n14728), .ZN(n9827) );
  AND2_X1 U12626 ( .A1(n12915), .A2(n10250), .ZN(n13049) );
  NOR2_X1 U12627 ( .A1(n12940), .A2(n10216), .ZN(n9828) );
  AND2_X1 U12628 ( .A1(n14105), .A2(n14192), .ZN(n9829) );
  INV_X1 U12629 ( .A(n14019), .ZN(n10069) );
  INV_X1 U12630 ( .A(n10202), .ZN(n13447) );
  OR2_X1 U12631 ( .A1(n13136), .A2(n13137), .ZN(n10202) );
  INV_X1 U12632 ( .A(n10001), .ZN(n12057) );
  NOR2_X1 U12633 ( .A1(n12055), .A2(n16078), .ZN(n10001) );
  NAND2_X1 U12634 ( .A1(n9911), .A2(n9912), .ZN(n13349) );
  OR2_X1 U12635 ( .A1(n17537), .A2(n17550), .ZN(n9830) );
  INV_X1 U12636 ( .A(n10019), .ZN(n10018) );
  NAND2_X1 U12637 ( .A1(n9755), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10019) );
  AND2_X1 U12638 ( .A1(n10199), .A2(n10207), .ZN(n9831) );
  AND2_X1 U12639 ( .A1(n9826), .A2(n15154), .ZN(n9832) );
  NOR2_X1 U12640 ( .A1(n13902), .A2(n10208), .ZN(n9833) );
  AND2_X1 U12641 ( .A1(n9980), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9834) );
  AND2_X1 U12642 ( .A1(n10112), .A2(n10109), .ZN(n9835) );
  AND2_X1 U12643 ( .A1(n9823), .A2(n10220), .ZN(n9836) );
  AND2_X1 U12644 ( .A1(n10004), .A2(n16815), .ZN(n9837) );
  AND2_X1 U12645 ( .A1(n10008), .A2(n17507), .ZN(n9838) );
  AND2_X1 U12646 ( .A1(n10018), .A2(n16544), .ZN(n9839) );
  AND2_X1 U12647 ( .A1(n9770), .A2(n12282), .ZN(n9840) );
  INV_X1 U12648 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n9983) );
  INV_X1 U12649 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9987) );
  INV_X1 U12650 ( .A(n17761), .ZN(n17598) );
  AND2_X1 U12651 ( .A1(n16528), .A2(n9755), .ZN(n9841) );
  NAND2_X1 U12652 ( .A1(n9729), .A2(n20189), .ZN(n12010) );
  INV_X1 U12653 ( .A(n12010), .ZN(n11926) );
  OR2_X1 U12654 ( .A1(n17218), .A2(n16937), .ZN(n9842) );
  OR2_X1 U12655 ( .A1(n16728), .A2(n16547), .ZN(n9843) );
  AND2_X1 U12656 ( .A1(n11133), .A2(n12388), .ZN(n9844) );
  INV_X1 U12657 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n9986) );
  INV_X1 U12658 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n9982) );
  NOR2_X1 U12659 ( .A1(n13495), .A2(n13494), .ZN(n9845) );
  AND2_X1 U12660 ( .A1(n9940), .A2(n9773), .ZN(n9846) );
  OR2_X1 U12661 ( .A1(n12519), .A2(n10037), .ZN(n9847) );
  INV_X1 U12662 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10114) );
  INV_X1 U12663 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10056) );
  INV_X1 U12664 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10020) );
  INV_X1 U12665 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10039) );
  INV_X1 U12666 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10038) );
  INV_X1 U12667 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10002) );
  INV_X1 U12668 ( .A(n14468), .ZN(n10053) );
  INV_X1 U12669 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10115) );
  INV_X1 U12670 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18787) );
  AOI22_X2 U12671 ( .A1(DATAI_18_), .A2(n20207), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n20208), .ZN(n20671) );
  AOI22_X2 U12672 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20208), .B1(DATAI_19_), 
        .B2(n20207), .ZN(n20678) );
  AOI22_X2 U12673 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20208), .B1(DATAI_21_), 
        .B2(n20207), .ZN(n20690) );
  NOR3_X2 U12674 ( .A1(n9722), .A2(n18527), .A3(n18452), .ZN(n18447) );
  NOR3_X2 U12675 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n9722), .A3(
        n18452), .ZN(n18420) );
  NOR3_X2 U12676 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n9722), .A3(
        n18332), .ZN(n18327) );
  NOR3_X2 U12677 ( .A1(n9722), .A2(n18527), .A3(n18526), .ZN(n18553) );
  AOI22_X2 U12678 ( .A1(DATAI_23_), .A2(n20207), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n20208), .ZN(n20706) );
  AOI22_X2 U12679 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20208), .B1(DATAI_22_), 
        .B2(n20207), .ZN(n20760) );
  NOR2_X2 U12680 ( .A1(n20161), .A2(n20160), .ZN(n20208) );
  NOR2_X2 U12681 ( .A1(n20159), .A2(n20161), .ZN(n20207) );
  NOR3_X2 U12682 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n9722), .A3(
        n18245), .ZN(n18241) );
  NOR2_X2 U12683 ( .A1(n12411), .A2(n11204), .ZN(n11136) );
  NOR2_X1 U12684 ( .A1(n9850), .A2(n9849), .ZN(n9848) );
  OR2_X2 U12685 ( .A1(n20285), .A2(n11163), .ZN(n20219) );
  NAND4_X1 U12686 ( .A1(n9868), .A2(n9870), .A3(n9856), .A4(n9854), .ZN(n13197) );
  NAND3_X1 U12687 ( .A1(n13126), .A2(n13125), .A3(n12448), .ZN(n9856) );
  NAND2_X1 U12689 ( .A1(n9858), .A2(n15923), .ZN(n14341) );
  NAND2_X1 U12690 ( .A1(n14371), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9858) );
  NAND4_X1 U12691 ( .A1(n9862), .A2(n15435), .A3(n15436), .A4(n9861), .ZN(
        n9860) );
  INV_X2 U12692 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18811) );
  NAND2_X1 U12693 ( .A1(n13125), .A2(n13126), .ZN(n13124) );
  NAND2_X1 U12694 ( .A1(n9869), .A2(n9789), .ZN(n9868) );
  INV_X1 U12695 ( .A(n13125), .ZN(n9869) );
  NAND2_X1 U12696 ( .A1(n13124), .A2(n12447), .ZN(n12453) );
  OAI21_X1 U12697 ( .B1(n14451), .B2(n15986), .A(n9878), .ZN(P1_U3000) );
  NAND3_X1 U12698 ( .A1(n9900), .A2(n9899), .A3(n9897), .ZN(n9896) );
  NAND3_X2 U12699 ( .A1(n15415), .A2(n15417), .A3(n15416), .ZN(n17263) );
  NOR2_X2 U12700 ( .A1(n18641), .A2(n18639), .ZN(n17947) );
  NAND2_X2 U12701 ( .A1(n12943), .A2(n12902), .ZN(n12915) );
  OAI21_X2 U12702 ( .B1(n14760), .B2(n9916), .A(n9915), .ZN(n13735) );
  XNOR2_X2 U12703 ( .A(n9918), .B(n10745), .ZN(n12889) );
  NAND2_X1 U12704 ( .A1(n10456), .A2(n10455), .ZN(n9918) );
  AOI21_X1 U12705 ( .B1(n10745), .B2(n9918), .A(n10744), .ZN(n12918) );
  NAND3_X1 U12706 ( .A1(n10504), .A2(n10505), .A3(n13832), .ZN(n10137) );
  NAND4_X1 U12707 ( .A1(n10270), .A2(n10539), .A3(n10271), .A4(n10538), .ZN(
        n10138) );
  AOI21_X2 U12708 ( .B1(n14925), .B2(n9964), .A(n12036), .ZN(n12039) );
  NAND2_X1 U12709 ( .A1(n9925), .A2(n9800), .ZN(n9972) );
  NAND2_X1 U12710 ( .A1(n10162), .A2(n9818), .ZN(n9925) );
  NAND2_X1 U12711 ( .A1(n10162), .A2(n10159), .ZN(n9930) );
  NAND2_X1 U12712 ( .A1(n9932), .A2(n9931), .ZN(n18119) );
  NAND2_X1 U12713 ( .A1(n17814), .A2(n17815), .ZN(n9931) );
  OR2_X1 U12714 ( .A1(n17814), .A2(n17815), .ZN(n9932) );
  INV_X1 U12715 ( .A(n17759), .ZN(n17693) );
  INV_X2 U12716 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18803) );
  XNOR2_X2 U12717 ( .A(n10658), .B(n9938), .ZN(n10659) );
  AND2_X2 U12718 ( .A1(n10146), .A2(n9940), .ZN(n14919) );
  NAND2_X2 U12719 ( .A1(n19212), .A2(n10411), .ZN(n12338) );
  NAND4_X1 U12720 ( .A1(n10361), .A2(n10358), .A3(n10359), .A4(n10360), .ZN(
        n9943) );
  NAND4_X1 U12721 ( .A1(n10365), .A2(n10362), .A3(n10363), .A4(n10364), .ZN(
        n9945) );
  NAND2_X1 U12722 ( .A1(n9947), .A2(n12956), .ZN(n9946) );
  NAND4_X1 U12723 ( .A1(n10373), .A2(n10370), .A3(n10371), .A4(n10372), .ZN(
        n9947) );
  NAND2_X1 U12724 ( .A1(n9949), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9948) );
  NAND4_X1 U12725 ( .A1(n10377), .A2(n10374), .A3(n10376), .A4(n10375), .ZN(
        n9949) );
  INV_X1 U12726 ( .A(n10658), .ZN(n10616) );
  NAND3_X1 U12727 ( .A1(n13443), .A2(n13439), .A3(n10889), .ZN(n9950) );
  NAND3_X1 U12728 ( .A1(n9954), .A2(n9953), .A3(n9951), .ZN(n15302) );
  AND2_X1 U12729 ( .A1(n15273), .A2(n9958), .ZN(n15217) );
  NAND2_X1 U12730 ( .A1(n15273), .A2(n9956), .ZN(n15221) );
  NAND2_X1 U12731 ( .A1(n15221), .A2(n9959), .ZN(n15225) );
  NOR2_X2 U12732 ( .A1(n9960), .A2(n10491), .ZN(n19325) );
  NOR2_X2 U12733 ( .A1(n9960), .A2(n10493), .ZN(n10589) );
  NOR2_X2 U12734 ( .A1(n10494), .A2(n9960), .ZN(n10590) );
  NOR2_X2 U12735 ( .A1(n10492), .A2(n9960), .ZN(n19291) );
  INV_X1 U12736 ( .A(n12889), .ZN(n9961) );
  NAND2_X1 U12737 ( .A1(n14925), .A2(n9963), .ZN(n9962) );
  NAND3_X1 U12738 ( .A1(n10138), .A2(n10137), .A3(n10136), .ZN(n10646) );
  AND2_X1 U12739 ( .A1(n10646), .A2(n10981), .ZN(n9967) );
  NAND2_X1 U12740 ( .A1(n9967), .A2(n9971), .ZN(n9966) );
  AOI21_X1 U12741 ( .B1(n9969), .B2(n9971), .A(n9968), .ZN(n13252) );
  NOR2_X1 U12742 ( .A1(n13851), .A2(n21153), .ZN(n9968) );
  AND2_X1 U12743 ( .A1(n10646), .A2(n9970), .ZN(n9969) );
  NAND2_X1 U12744 ( .A1(n9971), .A2(n10646), .ZN(n13257) );
  NAND2_X1 U12745 ( .A1(n9972), .A2(n9973), .ZN(n10983) );
  NAND2_X1 U12746 ( .A1(n10924), .A2(n9978), .ZN(n9977) );
  NAND2_X1 U12747 ( .A1(n12063), .A2(n9834), .ZN(n12060) );
  NAND2_X1 U12748 ( .A1(n12067), .A2(n9984), .ZN(n12086) );
  XNOR2_X1 U12749 ( .A(n9997), .B(n9996), .ZN(n12092) );
  INV_X1 U12750 ( .A(n16058), .ZN(n9996) );
  NOR2_X1 U12751 ( .A1(n14664), .A2(n9753), .ZN(n16065) );
  NAND2_X1 U12752 ( .A1(n12053), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10856) );
  NAND2_X1 U12753 ( .A1(n10003), .A2(n10004), .ZN(n16597) );
  INV_X1 U12754 ( .A(n10005), .ZN(n16609) );
  AOI21_X1 U12755 ( .B1(n16585), .B2(n17507), .A(n10010), .ZN(n10009) );
  NAND2_X1 U12756 ( .A1(n10007), .A2(n10006), .ZN(n16564) );
  NAND2_X1 U12757 ( .A1(n16585), .A2(n9838), .ZN(n10007) );
  NAND2_X1 U12758 ( .A1(n16528), .A2(n9839), .ZN(n10015) );
  NAND2_X1 U12759 ( .A1(n9757), .A2(n10021), .ZN(n16537) );
  NAND3_X1 U12760 ( .A1(n16543), .A2(n10030), .A3(n9812), .ZN(n10029) );
  NOR2_X1 U12761 ( .A1(n16554), .A2(n16852), .ZN(n16546) );
  INV_X2 U12762 ( .A(n11815), .ZN(n11794) );
  INV_X1 U12763 ( .A(n11116), .ZN(n10034) );
  INV_X1 U12764 ( .A(n11118), .ZN(n10036) );
  XNOR2_X2 U12765 ( .A(n11252), .B(n20322), .ZN(n12753) );
  NAND2_X1 U12766 ( .A1(n12620), .A2(n11134), .ZN(n10042) );
  NAND4_X1 U12767 ( .A1(n11133), .A2(n10047), .A3(n12388), .A4(n10042), .ZN(
        n11135) );
  INV_X1 U12768 ( .A(n10047), .ZN(n13001) );
  AND2_X2 U12769 ( .A1(n14323), .A2(n10048), .ZN(n14301) );
  INV_X1 U12770 ( .A(n10054), .ZN(n12522) );
  NAND3_X1 U12771 ( .A1(n11268), .A2(n10057), .A3(n11312), .ZN(n11374) );
  NAND3_X1 U12772 ( .A1(n11268), .A2(n11312), .A3(n11355), .ZN(n11368) );
  NAND2_X1 U12773 ( .A1(n10072), .A2(n9791), .ZN(n10071) );
  NAND2_X1 U12774 ( .A1(n10076), .A2(n10074), .ZN(n15893) );
  NAND2_X1 U12775 ( .A1(n10086), .A2(n10083), .ZN(P2_U2983) );
  NAND2_X1 U12776 ( .A1(n16057), .A2(n19156), .ZN(n10086) );
  AND2_X1 U12777 ( .A1(n14740), .A2(n9770), .ZN(n13573) );
  NAND2_X1 U12778 ( .A1(n14740), .A2(n9840), .ZN(n12281) );
  NAND2_X1 U12779 ( .A1(n14740), .A2(n9827), .ZN(n13572) );
  NAND2_X1 U12780 ( .A1(n14740), .A2(n14728), .ZN(n14730) );
  INV_X1 U12781 ( .A(n14788), .ZN(n10094) );
  NAND2_X1 U12782 ( .A1(n10943), .A2(n9817), .ZN(n10939) );
  NAND2_X1 U12783 ( .A1(n10891), .A2(n10107), .ZN(n10908) );
  AND2_X1 U12784 ( .A1(n10936), .A2(n10110), .ZN(n10948) );
  NAND2_X1 U12785 ( .A1(n10936), .A2(n10112), .ZN(n10950) );
  NAND2_X1 U12786 ( .A1(n10936), .A2(n9835), .ZN(n10977) );
  NAND2_X1 U12787 ( .A1(n10936), .A2(n10935), .ZN(n10952) );
  NOR2_X2 U12788 ( .A1(n10277), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10278) );
  NAND4_X1 U12789 ( .A1(n11131), .A2(n11204), .A3(n20209), .A4(n11328), .ZN(
        n11138) );
  NAND2_X1 U12790 ( .A1(n11132), .A2(n11136), .ZN(n12764) );
  NAND3_X1 U12791 ( .A1(n11132), .A2(n11136), .A3(n20166), .ZN(n12627) );
  INV_X1 U12792 ( .A(n12510), .ZN(n10127) );
  NAND2_X1 U12793 ( .A1(n11151), .A2(n10133), .ZN(n10132) );
  NAND2_X1 U12794 ( .A1(n10132), .A2(n11203), .ZN(n10128) );
  OAI211_X1 U12795 ( .C1(n10132), .C2(n10131), .A(n10135), .B(n10129), .ZN(
        n12442) );
  NAND2_X1 U12796 ( .A1(n11151), .A2(n11150), .ZN(n11332) );
  AND3_X1 U12797 ( .A1(n11027), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11024) );
  NAND2_X1 U12798 ( .A1(n10143), .A2(n10140), .ZN(n13274) );
  NAND2_X1 U12799 ( .A1(n13273), .A2(n13445), .ZN(n10144) );
  NAND2_X1 U12800 ( .A1(n10145), .A2(n10656), .ZN(n13273) );
  INV_X1 U12801 ( .A(n10656), .ZN(n10140) );
  NAND2_X1 U12802 ( .A1(n10143), .A2(n10142), .ZN(n10141) );
  NAND2_X1 U12803 ( .A1(n10656), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10142) );
  INV_X2 U12804 ( .A(n15142), .ZN(n10146) );
  OR2_X2 U12805 ( .A1(n15159), .A2(n10697), .ZN(n15142) );
  NAND2_X1 U12806 ( .A1(n14919), .A2(n9771), .ZN(n14900) );
  AND2_X1 U12807 ( .A1(n14919), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14905) );
  AND2_X2 U12808 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13150) );
  NAND2_X1 U12809 ( .A1(n10150), .A2(n10258), .ZN(n11022) );
  NAND3_X1 U12810 ( .A1(n14896), .A2(n14899), .A3(n10151), .ZN(n10150) );
  NAND2_X1 U12811 ( .A1(n10152), .A2(n14897), .ZN(n14890) );
  NAND4_X1 U12812 ( .A1(n10153), .A2(n10154), .A3(n13474), .A4(n11385), .ZN(
        n13475) );
  NAND2_X1 U12813 ( .A1(n11385), .A2(n11384), .ZN(n13409) );
  AOI21_X1 U12814 ( .B1(n12486), .B2(n11500), .A(n11311), .ZN(n13458) );
  INV_X1 U12815 ( .A(n11311), .ZN(n10156) );
  NAND3_X1 U12816 ( .A1(n10664), .A2(n10643), .A3(n10981), .ZN(n10157) );
  XNOR2_X1 U12817 ( .A(n10893), .B(n15354), .ZN(n15347) );
  NAND2_X1 U12818 ( .A1(n10895), .A2(n9763), .ZN(n10162) );
  CLKBUF_X1 U12819 ( .A(n10162), .Z(n10158) );
  NAND2_X1 U12820 ( .A1(n10895), .A2(n10894), .ZN(n15035) );
  OAI21_X1 U12821 ( .B1(n12426), .B2(n11315), .A(n10177), .ZN(n13121) );
  NOR2_X1 U12822 ( .A1(n13939), .A2(n13940), .ZN(n13923) );
  NOR3_X2 U12823 ( .A1(n13939), .A2(n13913), .A3(n10180), .ZN(n13912) );
  INV_X1 U12824 ( .A(n13529), .ZN(n10182) );
  NAND2_X1 U12825 ( .A1(n10182), .A2(n10183), .ZN(n14076) );
  INV_X1 U12826 ( .A(n15899), .ZN(n10187) );
  XNOR2_X1 U12827 ( .A(n12688), .B(n10188), .ZN(n19028) );
  INV_X1 U12828 ( .A(n12119), .ZN(n10189) );
  INV_X1 U12829 ( .A(n12120), .ZN(n10190) );
  NOR2_X1 U12830 ( .A1(n13018), .A2(n13017), .ZN(n13019) );
  NAND2_X1 U12831 ( .A1(n12120), .A2(n12119), .ZN(n10191) );
  NAND2_X1 U12832 ( .A1(n13136), .A2(n10193), .ZN(n10192) );
  NAND2_X1 U12833 ( .A1(n17836), .A2(n15738), .ZN(n10225) );
  INV_X1 U12834 ( .A(n10223), .ZN(n15740) );
  NAND2_X1 U12835 ( .A1(n17836), .A2(n9794), .ZN(n10223) );
  INV_X1 U12836 ( .A(n17823), .ZN(n10224) );
  NAND2_X1 U12837 ( .A1(n10225), .A2(n17823), .ZN(n17822) );
  NAND2_X1 U12838 ( .A1(n17772), .A2(n10235), .ZN(n17665) );
  AND2_X1 U12839 ( .A1(n15762), .A2(n18026), .ZN(n10239) );
  AND2_X4 U12840 ( .A1(n10510), .A2(n10277), .ZN(n13884) );
  AND2_X4 U12841 ( .A1(n12951), .A2(n10444), .ZN(n10518) );
  AND2_X2 U12842 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12951) );
  NAND2_X1 U12843 ( .A1(n14735), .A2(n9798), .ZN(n10248) );
  INV_X1 U12844 ( .A(n10243), .ZN(n10242) );
  NOR2_X1 U12845 ( .A1(n13899), .A2(n10102), .ZN(n14883) );
  INV_X1 U12846 ( .A(n12627), .ZN(n12620) );
  XNOR2_X1 U12847 ( .A(n12436), .B(n11317), .ZN(n11320) );
  NAND2_X1 U12848 ( .A1(n12442), .A2(n12441), .ZN(n12934) );
  INV_X1 U12849 ( .A(n12241), .ZN(n12225) );
  INV_X1 U12850 ( .A(n13264), .ZN(n11385) );
  INV_X1 U12851 ( .A(n13122), .ZN(n11340) );
  AND4_X1 U12852 ( .A1(n10503), .A2(n10502), .A3(n10501), .A4(n10500), .ZN(
        n10504) );
  INV_X1 U12853 ( .A(n12338), .ZN(n12313) );
  AOI22_X1 U12854 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10351) );
  AOI22_X1 U12855 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10340) );
  NAND2_X1 U12856 ( .A1(n10518), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10308) );
  NAND2_X1 U12857 ( .A1(n10518), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10276) );
  AOI22_X1 U12858 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10327) );
  NAND2_X1 U12859 ( .A1(n13976), .A2(n13978), .ZN(n13966) );
  NAND2_X1 U12860 ( .A1(n12889), .A2(n13322), .ZN(n10485) );
  INV_X1 U12861 ( .A(n14076), .ZN(n11508) );
  INV_X2 U12862 ( .A(n11815), .ZN(n11477) );
  NAND2_X1 U12863 ( .A1(n14743), .A2(n14746), .ZN(n14745) );
  NOR2_X1 U12864 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11338) );
  AND2_X1 U12865 ( .A1(n14888), .A2(n14897), .ZN(n10258) );
  AND2_X1 U12866 ( .A1(n10285), .A2(n10284), .ZN(n10259) );
  AND2_X1 U12867 ( .A1(n12537), .A2(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19205)
         );
  AND3_X1 U12868 ( .A1(n11249), .A2(n11248), .A3(n11247), .ZN(n10260) );
  AND2_X1 U12869 ( .A1(n11598), .A2(n11597), .ZN(n10261) );
  OR2_X1 U12870 ( .A1(n9753), .A2(n14973), .ZN(n10262) );
  OR2_X1 U12871 ( .A1(n14197), .A2(n12406), .ZN(n10263) );
  INV_X1 U12872 ( .A(n18773), .ZN(n18843) );
  AND3_X1 U12873 ( .A1(n20962), .A2(n16715), .A3(n16876), .ZN(n10264) );
  INV_X1 U12874 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10698) );
  AND2_X1 U12875 ( .A1(n18779), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18719) );
  OR3_X1 U12876 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17575), .ZN(n10265) );
  INV_X1 U12877 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n18855) );
  INV_X2 U12878 ( .A(n17216), .ZN(n17197) );
  NAND4_X1 U12879 ( .A1(n19234), .A2(n12851), .A3(n10860), .A4(n10399), .ZN(
        n10394) );
  NOR2_X1 U12880 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12682) );
  NAND2_X1 U12881 ( .A1(n10384), .A2(n12294), .ZN(n12675) );
  INV_X1 U12882 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15844) );
  INV_X2 U12883 ( .A(n13090), .ZN(n20104) );
  OR2_X1 U12884 ( .A1(n18334), .A2(n18528), .ZN(n18219) );
  CLKBUF_X1 U12885 ( .A(n16490), .Z(n16491) );
  NAND2_X1 U12886 ( .A1(n12882), .A2(n12588), .ZN(n18983) );
  OR2_X1 U12887 ( .A1(n12039), .A2(n12038), .ZN(n10266) );
  OR2_X1 U12888 ( .A1(n13585), .A2(n13584), .ZN(n10267) );
  AND2_X1 U12889 ( .A1(n15908), .A2(n13064), .ZN(n15906) );
  NAND2_X2 U12890 ( .A1(n13184), .A2(n13183), .ZN(n20040) );
  INV_X1 U12891 ( .A(n17563), .ZN(n17640) );
  OR3_X1 U12892 ( .A1(n15065), .A2(n15307), .A3(n10698), .ZN(n10268) );
  AND3_X1 U12893 ( .A1(n10385), .A2(n10414), .A3(n10384), .ZN(n10269) );
  INV_X1 U12894 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n21119) );
  AND3_X1 U12895 ( .A1(n10529), .A2(n10528), .A3(n10527), .ZN(n10270) );
  AND3_X1 U12896 ( .A1(n10532), .A2(n10531), .A3(n10530), .ZN(n10271) );
  AND4_X1 U12897 ( .A1(n11099), .A2(n11098), .A3(n11097), .A4(n11096), .ZN(
        n10272) );
  AND4_X1 U12898 ( .A1(n11075), .A2(n11074), .A3(n11073), .A4(n11072), .ZN(
        n10273) );
  NAND2_X1 U12899 ( .A1(n11091), .A2(n12970), .ZN(n10274) );
  INV_X1 U12900 ( .A(n11638), .ZN(n11825) );
  AND2_X1 U12901 ( .A1(n11868), .A2(n11867), .ZN(n11871) );
  NAND2_X1 U12902 ( .A1(n19635), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10535) );
  NAND2_X1 U12903 ( .A1(n10535), .A2(n13832), .ZN(n10536) );
  INV_X1 U12904 ( .A(n11876), .ZN(n11853) );
  NAND2_X1 U12905 ( .A1(n11767), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11036) );
  OR2_X1 U12906 ( .A1(n11290), .A2(n11289), .ZN(n12475) );
  NAND2_X1 U12907 ( .A1(n12686), .A2(n10413), .ZN(n10415) );
  INV_X1 U12908 ( .A(n13761), .ZN(n13762) );
  INV_X1 U12909 ( .A(n10714), .ZN(n10701) );
  NAND2_X1 U12910 ( .A1(n10518), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10288) );
  NAND2_X1 U12911 ( .A1(n11853), .A2(n11852), .ZN(n11877) );
  INV_X1 U12912 ( .A(n11265), .ZN(n11210) );
  OAI21_X1 U12913 ( .B1(n10416), .B2(n10415), .A(n12302), .ZN(n10417) );
  INV_X1 U12914 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10277) );
  NAND2_X1 U12915 ( .A1(n13760), .A2(n13762), .ZN(n13763) );
  NAND2_X1 U12916 ( .A1(n10525), .A2(n16316), .ZN(n10526) );
  AOI21_X1 U12917 ( .B1(n12312), .B2(n10701), .A(n10700), .ZN(n10706) );
  AOI22_X1 U12918 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10346) );
  INV_X1 U12919 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n21030) );
  NAND2_X1 U12920 ( .A1(n11280), .A2(n11279), .ZN(n11355) );
  OR2_X1 U12921 ( .A1(n11303), .A2(n11302), .ZN(n12488) );
  AOI21_X1 U12922 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20565), .A(
        n11888), .ZN(n11894) );
  AOI22_X1 U12923 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11092) );
  AND2_X1 U12924 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15844), .ZN(
        n10710) );
  INV_X1 U12925 ( .A(n14786), .ZN(n13606) );
  AND4_X1 U12926 ( .A1(n10680), .A2(n10679), .A3(n10678), .A4(n10677), .ZN(
        n10681) );
  INV_X1 U12927 ( .A(n10407), .ZN(n10403) );
  AND3_X1 U12928 ( .A1(n10276), .A2(n10275), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10283) );
  OAI21_X1 U12929 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18811), .A(
        n15469), .ZN(n15477) );
  INV_X1 U12930 ( .A(n12002), .ZN(n11959) );
  INV_X1 U12931 ( .A(n13991), .ZN(n11696) );
  INV_X1 U12932 ( .A(n13411), .ZN(n11384) );
  INV_X1 U12933 ( .A(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11123) );
  INV_X1 U12934 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n13994) );
  INV_X1 U12935 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11400) );
  INV_X1 U12936 ( .A(n11333), .ZN(n11689) );
  NAND2_X1 U12937 ( .A1(n13123), .A2(n11342), .ZN(n13198) );
  INV_X1 U12938 ( .A(n11155), .ZN(n11328) );
  NOR2_X1 U12939 ( .A1(n11034), .A2(n11033), .ZN(n11052) );
  INV_X1 U12940 ( .A(n11898), .ZN(n11889) );
  INV_X1 U12942 ( .A(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n20976) );
  OR2_X1 U12943 ( .A1(n10711), .A2(n10710), .ZN(n10713) );
  INV_X1 U12944 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10855) );
  INV_X1 U12945 ( .A(n13734), .ZN(n13731) );
  INV_X1 U12946 ( .A(n13351), .ZN(n13350) );
  NAND2_X1 U12947 ( .A1(n10343), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10344) );
  AND2_X1 U12948 ( .A1(n10822), .A2(n10821), .ZN(n14753) );
  AND2_X1 U12949 ( .A1(n16294), .A2(n13832), .ZN(n19072) );
  INV_X1 U12950 ( .A(n10485), .ZN(n10496) );
  NOR2_X1 U12951 ( .A1(n16884), .A2(n15389), .ZN(n15648) );
  NAND2_X1 U12952 ( .A1(n13179), .A2(n13909), .ZN(n12002) );
  INV_X1 U12953 ( .A(n13186), .ZN(n11935) );
  OR2_X1 U12954 ( .A1(n11918), .A2(n11917), .ZN(n11920) );
  OR2_X1 U12955 ( .A1(n11692), .A2(n13994), .ZN(n11720) );
  NAND2_X1 U12956 ( .A1(n9743), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11842) );
  AND2_X1 U12957 ( .A1(n11562), .A2(n11561), .ZN(n14173) );
  OR2_X1 U12958 ( .A1(n11401), .A2(n11400), .ZN(n11426) );
  OAI211_X1 U12959 ( .C1(n11889), .C2(n11207), .A(n11206), .B(n11205), .ZN(
        n11327) );
  OAI21_X1 U12960 ( .B1(n20859), .B2(n16047), .A(n14661), .ZN(n20165) );
  NAND2_X1 U12961 ( .A1(n10713), .A2(n10712), .ZN(n12328) );
  INV_X1 U12962 ( .A(n15153), .ZN(n12571) );
  AND2_X1 U12963 ( .A1(n10798), .A2(n10797), .ZN(n14797) );
  OR2_X1 U12964 ( .A1(n13834), .A2(n13833), .ZN(n13835) );
  OR2_X1 U12965 ( .A1(n13785), .A2(n13784), .ZN(n13787) );
  OAI21_X1 U12966 ( .B1(n12040), .B2(n11008), .A(n11007), .ZN(n11009) );
  AND2_X1 U12967 ( .A1(n15180), .A2(n10696), .ZN(n12372) );
  INV_X1 U12968 ( .A(n13322), .ZN(n19169) );
  OR2_X1 U12969 ( .A1(n19077), .A2(n12328), .ZN(n12329) );
  AND2_X1 U12970 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12839), .ZN(
        n12883) );
  AOI21_X1 U12971 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18665), .A(
        n15475), .ZN(n15579) );
  INV_X1 U12972 ( .A(n17976), .ZN(n15760) );
  AOI21_X1 U12973 ( .B1(n15574), .B2(n15573), .A(n15572), .ZN(n15599) );
  NAND2_X1 U12974 ( .A1(n18206), .A2(n18215), .ZN(n15564) );
  OR3_X1 U12975 ( .A1(n13955), .A2(n13959), .A3(n14316), .ZN(n13929) );
  OR2_X1 U12976 ( .A1(n14025), .A2(n12018), .ZN(n13997) );
  NOR2_X1 U12977 ( .A1(n11592), .A2(n14399), .ZN(n11593) );
  INV_X1 U12978 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14111) );
  INV_X1 U12979 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13521) );
  AND2_X1 U12980 ( .A1(n13364), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13365) );
  INV_X1 U12981 ( .A(n20021), .ZN(n20009) );
  NOR2_X1 U12982 ( .A1(n12014), .A2(n9731), .ZN(n12023) );
  AND2_X1 U12983 ( .A1(n11955), .A2(n11954), .ZN(n13517) );
  INV_X1 U12984 ( .A(n14198), .ZN(n14276) );
  AOI22_X1 U12985 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11130) );
  INV_X1 U12986 ( .A(n13990), .ZN(n14005) );
  INV_X1 U12987 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n14083) );
  OR2_X1 U12988 ( .A1(n10179), .A2(n11440), .ZN(n15899) );
  INV_X1 U12989 ( .A(n13212), .ZN(n13266) );
  AND2_X1 U12990 ( .A1(n12414), .A2(n12757), .ZN(n12790) );
  NOR2_X1 U12991 ( .A1(n13005), .A2(n12994), .ZN(n14557) );
  OR3_X1 U12992 ( .A1(n12798), .A2(n12797), .A3(n12796), .ZN(n15790) );
  INV_X1 U12993 ( .A(n11344), .ZN(n13404) );
  OR2_X1 U12994 ( .A1(n20247), .A2(n12437), .ZN(n20610) );
  OR2_X1 U12995 ( .A1(n20162), .A2(n13405), .ZN(n20536) );
  INV_X1 U12996 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20602) );
  NAND2_X1 U12997 ( .A1(n20772), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15820) );
  NAND2_X1 U12998 ( .A1(n12328), .A2(n10715), .ZN(n16291) );
  AND2_X1 U12999 ( .A1(n10842), .A2(n10841), .ZN(n13571) );
  NAND2_X1 U13000 ( .A1(n12938), .A2(n12939), .ZN(n12940) );
  NAND2_X1 U13001 ( .A1(n12679), .A2(n12678), .ZN(n12680) );
  OR2_X1 U13002 ( .A1(n12633), .A2(n9740), .ZN(n19073) );
  NAND2_X1 U13003 ( .A1(n12073), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12070) );
  INV_X1 U13004 ( .A(n11009), .ZN(n11010) );
  AND2_X1 U13005 ( .A1(n10793), .A2(n10792), .ZN(n14807) );
  INV_X1 U13006 ( .A(n16243), .ZN(n16226) );
  NOR2_X1 U13007 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12588) );
  INV_X1 U13008 ( .A(n19155), .ZN(n19035) );
  OR2_X1 U13009 ( .A1(n10719), .A2(n16323), .ZN(n15840) );
  NAND2_X1 U13010 ( .A1(n12330), .A2(n12329), .ZN(n16294) );
  INV_X1 U13011 ( .A(n12682), .ZN(n19679) );
  OR3_X1 U13012 ( .A1(n19442), .A2(n19476), .A3(n19441), .ZN(n19446) );
  NAND2_X1 U13013 ( .A1(n19909), .A2(n19920), .ZN(n19572) );
  INV_X1 U13014 ( .A(n19246), .ZN(n19253) );
  OR2_X1 U13015 ( .A1(n19750), .A2(n19744), .ZN(n19806) );
  OAI21_X1 U13016 ( .B1(n15581), .B2(n15580), .A(n15579), .ZN(n18654) );
  NOR2_X1 U13017 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16734), .ZN(n16719) );
  NOR2_X1 U13018 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16829), .ZN(n16811) );
  OR2_X1 U13019 ( .A1(n18846), .A2(n18183), .ZN(n16525) );
  INV_X1 U13020 ( .A(n16876), .ZN(n16894) );
  AOI211_X1 U13021 ( .C1(n17156), .C2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n15414), .B(n15413), .ZN(n15415) );
  NOR3_X1 U13022 ( .A1(n15468), .A2(n15611), .A3(n18621), .ZN(n15602) );
  NOR2_X1 U13023 ( .A1(n17494), .A2(n17493), .ZN(n17492) );
  NOR2_X1 U13024 ( .A1(n17998), .A2(n17552), .ZN(n17898) );
  INV_X1 U13025 ( .A(n16406), .ZN(n16409) );
  NAND2_X1 U13026 ( .A1(n15766), .A2(n10265), .ZN(n15767) );
  INV_X1 U13027 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17699) );
  INV_X1 U13028 ( .A(n15743), .ZN(n15744) );
  INV_X1 U13029 ( .A(n18186), .ZN(n18425) );
  NOR2_X1 U13030 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20859) );
  NAND2_X1 U13031 ( .A1(n11593), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11631) );
  NAND2_X1 U13032 ( .A1(n11560), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11592) );
  AND2_X1 U13033 ( .A1(n19982), .A2(n11921), .ZN(n19980) );
  AND2_X1 U13034 ( .A1(n19982), .A2(n13365), .ZN(n20027) );
  INV_X1 U13035 ( .A(n14196), .ZN(n20036) );
  BUF_X1 U13036 ( .A(n13966), .Z(n13977) );
  INV_X1 U13037 ( .A(n12405), .ZN(n13069) );
  INV_X1 U13038 ( .A(n13100), .ZN(n20101) );
  INV_X1 U13039 ( .A(n13091), .ZN(n20093) );
  INV_X1 U13040 ( .A(n15870), .ZN(n15915) );
  NAND2_X1 U13041 ( .A1(n11442), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11471) );
  AND2_X1 U13042 ( .A1(n13266), .A2(n13215), .ZN(n20116) );
  INV_X1 U13043 ( .A(n19955), .ZN(n20118) );
  NAND2_X1 U13044 ( .A1(n14657), .A2(n20773), .ZN(n12416) );
  INV_X1 U13045 ( .A(n20147), .ZN(n14618) );
  INV_X1 U13046 ( .A(n15986), .ZN(n20152) );
  INV_X1 U13047 ( .A(n15823), .ZN(n14661) );
  OAI22_X1 U13048 ( .A1(n20177), .A2(n20176), .B1(n20444), .B2(n20324), .ZN(
        n20215) );
  INV_X1 U13049 ( .A(n20230), .ZN(n20243) );
  OAI22_X1 U13050 ( .A1(n20254), .A2(n20253), .B1(n20383), .B2(n20444), .ZN(
        n20278) );
  AND2_X1 U13051 ( .A1(n20163), .A2(n20162), .ZN(n20289) );
  INV_X1 U13052 ( .A(n20412), .ZN(n20373) );
  OAI22_X1 U13053 ( .A1(n20385), .A2(n20384), .B1(n20563), .B2(n20383), .ZN(
        n20408) );
  INV_X1 U13054 ( .A(n20610), .ZN(n20350) );
  AND2_X1 U13055 ( .A1(n13405), .A2(n13404), .ZN(n20420) );
  NOR2_X1 U13056 ( .A1(n20247), .A2(n20164), .ZN(n20557) );
  NOR2_X2 U13057 ( .A1(n20536), .A2(n20610), .ZN(n21200) );
  AND2_X1 U13058 ( .A1(n20247), .A2(n12437), .ZN(n20637) );
  NOR2_X2 U13059 ( .A1(n20536), .A2(n20535), .ZN(n20597) );
  INV_X1 U13060 ( .A(n20327), .ZN(n20213) );
  INV_X1 U13061 ( .A(n20650), .ZN(n20702) );
  INV_X1 U13062 ( .A(n20660), .ZN(n20723) );
  INV_X1 U13063 ( .A(n20679), .ZN(n20741) );
  OAI211_X1 U13064 ( .C1(n20718), .C2(n20717), .A(n20716), .B(n20715), .ZN(
        n20767) );
  NAND2_X1 U13065 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20856) );
  INV_X1 U13066 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20794) );
  INV_X1 U13067 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20786) );
  INV_X1 U13068 ( .A(n20835), .ZN(n20829) );
  AND2_X1 U13069 ( .A1(n18853), .A2(n12272), .ZN(n19025) );
  OR2_X1 U13070 ( .A1(n14891), .A2(n19034), .ZN(n12287) );
  NAND2_X1 U13071 ( .A1(n14690), .A2(n10262), .ZN(n12564) );
  INV_X1 U13072 ( .A(n19026), .ZN(n19012) );
  INV_X1 U13073 ( .A(n19025), .ZN(n19010) );
  NAND2_X1 U13074 ( .A1(n12849), .A2(n12949), .ZN(n12850) );
  CLKBUF_X1 U13075 ( .A(n13111), .Z(n13109) );
  INV_X1 U13076 ( .A(n10414), .ZN(n12851) );
  NOR2_X1 U13077 ( .A1(n13899), .A2(n13898), .ZN(n19046) );
  INV_X1 U13078 ( .A(n16132), .ZN(n19055) );
  NOR2_X1 U13079 ( .A1(n12748), .A2(n12634), .ZN(n12693) );
  AND2_X1 U13080 ( .A1(n16225), .A2(n19153), .ZN(n16217) );
  OR2_X1 U13081 ( .A1(n14908), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15087) );
  AND2_X1 U13082 ( .A1(n18974), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16196) );
  INV_X1 U13083 ( .A(n16251), .ZN(n19187) );
  INV_X1 U13084 ( .A(n19682), .ZN(n19753) );
  AND2_X1 U13085 ( .A1(n16294), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16327) );
  INV_X1 U13086 ( .A(n19289), .ZN(n19281) );
  NOR2_X1 U13087 ( .A1(n19506), .A2(n19450), .ZN(n19293) );
  NOR2_X1 U13088 ( .A1(n19450), .A2(n19572), .ZN(n19375) );
  NOR2_X1 U13089 ( .A1(n19413), .A2(n19640), .ZN(n19398) );
  NOR2_X1 U13090 ( .A1(n19450), .A2(n19640), .ZN(n19431) );
  AND2_X1 U13091 ( .A1(n19446), .A2(n19444), .ZN(n19466) );
  OAI21_X1 U13092 ( .B1(n19480), .B2(n19479), .A(n19478), .ZN(n19500) );
  INV_X1 U13093 ( .A(n19537), .ZN(n19530) );
  NOR2_X1 U13094 ( .A1(n19633), .A2(n19506), .ZN(n19542) );
  INV_X1 U13095 ( .A(n19759), .ZN(n19609) );
  NOR2_X1 U13096 ( .A1(n19633), .A2(n19572), .ZN(n19602) );
  AND2_X1 U13097 ( .A1(n19243), .A2(n19249), .ZN(n19727) );
  OAI22_X1 U13098 ( .A1(n19231), .A2(n19255), .B1(n19230), .B2(n19253), .ZN(
        n19716) );
  OAI22_X1 U13099 ( .A1(n19241), .A2(n19255), .B1(n19240), .B2(n19253), .ZN(
        n19797) );
  NAND2_X1 U13100 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n15841) );
  INV_X1 U13101 ( .A(n16328), .ZN(n19834) );
  INV_X1 U13102 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19842) );
  NAND2_X1 U13103 ( .A1(n18653), .A2(n17415), .ZN(n18846) );
  OR2_X1 U13104 ( .A1(n16569), .A2(P3_EBX_REG_29__SCAN_IN), .ZN(n16545) );
  NOR2_X1 U13105 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16623), .ZN(n16608) );
  NOR2_X1 U13106 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16664), .ZN(n16648) );
  NOR2_X1 U13107 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16687), .ZN(n16673) );
  NOR2_X1 U13108 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16757), .ZN(n16742) );
  INV_X1 U13109 ( .A(n16897), .ZN(n16768) );
  INV_X1 U13110 ( .A(n16893), .ZN(n16888) );
  NAND2_X1 U13111 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17193), .ZN(n17187) );
  NOR2_X1 U13112 ( .A1(n17440), .A2(n17244), .ZN(n17238) );
  NOR3_X1 U13113 ( .A1(n17298), .A2(n17264), .A3(n17221), .ZN(n17259) );
  NOR2_X1 U13114 ( .A1(n15446), .A2(n15445), .ZN(n18210) );
  NOR2_X1 U13115 ( .A1(n17483), .A2(n17307), .ZN(n17302) );
  INV_X1 U13116 ( .A(n17325), .ZN(n17362) );
  AND2_X1 U13117 ( .A1(n18642), .A2(n15850), .ZN(n17335) );
  INV_X1 U13118 ( .A(n18183), .ZN(n17377) );
  INV_X1 U13119 ( .A(n17709), .ZN(n17692) );
  NOR2_X1 U13120 ( .A1(n17860), .A2(n17342), .ZN(n17752) );
  OAI21_X1 U13121 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18829), .A(n16498), 
        .ZN(n17857) );
  INV_X1 U13122 ( .A(n17857), .ZN(n17843) );
  NAND2_X1 U13123 ( .A1(n17709), .A2(n17640), .ZN(n17850) );
  NOR2_X1 U13124 ( .A1(n9736), .A2(n17490), .ZN(n16411) );
  INV_X1 U13125 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17992) );
  NOR2_X1 U13126 ( .A1(n18162), .A2(n17342), .ZN(n18073) );
  OAI21_X1 U13127 ( .B1(n15614), .B2(n15613), .A(n18830), .ZN(n18170) );
  NAND2_X1 U13128 ( .A1(n16516), .A2(n18181), .ZN(n18334) );
  NOR2_X1 U13129 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18787), .ZN(
        n18815) );
  INV_X1 U13130 ( .A(n18558), .ZN(n18540) );
  INV_X1 U13131 ( .A(n18439), .ZN(n18584) );
  NOR2_X1 U13132 ( .A1(n16516), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n16517) );
  INV_X1 U13133 ( .A(n18685), .ZN(n18830) );
  INV_X1 U13134 ( .A(n18836), .ZN(n18707) );
  INV_X1 U13135 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18700) );
  NAND2_X1 U13136 ( .A1(n12404), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14221)
         );
  NOR2_X1 U13137 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12538), .ZN(n16484)
         );
  OR2_X1 U13138 ( .A1(n12805), .A2(n12627), .ZN(n12854) );
  NAND2_X1 U13139 ( .A1(n12854), .A2(n12605), .ZN(n20854) );
  INV_X1 U13140 ( .A(n20025), .ZN(n19978) );
  AND2_X1 U13141 ( .A1(n12407), .A2(n10263), .ZN(n12408) );
  INV_X1 U13142 ( .A(n20116), .ZN(n13218) );
  OR2_X1 U13143 ( .A1(n20077), .A2(n9731), .ZN(n20044) );
  OR2_X1 U13144 ( .A1(n12805), .A2(n12804), .ZN(n20077) );
  NOR2_X1 U13145 ( .A1(n12854), .A2(n12853), .ZN(n13100) );
  INV_X1 U13146 ( .A(n15866), .ZN(n14408) );
  INV_X1 U13147 ( .A(n15932), .ZN(n20122) );
  OR2_X1 U13148 ( .A1(n12805), .A2(n15802), .ZN(n19955) );
  OR2_X1 U13149 ( .A1(n13005), .A2(n13004), .ZN(n20149) );
  OR2_X1 U13150 ( .A1(n13005), .A2(n12986), .ZN(n15986) );
  AOI21_X1 U13151 ( .B1(n13168), .B2(n13167), .A(n20213), .ZN(n20158) );
  AND2_X1 U13152 ( .A1(n12860), .A2(n12800), .ZN(n14662) );
  NAND2_X1 U13153 ( .A1(n20289), .A2(n20557), .ZN(n20230) );
  NAND2_X1 U13154 ( .A1(n20289), .A2(n20350), .ZN(n20276) );
  NAND2_X1 U13155 ( .A1(n20289), .A2(n20637), .ZN(n20316) );
  NAND2_X1 U13156 ( .A1(n20289), .A2(n20419), .ZN(n20329) );
  NAND2_X1 U13157 ( .A1(n20420), .A2(n20557), .ZN(n20377) );
  NAND2_X1 U13158 ( .A1(n20420), .A2(n20350), .ZN(n20412) );
  NAND2_X1 U13159 ( .A1(n20420), .A2(n20637), .ZN(n20435) );
  NAND2_X1 U13160 ( .A1(n20488), .A2(n20557), .ZN(n21204) );
  AOI22_X1 U13161 ( .A1(n20494), .A2(n20499), .B1(n20491), .B2(n20642), .ZN(
        n20527) );
  NAND2_X1 U13162 ( .A1(n20488), .A2(n20637), .ZN(n20556) );
  AOI22_X1 U13163 ( .A1(n20571), .A2(n20568), .B1(n20643), .B2(n20564), .ZN(
        n20601) );
  OR2_X1 U13164 ( .A1(n20639), .A2(n20558), .ZN(n20636) );
  OR2_X1 U13165 ( .A1(n20639), .A2(n20638), .ZN(n20770) );
  INV_X1 U13166 ( .A(n20844), .ZN(n20777) );
  INV_X1 U13167 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20795) );
  AND2_X1 U13168 ( .A1(n20786), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20853) );
  INV_X1 U13169 ( .A(n20827), .ZN(n20831) );
  NAND2_X1 U13170 ( .A1(n16292), .A2(n12578), .ZN(n18853) );
  INV_X1 U13171 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19898) );
  AND2_X1 U13172 ( .A1(n12288), .A2(n12287), .ZN(n12289) );
  NAND2_X1 U13173 ( .A1(n12286), .A2(n12285), .ZN(n19034) );
  NAND2_X1 U13174 ( .A1(n19010), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19037) );
  INV_X1 U13175 ( .A(n19032), .ZN(n19018) );
  NAND2_X1 U13176 ( .A1(n12850), .A2(n19815), .ZN(n14804) );
  NAND2_X1 U13177 ( .A1(n12943), .A2(n12946), .ZN(n19266) );
  INV_X1 U13178 ( .A(n19046), .ZN(n19051) );
  NAND2_X1 U13179 ( .A1(n13901), .A2(n13900), .ZN(n19059) );
  INV_X1 U13180 ( .A(n19053), .ZN(n19060) );
  AND2_X1 U13181 ( .A1(n12651), .A2(n12650), .ZN(n19232) );
  NAND2_X1 U13182 ( .A1(n13901), .A2(n12104), .ZN(n19061) );
  INV_X1 U13183 ( .A(n19081), .ZN(n19105) );
  OR2_X1 U13184 ( .A1(n19131), .A2(n19139), .ZN(n19133) );
  INV_X1 U13185 ( .A(n19131), .ZN(n19141) );
  AND2_X1 U13186 ( .A1(n12048), .A2(n12047), .ZN(n12049) );
  INV_X1 U13187 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16195) );
  NAND2_X1 U13188 ( .A1(n12587), .A2(n10852), .ZN(n16225) );
  XNOR2_X1 U13189 ( .A(n10699), .B(n10698), .ZN(n15062) );
  INV_X1 U13190 ( .A(n19182), .ZN(n19190) );
  INV_X1 U13191 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21153) );
  AND2_X1 U13192 ( .A1(n19262), .A2(n19261), .ZN(n19289) );
  INV_X1 U13193 ( .A(n19293), .ZN(n19317) );
  AND2_X1 U13194 ( .A1(n19324), .A2(n19323), .ZN(n19352) );
  INV_X1 U13195 ( .A(n19375), .ZN(n19383) );
  INV_X1 U13196 ( .A(n19398), .ZN(n19410) );
  INV_X1 U13197 ( .A(n19431), .ZN(n19439) );
  INV_X1 U13198 ( .A(n19459), .ZN(n19470) );
  INV_X1 U13199 ( .A(n19471), .ZN(n19504) );
  OR2_X1 U13200 ( .A1(n19678), .A2(n19506), .ZN(n19537) );
  INV_X1 U13201 ( .A(n19542), .ZN(n19565) );
  INV_X1 U13202 ( .A(n19797), .ZN(n19626) );
  AND2_X1 U13203 ( .A1(n19686), .A2(n19685), .ZN(n19705) );
  OR2_X1 U13204 ( .A1(n19633), .A2(n19640), .ZN(n19739) );
  INV_X1 U13205 ( .A(n19716), .ZN(n19786) );
  OR2_X1 U13206 ( .A1(n19678), .A2(n19899), .ZN(n19813) );
  INV_X1 U13207 ( .A(n19822), .ZN(n16336) );
  INV_X1 U13208 ( .A(n19896), .ZN(n19823) );
  INV_X1 U13209 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18834) );
  NAND2_X1 U13210 ( .A1(n18830), .A2(n18666), .ZN(n16498) );
  NOR2_X1 U13211 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16603), .ZN(n16596) );
  INV_X1 U13212 ( .A(n16880), .ZN(n16868) );
  OR2_X1 U13213 ( .A1(n17264), .A2(n17291), .ZN(n17282) );
  NOR3_X1 U13214 ( .A1(n17339), .A2(n17464), .A3(n17340), .ZN(n17338) );
  NOR2_X1 U13215 ( .A1(n15644), .A2(n15643), .ZN(n17358) );
  INV_X1 U13216 ( .A(n17371), .ZN(n17340) );
  NAND2_X1 U13217 ( .A1(n17394), .A2(n17377), .ZN(n17393) );
  INV_X1 U13218 ( .A(n17394), .ZN(n17413) );
  INV_X1 U13219 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17970) );
  INV_X1 U13220 ( .A(n17752), .ZN(n17764) );
  INV_X1 U13221 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17821) );
  INV_X1 U13222 ( .A(n16353), .ZN(n17860) );
  NAND2_X1 U13223 ( .A1(n16412), .A2(n16411), .ZN(n16413) );
  INV_X1 U13224 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17964) );
  INV_X1 U13225 ( .A(n18073), .ZN(n18078) );
  INV_X1 U13226 ( .A(n18149), .ZN(n18155) );
  NAND2_X1 U13227 ( .A1(n18656), .A2(n18154), .ZN(n18162) );
  AOI211_X1 U13228 ( .C1(n18830), .C2(n18640), .A(n18182), .B(n15594), .ZN(
        n18819) );
  INV_X1 U13229 ( .A(n18346), .ZN(n18355) );
  INV_X1 U13230 ( .A(n18369), .ZN(n18378) );
  INV_X1 U13231 ( .A(n18417), .ZN(n18424) );
  INV_X1 U13232 ( .A(n18444), .ZN(n18451) );
  INV_X1 U13233 ( .A(n18579), .ZN(n18539) );
  INV_X1 U13234 ( .A(n18554), .ZN(n18543) );
  INV_X1 U13235 ( .A(n18506), .ZN(n18576) );
  INV_X1 U13236 ( .A(n18548), .ZN(n18609) );
  INV_X1 U13237 ( .A(n16853), .ZN(n18693) );
  INV_X1 U13238 ( .A(n18784), .ZN(n18697) );
  INV_X1 U13239 ( .A(n16518), .ZN(n18833) );
  INV_X1 U13240 ( .A(n18843), .ZN(n18779) );
  INV_X1 U13241 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19847) );
  OR4_X1 U13242 ( .A1(n12562), .A2(n12561), .A3(n12560), .A4(n12559), .ZN(
        P2_U2832) );
  AND2_X4 U13243 ( .A1(n12951), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13885) );
  NOR2_X4 U13244 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13856) );
  AND2_X4 U13245 ( .A1(n13856), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10513) );
  AND2_X4 U13246 ( .A1(n13856), .A2(n10444), .ZN(n10509) );
  AOI22_X1 U13247 ( .A1(n10513), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10509), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10282) );
  AOI22_X1 U13248 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10281) );
  AND2_X4 U13249 ( .A1(n10279), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10512) );
  AOI22_X1 U13250 ( .A1(n9737), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10512), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10280) );
  NAND4_X1 U13251 ( .A1(n10283), .A2(n10282), .A3(n10281), .A4(n10280), .ZN(
        n10293) );
  AOI22_X1 U13252 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10512), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10285) );
  AOI22_X1 U13253 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10284) );
  AOI22_X1 U13254 ( .A1(n10513), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10509), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10286) );
  INV_X1 U13255 ( .A(n10286), .ZN(n10290) );
  NAND3_X1 U13256 ( .A1(n10288), .A2(n12956), .A3(n10287), .ZN(n10289) );
  NOR2_X1 U13257 ( .A1(n10290), .A2(n10289), .ZN(n10291) );
  NAND2_X1 U13258 ( .A1(n10259), .A2(n10291), .ZN(n10292) );
  NAND2_X1 U13259 ( .A1(n10509), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10295) );
  AOI22_X1 U13260 ( .A1(n10513), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10512), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10298) );
  AOI22_X1 U13261 ( .A1(n10506), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U13262 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10296) );
  NAND4_X1 U13263 ( .A1(n10299), .A2(n10298), .A3(n10297), .A4(n10296), .ZN(
        n10300) );
  NAND2_X1 U13264 ( .A1(n10300), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10307) );
  AOI22_X1 U13265 ( .A1(n10513), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10512), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U13266 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10509), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10303) );
  AOI22_X1 U13267 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10302) );
  AOI22_X1 U13268 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10301) );
  NAND4_X1 U13269 ( .A1(n10304), .A2(n10303), .A3(n10302), .A4(n10301), .ZN(
        n10305) );
  NAND2_X1 U13270 ( .A1(n10305), .A2(n12956), .ZN(n10306) );
  AOI22_X1 U13271 ( .A1(n10506), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10512), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10312) );
  AOI22_X1 U13272 ( .A1(n10509), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10311) );
  AOI22_X1 U13273 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10513), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10310) );
  NAND4_X1 U13274 ( .A1(n10313), .A2(n10312), .A3(n10311), .A4(n10310), .ZN(
        n10320) );
  AOI22_X1 U13275 ( .A1(n10513), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10512), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10314) );
  AOI22_X1 U13276 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U13277 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10509), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10316) );
  AOI22_X1 U13278 ( .A1(n10506), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10315) );
  NAND4_X1 U13279 ( .A1(n10318), .A2(n10317), .A3(n10316), .A4(n10315), .ZN(
        n10319) );
  NAND2_X1 U13280 ( .A1(n10320), .A2(n10319), .ZN(n10384) );
  INV_X1 U13281 ( .A(n10384), .ZN(n10381) );
  AOI22_X1 U13282 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10324) );
  AOI22_X1 U13283 ( .A1(n10506), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10323) );
  AOI22_X1 U13284 ( .A1(n10513), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10512), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10322) );
  AOI22_X1 U13285 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10509), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10321) );
  NAND4_X1 U13286 ( .A1(n10324), .A2(n10323), .A3(n10322), .A4(n10321), .ZN(
        n10325) );
  NAND2_X1 U13287 ( .A1(n10325), .A2(n12956), .ZN(n10332) );
  AOI22_X1 U13288 ( .A1(n10513), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10512), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10328) );
  AOI22_X1 U13289 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10326) );
  NAND4_X1 U13290 ( .A1(n10329), .A2(n10328), .A3(n10327), .A4(n10326), .ZN(
        n10330) );
  NAND2_X1 U13291 ( .A1(n10330), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10331) );
  AND2_X2 U13292 ( .A1(n10381), .A2(n10414), .ZN(n12300) );
  AND2_X2 U13293 ( .A1(n10333), .A2(n12300), .ZN(n10368) );
  AOI22_X1 U13294 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10337) );
  AOI22_X1 U13295 ( .A1(n10506), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U13296 ( .A1(n10513), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10512), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10335) );
  AOI22_X1 U13297 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10509), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10334) );
  NAND4_X1 U13298 ( .A1(n10337), .A2(n10336), .A3(n10335), .A4(n10334), .ZN(
        n10338) );
  AOI22_X1 U13299 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10509), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10342) );
  AOI22_X1 U13300 ( .A1(n10513), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10512), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10341) );
  AOI22_X1 U13301 ( .A1(n9737), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10339) );
  NAND4_X1 U13302 ( .A1(n10342), .A2(n10341), .A3(n10340), .A4(n10339), .ZN(
        n10343) );
  AOI22_X1 U13303 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10509), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10349) );
  AOI22_X1 U13304 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10348) );
  AOI22_X1 U13305 ( .A1(n10513), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10512), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10347) );
  NAND4_X1 U13306 ( .A1(n10349), .A2(n10348), .A3(n10347), .A4(n10346), .ZN(
        n10350) );
  NAND2_X1 U13307 ( .A1(n10350), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10357) );
  AOI22_X1 U13308 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10509), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10354) );
  AOI22_X1 U13309 ( .A1(n10513), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10512), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10353) );
  AOI22_X1 U13310 ( .A1(n9737), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10352) );
  NAND4_X1 U13311 ( .A1(n10354), .A2(n10353), .A3(n10352), .A4(n10351), .ZN(
        n10355) );
  NAND2_X1 U13312 ( .A1(n10355), .A2(n12956), .ZN(n10356) );
  NAND2_X1 U13313 ( .A1(n10368), .A2(n10386), .ZN(n10720) );
  AOI22_X1 U13314 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10509), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10361) );
  AOI22_X1 U13315 ( .A1(n10513), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10512), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10360) );
  AOI22_X1 U13316 ( .A1(n10506), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10359) );
  AOI22_X1 U13317 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10358) );
  AOI22_X1 U13318 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10509), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10365) );
  AOI22_X1 U13319 ( .A1(n10513), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10512), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10364) );
  AOI22_X1 U13320 ( .A1(n10506), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10363) );
  AOI22_X1 U13321 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10362) );
  INV_X4 U13322 ( .A(n10411), .ZN(n16316) );
  NOR2_X1 U13323 ( .A1(n16316), .A2(n19223), .ZN(n10366) );
  NAND2_X1 U13324 ( .A1(n10720), .A2(n10366), .ZN(n10369) );
  NAND2_X1 U13325 ( .A1(n10860), .A2(n10378), .ZN(n10391) );
  INV_X1 U13326 ( .A(n10391), .ZN(n10367) );
  NAND2_X1 U13327 ( .A1(n10368), .A2(n10367), .ZN(n10402) );
  NAND2_X1 U13328 ( .A1(n10369), .A2(n10402), .ZN(n12365) );
  AOI22_X1 U13329 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10509), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10373) );
  AOI22_X1 U13330 ( .A1(n10513), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10512), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10372) );
  AOI22_X1 U13331 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10371) );
  AOI22_X1 U13332 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10370) );
  AOI22_X1 U13333 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10509), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10377) );
  AOI22_X1 U13334 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10376) );
  AOI22_X1 U13335 ( .A1(n10513), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10512), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10375) );
  AOI22_X1 U13336 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10374) );
  NAND2_X1 U13337 ( .A1(n12365), .A2(n19212), .ZN(n10380) );
  INV_X1 U13338 ( .A(n10399), .ZN(n10378) );
  NAND2_X2 U13339 ( .A1(n10378), .A2(n10865), .ZN(n12104) );
  NAND2_X1 U13340 ( .A1(n12343), .A2(n16300), .ZN(n10379) );
  NAND2_X1 U13341 ( .A1(n10380), .A2(n10379), .ZN(n10389) );
  NAND2_X1 U13342 ( .A1(n12104), .A2(n19227), .ZN(n10410) );
  AND2_X1 U13343 ( .A1(n10390), .A2(n12294), .ZN(n10383) );
  NAND2_X1 U13344 ( .A1(n19234), .A2(n12686), .ZN(n10382) );
  NAND4_X1 U13345 ( .A1(n10410), .A2(n10383), .A3(n10382), .A4(n19250), .ZN(
        n10388) );
  INV_X1 U13346 ( .A(n10390), .ZN(n10386) );
  INV_X2 U13347 ( .A(n10413), .ZN(n19234) );
  INV_X1 U13348 ( .A(n10400), .ZN(n10387) );
  NAND2_X1 U13349 ( .A1(n10389), .A2(n12347), .ZN(n10424) );
  INV_X1 U13350 ( .A(n10424), .ZN(n10398) );
  NAND2_X1 U13351 ( .A1(n10391), .A2(n10390), .ZN(n12297) );
  INV_X1 U13352 ( .A(n12297), .ZN(n10392) );
  NAND2_X1 U13353 ( .A1(n10392), .A2(n19234), .ZN(n12305) );
  NAND2_X1 U13354 ( .A1(n12104), .A2(n10413), .ZN(n12295) );
  NAND2_X1 U13355 ( .A1(n12305), .A2(n10393), .ZN(n12349) );
  NAND2_X1 U13356 ( .A1(n12349), .A2(n19227), .ZN(n10396) );
  INV_X2 U13357 ( .A(n10865), .ZN(n10860) );
  NAND2_X1 U13358 ( .A1(n10423), .A2(n12313), .ZN(n10397) );
  NAND2_X1 U13359 ( .A1(n10457), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10405) );
  INV_X1 U13360 ( .A(n12675), .ZN(n12344) );
  NAND4_X1 U13361 ( .A1(n12094), .A2(n12344), .A3(n16300), .A4(n19243), .ZN(
        n10401) );
  INV_X1 U13362 ( .A(n10402), .ZN(n12292) );
  NAND2_X1 U13363 ( .A1(n12292), .A2(n19212), .ZN(n10406) );
  NAND2_X2 U13364 ( .A1(n10405), .A2(n10404), .ZN(n10471) );
  INV_X1 U13365 ( .A(n10471), .ZN(n10441) );
  NOR2_X1 U13366 ( .A1(n10408), .A2(n10407), .ZN(n10419) );
  NAND2_X1 U13367 ( .A1(n10409), .A2(n10412), .ZN(n12674) );
  NAND2_X1 U13368 ( .A1(n12674), .A2(n12338), .ZN(n12340) );
  INV_X1 U13369 ( .A(n10411), .ZN(n10412) );
  NAND3_X1 U13370 ( .A1(n10412), .A2(n10860), .A3(n19250), .ZN(n10416) );
  AND2_X1 U13371 ( .A1(n10414), .A2(n10413), .ZN(n12356) );
  NAND2_X1 U13372 ( .A1(n12356), .A2(n19227), .ZN(n12302) );
  AOI21_X2 U13373 ( .B1(n10419), .B2(n12377), .A(n16324), .ZN(n10447) );
  NAND2_X1 U13374 ( .A1(n10447), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10429) );
  NAND2_X1 U13375 ( .A1(n12344), .A2(n12313), .ZN(n10430) );
  INV_X1 U13376 ( .A(n12588), .ZN(n10434) );
  NAND2_X1 U13377 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10420) );
  NAND2_X1 U13378 ( .A1(n10434), .A2(n10420), .ZN(n10421) );
  AOI21_X1 U13379 ( .B1(n10733), .B2(P2_EBX_REG_0__SCAN_IN), .A(n10421), .ZN(
        n10428) );
  NAND2_X1 U13380 ( .A1(n10765), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10427) );
  INV_X1 U13381 ( .A(n12343), .ZN(n10422) );
  OAI21_X1 U13382 ( .B1(n10425), .B2(n10424), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n10426) );
  NAND4_X1 U13383 ( .A1(n10429), .A2(n10428), .A3(n10427), .A4(n10426), .ZN(
        n10474) );
  INV_X1 U13384 ( .A(n10430), .ZN(n10432) );
  AND2_X1 U13385 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n10431) );
  OAI22_X1 U13386 ( .A1(n12377), .A2(n16324), .B1(n10434), .B2(n19933), .ZN(
        n10435) );
  INV_X1 U13387 ( .A(n10435), .ZN(n10436) );
  NAND2_X1 U13388 ( .A1(n10437), .A2(n10436), .ZN(n10475) );
  NAND2_X1 U13389 ( .A1(n10474), .A2(n10475), .ZN(n10473) );
  BUF_X1 U13390 ( .A(n10447), .Z(n10736) );
  NAND2_X1 U13391 ( .A1(n10736), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10440) );
  NAND2_X1 U13392 ( .A1(n10765), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10439) );
  AOI22_X1 U13393 ( .A1(n10733), .A2(P2_EBX_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10438) );
  NAND2_X1 U13394 ( .A1(n10441), .A2(n10473), .ZN(n10442) );
  NAND2_X1 U13395 ( .A1(n10457), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10446) );
  AOI21_X1 U13396 ( .B1(n16324), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10445) );
  NAND2_X1 U13397 ( .A1(n10446), .A2(n10445), .ZN(n10453) );
  INV_X1 U13398 ( .A(n10453), .ZN(n10451) );
  INV_X1 U13399 ( .A(n10447), .ZN(n10460) );
  AOI22_X1 U13400 ( .A1(n10733), .A2(P2_EBX_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10449) );
  NAND2_X1 U13401 ( .A1(n10765), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10448) );
  OAI211_X2 U13402 ( .C1(n10460), .C2(n19185), .A(n10449), .B(n10448), .ZN(
        n10452) );
  INV_X1 U13403 ( .A(n10452), .ZN(n10450) );
  NAND2_X1 U13404 ( .A1(n10451), .A2(n10450), .ZN(n10455) );
  NAND2_X1 U13405 ( .A1(n10453), .A2(n10452), .ZN(n10454) );
  AND2_X2 U13406 ( .A1(n10455), .A2(n10454), .ZN(n10468) );
  NAND2_X1 U13407 ( .A1(n10469), .A2(n10468), .ZN(n10456) );
  INV_X1 U13408 ( .A(n10457), .ZN(n10459) );
  NAND2_X1 U13409 ( .A1(n12588), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10458) );
  OAI21_X1 U13410 ( .B1(n10459), .B2(n12956), .A(n10458), .ZN(n10463) );
  AOI22_X1 U13411 ( .A1(n10733), .A2(P2_EBX_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10462) );
  NAND2_X1 U13412 ( .A1(n10765), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10461) );
  OAI211_X1 U13413 ( .C1(n10460), .C2(n21153), .A(n10462), .B(n10461), .ZN(
        n10464) );
  NAND2_X1 U13414 ( .A1(n10463), .A2(n10464), .ZN(n10467) );
  INV_X1 U13415 ( .A(n10463), .ZN(n10466) );
  INV_X1 U13416 ( .A(n10464), .ZN(n10465) );
  XNOR2_X2 U13417 ( .A(n10469), .B(n10468), .ZN(n12838) );
  OR2_X2 U13418 ( .A1(n12889), .A2(n13322), .ZN(n10484) );
  INV_X1 U13419 ( .A(n10470), .ZN(n10472) );
  XNOR2_X2 U13420 ( .A(n10472), .B(n10471), .ZN(n10482) );
  INV_X1 U13421 ( .A(n10474), .ZN(n10477) );
  INV_X1 U13422 ( .A(n10475), .ZN(n10476) );
  NAND2_X1 U13423 ( .A1(n10477), .A2(n10476), .ZN(n10478) );
  NAND2_X1 U13424 ( .A1(n10482), .A2(n19155), .ZN(n10493) );
  NOR2_X2 U13425 ( .A1(n10484), .A2(n10493), .ZN(n19384) );
  INV_X1 U13426 ( .A(n10482), .ZN(n10479) );
  AOI22_X1 U13427 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19384), .B1(
        n19442), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10490) );
  INV_X1 U13428 ( .A(n10480), .ZN(n10481) );
  XNOR2_X2 U13429 ( .A(n10482), .B(n10481), .ZN(n12833) );
  NOR2_X2 U13430 ( .A1(n10484), .A2(n10492), .ZN(n10595) );
  AND2_X2 U13431 ( .A1(n19169), .A2(n12947), .ZN(n10499) );
  INV_X1 U13432 ( .A(n10491), .ZN(n10483) );
  AND2_X2 U13433 ( .A1(n10499), .A2(n10483), .ZN(n19741) );
  AOI22_X1 U13434 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10595), .B1(
        n19741), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10489) );
  NOR2_X2 U13435 ( .A1(n10484), .A2(n10494), .ZN(n19357) );
  INV_X1 U13436 ( .A(n10494), .ZN(n10497) );
  AOI22_X1 U13437 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19357), .B1(
        n19477), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10488) );
  INV_X1 U13438 ( .A(n19568), .ZN(n10486) );
  AOI22_X1 U13439 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n9730), .B1(
        n10486), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13440 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19325), .B1(
        n10589), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10503) );
  INV_X1 U13441 ( .A(n10493), .ZN(n10495) );
  AND2_X2 U13442 ( .A1(n10499), .A2(n10495), .ZN(n19635) );
  AOI22_X1 U13443 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19291), .B1(
        n19635), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10502) );
  AOI22_X1 U13444 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10590), .B1(
        n19510), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10501) );
  AND2_X2 U13445 ( .A1(n10499), .A2(n10497), .ZN(n19600) );
  AND2_X2 U13446 ( .A1(n10499), .A2(n10498), .ZN(n19690) );
  AOI22_X1 U13447 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19600), .B1(
        n19690), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10500) );
  AOI22_X1 U13448 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12162), .B1(
        n10574), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10517) );
  AND2_X2 U13449 ( .A1(n13880), .A2(n12956), .ZN(n10575) );
  AOI22_X1 U13450 ( .A1(n10575), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n10546), .ZN(n10516) );
  AND2_X2 U13451 ( .A1(n9738), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10545) );
  AND2_X2 U13452 ( .A1(n13886), .A2(n12956), .ZN(n10540) );
  AOI22_X1 U13453 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__3__SCAN_IN), .B2(n10540), .ZN(n10515) );
  AND2_X2 U13454 ( .A1(n13886), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13622) );
  AOI22_X1 U13455 ( .A1(n9728), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13622), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10514) );
  NAND4_X1 U13456 ( .A1(n10517), .A2(n10516), .A3(n10515), .A4(n10514), .ZN(
        n10524) );
  AOI22_X1 U13457 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n13652), .B1(
        n13647), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10522) );
  AND2_X2 U13458 ( .A1(n13879), .A2(n12956), .ZN(n13639) );
  AOI22_X1 U13459 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10521) );
  AND2_X2 U13460 ( .A1(n13884), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10582) );
  AOI22_X1 U13461 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10581), .B1(
        n10582), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10520) );
  AOI22_X1 U13462 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n10607), .B1(
        n12959), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10519) );
  NAND4_X1 U13463 ( .A1(n10522), .A2(n10521), .A3(n10520), .A4(n10519), .ZN(
        n10523) );
  INV_X1 U13464 ( .A(n12126), .ZN(n10525) );
  AOI22_X1 U13465 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19291), .B1(
        n19510), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10529) );
  AOI22_X1 U13466 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10590), .B1(
        n19690), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10528) );
  AOI22_X1 U13467 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10589), .B1(
        n19600), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10527) );
  AOI22_X1 U13468 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19442), .B1(
        n10486), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10532) );
  AOI22_X1 U13469 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19384), .B1(
        n19741), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10531) );
  AOI22_X1 U13470 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19325), .B1(
        n19357), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10530) );
  INV_X1 U13471 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13690) );
  INV_X1 U13472 ( .A(n19477), .ZN(n19474) );
  INV_X1 U13473 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10533) );
  OAI22_X1 U13474 ( .A1(n13690), .A2(n19544), .B1(n19474), .B2(n10533), .ZN(
        n10534) );
  INV_X1 U13475 ( .A(n10534), .ZN(n10539) );
  INV_X1 U13476 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13691) );
  NOR2_X1 U13477 ( .A1(n10537), .A2(n10536), .ZN(n10538) );
  AOI22_X1 U13478 ( .A1(n13647), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13622), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10544) );
  AOI22_X1 U13479 ( .A1(n10607), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10540), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10543) );
  AOI22_X1 U13480 ( .A1(n9728), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12959), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10542) );
  AOI22_X1 U13481 ( .A1(n13652), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10541) );
  NAND4_X1 U13482 ( .A1(n10544), .A2(n10543), .A3(n10542), .A4(n10541), .ZN(
        n10552) );
  AOI22_X1 U13483 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10575), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10550) );
  AOI22_X1 U13484 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10549) );
  AOI22_X1 U13485 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10545), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10548) );
  AOI22_X1 U13486 ( .A1(n10582), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10547) );
  NAND4_X1 U13487 ( .A1(n10550), .A2(n10549), .A3(n10548), .A4(n10547), .ZN(
        n10551) );
  OR2_X1 U13488 ( .A1(n16267), .A2(n13832), .ZN(n10647) );
  AOI22_X1 U13489 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n13621), .B1(
        n13647), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10556) );
  AOI22_X1 U13490 ( .A1(n10582), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n10546), .ZN(n10555) );
  AOI22_X1 U13491 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10607), .B1(
        n12959), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10554) );
  AOI22_X1 U13492 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n13622), .ZN(n10553) );
  NAND4_X1 U13493 ( .A1(n10556), .A2(n10555), .A3(n10554), .A4(n10553), .ZN(
        n10562) );
  AOI22_X1 U13494 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10560) );
  AOI22_X1 U13495 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10575), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10559) );
  AOI22_X1 U13496 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10558) );
  AOI22_X1 U13497 ( .A1(n13652), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10540), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10557) );
  NAND4_X1 U13498 ( .A1(n10560), .A2(n10559), .A3(n10558), .A4(n10557), .ZN(
        n10561) );
  NOR2_X1 U13499 ( .A1(n10647), .A2(n12109), .ZN(n10651) );
  AOI22_X1 U13500 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10575), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10566) );
  AOI22_X1 U13501 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n13652), .B1(
        n13621), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10565) );
  AOI22_X1 U13502 ( .A1(n10540), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n10546), .ZN(n10564) );
  AOI22_X1 U13503 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_11__2__SCAN_IN), .B2(n13622), .ZN(n10563) );
  NAND4_X1 U13504 ( .A1(n10566), .A2(n10565), .A3(n10564), .A4(n10563), .ZN(
        n10572) );
  AOI22_X1 U13505 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13647), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10570) );
  AOI22_X1 U13506 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12959), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10569) );
  AOI22_X1 U13507 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10580), .B1(
        n10582), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U13508 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10581), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10567) );
  NAND4_X1 U13509 ( .A1(n10570), .A2(n10569), .A3(n10568), .A4(n10567), .ZN(
        n10571) );
  OR2_X1 U13510 ( .A1(n10651), .A2(n10723), .ZN(n10573) );
  AOI22_X1 U13511 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12162), .B1(
        n10574), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10579) );
  AOI22_X1 U13512 ( .A1(n13647), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n10546), .ZN(n10578) );
  AOI22_X1 U13513 ( .A1(n10575), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13622), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10577) );
  AOI22_X1 U13514 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__4__SCAN_IN), .B2(n10540), .ZN(n10576) );
  NAND4_X1 U13515 ( .A1(n10579), .A2(n10578), .A3(n10577), .A4(n10576), .ZN(
        n10588) );
  AOI22_X1 U13516 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13652), .B1(
        n9728), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10586) );
  AOI22_X1 U13517 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10585) );
  AOI22_X1 U13518 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10581), .B1(
        n12959), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10584) );
  AOI22_X1 U13519 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n10582), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10583) );
  NAND4_X1 U13520 ( .A1(n10586), .A2(n10585), .A3(n10584), .A4(n10583), .ZN(
        n10587) );
  AOI22_X1 U13521 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19325), .B1(
        n10589), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10594) );
  AOI22_X1 U13522 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19600), .B1(
        n19690), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10593) );
  AOI22_X1 U13523 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n10590), .B1(
        n19510), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10592) );
  AOI22_X1 U13524 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19291), .B1(
        n19635), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10591) );
  NAND4_X1 U13525 ( .A1(n10594), .A2(n10593), .A3(n10592), .A4(n10591), .ZN(
        n10602) );
  AOI22_X1 U13526 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19384), .B1(
        n19442), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10600) );
  AOI22_X1 U13527 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n10595), .B1(
        n19741), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10599) );
  AOI22_X1 U13528 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19357), .B1(
        n19477), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10598) );
  INV_X1 U13529 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13798) );
  INV_X1 U13530 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13801) );
  OAI22_X1 U13531 ( .A1(n13798), .A2(n19544), .B1(n19568), .B2(n13801), .ZN(
        n10596) );
  INV_X1 U13532 ( .A(n10596), .ZN(n10597) );
  NAND4_X1 U13533 ( .A1(n10600), .A2(n10599), .A3(n10598), .A4(n10597), .ZN(
        n10601) );
  AOI22_X1 U13534 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10575), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10606) );
  AOI22_X1 U13535 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9728), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10605) );
  AOI22_X1 U13536 ( .A1(n13647), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10604) );
  AOI22_X1 U13537 ( .A1(n13652), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10540), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10603) );
  NAND4_X1 U13538 ( .A1(n10606), .A2(n10605), .A3(n10604), .A4(n10603), .ZN(
        n10613) );
  AOI22_X1 U13539 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13622), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10611) );
  AOI22_X1 U13540 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12959), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10610) );
  AOI22_X1 U13541 ( .A1(n10580), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10582), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10609) );
  AOI22_X1 U13542 ( .A1(n10581), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10608) );
  NAND4_X1 U13543 ( .A1(n10611), .A2(n10610), .A3(n10609), .A4(n10608), .ZN(
        n10612) );
  NAND2_X1 U13544 ( .A1(n12097), .A2(n16316), .ZN(n10614) );
  NAND2_X1 U13545 ( .A1(n10616), .A2(n10657), .ZN(n10642) );
  INV_X1 U13546 ( .A(n10642), .ZN(n10641) );
  AOI22_X1 U13547 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19384), .B1(
        n19442), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10620) );
  AOI22_X1 U13548 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19357), .B1(
        n9730), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U13549 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19325), .B1(
        n19477), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10618) );
  AOI22_X1 U13550 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10590), .B1(
        n19510), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10617) );
  NAND4_X1 U13551 ( .A1(n10620), .A2(n10619), .A3(n10618), .A4(n10617), .ZN(
        n10626) );
  AOI22_X1 U13552 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10595), .B1(
        n19741), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10624) );
  AOI22_X1 U13553 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10589), .B1(
        n10486), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10623) );
  AOI22_X1 U13554 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19600), .B1(
        n19690), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10622) );
  AOI22_X1 U13555 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19291), .B1(
        n19635), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10621) );
  NAND4_X1 U13556 ( .A1(n10624), .A2(n10623), .A3(n10622), .A4(n10621), .ZN(
        n10625) );
  AOI22_X1 U13557 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12162), .B1(
        n10574), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10630) );
  AOI22_X1 U13558 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12959), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10629) );
  AOI22_X1 U13559 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10581), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10628) );
  AOI22_X1 U13560 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10582), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10627) );
  NAND4_X1 U13561 ( .A1(n10630), .A2(n10629), .A3(n10628), .A4(n10627), .ZN(
        n10636) );
  AOI22_X1 U13562 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n13652), .B1(
        n13647), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10634) );
  AOI22_X1 U13563 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10575), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10633) );
  AOI22_X1 U13564 ( .A1(n10540), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n10546), .ZN(n10632) );
  AOI22_X1 U13565 ( .A1(n9728), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13622), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10631) );
  NAND4_X1 U13566 ( .A1(n10634), .A2(n10633), .A3(n10632), .A4(n10631), .ZN(
        n10635) );
  INV_X1 U13567 ( .A(n12134), .ZN(n10637) );
  NAND2_X1 U13568 ( .A1(n10637), .A2(n16316), .ZN(n10638) );
  NAND2_X1 U13569 ( .A1(n10641), .A2(n10640), .ZN(n10664) );
  NAND2_X1 U13570 ( .A1(n10642), .A2(n10660), .ZN(n10643) );
  XNOR2_X1 U13571 ( .A(n10646), .B(n12129), .ZN(n10656) );
  NAND2_X1 U13572 ( .A1(n10647), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16269) );
  INV_X1 U13573 ( .A(n16269), .ZN(n10648) );
  XOR2_X1 U13574 ( .A(n16267), .B(n12109), .Z(n10649) );
  NAND2_X1 U13575 ( .A1(n10648), .A2(n10649), .ZN(n10650) );
  XOR2_X1 U13576 ( .A(n10649), .B(n10648), .Z(n12600) );
  NAND2_X1 U13577 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12600), .ZN(
        n12599) );
  NAND2_X1 U13578 ( .A1(n10650), .A2(n12599), .ZN(n10652) );
  XNOR2_X1 U13579 ( .A(n19185), .B(n10652), .ZN(n12609) );
  XNOR2_X1 U13580 ( .A(n10723), .B(n10651), .ZN(n12608) );
  NAND2_X1 U13581 ( .A1(n12609), .A2(n12608), .ZN(n12607) );
  NAND2_X1 U13582 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10652), .ZN(
        n10653) );
  NAND2_X1 U13583 ( .A1(n12607), .A2(n10653), .ZN(n10654) );
  XNOR2_X1 U13584 ( .A(n10654), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13256) );
  INV_X1 U13585 ( .A(n10654), .ZN(n10655) );
  INV_X1 U13586 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13445) );
  INV_X1 U13587 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13449) );
  NAND2_X1 U13588 ( .A1(n10659), .A2(n13449), .ZN(n13438) );
  NAND2_X1 U13589 ( .A1(n10859), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13439) );
  INV_X1 U13590 ( .A(n13439), .ZN(n13442) );
  NAND2_X1 U13591 ( .A1(n13442), .A2(n10660), .ZN(n10661) );
  NAND2_X1 U13592 ( .A1(n13443), .A2(n13439), .ZN(n10662) );
  NAND2_X1 U13593 ( .A1(n10662), .A2(n10889), .ZN(n10663) );
  NAND2_X1 U13594 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10668) );
  NAND2_X1 U13595 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10667) );
  NAND2_X1 U13596 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10666) );
  NAND2_X1 U13597 ( .A1(n12959), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10665) );
  NAND2_X1 U13598 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10672) );
  NAND2_X1 U13599 ( .A1(n13652), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10671) );
  NAND2_X1 U13600 ( .A1(n13647), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10670) );
  NAND2_X1 U13601 ( .A1(n10575), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10669) );
  NAND2_X1 U13602 ( .A1(n9728), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10676) );
  NAND2_X1 U13603 ( .A1(n10540), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10675) );
  NAND2_X1 U13604 ( .A1(n10546), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10674) );
  NAND2_X1 U13605 ( .A1(n13622), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10673) );
  NAND2_X1 U13606 ( .A1(n10580), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10680) );
  NAND2_X1 U13607 ( .A1(n10581), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10679) );
  NAND2_X1 U13608 ( .A1(n10582), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10678) );
  NAND2_X1 U13609 ( .A1(n10607), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10677) );
  AND4_X2 U13610 ( .A1(n10684), .A2(n10683), .A3(n10682), .A4(n10681), .ZN(
        n10981) );
  NAND2_X1 U13611 ( .A1(n10664), .A2(n10981), .ZN(n10686) );
  NAND2_X1 U13612 ( .A1(n10691), .A2(n10686), .ZN(n10687) );
  INV_X1 U13613 ( .A(n10687), .ZN(n10688) );
  NAND2_X1 U13614 ( .A1(n10689), .A2(n10688), .ZN(n10690) );
  XNOR2_X1 U13615 ( .A(n10691), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16204) );
  INV_X1 U13616 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16246) );
  AND2_X1 U13617 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15309) );
  AND2_X1 U13618 ( .A1(n15309), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15258) );
  NAND2_X1 U13619 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15259) );
  INV_X1 U13620 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15260) );
  NOR2_X1 U13621 ( .A1(n15259), .A2(n15260), .ZN(n10693) );
  NAND2_X1 U13622 ( .A1(n15258), .A2(n10693), .ZN(n15224) );
  NAND3_X1 U13623 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10694) );
  NOR2_X1 U13624 ( .A1(n15224), .A2(n10694), .ZN(n15207) );
  AND2_X1 U13625 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10695) );
  AND2_X1 U13626 ( .A1(n15207), .A2(n10695), .ZN(n15180) );
  AND2_X1 U13627 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10696) );
  AND2_X1 U13628 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15134) );
  INV_X1 U13629 ( .A(n15134), .ZN(n10697) );
  INV_X1 U13630 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15124) );
  INV_X1 U13631 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21137) );
  INV_X1 U13632 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15076) );
  NAND2_X1 U13633 ( .A1(n19933), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10714) );
  OAI21_X1 U13634 ( .B1(n19933), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n10714), .ZN(n12314) );
  INV_X1 U13635 ( .A(n12314), .ZN(n12311) );
  MUX2_X1 U13636 ( .A(n19924), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n12312) );
  NAND2_X1 U13637 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19915), .ZN(
        n10702) );
  NAND2_X1 U13638 ( .A1(n10706), .A2(n10702), .ZN(n10703) );
  NAND2_X1 U13639 ( .A1(n10444), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10704) );
  NAND2_X1 U13640 ( .A1(n10703), .A2(n10704), .ZN(n10708) );
  MUX2_X1 U13641 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n19908), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10707) );
  OAI22_X1 U13642 ( .A1(n10708), .A2(n10707), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n12956), .ZN(n10711) );
  OR3_X1 U13643 ( .A1(n10711), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n15844), .ZN(n12322) );
  INV_X1 U13644 ( .A(n12322), .ZN(n10709) );
  OAI21_X1 U13645 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n10444), .A(
        n10704), .ZN(n10705) );
  XNOR2_X1 U13646 ( .A(n10706), .B(n10705), .ZN(n12317) );
  XNOR2_X1 U13647 ( .A(n10708), .B(n10707), .ZN(n10725) );
  NOR3_X1 U13648 ( .A1(n10709), .A2(n12317), .A3(n10725), .ZN(n10716) );
  NAND2_X1 U13649 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n21098), .ZN(
        n10712) );
  XNOR2_X1 U13650 ( .A(n12312), .B(n10714), .ZN(n12310) );
  NAND2_X1 U13651 ( .A1(n12310), .A2(n10716), .ZN(n10715) );
  AOI211_X1 U13652 ( .C1(n12311), .C2(n10716), .A(P2_STATE2_REG_1__SCAN_IN), 
        .B(n16291), .ZN(n10719) );
  NAND2_X1 U13653 ( .A1(n10510), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10717) );
  NAND2_X1 U13654 ( .A1(n10717), .A2(n21098), .ZN(n16299) );
  INV_X1 U13655 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12668) );
  OAI21_X1 U13656 ( .B1(n10574), .B2(n16299), .A(n12668), .ZN(n10718) );
  AND2_X1 U13657 ( .A1(n10718), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16323) );
  NOR2_X1 U13658 ( .A1(n10721), .A2(n16316), .ZN(n10722) );
  NAND2_X1 U13659 ( .A1(n15840), .A2(n10722), .ZN(n10731) );
  MUX2_X1 U13660 ( .A(n16267), .B(n12314), .S(n12338), .Z(n10870) );
  INV_X1 U13661 ( .A(n12312), .ZN(n10724) );
  OAI21_X1 U13662 ( .B1(n10870), .B2(n10724), .A(n10862), .ZN(n10728) );
  MUX2_X1 U13663 ( .A(n12129), .B(n12322), .S(n12338), .Z(n10864) );
  INV_X1 U13664 ( .A(n10725), .ZN(n12320) );
  MUX2_X1 U13665 ( .A(n12126), .B(n12320), .S(n12338), .Z(n10863) );
  NAND2_X1 U13666 ( .A1(n10864), .A2(n10863), .ZN(n12308) );
  INV_X1 U13667 ( .A(n12308), .ZN(n10727) );
  INV_X1 U13668 ( .A(n12328), .ZN(n10726) );
  AOI21_X1 U13669 ( .B1(n10728), .B2(n10727), .A(n10726), .ZN(n19935) );
  AND2_X1 U13670 ( .A1(n16316), .A2(n19212), .ZN(n12298) );
  INV_X1 U13671 ( .A(n12298), .ZN(n10729) );
  NAND2_X1 U13672 ( .A1(n19935), .A2(n19937), .ZN(n10730) );
  NAND2_X1 U13673 ( .A1(n10731), .A2(n10730), .ZN(n12291) );
  NAND2_X1 U13674 ( .A1(n21119), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12270) );
  AND2_X1 U13675 ( .A1(n19212), .A2(n19815), .ZN(n10732) );
  AOI22_X1 U13676 ( .A1(n10847), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n10735) );
  NAND2_X1 U13677 ( .A1(n10765), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n10734) );
  AND2_X1 U13678 ( .A1(n10735), .A2(n10734), .ZN(n10738) );
  NAND2_X1 U13679 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10737) );
  NAND2_X1 U13680 ( .A1(n10738), .A2(n10737), .ZN(n13241) );
  AOI22_X1 U13681 ( .A1(n10847), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10740) );
  NAND2_X1 U13682 ( .A1(n10848), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n10739) );
  AND2_X1 U13683 ( .A1(n10740), .A2(n10739), .ZN(n10742) );
  NAND2_X1 U13684 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10741) );
  INV_X1 U13685 ( .A(n10743), .ZN(n10744) );
  AOI22_X1 U13686 ( .A1(n10847), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10747) );
  NAND2_X1 U13687 ( .A1(n10848), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n10746) );
  AND2_X1 U13688 ( .A1(n10747), .A2(n10746), .ZN(n10749) );
  NAND2_X1 U13689 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10748) );
  NAND2_X1 U13690 ( .A1(n10749), .A2(n10748), .ZN(n12917) );
  NAND2_X1 U13691 ( .A1(n12918), .A2(n12917), .ZN(n12919) );
  AOI22_X1 U13692 ( .A1(n10847), .A2(P2_EBX_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10751) );
  NAND2_X1 U13693 ( .A1(n10848), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n10750) );
  AND2_X1 U13694 ( .A1(n10751), .A2(n10750), .ZN(n10753) );
  NAND2_X1 U13695 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10752) );
  NOR2_X2 U13696 ( .A1(n12919), .A2(n12904), .ZN(n13042) );
  INV_X1 U13697 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15354) );
  AOI22_X1 U13698 ( .A1(n10847), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10755) );
  NAND2_X1 U13699 ( .A1(n10848), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n10754) );
  OAI211_X1 U13700 ( .C1(n10460), .C2(n15354), .A(n10755), .B(n10754), .ZN(
        n13043) );
  AOI22_X1 U13701 ( .A1(n10847), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10757) );
  NAND2_X1 U13702 ( .A1(n10765), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10756) );
  AND2_X1 U13703 ( .A1(n10757), .A2(n10756), .ZN(n10759) );
  NAND2_X1 U13704 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10758) );
  NAND2_X1 U13705 ( .A1(n10759), .A2(n10758), .ZN(n13047) );
  AOI22_X1 U13706 ( .A1(n10847), .A2(P2_EBX_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10761) );
  NAND2_X1 U13707 ( .A1(n10765), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n10760) );
  AND2_X1 U13708 ( .A1(n10761), .A2(n10760), .ZN(n10764) );
  NAND2_X1 U13709 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10763) );
  NAND2_X1 U13710 ( .A1(n13241), .A2(n13240), .ZN(n13239) );
  AOI22_X1 U13711 ( .A1(n10847), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n10767) );
  NAND2_X1 U13712 ( .A1(n10765), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n10766) );
  AND2_X1 U13713 ( .A1(n10767), .A2(n10766), .ZN(n10769) );
  NAND2_X1 U13714 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10768) );
  AOI22_X1 U13715 ( .A1(n10847), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n10771) );
  NAND2_X1 U13716 ( .A1(n10848), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n10770) );
  AND2_X1 U13717 ( .A1(n10771), .A2(n10770), .ZN(n10773) );
  NAND2_X1 U13718 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10772) );
  NAND2_X1 U13719 ( .A1(n10773), .A2(n10772), .ZN(n13247) );
  NAND2_X1 U13720 ( .A1(n13229), .A2(n13247), .ZN(n13347) );
  AOI22_X1 U13721 ( .A1(n10847), .A2(P2_EBX_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n10775) );
  NAND2_X1 U13722 ( .A1(n10848), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n10774) );
  AND2_X1 U13723 ( .A1(n10775), .A2(n10774), .ZN(n10777) );
  NAND2_X1 U13724 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10776) );
  AOI22_X1 U13725 ( .A1(n10847), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n10779) );
  NAND2_X1 U13726 ( .A1(n10848), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n10778) );
  AND2_X1 U13727 ( .A1(n10779), .A2(n10778), .ZN(n10781) );
  NAND2_X1 U13728 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10780) );
  AOI22_X1 U13729 ( .A1(n10847), .A2(P2_EBX_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n10783) );
  NAND2_X1 U13730 ( .A1(n10848), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n10782) );
  AND2_X1 U13731 ( .A1(n10783), .A2(n10782), .ZN(n10785) );
  NAND2_X1 U13732 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10784) );
  AOI22_X1 U13733 ( .A1(n10847), .A2(P2_EBX_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n10787) );
  NAND2_X1 U13734 ( .A1(n10848), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n10786) );
  AND2_X1 U13735 ( .A1(n10787), .A2(n10786), .ZN(n10789) );
  NAND2_X1 U13736 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10788) );
  NAND2_X1 U13737 ( .A1(n10789), .A2(n10788), .ZN(n13483) );
  AOI22_X1 U13738 ( .A1(n10847), .A2(P2_EBX_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n10791) );
  NAND2_X1 U13739 ( .A1(n10848), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n10790) );
  AND2_X1 U13740 ( .A1(n10791), .A2(n10790), .ZN(n10793) );
  NAND2_X1 U13741 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10792) );
  INV_X1 U13742 ( .A(n10794), .ZN(n14805) );
  AOI22_X1 U13743 ( .A1(n10847), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n10796) );
  NAND2_X1 U13744 ( .A1(n10848), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n10795) );
  AND2_X1 U13745 ( .A1(n10796), .A2(n10795), .ZN(n10798) );
  NAND2_X1 U13746 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10797) );
  AOI22_X1 U13747 ( .A1(n10847), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n10800) );
  NAND2_X1 U13748 ( .A1(n10848), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n10799) );
  AND2_X1 U13749 ( .A1(n10800), .A2(n10799), .ZN(n10802) );
  NAND2_X1 U13750 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10801) );
  NAND2_X1 U13751 ( .A1(n10802), .A2(n10801), .ZN(n14788) );
  AOI22_X1 U13752 ( .A1(n10847), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n10804) );
  NAND2_X1 U13753 ( .A1(n10848), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n10803) );
  AND2_X1 U13754 ( .A1(n10804), .A2(n10803), .ZN(n10806) );
  NAND2_X1 U13755 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10805) );
  NAND2_X1 U13756 ( .A1(n10806), .A2(n10805), .ZN(n14693) );
  AOI22_X1 U13757 ( .A1(n10847), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n10808) );
  NAND2_X1 U13758 ( .A1(n10848), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n10807) );
  AND2_X1 U13759 ( .A1(n10808), .A2(n10807), .ZN(n10810) );
  NAND2_X1 U13760 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10809) );
  AOI22_X1 U13761 ( .A1(n10847), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n10812) );
  NAND2_X1 U13762 ( .A1(n10848), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n10811) );
  AND2_X1 U13763 ( .A1(n10812), .A2(n10811), .ZN(n10814) );
  NAND2_X1 U13764 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10813) );
  AOI22_X1 U13765 ( .A1(n10847), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n10816) );
  NAND2_X1 U13766 ( .A1(n10848), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n10815) );
  AND2_X1 U13767 ( .A1(n10816), .A2(n10815), .ZN(n10818) );
  NAND2_X1 U13768 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10817) );
  NAND2_X1 U13769 ( .A1(n10818), .A2(n10817), .ZN(n12554) );
  NAND2_X1 U13770 ( .A1(n14767), .A2(n12554), .ZN(n14754) );
  AOI22_X1 U13771 ( .A1(n10847), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n10820) );
  NAND2_X1 U13772 ( .A1(n10848), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n10819) );
  AND2_X1 U13773 ( .A1(n10820), .A2(n10819), .ZN(n10822) );
  NAND2_X1 U13774 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10821) );
  AOI22_X1 U13775 ( .A1(n10847), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n10824) );
  NAND2_X1 U13776 ( .A1(n10848), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n10823) );
  AND2_X1 U13777 ( .A1(n10824), .A2(n10823), .ZN(n10826) );
  NAND2_X1 U13778 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10825) );
  AOI22_X1 U13779 ( .A1(n10847), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n10828) );
  NAND2_X1 U13780 ( .A1(n10848), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n10827) );
  AND2_X1 U13781 ( .A1(n10828), .A2(n10827), .ZN(n10830) );
  NAND2_X1 U13782 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10829) );
  AOI22_X1 U13783 ( .A1(n10847), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n10832) );
  NAND2_X1 U13784 ( .A1(n10848), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n10831) );
  AND2_X1 U13785 ( .A1(n10832), .A2(n10831), .ZN(n10834) );
  NAND2_X1 U13786 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10833) );
  NAND2_X1 U13787 ( .A1(n10834), .A2(n10833), .ZN(n14728) );
  AOI22_X1 U13788 ( .A1(n10847), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n10836) );
  NAND2_X1 U13789 ( .A1(n10848), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n10835) );
  AND2_X1 U13790 ( .A1(n10836), .A2(n10835), .ZN(n10838) );
  NAND2_X1 U13791 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10837) );
  AND2_X1 U13792 ( .A1(n10838), .A2(n10837), .ZN(n12043) );
  AOI22_X1 U13793 ( .A1(n10847), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n10840) );
  NAND2_X1 U13794 ( .A1(n10848), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n10839) );
  AND2_X1 U13795 ( .A1(n10840), .A2(n10839), .ZN(n10842) );
  NAND2_X1 U13796 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10841) );
  AOI22_X1 U13797 ( .A1(n10847), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n10844) );
  NAND2_X1 U13798 ( .A1(n10848), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n10843) );
  AND2_X1 U13799 ( .A1(n10844), .A2(n10843), .ZN(n10846) );
  NAND2_X1 U13800 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10845) );
  NAND2_X1 U13801 ( .A1(n10846), .A2(n10845), .ZN(n12282) );
  AOI22_X1 U13802 ( .A1(n10847), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n10850) );
  NAND2_X1 U13803 ( .A1(n10848), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n10849) );
  OAI211_X1 U13804 ( .C1(n10460), .C2(n10698), .A(n10850), .B(n10849), .ZN(
        n10851) );
  NAND2_X1 U13805 ( .A1(n21119), .A2(n19576), .ZN(n19900) );
  INV_X1 U13806 ( .A(n19900), .ZN(n19817) );
  OR2_X1 U13807 ( .A1(n12882), .A2(n19817), .ZN(n19925) );
  NAND2_X1 U13808 ( .A1(n19925), .A2(n16324), .ZN(n10852) );
  AND2_X1 U13809 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19916) );
  INV_X1 U13810 ( .A(n12888), .ZN(n10854) );
  NAND2_X1 U13811 ( .A1(n19898), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n10853) );
  NAND2_X1 U13812 ( .A1(n10854), .A2(n10853), .ZN(n19153) );
  NAND2_X1 U13813 ( .A1(n12078), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12076) );
  INV_X1 U13814 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16224) );
  NAND2_X1 U13815 ( .A1(n12077), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12074) );
  INV_X1 U13816 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15041) );
  NAND2_X1 U13817 ( .A1(n12075), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12072) );
  NAND2_X1 U13818 ( .A1(n12071), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12068) );
  NAND2_X1 U13819 ( .A1(n12069), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12066) );
  NOR2_X2 U13820 ( .A1(n12086), .A2(n14984), .ZN(n12088) );
  NAND2_X1 U13821 ( .A1(n12088), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12064) );
  NAND2_X1 U13822 ( .A1(n12058), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12055) );
  INV_X1 U13823 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16078) );
  INV_X1 U13824 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19888) );
  NOR2_X1 U13825 ( .A1(n16226), .A2(n19888), .ZN(n15053) );
  AOI21_X1 U13826 ( .B1(n19154), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15053), .ZN(n10857) );
  OAI21_X1 U13827 ( .B1(n19152), .B2(n12051), .A(n10857), .ZN(n10858) );
  OR2_X1 U13828 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(
        n10861) );
  BUF_X4 U13829 ( .A(n10860), .Z(n11016) );
  MUX2_X1 U13830 ( .A(n12109), .B(n10861), .S(n11016), .Z(n10875) );
  INV_X1 U13831 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13847) );
  MUX2_X1 U13832 ( .A(n10863), .B(n13847), .S(n11016), .Z(n10869) );
  INV_X1 U13833 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n21092) );
  MUX2_X1 U13834 ( .A(n10864), .B(n21092), .S(n11016), .Z(n10884) );
  MUX2_X1 U13835 ( .A(P2_EBX_REG_5__SCAN_IN), .B(n12097), .S(n10102), .Z(
        n10866) );
  AND2_X1 U13836 ( .A1(n10883), .A2(n10866), .ZN(n10867) );
  OR2_X1 U13837 ( .A1(n10867), .A2(n10891), .ZN(n18998) );
  INV_X1 U13838 ( .A(n10885), .ZN(n10868) );
  OAI21_X1 U13839 ( .B1(n10869), .B2(n10874), .A(n10868), .ZN(n13851) );
  INV_X1 U13840 ( .A(n10870), .ZN(n10871) );
  MUX2_X1 U13841 ( .A(n10871), .B(P2_EBX_REG_0__SCAN_IN), .S(n11016), .Z(
        n19031) );
  NAND2_X1 U13842 ( .A1(n19031), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16264) );
  NAND3_X1 U13843 ( .A1(n11016), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n10872) );
  NAND2_X1 U13844 ( .A1(n10875), .A2(n10872), .ZN(n19017) );
  NOR2_X1 U13845 ( .A1(n16264), .A2(n19017), .ZN(n10873) );
  NAND2_X1 U13846 ( .A1(n16264), .A2(n19017), .ZN(n12597) );
  OAI21_X1 U13847 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10873), .A(
        n12597), .ZN(n12613) );
  INV_X1 U13848 ( .A(n10874), .ZN(n10878) );
  NAND2_X1 U13849 ( .A1(n10876), .A2(n10875), .ZN(n10877) );
  NAND2_X1 U13850 ( .A1(n10878), .A2(n10877), .ZN(n13318) );
  XNOR2_X1 U13851 ( .A(n13318), .B(n19185), .ZN(n12612) );
  OR2_X1 U13852 ( .A1(n12613), .A2(n12612), .ZN(n12615) );
  INV_X1 U13853 ( .A(n13318), .ZN(n10879) );
  NAND2_X1 U13854 ( .A1(n10879), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10880) );
  NAND2_X1 U13855 ( .A1(n12615), .A2(n10880), .ZN(n13254) );
  INV_X1 U13856 ( .A(n13254), .ZN(n10881) );
  NAND2_X1 U13857 ( .A1(n13252), .A2(n10881), .ZN(n10882) );
  NAND2_X1 U13858 ( .A1(n9795), .A2(n21153), .ZN(n13253) );
  NAND2_X1 U13859 ( .A1(n10882), .A2(n13253), .ZN(n13278) );
  OAI21_X1 U13860 ( .B1(n10885), .B2(n10884), .A(n10883), .ZN(n13301) );
  XNOR2_X1 U13861 ( .A(n13301), .B(n13445), .ZN(n13276) );
  OAI22_X1 U13862 ( .A1(n13278), .A2(n13276), .B1(n13301), .B2(n13445), .ZN(
        n13436) );
  NAND2_X1 U13863 ( .A1(n13437), .A2(n13436), .ZN(n10888) );
  NAND2_X1 U13864 ( .A1(n10886), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10887) );
  INV_X1 U13865 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n18984) );
  MUX2_X1 U13866 ( .A(n12134), .B(n18984), .S(n11016), .Z(n10890) );
  OR2_X1 U13867 ( .A1(n10891), .A2(n10890), .ZN(n10892) );
  NAND2_X1 U13868 ( .A1(n10902), .A2(n10892), .ZN(n18985) );
  NAND2_X1 U13869 ( .A1(n15348), .A2(n15347), .ZN(n10895) );
  NAND2_X1 U13870 ( .A1(n10893), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10894) );
  MUX2_X1 U13871 ( .A(P2_EBX_REG_7__SCAN_IN), .B(n10981), .S(n10102), .Z(
        n10900) );
  INV_X1 U13872 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n10896) );
  NOR2_X1 U13873 ( .A1(n10102), .A2(n10896), .ZN(n10897) );
  AND2_X1 U13874 ( .A1(n10908), .A2(n10897), .ZN(n10898) );
  OR2_X1 U13875 ( .A1(n10907), .A2(n10898), .ZN(n13313) );
  OR2_X1 U13876 ( .A1(n10981), .A2(n16246), .ZN(n10899) );
  NOR2_X1 U13877 ( .A1(n13313), .A2(n10899), .ZN(n16198) );
  INV_X1 U13878 ( .A(n10900), .ZN(n10901) );
  XNOR2_X1 U13879 ( .A(n10902), .B(n10901), .ZN(n18974) );
  OAI21_X1 U13880 ( .B1(n13313), .B2(n10981), .A(n16246), .ZN(n16199) );
  INV_X1 U13881 ( .A(n18974), .ZN(n10903) );
  INV_X1 U13882 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16245) );
  NAND2_X1 U13883 ( .A1(n10903), .A2(n16245), .ZN(n15036) );
  AND2_X1 U13884 ( .A1(n16199), .A2(n15036), .ZN(n10904) );
  INV_X1 U13885 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10906) );
  NOR2_X1 U13886 ( .A1(n10102), .A2(n10906), .ZN(n10905) );
  XNOR2_X1 U13887 ( .A(n10907), .B(n10905), .ZN(n18963) );
  NAND2_X1 U13888 ( .A1(n18963), .A2(n9924), .ZN(n10911) );
  INV_X1 U13889 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15328) );
  AND2_X1 U13890 ( .A1(n10911), .A2(n15328), .ZN(n15322) );
  NAND3_X1 U13891 ( .A1(n10913), .A2(P2_EBX_REG_10__SCAN_IN), .A3(n11016), 
        .ZN(n10909) );
  OR2_X2 U13892 ( .A1(n10908), .A2(n11016), .ZN(n11018) );
  OAI211_X1 U13893 ( .C1(n10913), .C2(P2_EBX_REG_10__SCAN_IN), .A(n10909), .B(
        n11018), .ZN(n18949) );
  OR2_X1 U13894 ( .A1(n18949), .A2(n10981), .ZN(n10910) );
  INV_X1 U13895 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16177) );
  OR3_X1 U13896 ( .A1(n18949), .A2(n10981), .A3(n16177), .ZN(n16180) );
  OR2_X1 U13897 ( .A1(n10911), .A2(n15328), .ZN(n15321) );
  AND2_X1 U13898 ( .A1(n16180), .A2(n15321), .ZN(n10912) );
  NOR2_X2 U13899 ( .A1(n10913), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n14709) );
  INV_X1 U13900 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13233) );
  NAND2_X1 U13901 ( .A1(n14709), .A2(n13233), .ZN(n10917) );
  NAND2_X2 U13902 ( .A1(n10917), .A2(n11018), .ZN(n14710) );
  NOR2_X1 U13903 ( .A1(n14710), .A2(n10981), .ZN(n15305) );
  INV_X1 U13904 ( .A(n15305), .ZN(n10914) );
  INV_X1 U13905 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15310) );
  NAND2_X1 U13906 ( .A1(n10914), .A2(n15310), .ZN(n10915) );
  NAND2_X1 U13907 ( .A1(n11016), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10916) );
  NAND3_X1 U13908 ( .A1(n11016), .A2(P2_EBX_REG_12__SCAN_IN), .A3(n10917), 
        .ZN(n10918) );
  AND2_X1 U13909 ( .A1(n10926), .A2(n10918), .ZN(n10923) );
  INV_X1 U13910 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15216) );
  NOR2_X1 U13911 ( .A1(n10981), .A2(n15216), .ZN(n10919) );
  NAND2_X1 U13912 ( .A1(n10923), .A2(n10919), .ZN(n15290) );
  INV_X1 U13913 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10920) );
  NOR2_X1 U13914 ( .A1(n10102), .A2(n10920), .ZN(n10925) );
  INV_X1 U13915 ( .A(n10925), .ZN(n10921) );
  XNOR2_X1 U13916 ( .A(n10926), .B(n10921), .ZN(n18925) );
  NAND2_X1 U13917 ( .A1(n18925), .A2(n9924), .ZN(n10922) );
  INV_X1 U13918 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15282) );
  NAND2_X1 U13919 ( .A1(n10922), .A2(n15282), .ZN(n15277) );
  INV_X1 U13920 ( .A(n10923), .ZN(n18937) );
  OAI21_X1 U13921 ( .B1(n18937), .B2(n10981), .A(n15216), .ZN(n15291) );
  AND2_X1 U13922 ( .A1(n15277), .A2(n15291), .ZN(n10924) );
  NOR2_X2 U13923 ( .A1(n10926), .A2(n10925), .ZN(n10943) );
  NAND2_X1 U13924 ( .A1(n11016), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10941) );
  INV_X1 U13925 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n10927) );
  NAND2_X2 U13926 ( .A1(n10939), .A2(n11018), .ZN(n10936) );
  NAND2_X1 U13927 ( .A1(n11016), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10935) );
  NOR2_X1 U13928 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(P2_EBX_REG_18__SCAN_IN), 
        .ZN(n10928) );
  NOR2_X1 U13929 ( .A1(n10102), .A2(n10928), .ZN(n10929) );
  INV_X1 U13930 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10930) );
  NAND2_X1 U13931 ( .A1(n10977), .A2(n11018), .ZN(n10974) );
  AND3_X1 U13932 ( .A1(n10950), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n11016), .ZN(
        n10931) );
  OR2_X1 U13933 ( .A1(n10974), .A2(n10931), .ZN(n12565) );
  INV_X1 U13934 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15169) );
  OAI21_X1 U13935 ( .B1(n12565), .B2(n10981), .A(n15169), .ZN(n14955) );
  INV_X1 U13936 ( .A(n10948), .ZN(n10934) );
  INV_X1 U13937 ( .A(n10952), .ZN(n10932) );
  INV_X1 U13938 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n14800) );
  NAND2_X1 U13939 ( .A1(n10932), .A2(n14800), .ZN(n10954) );
  NAND3_X1 U13940 ( .A1(n10954), .A2(P2_EBX_REG_19__SCAN_IN), .A3(n11016), 
        .ZN(n10933) );
  NAND2_X1 U13941 ( .A1(n10934), .A2(n10933), .ZN(n18879) );
  OR2_X2 U13942 ( .A1(n18879), .A2(n10981), .ZN(n10959) );
  INV_X1 U13943 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15195) );
  NAND2_X1 U13944 ( .A1(n10959), .A2(n15195), .ZN(n14979) );
  OAI21_X1 U13945 ( .B1(n10936), .B2(n10935), .A(n10952), .ZN(n18901) );
  INV_X1 U13946 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15004) );
  OAI21_X1 U13947 ( .B1(n18901), .B2(n10981), .A(n15004), .ZN(n14950) );
  NAND3_X1 U13948 ( .A1(n10937), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n11016), 
        .ZN(n10938) );
  AND3_X1 U13949 ( .A1(n10939), .A2(n11018), .A3(n10938), .ZN(n18915) );
  NAND2_X1 U13950 ( .A1(n18915), .A2(n9924), .ZN(n10940) );
  INV_X1 U13951 ( .A(n10941), .ZN(n10942) );
  XNOR2_X1 U13952 ( .A(n10943), .B(n10942), .ZN(n13396) );
  NAND2_X1 U13953 ( .A1(n13396), .A2(n9924), .ZN(n10944) );
  NAND2_X1 U13954 ( .A1(n10944), .A2(n15260), .ZN(n15027) );
  XNOR2_X1 U13955 ( .A(n10945), .B(n9825), .ZN(n12540) );
  NAND2_X1 U13956 ( .A1(n12540), .A2(n9924), .ZN(n10946) );
  INV_X1 U13957 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15252) );
  NAND2_X1 U13958 ( .A1(n10946), .A2(n15252), .ZN(n15016) );
  AND4_X1 U13959 ( .A1(n14950), .A2(n15008), .A3(n15027), .A4(n15016), .ZN(
        n10947) );
  AND2_X1 U13960 ( .A1(n14979), .A2(n10947), .ZN(n10956) );
  NAND2_X1 U13961 ( .A1(n11016), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10949) );
  MUX2_X1 U13962 ( .A(n10949), .B(n11016), .S(n10948), .Z(n10951) );
  NAND2_X1 U13963 ( .A1(n10951), .A2(n10950), .ZN(n14704) );
  INV_X1 U13964 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15179) );
  NAND2_X1 U13965 ( .A1(n10957), .A2(n15179), .ZN(n14970) );
  NAND2_X1 U13966 ( .A1(n11016), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10953) );
  MUX2_X1 U13967 ( .A(n11016), .B(n10953), .S(n10952), .Z(n10955) );
  NAND2_X1 U13968 ( .A1(n10955), .A2(n10954), .ZN(n18893) );
  INV_X1 U13969 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n20943) );
  OAI21_X1 U13970 ( .B1(n18893), .B2(n10981), .A(n20943), .ZN(n14990) );
  NAND4_X1 U13971 ( .A1(n14955), .A2(n10956), .A3(n14970), .A4(n14990), .ZN(
        n10973) );
  INV_X1 U13972 ( .A(n10957), .ZN(n10958) );
  NAND2_X1 U13973 ( .A1(n10958), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14968) );
  INV_X1 U13974 ( .A(n10959), .ZN(n10960) );
  NAND2_X1 U13975 ( .A1(n10960), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14980) );
  INV_X1 U13976 ( .A(n18893), .ZN(n10962) );
  NOR2_X1 U13977 ( .A1(n10981), .A2(n20943), .ZN(n10961) );
  NAND2_X1 U13978 ( .A1(n10962), .A2(n10961), .ZN(n14989) );
  AND2_X1 U13979 ( .A1(n14980), .A2(n14989), .ZN(n14952) );
  OR2_X1 U13980 ( .A1(n10981), .A2(n15004), .ZN(n10963) );
  NOR2_X1 U13981 ( .A1(n18901), .A2(n10963), .ZN(n14948) );
  INV_X1 U13982 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15218) );
  NOR2_X1 U13983 ( .A1(n10981), .A2(n15218), .ZN(n10964) );
  NAND2_X1 U13984 ( .A1(n18915), .A2(n10964), .ZN(n14946) );
  INV_X1 U13985 ( .A(n12540), .ZN(n10965) );
  OR3_X1 U13986 ( .A1(n10965), .A2(n10981), .A3(n15252), .ZN(n15015) );
  NOR2_X1 U13987 ( .A1(n10981), .A2(n15260), .ZN(n10966) );
  NAND2_X1 U13988 ( .A1(n13396), .A2(n10966), .ZN(n15026) );
  NOR2_X1 U13989 ( .A1(n10981), .A2(n15282), .ZN(n10967) );
  NAND2_X1 U13990 ( .A1(n18925), .A2(n10967), .ZN(n15276) );
  NAND4_X1 U13991 ( .A1(n14946), .A2(n15015), .A3(n15026), .A4(n15276), .ZN(
        n10968) );
  NOR2_X1 U13992 ( .A1(n14948), .A2(n10968), .ZN(n10971) );
  INV_X1 U13993 ( .A(n12565), .ZN(n10970) );
  NOR2_X1 U13994 ( .A1(n10981), .A2(n15169), .ZN(n10969) );
  NAND2_X1 U13995 ( .A1(n10970), .A2(n10969), .ZN(n14954) );
  AND4_X1 U13996 ( .A1(n14968), .A2(n14952), .A3(n10971), .A4(n14954), .ZN(
        n10972) );
  NAND2_X1 U13997 ( .A1(n11016), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10975) );
  NAND2_X1 U13998 ( .A1(n10974), .A2(n10975), .ZN(n10986) );
  INV_X1 U13999 ( .A(n10975), .ZN(n10976) );
  NAND2_X1 U14000 ( .A1(n10977), .A2(n10976), .ZN(n10978) );
  NAND2_X1 U14001 ( .A1(n10986), .A2(n10978), .ZN(n15781) );
  OR2_X1 U14002 ( .A1(n15781), .A2(n10981), .ZN(n10979) );
  INV_X1 U14003 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10980) );
  NAND2_X1 U14004 ( .A1(n10979), .A2(n10980), .ZN(n15149) );
  OR2_X1 U14005 ( .A1(n10981), .A2(n10980), .ZN(n10982) );
  NAND2_X1 U14006 ( .A1(n10983), .A2(n15148), .ZN(n15131) );
  INV_X1 U14007 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10984) );
  NOR2_X1 U14008 ( .A1(n10102), .A2(n10984), .ZN(n10985) );
  NAND2_X1 U14009 ( .A1(n10986), .A2(n10985), .ZN(n10987) );
  NAND2_X1 U14010 ( .A1(n12552), .A2(n9924), .ZN(n10988) );
  XNOR2_X1 U14011 ( .A(n10988), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15132) );
  NAND2_X1 U14012 ( .A1(n15131), .A2(n15132), .ZN(n10990) );
  NAND3_X1 U14013 ( .A1(n12552), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n9924), .ZN(n10989) );
  INV_X1 U14014 ( .A(n14935), .ZN(n10993) );
  NAND2_X1 U14015 ( .A1(n11016), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10991) );
  MUX2_X1 U14016 ( .A(P2_EBX_REG_24__SCAN_IN), .B(n10991), .S(n10994), .Z(
        n10992) );
  NAND2_X1 U14017 ( .A1(n10992), .A2(n11018), .ZN(n16107) );
  NOR2_X1 U14018 ( .A1(n16107), .A2(n10981), .ZN(n14933) );
  INV_X1 U14019 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14747) );
  NAND2_X1 U14020 ( .A1(n10995), .A2(n14747), .ZN(n16097) );
  NOR2_X1 U14021 ( .A1(n10995), .A2(n14747), .ZN(n10996) );
  NAND2_X1 U14022 ( .A1(n11016), .A2(n10996), .ZN(n10997) );
  AND2_X1 U14023 ( .A1(n11018), .A2(n10997), .ZN(n10998) );
  NAND2_X1 U14024 ( .A1(n16097), .A2(n10998), .ZN(n14689) );
  OAI21_X1 U14025 ( .B1(n14689), .B2(n10981), .A(n21137), .ZN(n14924) );
  INV_X1 U14026 ( .A(n16082), .ZN(n10999) );
  NOR2_X1 U14027 ( .A1(n16096), .A2(n10981), .ZN(n11005) );
  XNOR2_X1 U14028 ( .A(n11005), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14915) );
  NAND2_X1 U14029 ( .A1(n11016), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16081) );
  INV_X1 U14030 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n11000) );
  NOR2_X1 U14031 ( .A1(n10102), .A2(n11000), .ZN(n11001) );
  AND2_X1 U14032 ( .A1(n16080), .A2(n11001), .ZN(n11002) );
  NAND2_X1 U14033 ( .A1(n14672), .A2(n9924), .ZN(n12040) );
  INV_X1 U14034 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11004) );
  INV_X1 U14035 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15088) );
  NAND2_X1 U14036 ( .A1(n16080), .A2(n9924), .ZN(n12038) );
  AOI22_X1 U14037 ( .A1(n12040), .A2(n11004), .B1(n15088), .B2(n12038), .ZN(
        n11003) );
  NAND2_X1 U14038 ( .A1(n11004), .A2(n15088), .ZN(n12374) );
  INV_X1 U14039 ( .A(n12374), .ZN(n11008) );
  NAND2_X1 U14040 ( .A1(n11005), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11006) );
  NAND2_X1 U14041 ( .A1(n14923), .A2(n11006), .ZN(n12036) );
  INV_X1 U14042 ( .A(n12036), .ZN(n11007) );
  NAND2_X1 U14043 ( .A1(n11016), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11011) );
  NAND2_X1 U14044 ( .A1(n11012), .A2(n11011), .ZN(n11017) );
  NAND2_X1 U14045 ( .A1(n11016), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11013) );
  XNOR2_X1 U14046 ( .A(n11017), .B(n11013), .ZN(n12280) );
  AOI21_X1 U14047 ( .B1(n12280), .B2(n9924), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14887) );
  INV_X1 U14048 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15048) );
  NOR2_X1 U14049 ( .A1(n10981), .A2(n15048), .ZN(n11014) );
  NAND2_X1 U14050 ( .A1(n12280), .A2(n11014), .ZN(n14888) );
  INV_X1 U14051 ( .A(n16066), .ZN(n11015) );
  NAND3_X1 U14052 ( .A1(n11015), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n9924), .ZN(n14897) );
  OAI21_X1 U14053 ( .B1(n11017), .B2(P2_EBX_REG_30__SCAN_IN), .A(n11016), .ZN(
        n11019) );
  NAND2_X1 U14054 ( .A1(n11019), .A2(n11018), .ZN(n16054) );
  NOR2_X1 U14055 ( .A1(n16054), .A2(n10981), .ZN(n11020) );
  XNOR2_X1 U14056 ( .A(n11020), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11021) );
  INV_X1 U14057 ( .A(n12587), .ZN(n11023) );
  AND2_X2 U14058 ( .A1(n11024), .A2(n12774), .ZN(n11728) );
  OAI22_X1 U14059 ( .A1(n11189), .A2(n11026), .B1(n11787), .B2(n11025), .ZN(
        n11034) );
  AND2_X2 U14060 ( .A1(n11038), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12780) );
  NAND2_X1 U14061 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11032) );
  NAND2_X1 U14062 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11031) );
  INV_X2 U14063 ( .A(n11700), .ZN(n11651) );
  NAND2_X1 U14064 ( .A1(n11651), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11030) );
  NAND2_X1 U14065 ( .A1(n11794), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11029) );
  NAND4_X1 U14066 ( .A1(n11032), .A2(n11031), .A3(n11030), .A4(n11029), .ZN(
        n11033) );
  AND2_X4 U14067 ( .A1(n14646), .A2(n12777), .ZN(n11819) );
  AOI22_X1 U14068 ( .A1(n11547), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11043) );
  AND2_X4 U14069 ( .A1(n13147), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11121) );
  NOR2_X1 U14070 ( .A1(n11038), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11039) );
  AOI22_X1 U14071 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11041) );
  NAND3_X1 U14072 ( .A1(n11043), .A2(n11042), .A3(n11041), .ZN(n11050) );
  AND2_X2 U14073 ( .A1(n11044), .A2(n12777), .ZN(n11057) );
  AOI22_X1 U14074 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11057), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11048) );
  AOI22_X1 U14075 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11047) );
  NAND2_X1 U14076 ( .A1(n11048), .A2(n11047), .ZN(n11049) );
  NOR2_X1 U14077 ( .A1(n11050), .A2(n11049), .ZN(n11051) );
  AOI22_X1 U14078 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11056) );
  INV_X2 U14079 ( .A(n11787), .ZN(n11615) );
  AOI22_X1 U14080 ( .A1(n11728), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11615), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11055) );
  INV_X2 U14081 ( .A(n11815), .ZN(n11652) );
  AOI22_X1 U14082 ( .A1(n11652), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11054) );
  AOI22_X1 U14083 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11053) );
  AOI22_X1 U14084 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11057), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11061) );
  AOI22_X1 U14085 ( .A1(n11547), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11060) );
  AOI22_X1 U14086 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11059) );
  AOI22_X1 U14087 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11058) );
  AOI22_X1 U14088 ( .A1(n11767), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11065) );
  AOI22_X1 U14089 ( .A1(n11728), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11064) );
  AOI22_X1 U14090 ( .A1(n11794), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11063) );
  AOI22_X1 U14091 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11062) );
  NAND4_X1 U14092 ( .A1(n11065), .A2(n11064), .A3(n11063), .A4(n11062), .ZN(
        n11071) );
  AOI22_X1 U14093 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11820), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11069) );
  AOI22_X1 U14094 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11068) );
  AOI22_X1 U14095 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9745), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11067) );
  AOI22_X1 U14096 ( .A1(n11547), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11066) );
  NAND4_X1 U14097 ( .A1(n11069), .A2(n11068), .A3(n11067), .A4(n11066), .ZN(
        n11070) );
  OR2_X2 U14098 ( .A1(n11071), .A2(n11070), .ZN(n11131) );
  INV_X2 U14099 ( .A(n11787), .ZN(n11527) );
  AOI22_X1 U14100 ( .A1(n11728), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11615), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11075) );
  AOI22_X1 U14101 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11820), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11074) );
  AOI22_X1 U14102 ( .A1(n11794), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11073) );
  AOI22_X1 U14103 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11072) );
  AOI22_X1 U14104 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11079) );
  AOI22_X1 U14105 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11057), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11078) );
  AOI22_X1 U14106 ( .A1(n11547), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11077) );
  AOI22_X1 U14107 ( .A1(n9746), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11076) );
  AOI22_X1 U14108 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11084) );
  AOI22_X1 U14109 ( .A1(n11728), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11083) );
  AOI22_X1 U14110 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11082) );
  AOI22_X1 U14111 ( .A1(n11547), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11081) );
  NAND4_X1 U14112 ( .A1(n11084), .A2(n11083), .A3(n11082), .A4(n11081), .ZN(
        n11090) );
  AOI22_X1 U14113 ( .A1(n11057), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11820), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11088) );
  AOI22_X1 U14114 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11087) );
  AOI22_X1 U14115 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9745), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11086) );
  INV_X1 U14116 ( .A(n11813), .ZN(n11707) );
  AOI22_X1 U14117 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11085) );
  NAND4_X1 U14118 ( .A1(n11088), .A2(n11087), .A3(n11086), .A4(n11085), .ZN(
        n11089) );
  OR2_X2 U14119 ( .A1(n11090), .A2(n11089), .ZN(n20189) );
  NAND2_X1 U14120 ( .A1(n11131), .A2(n11155), .ZN(n11101) );
  NAND2_X2 U14121 ( .A1(n11131), .A2(n11139), .ZN(n11104) );
  INV_X1 U14122 ( .A(n11104), .ZN(n12415) );
  AOI22_X1 U14123 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11095) );
  AOI22_X1 U14124 ( .A1(n11728), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11615), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11094) );
  AOI22_X1 U14125 ( .A1(n11652), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11093) );
  AOI22_X1 U14126 ( .A1(n11547), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11057), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11099) );
  AOI22_X1 U14127 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11098) );
  AOI22_X1 U14128 ( .A1(n11819), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11097) );
  AOI22_X1 U14129 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11096) );
  MUX2_X1 U14130 ( .A(n11101), .B(n12415), .S(n20184), .Z(n11102) );
  AND3_X2 U14131 ( .A1(n11103), .A2(n10274), .A3(n11102), .ZN(n11143) );
  AOI22_X1 U14132 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11108) );
  AOI22_X1 U14133 ( .A1(n11728), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11615), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11107) );
  AOI22_X1 U14134 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11651), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11106) );
  AOI22_X1 U14135 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n11789), .B1(
        n11176), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11105) );
  NAND4_X1 U14136 ( .A1(n11108), .A2(n11107), .A3(n11106), .A4(n11105), .ZN(
        n11114) );
  AOI22_X1 U14137 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11057), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11112) );
  AOI22_X1 U14138 ( .A1(n11547), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11111) );
  AOI22_X1 U14139 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9745), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11110) );
  AOI22_X1 U14140 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11109) );
  NAND4_X1 U14141 ( .A1(n11112), .A2(n11111), .A3(n11110), .A4(n11109), .ZN(
        n11113) );
  NOR2_X1 U14142 ( .A1(n11104), .A2(n20166), .ZN(n11115) );
  AOI22_X1 U14143 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11057), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11119) );
  AOI22_X1 U14144 ( .A1(n11799), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11118) );
  AOI22_X1 U14145 ( .A1(n11176), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11117) );
  AOI22_X1 U14146 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11116) );
  OAI22_X1 U14147 ( .A1(n11189), .A2(n11123), .B1(n11787), .B2(n11122), .ZN(
        n11129) );
  NAND2_X1 U14148 ( .A1(n11789), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11127) );
  NAND2_X1 U14149 ( .A1(n11547), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11126) );
  NAND2_X1 U14150 ( .A1(n11651), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11125) );
  NAND2_X1 U14151 ( .A1(n11794), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11124) );
  NAND4_X1 U14152 ( .A1(n11127), .A2(n11126), .A3(n11125), .A4(n11124), .ZN(
        n11128) );
  NAND2_X1 U14154 ( .A1(n12620), .A2(n9729), .ZN(n11133) );
  NAND2_X1 U14155 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20784) );
  OAI21_X1 U14156 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(P1_STATE_REG_2__SCAN_IN), 
        .A(n20784), .ZN(n12016) );
  INV_X1 U14157 ( .A(n12016), .ZN(n11134) );
  NAND2_X2 U14158 ( .A1(n11135), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11218) );
  NAND2_X1 U14159 ( .A1(n11136), .A2(n11137), .ZN(n12761) );
  NAND2_X1 U14160 ( .A1(n12761), .A2(n9744), .ZN(n11142) );
  OR2_X1 U14161 ( .A1(n11104), .A2(n12010), .ZN(n12991) );
  NAND2_X1 U14162 ( .A1(n20166), .A2(n20184), .ZN(n12990) );
  NAND2_X1 U14163 ( .A1(n12991), .A2(n12990), .ZN(n12765) );
  NAND2_X1 U14164 ( .A1(n12626), .A2(n20166), .ZN(n20858) );
  NAND2_X1 U14165 ( .A1(n9731), .A2(n9729), .ZN(n12792) );
  INV_X1 U14166 ( .A(n13180), .ZN(n11156) );
  OAI211_X1 U14167 ( .C1(n20858), .C2(n13000), .A(n12792), .B(n11156), .ZN(
        n11140) );
  NOR2_X1 U14168 ( .A1(n12765), .A2(n11140), .ZN(n11141) );
  NAND2_X1 U14169 ( .A1(n11142), .A2(n11141), .ZN(n11144) );
  NAND2_X1 U14170 ( .A1(n11219), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11148) );
  NAND2_X1 U14171 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11221) );
  OAI21_X1 U14172 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11221), .ZN(n20490) );
  NAND2_X1 U14173 ( .A1(n15820), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11216) );
  OAI21_X1 U14174 ( .B1(n12416), .B2(n20490), .A(n11216), .ZN(n11146) );
  INV_X1 U14175 ( .A(n11146), .ZN(n11147) );
  NAND2_X1 U14176 ( .A1(n11148), .A2(n11147), .ZN(n11149) );
  NAND2_X1 U14177 ( .A1(n11219), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11151) );
  INV_X1 U14178 ( .A(n15820), .ZN(n15815) );
  MUX2_X1 U14179 ( .A(n15815), .B(n12416), .S(n20602), .Z(n11150) );
  NAND3_X1 U14180 ( .A1(n12761), .A2(n9729), .A3(n9744), .ZN(n11162) );
  NAND3_X1 U14181 ( .A1(n12763), .A2(n11137), .A3(n20189), .ZN(n11153) );
  NAND2_X1 U14182 ( .A1(n11154), .A2(n11153), .ZN(n11161) );
  OR2_X1 U14183 ( .A1(n11156), .A2(n11155), .ZN(n12989) );
  NAND4_X1 U14184 ( .A1(n12989), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n14657), 
        .A4(n12792), .ZN(n11157) );
  NOR2_X1 U14185 ( .A1(n11157), .A2(n12765), .ZN(n11160) );
  INV_X1 U14186 ( .A(n11136), .ZN(n11158) );
  NAND2_X1 U14187 ( .A1(n11158), .A2(n13002), .ZN(n11159) );
  NAND4_X1 U14188 ( .A1(n11162), .A2(n11161), .A3(n11160), .A4(n11159), .ZN(
        n11330) );
  INV_X1 U14189 ( .A(n11263), .ZN(n11188) );
  AOI22_X1 U14190 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11167) );
  AOI22_X1 U14191 ( .A1(n11728), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11166) );
  AOI22_X1 U14192 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11165) );
  AOI22_X1 U14193 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11460), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11164) );
  NAND4_X1 U14194 ( .A1(n11167), .A2(n11166), .A3(n11165), .A4(n11164), .ZN(
        n11174) );
  AOI22_X1 U14195 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11800), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11172) );
  AOI22_X1 U14196 ( .A1(n11547), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11171) );
  AOI22_X1 U14197 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11170) );
  AOI22_X1 U14198 ( .A1(n9751), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11169) );
  NAND4_X1 U14199 ( .A1(n11172), .A2(n11171), .A3(n11170), .A4(n11169), .ZN(
        n11173) );
  NAND2_X1 U14200 ( .A1(n11188), .A2(n12431), .ZN(n11175) );
  OAI21_X2 U14201 ( .B1(n13170), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11175), 
        .ZN(n12436) );
  AOI22_X1 U14202 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11180) );
  AOI22_X1 U14203 ( .A1(n11728), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11615), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11179) );
  AOI22_X1 U14204 ( .A1(n11652), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11178) );
  AOI22_X1 U14205 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11460), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11177) );
  NAND4_X1 U14206 ( .A1(n11180), .A2(n11179), .A3(n11178), .A4(n11177), .ZN(
        n11186) );
  AOI22_X1 U14207 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11184) );
  INV_X1 U14208 ( .A(n11547), .ZN(n11661) );
  INV_X2 U14209 ( .A(n11661), .ZN(n11644) );
  AOI22_X1 U14210 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11183) );
  AOI22_X1 U14211 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11182) );
  AOI22_X1 U14212 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11181) );
  NAND4_X1 U14213 ( .A1(n11184), .A2(n11183), .A3(n11182), .A4(n11181), .ZN(
        n11185) );
  INV_X1 U14214 ( .A(n12496), .ZN(n11187) );
  NAND2_X1 U14215 ( .A1(n13000), .A2(n12496), .ZN(n11205) );
  AOI22_X1 U14216 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n11121), .B1(
        n11120), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11193) );
  INV_X2 U14217 ( .A(n11189), .ZN(n11829) );
  AOI22_X1 U14218 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n11615), .B1(
        n11829), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11192) );
  AOI22_X1 U14219 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11191) );
  AOI22_X1 U14220 ( .A1(n11460), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9745), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11190) );
  NAND4_X1 U14221 ( .A1(n11193), .A2(n11192), .A3(n11191), .A4(n11190), .ZN(
        n11200) );
  AOI22_X1 U14222 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11820), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11198) );
  AOI22_X1 U14223 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n11644), .B1(
        n11800), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11197) );
  AOI22_X1 U14224 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n9747), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11196) );
  AOI22_X1 U14225 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11195) );
  NAND4_X1 U14226 ( .A1(n11198), .A2(n11197), .A3(n11196), .A4(n11195), .ZN(
        n11199) );
  INV_X1 U14227 ( .A(n12439), .ZN(n11201) );
  MUX2_X1 U14228 ( .A(n11209), .B(n11208), .S(n11201), .Z(n11202) );
  INV_X1 U14229 ( .A(n11202), .ZN(n11203) );
  INV_X1 U14230 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11207) );
  AOI21_X1 U14231 ( .B1(n9731), .B2(n12439), .A(n20773), .ZN(n11206) );
  NAND2_X1 U14232 ( .A1(n11326), .A2(n12424), .ZN(n11317) );
  INV_X1 U14233 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11213) );
  INV_X1 U14234 ( .A(n11209), .ZN(n11212) );
  NAND2_X1 U14235 ( .A1(n11210), .A2(n12431), .ZN(n11211) );
  OAI211_X1 U14236 ( .C1(n11213), .C2(n11889), .A(n11212), .B(n11211), .ZN(
        n11318) );
  NAND2_X1 U14237 ( .A1(n12436), .A2(n11317), .ZN(n11214) );
  AND2_X1 U14238 ( .A1(n11216), .A2(n11027), .ZN(n11217) );
  NAND2_X1 U14239 ( .A1(n11250), .A2(n11247), .ZN(n11226) );
  NAND2_X1 U14240 ( .A1(n11219), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11224) );
  INV_X1 U14241 ( .A(n12416), .ZN(n11229) );
  INV_X1 U14242 ( .A(n11221), .ZN(n11220) );
  NAND2_X1 U14243 ( .A1(n11220), .A2(n20566), .ZN(n20528) );
  NAND2_X1 U14244 ( .A1(n11221), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11222) );
  NAND2_X1 U14245 ( .A1(n20528), .A2(n11222), .ZN(n20174) );
  NAND2_X1 U14246 ( .A1(n11229), .A2(n20174), .ZN(n11223) );
  NAND2_X1 U14247 ( .A1(n11224), .A2(n11223), .ZN(n11245) );
  NAND2_X1 U14248 ( .A1(n11219), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11231) );
  NAND3_X1 U14249 ( .A1(n20565), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20415) );
  INV_X1 U14250 ( .A(n20415), .ZN(n11227) );
  NAND2_X1 U14251 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11227), .ZN(
        n20413) );
  NAND2_X1 U14252 ( .A1(n20565), .A2(n20413), .ZN(n11228) );
  NOR3_X1 U14253 ( .A1(n20565), .A2(n20566), .A3(n20492), .ZN(n20718) );
  NAND2_X1 U14254 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20718), .ZN(
        n20707) );
  AOI22_X1 U14255 ( .A1(n11229), .A2(n20443), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15820), .ZN(n11230) );
  AOI22_X1 U14256 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11236) );
  AOI22_X1 U14257 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11615), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11235) );
  AOI22_X1 U14258 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11234) );
  AOI22_X1 U14259 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11460), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11233) );
  NAND4_X1 U14260 ( .A1(n11236), .A2(n11235), .A3(n11234), .A4(n11233), .ZN(
        n11242) );
  AOI22_X1 U14261 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11800), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11240) );
  AOI22_X1 U14262 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11239) );
  AOI22_X1 U14263 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9745), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11238) );
  AOI22_X1 U14264 ( .A1(n9751), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11237) );
  NAND4_X1 U14265 ( .A1(n11240), .A2(n11239), .A3(n11238), .A4(n11237), .ZN(
        n11241) );
  AOI22_X1 U14266 ( .A1(n11895), .A2(n12465), .B1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n11898), .ZN(n11243) );
  INV_X1 U14267 ( .A(n11245), .ZN(n11249) );
  INV_X1 U14268 ( .A(n11246), .ZN(n11248) );
  NAND2_X1 U14269 ( .A1(n10260), .A2(n11250), .ZN(n11251) );
  AOI22_X1 U14270 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11256) );
  AOI22_X1 U14271 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11255) );
  AOI22_X1 U14272 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11651), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11254) );
  AOI22_X1 U14273 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11460), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11253) );
  NAND4_X1 U14274 ( .A1(n11256), .A2(n11255), .A3(n11254), .A4(n11253), .ZN(
        n11262) );
  AOI22_X1 U14275 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11800), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11260) );
  AOI22_X1 U14276 ( .A1(n11547), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11259) );
  AOI22_X1 U14277 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9745), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11258) );
  AOI22_X1 U14278 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11257) );
  NAND4_X1 U14279 ( .A1(n11260), .A2(n11259), .A3(n11258), .A4(n11257), .ZN(
        n11261) );
  INV_X1 U14280 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11264) );
  OAI22_X1 U14281 ( .A1(n12449), .A2(n11265), .B1(n11889), .B2(n11264), .ZN(
        n11266) );
  INV_X1 U14282 ( .A(n11343), .ZN(n11267) );
  AND2_X2 U14283 ( .A1(n11344), .A2(n11267), .ZN(n11268) );
  AOI22_X1 U14284 ( .A1(n11767), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11272) );
  AOI22_X1 U14285 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11271) );
  AOI22_X1 U14286 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11270) );
  AOI22_X1 U14287 ( .A1(n11460), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11269) );
  NAND4_X1 U14288 ( .A1(n11272), .A2(n11271), .A3(n11270), .A4(n11269), .ZN(
        n11278) );
  AOI22_X1 U14289 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11276) );
  AOI22_X1 U14290 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11275) );
  AOI22_X1 U14291 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9745), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11274) );
  AOI22_X1 U14292 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11273) );
  NAND4_X1 U14293 ( .A1(n11276), .A2(n11275), .A3(n11274), .A4(n11273), .ZN(
        n11277) );
  NAND2_X1 U14294 ( .A1(n11895), .A2(n12464), .ZN(n11280) );
  NAND2_X1 U14295 ( .A1(n11898), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11279) );
  AOI22_X1 U14296 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11284) );
  AOI22_X1 U14297 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11615), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11283) );
  AOI22_X1 U14298 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11282) );
  AOI22_X1 U14299 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11460), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11281) );
  NAND4_X1 U14300 ( .A1(n11284), .A2(n11283), .A3(n11282), .A4(n11281), .ZN(
        n11290) );
  AOI22_X1 U14301 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11800), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11288) );
  AOI22_X1 U14302 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11287) );
  AOI22_X1 U14303 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9746), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11286) );
  INV_X1 U14304 ( .A(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n21008) );
  AOI22_X1 U14305 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11285) );
  NAND4_X1 U14306 ( .A1(n11288), .A2(n11287), .A3(n11286), .A4(n11285), .ZN(
        n11289) );
  NAND2_X1 U14307 ( .A1(n11895), .A2(n12475), .ZN(n11292) );
  NAND2_X1 U14308 ( .A1(n11898), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11291) );
  NAND2_X1 U14309 ( .A1(n11292), .A2(n11291), .ZN(n11367) );
  INV_X1 U14310 ( .A(n11367), .ZN(n11293) );
  AOI22_X1 U14311 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11297) );
  AOI22_X1 U14312 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11615), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11296) );
  AOI22_X1 U14313 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11651), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11295) );
  AOI22_X1 U14314 ( .A1(n11460), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9745), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11294) );
  NAND4_X1 U14315 ( .A1(n11297), .A2(n11296), .A3(n11295), .A4(n11294), .ZN(
        n11303) );
  AOI22_X1 U14316 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9747), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11301) );
  AOI22_X1 U14317 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11300) );
  AOI22_X1 U14318 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9752), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11299) );
  AOI22_X1 U14319 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11298) );
  NAND4_X1 U14320 ( .A1(n11301), .A2(n11300), .A3(n11299), .A4(n11298), .ZN(
        n11302) );
  AOI22_X1 U14321 ( .A1(n11895), .A2(n12488), .B1(n11898), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11373) );
  NAND2_X1 U14322 ( .A1(n11895), .A2(n12496), .ZN(n11305) );
  NAND2_X1 U14323 ( .A1(n11898), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11304) );
  NAND2_X1 U14324 ( .A1(n11305), .A2(n11304), .ZN(n11306) );
  INV_X2 U14325 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n11307) );
  INV_X1 U14326 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11310) );
  NAND2_X1 U14327 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11348) );
  INV_X1 U14328 ( .A(n11348), .ZN(n11308) );
  OAI21_X1 U14329 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n11376), .A(
        n11401), .ZN(n19986) );
  AOI22_X1 U14330 ( .A1(n11914), .A2(n19986), .B1(n11846), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11309) );
  OAI21_X1 U14331 ( .B1(n11689), .B2(n11310), .A(n11309), .ZN(n11311) );
  INV_X1 U14332 ( .A(n12970), .ZN(n12394) );
  NAND2_X1 U14333 ( .A1(n12394), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11364) );
  XNOR2_X1 U14334 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13379) );
  AOI21_X1 U14335 ( .B1(n11338), .B2(n13379), .A(n11846), .ZN(n11314) );
  NAND2_X1 U14336 ( .A1(n11847), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11313) );
  OAI211_X1 U14337 ( .C1(n11364), .C2(n11038), .A(n11314), .B(n11313), .ZN(
        n11315) );
  INV_X1 U14338 ( .A(n11315), .ZN(n11316) );
  NAND2_X1 U14339 ( .A1(n11846), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11342) );
  INV_X1 U14340 ( .A(n13121), .ZN(n11341) );
  INV_X1 U14341 ( .A(n11318), .ZN(n11319) );
  NAND2_X1 U14342 ( .A1(n20247), .A2(n11500), .ZN(n11325) );
  AOI22_X1 U14343 ( .A1(n11847), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n11307), .ZN(n11323) );
  INV_X1 U14344 ( .A(n11364), .ZN(n11321) );
  NAND2_X1 U14345 ( .A1(n11321), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11322) );
  AND2_X1 U14346 ( .A1(n11323), .A2(n11322), .ZN(n11324) );
  NAND2_X1 U14347 ( .A1(n11325), .A2(n11324), .ZN(n13054) );
  NAND2_X1 U14348 ( .A1(n12437), .A2(n11328), .ZN(n11329) );
  NAND2_X1 U14349 ( .A1(n11329), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12928) );
  INV_X1 U14350 ( .A(n11330), .ZN(n11331) );
  XNOR2_X1 U14351 ( .A(n11332), .B(n11331), .ZN(n20284) );
  NAND2_X1 U14352 ( .A1(n11307), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11335) );
  NAND2_X1 U14353 ( .A1(n11333), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11334) );
  OAI211_X1 U14354 ( .C1(n11364), .C2(n13568), .A(n11335), .B(n11334), .ZN(
        n11336) );
  AOI21_X1 U14355 ( .B1(n20284), .B2(n11500), .A(n11336), .ZN(n11337) );
  OR2_X1 U14356 ( .A1(n12928), .A2(n11337), .ZN(n12929) );
  INV_X1 U14357 ( .A(n11337), .ZN(n12930) );
  OR2_X1 U14358 ( .A1(n12930), .A2(n11845), .ZN(n11339) );
  NAND2_X1 U14359 ( .A1(n12929), .A2(n11339), .ZN(n13053) );
  NAND2_X1 U14360 ( .A1(n13054), .A2(n13053), .ZN(n13122) );
  NAND2_X1 U14361 ( .A1(n11341), .A2(n11340), .ZN(n13123) );
  NAND2_X1 U14362 ( .A1(n11267), .A2(n11312), .ZN(n11345) );
  NAND2_X1 U14363 ( .A1(n11345), .A2(n13404), .ZN(n11346) );
  INV_X1 U14364 ( .A(n11347), .ZN(n11358) );
  INV_X1 U14365 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11349) );
  NAND2_X1 U14366 ( .A1(n11349), .A2(n11348), .ZN(n11350) );
  NAND2_X1 U14367 ( .A1(n11358), .A2(n11350), .ZN(n13366) );
  AOI22_X1 U14368 ( .A1(n13366), .A2(n11914), .B1(n11846), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11352) );
  NAND2_X1 U14369 ( .A1(n11847), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11351) );
  OAI211_X1 U14370 ( .C1(n11364), .C2(n12774), .A(n11352), .B(n11351), .ZN(
        n11353) );
  INV_X1 U14371 ( .A(n11353), .ZN(n11354) );
  NAND2_X1 U14372 ( .A1(n13198), .A2(n13199), .ZN(n13214) );
  XNOR2_X1 U14373 ( .A(n11356), .B(n11355), .ZN(n12455) );
  INV_X1 U14374 ( .A(n11369), .ZN(n11360) );
  INV_X1 U14375 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11357) );
  NAND2_X1 U14376 ( .A1(n11358), .A2(n11357), .ZN(n11359) );
  NAND2_X1 U14377 ( .A1(n11360), .A2(n11359), .ZN(n20121) );
  INV_X1 U14378 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n11363) );
  NAND2_X1 U14379 ( .A1(n11307), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11362) );
  NAND2_X1 U14380 ( .A1(n11847), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11361) );
  OAI211_X1 U14381 ( .C1(n11364), .C2(n11363), .A(n11362), .B(n11361), .ZN(
        n11365) );
  MUX2_X1 U14382 ( .A(n20121), .B(n11365), .S(n11845), .Z(n11366) );
  AOI21_X1 U14383 ( .B1(n12455), .B2(n11500), .A(n11366), .ZN(n13213) );
  XNOR2_X1 U14384 ( .A(n11368), .B(n11367), .ZN(n12463) );
  INV_X1 U14385 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13268) );
  OAI21_X1 U14386 ( .B1(n11369), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n11375), .ZN(n20017) );
  AOI22_X1 U14387 ( .A1(n20017), .A2(n11914), .B1(n11846), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11370) );
  OAI21_X1 U14388 ( .B1(n11689), .B2(n13268), .A(n11370), .ZN(n11371) );
  AOI21_X1 U14389 ( .B1(n12463), .B2(n11500), .A(n11371), .ZN(n13265) );
  NAND2_X1 U14390 ( .A1(n13212), .A2(n11372), .ZN(n13264) );
  NAND2_X1 U14391 ( .A1(n11374), .A2(n11373), .ZN(n12473) );
  INV_X1 U14392 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11382) );
  NAND2_X1 U14393 ( .A1(n11375), .A2(n11379), .ZN(n11378) );
  INV_X1 U14394 ( .A(n11376), .ZN(n11377) );
  NAND2_X1 U14395 ( .A1(n11378), .A2(n11377), .ZN(n19995) );
  INV_X1 U14396 ( .A(n11846), .ZN(n11539) );
  NOR2_X1 U14397 ( .A1(n11539), .A2(n11379), .ZN(n11380) );
  AOI21_X1 U14398 ( .B1(n19995), .B2(n11914), .A(n11380), .ZN(n11381) );
  OAI21_X1 U14399 ( .B1(n11689), .B2(n11382), .A(n11381), .ZN(n11383) );
  AOI22_X1 U14400 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11389) );
  AOI22_X1 U14401 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n11829), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11388) );
  AOI22_X1 U14402 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n11652), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11387) );
  AOI22_X1 U14403 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n9747), .B1(
        n11460), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11386) );
  NAND4_X1 U14404 ( .A1(n11389), .A2(n11388), .A3(n11387), .A4(n11386), .ZN(
        n11395) );
  AOI22_X1 U14405 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11393) );
  AOI22_X1 U14406 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n11644), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11392) );
  AOI22_X1 U14407 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9752), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11391) );
  AOI22_X1 U14408 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11390) );
  NAND4_X1 U14409 ( .A1(n11393), .A2(n11392), .A3(n11391), .A4(n11390), .ZN(
        n11394) );
  NOR2_X1 U14410 ( .A1(n11395), .A2(n11394), .ZN(n11399) );
  INV_X1 U14411 ( .A(n11401), .ZN(n11396) );
  XNOR2_X1 U14412 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n11396), .ZN(
        n14131) );
  AOI22_X1 U14413 ( .A1(n11914), .A2(n14131), .B1(n11846), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11398) );
  NAND2_X1 U14414 ( .A1(n11847), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11397) );
  OAI211_X1 U14415 ( .C1(n10179), .C2(n11399), .A(n11398), .B(n11397), .ZN(
        n13474) );
  XOR2_X1 U14416 ( .A(n13521), .B(n11426), .Z(n13552) );
  AOI22_X1 U14417 ( .A1(n11767), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11405) );
  AOI22_X1 U14418 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11404) );
  AOI22_X1 U14419 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11403) );
  AOI22_X1 U14420 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11460), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11402) );
  NAND4_X1 U14421 ( .A1(n11405), .A2(n11404), .A3(n11403), .A4(n11402), .ZN(
        n11411) );
  AOI22_X1 U14422 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11409) );
  AOI22_X1 U14423 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11408) );
  AOI22_X1 U14424 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11638), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11407) );
  AOI22_X1 U14425 ( .A1(n9751), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11406) );
  NAND4_X1 U14426 ( .A1(n11409), .A2(n11408), .A3(n11407), .A4(n11406), .ZN(
        n11410) );
  OR2_X1 U14427 ( .A1(n11411), .A2(n11410), .ZN(n11412) );
  AOI22_X1 U14428 ( .A1(n11500), .A2(n11412), .B1(n11846), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11414) );
  NAND2_X1 U14429 ( .A1(n11847), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11413) );
  OAI211_X1 U14430 ( .C1(n13552), .C2(n11845), .A(n11414), .B(n11413), .ZN(
        n13511) );
  AOI22_X1 U14431 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11419) );
  AOI22_X1 U14432 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11418) );
  AOI22_X1 U14433 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11651), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11417) );
  AOI22_X1 U14434 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11416) );
  NAND4_X1 U14435 ( .A1(n11419), .A2(n11418), .A3(n11417), .A4(n11416), .ZN(
        n11425) );
  AOI22_X1 U14436 ( .A1(n11460), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U14437 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9752), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11422) );
  AOI22_X1 U14438 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11638), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11421) );
  AOI22_X1 U14439 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11420) );
  NAND4_X1 U14440 ( .A1(n11423), .A2(n11422), .A3(n11421), .A4(n11420), .ZN(
        n11424) );
  NOR2_X1 U14441 ( .A1(n11425), .A2(n11424), .ZN(n11429) );
  XNOR2_X1 U14442 ( .A(n11441), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14446) );
  NAND2_X1 U14443 ( .A1(n14446), .A2(n11914), .ZN(n11428) );
  AOI22_X1 U14444 ( .A1(n11847), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n11846), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11427) );
  OAI211_X1 U14445 ( .C1(n11429), .C2(n10179), .A(n11428), .B(n11427), .ZN(
        n13531) );
  NAND2_X1 U14446 ( .A1(n13510), .A2(n13531), .ZN(n13529) );
  AOI22_X1 U14447 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11433) );
  AOI22_X1 U14448 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11432) );
  AOI22_X1 U14449 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11651), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11431) );
  AOI22_X1 U14450 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11460), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11430) );
  NAND4_X1 U14451 ( .A1(n11433), .A2(n11432), .A3(n11431), .A4(n11430), .ZN(
        n11439) );
  AOI22_X1 U14452 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11437) );
  AOI22_X1 U14453 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11436) );
  AOI22_X1 U14454 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11638), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U14455 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11790), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11434) );
  NAND4_X1 U14456 ( .A1(n11437), .A2(n11436), .A3(n11435), .A4(n11434), .ZN(
        n11438) );
  NOR2_X1 U14457 ( .A1(n11439), .A2(n11438), .ZN(n11440) );
  INV_X1 U14458 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11444) );
  OAI21_X1 U14459 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11442), .A(
        n11471), .ZN(n15945) );
  NAND2_X1 U14460 ( .A1(n15945), .A2(n11914), .ZN(n11443) );
  OAI21_X1 U14461 ( .B1(n11444), .B2(n11539), .A(n11443), .ZN(n11445) );
  AOI21_X1 U14462 ( .B1(n11847), .B2(P1_EAX_REG_11__SCAN_IN), .A(n11445), .ZN(
        n14103) );
  INV_X1 U14463 ( .A(n14103), .ZN(n11446) );
  INV_X1 U14464 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14284) );
  AOI22_X1 U14465 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11450) );
  AOI22_X1 U14466 ( .A1(n9751), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n9723), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11449) );
  AOI22_X1 U14467 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11638), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11448) );
  AOI22_X1 U14468 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11447) );
  NAND4_X1 U14469 ( .A1(n11450), .A2(n11449), .A3(n11448), .A4(n11447), .ZN(
        n11456) );
  AOI22_X1 U14470 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11454) );
  AOI22_X1 U14471 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11615), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11453) );
  AOI22_X1 U14472 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11452) );
  AOI22_X1 U14473 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11460), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11451) );
  NAND4_X1 U14474 ( .A1(n11454), .A2(n11453), .A3(n11452), .A4(n11451), .ZN(
        n11455) );
  OAI21_X1 U14475 ( .B1(n11456), .B2(n11455), .A(n11500), .ZN(n11459) );
  INV_X1 U14476 ( .A(n11476), .ZN(n11457) );
  XNOR2_X1 U14477 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n11457), .ZN(
        n14440) );
  AOI22_X1 U14478 ( .A1(n11914), .A2(n14440), .B1(n11846), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11458) );
  OAI211_X1 U14479 ( .C1(n11689), .C2(n14284), .A(n11459), .B(n11458), .ZN(
        n14105) );
  AOI22_X1 U14480 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11460), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U14481 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9752), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11463) );
  AOI22_X1 U14482 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11462) );
  AOI22_X1 U14483 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11461) );
  NAND4_X1 U14484 ( .A1(n11464), .A2(n11463), .A3(n11462), .A4(n11461), .ZN(
        n11470) );
  AOI22_X1 U14485 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11468) );
  AOI22_X1 U14486 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11467) );
  AOI22_X1 U14487 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11651), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11466) );
  AOI22_X1 U14488 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11638), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11465) );
  NAND4_X1 U14489 ( .A1(n11468), .A2(n11467), .A3(n11466), .A4(n11465), .ZN(
        n11469) );
  OAI21_X1 U14490 ( .B1(n11470), .B2(n11469), .A(n11500), .ZN(n11475) );
  NAND2_X1 U14491 ( .A1(n11847), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11474) );
  XNOR2_X1 U14492 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11471), .ZN(
        n15931) );
  OAI22_X1 U14493 ( .A1(n15931), .A2(n11845), .B1(n11539), .B2(n15881), .ZN(
        n11472) );
  INV_X1 U14494 ( .A(n11472), .ZN(n11473) );
  NAND3_X1 U14495 ( .A1(n11475), .A2(n11474), .A3(n11473), .ZN(n14192) );
  XOR2_X1 U14496 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n11491), .Z(
        n15926) );
  AOI22_X1 U14497 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11481) );
  AOI22_X1 U14498 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11615), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U14499 ( .A1(n11477), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11651), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11479) );
  AOI22_X1 U14500 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11638), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11478) );
  NAND4_X1 U14501 ( .A1(n11481), .A2(n11480), .A3(n11479), .A4(n11478), .ZN(
        n11487) );
  AOI22_X1 U14502 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11485) );
  AOI22_X1 U14503 ( .A1(n11460), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11057), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11484) );
  AOI22_X1 U14504 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11483) );
  AOI22_X1 U14505 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11482) );
  NAND4_X1 U14506 ( .A1(n11485), .A2(n11484), .A3(n11483), .A4(n11482), .ZN(
        n11486) );
  OR2_X1 U14507 ( .A1(n11487), .A2(n11486), .ZN(n11488) );
  AOI22_X1 U14508 ( .A1(n11500), .A2(n11488), .B1(n11846), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11490) );
  NAND2_X1 U14509 ( .A1(n11847), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11489) );
  OAI211_X1 U14510 ( .C1(n15926), .C2(n11845), .A(n11490), .B(n11489), .ZN(
        n14091) );
  XNOR2_X1 U14511 ( .A(n11523), .B(n14083), .ZN(n14427) );
  AOI22_X1 U14512 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11057), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11495) );
  AOI22_X1 U14513 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n9723), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11494) );
  AOI22_X1 U14514 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11638), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11493) );
  AOI22_X1 U14515 ( .A1(n11460), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11492) );
  NAND4_X1 U14516 ( .A1(n11495), .A2(n11494), .A3(n11493), .A4(n11492), .ZN(
        n11502) );
  AOI22_X1 U14517 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11499) );
  AOI22_X1 U14518 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11615), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11498) );
  AOI22_X1 U14519 ( .A1(n11652), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11651), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11497) );
  AOI22_X1 U14520 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11496) );
  NAND4_X1 U14521 ( .A1(n11499), .A2(n11498), .A3(n11497), .A4(n11496), .ZN(
        n11501) );
  OAI21_X1 U14522 ( .B1(n11502), .B2(n11501), .A(n11500), .ZN(n11505) );
  NAND2_X1 U14523 ( .A1(n11847), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11504) );
  NAND2_X1 U14524 ( .A1(n11846), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11503) );
  NAND3_X1 U14525 ( .A1(n11505), .A2(n11504), .A3(n11503), .ZN(n11506) );
  AOI21_X1 U14526 ( .B1(n14427), .B2(n11914), .A(n11506), .ZN(n14078) );
  AOI22_X1 U14527 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n11767), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U14528 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n11615), .B1(
        n11829), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11511) );
  AOI22_X1 U14529 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n11652), .B1(
        n11651), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11510) );
  AOI22_X1 U14530 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n9747), .B1(
        n11460), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11509) );
  NAND4_X1 U14531 ( .A1(n11512), .A2(n11511), .A3(n11510), .A4(n11509), .ZN(
        n11518) );
  AOI22_X1 U14532 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11516) );
  AOI22_X1 U14533 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n11194), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11515) );
  AOI22_X1 U14534 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11514) );
  AOI22_X1 U14535 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11513) );
  NAND4_X1 U14536 ( .A1(n11516), .A2(n11515), .A3(n11514), .A4(n11513), .ZN(
        n11517) );
  NOR2_X1 U14537 ( .A1(n11518), .A2(n11517), .ZN(n11522) );
  NAND2_X1 U14538 ( .A1(n11307), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11519) );
  NAND2_X1 U14539 ( .A1(n11845), .A2(n11519), .ZN(n11520) );
  AOI21_X1 U14540 ( .B1(n11847), .B2(P1_EAX_REG_16__SCAN_IN), .A(n11520), .ZN(
        n11521) );
  OAI21_X1 U14541 ( .B1(n11842), .B2(n11522), .A(n11521), .ZN(n11526) );
  OAI21_X1 U14542 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n11524), .A(
        n11558), .ZN(n15918) );
  OR2_X1 U14543 ( .A1(n11845), .A2(n15918), .ZN(n11525) );
  NAND2_X1 U14544 ( .A1(n11526), .A2(n11525), .ZN(n14271) );
  AOI22_X1 U14545 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11531) );
  AOI22_X1 U14546 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11530) );
  AOI22_X1 U14547 ( .A1(n11652), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11651), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11529) );
  AOI22_X1 U14548 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11638), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11528) );
  NAND4_X1 U14549 ( .A1(n11531), .A2(n11530), .A3(n11529), .A4(n11528), .ZN(
        n11537) );
  AOI22_X1 U14550 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11535) );
  AOI22_X1 U14551 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11534) );
  AOI22_X1 U14552 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11533) );
  AOI22_X1 U14553 ( .A1(n11460), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11532) );
  NAND4_X1 U14554 ( .A1(n11535), .A2(n11534), .A3(n11533), .A4(n11532), .ZN(
        n11536) );
  OR2_X1 U14555 ( .A1(n11537), .A2(n11536), .ZN(n11538) );
  NAND2_X1 U14556 ( .A1(n11806), .A2(n11538), .ZN(n11542) );
  XNOR2_X1 U14557 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11558), .ZN(
        n14420) );
  INV_X1 U14558 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14415) );
  OAI22_X1 U14559 ( .A1(n11845), .A2(n14420), .B1(n11539), .B2(n14415), .ZN(
        n11540) );
  AOI21_X1 U14560 ( .B1(n11847), .B2(P1_EAX_REG_17__SCAN_IN), .A(n11540), .ZN(
        n11541) );
  NAND2_X1 U14561 ( .A1(n11542), .A2(n11541), .ZN(n14066) );
  AOI22_X1 U14562 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U14563 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11615), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11545) );
  AOI22_X1 U14564 ( .A1(n11652), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11651), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11544) );
  AOI22_X1 U14565 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11638), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11543) );
  NAND4_X1 U14566 ( .A1(n11546), .A2(n11545), .A3(n11544), .A4(n11543), .ZN(
        n11553) );
  AOI22_X1 U14567 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11644), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U14568 ( .A1(n11460), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11550) );
  AOI22_X1 U14569 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9752), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11549) );
  AOI22_X1 U14570 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11548) );
  NAND4_X1 U14571 ( .A1(n11551), .A2(n11550), .A3(n11549), .A4(n11548), .ZN(
        n11552) );
  NOR2_X1 U14572 ( .A1(n11553), .A2(n11552), .ZN(n11557) );
  NAND2_X1 U14573 ( .A1(n11307), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11554) );
  NAND2_X1 U14574 ( .A1(n11845), .A2(n11554), .ZN(n11555) );
  AOI21_X1 U14575 ( .B1(n11847), .B2(P1_EAX_REG_18__SCAN_IN), .A(n11555), .ZN(
        n11556) );
  OAI21_X1 U14576 ( .B1(n11842), .B2(n11557), .A(n11556), .ZN(n11562) );
  OAI21_X1 U14577 ( .B1(n11560), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n11592), .ZN(n15868) );
  OR2_X1 U14578 ( .A1(n15868), .A2(n11845), .ZN(n11561) );
  AOI22_X1 U14579 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11566) );
  AOI22_X1 U14580 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11565) );
  AOI22_X1 U14581 ( .A1(n11652), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11651), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U14582 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11563) );
  NAND4_X1 U14583 ( .A1(n11566), .A2(n11565), .A3(n11564), .A4(n11563), .ZN(
        n11572) );
  AOI22_X1 U14584 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11460), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U14585 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U14586 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9752), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11568) );
  AOI22_X1 U14587 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11567) );
  NAND4_X1 U14588 ( .A1(n11570), .A2(n11569), .A3(n11568), .A4(n11567), .ZN(
        n11571) );
  NOR2_X1 U14589 ( .A1(n11572), .A2(n11571), .ZN(n11575) );
  OAI21_X1 U14590 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14399), .A(n11845), 
        .ZN(n11573) );
  AOI21_X1 U14591 ( .B1(n11847), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11573), .ZN(
        n11574) );
  OAI21_X1 U14592 ( .B1(n11842), .B2(n11575), .A(n11574), .ZN(n11577) );
  XNOR2_X1 U14593 ( .A(n11592), .B(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14397) );
  NAND2_X1 U14594 ( .A1(n14397), .A2(n11914), .ZN(n11576) );
  NAND2_X1 U14595 ( .A1(n11577), .A2(n11576), .ZN(n14049) );
  AOI22_X1 U14596 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11581) );
  AOI22_X1 U14597 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11580) );
  AOI22_X1 U14598 ( .A1(n11652), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11651), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U14599 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11460), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11578) );
  NAND4_X1 U14600 ( .A1(n11581), .A2(n11580), .A3(n11579), .A4(n11578), .ZN(
        n11587) );
  AOI22_X1 U14601 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9752), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11585) );
  AOI22_X1 U14602 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U14603 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11638), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U14604 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11582) );
  NAND4_X1 U14605 ( .A1(n11585), .A2(n11584), .A3(n11583), .A4(n11582), .ZN(
        n11586) );
  NOR2_X1 U14606 ( .A1(n11587), .A2(n11586), .ZN(n11591) );
  NAND2_X1 U14607 ( .A1(n11307), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11588) );
  NAND2_X1 U14608 ( .A1(n11845), .A2(n11588), .ZN(n11589) );
  AOI21_X1 U14609 ( .B1(n11847), .B2(P1_EAX_REG_20__SCAN_IN), .A(n11589), .ZN(
        n11590) );
  OAI21_X1 U14610 ( .B1(n11842), .B2(n11591), .A(n11590), .ZN(n11598) );
  INV_X1 U14611 ( .A(n11593), .ZN(n11595) );
  INV_X1 U14612 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11594) );
  NAND2_X1 U14613 ( .A1(n11595), .A2(n11594), .ZN(n11596) );
  NAND2_X1 U14614 ( .A1(n11631), .A2(n11596), .ZN(n15859) );
  OR2_X1 U14615 ( .A1(n15859), .A2(n11845), .ZN(n11597) );
  NAND2_X1 U14616 ( .A1(n14047), .A2(n10261), .ZN(n14030) );
  AOI22_X1 U14617 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11602) );
  AOI22_X1 U14618 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11615), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11601) );
  AOI22_X1 U14619 ( .A1(n11652), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11651), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U14620 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11460), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11599) );
  NAND4_X1 U14621 ( .A1(n11602), .A2(n11601), .A3(n11600), .A4(n11599), .ZN(
        n11608) );
  AOI22_X1 U14622 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11800), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11606) );
  AOI22_X1 U14623 ( .A1(n9751), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U14624 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11638), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U14625 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11603) );
  NAND4_X1 U14626 ( .A1(n11606), .A2(n11605), .A3(n11604), .A4(n11603), .ZN(
        n11607) );
  NOR2_X1 U14627 ( .A1(n11608), .A2(n11607), .ZN(n11612) );
  NAND2_X1 U14628 ( .A1(n11307), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11609) );
  NAND2_X1 U14629 ( .A1(n11845), .A2(n11609), .ZN(n11610) );
  AOI21_X1 U14630 ( .B1(n11847), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11610), .ZN(
        n11611) );
  OAI21_X1 U14631 ( .B1(n11842), .B2(n11612), .A(n11611), .ZN(n11614) );
  XNOR2_X1 U14632 ( .A(n11631), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14384) );
  NAND2_X1 U14633 ( .A1(n14384), .A2(n11914), .ZN(n11613) );
  NAND2_X1 U14634 ( .A1(n11614), .A2(n11613), .ZN(n14032) );
  AOI22_X1 U14635 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11619) );
  AOI22_X1 U14636 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U14637 ( .A1(n11652), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U14638 ( .A1(n11460), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11616) );
  NAND4_X1 U14639 ( .A1(n11619), .A2(n11618), .A3(n11617), .A4(n11616), .ZN(
        n11625) );
  AOI22_X1 U14640 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11644), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11623) );
  AOI22_X1 U14641 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U14642 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11638), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11621) );
  AOI22_X1 U14643 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11620) );
  NAND4_X1 U14644 ( .A1(n11623), .A2(n11622), .A3(n11621), .A4(n11620), .ZN(
        n11624) );
  NOR2_X1 U14645 ( .A1(n11625), .A2(n11624), .ZN(n11629) );
  NAND2_X1 U14646 ( .A1(n11307), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11626) );
  NAND2_X1 U14647 ( .A1(n11845), .A2(n11626), .ZN(n11627) );
  AOI21_X1 U14648 ( .B1(n11847), .B2(P1_EAX_REG_22__SCAN_IN), .A(n11627), .ZN(
        n11628) );
  OAI21_X1 U14649 ( .B1(n11842), .B2(n11629), .A(n11628), .ZN(n11634) );
  INV_X1 U14650 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14382) );
  INV_X1 U14651 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14022) );
  OAI21_X1 U14652 ( .B1(n11631), .B2(n14382), .A(n14022), .ZN(n11632) );
  NAND2_X1 U14653 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11630) );
  NAND2_X1 U14654 ( .A1(n11632), .A2(n11636), .ZN(n14368) );
  INV_X1 U14655 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n21122) );
  NAND2_X1 U14656 ( .A1(n11636), .A2(n21122), .ZN(n11637) );
  NAND2_X1 U14657 ( .A1(n11692), .A2(n11637), .ZN(n14363) );
  INV_X1 U14658 ( .A(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11812) );
  INV_X1 U14659 ( .A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11814) );
  INV_X1 U14660 ( .A(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11826) );
  OAI22_X1 U14661 ( .A1(n11703), .A2(n11814), .B1(n11700), .B2(n11826), .ZN(
        n11641) );
  INV_X1 U14662 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11816) );
  INV_X1 U14663 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11639) );
  OAI22_X1 U14664 ( .A1(n11827), .A2(n11816), .B1(n11825), .B2(n11639), .ZN(
        n11640) );
  AOI211_X1 U14665 ( .C1(n11121), .C2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n11641), .B(n11640), .ZN(n11643) );
  AOI22_X1 U14666 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11642) );
  OAI211_X1 U14667 ( .C1(n11232), .C2(n11812), .A(n11643), .B(n11642), .ZN(
        n11650) );
  AOI22_X1 U14668 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11615), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11648) );
  AOI22_X1 U14669 ( .A1(n9751), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11794), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11647) );
  AOI22_X1 U14670 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11800), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14671 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11645) );
  NAND4_X1 U14672 ( .A1(n11648), .A2(n11647), .A3(n11646), .A4(n11645), .ZN(
        n11649) );
  NOR2_X1 U14673 ( .A1(n11650), .A2(n11649), .ZN(n11674) );
  INV_X1 U14674 ( .A(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11655) );
  AOI22_X1 U14675 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n11652), .B1(
        n11651), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11654) );
  NAND2_X1 U14676 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11653) );
  OAI211_X1 U14677 ( .C1(n11711), .C2(n11655), .A(n11654), .B(n11653), .ZN(
        n11656) );
  INV_X1 U14678 ( .A(n11656), .ZN(n11659) );
  AOI22_X1 U14679 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11638), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U14680 ( .A1(n11819), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11657) );
  NAND3_X1 U14681 ( .A1(n11659), .A2(n11658), .A3(n11657), .ZN(n11668) );
  INV_X1 U14682 ( .A(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11660) );
  INV_X1 U14683 ( .A(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n21097) );
  OAI22_X1 U14684 ( .A1(n11661), .A2(n11660), .B1(n9779), .B2(n21097), .ZN(
        n11662) );
  AOI21_X1 U14685 ( .B1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B2(n11767), .A(
        n11662), .ZN(n11666) );
  AOI22_X1 U14686 ( .A1(n11728), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11057), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11665) );
  AOI22_X1 U14687 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n11460), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11664) );
  NAND2_X1 U14688 ( .A1(n11527), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11663) );
  NAND4_X1 U14689 ( .A1(n11666), .A2(n11665), .A3(n11664), .A4(n11663), .ZN(
        n11667) );
  NOR2_X1 U14690 ( .A1(n11668), .A2(n11667), .ZN(n11675) );
  XOR2_X1 U14691 ( .A(n11674), .B(n11675), .Z(n11669) );
  NAND2_X1 U14692 ( .A1(n11669), .A2(n11806), .ZN(n11672) );
  OAI21_X1 U14693 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n21122), .A(n11845), 
        .ZN(n11670) );
  AOI21_X1 U14694 ( .B1(n11847), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11670), .ZN(
        n11671) );
  NAND2_X1 U14695 ( .A1(n11672), .A2(n11671), .ZN(n11673) );
  OAI21_X1 U14696 ( .B1(n11845), .B2(n14363), .A(n11673), .ZN(n14006) );
  NOR2_X1 U14697 ( .A1(n11675), .A2(n11674), .ZN(n11698) );
  AOI22_X1 U14698 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U14699 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11615), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U14700 ( .A1(n11794), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11677) );
  AOI22_X1 U14701 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11460), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11676) );
  NAND4_X1 U14702 ( .A1(n11679), .A2(n11678), .A3(n11677), .A4(n11676), .ZN(
        n11685) );
  AOI22_X1 U14703 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11800), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U14704 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11682) );
  AOI22_X1 U14705 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11638), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11681) );
  AOI22_X1 U14706 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11680) );
  NAND4_X1 U14707 ( .A1(n11683), .A2(n11682), .A3(n11681), .A4(n11680), .ZN(
        n11684) );
  OR2_X1 U14708 ( .A1(n11685), .A2(n11684), .ZN(n11697) );
  INV_X1 U14709 ( .A(n11697), .ZN(n11686) );
  XNOR2_X1 U14710 ( .A(n11698), .B(n11686), .ZN(n11691) );
  INV_X1 U14711 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n11688) );
  NAND2_X1 U14712 ( .A1(n11307), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11687) );
  OAI211_X1 U14713 ( .C1(n11689), .C2(n11688), .A(n11845), .B(n11687), .ZN(
        n11690) );
  AOI21_X1 U14714 ( .B1(n11691), .B2(n11806), .A(n11690), .ZN(n11695) );
  NAND2_X1 U14715 ( .A1(n11692), .A2(n13994), .ZN(n11693) );
  NAND2_X1 U14716 ( .A1(n11720), .A2(n11693), .ZN(n14356) );
  NOR2_X1 U14717 ( .A1(n14356), .A2(n11845), .ZN(n11694) );
  NAND2_X1 U14718 ( .A1(n11698), .A2(n11697), .ZN(n11726) );
  INV_X1 U14719 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11710) );
  INV_X1 U14720 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11701) );
  INV_X1 U14721 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11699) );
  OAI22_X1 U14722 ( .A1(n11815), .A2(n11701), .B1(n11700), .B2(n11699), .ZN(
        n11706) );
  INV_X1 U14723 ( .A(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11704) );
  INV_X1 U14724 ( .A(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11702) );
  OAI22_X1 U14725 ( .A1(n11827), .A2(n11704), .B1(n11703), .B2(n11702), .ZN(
        n11705) );
  AOI211_X1 U14726 ( .C1(n11120), .C2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n11706), .B(n11705), .ZN(n11709) );
  AOI22_X1 U14727 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11708) );
  OAI211_X1 U14728 ( .C1(n11711), .C2(n11710), .A(n11709), .B(n11708), .ZN(
        n11717) );
  AOI22_X1 U14729 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11615), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U14730 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11638), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11714) );
  AOI22_X1 U14731 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11057), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11713) );
  AOI22_X1 U14732 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11712) );
  NAND4_X1 U14733 ( .A1(n11715), .A2(n11714), .A3(n11713), .A4(n11712), .ZN(
        n11716) );
  NOR2_X1 U14734 ( .A1(n11717), .A2(n11716), .ZN(n11727) );
  XOR2_X1 U14735 ( .A(n11726), .B(n11727), .Z(n11718) );
  NAND2_X1 U14736 ( .A1(n11718), .A2(n11806), .ZN(n11722) );
  INV_X1 U14737 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14346) );
  NOR2_X1 U14738 ( .A1(n14346), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11719) );
  AOI211_X1 U14739 ( .C1(n11847), .C2(P1_EAX_REG_25__SCAN_IN), .A(n11914), .B(
        n11719), .ZN(n11721) );
  XOR2_X1 U14740 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B(n11723), .Z(
        n14350) );
  AOI22_X1 U14741 ( .A1(n11722), .A2(n11721), .B1(n11914), .B2(n14350), .ZN(
        n13978) );
  INV_X1 U14742 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13968) );
  NAND2_X1 U14743 ( .A1(n11724), .A2(n13968), .ZN(n11725) );
  NAND2_X1 U14744 ( .A1(n11760), .A2(n11725), .ZN(n14337) );
  NOR2_X1 U14745 ( .A1(n11727), .A2(n11726), .ZN(n11745) );
  AOI22_X1 U14746 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11733) );
  AOI22_X1 U14747 ( .A1(n11728), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11732) );
  AOI22_X1 U14748 ( .A1(n11794), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11731) );
  AOI22_X1 U14749 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11460), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11730) );
  NAND4_X1 U14750 ( .A1(n11733), .A2(n11732), .A3(n11731), .A4(n11730), .ZN(
        n11739) );
  AOI22_X1 U14751 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11057), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U14752 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11736) );
  AOI22_X1 U14753 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11638), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11735) );
  AOI22_X1 U14754 ( .A1(n9751), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(n9748), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11734) );
  NAND4_X1 U14755 ( .A1(n11737), .A2(n11736), .A3(n11735), .A4(n11734), .ZN(
        n11738) );
  OR2_X1 U14756 ( .A1(n11739), .A2(n11738), .ZN(n11744) );
  XNOR2_X1 U14757 ( .A(n11745), .B(n11744), .ZN(n11742) );
  AOI21_X1 U14758 ( .B1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n11307), .A(
        n11914), .ZN(n11741) );
  NAND2_X1 U14759 ( .A1(n11847), .A2(P1_EAX_REG_26__SCAN_IN), .ZN(n11740) );
  OAI211_X1 U14760 ( .C1(n11742), .C2(n11842), .A(n11741), .B(n11740), .ZN(
        n11743) );
  OAI21_X1 U14761 ( .B1(n11845), .B2(n14337), .A(n11743), .ZN(n13967) );
  NAND2_X1 U14762 ( .A1(n11745), .A2(n11744), .ZN(n11765) );
  AOI22_X1 U14763 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11057), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11749) );
  AOI22_X1 U14764 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11748) );
  AOI22_X1 U14765 ( .A1(n11794), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11638), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11747) );
  AOI22_X1 U14766 ( .A1(n11460), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11746) );
  NAND4_X1 U14767 ( .A1(n11749), .A2(n11748), .A3(n11747), .A4(n11746), .ZN(
        n11755) );
  AOI22_X1 U14768 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11753) );
  AOI22_X1 U14769 ( .A1(n11527), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11644), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11752) );
  AOI22_X1 U14770 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11651), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U14771 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11750) );
  NAND4_X1 U14772 ( .A1(n11753), .A2(n11752), .A3(n11751), .A4(n11750), .ZN(
        n11754) );
  NOR2_X1 U14773 ( .A1(n11755), .A2(n11754), .ZN(n11766) );
  XOR2_X1 U14774 ( .A(n11765), .B(n11766), .Z(n11756) );
  NAND2_X1 U14775 ( .A1(n11756), .A2(n11806), .ZN(n11759) );
  NOR2_X1 U14776 ( .A1(n14325), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11757) );
  AOI211_X1 U14777 ( .C1(n11847), .C2(P1_EAX_REG_27__SCAN_IN), .A(n11914), .B(
        n11757), .ZN(n11758) );
  XNOR2_X1 U14778 ( .A(n11760), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14329) );
  AOI22_X1 U14779 ( .A1(n11759), .A2(n11758), .B1(n11914), .B2(n14329), .ZN(
        n13953) );
  INV_X1 U14780 ( .A(n11761), .ZN(n11763) );
  INV_X1 U14781 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11762) );
  NAND2_X1 U14782 ( .A1(n11763), .A2(n11762), .ZN(n11764) );
  NAND2_X1 U14783 ( .A1(n11811), .A2(n11764), .ZN(n14318) );
  NOR2_X1 U14784 ( .A1(n11766), .A2(n11765), .ZN(n11783) );
  AOI22_X1 U14785 ( .A1(n11120), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11121), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11771) );
  AOI22_X1 U14786 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11615), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11770) );
  AOI22_X1 U14787 ( .A1(n11794), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11651), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11769) );
  AOI22_X1 U14788 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11460), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11768) );
  NAND4_X1 U14789 ( .A1(n11771), .A2(n11770), .A3(n11769), .A4(n11768), .ZN(
        n11777) );
  AOI22_X1 U14790 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11057), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U14791 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11774) );
  AOI22_X1 U14792 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11638), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11773) );
  AOI22_X1 U14793 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11772) );
  NAND4_X1 U14794 ( .A1(n11775), .A2(n11774), .A3(n11773), .A4(n11772), .ZN(
        n11776) );
  OR2_X1 U14795 ( .A1(n11777), .A2(n11776), .ZN(n11782) );
  XNOR2_X1 U14796 ( .A(n11783), .B(n11782), .ZN(n11780) );
  AOI21_X1 U14797 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n11307), .A(
        n11914), .ZN(n11779) );
  NAND2_X1 U14798 ( .A1(n11847), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n11778) );
  OAI211_X1 U14799 ( .C1(n11780), .C2(n11842), .A(n11779), .B(n11778), .ZN(
        n11781) );
  OAI21_X1 U14800 ( .B1(n11845), .B2(n14318), .A(n11781), .ZN(n13940) );
  NAND2_X1 U14801 ( .A1(n11783), .A2(n11782), .ZN(n11836) );
  INV_X1 U14802 ( .A(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11786) );
  AOI22_X1 U14803 ( .A1(n11460), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11785) );
  NAND2_X1 U14804 ( .A1(n11121), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11784) );
  OAI211_X1 U14805 ( .C1(n11787), .C2(n11786), .A(n11785), .B(n11784), .ZN(
        n11788) );
  INV_X1 U14806 ( .A(n11788), .ZN(n11793) );
  AOI22_X1 U14807 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11638), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11792) );
  AOI22_X1 U14808 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11791) );
  NAND3_X1 U14809 ( .A1(n11793), .A2(n11792), .A3(n11791), .ZN(n11805) );
  INV_X1 U14810 ( .A(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11797) );
  AOI22_X1 U14811 ( .A1(n11168), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11794), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11796) );
  NAND2_X1 U14812 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11795) );
  OAI211_X1 U14813 ( .C1(n11232), .C2(n11797), .A(n11796), .B(n11795), .ZN(
        n11798) );
  INV_X1 U14814 ( .A(n11798), .ZN(n11803) );
  AOI22_X1 U14815 ( .A1(n11644), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9751), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11802) );
  AOI22_X1 U14816 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11801) );
  NAND3_X1 U14817 ( .A1(n11803), .A2(n11802), .A3(n11801), .ZN(n11804) );
  NOR2_X1 U14818 ( .A1(n11805), .A2(n11804), .ZN(n11837) );
  XOR2_X1 U14819 ( .A(n11836), .B(n11837), .Z(n11807) );
  NAND2_X1 U14820 ( .A1(n11807), .A2(n11806), .ZN(n11810) );
  INV_X1 U14821 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14298) );
  NOR2_X1 U14822 ( .A1(n14298), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11808) );
  AOI211_X1 U14823 ( .C1(n11847), .C2(P1_EAX_REG_29__SCAN_IN), .A(n11914), .B(
        n11808), .ZN(n11809) );
  XNOR2_X1 U14824 ( .A(n11811), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14300) );
  AOI22_X1 U14825 ( .A1(n11810), .A2(n11809), .B1(n11914), .B2(n14300), .ZN(
        n13924) );
  INV_X1 U14826 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11917) );
  XNOR2_X1 U14827 ( .A(n11918), .B(n11917), .ZN(n14294) );
  OAI22_X1 U14828 ( .A1(n11815), .A2(n11814), .B1(n11813), .B2(n11812), .ZN(
        n11818) );
  NOR2_X1 U14829 ( .A1(n11232), .A2(n11816), .ZN(n11817) );
  AOI211_X1 U14830 ( .C1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .C2(n11800), .A(
        n11818), .B(n11817), .ZN(n11823) );
  AOI22_X1 U14831 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11644), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11822) );
  AOI22_X1 U14832 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11821) );
  NAND3_X1 U14833 ( .A1(n11823), .A2(n11822), .A3(n11821), .ZN(n11835) );
  INV_X1 U14834 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11824) );
  OAI22_X1 U14835 ( .A1(n11827), .A2(n11826), .B1(n11825), .B2(n11824), .ZN(
        n11828) );
  AOI21_X1 U14836 ( .B1(n11121), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n11828), .ZN(n11833) );
  AOI22_X1 U14837 ( .A1(n11615), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11168), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11832) );
  AOI22_X1 U14838 ( .A1(n11460), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11729), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11831) );
  NAND2_X1 U14839 ( .A1(n11829), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11830) );
  NAND4_X1 U14840 ( .A1(n11833), .A2(n11832), .A3(n11831), .A4(n11830), .ZN(
        n11834) );
  NOR2_X1 U14841 ( .A1(n11835), .A2(n11834), .ZN(n11839) );
  NOR2_X1 U14842 ( .A1(n11837), .A2(n11836), .ZN(n11838) );
  XOR2_X1 U14843 ( .A(n11839), .B(n11838), .Z(n11843) );
  AOI21_X1 U14844 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n11307), .A(
        n11914), .ZN(n11841) );
  NAND2_X1 U14845 ( .A1(n11847), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n11840) );
  OAI211_X1 U14846 ( .C1(n11843), .C2(n11842), .A(n11841), .B(n11840), .ZN(
        n11844) );
  OAI21_X1 U14847 ( .B1(n11845), .B2(n14294), .A(n11844), .ZN(n13913) );
  AOI22_X1 U14848 ( .A1(n11847), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n11846), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11848) );
  NAND2_X1 U14849 ( .A1(n20492), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11850) );
  NAND2_X1 U14850 ( .A1(n11027), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11849) );
  NAND2_X1 U14851 ( .A1(n11850), .A2(n11849), .ZN(n11857) );
  NAND2_X1 U14852 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20602), .ZN(
        n11863) );
  NAND2_X1 U14853 ( .A1(n20566), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11854) );
  NAND2_X1 U14854 ( .A1(n11038), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11851) );
  NAND2_X1 U14855 ( .A1(n11854), .A2(n11851), .ZN(n11875) );
  INV_X1 U14856 ( .A(n11875), .ZN(n11852) );
  XNOR2_X1 U14857 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11885) );
  AND2_X1 U14858 ( .A1(n11363), .A2(n11894), .ZN(n11855) );
  NOR2_X1 U14859 ( .A1(n20198), .A2(n20773), .ZN(n11856) );
  NAND2_X1 U14860 ( .A1(n12626), .A2(n20198), .ZN(n11862) );
  NAND2_X1 U14861 ( .A1(n11896), .A2(n11862), .ZN(n11861) );
  NAND2_X1 U14862 ( .A1(n11857), .A2(n11863), .ZN(n11858) );
  NAND2_X1 U14863 ( .A1(n11859), .A2(n11858), .ZN(n11910) );
  NAND2_X1 U14864 ( .A1(n11898), .A2(n11910), .ZN(n11860) );
  NAND2_X1 U14865 ( .A1(n11861), .A2(n11860), .ZN(n11870) );
  INV_X1 U14866 ( .A(n11870), .ZN(n11874) );
  AND2_X1 U14867 ( .A1(n12763), .A2(n11862), .ZN(n11880) );
  OAI21_X1 U14868 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20602), .A(
        n11863), .ZN(n11864) );
  INV_X1 U14869 ( .A(n11864), .ZN(n11865) );
  OAI211_X1 U14870 ( .C1(n9731), .C2(n11104), .A(n11880), .B(n11865), .ZN(
        n11868) );
  NAND2_X1 U14871 ( .A1(n11895), .A2(n11865), .ZN(n11866) );
  NAND2_X1 U14872 ( .A1(n11866), .A2(n11904), .ZN(n11867) );
  INV_X1 U14873 ( .A(n11871), .ZN(n11873) );
  OAI21_X1 U14874 ( .B1(n11896), .B2(n12626), .A(n11910), .ZN(n11869) );
  OAI21_X1 U14875 ( .B1(n11871), .B2(n11870), .A(n11869), .ZN(n11872) );
  OAI21_X1 U14876 ( .B1(n11874), .B2(n11873), .A(n11872), .ZN(n11884) );
  NAND2_X1 U14877 ( .A1(n11876), .A2(n11875), .ZN(n11878) );
  NAND2_X1 U14878 ( .A1(n11878), .A2(n11877), .ZN(n11909) );
  INV_X1 U14879 ( .A(n11909), .ZN(n11879) );
  NAND2_X1 U14880 ( .A1(n11895), .A2(n11879), .ZN(n11881) );
  OAI211_X1 U14881 ( .C1(n11879), .C2(n11889), .A(n11881), .B(n11880), .ZN(
        n11883) );
  NOR2_X1 U14882 ( .A1(n11881), .A2(n11880), .ZN(n11882) );
  AOI21_X1 U14883 ( .B1(n11884), .B2(n11883), .A(n11882), .ZN(n11892) );
  NOR2_X1 U14884 ( .A1(n11886), .A2(n11885), .ZN(n11887) );
  OR2_X1 U14885 ( .A1(n11888), .A2(n11887), .ZN(n11908) );
  AND2_X1 U14886 ( .A1(n11889), .A2(n11908), .ZN(n11891) );
  INV_X1 U14887 ( .A(n11908), .ZN(n11890) );
  OAI22_X1 U14888 ( .A1(n11892), .A2(n11891), .B1(n11890), .B2(n11904), .ZN(
        n11893) );
  OAI21_X1 U14889 ( .B1(n11898), .B2(n11911), .A(n11893), .ZN(n11903) );
  AOI222_X1 U14890 ( .A1(n11894), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .B1(n11894), .B2(n11363), .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .C2(n11363), .ZN(n11912) );
  NAND2_X1 U14891 ( .A1(n11912), .A2(n11895), .ZN(n11902) );
  NAND2_X1 U14892 ( .A1(n20773), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11901) );
  INV_X1 U14893 ( .A(n11911), .ZN(n11899) );
  INV_X1 U14894 ( .A(n11896), .ZN(n11897) );
  NAND4_X1 U14895 ( .A1(n11899), .A2(n11898), .A3(n11897), .A4(n9729), .ZN(
        n11900) );
  NAND4_X1 U14896 ( .A1(n11903), .A2(n11902), .A3(n11901), .A4(n11900), .ZN(
        n11907) );
  INV_X1 U14897 ( .A(n11904), .ZN(n11905) );
  NAND2_X1 U14898 ( .A1(n11912), .A2(n11905), .ZN(n11906) );
  NOR3_X1 U14899 ( .A1(n11910), .A2(n11909), .A3(n11908), .ZN(n11913) );
  OAI21_X1 U14900 ( .B1(n11913), .B2(n11912), .A(n11911), .ZN(n12968) );
  NAND2_X1 U14901 ( .A1(n12968), .A2(n9805), .ZN(n12618) );
  INV_X1 U14902 ( .A(n20859), .ZN(n16049) );
  NOR3_X1 U14903 ( .A1(n20773), .A2(n20573), .A3(n16049), .ZN(n15817) );
  AND2_X1 U14904 ( .A1(n20773), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12410) );
  NAND2_X1 U14905 ( .A1(n12410), .A2(n11914), .ZN(n11915) );
  NAND2_X1 U14906 ( .A1(n19990), .A2(n11915), .ZN(n11916) );
  INV_X1 U14907 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11919) );
  NOR2_X1 U14908 ( .A1(n13364), .A2(n20772), .ZN(n11921) );
  NAND2_X1 U14909 ( .A1(n12423), .A2(n19980), .ZN(n12035) );
  INV_X1 U14910 ( .A(n20189), .ZN(n11922) );
  INV_X2 U14911 ( .A(n11926), .ZN(n13909) );
  OR2_X2 U14912 ( .A1(n9731), .A2(n12626), .ZN(n11929) );
  AOI22_X1 U14913 ( .A1(n13006), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n11929), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U14914 ( .A1(n13006), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n11929), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13910) );
  INV_X1 U14915 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n14139) );
  NAND2_X1 U14916 ( .A1(n12004), .A2(n14139), .ZN(n11925) );
  INV_X1 U14917 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20973) );
  NAND2_X1 U14918 ( .A1(n12005), .A2(n20973), .ZN(n11923) );
  OAI211_X1 U14919 ( .C1(n11929), .C2(P1_EBX_REG_1__SCAN_IN), .A(n13909), .B(
        n11923), .ZN(n11924) );
  NAND2_X1 U14920 ( .A1(n11925), .A2(n11924), .ZN(n11930) );
  NAND2_X1 U14921 ( .A1(n12005), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n11928) );
  INV_X1 U14922 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13211) );
  NAND2_X1 U14923 ( .A1(n13909), .A2(n13211), .ZN(n11927) );
  NAND2_X1 U14924 ( .A1(n11928), .A2(n11927), .ZN(n13007) );
  XNOR2_X1 U14925 ( .A(n11930), .B(n13007), .ZN(n13192) );
  NAND2_X1 U14926 ( .A1(n13192), .A2(n13179), .ZN(n11931) );
  INV_X1 U14927 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13189) );
  NAND2_X1 U14928 ( .A1(n12004), .A2(n13189), .ZN(n11934) );
  INV_X1 U14929 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20156) );
  NAND2_X1 U14930 ( .A1(n12005), .A2(n20156), .ZN(n11932) );
  OAI211_X1 U14931 ( .C1(n11929), .C2(P1_EBX_REG_2__SCAN_IN), .A(n13909), .B(
        n11932), .ZN(n11933) );
  AND2_X1 U14932 ( .A1(n11934), .A2(n11933), .ZN(n13186) );
  MUX2_X1 U14933 ( .A(n12002), .B(n13909), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n11936) );
  OAI21_X1 U14934 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13006), .A(
        n11936), .ZN(n13234) );
  INV_X1 U14935 ( .A(n12005), .ZN(n11982) );
  MUX2_X1 U14936 ( .A(n12004), .B(n11982), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n11937) );
  INV_X1 U14937 ( .A(n11937), .ZN(n11940) );
  NAND2_X1 U14938 ( .A1(n11982), .A2(n11929), .ZN(n11985) );
  NAND2_X1 U14939 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11929), .ZN(
        n11938) );
  AND2_X1 U14940 ( .A1(n11985), .A2(n11938), .ZN(n11939) );
  NAND2_X1 U14941 ( .A1(n11940), .A2(n11939), .ZN(n16034) );
  NAND2_X1 U14942 ( .A1(n11959), .A2(n20008), .ZN(n11943) );
  NAND2_X1 U14943 ( .A1(n13909), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11941) );
  OAI211_X1 U14944 ( .C1(n11929), .C2(P1_EBX_REG_5__SCAN_IN), .A(n12005), .B(
        n11941), .ZN(n11942) );
  AND2_X1 U14945 ( .A1(n11943), .A2(n11942), .ZN(n16033) );
  INV_X1 U14946 ( .A(n12004), .ZN(n11994) );
  MUX2_X1 U14947 ( .A(n11994), .B(n12005), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n11946) );
  NAND2_X1 U14948 ( .A1(n11929), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11944) );
  AND2_X1 U14949 ( .A1(n11985), .A2(n11944), .ZN(n11945) );
  NAND2_X1 U14950 ( .A1(n11946), .A2(n11945), .ZN(n13418) );
  NAND2_X1 U14951 ( .A1(n16036), .A2(n13418), .ZN(n13469) );
  INV_X1 U14952 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13471) );
  NAND2_X1 U14953 ( .A1(n11959), .A2(n13471), .ZN(n11949) );
  NAND2_X1 U14954 ( .A1(n13909), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11947) );
  OAI211_X1 U14955 ( .C1(n11929), .C2(P1_EBX_REG_7__SCAN_IN), .A(n12005), .B(
        n11947), .ZN(n11948) );
  NAND2_X1 U14956 ( .A1(n11949), .A2(n11948), .ZN(n13468) );
  MUX2_X1 U14957 ( .A(n12004), .B(n11982), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n11952) );
  NAND2_X1 U14958 ( .A1(n11929), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11950) );
  NAND2_X1 U14959 ( .A1(n11985), .A2(n11950), .ZN(n11951) );
  NOR2_X1 U14960 ( .A1(n11952), .A2(n11951), .ZN(n13500) );
  INV_X1 U14961 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n13524) );
  NAND2_X1 U14962 ( .A1(n11959), .A2(n13524), .ZN(n11955) );
  NAND2_X1 U14963 ( .A1(n13909), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11953) );
  OAI211_X1 U14964 ( .C1(n11929), .C2(P1_EBX_REG_9__SCAN_IN), .A(n12005), .B(
        n11953), .ZN(n11954) );
  INV_X1 U14965 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14122) );
  NAND2_X1 U14966 ( .A1(n12004), .A2(n14122), .ZN(n11958) );
  INV_X1 U14967 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12514) );
  NAND2_X1 U14968 ( .A1(n12005), .A2(n12514), .ZN(n11956) );
  OAI211_X1 U14969 ( .C1(n11929), .C2(P1_EBX_REG_10__SCAN_IN), .A(n13909), .B(
        n11956), .ZN(n11957) );
  NAND2_X1 U14970 ( .A1(n11958), .A2(n11957), .ZN(n13536) );
  INV_X1 U14971 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15904) );
  NAND2_X1 U14972 ( .A1(n11959), .A2(n15904), .ZN(n11962) );
  NAND2_X1 U14973 ( .A1(n13909), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11960) );
  OAI211_X1 U14974 ( .C1(n11929), .C2(P1_EBX_REG_11__SCAN_IN), .A(n12005), .B(
        n11960), .ZN(n11961) );
  NAND2_X1 U14975 ( .A1(n11962), .A2(n11961), .ZN(n15890) );
  MUX2_X1 U14976 ( .A(n12004), .B(n11982), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n11965) );
  NAND2_X1 U14977 ( .A1(n11929), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11963) );
  NAND2_X1 U14978 ( .A1(n11985), .A2(n11963), .ZN(n11964) );
  NOR2_X1 U14979 ( .A1(n11965), .A2(n11964), .ZN(n14188) );
  MUX2_X1 U14980 ( .A(n12002), .B(n13909), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n11966) );
  OAI21_X1 U14981 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n13006), .A(
        n11966), .ZN(n14107) );
  INV_X1 U14982 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14183) );
  NAND2_X1 U14983 ( .A1(n12004), .A2(n14183), .ZN(n11969) );
  INV_X1 U14984 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15992) );
  NAND2_X1 U14985 ( .A1(n12005), .A2(n15992), .ZN(n11967) );
  OAI211_X1 U14986 ( .C1(n11929), .C2(P1_EBX_REG_14__SCAN_IN), .A(n13909), .B(
        n11967), .ZN(n11968) );
  NAND2_X1 U14987 ( .A1(n11969), .A2(n11968), .ZN(n14094) );
  MUX2_X1 U14988 ( .A(n12002), .B(n13909), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n11970) );
  OAI21_X1 U14989 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n13006), .A(
        n11970), .ZN(n14086) );
  MUX2_X1 U14990 ( .A(n12002), .B(n13909), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n11971) );
  OAI21_X1 U14991 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n13006), .A(
        n11971), .ZN(n11972) );
  INV_X1 U14992 ( .A(n11972), .ZN(n14068) );
  INV_X1 U14993 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n21002) );
  NAND2_X1 U14994 ( .A1(n12004), .A2(n21002), .ZN(n11975) );
  INV_X1 U14995 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15971) );
  NAND2_X1 U14996 ( .A1(n12005), .A2(n15971), .ZN(n11973) );
  OAI211_X1 U14997 ( .C1(n11929), .C2(P1_EBX_REG_16__SCAN_IN), .A(n13909), .B(
        n11973), .ZN(n11974) );
  NAND2_X1 U14998 ( .A1(n11975), .A2(n11974), .ZN(n15871) );
  INV_X1 U14999 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14179) );
  NAND2_X1 U15000 ( .A1(n12004), .A2(n14179), .ZN(n11978) );
  INV_X1 U15001 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14609) );
  NAND2_X1 U15002 ( .A1(n12005), .A2(n14609), .ZN(n11976) );
  OAI211_X1 U15003 ( .C1(n11929), .C2(P1_EBX_REG_18__SCAN_IN), .A(n13909), .B(
        n11976), .ZN(n11977) );
  NAND2_X1 U15004 ( .A1(n11978), .A2(n11977), .ZN(n14175) );
  NAND2_X1 U15005 ( .A1(n14176), .A2(n14175), .ZN(n14178) );
  MUX2_X1 U15006 ( .A(n12002), .B(n13909), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n11979) );
  OAI21_X1 U15007 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n13006), .A(
        n11979), .ZN(n14056) );
  OR2_X2 U15008 ( .A1(n14178), .A2(n14056), .ZN(n14170) );
  MUX2_X1 U15009 ( .A(n12002), .B(n13909), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n11980) );
  OAI21_X1 U15010 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n13006), .A(
        n11980), .ZN(n11981) );
  INV_X1 U15011 ( .A(n11981), .ZN(n14033) );
  MUX2_X1 U15012 ( .A(n12004), .B(n11982), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n11983) );
  INV_X1 U15013 ( .A(n11983), .ZN(n11987) );
  NAND2_X1 U15014 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n11929), .ZN(
        n11984) );
  AND2_X1 U15015 ( .A1(n11985), .A2(n11984), .ZN(n11986) );
  NAND2_X1 U15016 ( .A1(n11987), .A2(n11986), .ZN(n14169) );
  NAND2_X1 U15017 ( .A1(n14033), .A2(n14169), .ZN(n11988) );
  INV_X1 U15018 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14167) );
  NAND2_X1 U15019 ( .A1(n12004), .A2(n14167), .ZN(n11991) );
  INV_X1 U15020 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14567) );
  NAND2_X1 U15021 ( .A1(n12005), .A2(n14567), .ZN(n11989) );
  OAI211_X1 U15022 ( .C1(n11929), .C2(P1_EBX_REG_22__SCAN_IN), .A(n13909), .B(
        n11989), .ZN(n11990) );
  NAND2_X1 U15023 ( .A1(n11991), .A2(n11990), .ZN(n14019) );
  MUX2_X1 U15024 ( .A(n12002), .B(n13909), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n11992) );
  OAI21_X1 U15025 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n13006), .A(
        n11992), .ZN(n11993) );
  INV_X1 U15026 ( .A(n11993), .ZN(n14003) );
  MUX2_X1 U15027 ( .A(n11994), .B(n12005), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n11996) );
  NAND2_X1 U15028 ( .A1(n11929), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11995) );
  AND2_X1 U15029 ( .A1(n11996), .A2(n11995), .ZN(n13998) );
  NAND2_X1 U15030 ( .A1(n13909), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11997) );
  OAI211_X1 U15031 ( .C1(n11929), .C2(P1_EBX_REG_25__SCAN_IN), .A(n12005), .B(
        n11997), .ZN(n11998) );
  OAI21_X1 U15032 ( .B1(n12002), .B2(P1_EBX_REG_25__SCAN_IN), .A(n11998), .ZN(
        n13979) );
  NOR2_X2 U15033 ( .A1(n9777), .A2(n13979), .ZN(n13980) );
  INV_X1 U15034 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14163) );
  NAND2_X1 U15035 ( .A1(n12004), .A2(n14163), .ZN(n12001) );
  INV_X1 U15036 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14512) );
  NAND2_X1 U15037 ( .A1(n12005), .A2(n14512), .ZN(n11999) );
  OAI211_X1 U15038 ( .C1(n11929), .C2(P1_EBX_REG_26__SCAN_IN), .A(n13909), .B(
        n11999), .ZN(n12000) );
  NAND2_X1 U15039 ( .A1(n12001), .A2(n12000), .ZN(n13963) );
  NAND2_X1 U15040 ( .A1(n13980), .A2(n13963), .ZN(n13965) );
  MUX2_X1 U15041 ( .A(n12002), .B(n13909), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12003) );
  OAI21_X1 U15042 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n13006), .A(
        n12003), .ZN(n13949) );
  INV_X1 U15043 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14161) );
  NAND2_X1 U15044 ( .A1(n12004), .A2(n14161), .ZN(n12008) );
  INV_X1 U15045 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14314) );
  NAND2_X1 U15046 ( .A1(n12005), .A2(n14314), .ZN(n12006) );
  OAI211_X1 U15047 ( .C1(n11929), .C2(P1_EBX_REG_28__SCAN_IN), .A(n13909), .B(
        n12006), .ZN(n12007) );
  AND2_X1 U15048 ( .A1(n12008), .A2(n12007), .ZN(n13936) );
  INV_X1 U15049 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14160) );
  NAND2_X1 U15050 ( .A1(n13179), .A2(n14160), .ZN(n12011) );
  OR2_X1 U15051 ( .A1(n13006), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12009) );
  NAND2_X1 U15052 ( .A1(n12011), .A2(n12009), .ZN(n13908) );
  MUX2_X1 U15053 ( .A(n13908), .B(n12011), .S(n11926), .Z(n13926) );
  MUX2_X1 U15054 ( .A(n13909), .B(n13910), .S(n13925), .Z(n12012) );
  XOR2_X1 U15055 ( .A(n12013), .B(n12012), .Z(n14472) );
  INV_X1 U15056 ( .A(n20854), .ZN(n12014) );
  INV_X1 U15057 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14157) );
  OR2_X1 U15058 ( .A1(n12626), .A2(n14157), .ZN(n12019) );
  INV_X1 U15059 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20649) );
  NAND2_X1 U15060 ( .A1(n20856), .A2(n20649), .ZN(n15812) );
  INV_X1 U15061 ( .A(n15812), .ZN(n12017) );
  NOR2_X1 U15062 ( .A1(n12019), .A2(n12017), .ZN(n12015) );
  OR2_X1 U15063 ( .A1(n12016), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n12966) );
  NAND2_X1 U15064 ( .A1(n12626), .A2(n12966), .ZN(n12969) );
  AND2_X1 U15065 ( .A1(n12969), .A2(n12017), .ZN(n12021) );
  INV_X1 U15066 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n14043) );
  INV_X1 U15067 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20814) );
  INV_X1 U15068 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n15976) );
  INV_X1 U15069 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20803) );
  INV_X1 U15070 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20928) );
  INV_X1 U15071 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20012) );
  NAND4_X1 U15072 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n20004)
         );
  NOR3_X1 U15073 ( .A1(n20928), .A2(n20012), .A3(n20004), .ZN(n19983) );
  NAND2_X1 U15074 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19983), .ZN(n14129) );
  NOR2_X1 U15075 ( .A1(n20803), .A2(n14129), .ZN(n14123) );
  NAND3_X1 U15076 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(n14123), .ZN(n14079) );
  NAND4_X1 U15077 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(P1_REIP_REG_12__SCAN_IN), .A4(P1_REIP_REG_11__SCAN_IN), .ZN(n14080) );
  NOR3_X1 U15078 ( .A1(n15976), .A2(n14079), .A3(n14080), .ZN(n15875) );
  NAND2_X1 U15079 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n15875), .ZN(n14067) );
  NOR2_X1 U15080 ( .A1(n20814), .A2(n14067), .ZN(n14051) );
  NAND4_X1 U15081 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .A3(P1_REIP_REG_18__SCAN_IN), .A4(n14051), .ZN(n14038) );
  NOR2_X1 U15082 ( .A1(n14043), .A2(n14038), .ZN(n12024) );
  NAND2_X1 U15083 ( .A1(n20005), .A2(n12024), .ZN(n14025) );
  NAND2_X1 U15084 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n12018) );
  NAND2_X1 U15085 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n13982) );
  NOR2_X1 U15086 ( .A1(n13997), .A2(n13982), .ZN(n13969) );
  NAND2_X1 U15087 ( .A1(n13969), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n13955) );
  INV_X1 U15088 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n13959) );
  INV_X1 U15089 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14316) );
  INV_X1 U15090 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20832) );
  NOR2_X1 U15091 ( .A1(n13929), .A2(n20832), .ZN(n13920) );
  INV_X1 U15092 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20836) );
  NAND3_X1 U15093 ( .A1(n13920), .A2(P1_REIP_REG_30__SCAN_IN), .A3(n20836), 
        .ZN(n12032) );
  INV_X1 U15094 ( .A(n12019), .ZN(n12020) );
  NOR2_X1 U15095 ( .A1(n12021), .A2(n12020), .ZN(n12022) );
  AOI22_X1 U15096 ( .A1(n20021), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20024), .ZN(n12031) );
  INV_X1 U15097 ( .A(n19982), .ZN(n20003) );
  NAND4_X1 U15098 ( .A1(n19982), .A2(n12024), .A3(P1_REIP_REG_23__SCAN_IN), 
        .A4(P1_REIP_REG_22__SCAN_IN), .ZN(n13992) );
  NOR2_X1 U15099 ( .A1(n13982), .A2(n13992), .ZN(n12025) );
  NAND2_X1 U15100 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n12025), .ZN(n12026) );
  NAND2_X1 U15101 ( .A1(n14112), .A2(n12026), .ZN(n13970) );
  NAND2_X1 U15102 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n12027) );
  NAND2_X1 U15103 ( .A1(n14112), .A2(n12027), .ZN(n12028) );
  AND2_X1 U15104 ( .A1(n13970), .A2(n12028), .ZN(n13941) );
  NAND2_X1 U15105 ( .A1(n14112), .A2(n20832), .ZN(n12029) );
  NAND2_X1 U15106 ( .A1(n13941), .A2(n12029), .ZN(n13914) );
  INV_X1 U15107 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14292) );
  AND2_X1 U15108 ( .A1(n14112), .A2(n14292), .ZN(n13919) );
  OAI21_X1 U15109 ( .B1(n13914), .B2(n13919), .A(P1_REIP_REG_31__SCAN_IN), 
        .ZN(n12030) );
  NAND3_X1 U15110 ( .A1(n12032), .A2(n12031), .A3(n12030), .ZN(n12033) );
  AOI21_X1 U15111 ( .B1(n14472), .B2(n20025), .A(n12033), .ZN(n12034) );
  NAND2_X1 U15112 ( .A1(n12035), .A2(n12034), .ZN(P1_U2809) );
  INV_X1 U15113 ( .A(n12038), .ZN(n12037) );
  XNOR2_X1 U15114 ( .A(n12039), .B(n12037), .ZN(n14908) );
  NAND2_X1 U15115 ( .A1(n14908), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14907) );
  NAND2_X1 U15116 ( .A1(n14907), .A2(n10266), .ZN(n12042) );
  XOR2_X1 U15117 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n12040), .Z(
        n12041) );
  XNOR2_X1 U15118 ( .A(n12042), .B(n12041), .ZN(n12339) );
  NAND2_X1 U15119 ( .A1(n12339), .A2(n19162), .ZN(n12050) );
  AOI21_X1 U15120 ( .B1(n14668), .B2(n12057), .A(n12052), .ZN(n14665) );
  NAND2_X1 U15121 ( .A1(n19000), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12376) );
  OAI21_X1 U15122 ( .B1(n16225), .B2(n14668), .A(n12376), .ZN(n12046) );
  NAND2_X1 U15123 ( .A1(n14730), .A2(n12043), .ZN(n12044) );
  NAND2_X1 U15124 ( .A1(n13572), .A2(n12044), .ZN(n14723) );
  NOR2_X1 U15125 ( .A1(n14723), .A2(n16211), .ZN(n12045) );
  AOI211_X1 U15126 ( .C1(n16217), .C2(n14665), .A(n12046), .B(n12045), .ZN(
        n12048) );
  OAI21_X1 U15127 ( .B1(n14905), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14900), .ZN(n12383) );
  OR2_X1 U15128 ( .A1(n12383), .A2(n19159), .ZN(n12047) );
  NAND2_X1 U15129 ( .A1(n12050), .A2(n12049), .ZN(P2_U2986) );
  INV_X1 U15130 ( .A(n12052), .ZN(n12054) );
  AOI21_X1 U15131 ( .B1(n10002), .B2(n12054), .A(n12053), .ZN(n16064) );
  AOI21_X1 U15132 ( .B1(n16078), .B2(n12056), .A(n10001), .ZN(n16076) );
  OR2_X1 U15133 ( .A1(n12058), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12059) );
  NAND2_X1 U15134 ( .A1(n12056), .A2(n12059), .ZN(n14917) );
  INV_X1 U15135 ( .A(n14917), .ZN(n16092) );
  AOI21_X1 U15136 ( .B1(n14927), .B2(n12061), .A(n12058), .ZN(n14930) );
  OAI21_X1 U15137 ( .B1(n9803), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n12061), .ZN(n14939) );
  INV_X1 U15138 ( .A(n14939), .ZN(n16114) );
  AOI21_X1 U15139 ( .B1(n9983), .B2(n12062), .A(n9803), .ZN(n16138) );
  OAI21_X1 U15140 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12063), .A(
        n12062), .ZN(n16153) );
  INV_X1 U15141 ( .A(n16153), .ZN(n15779) );
  AOI21_X1 U15142 ( .B1(n14960), .B2(n12090), .A(n12063), .ZN(n14962) );
  AOI21_X1 U15143 ( .B1(n12065), .B2(n9987), .A(n9754), .ZN(n18905) );
  AOI21_X1 U15144 ( .B1(n12085), .B2(n15019), .A(n12067), .ZN(n15022) );
  AOI21_X1 U15145 ( .B1(n16159), .B2(n12084), .A(n12069), .ZN(n18932) );
  AOI21_X1 U15146 ( .B1(n16174), .B2(n12083), .A(n12071), .ZN(n16167) );
  AOI21_X1 U15147 ( .B1(n16195), .B2(n12082), .A(n12073), .ZN(n18961) );
  AOI21_X1 U15148 ( .B1(n15041), .B2(n12081), .A(n12075), .ZN(n18972) );
  AOI21_X1 U15149 ( .B1(n16224), .B2(n12080), .A(n12077), .ZN(n19004) );
  AOI21_X1 U15150 ( .B1(n21074), .B2(n12079), .A(n12078), .ZN(n13845) );
  OAI22_X1 U15151 ( .A1(n16324), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n19043) );
  INV_X1 U15152 ( .A(n19043), .ZN(n13866) );
  INV_X1 U15153 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19195) );
  AOI22_X1 U15154 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19195), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16324), .ZN(n13865) );
  NOR2_X1 U15155 ( .A1(n13866), .A2(n13865), .ZN(n13864) );
  OAI21_X1 U15156 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n12079), .ZN(n13314) );
  NAND2_X1 U15157 ( .A1(n13864), .A2(n13314), .ZN(n13843) );
  NOR2_X1 U15158 ( .A1(n13845), .A2(n13843), .ZN(n13293) );
  OAI21_X1 U15159 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12078), .A(
        n12080), .ZN(n19151) );
  NAND2_X1 U15160 ( .A1(n13293), .A2(n19151), .ZN(n19001) );
  NOR2_X1 U15161 ( .A1(n19004), .A2(n19001), .ZN(n18988) );
  OAI21_X1 U15162 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n12077), .A(
        n12081), .ZN(n18989) );
  NAND2_X1 U15163 ( .A1(n18988), .A2(n18989), .ZN(n18971) );
  NOR2_X1 U15164 ( .A1(n18972), .A2(n18971), .ZN(n13305) );
  OAI21_X1 U15165 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n12075), .A(
        n12082), .ZN(n16209) );
  NAND2_X1 U15166 ( .A1(n13305), .A2(n16209), .ZN(n18960) );
  NOR2_X1 U15167 ( .A1(n18961), .A2(n18960), .ZN(n18952) );
  OAI21_X1 U15168 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12073), .A(
        n12083), .ZN(n18953) );
  NAND2_X1 U15169 ( .A1(n18952), .A2(n18953), .ZN(n14706) );
  NOR2_X1 U15170 ( .A1(n16167), .A2(n14706), .ZN(n14705) );
  OAI21_X1 U15171 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n12071), .A(
        n12084), .ZN(n18940) );
  NAND2_X1 U15172 ( .A1(n14705), .A2(n18940), .ZN(n18924) );
  NOR2_X1 U15173 ( .A1(n18932), .A2(n18924), .ZN(n18923) );
  OAI21_X1 U15174 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n12069), .A(
        n12085), .ZN(n15030) );
  NAND2_X1 U15175 ( .A1(n18923), .A2(n15030), .ZN(n12539) );
  NOR2_X1 U15176 ( .A1(n15022), .A2(n12539), .ZN(n18912) );
  OAI21_X1 U15177 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12067), .A(
        n12065), .ZN(n18913) );
  NAND2_X1 U15178 ( .A1(n18912), .A2(n18913), .ZN(n18904) );
  NOR2_X1 U15179 ( .A1(n18905), .A2(n18904), .ZN(n18889) );
  OAI21_X1 U15180 ( .B1(n9754), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n12086), .ZN(n18890) );
  AOI21_X1 U15181 ( .B1(n18889), .B2(n18890), .A(n12087), .ZN(n18882) );
  AOI21_X1 U15182 ( .B1(n14984), .B2(n12086), .A(n12091), .ZN(n18881) );
  OAI21_X1 U15183 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12091), .A(
        n12090), .ZN(n14973) );
  NOR2_X1 U15184 ( .A1(n14962), .A2(n12564), .ZN(n12563) );
  NOR2_X1 U15185 ( .A1(n16114), .A2(n16113), .ZN(n16112) );
  NOR2_X1 U15186 ( .A1(n9753), .A2(n16090), .ZN(n16077) );
  NOR2_X1 U15187 ( .A1(n16076), .A2(n16077), .ZN(n16075) );
  NOR2_X1 U15188 ( .A1(n9753), .A2(n16075), .ZN(n14666) );
  NOR2_X1 U15189 ( .A1(n14665), .A2(n14666), .ZN(n14664) );
  XNOR2_X1 U15190 ( .A(n12053), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16058) );
  INV_X1 U15191 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19441) );
  NAND4_X1 U15192 ( .A1(n19441), .A2(n16324), .A3(n19898), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19820) );
  NAND2_X1 U15193 ( .A1(n12092), .A2(n19021), .ZN(n12290) );
  OR2_X1 U15194 ( .A1(n18853), .A2(n12338), .ZN(n12283) );
  NAND2_X1 U15195 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n16328) );
  NAND2_X1 U15196 ( .A1(n19898), .A2(n16328), .ZN(n12284) );
  NAND2_X1 U15197 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n12284), .ZN(n12093) );
  INV_X1 U15198 ( .A(n12121), .ZN(n12095) );
  INV_X1 U15199 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n12101) );
  AOI22_X1 U15200 ( .A1(n12264), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12253), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12100) );
  AND2_X1 U15201 ( .A1(n10102), .A2(n19576), .ZN(n12096) );
  INV_X1 U15202 ( .A(n12097), .ZN(n12098) );
  NAND2_X1 U15203 ( .A1(n12225), .A2(n12098), .ZN(n12099) );
  OAI211_X1 U15204 ( .C1(n12121), .C2(n12101), .A(n12100), .B(n12099), .ZN(
        n13446) );
  INV_X1 U15205 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18870) );
  AOI21_X1 U15206 ( .B1(n13832), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12103) );
  NAND2_X1 U15207 ( .A1(n12851), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n12102) );
  OAI211_X1 U15208 ( .C1(n12121), .C2(n18870), .A(n12103), .B(n12102), .ZN(
        n12688) );
  MUX2_X1 U15209 ( .A(n19250), .B(n19933), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12106) );
  INV_X1 U15210 ( .A(n12104), .ZN(n12105) );
  NAND2_X1 U15211 ( .A1(n12105), .A2(n12253), .ZN(n12117) );
  AND2_X1 U15212 ( .A1(n12106), .A2(n12117), .ZN(n12107) );
  INV_X1 U15213 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19138) );
  INV_X1 U15214 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19843) );
  OAI222_X1 U15215 ( .A1(n12260), .A2(n19195), .B1(n9775), .B2(n19138), .C1(
        n12121), .C2(n19843), .ZN(n12113) );
  XNOR2_X1 U15216 ( .A(n12114), .B(n12113), .ZN(n12865) );
  OR2_X1 U15217 ( .A1(n12109), .A2(n12241), .ZN(n12112) );
  NAND2_X1 U15218 ( .A1(n12104), .A2(n19250), .ZN(n12110) );
  MUX2_X1 U15219 ( .A(n12110), .B(n19924), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12111) );
  NAND2_X1 U15220 ( .A1(n12112), .A2(n12111), .ZN(n12866) );
  NOR2_X1 U15221 ( .A1(n12114), .A2(n12113), .ZN(n12115) );
  NAND2_X1 U15222 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12116) );
  OAI211_X1 U15223 ( .C1(n12118), .C2(n12241), .A(n12117), .B(n12116), .ZN(
        n12119) );
  INV_X1 U15224 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19845) );
  OR2_X1 U15225 ( .A1(n12121), .A2(n19845), .ZN(n12123) );
  INV_X2 U15226 ( .A(n9775), .ZN(n12264) );
  AOI22_X1 U15227 ( .A1(n12264), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12253), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12122) );
  NAND2_X1 U15228 ( .A1(n12123), .A2(n12122), .ZN(n13017) );
  INV_X1 U15229 ( .A(n12124), .ZN(n12125) );
  INV_X1 U15230 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n13258) );
  AOI22_X1 U15231 ( .A1(n12253), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12128) );
  AOI22_X1 U15232 ( .A1(n12225), .A2(n12126), .B1(n12264), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n12127) );
  OAI211_X1 U15233 ( .C1(n12121), .C2(n13258), .A(n12128), .B(n12127), .ZN(
        n13079) );
  NAND2_X1 U15234 ( .A1(n13078), .A2(n13079), .ZN(n13136) );
  INV_X1 U15235 ( .A(n12129), .ZN(n12132) );
  NAND2_X1 U15236 ( .A1(n12264), .A2(P2_EAX_REG_4__SCAN_IN), .ZN(n12131) );
  NAND2_X1 U15237 ( .A1(n12253), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12130) );
  OAI211_X1 U15238 ( .C1(n12241), .C2(n12132), .A(n12131), .B(n12130), .ZN(
        n12133) );
  AOI21_X1 U15239 ( .B1(n12095), .B2(P2_REIP_REG_4__SCAN_IN), .A(n12133), .ZN(
        n13137) );
  AOI222_X1 U15240 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n12095), .B1(n12253), 
        .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(P2_EAX_REG_6__SCAN_IN), 
        .C2(n12264), .ZN(n12692) );
  INV_X1 U15241 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19123) );
  INV_X1 U15242 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19853) );
  OAI222_X1 U15243 ( .A1(n16245), .A2(n12260), .B1(n9775), .B2(n19123), .C1(
        n12121), .C2(n19853), .ZN(n12751) );
  AOI22_X1 U15244 ( .A1(n13647), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9728), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12138) );
  AOI22_X1 U15245 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10575), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12137) );
  AOI22_X1 U15246 ( .A1(n13652), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12136) );
  AOI22_X1 U15247 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10540), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12135) );
  NAND4_X1 U15248 ( .A1(n12138), .A2(n12137), .A3(n12136), .A4(n12135), .ZN(
        n12144) );
  AOI22_X1 U15249 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13622), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12142) );
  AOI22_X1 U15250 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U15251 ( .A1(n12959), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12140) );
  AOI22_X1 U15252 ( .A1(n10582), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12139) );
  NAND4_X1 U15253 ( .A1(n12142), .A2(n12141), .A3(n12140), .A4(n12139), .ZN(
        n12143) );
  INV_X1 U15254 ( .A(n13050), .ZN(n12147) );
  NAND2_X1 U15255 ( .A1(n12264), .A2(P2_EAX_REG_8__SCAN_IN), .ZN(n12146) );
  NAND2_X1 U15256 ( .A1(n12253), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12145) );
  OAI211_X1 U15257 ( .C1(n12241), .C2(n12147), .A(n12146), .B(n12145), .ZN(
        n12148) );
  AOI21_X1 U15258 ( .B1(n12095), .B2(P2_REIP_REG_8__SCAN_IN), .A(n12148), .ZN(
        n12924) );
  NOR2_X2 U15259 ( .A1(n12923), .A2(n12924), .ZN(n12938) );
  INV_X1 U15260 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n12161) );
  AOI22_X1 U15261 ( .A1(n12264), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12253), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12160) );
  AOI22_X1 U15262 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12162), .B1(
        n10574), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U15263 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12959), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12151) );
  AOI22_X1 U15264 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10580), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12150) );
  AOI22_X1 U15265 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10582), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12149) );
  NAND4_X1 U15266 ( .A1(n12152), .A2(n12151), .A3(n12150), .A4(n12149), .ZN(
        n12158) );
  AOI22_X1 U15267 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n13652), .B1(
        n13647), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12156) );
  AOI22_X1 U15268 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10575), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12155) );
  AOI22_X1 U15269 ( .A1(n10540), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n10546), .ZN(n12154) );
  AOI22_X1 U15270 ( .A1(n9728), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13622), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12153) );
  NAND4_X1 U15271 ( .A1(n12156), .A2(n12155), .A3(n12154), .A4(n12153), .ZN(
        n12157) );
  NAND2_X1 U15272 ( .A1(n12225), .A2(n13113), .ZN(n12159) );
  OAI211_X1 U15273 ( .C1(n12121), .C2(n12161), .A(n12160), .B(n12159), .ZN(
        n12939) );
  AOI22_X1 U15274 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12162), .B1(
        n10574), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12166) );
  AOI22_X1 U15275 ( .A1(n13647), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n10546), .ZN(n12165) );
  AOI22_X1 U15276 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10575), .B1(
        n9728), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12164) );
  AOI22_X1 U15277 ( .A1(n13652), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10540), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12163) );
  NAND4_X1 U15278 ( .A1(n12166), .A2(n12165), .A3(n12164), .A4(n12163), .ZN(
        n12172) );
  AOI22_X1 U15279 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__2__SCAN_IN), .B2(n13622), .ZN(n12170) );
  AOI22_X1 U15280 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12169) );
  AOI22_X1 U15281 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10582), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12168) );
  AOI22_X1 U15282 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n12959), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12167) );
  NAND4_X1 U15283 ( .A1(n12170), .A2(n12169), .A3(n12168), .A4(n12167), .ZN(
        n12171) );
  AOI22_X1 U15284 ( .A1(n12264), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12253), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12173) );
  OAI21_X1 U15285 ( .B1(n13243), .B2(n12241), .A(n12173), .ZN(n12174) );
  AOI21_X1 U15286 ( .B1(P2_REIP_REG_10__SCAN_IN), .B2(n12095), .A(n12174), 
        .ZN(n13037) );
  INV_X1 U15287 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n12187) );
  AOI22_X1 U15288 ( .A1(n12264), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12253), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12186) );
  AOI22_X1 U15289 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12162), .B1(
        n10574), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12178) );
  AOI22_X1 U15290 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12959), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12177) );
  AOI22_X1 U15291 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10580), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12176) );
  AOI22_X1 U15292 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10582), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12175) );
  NAND4_X1 U15293 ( .A1(n12178), .A2(n12177), .A3(n12176), .A4(n12175), .ZN(
        n12184) );
  AOI22_X1 U15294 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n13652), .B1(
        n13647), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12182) );
  AOI22_X1 U15295 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10575), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15296 ( .A1(n10540), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n10546), .ZN(n12180) );
  AOI22_X1 U15297 ( .A1(n9728), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13622), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12179) );
  NAND4_X1 U15298 ( .A1(n12182), .A2(n12181), .A3(n12180), .A4(n12179), .ZN(
        n12183) );
  NAND2_X1 U15299 ( .A1(n12225), .A2(n13227), .ZN(n12185) );
  OAI211_X1 U15300 ( .C1(n12121), .C2(n12187), .A(n12186), .B(n12185), .ZN(
        n13061) );
  AOI22_X1 U15301 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13652), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12191) );
  AOI22_X1 U15302 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10575), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U15303 ( .A1(n10540), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n10546), .ZN(n12189) );
  AOI22_X1 U15304 ( .A1(n9728), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13622), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12188) );
  NAND4_X1 U15305 ( .A1(n12191), .A2(n12190), .A3(n12189), .A4(n12188), .ZN(
        n12197) );
  AOI22_X1 U15306 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13647), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U15307 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12959), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U15308 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10580), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12193) );
  AOI22_X1 U15309 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10582), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12192) );
  NAND4_X1 U15310 ( .A1(n12195), .A2(n12194), .A3(n12193), .A4(n12192), .ZN(
        n12196) );
  AOI22_X1 U15311 ( .A1(n12264), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12253), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12198) );
  OAI21_X1 U15312 ( .B1(n9913), .B2(n12241), .A(n12198), .ZN(n12199) );
  AOI21_X1 U15313 ( .B1(P2_REIP_REG_12__SCAN_IN), .B2(n12095), .A(n12199), 
        .ZN(n13088) );
  INV_X1 U15314 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n15283) );
  OR2_X1 U15315 ( .A1(n12121), .A2(n15283), .ZN(n12214) );
  AOI22_X1 U15316 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10574), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U15317 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12959), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12202) );
  AOI22_X1 U15318 ( .A1(n10580), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12201) );
  AOI22_X1 U15319 ( .A1(n10582), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12200) );
  NAND4_X1 U15320 ( .A1(n12203), .A2(n12202), .A3(n12201), .A4(n12200), .ZN(
        n12209) );
  AOI22_X1 U15321 ( .A1(n13647), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13652), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12207) );
  AOI22_X1 U15322 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10575), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12206) );
  AOI22_X1 U15323 ( .A1(n10540), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12205) );
  AOI22_X1 U15324 ( .A1(n9728), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13622), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12204) );
  NAND4_X1 U15325 ( .A1(n12207), .A2(n12206), .A3(n12205), .A4(n12204), .ZN(
        n12208) );
  NAND2_X1 U15326 ( .A1(n12264), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n12211) );
  NAND2_X1 U15327 ( .A1(n12253), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12210) );
  OAI211_X1 U15328 ( .C1(n12241), .C2(n13350), .A(n12211), .B(n12210), .ZN(
        n12212) );
  INV_X1 U15329 ( .A(n12212), .ZN(n12213) );
  NAND2_X1 U15330 ( .A1(n12214), .A2(n12213), .ZN(n13209) );
  INV_X1 U15331 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19864) );
  AOI22_X1 U15332 ( .A1(n12264), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12253), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12227) );
  AOI22_X1 U15333 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12162), .B1(
        n10574), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12218) );
  AOI22_X1 U15334 ( .A1(n13647), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n10546), .ZN(n12217) );
  AOI22_X1 U15335 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n13652), .B1(
        n13621), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12216) );
  AOI22_X1 U15336 ( .A1(n10575), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10540), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12215) );
  NAND4_X1 U15337 ( .A1(n12218), .A2(n12217), .A3(n12216), .A4(n12215), .ZN(
        n12224) );
  AOI22_X1 U15338 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n13622), .ZN(n12222) );
  AOI22_X1 U15339 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12221) );
  AOI22_X1 U15340 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10582), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12220) );
  AOI22_X1 U15341 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n12959), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12219) );
  NAND4_X1 U15342 ( .A1(n12222), .A2(n12221), .A3(n12220), .A4(n12219), .ZN(
        n12223) );
  NAND2_X1 U15343 ( .A1(n12225), .A2(n9820), .ZN(n12226) );
  OAI211_X1 U15344 ( .C1(n12121), .C2(n19864), .A(n12227), .B(n12226), .ZN(
        n13220) );
  AOI22_X1 U15345 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12162), .B1(
        n10574), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12231) );
  AOI22_X1 U15346 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12959), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12230) );
  AOI22_X1 U15347 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10580), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12229) );
  AOI22_X1 U15348 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10582), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12228) );
  NAND4_X1 U15349 ( .A1(n12231), .A2(n12230), .A3(n12229), .A4(n12228), .ZN(
        n12237) );
  AOI22_X1 U15350 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n13652), .B1(
        n13647), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12235) );
  AOI22_X1 U15351 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10575), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12234) );
  AOI22_X1 U15352 ( .A1(n10540), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n10546), .ZN(n12233) );
  AOI22_X1 U15353 ( .A1(n9728), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13622), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12232) );
  NAND4_X1 U15354 ( .A1(n12235), .A2(n12234), .A3(n12233), .A4(n12232), .ZN(
        n12236) );
  INV_X1 U15355 ( .A(n13463), .ZN(n12240) );
  NAND2_X1 U15356 ( .A1(n12264), .A2(P2_EAX_REG_15__SCAN_IN), .ZN(n12239) );
  NAND2_X1 U15357 ( .A1(n12253), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12238) );
  OAI211_X1 U15358 ( .C1(n12241), .C2(n12240), .A(n12239), .B(n12238), .ZN(
        n12242) );
  AOI21_X1 U15359 ( .B1(n12095), .B2(P2_REIP_REG_15__SCAN_IN), .A(n12242), 
        .ZN(n12544) );
  INV_X1 U15360 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n15235) );
  AOI22_X1 U15361 ( .A1(n12264), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12253), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12243) );
  OAI21_X1 U15362 ( .B1(n12121), .B2(n15235), .A(n12243), .ZN(n15231) );
  NAND2_X1 U15363 ( .A1(n15232), .A2(n15231), .ZN(n15234) );
  INV_X1 U15364 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n21170) );
  OR2_X1 U15365 ( .A1(n12121), .A2(n21170), .ZN(n12245) );
  AOI22_X1 U15366 ( .A1(n12264), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12253), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12244) );
  NAND2_X1 U15367 ( .A1(n12245), .A2(n12244), .ZN(n14880) );
  INV_X1 U15368 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19869) );
  OR2_X1 U15369 ( .A1(n12121), .A2(n19869), .ZN(n12248) );
  AOI22_X1 U15370 ( .A1(n12264), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12253), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12247) );
  INV_X1 U15371 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19871) );
  AOI22_X1 U15372 ( .A1(n12264), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12253), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12249) );
  OAI21_X1 U15373 ( .B1(n12121), .B2(n19871), .A(n12249), .ZN(n14873) );
  INV_X1 U15374 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n14972) );
  AOI22_X1 U15375 ( .A1(n12264), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12253), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12250) );
  OAI21_X1 U15376 ( .B1(n12121), .B2(n14972), .A(n12250), .ZN(n14696) );
  INV_X1 U15377 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19874) );
  OR2_X1 U15378 ( .A1(n12121), .A2(n19874), .ZN(n12252) );
  AOI22_X1 U15379 ( .A1(n12264), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12253), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12251) );
  NAND2_X1 U15380 ( .A1(n12252), .A2(n12251), .ZN(n12570) );
  INV_X1 U15381 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n12255) );
  AOI22_X1 U15382 ( .A1(n12264), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12253), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12254) );
  OAI21_X1 U15383 ( .B1(n12121), .B2(n12255), .A(n12254), .ZN(n15154) );
  INV_X1 U15384 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n21110) );
  AOI22_X1 U15385 ( .A1(n12264), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12253), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12256) );
  OAI21_X1 U15386 ( .B1(n12121), .B2(n21110), .A(n12256), .ZN(n12557) );
  AND2_X2 U15387 ( .A1(n15156), .A2(n12557), .ZN(n14852) );
  INV_X1 U15388 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n16106) );
  AOI22_X1 U15389 ( .A1(n12264), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12253), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12257) );
  OAI21_X1 U15390 ( .B1(n12121), .B2(n16106), .A(n12257), .ZN(n14851) );
  INV_X1 U15391 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n19089) );
  OAI22_X1 U15392 ( .A1(n9775), .A2(n19089), .B1(n21137), .B2(n12260), .ZN(
        n12258) );
  AOI21_X1 U15393 ( .B1(n12095), .B2(P2_REIP_REG_25__SCAN_IN), .A(n12258), 
        .ZN(n14680) );
  INV_X1 U15394 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n20996) );
  INV_X1 U15395 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15103) );
  OAI22_X1 U15396 ( .A1(n9775), .A2(n20996), .B1(n15103), .B2(n12260), .ZN(
        n12259) );
  AOI21_X1 U15397 ( .B1(n12095), .B2(P2_REIP_REG_26__SCAN_IN), .A(n12259), 
        .ZN(n14836) );
  INV_X1 U15398 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n19086) );
  OAI22_X1 U15399 ( .A1(n9775), .A2(n19086), .B1(n15088), .B2(n12260), .ZN(
        n12261) );
  AOI21_X1 U15400 ( .B1(n12095), .B2(P2_REIP_REG_27__SCAN_IN), .A(n12261), 
        .ZN(n14829) );
  INV_X1 U15401 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19882) );
  AOI22_X1 U15402 ( .A1(n12264), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12253), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12262) );
  OAI21_X1 U15403 ( .B1(n12121), .B2(n19882), .A(n12262), .ZN(n12369) );
  INV_X1 U15404 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19884) );
  AOI22_X1 U15405 ( .A1(n12264), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12253), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12263) );
  OAI21_X1 U15406 ( .B1(n12121), .B2(n19884), .A(n12263), .ZN(n14814) );
  INV_X1 U15407 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n12266) );
  AOI22_X1 U15408 ( .A1(n12264), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n12253), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12265) );
  OAI21_X1 U15409 ( .B1(n12121), .B2(n12266), .A(n12265), .ZN(n12267) );
  NAND2_X1 U15410 ( .A1(n12269), .A2(n12578), .ZN(n12633) );
  INV_X1 U15411 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19832) );
  NAND2_X1 U15412 ( .A1(n19832), .A2(n19842), .ZN(n19837) );
  INV_X1 U15413 ( .A(n19837), .ZN(n19824) );
  AOI211_X1 U15414 ( .C1(P2_STATE_REG_1__SCAN_IN), .C2(P2_STATE_REG_2__SCAN_IN), .A(P2_STATE_REG_0__SCAN_IN), .B(n19824), .ZN(n19828) );
  NAND2_X1 U15415 ( .A1(n19828), .A2(n16328), .ZN(n12293) );
  NOR2_X1 U15416 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n12293), .ZN(n16315) );
  INV_X1 U15417 ( .A(n16315), .ZN(n12275) );
  INV_X2 U15418 ( .A(n19015), .ZN(n19029) );
  NOR3_X1 U15419 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n12270), .A3(n19576), 
        .ZN(n16325) );
  NOR2_X1 U15420 ( .A1(n19021), .A2(n16325), .ZN(n12271) );
  AND2_X1 U15421 ( .A1(n16226), .A2(n12271), .ZN(n12272) );
  AOI22_X1 U15422 ( .A1(n19025), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18996), .ZN(n12278) );
  INV_X1 U15423 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n14718) );
  NAND2_X1 U15424 ( .A1(n12284), .A2(n14718), .ZN(n12273) );
  OR2_X1 U15425 ( .A1(n12633), .A2(n12273), .ZN(n12274) );
  NAND2_X1 U15426 ( .A1(n19073), .A2(n12274), .ZN(n12276) );
  NAND2_X1 U15427 ( .A1(n19026), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12277) );
  OAI211_X1 U15428 ( .C1(n15067), .C2(n19029), .A(n12278), .B(n12277), .ZN(
        n12279) );
  AOI21_X1 U15429 ( .B1(n12280), .B2(n19032), .A(n12279), .ZN(n12288) );
  OAI21_X1 U15430 ( .B1(n13573), .B2(n12282), .A(n12281), .ZN(n14891) );
  INV_X1 U15431 ( .A(n12283), .ZN(n12286) );
  INV_X1 U15432 ( .A(n12284), .ZN(n12285) );
  NAND2_X1 U15433 ( .A1(n12290), .A2(n12289), .ZN(P2_U2825) );
  INV_X1 U15434 ( .A(n12291), .ZN(n12336) );
  NOR2_X1 U15435 ( .A1(n16291), .A2(n19834), .ZN(n12662) );
  MUX2_X1 U15436 ( .A(n12292), .B(n19223), .S(n16316), .Z(n12307) );
  INV_X1 U15437 ( .A(n16291), .ZN(n12584) );
  INV_X1 U15438 ( .A(n12293), .ZN(n12660) );
  AND3_X1 U15439 ( .A1(n12292), .A2(n12584), .A3(n12660), .ZN(n12306) );
  NAND2_X1 U15440 ( .A1(n12295), .A2(n12294), .ZN(n12296) );
  NAND2_X1 U15441 ( .A1(n16302), .A2(n12296), .ZN(n12304) );
  NAND2_X1 U15442 ( .A1(n12297), .A2(n19250), .ZN(n12299) );
  NAND2_X1 U15443 ( .A1(n12299), .A2(n12298), .ZN(n12350) );
  AOI21_X1 U15444 ( .B1(n12300), .B2(n19212), .A(n19223), .ZN(n12301) );
  OAI21_X1 U15445 ( .B1(n12302), .B2(n13832), .A(n12301), .ZN(n12303) );
  NAND4_X1 U15446 ( .A1(n12305), .A2(n12304), .A3(n12350), .A4(n12303), .ZN(
        n12358) );
  OR2_X1 U15447 ( .A1(n12306), .A2(n12358), .ZN(n12665) );
  AOI21_X1 U15448 ( .B1(n12662), .B2(n12307), .A(n12665), .ZN(n12335) );
  NAND2_X1 U15449 ( .A1(n12308), .A2(n12338), .ZN(n12325) );
  NAND2_X1 U15450 ( .A1(n19212), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19077) );
  NAND2_X1 U15451 ( .A1(n19077), .A2(n13832), .ZN(n12309) );
  MUX2_X1 U15452 ( .A(n12338), .B(n12309), .S(n12317), .Z(n12319) );
  OAI211_X1 U15453 ( .C1(n13832), .C2(n12311), .A(n16300), .B(n12310), .ZN(
        n12316) );
  OAI21_X1 U15454 ( .B1(n12314), .B2(n10724), .A(n12313), .ZN(n12315) );
  OAI211_X1 U15455 ( .C1(n12674), .C2(n12317), .A(n12316), .B(n12315), .ZN(
        n12318) );
  NAND2_X1 U15456 ( .A1(n12319), .A2(n12318), .ZN(n12321) );
  NAND2_X1 U15457 ( .A1(n12321), .A2(n12320), .ZN(n12324) );
  OAI21_X1 U15458 ( .B1(n12322), .B2(n12338), .A(n12328), .ZN(n12323) );
  AOI21_X1 U15459 ( .B1(n12325), .B2(n12324), .A(n12323), .ZN(n12326) );
  MUX2_X1 U15460 ( .A(n21098), .B(n12326), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n12327) );
  INV_X1 U15461 ( .A(n19072), .ZN(n12332) );
  AOI21_X1 U15462 ( .B1(n12330), .B2(n16300), .A(n19234), .ZN(n12331) );
  NAND2_X1 U15463 ( .A1(n12332), .A2(n12331), .ZN(n12334) );
  NAND3_X1 U15464 ( .A1(n19072), .A2(n19223), .A3(n12660), .ZN(n12333) );
  NAND4_X1 U15465 ( .A1(n12336), .A2(n12335), .A3(n12334), .A4(n12333), .ZN(
        n12337) );
  NOR2_X1 U15466 ( .A1(n10721), .A2(n12338), .ZN(n19938) );
  NAND2_X1 U15467 ( .A1(n12339), .A2(n19182), .ZN(n12387) );
  NAND2_X1 U15468 ( .A1(n19223), .A2(n19212), .ZN(n12341) );
  OAI21_X1 U15469 ( .B1(n19234), .B2(n12661), .A(n12341), .ZN(n12342) );
  INV_X1 U15470 ( .A(n12342), .ZN(n12348) );
  INV_X1 U15471 ( .A(n10394), .ZN(n12676) );
  OAI21_X1 U15472 ( .B1(n12676), .B2(n12343), .A(n12661), .ZN(n12345) );
  NAND2_X1 U15473 ( .A1(n12345), .A2(n12344), .ZN(n12346) );
  AND3_X1 U15474 ( .A1(n12348), .A2(n12347), .A3(n12346), .ZN(n12353) );
  NAND2_X1 U15475 ( .A1(n12349), .A2(n13832), .ZN(n13288) );
  NAND2_X1 U15476 ( .A1(n13288), .A2(n12350), .ZN(n12351) );
  NAND2_X1 U15477 ( .A1(n12351), .A2(n19227), .ZN(n12352) );
  NAND2_X1 U15478 ( .A1(n12353), .A2(n12352), .ZN(n15358) );
  OR2_X1 U15479 ( .A1(n15358), .A2(n12848), .ZN(n12354) );
  NAND2_X1 U15480 ( .A1(n12382), .A2(n12354), .ZN(n15226) );
  INV_X1 U15481 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19194) );
  NOR2_X1 U15482 ( .A1(n19194), .A2(n19195), .ZN(n19193) );
  OR2_X1 U15483 ( .A1(n15226), .A2(n19193), .ZN(n12355) );
  OR2_X1 U15484 ( .A1(n12382), .A2(n16243), .ZN(n16262) );
  NAND2_X1 U15485 ( .A1(n12356), .A2(n16316), .ZN(n12357) );
  NAND2_X1 U15486 ( .A1(n12382), .A2(n16295), .ZN(n19175) );
  OR2_X1 U15487 ( .A1(n15226), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19176) );
  NAND2_X1 U15488 ( .A1(n19186), .A2(n19176), .ZN(n13279) );
  NOR2_X1 U15489 ( .A1(n13449), .A2(n13445), .ZN(n13444) );
  INV_X1 U15490 ( .A(n13444), .ZN(n15350) );
  NOR3_X1 U15491 ( .A1(n21153), .A2(n15354), .A3(n15350), .ZN(n15338) );
  AND3_X1 U15492 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n15338), .ZN(n12371) );
  INV_X1 U15493 ( .A(n19193), .ZN(n19177) );
  NAND2_X1 U15494 ( .A1(n19185), .A2(n19177), .ZN(n19174) );
  AND2_X1 U15495 ( .A1(n12371), .A2(n19174), .ZN(n12359) );
  NOR2_X1 U15496 ( .A1(n19192), .A2(n12359), .ZN(n12360) );
  INV_X1 U15497 ( .A(n15330), .ZN(n15308) );
  AND2_X1 U15498 ( .A1(n12372), .A2(n15308), .ZN(n15133) );
  AND2_X1 U15499 ( .A1(n15134), .A2(n15133), .ZN(n12361) );
  OR2_X1 U15500 ( .A1(n15307), .A2(n12361), .ZN(n15123) );
  OR2_X1 U15501 ( .A1(n15307), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12362) );
  NAND2_X1 U15502 ( .A1(n15123), .A2(n12362), .ZN(n15116) );
  INV_X1 U15503 ( .A(n15116), .ZN(n15104) );
  AND2_X1 U15504 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12373) );
  OR2_X1 U15505 ( .A1(n19192), .A2(n12373), .ZN(n12363) );
  NAND2_X1 U15506 ( .A1(n15104), .A2(n12363), .ZN(n15094) );
  INV_X1 U15507 ( .A(n16293), .ZN(n12955) );
  NAND2_X1 U15508 ( .A1(n16292), .A2(n13832), .ZN(n12366) );
  NAND2_X1 U15509 ( .A1(n12955), .A2(n12366), .ZN(n12367) );
  INV_X1 U15510 ( .A(n14815), .ZN(n12368) );
  OAI21_X1 U15511 ( .B1(n14828), .B2(n12369), .A(n12368), .ZN(n14822) );
  INV_X1 U15512 ( .A(n19174), .ZN(n13280) );
  OR2_X1 U15513 ( .A1(n19175), .A2(n13280), .ZN(n16252) );
  NAND2_X1 U15514 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19193), .ZN(
        n19172) );
  OR2_X1 U15515 ( .A1(n15226), .A2(n19172), .ZN(n12370) );
  NAND2_X1 U15516 ( .A1(n16252), .A2(n12370), .ZN(n15337) );
  NAND2_X1 U15517 ( .A1(n12372), .A2(n15329), .ZN(n15152) );
  INV_X1 U15518 ( .A(n15152), .ZN(n15138) );
  NAND2_X1 U15519 ( .A1(n15134), .A2(n15138), .ZN(n15125) );
  NOR2_X1 U15520 ( .A1(n15125), .A2(n15124), .ZN(n15110) );
  NAND2_X1 U15521 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15077) );
  NAND3_X1 U15522 ( .A1(n15089), .A2(n15077), .A3(n12374), .ZN(n12375) );
  OAI211_X1 U15523 ( .C1(n16251), .C2(n14822), .A(n12376), .B(n12375), .ZN(
        n12381) );
  NAND2_X1 U15524 ( .A1(n13859), .A2(n16316), .ZN(n12378) );
  NAND2_X1 U15525 ( .A1(n12378), .A2(n12950), .ZN(n12379) );
  NOR2_X1 U15526 ( .A1(n14723), .A2(n16266), .ZN(n12380) );
  AOI211_X1 U15527 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n15094), .A(
        n12381), .B(n12380), .ZN(n12385) );
  OR2_X1 U15528 ( .A1(n12383), .A2(n19202), .ZN(n12384) );
  NAND2_X1 U15529 ( .A1(n12387), .A2(n12386), .ZN(P2_U3018) );
  AOI21_X1 U15530 ( .B1(n9744), .B2(n9731), .A(n12623), .ZN(n12414) );
  NAND2_X1 U15531 ( .A1(n12414), .A2(n13357), .ZN(n12771) );
  OR2_X1 U15532 ( .A1(n12979), .A2(n12771), .ZN(n12390) );
  INV_X1 U15533 ( .A(n12388), .ZN(n12859) );
  NAND3_X1 U15534 ( .A1(n12859), .A2(n12968), .A3(n20856), .ZN(n12389) );
  NAND2_X1 U15535 ( .A1(n12390), .A2(n12389), .ZN(n12797) );
  INV_X1 U15536 ( .A(n20209), .ZN(n13185) );
  NAND4_X1 U15537 ( .A1(n13185), .A2(n13000), .A3(n12982), .A4(n11155), .ZN(
        n13178) );
  NOR2_X1 U15538 ( .A1(n12766), .A2(n13178), .ZN(n12391) );
  INV_X1 U15539 ( .A(n20856), .ZN(n20783) );
  OR3_X1 U15540 ( .A1(n12854), .A2(n12626), .A3(n20783), .ZN(n13091) );
  AND2_X1 U15541 ( .A1(n15908), .A2(n13185), .ZN(n12393) );
  NAND2_X1 U15542 ( .A1(n12423), .A2(n12393), .ZN(n12409) );
  NAND2_X1 U15543 ( .A1(n15908), .A2(n12394), .ZN(n12405) );
  NOR4_X1 U15544 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n12398) );
  NOR4_X1 U15545 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(
        P1_ADDRESS_REG_19__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_18__SCAN_IN), .ZN(n12397) );
  NOR4_X1 U15546 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12396) );
  NOR4_X1 U15547 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_8__SCAN_IN), .A3(P1_ADDRESS_REG_10__SCAN_IN), .A4(
        P1_ADDRESS_REG_9__SCAN_IN), .ZN(n12395) );
  AND4_X1 U15548 ( .A1(n12398), .A2(n12397), .A3(n12396), .A4(n12395), .ZN(
        n12403) );
  NOR4_X1 U15549 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12401) );
  NOR4_X1 U15550 ( .A1(P1_ADDRESS_REG_24__SCAN_IN), .A2(
        P1_ADDRESS_REG_23__SCAN_IN), .A3(P1_ADDRESS_REG_22__SCAN_IN), .A4(
        P1_ADDRESS_REG_21__SCAN_IN), .ZN(n12400) );
  NOR4_X1 U15551 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_27__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_25__SCAN_IN), .ZN(n12399) );
  AND4_X1 U15552 ( .A1(n12401), .A2(n12400), .A3(n12399), .A4(n20795), .ZN(
        n12402) );
  NAND2_X1 U15553 ( .A1(n12403), .A2(n12402), .ZN(n12404) );
  NOR2_X1 U15554 ( .A1(n12405), .A2(n14221), .ZN(n14198) );
  AOI22_X1 U15555 ( .A1(n14198), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(n14289), .ZN(n12407) );
  NAND2_X1 U15556 ( .A1(n13069), .A2(n14221), .ZN(n14197) );
  INV_X1 U15557 ( .A(DATAI_31_), .ZN(n12406) );
  NAND2_X1 U15558 ( .A1(n12409), .A2(n12408), .ZN(P1_U2873) );
  NAND2_X1 U15559 ( .A1(n12410), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n16045) );
  INV_X1 U15560 ( .A(n12411), .ZN(n12413) );
  OR2_X1 U15561 ( .A1(n11137), .A2(n11204), .ZN(n12412) );
  AND2_X1 U15562 ( .A1(n12413), .A2(n12412), .ZN(n12757) );
  NAND2_X1 U15563 ( .A1(n12790), .A2(n12415), .ZN(n15802) );
  NAND2_X1 U15564 ( .A1(n20711), .A2(n12416), .ZN(n20855) );
  NAND2_X1 U15565 ( .A1(n20855), .A2(n20773), .ZN(n12417) );
  NAND2_X1 U15566 ( .A1(n20773), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12419) );
  NAND2_X1 U15567 ( .A1(n20649), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12418) );
  AND2_X1 U15568 ( .A1(n12419), .A2(n12418), .ZN(n12932) );
  INV_X1 U15569 ( .A(n12932), .ZN(n12420) );
  NOR2_X1 U15570 ( .A1(n19990), .A2(n20836), .ZN(n14470) );
  AOI21_X1 U15571 ( .B1(n20111), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14470), .ZN(n12421) );
  OAI21_X1 U15572 ( .B1(n20122), .B2(n13364), .A(n12421), .ZN(n12422) );
  AOI21_X1 U15573 ( .B1(n12423), .B2(n20117), .A(n12422), .ZN(n12523) );
  INV_X1 U15574 ( .A(n12485), .ZN(n12452) );
  NOR2_X1 U15575 ( .A1(n12424), .A2(n12452), .ZN(n12425) );
  INV_X4 U15576 ( .A(n14342), .ZN(n15923) );
  NAND2_X1 U15577 ( .A1(n12426), .A2(n12485), .ZN(n12430) );
  NAND2_X1 U15578 ( .A1(n12431), .A2(n12439), .ZN(n12450) );
  XNOR2_X1 U15579 ( .A(n12450), .B(n12449), .ZN(n12428) );
  NAND2_X1 U15580 ( .A1(n9731), .A2(n20189), .ZN(n12438) );
  INV_X1 U15581 ( .A(n12438), .ZN(n12427) );
  AOI21_X1 U15582 ( .B1(n12428), .B2(n13002), .A(n12427), .ZN(n12429) );
  NAND2_X1 U15583 ( .A1(n12430), .A2(n12429), .ZN(n13125) );
  XNOR2_X1 U15584 ( .A(n12431), .B(n12439), .ZN(n12433) );
  INV_X1 U15585 ( .A(n12623), .ZN(n12432) );
  OAI211_X1 U15586 ( .C1(n12433), .C2(n20858), .A(n12432), .B(n20198), .ZN(
        n12434) );
  INV_X1 U15587 ( .A(n12434), .ZN(n12435) );
  OAI21_X1 U15588 ( .B1(n12436), .B2(n12626), .A(n12435), .ZN(n12444) );
  OAI21_X1 U15589 ( .B1(n20858), .B2(n12439), .A(n12438), .ZN(n12440) );
  INV_X1 U15590 ( .A(n12440), .ZN(n12441) );
  XNOR2_X1 U15591 ( .A(n12444), .B(n12933), .ZN(n13056) );
  NAND2_X1 U15592 ( .A1(n13056), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13057) );
  INV_X1 U15593 ( .A(n12933), .ZN(n12443) );
  NAND2_X1 U15594 ( .A1(n12444), .A2(n12443), .ZN(n12445) );
  NAND2_X1 U15595 ( .A1(n12446), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12447) );
  INV_X1 U15596 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12448) );
  NAND2_X1 U15597 ( .A1(n12450), .A2(n12449), .ZN(n12467) );
  XNOR2_X1 U15598 ( .A(n12467), .B(n12465), .ZN(n12451) );
  OAI22_X1 U15599 ( .A1(n20162), .A2(n12452), .B1(n20858), .B2(n12451), .ZN(
        n13196) );
  NAND2_X1 U15600 ( .A1(n12453), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12454) );
  NAND2_X1 U15601 ( .A1(n12455), .A2(n12485), .ZN(n12459) );
  NAND2_X1 U15602 ( .A1(n12467), .A2(n12465), .ZN(n12456) );
  XNOR2_X1 U15603 ( .A(n12456), .B(n12464), .ZN(n12457) );
  NAND2_X1 U15604 ( .A1(n12457), .A2(n13002), .ZN(n12458) );
  NAND2_X1 U15605 ( .A1(n12459), .A2(n12458), .ZN(n12461) );
  INV_X1 U15606 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12460) );
  XNOR2_X1 U15607 ( .A(n12461), .B(n12460), .ZN(n20113) );
  NAND2_X1 U15608 ( .A1(n12461), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12462) );
  NAND2_X1 U15609 ( .A1(n12463), .A2(n12485), .ZN(n12470) );
  AND2_X1 U15610 ( .A1(n12465), .A2(n12464), .ZN(n12466) );
  NAND2_X1 U15611 ( .A1(n12467), .A2(n12466), .ZN(n12477) );
  XNOR2_X1 U15612 ( .A(n12477), .B(n12475), .ZN(n12468) );
  NAND2_X1 U15613 ( .A1(n12468), .A2(n13002), .ZN(n12469) );
  NAND2_X1 U15614 ( .A1(n12470), .A2(n12469), .ZN(n12471) );
  INV_X1 U15615 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16042) );
  XNOR2_X1 U15616 ( .A(n12471), .B(n16042), .ZN(n15953) );
  NAND2_X1 U15617 ( .A1(n12471), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12472) );
  NAND3_X1 U15618 ( .A1(n12474), .A2(n12473), .A3(n12485), .ZN(n12480) );
  INV_X1 U15619 ( .A(n12475), .ZN(n12476) );
  OR2_X1 U15620 ( .A1(n12477), .A2(n12476), .ZN(n12487) );
  XNOR2_X1 U15621 ( .A(n12487), .B(n12488), .ZN(n12478) );
  NAND2_X1 U15622 ( .A1(n12478), .A2(n13002), .ZN(n12479) );
  INV_X1 U15623 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12481) );
  NAND2_X1 U15624 ( .A1(n13422), .A2(n12481), .ZN(n12482) );
  INV_X1 U15625 ( .A(n13422), .ZN(n12483) );
  NAND2_X1 U15626 ( .A1(n12483), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12484) );
  NAND2_X1 U15627 ( .A1(n12486), .A2(n12485), .ZN(n12492) );
  INV_X1 U15628 ( .A(n12487), .ZN(n12489) );
  NAND2_X1 U15629 ( .A1(n12489), .A2(n12488), .ZN(n12495) );
  XNOR2_X1 U15630 ( .A(n12495), .B(n12496), .ZN(n12490) );
  NAND2_X1 U15631 ( .A1(n12490), .A2(n13002), .ZN(n12491) );
  NAND2_X1 U15632 ( .A1(n12492), .A2(n12491), .ZN(n12493) );
  OR2_X1 U15633 ( .A1(n12493), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15948) );
  NAND2_X1 U15634 ( .A1(n15946), .A2(n15948), .ZN(n12494) );
  NAND2_X1 U15635 ( .A1(n12493), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15947) );
  INV_X1 U15636 ( .A(n12495), .ZN(n12497) );
  NAND3_X1 U15637 ( .A1(n12497), .A2(n13002), .A3(n12496), .ZN(n12498) );
  NAND2_X1 U15638 ( .A1(n15937), .A2(n12498), .ZN(n13504) );
  OR2_X1 U15639 ( .A1(n13504), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12499) );
  NAND2_X1 U15640 ( .A1(n13504), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12500) );
  INV_X1 U15641 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n13542) );
  NAND2_X1 U15642 ( .A1(n15923), .A2(n13542), .ZN(n12501) );
  NAND2_X1 U15643 ( .A1(n14411), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15921) );
  INV_X1 U15644 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15999) );
  NAND2_X1 U15645 ( .A1(n15923), .A2(n15999), .ZN(n12503) );
  NAND2_X1 U15646 ( .A1(n15921), .A2(n12503), .ZN(n14437) );
  INV_X1 U15647 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15984) );
  NAND2_X1 U15648 ( .A1(n15923), .A2(n15984), .ZN(n14436) );
  NAND2_X1 U15649 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12504) );
  NAND2_X1 U15650 ( .A1(n15923), .A2(n12504), .ZN(n14434) );
  NAND2_X1 U15651 ( .A1(n14436), .A2(n14434), .ZN(n12505) );
  NOR2_X1 U15652 ( .A1(n14437), .A2(n12505), .ZN(n15919) );
  NAND2_X1 U15653 ( .A1(n15923), .A2(n15992), .ZN(n12506) );
  NAND2_X1 U15654 ( .A1(n15919), .A2(n12506), .ZN(n14422) );
  NAND2_X1 U15655 ( .A1(n14411), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12507) );
  NAND2_X1 U15656 ( .A1(n15921), .A2(n12507), .ZN(n14423) );
  INV_X1 U15657 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21157) );
  NAND2_X1 U15658 ( .A1(n14422), .A2(n12513), .ZN(n12509) );
  XNOR2_X1 U15659 ( .A(n15923), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15913) );
  NAND2_X1 U15660 ( .A1(n15923), .A2(n21157), .ZN(n15910) );
  AND2_X1 U15661 ( .A1(n15913), .A2(n15910), .ZN(n12508) );
  NAND2_X1 U15662 ( .A1(n12509), .A2(n12508), .ZN(n14410) );
  OAI21_X1 U15663 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(n14411), .ZN(n12510) );
  INV_X1 U15664 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12511) );
  NAND2_X1 U15665 ( .A1(n15923), .A2(n12511), .ZN(n12512) );
  INV_X1 U15666 ( .A(n12513), .ZN(n12516) );
  INV_X1 U15667 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15940) );
  NAND2_X1 U15668 ( .A1(n12514), .A2(n15940), .ZN(n12515) );
  NAND2_X1 U15669 ( .A1(n14411), .A2(n12515), .ZN(n14432) );
  NAND2_X1 U15670 ( .A1(n14411), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14435) );
  NAND2_X1 U15671 ( .A1(n14432), .A2(n14435), .ZN(n15920) );
  XNOR2_X1 U15672 ( .A(n15923), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14404) );
  NAND2_X1 U15673 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14564) );
  INV_X1 U15674 ( .A(n14564), .ZN(n12517) );
  NAND2_X1 U15675 ( .A1(n12517), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12518) );
  INV_X1 U15676 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14377) );
  NAND2_X1 U15677 ( .A1(n14377), .A2(n14609), .ZN(n12519) );
  NAND2_X1 U15678 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14530) );
  INV_X1 U15679 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14525) );
  NOR2_X1 U15680 ( .A1(n14530), .A2(n14525), .ZN(n14310) );
  INV_X1 U15681 ( .A(n14310), .ZN(n12521) );
  OR3_X1 U15682 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14309) );
  AND2_X1 U15683 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14468) );
  INV_X1 U15684 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14476) );
  NOR2_X1 U15685 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12525) );
  NOR4_X1 U15686 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12524) );
  NAND4_X1 U15687 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12525), .A4(n12524), .ZN(n12538) );
  INV_X1 U15688 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20852) );
  NOR3_X1 U15689 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n20852), .ZN(n12527) );
  NOR4_X1 U15690 ( .A1(P1_BE_N_REG_1__SCAN_IN), .A2(P1_BE_N_REG_2__SCAN_IN), 
        .A3(P1_BE_N_REG_3__SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12526) );
  NAND4_X1 U15691 ( .A1(n20159), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12527), .A4(
        n12526), .ZN(U214) );
  NOR4_X1 U15692 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12531) );
  NOR4_X1 U15693 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12530) );
  NOR4_X1 U15694 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12529) );
  NOR4_X1 U15695 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12528) );
  AND4_X1 U15696 ( .A1(n12531), .A2(n12530), .A3(n12529), .A4(n12528), .ZN(
        n12536) );
  NOR4_X1 U15697 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n12534) );
  NOR4_X1 U15698 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12533) );
  NOR4_X1 U15699 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n12532) );
  AND4_X1 U15700 ( .A1(n12534), .A2(n12533), .A3(n12532), .A4(n19847), .ZN(
        n12535) );
  NAND2_X1 U15701 ( .A1(n12536), .A2(n12535), .ZN(n12537) );
  NOR2_X1 U15702 ( .A1(n13897), .A2(n12538), .ZN(n16419) );
  NAND2_X1 U15703 ( .A1(n16419), .A2(U214), .ZN(U212) );
  NAND2_X1 U15704 ( .A1(n19021), .A2(n19002), .ZN(n19042) );
  AOI211_X1 U15705 ( .C1(n15022), .C2(n12539), .A(n18912), .B(n19042), .ZN(
        n12550) );
  OAI22_X1 U15706 ( .A1(n15019), .A2(n19037), .B1(n10927), .B2(n19012), .ZN(
        n12549) );
  INV_X1 U15707 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n21120) );
  NAND2_X1 U15708 ( .A1(n19021), .A2(n9753), .ZN(n19036) );
  INV_X1 U15709 ( .A(n19036), .ZN(n18931) );
  AOI22_X1 U15710 ( .A1(n12540), .A2(n19032), .B1(n15022), .B2(n18931), .ZN(
        n12541) );
  OAI211_X1 U15711 ( .C1(n21120), .C2(n19010), .A(n12541), .B(n18983), .ZN(
        n12548) );
  AND2_X1 U15712 ( .A1(n13393), .A2(n12542), .ZN(n12543) );
  OR2_X1 U15713 ( .A1(n12543), .A2(n13484), .ZN(n15248) );
  INV_X1 U15714 ( .A(n15232), .ZN(n12546) );
  NAND2_X1 U15715 ( .A1(n13219), .A2(n12544), .ZN(n12545) );
  NAND2_X1 U15716 ( .A1(n12546), .A2(n12545), .ZN(n15245) );
  OAI22_X1 U15717 ( .A1(n15248), .A2(n19034), .B1(n19029), .B2(n15245), .ZN(
        n12547) );
  OR4_X1 U15718 ( .A1(n12550), .A2(n12549), .A3(n12548), .A4(n12547), .ZN(
        P2_U2840) );
  AOI211_X1 U15719 ( .C1(n16138), .C2(n9762), .A(n12551), .B(n19820), .ZN(
        n12562) );
  INV_X1 U15720 ( .A(n12552), .ZN(n12553) );
  OAI22_X1 U15721 ( .A1(n12553), .A2(n19018), .B1(n10984), .B2(n19012), .ZN(
        n12561) );
  OAI22_X1 U15722 ( .A1(n9983), .A2(n19037), .B1(n21110), .B2(n19010), .ZN(
        n12560) );
  OR2_X1 U15723 ( .A1(n14767), .A2(n12554), .ZN(n12555) );
  AND2_X1 U15724 ( .A1(n14754), .A2(n12555), .ZN(n16142) );
  INV_X1 U15725 ( .A(n16142), .ZN(n12558) );
  INV_X1 U15726 ( .A(n14852), .ZN(n12556) );
  OAI21_X1 U15727 ( .B1(n15156), .B2(n12557), .A(n12556), .ZN(n15135) );
  OAI22_X1 U15728 ( .A1(n12558), .A2(n19034), .B1(n19029), .B2(n15135), .ZN(
        n12559) );
  AOI211_X1 U15729 ( .C1(n14962), .C2(n12564), .A(n12563), .B(n19820), .ZN(
        n12577) );
  OAI22_X1 U15730 ( .A1(n12565), .A2(n19018), .B1(n19874), .B2(n19010), .ZN(
        n12576) );
  AOI22_X1 U15731 ( .A1(P2_EBX_REG_21__SCAN_IN), .A2(n19026), .B1(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n18996), .ZN(n12566) );
  INV_X1 U15732 ( .A(n12566), .ZN(n12575) );
  NAND2_X1 U15733 ( .A1(n9807), .A2(n12567), .ZN(n12568) );
  NAND2_X1 U15734 ( .A1(n9778), .A2(n12568), .ZN(n15163) );
  OR2_X1 U15735 ( .A1(n12569), .A2(n12570), .ZN(n12572) );
  AND2_X1 U15736 ( .A1(n12572), .A2(n12571), .ZN(n15166) );
  INV_X1 U15737 ( .A(n15166), .ZN(n12573) );
  OAI22_X1 U15738 ( .A1(n15163), .A2(n19034), .B1(n12573), .B2(n19029), .ZN(
        n12574) );
  OR4_X1 U15739 ( .A1(n12577), .A2(n12576), .A3(n12575), .A4(n12574), .ZN(
        P2_U2834) );
  INV_X1 U15740 ( .A(n16302), .ZN(n19071) );
  AND2_X1 U15741 ( .A1(n19071), .A2(n12578), .ZN(n19040) );
  INV_X1 U15742 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n12580) );
  AND2_X1 U15743 ( .A1(n12682), .A2(n21119), .ZN(n12581) );
  INV_X1 U15744 ( .A(n12581), .ZN(n12579) );
  OAI211_X1 U15745 ( .C1(n19040), .C2(n12580), .A(n12633), .B(n12579), .ZN(
        P2_U2814) );
  INV_X1 U15746 ( .A(n12661), .ZN(n12583) );
  OAI21_X1 U15747 ( .B1(n12581), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n18853), 
        .ZN(n12582) );
  OAI21_X1 U15748 ( .B1(n12583), .B2(n18853), .A(n12582), .ZN(P2_U3612) );
  AOI21_X1 U15749 ( .B1(n12661), .B2(n16328), .A(n12660), .ZN(n12585) );
  AND2_X1 U15750 ( .A1(n12585), .A2(n12584), .ZN(n12586) );
  AND2_X1 U15751 ( .A1(n16292), .A2(n12586), .ZN(n16304) );
  NOR2_X1 U15752 ( .A1(n16304), .A2(n16333), .ZN(n19942) );
  OAI21_X1 U15753 ( .B1(n12668), .B2(n19942), .A(n12587), .ZN(P2_U2819) );
  INV_X1 U15754 ( .A(n18853), .ZN(n12590) );
  NOR2_X1 U15755 ( .A1(n15841), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19130) );
  INV_X1 U15756 ( .A(n19130), .ZN(n19076) );
  NOR2_X1 U15757 ( .A1(n12588), .A2(n19441), .ZN(n16317) );
  OAI22_X1 U15758 ( .A1(n19834), .A2(n19076), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n16317), .ZN(n12589) );
  NOR2_X1 U15759 ( .A1(n12590), .A2(n12589), .ZN(n12596) );
  NAND2_X1 U15760 ( .A1(n19212), .A2(n19898), .ZN(n12591) );
  AOI211_X1 U15761 ( .C1(n19828), .C2(n12591), .A(n16324), .B(n12661), .ZN(
        n12593) );
  AOI21_X1 U15762 ( .B1(n19441), .B2(n21119), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n16330) );
  AOI21_X1 U15763 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n16328), .A(n16330), 
        .ZN(n12592) );
  NOR2_X1 U15764 ( .A1(n12593), .A2(n12592), .ZN(n12595) );
  NAND2_X1 U15765 ( .A1(n12596), .A2(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n12594) );
  OAI21_X1 U15766 ( .B1(n12596), .B2(n12595), .A(n12594), .ZN(P2_U3610) );
  OAI21_X1 U15767 ( .B1(n16264), .B2(n19017), .A(n12597), .ZN(n12598) );
  XOR2_X1 U15768 ( .A(n12598), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n19191) );
  INV_X1 U15769 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19009) );
  NOR2_X1 U15770 ( .A1(n16225), .A2(n19009), .ZN(n12602) );
  OAI21_X1 U15771 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12600), .A(
        n12599), .ZN(n19203) );
  OR2_X1 U15772 ( .A1(n18983), .A2(n19843), .ZN(n19200) );
  OAI21_X1 U15773 ( .B1(n19159), .B2(n19203), .A(n19200), .ZN(n12601) );
  AOI211_X1 U15774 ( .C1(n19009), .C2(n16217), .A(n12602), .B(n12601), .ZN(
        n12604) );
  INV_X1 U15775 ( .A(n12833), .ZN(n13862) );
  INV_X1 U15776 ( .A(n13862), .ZN(n19198) );
  NAND2_X1 U15777 ( .A1(n19156), .A2(n19198), .ZN(n12603) );
  OAI211_X1 U15778 ( .C1(n19191), .C2(n16219), .A(n12604), .B(n12603), .ZN(
        P2_U3013) );
  NAND2_X1 U15779 ( .A1(n20717), .A2(n20772), .ZN(n19952) );
  INV_X1 U15780 ( .A(n19952), .ZN(n12657) );
  AOI21_X1 U15781 ( .B1(n12605), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n12657), 
        .ZN(n12606) );
  NAND2_X1 U15782 ( .A1(n12854), .A2(n12606), .ZN(P1_U2801) );
  OAI21_X1 U15783 ( .B1(n12609), .B2(n12608), .A(n12607), .ZN(n19178) );
  OR2_X1 U15784 ( .A1(n18983), .A2(n19845), .ZN(n19170) );
  OAI21_X1 U15785 ( .B1(n19178), .B2(n19159), .A(n19170), .ZN(n12611) );
  NOR2_X1 U15786 ( .A1(n19152), .A2(n13314), .ZN(n12610) );
  AOI211_X1 U15787 ( .C1(n19154), .C2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n12611), .B(n12610), .ZN(n12617) );
  NAND2_X1 U15788 ( .A1(n12613), .A2(n12612), .ZN(n12614) );
  AND2_X1 U15789 ( .A1(n12615), .A2(n12614), .ZN(n19181) );
  NAND2_X1 U15790 ( .A1(n19181), .A2(n19162), .ZN(n12616) );
  OAI211_X1 U15791 ( .C1(n16211), .C2(n13322), .A(n12617), .B(n12616), .ZN(
        P2_U3012) );
  INV_X1 U15792 ( .A(n12979), .ZN(n12621) );
  INV_X1 U15793 ( .A(n12618), .ZN(n12619) );
  OAI22_X1 U15794 ( .A1(n12621), .A2(n13357), .B1(n12620), .B2(n12619), .ZN(
        n19950) );
  INV_X1 U15795 ( .A(n12966), .ZN(n15835) );
  NOR3_X1 U15796 ( .A1(n13179), .A2(n13357), .A3(n15835), .ZN(n12622) );
  NOR2_X1 U15797 ( .A1(n12622), .A2(n20783), .ZN(n20857) );
  NOR2_X1 U15798 ( .A1(n19950), .A2(n20857), .ZN(n15805) );
  NOR2_X1 U15799 ( .A1(n15805), .A2(n19949), .ZN(n19957) );
  INV_X1 U15800 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n12632) );
  NAND2_X1 U15801 ( .A1(n13006), .A2(n12623), .ZN(n12625) );
  INV_X1 U15802 ( .A(n12792), .ZN(n13356) );
  NAND2_X1 U15803 ( .A1(n13356), .A2(n11104), .ZN(n12624) );
  NOR2_X1 U15804 ( .A1(n9744), .A2(n12626), .ZN(n12978) );
  INV_X1 U15805 ( .A(n12786), .ZN(n12988) );
  AND2_X1 U15806 ( .A1(n15802), .A2(n12771), .ZN(n12984) );
  NAND2_X1 U15807 ( .A1(n12984), .A2(n12627), .ZN(n12629) );
  INV_X1 U15808 ( .A(n12968), .ZN(n12628) );
  AOI22_X1 U15809 ( .A1(n12979), .A2(n12629), .B1(n9805), .B2(n12628), .ZN(
        n12630) );
  OAI21_X1 U15810 ( .B1(n12979), .B2(n12988), .A(n12630), .ZN(n15804) );
  NAND2_X1 U15811 ( .A1(n19957), .A2(n15804), .ZN(n12631) );
  OAI21_X1 U15812 ( .B1(n19957), .B2(n12632), .A(n12631), .ZN(P1_U3484) );
  NOR2_X1 U15813 ( .A1(n12633), .A2(n19834), .ZN(n12634) );
  AOI22_X1 U15814 ( .A1(n12693), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_17__SCAN_IN), .B2(n12748), .ZN(n12638) );
  INV_X1 U15815 ( .A(n12634), .ZN(n12635) );
  NOR2_X2 U15816 ( .A1(n12635), .A2(n16316), .ZN(n12880) );
  INV_X2 U15817 ( .A(n19205), .ZN(n13897) );
  INV_X1 U15818 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n13071) );
  OR2_X1 U15819 ( .A1(n13897), .A2(n13071), .ZN(n12637) );
  NAND2_X1 U15820 ( .A1(n13897), .A2(BUF2_REG_1__SCAN_IN), .ZN(n12636) );
  AND2_X1 U15821 ( .A1(n12637), .A2(n12636), .ZN(n19219) );
  INV_X1 U15822 ( .A(n19219), .ZN(n14882) );
  NAND2_X1 U15823 ( .A1(n12880), .A2(n14882), .ZN(n12728) );
  NAND2_X1 U15824 ( .A1(n12638), .A2(n12728), .ZN(P2_U2953) );
  AOI22_X1 U15825 ( .A1(n12693), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n12748), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n12641) );
  INV_X1 U15826 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n13203) );
  OR2_X1 U15827 ( .A1(n13897), .A2(n13203), .ZN(n12640) );
  NAND2_X1 U15828 ( .A1(n13897), .A2(BUF2_REG_3__SCAN_IN), .ZN(n12639) );
  AND2_X1 U15829 ( .A1(n12640), .A2(n12639), .ZN(n19226) );
  INV_X1 U15830 ( .A(n19226), .ZN(n14876) );
  NAND2_X1 U15831 ( .A1(n12880), .A2(n14876), .ZN(n12724) );
  NAND2_X1 U15832 ( .A1(n12641), .A2(n12724), .ZN(P2_U2955) );
  AOI22_X1 U15833 ( .A1(n12693), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n12748), .ZN(n12645) );
  INV_X1 U15834 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n13092) );
  OR2_X1 U15835 ( .A1(n13897), .A2(n13092), .ZN(n12643) );
  NAND2_X1 U15836 ( .A1(n13897), .A2(BUF2_REG_6__SCAN_IN), .ZN(n12642) );
  AND2_X1 U15837 ( .A1(n12643), .A2(n12642), .ZN(n19242) );
  INV_X1 U15838 ( .A(n19242), .ZN(n12644) );
  NAND2_X1 U15839 ( .A1(n12880), .A2(n12644), .ZN(n12718) );
  NAND2_X1 U15840 ( .A1(n12645), .A2(n12718), .ZN(P2_U2958) );
  AOI22_X1 U15841 ( .A1(n12693), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n12748), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n12649) );
  INV_X1 U15842 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n13105) );
  OR2_X1 U15843 ( .A1(n13897), .A2(n13105), .ZN(n12647) );
  NAND2_X1 U15844 ( .A1(n13897), .A2(BUF2_REG_5__SCAN_IN), .ZN(n12646) );
  AND2_X1 U15845 ( .A1(n12647), .A2(n12646), .ZN(n19237) );
  INV_X1 U15846 ( .A(n19237), .ZN(n12648) );
  NAND2_X1 U15847 ( .A1(n12880), .A2(n12648), .ZN(n12720) );
  NAND2_X1 U15848 ( .A1(n12649), .A2(n12720), .ZN(P2_U2957) );
  AOI22_X1 U15849 ( .A1(n12693), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n12748), .ZN(n12653) );
  INV_X1 U15850 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n13096) );
  OR2_X1 U15851 ( .A1(n13897), .A2(n13096), .ZN(n12651) );
  NAND2_X1 U15852 ( .A1(n13897), .A2(BUF2_REG_4__SCAN_IN), .ZN(n12650) );
  INV_X1 U15853 ( .A(n19232), .ZN(n12652) );
  NAND2_X1 U15854 ( .A1(n12880), .A2(n12652), .ZN(n12697) );
  NAND2_X1 U15855 ( .A1(n12653), .A2(n12697), .ZN(P2_U2956) );
  AOI22_X1 U15856 ( .A1(n12693), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n12748), .ZN(n12656) );
  INV_X1 U15857 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n13131) );
  OR2_X1 U15858 ( .A1(n13897), .A2(n13131), .ZN(n12655) );
  NAND2_X1 U15859 ( .A1(n13897), .A2(BUF2_REG_2__SCAN_IN), .ZN(n12654) );
  AND2_X1 U15860 ( .A1(n12655), .A2(n12654), .ZN(n19222) );
  INV_X1 U15861 ( .A(n19222), .ZN(n13025) );
  NAND2_X1 U15862 ( .A1(n12880), .A2(n13025), .ZN(n12726) );
  NAND2_X1 U15863 ( .A1(n12656), .A2(n12726), .ZN(P2_U2954) );
  NOR2_X1 U15864 ( .A1(n12657), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n12659)
         );
  OAI21_X1 U15865 ( .B1(n13357), .B2(n11926), .A(n20854), .ZN(n12658) );
  OAI21_X1 U15866 ( .B1(n12659), .B2(n20854), .A(n12658), .ZN(P1_U3487) );
  NAND3_X1 U15867 ( .A1(n19072), .A2(n19071), .A3(n12660), .ZN(n12667) );
  NAND2_X1 U15868 ( .A1(n16294), .A2(n16295), .ZN(n12664) );
  NAND3_X1 U15869 ( .A1(n16292), .A2(n12662), .A3(n12661), .ZN(n12663) );
  INV_X1 U15870 ( .A(n12665), .ZN(n12666) );
  INV_X1 U15871 ( .A(n16294), .ZN(n16296) );
  AND4_X1 U15872 ( .A1(n12667), .A2(n12679), .A3(n12666), .A4(n12849), .ZN(
        n16308) );
  NOR2_X1 U15873 ( .A1(n16324), .A2(n15841), .ZN(n15843) );
  INV_X1 U15874 ( .A(n15843), .ZN(n16335) );
  OAI22_X1 U15875 ( .A1(n16308), .A2(n16333), .B1(n12668), .B2(n16335), .ZN(
        n12669) );
  NAND4_X1 U15876 ( .A1(n19071), .A2(n16316), .A3(n16299), .A4(n19817), .ZN(
        n12671) );
  NAND2_X1 U15877 ( .A1(n15376), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12670) );
  OAI21_X1 U15878 ( .B1(n15376), .B2(n12671), .A(n12670), .ZN(P2_U3595) );
  INV_X1 U15879 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n13065) );
  OR2_X1 U15880 ( .A1(n13897), .A2(n13065), .ZN(n12673) );
  NAND2_X1 U15881 ( .A1(n13897), .A2(BUF2_REG_0__SCAN_IN), .ZN(n12672) );
  AND2_X1 U15882 ( .A1(n12673), .A2(n12672), .ZN(n19211) );
  NOR2_X1 U15883 ( .A1(n12675), .A2(n12674), .ZN(n12677) );
  NAND2_X1 U15884 ( .A1(n12677), .A2(n12676), .ZN(n12678) );
  OR2_X1 U15885 ( .A1(n19053), .A2(n12851), .ZN(n13899) );
  INV_X1 U15886 ( .A(n13899), .ZN(n13901) );
  NAND2_X1 U15887 ( .A1(n19243), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12681) );
  AOI22_X1 U15888 ( .A1(n12885), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n12682), .B2(n19933), .ZN(n12683) );
  NAND2_X1 U15889 ( .A1(n13832), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12685) );
  INV_X1 U15890 ( .A(n19028), .ZN(n16263) );
  NOR2_X1 U15891 ( .A1(n19928), .A2(n19028), .ZN(n12872) );
  OAI22_X1 U15892 ( .A1(n12872), .A2(n16133), .B1(n16132), .B2(n19028), .ZN(
        n12689) );
  OAI21_X1 U15893 ( .B1(n19265), .B2(n16263), .A(n12689), .ZN(n12691) );
  NAND2_X1 U15894 ( .A1(n19053), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n12690) );
  OAI211_X1 U15895 ( .C1(n19211), .C2(n19061), .A(n12691), .B(n12690), .ZN(
        P2_U2919) );
  XNOR2_X1 U15896 ( .A(n12692), .B(n9831), .ZN(n18995) );
  INV_X1 U15897 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19125) );
  OAI222_X1 U15898 ( .A1(n19061), .A2(n19242), .B1(n18995), .B2(n19070), .C1(
        n19125), .C2(n19060), .ZN(P2_U2913) );
  AOI22_X1 U15899 ( .A1(n12879), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n12748), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n12696) );
  INV_X1 U15900 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n13101) );
  OR2_X1 U15901 ( .A1(n13897), .A2(n13101), .ZN(n12695) );
  NAND2_X1 U15902 ( .A1(n13897), .A2(BUF2_REG_7__SCAN_IN), .ZN(n12694) );
  AND2_X1 U15903 ( .A1(n12695), .A2(n12694), .ZN(n19248) );
  INV_X1 U15904 ( .A(n19248), .ZN(n14862) );
  NAND2_X1 U15905 ( .A1(n12880), .A2(n14862), .ZN(n12716) );
  NAND2_X1 U15906 ( .A1(n12696), .A2(n12716), .ZN(P2_U2974) );
  AOI22_X1 U15907 ( .A1(n12879), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n12748), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n12698) );
  NAND2_X1 U15908 ( .A1(n12698), .A2(n12697), .ZN(P2_U2971) );
  AOI22_X1 U15909 ( .A1(n12879), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n12748), .ZN(n12701) );
  INV_X1 U15910 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14199) );
  OR2_X1 U15911 ( .A1(n13897), .A2(n14199), .ZN(n12700) );
  NAND2_X1 U15912 ( .A1(n13897), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12699) );
  NAND2_X1 U15913 ( .A1(n12700), .A2(n12699), .ZN(n13903) );
  NAND2_X1 U15914 ( .A1(n12880), .A2(n13903), .ZN(n12744) );
  NAND2_X1 U15915 ( .A1(n12701), .A2(n12744), .ZN(P2_U2966) );
  AOI22_X1 U15916 ( .A1(n12879), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n12748), 
        .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n12704) );
  INV_X1 U15917 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n13479) );
  OR2_X1 U15918 ( .A1(n13897), .A2(n13479), .ZN(n12703) );
  NAND2_X1 U15919 ( .A1(n13897), .A2(BUF2_REG_8__SCAN_IN), .ZN(n12702) );
  NAND2_X1 U15920 ( .A1(n12703), .A2(n12702), .ZN(n14858) );
  NAND2_X1 U15921 ( .A1(n12880), .A2(n14858), .ZN(n12714) );
  NAND2_X1 U15922 ( .A1(n12704), .A2(n12714), .ZN(P2_U2975) );
  AOI22_X1 U15923 ( .A1(n12879), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n12748), .ZN(n12707) );
  INV_X1 U15924 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n14220) );
  OR2_X1 U15925 ( .A1(n13897), .A2(n14220), .ZN(n12706) );
  NAND2_X1 U15926 ( .A1(n13897), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12705) );
  NAND2_X1 U15927 ( .A1(n12706), .A2(n12705), .ZN(n14832) );
  NAND2_X1 U15928 ( .A1(n12880), .A2(n14832), .ZN(n12742) );
  NAND2_X1 U15929 ( .A1(n12707), .A2(n12742), .ZN(P2_U2963) );
  AOI22_X1 U15930 ( .A1(n12879), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_26__SCAN_IN), .B2(n12748), .ZN(n12710) );
  INV_X1 U15931 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n13532) );
  OR2_X1 U15932 ( .A1(n13897), .A2(n13532), .ZN(n12709) );
  NAND2_X1 U15933 ( .A1(n13897), .A2(BUF2_REG_10__SCAN_IN), .ZN(n12708) );
  NAND2_X1 U15934 ( .A1(n12709), .A2(n12708), .ZN(n14842) );
  NAND2_X1 U15935 ( .A1(n12880), .A2(n14842), .ZN(n12722) );
  NAND2_X1 U15936 ( .A1(n12710), .A2(n12722), .ZN(P2_U2962) );
  AOI22_X1 U15937 ( .A1(n12879), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n12748), .ZN(n12713) );
  INV_X1 U15938 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n13513) );
  OR2_X1 U15939 ( .A1(n13897), .A2(n13513), .ZN(n12712) );
  NAND2_X1 U15940 ( .A1(n13897), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12711) );
  NAND2_X1 U15941 ( .A1(n12712), .A2(n12711), .ZN(n14847) );
  NAND2_X1 U15942 ( .A1(n12880), .A2(n14847), .ZN(n12732) );
  NAND2_X1 U15943 ( .A1(n12713), .A2(n12732), .ZN(P2_U2961) );
  AOI22_X1 U15944 ( .A1(n12879), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_24__SCAN_IN), .B2(n12748), .ZN(n12715) );
  NAND2_X1 U15945 ( .A1(n12715), .A2(n12714), .ZN(P2_U2960) );
  AOI22_X1 U15946 ( .A1(n12879), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n12748), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n12717) );
  NAND2_X1 U15947 ( .A1(n12717), .A2(n12716), .ZN(P2_U2959) );
  AOI22_X1 U15948 ( .A1(n12879), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n12748), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n12719) );
  NAND2_X1 U15949 ( .A1(n12719), .A2(n12718), .ZN(P2_U2973) );
  AOI22_X1 U15950 ( .A1(n12879), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n12748), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n12721) );
  NAND2_X1 U15951 ( .A1(n12721), .A2(n12720), .ZN(P2_U2972) );
  AOI22_X1 U15952 ( .A1(n12879), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n12748), 
        .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n12723) );
  NAND2_X1 U15953 ( .A1(n12723), .A2(n12722), .ZN(P2_U2977) );
  AOI22_X1 U15954 ( .A1(n12879), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n12748), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n12725) );
  NAND2_X1 U15955 ( .A1(n12725), .A2(n12724), .ZN(P2_U2970) );
  AOI22_X1 U15956 ( .A1(n12879), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n12748), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n12727) );
  NAND2_X1 U15957 ( .A1(n12727), .A2(n12726), .ZN(P2_U2969) );
  AOI22_X1 U15958 ( .A1(n12879), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n12748), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n12729) );
  NAND2_X1 U15959 ( .A1(n12729), .A2(n12728), .ZN(P2_U2968) );
  AOI22_X1 U15960 ( .A1(n12879), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n12748), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n12731) );
  INV_X1 U15961 ( .A(n19211), .ZN(n12730) );
  NAND2_X1 U15962 ( .A1(n12880), .A2(n12730), .ZN(n12737) );
  NAND2_X1 U15963 ( .A1(n12731), .A2(n12737), .ZN(P2_U2967) );
  AOI22_X1 U15964 ( .A1(n12879), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n12748), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n12733) );
  NAND2_X1 U15965 ( .A1(n12733), .A2(n12732), .ZN(P2_U2976) );
  AOI22_X1 U15966 ( .A1(n12879), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n12748), .ZN(n12736) );
  INV_X1 U15967 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n14206) );
  OR2_X1 U15968 ( .A1(n13897), .A2(n14206), .ZN(n12735) );
  NAND2_X1 U15969 ( .A1(n13897), .A2(BUF2_REG_13__SCAN_IN), .ZN(n12734) );
  NAND2_X1 U15970 ( .A1(n12735), .A2(n12734), .ZN(n14817) );
  NAND2_X1 U15971 ( .A1(n12880), .A2(n14817), .ZN(n12749) );
  NAND2_X1 U15972 ( .A1(n12736), .A2(n12749), .ZN(P2_U2965) );
  AOI22_X1 U15973 ( .A1(n12879), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n12748), .ZN(n12738) );
  NAND2_X1 U15974 ( .A1(n12738), .A2(n12737), .ZN(P2_U2952) );
  AOI22_X1 U15975 ( .A1(n12879), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(n12748), .ZN(n12741) );
  INV_X1 U15976 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n14213) );
  OR2_X1 U15977 ( .A1(n13897), .A2(n14213), .ZN(n12740) );
  NAND2_X1 U15978 ( .A1(n13897), .A2(BUF2_REG_12__SCAN_IN), .ZN(n12739) );
  NAND2_X1 U15979 ( .A1(n12740), .A2(n12739), .ZN(n14825) );
  NAND2_X1 U15980 ( .A1(n12880), .A2(n14825), .ZN(n12746) );
  NAND2_X1 U15981 ( .A1(n12741), .A2(n12746), .ZN(P2_U2964) );
  AOI22_X1 U15982 ( .A1(n12879), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n12748), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n12743) );
  NAND2_X1 U15983 ( .A1(n12743), .A2(n12742), .ZN(P2_U2978) );
  AOI22_X1 U15984 ( .A1(n12879), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_14__SCAN_IN), .B2(n12748), .ZN(n12745) );
  NAND2_X1 U15985 ( .A1(n12745), .A2(n12744), .ZN(P2_U2981) );
  AOI22_X1 U15986 ( .A1(n12879), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n12748), 
        .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n12747) );
  NAND2_X1 U15987 ( .A1(n12747), .A2(n12746), .ZN(P2_U2979) );
  AOI22_X1 U15988 ( .A1(n12879), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n12748), .ZN(n12750) );
  NAND2_X1 U15989 ( .A1(n12750), .A2(n12749), .ZN(P2_U2980) );
  OAI21_X1 U15990 ( .B1(n12752), .B2(n12751), .A(n12923), .ZN(n18977) );
  OAI222_X1 U15991 ( .A1(n19061), .A2(n19248), .B1(n18977), .B2(n19070), .C1(
        n19123), .C2(n19060), .ZN(P2_U2912) );
  OAI21_X1 U15992 ( .B1(n12974), .B2(n11155), .A(n20209), .ZN(n12754) );
  OAI21_X1 U15993 ( .B1(n12754), .B2(n13180), .A(n9729), .ZN(n12755) );
  OAI211_X1 U15994 ( .C1(n12757), .C2(n13909), .A(n12756), .B(n12755), .ZN(
        n12758) );
  INV_X1 U15995 ( .A(n12758), .ZN(n12762) );
  INV_X1 U15996 ( .A(n11137), .ZN(n12759) );
  AOI21_X1 U15997 ( .B1(n12759), .B2(n9729), .A(n9731), .ZN(n12760) );
  NAND2_X1 U15998 ( .A1(n12761), .A2(n12760), .ZN(n12789) );
  INV_X1 U15999 ( .A(n12765), .ZN(n12767) );
  NAND3_X1 U16000 ( .A1(n12764), .A2(n12767), .A3(n12766), .ZN(n12768) );
  NOR2_X1 U16001 ( .A1(n12993), .A2(n12768), .ZN(n12769) );
  NAND2_X1 U16002 ( .A1(n12769), .A2(n12388), .ZN(n13565) );
  NAND2_X1 U16003 ( .A1(n12753), .A2(n13565), .ZN(n12784) );
  NAND2_X1 U16004 ( .A1(n9805), .A2(n9729), .ZN(n12987) );
  INV_X1 U16005 ( .A(n13150), .ZN(n12770) );
  NAND2_X1 U16006 ( .A1(n15787), .A2(n12770), .ZN(n12776) );
  INV_X1 U16007 ( .A(n12771), .ZN(n12772) );
  OR2_X1 U16008 ( .A1(n12772), .A2(n12786), .ZN(n13152) );
  NAND2_X1 U16009 ( .A1(n12773), .A2(n11038), .ZN(n13146) );
  AOI22_X1 U16010 ( .A1(n15787), .A2(n13150), .B1(n13152), .B2(n13146), .ZN(
        n12775) );
  MUX2_X1 U16011 ( .A(n12776), .B(n12775), .S(n12774), .Z(n12783) );
  INV_X1 U16012 ( .A(n13565), .ZN(n14650) );
  INV_X1 U16013 ( .A(n12777), .ZN(n12778) );
  OAI21_X1 U16014 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n14646), .A(
        n12778), .ZN(n12779) );
  NOR2_X1 U16015 ( .A1(n11121), .A2(n12779), .ZN(n12785) );
  NAND3_X1 U16016 ( .A1(n14650), .A2(n13180), .A3(n12785), .ZN(n12782) );
  NAND3_X1 U16017 ( .A1(n13152), .A2(n12780), .A3(n12773), .ZN(n12781) );
  NAND4_X1 U16018 ( .A1(n12784), .A2(n12783), .A3(n12782), .A4(n12781), .ZN(
        n13159) );
  AOI22_X1 U16019 ( .A1(n14657), .A2(n13159), .B1(n15823), .B2(n12785), .ZN(
        n12802) );
  NAND2_X1 U16020 ( .A1(n12979), .A2(n12786), .ZN(n13177) );
  INV_X1 U16021 ( .A(n13177), .ZN(n12798) );
  AND2_X1 U16022 ( .A1(n11929), .A2(n12966), .ZN(n12787) );
  NAND2_X1 U16023 ( .A1(n15787), .A2(n15835), .ZN(n12803) );
  OAI21_X1 U16024 ( .B1(n12787), .B2(n12764), .A(n12803), .ZN(n12788) );
  NAND2_X1 U16025 ( .A1(n12788), .A2(n20856), .ZN(n12795) );
  AND2_X1 U16026 ( .A1(n12790), .A2(n12789), .ZN(n12791) );
  NOR2_X1 U16027 ( .A1(n12791), .A2(n9805), .ZN(n12977) );
  NOR2_X1 U16028 ( .A1(n12792), .A2(n20184), .ZN(n12793) );
  NOR2_X1 U16029 ( .A1(n12977), .A2(n12793), .ZN(n12794) );
  OAI21_X1 U16030 ( .B1(n12979), .B2(n12795), .A(n12794), .ZN(n12796) );
  NAND2_X1 U16031 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16047), .ZN(n16052) );
  INV_X1 U16032 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19956) );
  NOR2_X1 U16033 ( .A1(n16052), .A2(n19956), .ZN(n12799) );
  AOI21_X1 U16034 ( .B1(n15790), .B2(n12982), .A(n12799), .ZN(n12860) );
  NAND2_X1 U16035 ( .A1(n20773), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n12800) );
  NAND2_X1 U16036 ( .A1(n14662), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12801) );
  OAI21_X1 U16037 ( .B1(n12802), .B2(n14662), .A(n12801), .ZN(P1_U3469) );
  INV_X1 U16038 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n12807) );
  OR3_X1 U16039 ( .A1(n12764), .A2(n20858), .A3(n12966), .ZN(n15813) );
  AND2_X1 U16040 ( .A1(n12803), .A2(n15813), .ZN(n12804) );
  NAND2_X1 U16041 ( .A1(n16047), .A2(n20773), .ZN(n20050) );
  INV_X2 U16042 ( .A(n20050), .ZN(n20075) );
  AOI22_X1 U16043 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n20074), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20075), .ZN(n12806) );
  OAI21_X1 U16044 ( .B1(n12807), .B2(n20044), .A(n12806), .ZN(P1_U2916) );
  INV_X1 U16045 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n12809) );
  AOI22_X1 U16046 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n12808) );
  OAI21_X1 U16047 ( .B1(n12809), .B2(n20044), .A(n12808), .ZN(P1_U2914) );
  INV_X1 U16048 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n12811) );
  AOI22_X1 U16049 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n12810) );
  OAI21_X1 U16050 ( .B1(n12811), .B2(n20044), .A(n12810), .ZN(P1_U2913) );
  INV_X1 U16051 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n12813) );
  AOI22_X1 U16052 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n12812) );
  OAI21_X1 U16053 ( .B1(n12813), .B2(n20044), .A(n12812), .ZN(P1_U2915) );
  INV_X1 U16054 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n12815) );
  AOI22_X1 U16055 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n12814) );
  OAI21_X1 U16056 ( .B1(n12815), .B2(n20044), .A(n12814), .ZN(P1_U2920) );
  INV_X1 U16057 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n12817) );
  AOI22_X1 U16058 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n12816) );
  OAI21_X1 U16059 ( .B1(n12817), .B2(n20044), .A(n12816), .ZN(P1_U2917) );
  AOI22_X1 U16060 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n12818) );
  OAI21_X1 U16061 ( .B1(n11688), .B2(n20044), .A(n12818), .ZN(P1_U2912) );
  INV_X1 U16062 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n12820) );
  AOI22_X1 U16063 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n12819) );
  OAI21_X1 U16064 ( .B1(n12820), .B2(n20044), .A(n12819), .ZN(P1_U2910) );
  INV_X1 U16065 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n12822) );
  AOI22_X1 U16066 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12821) );
  OAI21_X1 U16067 ( .B1(n12822), .B2(n20044), .A(n12821), .ZN(P1_U2908) );
  INV_X1 U16068 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n12824) );
  AOI22_X1 U16069 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12823) );
  OAI21_X1 U16070 ( .B1(n12824), .B2(n20044), .A(n12823), .ZN(P1_U2907) );
  INV_X1 U16071 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n12826) );
  AOI22_X1 U16072 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n12825) );
  OAI21_X1 U16073 ( .B1(n12826), .B2(n20044), .A(n12825), .ZN(P1_U2919) );
  INV_X1 U16074 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n12828) );
  AOI22_X1 U16075 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12827) );
  OAI21_X1 U16076 ( .B1(n12828), .B2(n20044), .A(n12827), .ZN(P1_U2911) );
  INV_X1 U16077 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n12830) );
  AOI22_X1 U16078 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12829) );
  OAI21_X1 U16079 ( .B1(n12830), .B2(n20044), .A(n12829), .ZN(P1_U2909) );
  NAND2_X1 U16080 ( .A1(n13757), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12834) );
  NAND2_X1 U16081 ( .A1(n12885), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12831) );
  NAND2_X1 U16082 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19924), .ZN(
        n19505) );
  NAND2_X1 U16083 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19933), .ZN(
        n19538) );
  NAND2_X1 U16084 ( .A1(n19505), .A2(n19538), .ZN(n19414) );
  NAND2_X1 U16085 ( .A1(n12882), .A2(n19414), .ZN(n19540) );
  NAND2_X1 U16086 ( .A1(n12831), .A2(n19540), .ZN(n12832) );
  INV_X1 U16087 ( .A(n12834), .ZN(n12835) );
  NOR2_X1 U16088 ( .A1(n12836), .A2(n12835), .ZN(n12837) );
  NAND2_X1 U16089 ( .A1(n12838), .A2(n12888), .ZN(n12843) );
  NAND2_X1 U16090 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19566) );
  NAND2_X1 U16091 ( .A1(n19566), .A2(n19915), .ZN(n12841) );
  NAND2_X1 U16092 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19742) );
  INV_X1 U16093 ( .A(n19742), .ZN(n12839) );
  INV_X1 U16094 ( .A(n12883), .ZN(n12840) );
  AND2_X1 U16095 ( .A1(n12841), .A2(n12840), .ZN(n19354) );
  AOI22_X1 U16096 ( .A1(n12885), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n12882), .B2(n19354), .ZN(n12842) );
  NAND2_X1 U16097 ( .A1(n12843), .A2(n12842), .ZN(n12846) );
  INV_X1 U16098 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12844) );
  NOR2_X1 U16099 ( .A1(n13786), .A2(n12844), .ZN(n12845) );
  OR2_X1 U16100 ( .A1(n12846), .A2(n12845), .ZN(n12847) );
  NAND2_X1 U16101 ( .A1(n12846), .A2(n12845), .ZN(n12898) );
  INV_X1 U16102 ( .A(n12848), .ZN(n12949) );
  INV_X1 U16103 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13317) );
  MUX2_X1 U16104 ( .A(n13317), .B(n13322), .S(n14808), .Z(n12852) );
  OAI21_X1 U16105 ( .B1(n19909), .B2(n14811), .A(n12852), .ZN(P2_U2885) );
  AND2_X1 U16106 ( .A1(n20858), .A2(n20783), .ZN(n12853) );
  OR2_X1 U16107 ( .A1(n20083), .A2(n9729), .ZN(n13090) );
  INV_X1 U16108 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n12857) );
  INV_X1 U16109 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n12876) );
  NOR2_X1 U16110 ( .A1(n14221), .A2(n12876), .ZN(n12855) );
  AOI21_X1 U16111 ( .B1(DATAI_15_), .B2(n14221), .A(n12855), .ZN(n14280) );
  INV_X1 U16112 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n12856) );
  OAI222_X1 U16113 ( .A1(n13090), .A2(n12857), .B1(n13091), .B2(n14280), .C1(
        n12856), .C2(n13100), .ZN(P1_U2967) );
  INV_X1 U16114 ( .A(n14662), .ZN(n12862) );
  INV_X1 U16115 ( .A(n20322), .ZN(n20562) );
  XNOR2_X1 U16116 ( .A(n12858), .B(n11363), .ZN(n20019) );
  NAND2_X1 U16117 ( .A1(n20019), .A2(n12859), .ZN(n13166) );
  INV_X1 U16118 ( .A(n14657), .ZN(n13566) );
  OR3_X1 U16119 ( .A1(n13166), .A2(n12860), .A3(n13566), .ZN(n12861) );
  OAI21_X1 U16120 ( .B1(n11363), .B2(n12862), .A(n12861), .ZN(P1_U3468) );
  NAND2_X1 U16121 ( .A1(n12866), .A2(n12865), .ZN(n12869) );
  INV_X1 U16122 ( .A(n12867), .ZN(n12868) );
  NAND2_X1 U16123 ( .A1(n12869), .A2(n12868), .ZN(n19922) );
  INV_X1 U16124 ( .A(n19922), .ZN(n12870) );
  NAND2_X1 U16125 ( .A1(n19910), .A2(n12870), .ZN(n13014) );
  OAI21_X1 U16126 ( .B1(n19910), .B2(n12870), .A(n13014), .ZN(n12871) );
  NOR2_X1 U16127 ( .A1(n12871), .A2(n12872), .ZN(n13016) );
  AOI21_X1 U16128 ( .B1(n12872), .B2(n12871), .A(n13016), .ZN(n12875) );
  AOI22_X1 U16129 ( .A1(n19055), .A2(n19922), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19053), .ZN(n12874) );
  INV_X1 U16130 ( .A(n19061), .ZN(n13083) );
  NAND2_X1 U16131 ( .A1(n13083), .A2(n14882), .ZN(n12873) );
  OAI211_X1 U16132 ( .C1(n12875), .C2(n16133), .A(n12874), .B(n12873), .ZN(
        P2_U2918) );
  OR2_X1 U16133 ( .A1(n13897), .A2(n12876), .ZN(n12878) );
  NAND2_X1 U16134 ( .A1(n13897), .A2(BUF2_REG_15__SCAN_IN), .ZN(n12877) );
  NAND2_X1 U16135 ( .A1(n12878), .A2(n12877), .ZN(n13271) );
  AOI222_X1 U16136 ( .A1(n13271), .A2(n12880), .B1(n12879), .B2(
        P2_LWORD_REG_15__SCAN_IN), .C1(P2_EAX_REG_15__SCAN_IN), .C2(n12748), 
        .ZN(n12881) );
  INV_X1 U16137 ( .A(n12881), .ZN(P2_U2982) );
  NAND2_X1 U16138 ( .A1(n12883), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19804) );
  INV_X1 U16139 ( .A(n19679), .ZN(n12882) );
  OAI211_X1 U16140 ( .C1(n12883), .C2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n19804), .B(n12882), .ZN(n19599) );
  INV_X1 U16141 ( .A(n19599), .ZN(n12884) );
  INV_X1 U16142 ( .A(n12891), .ZN(n12887) );
  INV_X1 U16143 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12886) );
  NOR2_X1 U16144 ( .A1(n13786), .A2(n12886), .ZN(n12890) );
  NAND2_X1 U16145 ( .A1(n12887), .A2(n12890), .ZN(n12901) );
  NAND2_X1 U16146 ( .A1(n12889), .A2(n12888), .ZN(n12894) );
  INV_X1 U16147 ( .A(n12890), .ZN(n12892) );
  NAND2_X1 U16148 ( .A1(n12894), .A2(n12893), .ZN(n12895) );
  NAND2_X1 U16149 ( .A1(n12897), .A2(n12896), .ZN(n12899) );
  NAND2_X1 U16150 ( .A1(n19243), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12900) );
  INV_X1 U16151 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12903) );
  NOR2_X1 U16152 ( .A1(n13786), .A2(n12903), .ZN(n12914) );
  XOR2_X1 U16153 ( .A(n13029), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n12909)
         );
  NAND2_X1 U16154 ( .A1(n12904), .A2(n12919), .ZN(n12906) );
  INV_X1 U16155 ( .A(n13042), .ZN(n12905) );
  AND2_X1 U16156 ( .A1(n12906), .A2(n12905), .ZN(n19005) );
  INV_X1 U16157 ( .A(n19005), .ZN(n13453) );
  NOR2_X1 U16158 ( .A1(n14791), .A2(n13453), .ZN(n12907) );
  AOI21_X1 U16159 ( .B1(P2_EBX_REG_5__SCAN_IN), .B2(n14791), .A(n12907), .ZN(
        n12908) );
  OAI21_X1 U16160 ( .B1(n12909), .B2(n14811), .A(n12908), .ZN(P2_U2882) );
  NOR2_X1 U16161 ( .A1(n13862), .A2(n14791), .ZN(n12910) );
  AOI21_X1 U16162 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n14791), .A(n12910), .ZN(
        n12911) );
  OAI21_X1 U16163 ( .B1(n19910), .B2(n14811), .A(n12911), .ZN(P2_U2886) );
  NOR2_X1 U16164 ( .A1(n19035), .A2(n14791), .ZN(n12912) );
  AOI21_X1 U16165 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n14791), .A(n12912), .ZN(
        n12913) );
  OAI21_X1 U16166 ( .B1(n19928), .B2(n14811), .A(n12913), .ZN(P2_U2887) );
  OR2_X1 U16167 ( .A1(n12915), .A2(n12914), .ZN(n12916) );
  NAND2_X1 U16168 ( .A1(n13029), .A2(n12916), .ZN(n19063) );
  NAND2_X1 U16169 ( .A1(n14804), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n12922) );
  OR2_X1 U16170 ( .A1(n12918), .A2(n12917), .ZN(n12920) );
  AND2_X1 U16171 ( .A1(n12920), .A2(n12919), .ZN(n19144) );
  NAND2_X1 U16172 ( .A1(n19144), .A2(n14808), .ZN(n12921) );
  OAI211_X1 U16173 ( .C1(n19063), .C2(n14811), .A(n12922), .B(n12921), .ZN(
        P2_U2883) );
  INV_X1 U16174 ( .A(n14858), .ZN(n12927) );
  NAND2_X1 U16175 ( .A1(n12924), .A2(n12923), .ZN(n12926) );
  INV_X1 U16176 ( .A(n12938), .ZN(n12925) );
  NAND2_X1 U16177 ( .A1(n12926), .A2(n12925), .ZN(n16236) );
  INV_X1 U16178 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19121) );
  OAI222_X1 U16179 ( .A1(n19061), .A2(n12927), .B1(n16236), .B2(n19070), .C1(
        n19121), .C2(n19060), .ZN(P2_U2911) );
  INV_X1 U16180 ( .A(n12928), .ZN(n12931) );
  OAI21_X1 U16181 ( .B1(n12931), .B2(n12930), .A(n12929), .ZN(n14149) );
  NAND2_X1 U16182 ( .A1(n12932), .A2(n14416), .ZN(n12936) );
  INV_X1 U16183 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n14155) );
  NOR2_X1 U16184 ( .A1(n19990), .A2(n14155), .ZN(n13009) );
  OAI21_X1 U16185 ( .B1(n12934), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12933), .ZN(n13013) );
  NOR2_X1 U16186 ( .A1(n13013), .A2(n19955), .ZN(n12935) );
  AOI211_X1 U16187 ( .C1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n12936), .A(
        n13009), .B(n12935), .ZN(n12937) );
  OAI21_X1 U16188 ( .B1(n20161), .B2(n14149), .A(n12937), .ZN(P1_U2999) );
  INV_X1 U16189 ( .A(n14847), .ZN(n12942) );
  OR2_X1 U16190 ( .A1(n12939), .A2(n12938), .ZN(n12941) );
  NAND2_X1 U16191 ( .A1(n12941), .A2(n12940), .ZN(n18965) );
  INV_X1 U16192 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19119) );
  OAI222_X1 U16193 ( .A1(n19061), .A2(n12942), .B1(n18965), .B2(n19070), .C1(
        n19119), .C2(n19060), .ZN(P2_U2910) );
  NAND2_X1 U16194 ( .A1(n16255), .A2(n15358), .ZN(n12963) );
  INV_X1 U16195 ( .A(n10510), .ZN(n12948) );
  NAND2_X1 U16196 ( .A1(n13859), .A2(n12948), .ZN(n15364) );
  NAND2_X1 U16197 ( .A1(n12950), .A2(n12949), .ZN(n15361) );
  INV_X1 U16198 ( .A(n13885), .ZN(n15360) );
  NAND2_X1 U16199 ( .A1(n15361), .A2(n15360), .ZN(n12953) );
  INV_X1 U16200 ( .A(n12951), .ZN(n12952) );
  NAND2_X1 U16201 ( .A1(n12952), .A2(n10444), .ZN(n15359) );
  AND3_X1 U16202 ( .A1(n15364), .A2(n12953), .A3(n15359), .ZN(n12958) );
  NAND2_X1 U16203 ( .A1(n12955), .A2(n12954), .ZN(n15367) );
  AOI22_X1 U16204 ( .A1(n15367), .A2(n15359), .B1(n10510), .B2(n13859), .ZN(
        n12957) );
  MUX2_X1 U16205 ( .A(n12958), .B(n12957), .S(n12956), .Z(n12961) );
  INV_X1 U16206 ( .A(n12959), .ZN(n12960) );
  AND2_X1 U16207 ( .A1(n12961), .A2(n12960), .ZN(n12962) );
  NAND2_X1 U16208 ( .A1(n12963), .A2(n12962), .ZN(n16285) );
  AOI22_X1 U16209 ( .A1(n19902), .A2(n16327), .B1(n19817), .B2(n16285), .ZN(
        n12965) );
  NAND2_X1 U16210 ( .A1(n15376), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12964) );
  OAI21_X1 U16211 ( .B1(n12965), .B2(n15376), .A(n12964), .ZN(P2_U3596) );
  AOI21_X1 U16212 ( .B1(n9729), .B2(n12966), .A(n20783), .ZN(n12967) );
  NAND2_X1 U16213 ( .A1(n12968), .A2(n12967), .ZN(n12976) );
  NAND2_X1 U16214 ( .A1(n12969), .A2(n20856), .ZN(n12971) );
  OAI211_X1 U16215 ( .C1(n12764), .C2(n12971), .A(n20166), .B(n12970), .ZN(
        n12972) );
  INV_X1 U16216 ( .A(n12972), .ZN(n12973) );
  OR2_X1 U16217 ( .A1(n12979), .A2(n12973), .ZN(n12975) );
  MUX2_X1 U16218 ( .A(n12976), .B(n12975), .S(n12974), .Z(n12981) );
  AOI21_X1 U16219 ( .B1(n12979), .B2(n12978), .A(n12977), .ZN(n12980) );
  NAND2_X1 U16220 ( .A1(n12981), .A2(n12980), .ZN(n12983) );
  OAI211_X1 U16221 ( .C1(n13000), .C2(n10047), .A(n9844), .B(n12984), .ZN(
        n12985) );
  INV_X1 U16222 ( .A(n12985), .ZN(n12986) );
  INV_X1 U16223 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20143) );
  OAI211_X1 U16224 ( .C1(n12991), .C2(n20166), .A(n12990), .B(n12989), .ZN(
        n12992) );
  NOR2_X1 U16225 ( .A1(n12993), .A2(n12992), .ZN(n12994) );
  NAND2_X1 U16226 ( .A1(n14557), .A2(n20143), .ZN(n12996) );
  NAND2_X1 U16227 ( .A1(n13005), .A2(n19990), .ZN(n12995) );
  AOI21_X1 U16228 ( .B1(n14618), .B2(n20143), .A(n20141), .ZN(n14634) );
  INV_X1 U16229 ( .A(n14634), .ZN(n12999) );
  INV_X1 U16230 ( .A(n14557), .ZN(n12997) );
  NAND3_X1 U16231 ( .A1(n12997), .A2(n20143), .A3(n20147), .ZN(n12998) );
  OAI21_X1 U16232 ( .B1(n14555), .B2(n12999), .A(n12998), .ZN(n13012) );
  INV_X1 U16233 ( .A(n12764), .ZN(n13003) );
  AOI22_X1 U16234 ( .A1(n13003), .A2(n13002), .B1(n13001), .B2(n13000), .ZN(
        n13004) );
  OR2_X1 U16235 ( .A1(n13006), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13008) );
  NAND2_X1 U16236 ( .A1(n13008), .A2(n13007), .ZN(n14151) );
  INV_X1 U16237 ( .A(n14151), .ZN(n13010) );
  AOI21_X1 U16238 ( .B1(n20133), .B2(n13010), .A(n13009), .ZN(n13011) );
  OAI211_X1 U16239 ( .C1(n15986), .C2(n13013), .A(n13012), .B(n13011), .ZN(
        P1_U3031) );
  INV_X1 U16240 ( .A(n13014), .ZN(n13015) );
  NOR2_X1 U16241 ( .A1(n13016), .A2(n13015), .ZN(n13024) );
  NAND2_X1 U16242 ( .A1(n13018), .A2(n13017), .ZN(n13021) );
  INV_X1 U16243 ( .A(n13019), .ZN(n13020) );
  NAND2_X1 U16244 ( .A1(n13021), .A2(n13020), .ZN(n19913) );
  INV_X1 U16245 ( .A(n19913), .ZN(n13022) );
  NAND2_X1 U16246 ( .A1(n19909), .A2(n13022), .ZN(n13075) );
  OAI21_X1 U16247 ( .B1(n19909), .B2(n13022), .A(n13075), .ZN(n13023) );
  NOR2_X1 U16248 ( .A1(n13024), .A2(n13023), .ZN(n13077) );
  AOI21_X1 U16249 ( .B1(n13024), .B2(n13023), .A(n13077), .ZN(n13028) );
  AOI22_X1 U16250 ( .A1(n13083), .A2(n13025), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19053), .ZN(n13027) );
  NAND2_X1 U16251 ( .A1(n19913), .A2(n19055), .ZN(n13026) );
  OAI211_X1 U16252 ( .C1(n13028), .C2(n16133), .A(n13027), .B(n13026), .ZN(
        P2_U2917) );
  INV_X1 U16253 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13030) );
  INV_X1 U16254 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13039) );
  XOR2_X1 U16255 ( .A(n13048), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13036)
         );
  AOI21_X1 U16256 ( .B1(n13032), .B2(n13041), .A(n13046), .ZN(n18976) );
  INV_X1 U16257 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13033) );
  NOR2_X1 U16258 ( .A1(n14808), .A2(n13033), .ZN(n13034) );
  AOI21_X1 U16259 ( .B1(n18976), .B2(n14808), .A(n13034), .ZN(n13035) );
  OAI21_X1 U16260 ( .B1(n13036), .B2(n14811), .A(n13035), .ZN(P2_U2880) );
  INV_X1 U16261 ( .A(n14842), .ZN(n13038) );
  XNOR2_X1 U16262 ( .A(n12940), .B(n13037), .ZN(n18959) );
  INV_X1 U16263 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n21013) );
  OAI222_X1 U16264 ( .A1(n19061), .A2(n13038), .B1(n18959), .B2(n19070), .C1(
        n21013), .C2(n19060), .ZN(P2_U2909) );
  NOR2_X1 U16265 ( .A1(n13029), .A2(n13039), .ZN(n13040) );
  OAI211_X1 U16266 ( .C1(n13040), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n14783), .B(n13048), .ZN(n13045) );
  OAI21_X1 U16267 ( .B1(n13043), .B2(n13042), .A(n13041), .ZN(n16210) );
  INV_X1 U16268 ( .A(n16210), .ZN(n18991) );
  NAND2_X1 U16269 ( .A1(n14808), .A2(n18991), .ZN(n13044) );
  OAI211_X1 U16270 ( .C1(n14808), .C2(n18984), .A(n13045), .B(n13044), .ZN(
        P2_U2881) );
  OAI21_X1 U16271 ( .B1(n13047), .B2(n13046), .A(n13115), .ZN(n16241) );
  NAND2_X1 U16272 ( .A1(n13049), .A2(n13050), .ZN(n13111) );
  OAI211_X1 U16273 ( .C1(n13049), .C2(n13050), .A(n13109), .B(n14783), .ZN(
        n13052) );
  NAND2_X1 U16274 ( .A1(n14804), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13051) );
  OAI211_X1 U16275 ( .C1(n16241), .C2(n14791), .A(n13052), .B(n13051), .ZN(
        P2_U2879) );
  OAI21_X1 U16276 ( .B1(n13054), .B2(n13053), .A(n13122), .ZN(n14146) );
  INV_X1 U16277 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n14140) );
  NOR2_X1 U16278 ( .A1(n19990), .A2(n14140), .ZN(n14636) );
  NOR2_X1 U16279 ( .A1(n20122), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13055) );
  AOI211_X1 U16280 ( .C1(n20111), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14636), .B(n13055), .ZN(n13059) );
  OR2_X1 U16281 ( .A1(n13056), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14632) );
  NAND3_X1 U16282 ( .A1(n14632), .A2(n20118), .A3(n13057), .ZN(n13058) );
  OAI211_X1 U16283 ( .C1(n14146), .C2(n20161), .A(n13059), .B(n13058), .ZN(
        P1_U2998) );
  INV_X1 U16284 ( .A(n14832), .ZN(n13063) );
  OR2_X1 U16285 ( .A1(n13061), .A2(n13060), .ZN(n13062) );
  NAND2_X1 U16286 ( .A1(n13062), .A2(n13087), .ZN(n15313) );
  INV_X1 U16287 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19116) );
  OAI222_X1 U16288 ( .A1(n19061), .A2(n13063), .B1(n15313), .B2(n19070), .C1(
        n19116), .C2(n19060), .ZN(P2_U2908) );
  NAND2_X1 U16289 ( .A1(n11137), .A2(n20209), .ZN(n13064) );
  OR2_X1 U16290 ( .A1(n20160), .A2(n13065), .ZN(n13067) );
  NAND2_X1 U16291 ( .A1(n20160), .A2(DATAI_0_), .ZN(n13066) );
  NAND2_X1 U16292 ( .A1(n13067), .A2(n13066), .ZN(n20172) );
  INV_X1 U16293 ( .A(n20172), .ZN(n13070) );
  AND2_X1 U16294 ( .A1(n13181), .A2(n20209), .ZN(n13068) );
  INV_X1 U16295 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20078) );
  OAI222_X1 U16296 ( .A1(n14149), .A2(n14287), .B1(n13070), .B2(n14285), .C1(
        n15908), .C2(n20078), .ZN(P1_U2904) );
  INV_X2 U16297 ( .A(n15906), .ZN(n14287) );
  OR2_X1 U16298 ( .A1(n14221), .A2(n13071), .ZN(n13073) );
  NAND2_X1 U16299 ( .A1(n20160), .A2(DATAI_1_), .ZN(n13072) );
  NAND2_X1 U16300 ( .A1(n13073), .A2(n13072), .ZN(n20181) );
  INV_X1 U16301 ( .A(n20181), .ZN(n13074) );
  INV_X1 U16302 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20073) );
  OAI222_X1 U16303 ( .A1(n14146), .A2(n14287), .B1(n13074), .B2(n14285), .C1(
        n15908), .C2(n20073), .ZN(P1_U2903) );
  INV_X1 U16304 ( .A(n13075), .ZN(n13076) );
  NOR2_X1 U16305 ( .A1(n13077), .A2(n13076), .ZN(n13082) );
  OR2_X1 U16306 ( .A1(n13079), .A2(n13078), .ZN(n13080) );
  NAND2_X1 U16307 ( .A1(n13080), .A2(n13136), .ZN(n19905) );
  XNOR2_X1 U16308 ( .A(n19266), .B(n19905), .ZN(n13081) );
  NOR2_X1 U16309 ( .A1(n13082), .A2(n13081), .ZN(n13140) );
  AOI21_X1 U16310 ( .B1(n13082), .B2(n13081), .A(n13140), .ZN(n13086) );
  INV_X1 U16311 ( .A(n19905), .ZN(n13135) );
  AOI22_X1 U16312 ( .A1(n19055), .A2(n13135), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19053), .ZN(n13085) );
  NAND2_X1 U16313 ( .A1(n13083), .A2(n14876), .ZN(n13084) );
  OAI211_X1 U16314 ( .C1(n13086), .C2(n16133), .A(n13085), .B(n13084), .ZN(
        P2_U2916) );
  INV_X1 U16315 ( .A(n14825), .ZN(n13089) );
  XNOR2_X1 U16316 ( .A(n13088), .B(n13087), .ZN(n18941) );
  INV_X1 U16317 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19114) );
  OAI222_X1 U16318 ( .A1(n19061), .A2(n13089), .B1(n18941), .B2(n19070), .C1(
        n19114), .C2(n19060), .ZN(P2_U2907) );
  AOI22_X1 U16319 ( .A1(n20104), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20101), .ZN(n13095) );
  OR2_X1 U16320 ( .A1(n14221), .A2(n13092), .ZN(n13094) );
  NAND2_X1 U16321 ( .A1(n20160), .A2(DATAI_6_), .ZN(n13093) );
  NAND2_X1 U16322 ( .A1(n13094), .A2(n13093), .ZN(n20204) );
  NAND2_X1 U16323 ( .A1(n20093), .A2(n20204), .ZN(n13330) );
  NAND2_X1 U16324 ( .A1(n13095), .A2(n13330), .ZN(P1_U2958) );
  AOI22_X1 U16325 ( .A1(n20104), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20101), .ZN(n13099) );
  OR2_X1 U16326 ( .A1(n14221), .A2(n13096), .ZN(n13098) );
  NAND2_X1 U16327 ( .A1(n20160), .A2(DATAI_4_), .ZN(n13097) );
  NAND2_X1 U16328 ( .A1(n13098), .A2(n13097), .ZN(n20195) );
  NAND2_X1 U16329 ( .A1(n20093), .A2(n20195), .ZN(n13333) );
  NAND2_X1 U16330 ( .A1(n13099), .A2(n13333), .ZN(P1_U2956) );
  AOI22_X1 U16331 ( .A1(n20104), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20083), .ZN(n13104) );
  OR2_X1 U16332 ( .A1(n14221), .A2(n13101), .ZN(n13103) );
  NAND2_X1 U16333 ( .A1(n14221), .A2(DATAI_7_), .ZN(n13102) );
  NAND2_X1 U16334 ( .A1(n13103), .A2(n13102), .ZN(n20214) );
  NAND2_X1 U16335 ( .A1(n20093), .A2(n20214), .ZN(n13335) );
  NAND2_X1 U16336 ( .A1(n13104), .A2(n13335), .ZN(P1_U2959) );
  AOI22_X1 U16337 ( .A1(n20104), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20101), .ZN(n13108) );
  OR2_X1 U16338 ( .A1(n14221), .A2(n13105), .ZN(n13107) );
  NAND2_X1 U16339 ( .A1(n20160), .A2(DATAI_5_), .ZN(n13106) );
  NAND2_X1 U16340 ( .A1(n13107), .A2(n13106), .ZN(n20200) );
  NAND2_X1 U16341 ( .A1(n20093), .A2(n20200), .ZN(n13339) );
  NAND2_X1 U16342 ( .A1(n13108), .A2(n13339), .ZN(P1_U2957) );
  INV_X1 U16343 ( .A(n13109), .ZN(n13114) );
  INV_X1 U16344 ( .A(n13113), .ZN(n13110) );
  NOR2_X2 U16345 ( .A1(n13111), .A2(n13110), .ZN(n13223) );
  INV_X1 U16346 ( .A(n13112), .ZN(n13242) );
  OAI211_X1 U16347 ( .C1(n13114), .C2(n13113), .A(n14783), .B(n13242), .ZN(
        n13120) );
  NAND2_X1 U16348 ( .A1(n13116), .A2(n13115), .ZN(n13118) );
  INV_X1 U16349 ( .A(n13240), .ZN(n13117) );
  AND2_X1 U16350 ( .A1(n13118), .A2(n13117), .ZN(n16192) );
  NAND2_X1 U16351 ( .A1(n14808), .A2(n16192), .ZN(n13119) );
  OAI211_X1 U16352 ( .C1(n14808), .C2(n10906), .A(n13120), .B(n13119), .ZN(
        P2_U2878) );
  OAI21_X1 U16353 ( .B1(n11341), .B2(n11340), .A(n13123), .ZN(n13389) );
  OAI21_X1 U16354 ( .B1(n13126), .B2(n13125), .A(n13124), .ZN(n13127) );
  INV_X1 U16355 ( .A(n13127), .ZN(n20153) );
  INV_X2 U16356 ( .A(n19990), .ZN(n20123) );
  AOI22_X1 U16357 ( .A1(n20111), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20123), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13128) );
  OAI21_X1 U16358 ( .B1(n20122), .B2(n13379), .A(n13128), .ZN(n13129) );
  AOI21_X1 U16359 ( .B1(n20153), .B2(n20118), .A(n13129), .ZN(n13130) );
  OAI21_X1 U16360 ( .B1(n20161), .B2(n13389), .A(n13130), .ZN(P1_U2997) );
  OR2_X1 U16361 ( .A1(n14221), .A2(n13131), .ZN(n13133) );
  NAND2_X1 U16362 ( .A1(n20160), .A2(DATAI_2_), .ZN(n13132) );
  NAND2_X1 U16363 ( .A1(n13133), .A2(n13132), .ZN(n20186) );
  INV_X1 U16364 ( .A(n20186), .ZN(n13134) );
  INV_X1 U16365 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20071) );
  OAI222_X1 U16366 ( .A1(n13389), .A2(n14287), .B1(n13134), .B2(n14285), .C1(
        n15908), .C2(n20071), .ZN(P1_U2902) );
  NOR2_X1 U16367 ( .A1(n19902), .A2(n13135), .ZN(n13139) );
  NAND2_X1 U16368 ( .A1(n13137), .A2(n13136), .ZN(n13138) );
  NAND2_X1 U16369 ( .A1(n13138), .A2(n10202), .ZN(n13298) );
  OAI21_X1 U16370 ( .B1(n13140), .B2(n13139), .A(n13298), .ZN(n19066) );
  XNOR2_X1 U16371 ( .A(n19066), .B(n19063), .ZN(n13141) );
  NAND2_X1 U16372 ( .A1(n13141), .A2(n19064), .ZN(n13144) );
  INV_X1 U16373 ( .A(n13298), .ZN(n13142) );
  AOI22_X1 U16374 ( .A1(n19055), .A2(n13142), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19053), .ZN(n13143) );
  OAI211_X1 U16375 ( .C1(n19232), .C2(n19061), .A(n13144), .B(n13143), .ZN(
        P2_U2915) );
  NOR2_X1 U16376 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20772), .ZN(n13160) );
  OR2_X1 U16377 ( .A1(n13145), .A2(n14650), .ZN(n13158) );
  INV_X1 U16378 ( .A(n13146), .ZN(n13148) );
  OR2_X1 U16379 ( .A1(n13148), .A2(n13147), .ZN(n14660) );
  INV_X1 U16380 ( .A(n14660), .ZN(n13149) );
  NAND2_X1 U16381 ( .A1(n13180), .A2(n13149), .ZN(n13155) );
  NOR2_X1 U16382 ( .A1(n13151), .A2(n13150), .ZN(n13153) );
  AOI22_X1 U16383 ( .A1(n15787), .A2(n13153), .B1(n13152), .B2(n14660), .ZN(
        n13154) );
  OAI21_X1 U16384 ( .B1(n13565), .B2(n13155), .A(n13154), .ZN(n13156) );
  INV_X1 U16385 ( .A(n13156), .ZN(n13157) );
  NAND2_X1 U16386 ( .A1(n13158), .A2(n13157), .ZN(n14658) );
  MUX2_X1 U16387 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14658), .S(
        n15790), .Z(n15786) );
  AOI22_X1 U16388 ( .A1(n13160), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n20772), .B2(n15786), .ZN(n13162) );
  MUX2_X1 U16389 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n13159), .S(
        n15790), .Z(n15800) );
  AOI22_X1 U16390 ( .A1(n13160), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n15800), .B2(n20772), .ZN(n13161) );
  NOR2_X1 U16391 ( .A1(n13162), .A2(n13161), .ZN(n15811) );
  INV_X1 U16392 ( .A(n11044), .ZN(n13163) );
  NAND2_X1 U16393 ( .A1(n15811), .A2(n13163), .ZN(n14642) );
  AND2_X1 U16394 ( .A1(n15790), .A2(n20772), .ZN(n13165) );
  OAI22_X1 U16395 ( .A1(n13165), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B1(
        n20772), .B2(n19956), .ZN(n13164) );
  AOI21_X1 U16396 ( .B1(n13166), .B2(n13165), .A(n13164), .ZN(n15810) );
  INV_X1 U16397 ( .A(n15810), .ZN(n14641) );
  NAND3_X1 U16398 ( .A1(n14642), .A2(n19956), .A3(n14641), .ZN(n13168) );
  INV_X1 U16399 ( .A(n16052), .ZN(n13167) );
  INV_X1 U16400 ( .A(n20247), .ZN(n13169) );
  AOI21_X1 U16401 ( .B1(n13169), .B2(n20649), .A(n20711), .ZN(n13171) );
  NAND2_X1 U16402 ( .A1(n20247), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20532) );
  INV_X1 U16403 ( .A(n9741), .ZN(n20652) );
  NAND2_X1 U16404 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20573), .ZN(n14643) );
  AOI22_X1 U16405 ( .A1(n13171), .A2(n20532), .B1(n20652), .B2(n14643), .ZN(
        n13173) );
  NAND2_X1 U16406 ( .A1(n20158), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13172) );
  OAI21_X1 U16407 ( .B1(n20158), .B2(n13173), .A(n13172), .ZN(P1_U3477) );
  INV_X1 U16408 ( .A(n20532), .ZN(n20288) );
  AOI21_X1 U16409 ( .B1(n13405), .B2(n20288), .A(n20711), .ZN(n20713) );
  INV_X1 U16410 ( .A(n13405), .ZN(n20163) );
  NAND2_X1 U16411 ( .A1(n20163), .A2(n20532), .ZN(n13174) );
  INV_X1 U16412 ( .A(n13145), .ZN(n20170) );
  AOI22_X1 U16413 ( .A1(n20713), .A2(n13174), .B1(n20170), .B2(n14643), .ZN(
        n13176) );
  NAND2_X1 U16414 ( .A1(n20158), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13175) );
  OAI21_X1 U16415 ( .B1(n20158), .B2(n13176), .A(n13175), .ZN(P1_U3476) );
  INV_X1 U16416 ( .A(n13178), .ZN(n13182) );
  NAND4_X1 U16417 ( .A1(n13182), .A2(n13181), .A3(n13180), .A4(n13179), .ZN(
        n13183) );
  NAND2_X1 U16418 ( .A1(n13187), .A2(n13186), .ZN(n13188) );
  NAND2_X1 U16419 ( .A1(n13235), .A2(n13188), .ZN(n20148) );
  OAI22_X1 U16420 ( .A1(n14196), .A2(n20148), .B1(n13189), .B2(n20040), .ZN(
        n13190) );
  INV_X1 U16421 ( .A(n13190), .ZN(n13191) );
  OAI21_X1 U16422 ( .B1(n13389), .B2(n14194), .A(n13191), .ZN(P1_U2870) );
  XNOR2_X1 U16423 ( .A(n13192), .B(n11929), .ZN(n14633) );
  OAI22_X1 U16424 ( .A1(n14196), .A2(n14633), .B1(n14139), .B2(n20040), .ZN(
        n13193) );
  INV_X1 U16425 ( .A(n13193), .ZN(n13194) );
  OAI21_X1 U16426 ( .B1(n14146), .B2(n14194), .A(n13194), .ZN(P1_U2871) );
  OAI21_X1 U16427 ( .B1(n13197), .B2(n13196), .A(n13195), .ZN(n20134) );
  XOR2_X1 U16428 ( .A(n13198), .B(n13199), .Z(n13359) );
  NOR2_X1 U16429 ( .A1(n19990), .A2(n13362), .ZN(n20131) );
  AOI21_X1 U16430 ( .B1(n20111), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20131), .ZN(n13200) );
  OAI21_X1 U16431 ( .B1(n20122), .B2(n13366), .A(n13200), .ZN(n13201) );
  AOI21_X1 U16432 ( .B1(n13359), .B2(n20117), .A(n13201), .ZN(n13202) );
  OAI21_X1 U16433 ( .B1(n19955), .B2(n20134), .A(n13202), .ZN(P1_U2996) );
  INV_X1 U16434 ( .A(n13359), .ZN(n13237) );
  OR2_X1 U16435 ( .A1(n14221), .A2(n13203), .ZN(n13205) );
  NAND2_X1 U16436 ( .A1(n20160), .A2(DATAI_3_), .ZN(n13204) );
  NAND2_X1 U16437 ( .A1(n13205), .A2(n13204), .ZN(n20191) );
  INV_X1 U16438 ( .A(n20191), .ZN(n13206) );
  INV_X1 U16439 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20069) );
  OAI222_X1 U16440 ( .A1(n13237), .A2(n14287), .B1(n13206), .B2(n14285), .C1(
        n15908), .C2(n20069), .ZN(P1_U2901) );
  INV_X1 U16441 ( .A(n14817), .ZN(n13210) );
  INV_X1 U16442 ( .A(n13207), .ZN(n13208) );
  OAI21_X1 U16443 ( .B1(n9828), .B2(n13209), .A(n13208), .ZN(n18936) );
  INV_X1 U16444 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19112) );
  OAI222_X1 U16445 ( .A1(n19061), .A2(n13210), .B1(n18936), .B2(n19070), .C1(
        n19112), .C2(n19060), .ZN(P2_U2906) );
  OAI222_X1 U16446 ( .A1(n14151), .A2(n14196), .B1(n20040), .B2(n13211), .C1(
        n14149), .C2(n14194), .ZN(P1_U2872) );
  NAND2_X1 U16447 ( .A1(n13214), .A2(n13213), .ZN(n13215) );
  XNOR2_X1 U16448 ( .A(n16032), .B(n16034), .ZN(n20124) );
  INV_X1 U16449 ( .A(n20040), .ZN(n14186) );
  AOI22_X1 U16450 ( .A1(n20036), .A2(n20124), .B1(n14186), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n13216) );
  OAI21_X1 U16451 ( .B1(n13218), .B2(n14194), .A(n13216), .ZN(P1_U2868) );
  INV_X1 U16452 ( .A(n20195), .ZN(n13217) );
  INV_X1 U16453 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20067) );
  OAI222_X1 U16454 ( .A1(n13218), .A2(n14287), .B1(n13217), .B2(n14285), .C1(
        n15908), .C2(n20067), .ZN(P1_U2900) );
  INV_X1 U16455 ( .A(n13903), .ZN(n13221) );
  OAI21_X1 U16456 ( .B1(n13207), .B2(n13220), .A(n13219), .ZN(n15267) );
  INV_X1 U16457 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19110) );
  OAI222_X1 U16458 ( .A1(n19061), .A2(n13221), .B1(n15267), .B2(n19070), .C1(
        n19110), .C2(n19060), .ZN(P2_U2905) );
  INV_X1 U16459 ( .A(n13243), .ZN(n13222) );
  NAND2_X1 U16460 ( .A1(n13223), .A2(n13222), .ZN(n13225) );
  INV_X1 U16461 ( .A(n13248), .ZN(n13226) );
  OAI211_X1 U16462 ( .C1(n9911), .C2(n13227), .A(n13226), .B(n14783), .ZN(
        n13232) );
  AND2_X1 U16463 ( .A1(n13239), .A2(n13228), .ZN(n13230) );
  OR2_X1 U16464 ( .A1(n13230), .A2(n13229), .ZN(n15314) );
  INV_X1 U16465 ( .A(n15314), .ZN(n16171) );
  NAND2_X1 U16466 ( .A1(n14808), .A2(n16171), .ZN(n13231) );
  OAI211_X1 U16467 ( .C1(n14808), .C2(n13233), .A(n13232), .B(n13231), .ZN(
        P2_U2876) );
  NAND2_X1 U16468 ( .A1(n13235), .A2(n13234), .ZN(n13236) );
  NAND2_X1 U16469 ( .A1(n16032), .A2(n13236), .ZN(n13363) );
  INV_X1 U16470 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13238) );
  OAI222_X1 U16471 ( .A1(n13363), .A2(n14196), .B1(n13238), .B2(n20040), .C1(
        n14194), .C2(n13237), .ZN(P1_U2869) );
  OAI21_X1 U16472 ( .B1(n13241), .B2(n13240), .A(n13239), .ZN(n16184) );
  INV_X1 U16473 ( .A(n16184), .ZN(n18955) );
  INV_X1 U16474 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n18948) );
  NOR2_X1 U16475 ( .A1(n14808), .A2(n18948), .ZN(n13245) );
  AOI211_X1 U16476 ( .C1(n13243), .C2(n13242), .A(n14811), .B(n9911), .ZN(
        n13244) );
  AOI211_X1 U16477 ( .C1(n18955), .C2(n14808), .A(n13245), .B(n13244), .ZN(
        n13246) );
  INV_X1 U16478 ( .A(n13246), .ZN(P2_U2877) );
  OAI21_X1 U16479 ( .B1(n13229), .B2(n13247), .A(n13347), .ZN(n18942) );
  OAI211_X1 U16480 ( .C1(n13248), .C2(n13249), .A(n13349), .B(n14783), .ZN(
        n13251) );
  NAND2_X1 U16481 ( .A1(n14804), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13250) );
  OAI211_X1 U16482 ( .C1(n18942), .C2(n14791), .A(n13251), .B(n13250), .ZN(
        P2_U2875) );
  NAND2_X1 U16483 ( .A1(n13253), .A2(n13252), .ZN(n13255) );
  XNOR2_X1 U16484 ( .A(n13255), .B(n13254), .ZN(n16259) );
  XNOR2_X1 U16485 ( .A(n13257), .B(n13256), .ZN(n16257) );
  OAI22_X1 U16486 ( .A1(n16225), .A2(n21074), .B1(n13258), .B2(n16226), .ZN(
        n13259) );
  AOI21_X1 U16487 ( .B1(n16217), .B2(n13845), .A(n13259), .ZN(n13261) );
  NAND2_X1 U16488 ( .A1(n16255), .A2(n19156), .ZN(n13260) );
  OAI211_X1 U16489 ( .C1(n16257), .C2(n19159), .A(n13261), .B(n13260), .ZN(
        n13262) );
  AOI21_X1 U16490 ( .B1(n16259), .B2(n19162), .A(n13262), .ZN(n13263) );
  INV_X1 U16491 ( .A(n13263), .ZN(P2_U3011) );
  NAND2_X1 U16492 ( .A1(n13266), .A2(n13265), .ZN(n13267) );
  AND2_X1 U16493 ( .A1(n13264), .A2(n13267), .ZN(n20038) );
  INV_X1 U16494 ( .A(n20038), .ZN(n13270) );
  INV_X1 U16495 ( .A(n20200), .ZN(n13269) );
  OAI222_X1 U16496 ( .A1(n13270), .A2(n14287), .B1(n13269), .B2(n14285), .C1(
        n13268), .C2(n15908), .ZN(P1_U2899) );
  INV_X1 U16497 ( .A(n13271), .ZN(n13272) );
  INV_X1 U16498 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19108) );
  OAI222_X1 U16499 ( .A1(n19061), .A2(n13272), .B1(n15245), .B2(n19070), .C1(
        n19108), .C2(n19060), .ZN(P2_U2904) );
  NAND2_X1 U16500 ( .A1(n13274), .A2(n13273), .ZN(n13275) );
  XNOR2_X1 U16501 ( .A(n13275), .B(n13445), .ZN(n19147) );
  INV_X1 U16502 ( .A(n13276), .ZN(n13277) );
  XNOR2_X1 U16503 ( .A(n13278), .B(n13277), .ZN(n19143) );
  NAND2_X1 U16504 ( .A1(n15337), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15349) );
  NOR2_X1 U16505 ( .A1(n16251), .A2(n13298), .ZN(n13283) );
  INV_X1 U16506 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19848) );
  INV_X1 U16507 ( .A(n19175), .ZN(n15222) );
  AOI21_X1 U16508 ( .B1(n15222), .B2(n13280), .A(n13279), .ZN(n16261) );
  OAI21_X1 U16509 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n19192), .A(
        n16261), .ZN(n13281) );
  INV_X1 U16510 ( .A(n13281), .ZN(n13448) );
  OAI22_X1 U16511 ( .A1(n16226), .A2(n19848), .B1(n13445), .B2(n13448), .ZN(
        n13282) );
  AOI211_X1 U16512 ( .C1(n19144), .C2(n19199), .A(n13283), .B(n13282), .ZN(
        n13284) );
  OAI21_X1 U16513 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15349), .A(
        n13284), .ZN(n13285) );
  AOI21_X1 U16514 ( .B1(n19143), .B2(n19182), .A(n13285), .ZN(n13286) );
  OAI21_X1 U16515 ( .B1(n19202), .B2(n19147), .A(n13286), .ZN(P2_U3042) );
  OAI22_X1 U16516 ( .A1(n19002), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n13866), .B2(n9753), .ZN(n13863) );
  INV_X1 U16517 ( .A(n12364), .ZN(n13287) );
  NAND2_X1 U16518 ( .A1(n13288), .A2(n13287), .ZN(n13858) );
  MUX2_X1 U16519 ( .A(n13858), .B(n13859), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n13289) );
  AOI21_X1 U16520 ( .B1(n19155), .B2(n15358), .A(n13289), .ZN(n16275) );
  INV_X1 U16521 ( .A(n16327), .ZN(n15375) );
  OAI22_X1 U16522 ( .A1(n16275), .A2(n19900), .B1(n12836), .B2(n15375), .ZN(
        n13290) );
  AOI21_X1 U16523 ( .B1(n13863), .B2(P2_STATE2_REG_1__SCAN_IN), .A(n13290), 
        .ZN(n13292) );
  NAND2_X1 U16524 ( .A1(n15376), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13291) );
  OAI21_X1 U16525 ( .B1(n13292), .B2(n15376), .A(n13291), .ZN(P2_U3601) );
  INV_X1 U16526 ( .A(n19040), .ZN(n13855) );
  INV_X1 U16527 ( .A(n19151), .ZN(n13296) );
  NOR2_X1 U16528 ( .A1(n9753), .A2(n13293), .ZN(n13295) );
  AOI21_X1 U16529 ( .B1(n13296), .B2(n13295), .A(n19820), .ZN(n13294) );
  OAI21_X1 U16530 ( .B1(n13296), .B2(n13295), .A(n13294), .ZN(n13304) );
  AOI22_X1 U16531 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18996), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19025), .ZN(n13297) );
  OAI211_X1 U16532 ( .C1(n19029), .C2(n13298), .A(n13297), .B(n18983), .ZN(
        n13299) );
  AOI21_X1 U16533 ( .B1(n19026), .B2(P2_EBX_REG_4__SCAN_IN), .A(n13299), .ZN(
        n13300) );
  OAI21_X1 U16534 ( .B1(n13301), .B2(n19018), .A(n13300), .ZN(n13302) );
  AOI21_X1 U16535 ( .B1(n19144), .B2(n19020), .A(n13302), .ZN(n13303) );
  OAI211_X1 U16536 ( .C1(n13855), .C2(n19063), .A(n13304), .B(n13303), .ZN(
        P2_U2851) );
  NOR2_X1 U16537 ( .A1(n9753), .A2(n13305), .ZN(n13306) );
  XNOR2_X1 U16538 ( .A(n13306), .B(n16209), .ZN(n13307) );
  NAND2_X1 U16539 ( .A1(n13307), .A2(n19021), .ZN(n13312) );
  AOI22_X1 U16540 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18996), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19025), .ZN(n13308) );
  OAI211_X1 U16541 ( .C1(n19029), .C2(n16236), .A(n13308), .B(n16226), .ZN(
        n13310) );
  NOR2_X1 U16542 ( .A1(n16241), .A2(n19034), .ZN(n13309) );
  AOI211_X1 U16543 ( .C1(n19026), .C2(P2_EBX_REG_8__SCAN_IN), .A(n13310), .B(
        n13309), .ZN(n13311) );
  OAI211_X1 U16544 ( .C1(n19018), .C2(n13313), .A(n13312), .B(n13311), .ZN(
        P2_U2847) );
  NOR2_X1 U16545 ( .A1(n9753), .A2(n13864), .ZN(n13315) );
  XNOR2_X1 U16546 ( .A(n13315), .B(n13314), .ZN(n13316) );
  NAND2_X1 U16547 ( .A1(n13316), .A2(n19021), .ZN(n13325) );
  OAI22_X1 U16548 ( .A1(n13317), .A2(n19012), .B1(n19845), .B2(n19010), .ZN(
        n13320) );
  NOR2_X1 U16549 ( .A1(n19018), .A2(n13318), .ZN(n13319) );
  AOI211_X1 U16550 ( .C1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .C2(n18996), .A(
        n13320), .B(n13319), .ZN(n13321) );
  OAI21_X1 U16551 ( .B1(n13322), .B2(n19034), .A(n13321), .ZN(n13323) );
  AOI21_X1 U16552 ( .B1(n19913), .B2(n19015), .A(n13323), .ZN(n13324) );
  OAI211_X1 U16553 ( .C1(n19909), .C2(n13855), .A(n13325), .B(n13324), .ZN(
        P2_U2853) );
  AOI22_X1 U16554 ( .A1(n20104), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20083), .ZN(n13326) );
  NAND2_X1 U16555 ( .A1(n20093), .A2(n20181), .ZN(n13328) );
  NAND2_X1 U16556 ( .A1(n13326), .A2(n13328), .ZN(P1_U2938) );
  AOI22_X1 U16557 ( .A1(n20104), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20083), .ZN(n13327) );
  NAND2_X1 U16558 ( .A1(n20093), .A2(n20191), .ZN(n13337) );
  NAND2_X1 U16559 ( .A1(n13327), .A2(n13337), .ZN(P1_U2940) );
  AOI22_X1 U16560 ( .A1(n20104), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20101), .ZN(n13329) );
  NAND2_X1 U16561 ( .A1(n13329), .A2(n13328), .ZN(P1_U2953) );
  AOI22_X1 U16562 ( .A1(n20104), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20101), .ZN(n13331) );
  NAND2_X1 U16563 ( .A1(n13331), .A2(n13330), .ZN(P1_U2943) );
  AOI22_X1 U16564 ( .A1(n20104), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20101), .ZN(n13332) );
  NAND2_X1 U16565 ( .A1(n20093), .A2(n20186), .ZN(n13342) );
  NAND2_X1 U16566 ( .A1(n13332), .A2(n13342), .ZN(P1_U2939) );
  AOI22_X1 U16567 ( .A1(n20104), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20101), .ZN(n13334) );
  NAND2_X1 U16568 ( .A1(n13334), .A2(n13333), .ZN(P1_U2941) );
  AOI22_X1 U16569 ( .A1(n20104), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20101), .ZN(n13336) );
  NAND2_X1 U16570 ( .A1(n13336), .A2(n13335), .ZN(P1_U2944) );
  AOI22_X1 U16571 ( .A1(n20104), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20101), .ZN(n13338) );
  NAND2_X1 U16572 ( .A1(n13338), .A2(n13337), .ZN(P1_U2955) );
  AOI22_X1 U16573 ( .A1(n20104), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20101), .ZN(n13340) );
  NAND2_X1 U16574 ( .A1(n13340), .A2(n13339), .ZN(P1_U2942) );
  AOI22_X1 U16575 ( .A1(n20104), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20101), .ZN(n13341) );
  NAND2_X1 U16576 ( .A1(n20093), .A2(n20172), .ZN(n13344) );
  NAND2_X1 U16577 ( .A1(n13341), .A2(n13344), .ZN(P1_U2937) );
  AOI22_X1 U16578 ( .A1(n20104), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20101), .ZN(n13343) );
  NAND2_X1 U16579 ( .A1(n13343), .A2(n13342), .ZN(P1_U2954) );
  AOI22_X1 U16580 ( .A1(n20104), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20101), .ZN(n13345) );
  NAND2_X1 U16581 ( .A1(n13345), .A2(n13344), .ZN(P1_U2952) );
  NAND2_X1 U16582 ( .A1(n13347), .A2(n13346), .ZN(n13348) );
  INV_X1 U16583 ( .A(n18933), .ZN(n13355) );
  INV_X1 U16584 ( .A(n13349), .ZN(n13352) );
  OAI211_X1 U16585 ( .C1(n13352), .C2(n13351), .A(n14783), .B(n13413), .ZN(
        n13354) );
  NAND2_X1 U16586 ( .A1(n14804), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13353) );
  OAI211_X1 U16587 ( .C1(n13355), .C2(n14791), .A(n13354), .B(n13353), .ZN(
        P2_U2874) );
  INV_X1 U16588 ( .A(n12753), .ZN(n13375) );
  NAND2_X1 U16589 ( .A1(n20854), .A2(n13356), .ZN(n20018) );
  NAND2_X1 U16590 ( .A1(n20854), .A2(n13357), .ZN(n13358) );
  NAND2_X1 U16591 ( .A1(n19996), .A2(n13358), .ZN(n20022) );
  NAND2_X1 U16592 ( .A1(n13359), .A2(n20022), .ZN(n13374) );
  AND2_X1 U16593 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n13360) );
  NAND2_X1 U16594 ( .A1(n19982), .A2(n13360), .ZN(n13361) );
  AND2_X1 U16595 ( .A1(n14112), .A2(n13361), .ZN(n13387) );
  INV_X1 U16596 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13362) );
  NAND4_X1 U16597 ( .A1(n20005), .A2(n13362), .A3(P1_REIP_REG_2__SCAN_IN), 
        .A4(P1_REIP_REG_1__SCAN_IN), .ZN(n13371) );
  INV_X1 U16598 ( .A(n13363), .ZN(n20132) );
  NAND2_X1 U16599 ( .A1(n20025), .A2(n20132), .ZN(n13370) );
  NAND2_X1 U16600 ( .A1(n20021), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n13369) );
  INV_X1 U16601 ( .A(n13366), .ZN(n13367) );
  AOI22_X1 U16602 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n20024), .B1(
        n20027), .B2(n13367), .ZN(n13368) );
  NAND4_X1 U16603 ( .A1(n13371), .A2(n13370), .A3(n13369), .A4(n13368), .ZN(
        n13372) );
  AOI21_X1 U16604 ( .B1(n13387), .B2(P1_REIP_REG_3__SCAN_IN), .A(n13372), .ZN(
        n13373) );
  OAI211_X1 U16605 ( .C1(n13375), .C2(n20018), .A(n13374), .B(n13373), .ZN(
        P1_U2837) );
  INV_X1 U16606 ( .A(n20022), .ZN(n14150) );
  NAND2_X1 U16607 ( .A1(n20005), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n13377) );
  INV_X1 U16608 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n13376) );
  NAND2_X1 U16609 ( .A1(n13377), .A2(n13376), .ZN(n13386) );
  INV_X1 U16610 ( .A(n20148), .ZN(n13378) );
  NAND2_X1 U16611 ( .A1(n20025), .A2(n13378), .ZN(n13384) );
  NAND2_X1 U16612 ( .A1(n20021), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n13383) );
  INV_X1 U16613 ( .A(n13379), .ZN(n13380) );
  AOI22_X1 U16614 ( .A1(n13380), .A2(n20027), .B1(n20024), .B2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13382) );
  OR2_X1 U16615 ( .A1(n20018), .A2(n13145), .ZN(n13381) );
  NAND4_X1 U16616 ( .A1(n13384), .A2(n13383), .A3(n13382), .A4(n13381), .ZN(
        n13385) );
  AOI21_X1 U16617 ( .B1(n13387), .B2(n13386), .A(n13385), .ZN(n13388) );
  OAI21_X1 U16618 ( .B1(n13389), .B2(n14150), .A(n13388), .ZN(P1_U2838) );
  NAND2_X1 U16619 ( .A1(n13391), .A2(n13390), .ZN(n13392) );
  NAND2_X1 U16620 ( .A1(n13393), .A2(n13392), .ZN(n15262) );
  NOR2_X1 U16621 ( .A1(n9753), .A2(n18923), .ZN(n13394) );
  XNOR2_X1 U16622 ( .A(n13394), .B(n15030), .ZN(n13395) );
  NAND2_X1 U16623 ( .A1(n13395), .A2(n19021), .ZN(n13402) );
  AOI22_X1 U16624 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18996), .B1(
        n19032), .B2(n13396), .ZN(n13397) );
  OAI21_X1 U16625 ( .B1(n19864), .B2(n19010), .A(n13397), .ZN(n13398) );
  NOR2_X1 U16626 ( .A1(n19000), .A2(n13398), .ZN(n13399) );
  OAI21_X1 U16627 ( .B1(n19029), .B2(n15267), .A(n13399), .ZN(n13400) );
  AOI21_X1 U16628 ( .B1(P2_EBX_REG_14__SCAN_IN), .B2(n19026), .A(n13400), .ZN(
        n13401) );
  OAI211_X1 U16629 ( .C1(n15262), .C2(n19034), .A(n13402), .B(n13401), .ZN(
        P2_U2841) );
  INV_X1 U16630 ( .A(n20162), .ZN(n13403) );
  OR2_X1 U16631 ( .A1(n20247), .A2(n20649), .ZN(n20471) );
  NOR2_X1 U16632 ( .A1(n20639), .A2(n20471), .ZN(n20605) );
  AOI211_X1 U16633 ( .C1(n13403), .C2(n20649), .A(n20488), .B(n20605), .ZN(
        n13406) );
  NAND2_X1 U16634 ( .A1(n20420), .A2(n20288), .ZN(n20417) );
  AOI21_X1 U16635 ( .B1(n13406), .B2(n20417), .A(n20711), .ZN(n20714) );
  AOI21_X1 U16636 ( .B1(n14643), .B2(n12753), .A(n20714), .ZN(n13408) );
  NAND2_X1 U16637 ( .A1(n20158), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13407) );
  OAI21_X1 U16638 ( .B1(n20158), .B2(n13408), .A(n13407), .ZN(P1_U3475) );
  INV_X1 U16639 ( .A(n13409), .ZN(n13410) );
  AOI21_X1 U16640 ( .B1(n13411), .B2(n13264), .A(n13410), .ZN(n13433) );
  INV_X1 U16641 ( .A(n13433), .ZN(n19997) );
  INV_X1 U16642 ( .A(n20204), .ZN(n13412) );
  OAI222_X1 U16643 ( .A1(n19997), .A2(n14287), .B1(n13412), .B2(n14285), .C1(
        n15908), .C2(n11382), .ZN(P1_U2898) );
  INV_X1 U16644 ( .A(n13413), .ZN(n13415) );
  INV_X1 U16645 ( .A(n13462), .ZN(n13414) );
  OAI211_X1 U16646 ( .C1(n13415), .C2(n9820), .A(n13414), .B(n14783), .ZN(
        n13417) );
  NAND2_X1 U16647 ( .A1(n14804), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13416) );
  OAI211_X1 U16648 ( .C1(n15262), .C2(n14804), .A(n13417), .B(n13416), .ZN(
        P2_U2873) );
  OR2_X1 U16649 ( .A1(n16036), .A2(n13418), .ZN(n13419) );
  NAND2_X1 U16650 ( .A1(n13469), .A2(n13419), .ZN(n19987) );
  INV_X1 U16651 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n13420) );
  OAI222_X1 U16652 ( .A1(n19987), .A2(n14196), .B1(n20040), .B2(n13420), .C1(
        n14194), .C2(n19997), .ZN(P1_U2866) );
  XNOR2_X1 U16653 ( .A(n13422), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13423) );
  XNOR2_X1 U16654 ( .A(n13421), .B(n13423), .ZN(n13435) );
  NOR2_X1 U16655 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n14555), .ZN(
        n14631) );
  INV_X1 U16656 ( .A(n20140), .ZN(n14619) );
  NAND2_X1 U16657 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20126) );
  NOR2_X1 U16658 ( .A1(n20126), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16038) );
  INV_X1 U16659 ( .A(n16038), .ZN(n13425) );
  NOR2_X1 U16660 ( .A1(n16042), .A2(n20126), .ZN(n16019) );
  NOR2_X1 U16661 ( .A1(n16019), .A2(n20147), .ZN(n13424) );
  OAI21_X1 U16662 ( .B1(n20143), .B2(n20973), .A(n20156), .ZN(n13544) );
  NAND2_X1 U16663 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14454) );
  AOI21_X1 U16664 ( .B1(n20142), .B2(n14454), .A(n20141), .ZN(n13545) );
  OAI21_X1 U16665 ( .B1(n20147), .B2(n13544), .A(n13545), .ZN(n20135) );
  AOI211_X1 U16666 ( .C1(n20142), .C2(n20126), .A(n13424), .B(n20135), .ZN(
        n16043) );
  OAI21_X1 U16667 ( .B1(n14619), .B2(n13425), .A(n16043), .ZN(n16016) );
  OAI21_X1 U16668 ( .B1(n14454), .B2(n14619), .A(n20147), .ZN(n14624) );
  NAND2_X1 U16669 ( .A1(n13544), .A2(n14624), .ZN(n20139) );
  NAND3_X1 U16670 ( .A1(n16019), .A2(n20127), .A3(n12481), .ZN(n13427) );
  NOR2_X1 U16671 ( .A1(n19990), .A2(n20928), .ZN(n13430) );
  INV_X1 U16672 ( .A(n13430), .ZN(n13426) );
  OAI211_X1 U16673 ( .C1(n20149), .C2(n19987), .A(n13427), .B(n13426), .ZN(
        n13428) );
  AOI21_X1 U16674 ( .B1(n16016), .B2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13428), .ZN(n13429) );
  OAI21_X1 U16675 ( .B1(n13435), .B2(n15986), .A(n13429), .ZN(P1_U3025) );
  AOI21_X1 U16676 ( .B1(n20111), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n13430), .ZN(n13431) );
  OAI21_X1 U16677 ( .B1(n20122), .B2(n19995), .A(n13431), .ZN(n13432) );
  AOI21_X1 U16678 ( .B1(n13433), .B2(n20117), .A(n13432), .ZN(n13434) );
  OAI21_X1 U16679 ( .B1(n13435), .B2(n19955), .A(n13434), .ZN(P1_U2993) );
  XNOR2_X1 U16680 ( .A(n13436), .B(n13437), .ZN(n16220) );
  AND2_X1 U16681 ( .A1(n13439), .A2(n13438), .ZN(n13440) );
  OAI22_X1 U16682 ( .A1(n13443), .A2(n13442), .B1(n13441), .B2(n13440), .ZN(
        n16218) );
  INV_X1 U16683 ( .A(n16218), .ZN(n13456) );
  AOI211_X1 U16684 ( .C1(n13449), .C2(n13445), .A(n13444), .B(n15349), .ZN(
        n13455) );
  XNOR2_X1 U16685 ( .A(n13447), .B(n13446), .ZN(n19069) );
  OR2_X1 U16686 ( .A1(n16251), .A2(n19069), .ZN(n13452) );
  OAI22_X1 U16687 ( .A1(n16226), .A2(n12101), .B1(n13449), .B2(n13448), .ZN(
        n13450) );
  INV_X1 U16688 ( .A(n13450), .ZN(n13451) );
  OAI211_X1 U16689 ( .C1(n16266), .C2(n13453), .A(n13452), .B(n13451), .ZN(
        n13454) );
  AOI211_X1 U16690 ( .C1(n13456), .C2(n16231), .A(n13455), .B(n13454), .ZN(
        n13457) );
  OAI21_X1 U16691 ( .B1(n19190), .B2(n16220), .A(n13457), .ZN(P2_U3041) );
  AND2_X1 U16692 ( .A1(n13409), .A2(n13458), .ZN(n13460) );
  OR2_X1 U16693 ( .A1(n13460), .A2(n13459), .ZN(n13467) );
  INV_X1 U16694 ( .A(n20214), .ZN(n13461) );
  OAI222_X1 U16695 ( .A1(n13467), .A2(n14287), .B1(n13461), .B2(n14285), .C1(
        n15908), .C2(n11310), .ZN(P1_U2897) );
  OAI211_X1 U16696 ( .C1(n13462), .C2(n13463), .A(n9914), .B(n14783), .ZN(
        n13466) );
  INV_X1 U16697 ( .A(n15248), .ZN(n13464) );
  NAND2_X1 U16698 ( .A1(n13464), .A2(n14808), .ZN(n13465) );
  OAI211_X1 U16699 ( .C1(n14808), .C2(n10927), .A(n13466), .B(n13465), .ZN(
        P2_U2872) );
  INV_X1 U16700 ( .A(n13467), .ZN(n19981) );
  INV_X1 U16701 ( .A(n14194), .ZN(n20037) );
  NAND2_X1 U16702 ( .A1(n13469), .A2(n13468), .ZN(n13470) );
  AND2_X1 U16703 ( .A1(n13499), .A2(n13470), .ZN(n16026) );
  INV_X1 U16704 ( .A(n16026), .ZN(n19977) );
  OAI22_X1 U16705 ( .A1(n14196), .A2(n19977), .B1(n13471), .B2(n20040), .ZN(
        n13472) );
  AOI21_X1 U16706 ( .B1(n19981), .B2(n20037), .A(n13472), .ZN(n13473) );
  INV_X1 U16707 ( .A(n13473), .ZN(P1_U2865) );
  INV_X1 U16708 ( .A(n13474), .ZN(n13478) );
  INV_X1 U16709 ( .A(n13459), .ZN(n13477) );
  INV_X1 U16710 ( .A(n13475), .ZN(n13476) );
  AOI21_X1 U16711 ( .B1(n13478), .B2(n13477), .A(n13476), .ZN(n13508) );
  INV_X1 U16712 ( .A(n13508), .ZN(n14138) );
  OR2_X1 U16713 ( .A1(n14221), .A2(n13479), .ZN(n13481) );
  NAND2_X1 U16714 ( .A1(n14221), .A2(DATAI_8_), .ZN(n13480) );
  NAND2_X1 U16715 ( .A1(n13481), .A2(n13480), .ZN(n20079) );
  AOI22_X1 U16716 ( .A1(n15905), .A2(n20079), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14289), .ZN(n13482) );
  OAI21_X1 U16717 ( .B1(n14138), .B2(n14287), .A(n13482), .ZN(P1_U2896) );
  OR2_X1 U16718 ( .A1(n13484), .A2(n13483), .ZN(n13485) );
  NAND2_X1 U16719 ( .A1(n14806), .A2(n13485), .ZN(n15236) );
  AOI22_X1 U16720 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10574), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13489) );
  AOI22_X1 U16721 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12959), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13488) );
  AOI22_X1 U16722 ( .A1(n10580), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13487) );
  AOI22_X1 U16723 ( .A1(n10582), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13486) );
  NAND4_X1 U16724 ( .A1(n13489), .A2(n13488), .A3(n13487), .A4(n13486), .ZN(
        n13495) );
  AOI22_X1 U16725 ( .A1(n13647), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13652), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13493) );
  AOI22_X1 U16726 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10575), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13492) );
  AOI22_X1 U16727 ( .A1(n10540), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10546), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13491) );
  AOI22_X1 U16728 ( .A1(n9728), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13622), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13490) );
  NAND4_X1 U16729 ( .A1(n13493), .A2(n13492), .A3(n13491), .A4(n13490), .ZN(
        n13494) );
  INV_X1 U16730 ( .A(n13496), .ZN(n14803) );
  AOI21_X1 U16731 ( .B1(n9845), .B2(n9914), .A(n14803), .ZN(n19056) );
  NAND2_X1 U16732 ( .A1(n19056), .A2(n14783), .ZN(n13498) );
  NAND2_X1 U16733 ( .A1(n14804), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n13497) );
  OAI211_X1 U16734 ( .C1(n15236), .C2(n14804), .A(n13498), .B(n13497), .ZN(
        P2_U2871) );
  AOI21_X1 U16735 ( .B1(n13500), .B2(n13499), .A(n13518), .ZN(n13501) );
  INV_X1 U16736 ( .A(n13501), .ZN(n16020) );
  INV_X1 U16737 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13502) );
  OAI222_X1 U16738 ( .A1(n16020), .A2(n14196), .B1(n20040), .B2(n13502), .C1(
        n14194), .C2(n14138), .ZN(P1_U2864) );
  XOR2_X1 U16739 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n13504), .Z(
        n13505) );
  XNOR2_X1 U16740 ( .A(n13503), .B(n13505), .ZN(n16018) );
  AOI22_X1 U16741 ( .A1(n20111), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n20123), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13506) );
  OAI21_X1 U16742 ( .B1(n20122), .B2(n14131), .A(n13506), .ZN(n13507) );
  AOI21_X1 U16743 ( .B1(n13508), .B2(n20117), .A(n13507), .ZN(n13509) );
  OAI21_X1 U16744 ( .B1(n16018), .B2(n19955), .A(n13509), .ZN(P1_U2991) );
  NOR2_X1 U16745 ( .A1(n13476), .A2(n13511), .ZN(n13512) );
  OR2_X1 U16746 ( .A1(n13510), .A2(n13512), .ZN(n13555) );
  OR2_X1 U16747 ( .A1(n14221), .A2(n13513), .ZN(n13515) );
  NAND2_X1 U16748 ( .A1(n14221), .A2(DATAI_9_), .ZN(n13514) );
  NAND2_X1 U16749 ( .A1(n13515), .A2(n13514), .ZN(n20081) );
  AOI22_X1 U16750 ( .A1(n15905), .A2(n20081), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14289), .ZN(n13516) );
  OAI21_X1 U16751 ( .B1(n13555), .B2(n14287), .A(n13516), .ZN(P1_U2895) );
  NOR2_X1 U16752 ( .A1(n13518), .A2(n13517), .ZN(n13519) );
  OR2_X1 U16753 ( .A1(n13537), .A2(n13519), .ZN(n13540) );
  INV_X1 U16754 ( .A(n13540), .ZN(n13548) );
  OAI21_X1 U16755 ( .B1(n14123), .B2(n19994), .A(n19982), .ZN(n14135) );
  AOI22_X1 U16756 ( .A1(n20025), .A2(n13548), .B1(P1_REIP_REG_9__SCAN_IN), 
        .B2(n14135), .ZN(n13520) );
  OAI211_X1 U16757 ( .C1(n20006), .C2(n13521), .A(n13520), .B(n19990), .ZN(
        n13527) );
  INV_X1 U16758 ( .A(n14123), .ZN(n13522) );
  NOR3_X1 U16759 ( .A1(n19994), .A2(P1_REIP_REG_9__SCAN_IN), .A3(n13522), .ZN(
        n13526) );
  INV_X1 U16760 ( .A(n13552), .ZN(n13523) );
  OAI22_X1 U16761 ( .A1(n20009), .A2(n13524), .B1(n13523), .B2(n20016), .ZN(
        n13525) );
  NOR3_X1 U16762 ( .A1(n13527), .A2(n13526), .A3(n13525), .ZN(n13528) );
  OAI21_X1 U16763 ( .B1(n13555), .B2(n19996), .A(n13528), .ZN(P1_U2831) );
  OAI21_X1 U16764 ( .B1(n13510), .B2(n13531), .A(n13530), .ZN(n14450) );
  OR2_X1 U16765 ( .A1(n14221), .A2(n13532), .ZN(n13534) );
  NAND2_X1 U16766 ( .A1(n14221), .A2(DATAI_10_), .ZN(n13533) );
  NAND2_X1 U16767 ( .A1(n13534), .A2(n13533), .ZN(n20084) );
  AOI22_X1 U16768 ( .A1(n15905), .A2(n20084), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14289), .ZN(n13535) );
  OAI21_X1 U16769 ( .B1(n14450), .B2(n14287), .A(n13535), .ZN(P1_U2894) );
  OAI21_X1 U16770 ( .B1(n13537), .B2(n13536), .A(n15891), .ZN(n13538) );
  INV_X1 U16771 ( .A(n13538), .ZN(n16009) );
  AOI22_X1 U16772 ( .A1(n16009), .A2(n20036), .B1(n14186), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n13539) );
  OAI21_X1 U16773 ( .B1(n14450), .B2(n14194), .A(n13539), .ZN(P1_U2862) );
  OAI222_X1 U16774 ( .A1(n13540), .A2(n14196), .B1(n13524), .B2(n20040), .C1(
        n13555), .C2(n14194), .ZN(P1_U2863) );
  MUX2_X1 U16775 ( .A(n13542), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .S(
        n15937), .Z(n13543) );
  XNOR2_X1 U16776 ( .A(n13541), .B(n13543), .ZN(n13558) );
  INV_X1 U16777 ( .A(n13544), .ZN(n20144) );
  NAND4_X1 U16778 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A4(n16019), .ZN(n14453) );
  NOR2_X1 U16779 ( .A1(n20144), .A2(n14453), .ZN(n14455) );
  OAI21_X1 U16780 ( .B1(n15969), .B2(n14455), .A(n13545), .ZN(n16011) );
  NAND2_X1 U16781 ( .A1(n14455), .A2(n14624), .ZN(n16015) );
  INV_X1 U16782 ( .A(n16015), .ZN(n13546) );
  AOI22_X1 U16783 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16011), .B1(
        n13546), .B2(n13542), .ZN(n13550) );
  INV_X1 U16784 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n13547) );
  NOR2_X1 U16785 ( .A1(n19990), .A2(n13547), .ZN(n13551) );
  AOI21_X1 U16786 ( .B1(n13548), .B2(n20133), .A(n13551), .ZN(n13549) );
  OAI211_X1 U16787 ( .C1(n13558), .C2(n15986), .A(n13550), .B(n13549), .ZN(
        P1_U3022) );
  AOI21_X1 U16788 ( .B1(n20111), .B2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n13551), .ZN(n13554) );
  NAND2_X1 U16789 ( .A1(n15932), .A2(n13552), .ZN(n13553) );
  OAI211_X1 U16790 ( .C1(n13555), .C2(n20161), .A(n13554), .B(n13553), .ZN(
        n13556) );
  INV_X1 U16791 ( .A(n13556), .ZN(n13557) );
  OAI21_X1 U16792 ( .B1(n13558), .B2(n19955), .A(n13557), .ZN(P1_U2990) );
  NOR2_X2 U16793 ( .A1(n18803), .A2(n18811), .ZN(n18635) );
  AOI21_X1 U16794 ( .B1(n18635), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15595) );
  INV_X1 U16795 ( .A(n15379), .ZN(n16981) );
  NAND2_X1 U16796 ( .A1(n15595), .A2(n16981), .ZN(n18174) );
  NOR2_X1 U16797 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18174), .ZN(n13560) );
  NAND3_X1 U16798 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18785)
         );
  INV_X1 U16799 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n20974) );
  INV_X1 U16800 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18687) );
  AOI221_X1 U16801 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n20974), .C1(n18687), 
        .C2(P3_STATE2_REG_1__SCAN_IN), .A(n18815), .ZN(n13559) );
  INV_X1 U16802 ( .A(n13559), .ZN(n18181) );
  OAI21_X1 U16803 ( .B1(n13560), .B2(n18785), .A(n18334), .ZN(n18180) );
  INV_X1 U16804 ( .A(n18180), .ZN(n13561) );
  NOR2_X1 U16805 ( .A1(n20974), .A2(n18834), .ZN(n17810) );
  NAND2_X1 U16806 ( .A1(n20974), .A2(n18787), .ZN(n18845) );
  NAND2_X1 U16807 ( .A1(n18687), .A2(n18787), .ZN(n16494) );
  AND2_X1 U16808 ( .A1(n18845), .A2(n16494), .ZN(n18829) );
  NOR2_X1 U16809 ( .A1(n17810), .A2(n18829), .ZN(n15556) );
  AOI21_X1 U16810 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15556), .ZN(n15557) );
  NOR2_X1 U16811 ( .A1(n13561), .A2(n15557), .ZN(n13563) );
  NAND3_X1 U16812 ( .A1(n18687), .A2(n18787), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18528) );
  INV_X1 U16813 ( .A(n18528), .ZN(n18267) );
  NOR2_X1 U16814 ( .A1(n18787), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18226) );
  OR2_X1 U16815 ( .A1(n18226), .A2(n13561), .ZN(n15555) );
  OR2_X1 U16816 ( .A1(n18267), .A2(n15555), .ZN(n13562) );
  MUX2_X1 U16817 ( .A(n13563), .B(n13562), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  NOR2_X1 U16818 ( .A1(n9744), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13564) );
  AOI21_X1 U16819 ( .B1(n20284), .B2(n13565), .A(n13564), .ZN(n15789) );
  OAI22_X1 U16820 ( .A1(n15789), .A2(n13566), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n20772), .ZN(n13567) );
  AOI21_X1 U16821 ( .B1(n15823), .B2(n13568), .A(n13567), .ZN(n13570) );
  AOI21_X1 U16822 ( .B1(n15787), .B2(n14657), .A(n14662), .ZN(n13569) );
  OAI22_X1 U16823 ( .A1(n13570), .A2(n14662), .B1(n13569), .B2(n13568), .ZN(
        P1_U3474) );
  AND2_X1 U16824 ( .A1(n13572), .A2(n13571), .ZN(n13574) );
  AOI22_X1 U16825 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12162), .B1(
        n10574), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13579) );
  AOI22_X1 U16826 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12959), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13578) );
  AOI22_X1 U16827 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10580), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13577) );
  AOI22_X1 U16828 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10582), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13576) );
  NAND4_X1 U16829 ( .A1(n13579), .A2(n13578), .A3(n13577), .A4(n13576), .ZN(
        n13585) );
  AOI22_X1 U16830 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n13652), .B1(
        n13647), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13583) );
  AOI22_X1 U16831 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10575), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13582) );
  AOI22_X1 U16832 ( .A1(n10540), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n10546), .ZN(n13581) );
  AOI22_X1 U16833 ( .A1(n13621), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13622), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13580) );
  NAND4_X1 U16834 ( .A1(n13583), .A2(n13582), .A3(n13581), .A4(n13580), .ZN(
        n13584) );
  AOI22_X1 U16835 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12162), .B1(
        n10574), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13589) );
  AOI22_X1 U16836 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12959), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13588) );
  AOI22_X1 U16837 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10580), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13587) );
  AOI22_X1 U16838 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10582), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13586) );
  NAND4_X1 U16839 ( .A1(n13589), .A2(n13588), .A3(n13587), .A4(n13586), .ZN(
        n13595) );
  AOI22_X1 U16840 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n13652), .B1(
        n13647), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13593) );
  AOI22_X1 U16841 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10575), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13592) );
  AOI22_X1 U16842 ( .A1(n10540), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n10546), .ZN(n13591) );
  AOI22_X1 U16843 ( .A1(n9728), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13622), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13590) );
  NAND4_X1 U16844 ( .A1(n13593), .A2(n13592), .A3(n13591), .A4(n13590), .ZN(
        n13594) );
  NOR2_X1 U16845 ( .A1(n13595), .A2(n13594), .ZN(n14795) );
  AOI22_X1 U16846 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12162), .B1(
        n10574), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13599) );
  AOI22_X1 U16847 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12959), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13598) );
  AOI22_X1 U16848 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10580), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13597) );
  AOI22_X1 U16849 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10582), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13596) );
  NAND4_X1 U16850 ( .A1(n13599), .A2(n13598), .A3(n13597), .A4(n13596), .ZN(
        n13605) );
  AOI22_X1 U16851 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n13652), .B1(
        n13647), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13603) );
  AOI22_X1 U16852 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10575), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13602) );
  AOI22_X1 U16853 ( .A1(n10540), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n10546), .ZN(n13601) );
  AOI22_X1 U16854 ( .A1(n13621), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13622), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13600) );
  NAND4_X1 U16855 ( .A1(n13603), .A2(n13602), .A3(n13601), .A4(n13600), .ZN(
        n13604) );
  NOR2_X1 U16856 ( .A1(n13605), .A2(n13604), .ZN(n14786) );
  AOI22_X1 U16857 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12162), .B1(
        n10574), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13610) );
  AOI22_X1 U16858 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12959), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13609) );
  AOI22_X1 U16859 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10580), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13608) );
  AOI22_X1 U16860 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10582), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13607) );
  NAND4_X1 U16861 ( .A1(n13610), .A2(n13609), .A3(n13608), .A4(n13607), .ZN(
        n13616) );
  AOI22_X1 U16862 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n13652), .B1(
        n13647), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13614) );
  AOI22_X1 U16863 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10575), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13613) );
  AOI22_X1 U16864 ( .A1(n10540), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n10546), .ZN(n13612) );
  AOI22_X1 U16865 ( .A1(n13621), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13622), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13611) );
  NAND4_X1 U16866 ( .A1(n13614), .A2(n13613), .A3(n13612), .A4(n13611), .ZN(
        n13615) );
  OR2_X1 U16867 ( .A1(n13616), .A2(n13615), .ZN(n14781) );
  AOI22_X1 U16868 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10574), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13620) );
  AOI22_X1 U16869 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12959), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13619) );
  AOI22_X1 U16870 ( .A1(n10580), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13618) );
  AOI22_X1 U16871 ( .A1(n10582), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13617) );
  NAND4_X1 U16872 ( .A1(n13620), .A2(n13619), .A3(n13618), .A4(n13617), .ZN(
        n13634) );
  AOI22_X1 U16873 ( .A1(n13647), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13652), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13632) );
  AOI22_X1 U16874 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10575), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13631) );
  INV_X1 U16875 ( .A(n13621), .ZN(n13624) );
  INV_X1 U16876 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13800) );
  INV_X1 U16877 ( .A(n13622), .ZN(n13623) );
  INV_X1 U16878 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13799) );
  OAI22_X1 U16879 ( .A1(n13624), .A2(n13800), .B1(n13623), .B2(n13799), .ZN(
        n13629) );
  INV_X1 U16880 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13790) );
  INV_X1 U16881 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13626) );
  OAI22_X1 U16882 ( .A1(n13627), .A2(n13790), .B1(n13626), .B2(n13625), .ZN(
        n13628) );
  NOR2_X1 U16883 ( .A1(n13629), .A2(n13628), .ZN(n13630) );
  NAND3_X1 U16884 ( .A1(n13632), .A2(n13631), .A3(n13630), .ZN(n13633) );
  NOR2_X1 U16885 ( .A1(n13634), .A2(n13633), .ZN(n14777) );
  NOR2_X2 U16886 ( .A1(n14776), .A2(n14777), .ZN(n14769) );
  AOI22_X1 U16887 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10574), .B1(
        n12162), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13638) );
  AOI22_X1 U16888 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12959), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13637) );
  AOI22_X1 U16889 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10580), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13636) );
  AOI22_X1 U16890 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10582), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13635) );
  NAND4_X1 U16891 ( .A1(n13638), .A2(n13637), .A3(n13636), .A4(n13635), .ZN(
        n13645) );
  AOI22_X1 U16892 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n13652), .B1(
        n13647), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13643) );
  AOI22_X1 U16893 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10575), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13642) );
  AOI22_X1 U16894 ( .A1(n10540), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n10546), .ZN(n13641) );
  AOI22_X1 U16895 ( .A1(n9728), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13622), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13640) );
  NAND4_X1 U16896 ( .A1(n13643), .A2(n13642), .A3(n13641), .A4(n13640), .ZN(
        n13644) );
  NOR2_X1 U16897 ( .A1(n13645), .A2(n13644), .ZN(n14773) );
  INV_X1 U16898 ( .A(n14773), .ZN(n13646) );
  AND2_X2 U16899 ( .A1(n14769), .A2(n13646), .ZN(n13679) );
  AOI22_X1 U16900 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13647), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13651) );
  AOI22_X1 U16901 ( .A1(n10574), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10575), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13650) );
  AOI22_X1 U16902 ( .A1(n13622), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n10546), .ZN(n13649) );
  AOI22_X1 U16903 ( .A1(n9728), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10540), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13648) );
  NAND4_X1 U16904 ( .A1(n13651), .A2(n13650), .A3(n13649), .A4(n13648), .ZN(
        n13658) );
  AOI22_X1 U16905 ( .A1(n13639), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13652), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13656) );
  AOI22_X1 U16906 ( .A1(n10545), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12959), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13655) );
  AOI22_X1 U16907 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10580), .B1(
        n10581), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13654) );
  AOI22_X1 U16908 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10582), .B1(
        n10607), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13653) );
  NAND4_X1 U16909 ( .A1(n13656), .A2(n13655), .A3(n13654), .A4(n13653), .ZN(
        n13657) );
  OR2_X1 U16910 ( .A1(n13658), .A2(n13657), .ZN(n13702) );
  INV_X1 U16911 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n19269) );
  INV_X1 U16912 ( .A(n13884), .ZN(n13819) );
  INV_X1 U16913 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13659) );
  OAI22_X1 U16914 ( .A1(n13660), .A2(n19269), .B1(n13819), .B2(n13659), .ZN(
        n13663) );
  INV_X1 U16915 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n19331) );
  INV_X1 U16916 ( .A(n10518), .ZN(n13874) );
  INV_X1 U16917 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13661) );
  OAI22_X1 U16918 ( .A1(n15360), .A2(n19331), .B1(n13874), .B2(n13661), .ZN(
        n13662) );
  NOR2_X1 U16919 ( .A1(n13663), .A2(n13662), .ZN(n13666) );
  AOI22_X1 U16920 ( .A1(n13880), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13665) );
  AOI22_X1 U16921 ( .A1(n10506), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13878), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13664) );
  XNOR2_X1 U16922 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13875) );
  NAND4_X1 U16923 ( .A1(n13666), .A2(n13665), .A3(n13664), .A4(n13875), .ZN(
        n13677) );
  INV_X1 U16924 ( .A(n10506), .ZN(n13821) );
  INV_X1 U16925 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13668) );
  INV_X1 U16926 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13667) );
  OAI22_X1 U16927 ( .A1(n13821), .A2(n13668), .B1(n15360), .B2(n13667), .ZN(
        n13672) );
  INV_X1 U16928 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13670) );
  INV_X1 U16929 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13669) );
  OAI22_X1 U16930 ( .A1(n13819), .A2(n13670), .B1(n13874), .B2(n13669), .ZN(
        n13671) );
  NOR2_X1 U16931 ( .A1(n13672), .A2(n13671), .ZN(n13675) );
  INV_X1 U16932 ( .A(n13875), .ZN(n13881) );
  AOI22_X1 U16933 ( .A1(n13878), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13674) );
  AOI22_X1 U16934 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13880), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13673) );
  NAND4_X1 U16935 ( .A1(n13675), .A2(n13881), .A3(n13674), .A4(n13673), .ZN(
        n13676) );
  NAND2_X1 U16936 ( .A1(n13677), .A2(n13676), .ZN(n13706) );
  NOR2_X1 U16937 ( .A1(n16316), .A2(n13706), .ZN(n13678) );
  XOR2_X1 U16938 ( .A(n13702), .B(n13678), .Z(n13704) );
  XNOR2_X1 U16939 ( .A(n13679), .B(n13704), .ZN(n14759) );
  INV_X1 U16940 ( .A(n13706), .ZN(n13701) );
  NAND2_X1 U16941 ( .A1(n16316), .A2(n13701), .ZN(n14762) );
  NOR2_X1 U16942 ( .A1(n14759), .A2(n14762), .ZN(n14760) );
  BUF_X1 U16943 ( .A(n13679), .Z(n14772) );
  AND2_X2 U16944 ( .A1(n14772), .A2(n13704), .ZN(n13680) );
  INV_X1 U16945 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13682) );
  INV_X1 U16946 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13681) );
  OAI22_X1 U16947 ( .A1(n13821), .A2(n13682), .B1(n13819), .B2(n13681), .ZN(
        n13686) );
  INV_X1 U16948 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13684) );
  INV_X1 U16949 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13683) );
  OAI22_X1 U16950 ( .A1(n15360), .A2(n13684), .B1(n13874), .B2(n13683), .ZN(
        n13685) );
  NOR2_X1 U16951 ( .A1(n13686), .A2(n13685), .ZN(n13689) );
  AOI22_X1 U16952 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13880), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13688) );
  AOI22_X1 U16953 ( .A1(n13878), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13687) );
  NAND4_X1 U16954 ( .A1(n13689), .A2(n13688), .A3(n13687), .A4(n13875), .ZN(
        n13700) );
  OAI22_X1 U16955 ( .A1(n13821), .A2(n13691), .B1(n13819), .B2(n13690), .ZN(
        n13695) );
  INV_X1 U16956 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13693) );
  INV_X1 U16957 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13692) );
  OAI22_X1 U16958 ( .A1(n15360), .A2(n13693), .B1(n13874), .B2(n13692), .ZN(
        n13694) );
  NOR2_X1 U16959 ( .A1(n13695), .A2(n13694), .ZN(n13698) );
  AOI22_X1 U16960 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13880), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13697) );
  AOI22_X1 U16961 ( .A1(n13878), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13696) );
  NAND4_X1 U16962 ( .A1(n13698), .A2(n13881), .A3(n13697), .A4(n13696), .ZN(
        n13699) );
  NAND2_X1 U16963 ( .A1(n13700), .A2(n13699), .ZN(n13708) );
  NAND2_X1 U16964 ( .A1(n13702), .A2(n13701), .ZN(n13709) );
  XOR2_X1 U16965 ( .A(n13708), .B(n13709), .Z(n13703) );
  NAND2_X1 U16966 ( .A1(n13703), .A2(n13757), .ZN(n14750) );
  INV_X1 U16967 ( .A(n13704), .ZN(n13707) );
  INV_X1 U16968 ( .A(n13708), .ZN(n13705) );
  NAND2_X1 U16969 ( .A1(n16316), .A2(n13705), .ZN(n14752) );
  NOR2_X1 U16970 ( .A1(n13709), .A2(n13708), .ZN(n13730) );
  INV_X1 U16971 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13711) );
  INV_X1 U16972 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13710) );
  OAI22_X1 U16973 ( .A1(n13821), .A2(n13711), .B1(n13819), .B2(n13710), .ZN(
        n13715) );
  INV_X1 U16974 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13713) );
  INV_X1 U16975 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13712) );
  OAI22_X1 U16976 ( .A1(n15360), .A2(n13713), .B1(n13874), .B2(n13712), .ZN(
        n13714) );
  NOR2_X1 U16977 ( .A1(n13715), .A2(n13714), .ZN(n13718) );
  AOI22_X1 U16978 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13880), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13717) );
  AOI22_X1 U16979 ( .A1(n13878), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13716) );
  NAND4_X1 U16980 ( .A1(n13718), .A2(n13717), .A3(n13716), .A4(n13875), .ZN(
        n13729) );
  INV_X1 U16981 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13720) );
  INV_X1 U16982 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13719) );
  OAI22_X1 U16983 ( .A1(n13821), .A2(n13720), .B1(n13819), .B2(n13719), .ZN(
        n13724) );
  INV_X1 U16984 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13722) );
  INV_X1 U16985 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13721) );
  OAI22_X1 U16986 ( .A1(n15360), .A2(n13722), .B1(n13874), .B2(n13721), .ZN(
        n13723) );
  NOR2_X1 U16987 ( .A1(n13724), .A2(n13723), .ZN(n13727) );
  AOI22_X1 U16988 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13880), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13726) );
  AOI22_X1 U16989 ( .A1(n13878), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13725) );
  NAND4_X1 U16990 ( .A1(n13727), .A2(n13881), .A3(n13726), .A4(n13725), .ZN(
        n13728) );
  AND2_X1 U16991 ( .A1(n13729), .A2(n13728), .ZN(n13732) );
  NAND2_X1 U16992 ( .A1(n13730), .A2(n13732), .ZN(n13785) );
  OAI211_X1 U16993 ( .C1(n13730), .C2(n13732), .A(n13757), .B(n13785), .ZN(
        n13734) );
  XNOR2_X1 U16994 ( .A(n13735), .B(n13731), .ZN(n14743) );
  INV_X1 U16995 ( .A(n13732), .ZN(n13733) );
  NOR2_X1 U16996 ( .A1(n9740), .A2(n13733), .ZN(n14746) );
  INV_X1 U16997 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13738) );
  INV_X1 U16998 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13737) );
  OAI22_X1 U16999 ( .A1(n13821), .A2(n13738), .B1(n13819), .B2(n13737), .ZN(
        n13742) );
  INV_X1 U17000 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13740) );
  INV_X1 U17001 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13739) );
  OAI22_X1 U17002 ( .A1(n15360), .A2(n13740), .B1(n13874), .B2(n13739), .ZN(
        n13741) );
  NOR2_X1 U17003 ( .A1(n13742), .A2(n13741), .ZN(n13745) );
  AOI22_X1 U17004 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13880), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13744) );
  AOI22_X1 U17005 ( .A1(n13878), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13743) );
  NAND4_X1 U17006 ( .A1(n13745), .A2(n13744), .A3(n13743), .A4(n13875), .ZN(
        n13756) );
  INV_X1 U17007 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13747) );
  INV_X1 U17008 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13746) );
  OAI22_X1 U17009 ( .A1(n13821), .A2(n13747), .B1(n13819), .B2(n13746), .ZN(
        n13751) );
  INV_X1 U17010 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13749) );
  INV_X1 U17011 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13748) );
  OAI22_X1 U17012 ( .A1(n15360), .A2(n13749), .B1(n13874), .B2(n13748), .ZN(
        n13750) );
  NOR2_X1 U17013 ( .A1(n13751), .A2(n13750), .ZN(n13754) );
  AOI22_X1 U17014 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13880), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13753) );
  AOI22_X1 U17015 ( .A1(n13878), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13752) );
  NAND4_X1 U17016 ( .A1(n13754), .A2(n13881), .A3(n13753), .A4(n13752), .ZN(
        n13755) );
  AND2_X1 U17017 ( .A1(n13756), .A2(n13755), .ZN(n13759) );
  XNOR2_X1 U17018 ( .A(n13785), .B(n13759), .ZN(n13758) );
  NAND2_X1 U17019 ( .A1(n13758), .A2(n13757), .ZN(n13761) );
  INV_X1 U17020 ( .A(n13759), .ZN(n13784) );
  NOR2_X1 U17021 ( .A1(n9740), .A2(n13784), .ZN(n14736) );
  INV_X1 U17022 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13765) );
  INV_X1 U17023 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13764) );
  OAI22_X1 U17024 ( .A1(n13821), .A2(n13765), .B1(n13819), .B2(n13764), .ZN(
        n13769) );
  INV_X1 U17025 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13767) );
  INV_X1 U17026 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13766) );
  OAI22_X1 U17027 ( .A1(n15360), .A2(n13767), .B1(n13874), .B2(n13766), .ZN(
        n13768) );
  NOR2_X1 U17028 ( .A1(n13769), .A2(n13768), .ZN(n13772) );
  AOI22_X1 U17029 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13880), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13771) );
  AOI22_X1 U17030 ( .A1(n13878), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13770) );
  NAND4_X1 U17031 ( .A1(n13772), .A2(n13771), .A3(n13770), .A4(n13875), .ZN(
        n13783) );
  INV_X1 U17032 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13774) );
  INV_X1 U17033 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13773) );
  OAI22_X1 U17034 ( .A1(n13821), .A2(n13774), .B1(n13819), .B2(n13773), .ZN(
        n13778) );
  INV_X1 U17035 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13776) );
  INV_X1 U17036 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13775) );
  OAI22_X1 U17037 ( .A1(n15360), .A2(n13776), .B1(n13874), .B2(n13775), .ZN(
        n13777) );
  NOR2_X1 U17038 ( .A1(n13778), .A2(n13777), .ZN(n13781) );
  AOI22_X1 U17039 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13880), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13780) );
  AOI22_X1 U17040 ( .A1(n13878), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13779) );
  NAND4_X1 U17041 ( .A1(n13781), .A2(n13881), .A3(n13780), .A4(n13779), .ZN(
        n13782) );
  NAND2_X1 U17042 ( .A1(n13783), .A2(n13782), .ZN(n13789) );
  NOR2_X1 U17043 ( .A1(n13787), .A2(n13789), .ZN(n14720) );
  AOI211_X1 U17044 ( .C1(n13789), .C2(n13787), .A(n13786), .B(n14720), .ZN(
        n13788) );
  NOR2_X1 U17045 ( .A1(n9740), .A2(n13789), .ZN(n14727) );
  OAI22_X1 U17046 ( .A1(n13821), .A2(n13790), .B1(n13819), .B2(n13626), .ZN(
        n13794) );
  INV_X1 U17047 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13792) );
  INV_X1 U17048 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13791) );
  OAI22_X1 U17049 ( .A1(n15360), .A2(n13792), .B1(n13874), .B2(n13791), .ZN(
        n13793) );
  NOR2_X1 U17050 ( .A1(n13794), .A2(n13793), .ZN(n13797) );
  AOI22_X1 U17051 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13880), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13796) );
  AOI22_X1 U17052 ( .A1(n13878), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13795) );
  NAND4_X1 U17053 ( .A1(n13797), .A2(n13796), .A3(n13795), .A4(n13875), .ZN(
        n13808) );
  OAI22_X1 U17054 ( .A1(n13821), .A2(n13799), .B1(n13819), .B2(n13798), .ZN(
        n13803) );
  OAI22_X1 U17055 ( .A1(n15360), .A2(n13801), .B1(n13874), .B2(n13800), .ZN(
        n13802) );
  NOR2_X1 U17056 ( .A1(n13803), .A2(n13802), .ZN(n13806) );
  AOI22_X1 U17057 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13880), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13805) );
  AOI22_X1 U17058 ( .A1(n13878), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13804) );
  NAND4_X1 U17059 ( .A1(n13806), .A2(n13881), .A3(n13805), .A4(n13804), .ZN(
        n13807) );
  NAND2_X1 U17060 ( .A1(n13808), .A2(n13807), .ZN(n14721) );
  INV_X1 U17061 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13810) );
  INV_X1 U17062 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13809) );
  OAI22_X1 U17063 ( .A1(n13821), .A2(n13810), .B1(n15360), .B2(n13809), .ZN(
        n13814) );
  INV_X1 U17064 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13812) );
  INV_X1 U17065 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13811) );
  OAI22_X1 U17066 ( .A1(n13819), .A2(n13812), .B1(n13874), .B2(n13811), .ZN(
        n13813) );
  NOR2_X1 U17067 ( .A1(n13814), .A2(n13813), .ZN(n13817) );
  AOI22_X1 U17068 ( .A1(n13878), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13816) );
  AOI22_X1 U17069 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13880), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13815) );
  NAND4_X1 U17070 ( .A1(n13817), .A2(n13816), .A3(n13815), .A4(n13875), .ZN(
        n13830) );
  INV_X1 U17071 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13820) );
  INV_X1 U17072 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13818) );
  OAI22_X1 U17073 ( .A1(n13821), .A2(n13820), .B1(n13819), .B2(n13818), .ZN(
        n13825) );
  INV_X1 U17074 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13823) );
  INV_X1 U17075 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13822) );
  OAI22_X1 U17076 ( .A1(n15360), .A2(n13823), .B1(n13874), .B2(n13822), .ZN(
        n13824) );
  NOR2_X1 U17077 ( .A1(n13825), .A2(n13824), .ZN(n13828) );
  AOI22_X1 U17078 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13880), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13827) );
  AOI22_X1 U17079 ( .A1(n13878), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13826) );
  NAND4_X1 U17080 ( .A1(n13828), .A2(n13881), .A3(n13827), .A4(n13826), .ZN(
        n13829) );
  NAND2_X1 U17081 ( .A1(n13830), .A2(n13829), .ZN(n13836) );
  INV_X1 U17082 ( .A(n14720), .ZN(n13834) );
  INV_X1 U17083 ( .A(n14721), .ZN(n13831) );
  NAND2_X1 U17084 ( .A1(n13832), .A2(n13831), .ZN(n13833) );
  NOR2_X1 U17085 ( .A1(n13835), .A2(n13836), .ZN(n13869) );
  AOI21_X1 U17086 ( .B1(n13836), .B2(n13835), .A(n13869), .ZN(n13837) );
  OR2_X1 U17087 ( .A1(n13838), .A2(n13837), .ZN(n14812) );
  NAND2_X1 U17088 ( .A1(n13838), .A2(n13837), .ZN(n13871) );
  NAND3_X1 U17089 ( .A1(n14812), .A2(n13871), .A3(n14783), .ZN(n13840) );
  NAND2_X1 U17090 ( .A1(n14804), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n13839) );
  OAI211_X1 U17091 ( .C1(n14804), .C2(n16070), .A(n13840), .B(n13839), .ZN(
        P2_U2858) );
  NAND2_X1 U17092 ( .A1(n16255), .A2(n14808), .ZN(n13842) );
  NAND2_X1 U17093 ( .A1(n14804), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n13841) );
  OAI211_X1 U17094 ( .C1(n19266), .C2(n14811), .A(n13842), .B(n13841), .ZN(
        P2_U2884) );
  NAND2_X1 U17095 ( .A1(n19002), .A2(n13843), .ZN(n13844) );
  XNOR2_X1 U17096 ( .A(n13845), .B(n13844), .ZN(n13846) );
  NAND2_X1 U17097 ( .A1(n13846), .A2(n19021), .ZN(n13854) );
  OAI22_X1 U17098 ( .A1(n13847), .A2(n19012), .B1(n13258), .B2(n19010), .ZN(
        n13849) );
  NOR2_X1 U17099 ( .A1(n19029), .A2(n19905), .ZN(n13848) );
  AOI211_X1 U17100 ( .C1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .C2(n18996), .A(
        n13849), .B(n13848), .ZN(n13850) );
  OAI21_X1 U17101 ( .B1(n13851), .B2(n19018), .A(n13850), .ZN(n13852) );
  AOI21_X1 U17102 ( .B1(n16255), .B2(n19020), .A(n13852), .ZN(n13853) );
  OAI211_X1 U17103 ( .C1(n19266), .C2(n13855), .A(n13854), .B(n13853), .ZN(
        P2_U2852) );
  INV_X1 U17104 ( .A(n15358), .ZN(n13861) );
  NOR2_X1 U17105 ( .A1(n13856), .A2(n12951), .ZN(n13857) );
  AOI22_X1 U17106 ( .A1(n10114), .A2(n13859), .B1(n13858), .B2(n13857), .ZN(
        n13860) );
  OAI21_X1 U17107 ( .B1(n13862), .B2(n13861), .A(n13860), .ZN(n16277) );
  NOR2_X1 U17108 ( .A1(n21119), .A2(n13863), .ZN(n15370) );
  AOI211_X1 U17109 ( .C1(n13866), .C2(n13865), .A(n9753), .B(n13864), .ZN(
        n19022) );
  AOI21_X1 U17110 ( .B1(n9753), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n19022), .ZN(n15371) );
  AOI22_X1 U17111 ( .A1(n16277), .A2(n19817), .B1(n15370), .B2(n15371), .ZN(
        n13867) );
  OAI21_X1 U17112 ( .B1(n19910), .B2(n15375), .A(n13867), .ZN(n13868) );
  MUX2_X1 U17113 ( .A(n13868), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n15376), .Z(P2_U3600) );
  INV_X1 U17114 ( .A(n13869), .ZN(n13870) );
  NAND2_X1 U17115 ( .A1(n13871), .A2(n13870), .ZN(n13895) );
  INV_X1 U17116 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n21069) );
  AOI22_X1 U17117 ( .A1(n13878), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13885), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13873) );
  NAND2_X1 U17118 ( .A1(n13884), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n13872) );
  OAI211_X1 U17119 ( .C1(n13874), .C2(n21069), .A(n13873), .B(n13872), .ZN(
        n13892) );
  AOI22_X1 U17120 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13880), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13877) );
  AOI22_X1 U17121 ( .A1(n10506), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13876) );
  NAND3_X1 U17122 ( .A1(n13877), .A2(n13876), .A3(n13875), .ZN(n13891) );
  AOI22_X1 U17123 ( .A1(n13879), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13878), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13883) );
  AOI22_X1 U17124 ( .A1(n9737), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13880), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13882) );
  NAND3_X1 U17125 ( .A1(n13883), .A2(n13882), .A3(n13881), .ZN(n13890) );
  AOI22_X1 U17126 ( .A1(n13885), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13884), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13888) );
  AOI22_X1 U17127 ( .A1(n10518), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13887) );
  NAND2_X1 U17128 ( .A1(n13888), .A2(n13887), .ZN(n13889) );
  OAI22_X1 U17129 ( .A1(n13892), .A2(n13891), .B1(n13890), .B2(n13889), .ZN(
        n13893) );
  INV_X1 U17130 ( .A(n13893), .ZN(n13894) );
  XNOR2_X1 U17131 ( .A(n13895), .B(n13894), .ZN(n13907) );
  INV_X1 U17132 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13896) );
  NAND2_X1 U17133 ( .A1(n19243), .A2(n13897), .ZN(n13898) );
  INV_X1 U17134 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n19240) );
  INV_X1 U17135 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n19241) );
  AND2_X1 U17136 ( .A1(n19243), .A2(n19205), .ZN(n13900) );
  OAI22_X1 U17137 ( .A1(n19051), .A2(n19240), .B1(n19241), .B2(n19059), .ZN(
        n13902) );
  OAI21_X1 U17138 ( .B1(n13907), .B2(n16133), .A(n13904), .ZN(P2_U2889) );
  NOR2_X1 U17139 ( .A1(n14891), .A2(n14791), .ZN(n13905) );
  AOI21_X1 U17140 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n14791), .A(n13905), .ZN(
        n13906) );
  OAI21_X1 U17141 ( .B1(n13907), .B2(n14811), .A(n13906), .ZN(P2_U2857) );
  OAI22_X1 U17142 ( .A1(n13925), .A2(n13909), .B1(n13938), .B2(n13908), .ZN(
        n13911) );
  NAND2_X1 U17143 ( .A1(n14296), .A2(n19980), .ZN(n13922) );
  INV_X1 U17144 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14159) );
  NAND2_X1 U17145 ( .A1(n13914), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n13917) );
  INV_X1 U17146 ( .A(n14294), .ZN(n13915) );
  AOI22_X1 U17147 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n20024), .B1(
        n20027), .B2(n13915), .ZN(n13916) );
  OAI211_X1 U17148 ( .C1(n20009), .C2(n14159), .A(n13917), .B(n13916), .ZN(
        n13918) );
  AOI21_X1 U17149 ( .B1(n13920), .B2(n13919), .A(n13918), .ZN(n13921) );
  OAI211_X1 U17150 ( .C1(n19978), .C2(n14477), .A(n13922), .B(n13921), .ZN(
        P1_U2810) );
  OAI21_X1 U17151 ( .B1(n13923), .B2(n13924), .A(n9787), .ZN(n14307) );
  INV_X1 U17152 ( .A(n13925), .ZN(n13928) );
  NAND2_X1 U17153 ( .A1(n13938), .A2(n13926), .ZN(n13927) );
  NAND2_X1 U17154 ( .A1(n13928), .A2(n13927), .ZN(n14490) );
  INV_X1 U17155 ( .A(n14490), .ZN(n13934) );
  NOR2_X1 U17156 ( .A1(n13929), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n13933) );
  AOI22_X1 U17157 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n20024), .B1(
        n20027), .B2(n14300), .ZN(n13931) );
  NAND2_X1 U17158 ( .A1(n20021), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n13930) );
  OAI211_X1 U17159 ( .C1(n13941), .C2(n20832), .A(n13931), .B(n13930), .ZN(
        n13932) );
  AOI211_X1 U17160 ( .C1(n13934), .C2(n20025), .A(n13933), .B(n13932), .ZN(
        n13935) );
  OAI21_X1 U17161 ( .B1(n14307), .B2(n19996), .A(n13935), .ZN(P1_U2811) );
  NAND2_X1 U17162 ( .A1(n13951), .A2(n13936), .ZN(n13937) );
  NAND2_X1 U17163 ( .A1(n13938), .A2(n13937), .ZN(n14491) );
  AOI21_X1 U17164 ( .B1(n13940), .B2(n13939), .A(n13923), .ZN(n14320) );
  NAND2_X1 U17165 ( .A1(n14320), .A2(n19980), .ZN(n13948) );
  INV_X1 U17166 ( .A(n13941), .ZN(n13946) );
  INV_X1 U17167 ( .A(n14318), .ZN(n13942) );
  AOI22_X1 U17168 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n20024), .B1(
        n20027), .B2(n13942), .ZN(n13943) );
  OAI21_X1 U17169 ( .B1(n20009), .B2(n14161), .A(n13943), .ZN(n13945) );
  NOR3_X1 U17170 ( .A1(n13955), .A2(P1_REIP_REG_28__SCAN_IN), .A3(n13959), 
        .ZN(n13944) );
  AOI211_X1 U17171 ( .C1(P1_REIP_REG_28__SCAN_IN), .C2(n13946), .A(n13945), 
        .B(n13944), .ZN(n13947) );
  OAI211_X1 U17172 ( .C1(n14491), .C2(n19978), .A(n13948), .B(n13947), .ZN(
        P1_U2812) );
  NAND2_X1 U17173 ( .A1(n13965), .A2(n13949), .ZN(n13950) );
  NAND2_X1 U17174 ( .A1(n13951), .A2(n13950), .ZN(n14503) );
  INV_X1 U17175 ( .A(n14326), .ZN(n13954) );
  NAND2_X1 U17176 ( .A1(n13954), .A2(n19980), .ZN(n13962) );
  INV_X1 U17177 ( .A(n13955), .ZN(n13960) );
  AOI22_X1 U17178 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n20024), .B1(
        n20027), .B2(n14329), .ZN(n13957) );
  NAND2_X1 U17179 ( .A1(n20021), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n13956) );
  OAI211_X1 U17180 ( .C1(n13970), .C2(n13959), .A(n13957), .B(n13956), .ZN(
        n13958) );
  AOI21_X1 U17181 ( .B1(n13960), .B2(n13959), .A(n13958), .ZN(n13961) );
  OAI211_X1 U17182 ( .C1(n19978), .C2(n14503), .A(n13962), .B(n13961), .ZN(
        P1_U2813) );
  OR2_X1 U17183 ( .A1(n13980), .A2(n13963), .ZN(n13964) );
  NAND2_X1 U17184 ( .A1(n13965), .A2(n13964), .ZN(n14517) );
  AOI21_X1 U17185 ( .B1(n13967), .B2(n13977), .A(n13952), .ZN(n14339) );
  NAND2_X1 U17186 ( .A1(n14339), .A2(n19980), .ZN(n13975) );
  OAI22_X1 U17187 ( .A1(n13968), .A2(n20006), .B1(n20016), .B2(n14337), .ZN(
        n13973) );
  INV_X1 U17188 ( .A(n13969), .ZN(n13971) );
  INV_X1 U17189 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n14335) );
  AOI21_X1 U17190 ( .B1(n13971), .B2(n14335), .A(n13970), .ZN(n13972) );
  AOI211_X1 U17191 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n20021), .A(n13973), .B(
        n13972), .ZN(n13974) );
  OAI211_X1 U17192 ( .C1(n14517), .C2(n19978), .A(n13975), .B(n13974), .ZN(
        P1_U2814) );
  OAI21_X1 U17193 ( .B1(n13976), .B2(n13978), .A(n13977), .ZN(n14347) );
  AND2_X1 U17194 ( .A1(n9777), .A2(n13979), .ZN(n13981) );
  OR2_X1 U17195 ( .A1(n13981), .A2(n13980), .ZN(n14164) );
  INV_X1 U17196 ( .A(n14164), .ZN(n14524) );
  INV_X1 U17197 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14165) );
  INV_X1 U17198 ( .A(n13997), .ZN(n13983) );
  OAI211_X1 U17199 ( .C1(P1_REIP_REG_24__SCAN_IN), .C2(P1_REIP_REG_25__SCAN_IN), .A(n13983), .B(n13982), .ZN(n13987) );
  NAND3_X1 U17200 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n14112), .A3(n13992), 
        .ZN(n13984) );
  OAI21_X1 U17201 ( .B1(n20006), .B2(n14346), .A(n13984), .ZN(n13985) );
  AOI21_X1 U17202 ( .B1(n14350), .B2(n20027), .A(n13985), .ZN(n13986) );
  OAI211_X1 U17203 ( .C1(n14165), .C2(n20009), .A(n13987), .B(n13986), .ZN(
        n13988) );
  AOI21_X1 U17204 ( .B1(n14524), .B2(n20025), .A(n13988), .ZN(n13989) );
  OAI21_X1 U17205 ( .B1(n14347), .B2(n19996), .A(n13989), .ZN(P1_U2815) );
  AOI21_X1 U17206 ( .B1(n13991), .B2(n14005), .A(n13976), .ZN(n14358) );
  INV_X1 U17207 ( .A(n14358), .ZN(n14239) );
  INV_X1 U17208 ( .A(n14112), .ZN(n14156) );
  INV_X1 U17209 ( .A(n13992), .ZN(n13993) );
  NOR2_X1 U17210 ( .A1(n14156), .A2(n13993), .ZN(n14007) );
  OAI22_X1 U17211 ( .A1(n13994), .A2(n20006), .B1(n20016), .B2(n14356), .ZN(
        n13995) );
  AOI21_X1 U17212 ( .B1(n20021), .B2(P1_EBX_REG_24__SCAN_IN), .A(n13995), .ZN(
        n13996) );
  OAI21_X1 U17213 ( .B1(n13997), .B2(P1_REIP_REG_24__SCAN_IN), .A(n13996), 
        .ZN(n14001) );
  NAND2_X1 U17214 ( .A1(n9806), .A2(n13998), .ZN(n13999) );
  NAND2_X1 U17215 ( .A1(n9777), .A2(n13999), .ZN(n14539) );
  NOR2_X1 U17216 ( .A1(n14539), .A2(n19978), .ZN(n14000) );
  AOI211_X1 U17217 ( .C1(P1_REIP_REG_24__SCAN_IN), .C2(n14007), .A(n14001), 
        .B(n14000), .ZN(n14002) );
  OAI21_X1 U17218 ( .B1(n14239), .B2(n19996), .A(n14002), .ZN(P1_U2816) );
  OR2_X1 U17219 ( .A1(n14017), .A2(n14003), .ZN(n14004) );
  NAND2_X1 U17220 ( .A1(n9806), .A2(n14004), .ZN(n14547) );
  AOI21_X1 U17221 ( .B1(n14006), .B2(n9756), .A(n13990), .ZN(n14365) );
  NAND2_X1 U17222 ( .A1(n14365), .A2(n19980), .ZN(n14014) );
  OAI22_X1 U17223 ( .A1(n21122), .A2(n20006), .B1(n20016), .B2(n14363), .ZN(
        n14012) );
  INV_X1 U17224 ( .A(n14007), .ZN(n14010) );
  INV_X1 U17225 ( .A(n14025), .ZN(n14008) );
  AOI21_X1 U17226 ( .B1(n14008), .B2(P1_REIP_REG_22__SCAN_IN), .A(
        P1_REIP_REG_23__SCAN_IN), .ZN(n14009) );
  NOR2_X1 U17227 ( .A1(n14010), .A2(n14009), .ZN(n14011) );
  AOI211_X1 U17228 ( .C1(n20021), .C2(P1_EBX_REG_23__SCAN_IN), .A(n14012), .B(
        n14011), .ZN(n14013) );
  OAI211_X1 U17229 ( .C1(n14547), .C2(n19978), .A(n14014), .B(n14013), .ZN(
        P1_U2817) );
  OAI21_X1 U17230 ( .B1(n14015), .B2(n14016), .A(n9756), .ZN(n14375) );
  INV_X1 U17231 ( .A(n14017), .ZN(n14018) );
  OAI21_X1 U17232 ( .B1(n14035), .B2(n14019), .A(n14018), .ZN(n14573) );
  INV_X1 U17233 ( .A(n14573), .ZN(n14028) );
  INV_X1 U17234 ( .A(n14038), .ZN(n14020) );
  NAND2_X1 U17235 ( .A1(n19982), .A2(n14020), .ZN(n14021) );
  NAND2_X1 U17236 ( .A1(n14112), .A2(n14021), .ZN(n15852) );
  NAND2_X1 U17237 ( .A1(n20005), .A2(n14043), .ZN(n14037) );
  INV_X1 U17238 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n14367) );
  AOI21_X1 U17239 ( .B1(n15852), .B2(n14037), .A(n14367), .ZN(n14027) );
  OAI22_X1 U17240 ( .A1(n14022), .A2(n20006), .B1(n20016), .B2(n14368), .ZN(
        n14023) );
  AOI21_X1 U17241 ( .B1(n20021), .B2(P1_EBX_REG_22__SCAN_IN), .A(n14023), .ZN(
        n14024) );
  OAI21_X1 U17242 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n14025), .A(n14024), 
        .ZN(n14026) );
  AOI211_X1 U17243 ( .C1(n14028), .C2(n20025), .A(n14027), .B(n14026), .ZN(
        n14029) );
  OAI21_X1 U17244 ( .B1(n14375), .B2(n19996), .A(n14029), .ZN(P1_U2818) );
  AOI21_X1 U17245 ( .B1(n14032), .B2(n14031), .A(n14015), .ZN(n14381) );
  INV_X1 U17246 ( .A(n14381), .ZN(n14253) );
  INV_X1 U17247 ( .A(n14170), .ZN(n14034) );
  AOI21_X1 U17248 ( .B1(n14034), .B2(n14169), .A(n14033), .ZN(n14036) );
  NOR2_X1 U17249 ( .A1(n14036), .A2(n14035), .ZN(n14579) );
  NOR2_X1 U17250 ( .A1(n14038), .A2(n14037), .ZN(n14040) );
  NOR2_X1 U17251 ( .A1(n20006), .A2(n14382), .ZN(n14039) );
  AOI211_X1 U17252 ( .C1(n20027), .C2(n14384), .A(n14040), .B(n14039), .ZN(
        n14042) );
  NAND2_X1 U17253 ( .A1(n20021), .A2(P1_EBX_REG_21__SCAN_IN), .ZN(n14041) );
  OAI211_X1 U17254 ( .C1(n14043), .C2(n15852), .A(n14042), .B(n14041), .ZN(
        n14044) );
  AOI21_X1 U17255 ( .B1(n14579), .B2(n20025), .A(n14044), .ZN(n14045) );
  OAI21_X1 U17256 ( .B1(n14253), .B2(n19996), .A(n14045), .ZN(P1_U2819) );
  AOI21_X1 U17257 ( .B1(n14049), .B2(n14046), .A(n14048), .ZN(n14401) );
  INV_X1 U17258 ( .A(n14401), .ZN(n14262) );
  INV_X1 U17259 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n14050) );
  NAND2_X1 U17260 ( .A1(n20005), .A2(n14051), .ZN(n14052) );
  NOR2_X1 U17261 ( .A1(n14050), .A2(n14052), .ZN(n15851) );
  INV_X1 U17262 ( .A(n15851), .ZN(n14054) );
  AOI21_X1 U17263 ( .B1(n14051), .B2(n19982), .A(n14156), .ZN(n15861) );
  NOR2_X1 U17264 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n14052), .ZN(n15860) );
  NOR2_X1 U17265 ( .A1(n15861), .A2(n15860), .ZN(n14053) );
  MUX2_X1 U17266 ( .A(n14054), .B(n14053), .S(P1_REIP_REG_19__SCAN_IN), .Z(
        n14062) );
  NAND2_X1 U17267 ( .A1(n20027), .A2(n14397), .ZN(n14055) );
  OAI211_X1 U17268 ( .C1(n20006), .C2(n14399), .A(n14055), .B(n19990), .ZN(
        n14060) );
  INV_X1 U17269 ( .A(n14178), .ZN(n14058) );
  INV_X1 U17270 ( .A(n14056), .ZN(n14057) );
  OAI21_X1 U17271 ( .B1(n14058), .B2(n14057), .A(n14170), .ZN(n14595) );
  NOR2_X1 U17272 ( .A1(n14595), .A2(n19978), .ZN(n14059) );
  AOI211_X1 U17273 ( .C1(P1_EBX_REG_19__SCAN_IN), .C2(n20021), .A(n14060), .B(
        n14059), .ZN(n14061) );
  OAI211_X1 U17274 ( .C1(n14262), .C2(n19996), .A(n14062), .B(n14061), .ZN(
        P1_U2821) );
  INV_X1 U17275 ( .A(n14064), .ZN(n14065) );
  OAI21_X1 U17276 ( .B1(n14063), .B2(n14066), .A(n14065), .ZN(n14417) );
  OAI21_X1 U17277 ( .B1(n19994), .B2(n14067), .A(n20814), .ZN(n14074) );
  INV_X1 U17278 ( .A(n15872), .ZN(n14085) );
  AOI21_X1 U17279 ( .B1(n14085), .B2(n15871), .A(n14068), .ZN(n14069) );
  OR2_X1 U17280 ( .A1(n14069), .A2(n14176), .ZN(n15959) );
  OAI21_X1 U17281 ( .B1(n20006), .B2(n14415), .A(n19990), .ZN(n14071) );
  INV_X1 U17282 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n21043) );
  NOR2_X1 U17283 ( .A1(n20009), .A2(n21043), .ZN(n14070) );
  AOI211_X1 U17284 ( .C1(n20027), .C2(n14420), .A(n14071), .B(n14070), .ZN(
        n14072) );
  OAI21_X1 U17285 ( .B1(n15959), .B2(n19978), .A(n14072), .ZN(n14073) );
  AOI21_X1 U17286 ( .B1(n14074), .B2(n15861), .A(n14073), .ZN(n14075) );
  OAI21_X1 U17287 ( .B1(n14417), .B2(n19996), .A(n14075), .ZN(P1_U2823) );
  AOI21_X1 U17288 ( .B1(n14078), .B2(n14076), .A(n10170), .ZN(n14429) );
  INV_X1 U17289 ( .A(n14429), .ZN(n14281) );
  INV_X1 U17290 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n14093) );
  INV_X1 U17291 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20810) );
  NAND2_X1 U17292 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14113) );
  NAND4_X1 U17293 ( .A1(n20005), .A2(P1_REIP_REG_10__SCAN_IN), .A3(
        P1_REIP_REG_9__SCAN_IN), .A4(n14123), .ZN(n15880) );
  OR3_X1 U17294 ( .A1(n20810), .A2(n14113), .A3(n15880), .ZN(n14092) );
  NOR3_X1 U17295 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n14093), .A3(n14092), 
        .ZN(n15874) );
  OAI21_X1 U17296 ( .B1(n14079), .B2(n20003), .A(n14112), .ZN(n14124) );
  INV_X1 U17297 ( .A(n14124), .ZN(n15897) );
  AOI21_X1 U17298 ( .B1(n14080), .B2(n14112), .A(n15897), .ZN(n14081) );
  INV_X1 U17299 ( .A(n14081), .ZN(n15873) );
  AOI22_X1 U17300 ( .A1(n15873), .A2(P1_REIP_REG_15__SCAN_IN), .B1(n20021), 
        .B2(P1_EBX_REG_15__SCAN_IN), .ZN(n14082) );
  OAI211_X1 U17301 ( .C1(n20006), .C2(n14083), .A(n14082), .B(n19990), .ZN(
        n14084) );
  NOR2_X1 U17302 ( .A1(n15874), .A2(n14084), .ZN(n14089) );
  AOI21_X1 U17303 ( .B1(n14086), .B2(n14096), .A(n14085), .ZN(n15981) );
  INV_X1 U17304 ( .A(n14427), .ZN(n14087) );
  AOI22_X1 U17305 ( .A1(n15981), .A2(n20025), .B1(n20027), .B2(n14087), .ZN(
        n14088) );
  OAI211_X1 U17306 ( .C1(n14281), .C2(n19996), .A(n14089), .B(n14088), .ZN(
        P1_U2825) );
  OAI21_X1 U17307 ( .B1(n14090), .B2(n14091), .A(n14076), .ZN(n14283) );
  NAND2_X1 U17308 ( .A1(n14093), .A2(n14092), .ZN(n14101) );
  OR2_X1 U17309 ( .A1(n14109), .A2(n14094), .ZN(n14095) );
  NAND2_X1 U17310 ( .A1(n14096), .A2(n14095), .ZN(n15985) );
  NOR2_X1 U17311 ( .A1(n15985), .A2(n19978), .ZN(n14100) );
  AOI21_X1 U17312 ( .B1(n20027), .B2(n15926), .A(n20123), .ZN(n14098) );
  NAND2_X1 U17313 ( .A1(n20024), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14097) );
  OAI211_X1 U17314 ( .C1(n20009), .C2(n14183), .A(n14098), .B(n14097), .ZN(
        n14099) );
  AOI211_X1 U17315 ( .C1(n15873), .C2(n14101), .A(n14100), .B(n14099), .ZN(
        n14102) );
  OAI21_X1 U17316 ( .B1(n14283), .B2(n19996), .A(n14102), .ZN(P1_U2826) );
  OAI21_X1 U17317 ( .B1(n10186), .B2(n11446), .A(n14104), .ZN(n15898) );
  OAI21_X1 U17318 ( .B1(n15898), .B2(n15899), .A(n14104), .ZN(n14193) );
  NAND2_X1 U17319 ( .A1(n14193), .A2(n14192), .ZN(n14191) );
  INV_X1 U17320 ( .A(n14105), .ZN(n14106) );
  AOI21_X1 U17321 ( .B1(n14191), .B2(n14106), .A(n14090), .ZN(n14442) );
  INV_X1 U17322 ( .A(n14442), .ZN(n14288) );
  INV_X1 U17323 ( .A(n14440), .ZN(n14118) );
  AND2_X1 U17324 ( .A1(n14190), .A2(n14107), .ZN(n14108) );
  NOR2_X1 U17325 ( .A1(n14109), .A2(n14108), .ZN(n15995) );
  AOI22_X1 U17326 ( .A1(n15995), .A2(n20025), .B1(n20021), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14110) );
  OAI211_X1 U17327 ( .C1(n20006), .C2(n14111), .A(n14110), .B(n19990), .ZN(
        n14117) );
  NOR2_X1 U17328 ( .A1(n14113), .A2(n15880), .ZN(n14115) );
  AOI21_X1 U17329 ( .B1(n14113), .B2(n14112), .A(n15897), .ZN(n15889) );
  INV_X1 U17330 ( .A(n15889), .ZN(n14114) );
  MUX2_X1 U17331 ( .A(n14115), .B(n14114), .S(P1_REIP_REG_13__SCAN_IN), .Z(
        n14116) );
  AOI211_X1 U17332 ( .C1(n20027), .C2(n14118), .A(n14117), .B(n14116), .ZN(
        n14119) );
  OAI21_X1 U17333 ( .B1(n14288), .B2(n19996), .A(n14119), .ZN(P1_U2827) );
  OAI21_X1 U17334 ( .B1(n20016), .B2(n14446), .A(n19990), .ZN(n14120) );
  AOI21_X1 U17335 ( .B1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n20024), .A(
        n14120), .ZN(n14121) );
  OAI21_X1 U17336 ( .B1(n14122), .B2(n20009), .A(n14121), .ZN(n14127) );
  INV_X1 U17337 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20805) );
  NAND3_X1 U17338 ( .A1(n20005), .A2(P1_REIP_REG_9__SCAN_IN), .A3(n14123), 
        .ZN(n14125) );
  AOI21_X1 U17339 ( .B1(n20805), .B2(n14125), .A(n14124), .ZN(n14126) );
  AOI211_X1 U17340 ( .C1(n16009), .C2(n20025), .A(n14127), .B(n14126), .ZN(
        n14128) );
  OAI21_X1 U17341 ( .B1(n14450), .B2(n19996), .A(n14128), .ZN(P1_U2830) );
  OAI21_X1 U17342 ( .B1(n19994), .B2(n14129), .A(n20803), .ZN(n14136) );
  AOI21_X1 U17343 ( .B1(n20024), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n20123), .ZN(n14130) );
  OAI21_X1 U17344 ( .B1(n14131), .B2(n20016), .A(n14130), .ZN(n14132) );
  AOI21_X1 U17345 ( .B1(P1_EBX_REG_8__SCAN_IN), .B2(n20021), .A(n14132), .ZN(
        n14133) );
  OAI21_X1 U17346 ( .B1(n19978), .B2(n16020), .A(n14133), .ZN(n14134) );
  AOI21_X1 U17347 ( .B1(n14136), .B2(n14135), .A(n14134), .ZN(n14137) );
  OAI21_X1 U17348 ( .B1(n14138), .B2(n19996), .A(n14137), .ZN(P1_U2832) );
  OAI22_X1 U17349 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n19994), .B1(n20009), 
        .B2(n14139), .ZN(n14144) );
  OAI22_X1 U17350 ( .A1(n20016), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n14140), .B2(n19982), .ZN(n14141) );
  AOI21_X1 U17351 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20024), .A(
        n14141), .ZN(n14142) );
  OAI21_X1 U17352 ( .B1(n9741), .B2(n20018), .A(n14142), .ZN(n14143) );
  AOI211_X1 U17353 ( .C1(n20025), .C2(n13192), .A(n14144), .B(n14143), .ZN(
        n14145) );
  OAI21_X1 U17354 ( .B1(n14150), .B2(n14146), .A(n14145), .ZN(P1_U2839) );
  INV_X1 U17355 ( .A(n20284), .ZN(n14148) );
  OAI21_X1 U17356 ( .B1(n20024), .B2(n20027), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14147) );
  OAI21_X1 U17357 ( .B1(n20018), .B2(n14148), .A(n14147), .ZN(n14153) );
  OAI22_X1 U17358 ( .A1(n19978), .A2(n14151), .B1(n14150), .B2(n14149), .ZN(
        n14152) );
  AOI211_X1 U17359 ( .C1(P1_EBX_REG_0__SCAN_IN), .C2(n20021), .A(n14153), .B(
        n14152), .ZN(n14154) );
  OAI21_X1 U17360 ( .B1(n14156), .B2(n14155), .A(n14154), .ZN(P1_U2840) );
  INV_X1 U17361 ( .A(n14472), .ZN(n14158) );
  OAI22_X1 U17362 ( .A1(n14158), .A2(n14196), .B1(n14157), .B2(n20040), .ZN(
        P1_U2841) );
  INV_X1 U17363 ( .A(n14296), .ZN(n14205) );
  OAI222_X1 U17364 ( .A1(n14194), .A2(n14205), .B1(n20040), .B2(n14159), .C1(
        n14477), .C2(n14196), .ZN(P1_U2842) );
  OAI222_X1 U17365 ( .A1(n14160), .A2(n20040), .B1(n14196), .B2(n14490), .C1(
        n14307), .C2(n14194), .ZN(P1_U2843) );
  INV_X1 U17366 ( .A(n14320), .ZN(n14219) );
  OAI222_X1 U17367 ( .A1(n14161), .A2(n20040), .B1(n14196), .B2(n14491), .C1(
        n14219), .C2(n14194), .ZN(P1_U2844) );
  INV_X1 U17368 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14162) );
  OAI222_X1 U17369 ( .A1(n14162), .A2(n20040), .B1(n14196), .B2(n14503), .C1(
        n14326), .C2(n14194), .ZN(P1_U2845) );
  INV_X1 U17370 ( .A(n14339), .ZN(n14231) );
  OAI222_X1 U17371 ( .A1(n14163), .A2(n20040), .B1(n14196), .B2(n14517), .C1(
        n14231), .C2(n14194), .ZN(P1_U2846) );
  OAI222_X1 U17372 ( .A1(n14165), .A2(n20040), .B1(n14196), .B2(n14164), .C1(
        n14347), .C2(n14194), .ZN(P1_U2847) );
  INV_X1 U17373 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14166) );
  OAI222_X1 U17374 ( .A1(n14166), .A2(n20040), .B1(n14196), .B2(n14539), .C1(
        n14239), .C2(n14194), .ZN(P1_U2848) );
  INV_X1 U17375 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n20958) );
  INV_X1 U17376 ( .A(n14365), .ZN(n14244) );
  OAI222_X1 U17377 ( .A1(n14547), .A2(n14196), .B1(n20040), .B2(n20958), .C1(
        n14194), .C2(n14244), .ZN(P1_U2849) );
  OAI222_X1 U17378 ( .A1(n14573), .A2(n14196), .B1(n14167), .B2(n20040), .C1(
        n14375), .C2(n14194), .ZN(P1_U2850) );
  AOI22_X1 U17379 ( .A1(n14579), .A2(n20036), .B1(n14186), .B2(
        P1_EBX_REG_21__SCAN_IN), .ZN(n14168) );
  OAI21_X1 U17380 ( .B1(n14253), .B2(n14194), .A(n14168), .ZN(P1_U2851) );
  OAI21_X1 U17381 ( .B1(n14048), .B2(n10261), .A(n14031), .ZN(n15854) );
  XNOR2_X1 U17382 ( .A(n14170), .B(n14169), .ZN(n15856) );
  AOI22_X1 U17383 ( .A1(n15856), .A2(n20036), .B1(n14186), .B2(
        P1_EBX_REG_20__SCAN_IN), .ZN(n14171) );
  OAI21_X1 U17384 ( .B1(n15854), .B2(n14194), .A(n14171), .ZN(P1_U2852) );
  INV_X1 U17385 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14172) );
  OAI222_X1 U17386 ( .A1(n14595), .A2(n14196), .B1(n14172), .B2(n20040), .C1(
        n14262), .C2(n14194), .ZN(P1_U2853) );
  OR2_X1 U17387 ( .A1(n14064), .A2(n14173), .ZN(n14174) );
  AND2_X1 U17388 ( .A1(n14046), .A2(n14174), .ZN(n15866) );
  OR2_X1 U17389 ( .A1(n14176), .A2(n14175), .ZN(n14177) );
  NAND2_X1 U17390 ( .A1(n14178), .A2(n14177), .ZN(n15864) );
  OAI22_X1 U17391 ( .A1(n15864), .A2(n14196), .B1(n14179), .B2(n20040), .ZN(
        n14180) );
  INV_X1 U17392 ( .A(n14180), .ZN(n14181) );
  OAI21_X1 U17393 ( .B1(n14408), .B2(n14194), .A(n14181), .ZN(P1_U2854) );
  OAI222_X1 U17394 ( .A1(n15959), .A2(n14196), .B1(n20040), .B2(n21043), .C1(
        n14194), .C2(n14417), .ZN(P1_U2855) );
  AOI22_X1 U17395 ( .A1(n15981), .A2(n20036), .B1(n14186), .B2(
        P1_EBX_REG_15__SCAN_IN), .ZN(n14182) );
  OAI21_X1 U17396 ( .B1(n14281), .B2(n14194), .A(n14182), .ZN(P1_U2857) );
  INV_X1 U17397 ( .A(n14283), .ZN(n15927) );
  OAI22_X1 U17398 ( .A1(n15985), .A2(n14196), .B1(n14183), .B2(n20040), .ZN(
        n14184) );
  AOI21_X1 U17399 ( .B1(n15927), .B2(n20037), .A(n14184), .ZN(n14185) );
  INV_X1 U17400 ( .A(n14185), .ZN(P1_U2858) );
  AOI22_X1 U17401 ( .A1(n15995), .A2(n20036), .B1(n14186), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14187) );
  OAI21_X1 U17402 ( .B1(n14288), .B2(n14194), .A(n14187), .ZN(P1_U2859) );
  NAND2_X1 U17403 ( .A1(n15893), .A2(n14188), .ZN(n14189) );
  NAND2_X1 U17404 ( .A1(n14190), .A2(n14189), .ZN(n15882) );
  INV_X1 U17405 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14195) );
  OAI21_X1 U17406 ( .B1(n14193), .B2(n14192), .A(n14191), .ZN(n15885) );
  OAI222_X1 U17407 ( .A1(n15882), .A2(n14196), .B1(n14195), .B2(n20040), .C1(
        n15885), .C2(n14194), .ZN(P1_U2860) );
  OR2_X1 U17408 ( .A1(n14221), .A2(n14199), .ZN(n14201) );
  NAND2_X1 U17409 ( .A1(n20160), .A2(DATAI_14_), .ZN(n14200) );
  NAND2_X1 U17410 ( .A1(n14201), .A2(n14200), .ZN(n20092) );
  AOI22_X1 U17411 ( .A1(n14273), .A2(n20092), .B1(n14289), .B2(
        P1_EAX_REG_30__SCAN_IN), .ZN(n14202) );
  OAI21_X1 U17412 ( .B1(n14276), .B2(n19241), .A(n14202), .ZN(n14203) );
  AOI21_X1 U17413 ( .B1(n14278), .B2(DATAI_30_), .A(n14203), .ZN(n14204) );
  OAI21_X1 U17414 ( .B1(n14205), .B2(n14287), .A(n14204), .ZN(P1_U2874) );
  INV_X1 U17415 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n14210) );
  OR2_X1 U17416 ( .A1(n14221), .A2(n14206), .ZN(n14208) );
  NAND2_X1 U17417 ( .A1(n20160), .A2(DATAI_13_), .ZN(n14207) );
  NAND2_X1 U17418 ( .A1(n14208), .A2(n14207), .ZN(n20090) );
  AOI22_X1 U17419 ( .A1(n14273), .A2(n20090), .B1(n14289), .B2(
        P1_EAX_REG_29__SCAN_IN), .ZN(n14209) );
  OAI21_X1 U17420 ( .B1(n14276), .B2(n14210), .A(n14209), .ZN(n14211) );
  AOI21_X1 U17421 ( .B1(n14278), .B2(DATAI_29_), .A(n14211), .ZN(n14212) );
  OAI21_X1 U17422 ( .B1(n14307), .B2(n14287), .A(n14212), .ZN(P1_U2875) );
  INV_X1 U17423 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n19231) );
  OR2_X1 U17424 ( .A1(n14221), .A2(n14213), .ZN(n14215) );
  NAND2_X1 U17425 ( .A1(n14221), .A2(DATAI_12_), .ZN(n14214) );
  NAND2_X1 U17426 ( .A1(n14215), .A2(n14214), .ZN(n20088) );
  AOI22_X1 U17427 ( .A1(n14273), .A2(n20088), .B1(n14289), .B2(
        P1_EAX_REG_28__SCAN_IN), .ZN(n14216) );
  OAI21_X1 U17428 ( .B1(n14276), .B2(n19231), .A(n14216), .ZN(n14217) );
  AOI21_X1 U17429 ( .B1(n14278), .B2(DATAI_28_), .A(n14217), .ZN(n14218) );
  OAI21_X1 U17430 ( .B1(n14219), .B2(n14287), .A(n14218), .ZN(P1_U2876) );
  INV_X1 U17431 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n14225) );
  OR2_X1 U17432 ( .A1(n14221), .A2(n14220), .ZN(n14223) );
  NAND2_X1 U17433 ( .A1(n14221), .A2(DATAI_11_), .ZN(n14222) );
  NAND2_X1 U17434 ( .A1(n14223), .A2(n14222), .ZN(n20086) );
  AOI22_X1 U17435 ( .A1(n14273), .A2(n20086), .B1(n14289), .B2(
        P1_EAX_REG_27__SCAN_IN), .ZN(n14224) );
  OAI21_X1 U17436 ( .B1(n14276), .B2(n14225), .A(n14224), .ZN(n14226) );
  AOI21_X1 U17437 ( .B1(n14278), .B2(DATAI_27_), .A(n14226), .ZN(n14227) );
  OAI21_X1 U17438 ( .B1(n14326), .B2(n14287), .A(n14227), .ZN(P1_U2877) );
  INV_X1 U17439 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16425) );
  AOI22_X1 U17440 ( .A1(n14273), .A2(n20084), .B1(n14289), .B2(
        P1_EAX_REG_26__SCAN_IN), .ZN(n14228) );
  OAI21_X1 U17441 ( .B1(n14276), .B2(n16425), .A(n14228), .ZN(n14229) );
  AOI21_X1 U17442 ( .B1(n14278), .B2(DATAI_26_), .A(n14229), .ZN(n14230) );
  OAI21_X1 U17443 ( .B1(n14231), .B2(n14287), .A(n14230), .ZN(P1_U2878) );
  INV_X1 U17444 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n14233) );
  AOI22_X1 U17445 ( .A1(n14273), .A2(n20081), .B1(n14289), .B2(
        P1_EAX_REG_25__SCAN_IN), .ZN(n14232) );
  OAI21_X1 U17446 ( .B1(n14276), .B2(n14233), .A(n14232), .ZN(n14234) );
  AOI21_X1 U17447 ( .B1(n14278), .B2(DATAI_25_), .A(n14234), .ZN(n14235) );
  OAI21_X1 U17448 ( .B1(n14347), .B2(n14287), .A(n14235), .ZN(P1_U2879) );
  INV_X1 U17449 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n19207) );
  AOI22_X1 U17450 ( .A1(n14273), .A2(n20079), .B1(n14289), .B2(
        P1_EAX_REG_24__SCAN_IN), .ZN(n14236) );
  OAI21_X1 U17451 ( .B1(n14276), .B2(n19207), .A(n14236), .ZN(n14237) );
  AOI21_X1 U17452 ( .B1(n14278), .B2(DATAI_24_), .A(n14237), .ZN(n14238) );
  OAI21_X1 U17453 ( .B1(n14239), .B2(n14287), .A(n14238), .ZN(P1_U2880) );
  INV_X1 U17454 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n14241) );
  AOI22_X1 U17455 ( .A1(n14273), .A2(n20214), .B1(n14289), .B2(
        P1_EAX_REG_23__SCAN_IN), .ZN(n14240) );
  OAI21_X1 U17456 ( .B1(n14276), .B2(n14241), .A(n14240), .ZN(n14242) );
  AOI21_X1 U17457 ( .B1(n14278), .B2(DATAI_23_), .A(n14242), .ZN(n14243) );
  OAI21_X1 U17458 ( .B1(n14244), .B2(n14287), .A(n14243), .ZN(P1_U2881) );
  INV_X1 U17459 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n14246) );
  AOI22_X1 U17460 ( .A1(n14273), .A2(n20204), .B1(n14289), .B2(
        P1_EAX_REG_22__SCAN_IN), .ZN(n14245) );
  OAI21_X1 U17461 ( .B1(n14276), .B2(n14246), .A(n14245), .ZN(n14247) );
  AOI21_X1 U17462 ( .B1(n14278), .B2(DATAI_22_), .A(n14247), .ZN(n14248) );
  OAI21_X1 U17463 ( .B1(n14375), .B2(n14287), .A(n14248), .ZN(P1_U2882) );
  INV_X1 U17464 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n14250) );
  AOI22_X1 U17465 ( .A1(n14273), .A2(n20200), .B1(n14289), .B2(
        P1_EAX_REG_21__SCAN_IN), .ZN(n14249) );
  OAI21_X1 U17466 ( .B1(n14276), .B2(n14250), .A(n14249), .ZN(n14251) );
  AOI21_X1 U17467 ( .B1(n14278), .B2(DATAI_21_), .A(n14251), .ZN(n14252) );
  OAI21_X1 U17468 ( .B1(n14253), .B2(n14287), .A(n14252), .ZN(P1_U2883) );
  INV_X1 U17469 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n14255) );
  AOI22_X1 U17470 ( .A1(n14273), .A2(n20195), .B1(n14289), .B2(
        P1_EAX_REG_20__SCAN_IN), .ZN(n14254) );
  OAI21_X1 U17471 ( .B1(n14276), .B2(n14255), .A(n14254), .ZN(n14256) );
  AOI21_X1 U17472 ( .B1(n14278), .B2(DATAI_20_), .A(n14256), .ZN(n14257) );
  OAI21_X1 U17473 ( .B1(n15854), .B2(n14287), .A(n14257), .ZN(P1_U2884) );
  INV_X1 U17474 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n14259) );
  AOI22_X1 U17475 ( .A1(n14273), .A2(n20191), .B1(n14289), .B2(
        P1_EAX_REG_19__SCAN_IN), .ZN(n14258) );
  OAI21_X1 U17476 ( .B1(n14276), .B2(n14259), .A(n14258), .ZN(n14260) );
  AOI21_X1 U17477 ( .B1(n14278), .B2(DATAI_19_), .A(n14260), .ZN(n14261) );
  OAI21_X1 U17478 ( .B1(n14262), .B2(n14287), .A(n14261), .ZN(P1_U2885) );
  INV_X1 U17479 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n14264) );
  AOI22_X1 U17480 ( .A1(n14273), .A2(n20186), .B1(n14289), .B2(
        P1_EAX_REG_18__SCAN_IN), .ZN(n14263) );
  OAI21_X1 U17481 ( .B1(n14276), .B2(n14264), .A(n14263), .ZN(n14265) );
  AOI21_X1 U17482 ( .B1(n14278), .B2(DATAI_18_), .A(n14265), .ZN(n14266) );
  OAI21_X1 U17483 ( .B1(n14408), .B2(n14287), .A(n14266), .ZN(P1_U2886) );
  INV_X1 U17484 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n14268) );
  AOI22_X1 U17485 ( .A1(n14273), .A2(n20181), .B1(n14289), .B2(
        P1_EAX_REG_17__SCAN_IN), .ZN(n14267) );
  OAI21_X1 U17486 ( .B1(n14276), .B2(n14268), .A(n14267), .ZN(n14269) );
  AOI21_X1 U17487 ( .B1(n14278), .B2(DATAI_17_), .A(n14269), .ZN(n14270) );
  OAI21_X1 U17488 ( .B1(n14417), .B2(n14287), .A(n14270), .ZN(P1_U2887) );
  AND2_X1 U17489 ( .A1(n14077), .A2(n14271), .ZN(n14272) );
  OR2_X1 U17490 ( .A1(n14272), .A2(n14063), .ZN(n15870) );
  INV_X1 U17491 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n14275) );
  AOI22_X1 U17492 ( .A1(n14273), .A2(n20172), .B1(n14289), .B2(
        P1_EAX_REG_16__SCAN_IN), .ZN(n14274) );
  OAI21_X1 U17493 ( .B1(n14276), .B2(n14275), .A(n14274), .ZN(n14277) );
  AOI21_X1 U17494 ( .B1(n14278), .B2(DATAI_16_), .A(n14277), .ZN(n14279) );
  OAI21_X1 U17495 ( .B1(n15870), .B2(n14287), .A(n14279), .ZN(P1_U2888) );
  OAI222_X1 U17496 ( .A1(n14281), .A2(n14287), .B1(n14285), .B2(n14280), .C1(
        n15908), .C2(n12857), .ZN(P1_U2889) );
  AOI22_X1 U17497 ( .A1(n15905), .A2(n20092), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14289), .ZN(n14282) );
  OAI21_X1 U17498 ( .B1(n14283), .B2(n14287), .A(n14282), .ZN(P1_U2890) );
  INV_X1 U17499 ( .A(n20090), .ZN(n14286) );
  OAI222_X1 U17500 ( .A1(n14288), .A2(n14287), .B1(n14286), .B2(n14285), .C1(
        n14284), .C2(n15908), .ZN(P1_U2891) );
  AOI22_X1 U17501 ( .A1(n15905), .A2(n20088), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n14289), .ZN(n14290) );
  OAI21_X1 U17502 ( .B1(n15885), .B2(n14287), .A(n14290), .ZN(P1_U2892) );
  NOR2_X1 U17503 ( .A1(n19990), .A2(n14292), .ZN(n14478) );
  AOI21_X1 U17504 ( .B1(n20111), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14478), .ZN(n14293) );
  OAI21_X1 U17505 ( .B1(n20122), .B2(n14294), .A(n14293), .ZN(n14295) );
  AOI21_X1 U17506 ( .B1(n14296), .B2(n20117), .A(n14295), .ZN(n14297) );
  OAI21_X1 U17507 ( .B1(n14481), .B2(n19955), .A(n14297), .ZN(P1_U2969) );
  NOR2_X1 U17508 ( .A1(n19990), .A2(n20832), .ZN(n14486) );
  NOR2_X1 U17509 ( .A1(n14416), .A2(n14298), .ZN(n14299) );
  AOI211_X1 U17510 ( .C1(n15932), .C2(n14300), .A(n14486), .B(n14299), .ZN(
        n14306) );
  INV_X1 U17511 ( .A(n14301), .ZN(n14302) );
  MUX2_X1 U17512 ( .A(n14303), .B(n14302), .S(n14411), .Z(n14304) );
  NAND2_X1 U17513 ( .A1(n14482), .A2(n20118), .ZN(n14305) );
  OAI211_X1 U17514 ( .C1(n14307), .C2(n20161), .A(n14306), .B(n14305), .ZN(
        P1_U2970) );
  NOR3_X1 U17515 ( .A1(n9721), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14309), .ZN(n14313) );
  NOR2_X1 U17516 ( .A1(n14411), .A2(n14310), .ZN(n14331) );
  NOR3_X1 U17517 ( .A1(n14361), .A2(n14331), .A3(n10056), .ZN(n14312) );
  MUX2_X1 U17518 ( .A(n10056), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n15937), .Z(n14311) );
  OAI21_X1 U17519 ( .B1(n14313), .B2(n14312), .A(n14311), .ZN(n14315) );
  XNOR2_X1 U17520 ( .A(n14315), .B(n14314), .ZN(n14499) );
  NOR2_X1 U17521 ( .A1(n19990), .A2(n14316), .ZN(n14492) );
  AOI21_X1 U17522 ( .B1(n20111), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14492), .ZN(n14317) );
  OAI21_X1 U17523 ( .B1(n20122), .B2(n14318), .A(n14317), .ZN(n14319) );
  AOI21_X1 U17524 ( .B1(n14320), .B2(n20117), .A(n14319), .ZN(n14321) );
  OAI21_X1 U17525 ( .B1(n19955), .B2(n14499), .A(n14321), .ZN(P1_U2971) );
  MUX2_X1 U17526 ( .A(n14323), .B(n14322), .S(n14411), .Z(n14324) );
  XNOR2_X1 U17527 ( .A(n14324), .B(n10056), .ZN(n14508) );
  NAND2_X1 U17528 ( .A1(n20123), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14501) );
  OAI21_X1 U17529 ( .B1(n14416), .B2(n14325), .A(n14501), .ZN(n14328) );
  NOR2_X1 U17530 ( .A1(n14326), .A2(n20161), .ZN(n14327) );
  OAI21_X1 U17531 ( .B1(n19955), .B2(n14508), .A(n14330), .ZN(P1_U2972) );
  INV_X1 U17532 ( .A(n14331), .ZN(n14332) );
  OAI211_X1 U17533 ( .C1(n9721), .C2(n14411), .A(n14333), .B(n14332), .ZN(
        n14334) );
  XNOR2_X1 U17534 ( .A(n14334), .B(n14512), .ZN(n14520) );
  NOR2_X1 U17535 ( .A1(n19990), .A2(n14335), .ZN(n14509) );
  AOI21_X1 U17536 ( .B1(n20111), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14509), .ZN(n14336) );
  OAI21_X1 U17537 ( .B1(n20122), .B2(n14337), .A(n14336), .ZN(n14338) );
  AOI21_X1 U17538 ( .B1(n14339), .B2(n20117), .A(n14338), .ZN(n14340) );
  OAI21_X1 U17539 ( .B1(n19955), .B2(n14520), .A(n14340), .ZN(P1_U2973) );
  NAND2_X1 U17540 ( .A1(n14341), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14353) );
  INV_X1 U17541 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14534) );
  NOR2_X1 U17542 ( .A1(n14353), .A2(n14534), .ZN(n14344) );
  NOR3_X1 U17543 ( .A1(n9721), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14343) );
  MUX2_X1 U17544 ( .A(n14344), .B(n14343), .S(n14342), .Z(n14345) );
  XNOR2_X1 U17545 ( .A(n14345), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14529) );
  NAND2_X1 U17546 ( .A1(n20123), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14521) );
  OAI21_X1 U17547 ( .B1(n14416), .B2(n14346), .A(n14521), .ZN(n14349) );
  NOR2_X1 U17548 ( .A1(n14347), .A2(n20161), .ZN(n14348) );
  AOI211_X1 U17549 ( .C1(n15932), .C2(n14350), .A(n14349), .B(n14348), .ZN(
        n14351) );
  OAI21_X1 U17550 ( .B1(n19955), .B2(n14529), .A(n14351), .ZN(P1_U2974) );
  NAND2_X1 U17551 ( .A1(n14353), .A2(n14361), .ZN(n14352) );
  MUX2_X1 U17552 ( .A(n14353), .B(n14352), .S(n14411), .Z(n14354) );
  XOR2_X1 U17553 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n14354), .Z(
        n14542) );
  NAND2_X1 U17554 ( .A1(n20123), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14538) );
  NAND2_X1 U17555 ( .A1(n20111), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14355) );
  OAI211_X1 U17556 ( .C1(n20122), .C2(n14356), .A(n14538), .B(n14355), .ZN(
        n14357) );
  AOI21_X1 U17557 ( .B1(n14358), .B2(n20117), .A(n14357), .ZN(n14359) );
  OAI21_X1 U17558 ( .B1(n19955), .B2(n14542), .A(n14359), .ZN(P1_U2975) );
  XNOR2_X1 U17559 ( .A(n14411), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14360) );
  XNOR2_X1 U17560 ( .A(n14361), .B(n14360), .ZN(n14552) );
  NAND2_X1 U17561 ( .A1(n20123), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14546) );
  NAND2_X1 U17562 ( .A1(n20111), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14362) );
  OAI211_X1 U17563 ( .C1(n20122), .C2(n14363), .A(n14546), .B(n14362), .ZN(
        n14364) );
  AOI21_X1 U17564 ( .B1(n14365), .B2(n20117), .A(n14364), .ZN(n14366) );
  OAI21_X1 U17565 ( .B1(n14552), .B2(n19955), .A(n14366), .ZN(P1_U2976) );
  NOR2_X1 U17566 ( .A1(n19990), .A2(n14367), .ZN(n14569) );
  NOR2_X1 U17567 ( .A1(n20122), .A2(n14368), .ZN(n14369) );
  AOI211_X1 U17568 ( .C1(n20111), .C2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n14569), .B(n14369), .ZN(n14374) );
  NAND2_X1 U17569 ( .A1(n9720), .A2(n14370), .ZN(n14372) );
  XNOR2_X1 U17570 ( .A(n14372), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14553) );
  NAND2_X1 U17571 ( .A1(n14553), .A2(n20118), .ZN(n14373) );
  OAI211_X1 U17572 ( .C1(n14375), .C2(n20161), .A(n14374), .B(n14373), .ZN(
        P1_U2977) );
  OAI21_X1 U17573 ( .B1(n15937), .B2(n14609), .A(n14601), .ZN(n14396) );
  NAND2_X1 U17574 ( .A1(n14411), .A2(n14377), .ZN(n14394) );
  NAND2_X1 U17575 ( .A1(n15923), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14393) );
  OAI22_X1 U17576 ( .A1(n14396), .A2(n14394), .B1(n14601), .B2(n14393), .ZN(
        n14390) );
  NAND2_X1 U17577 ( .A1(n14390), .A2(n10038), .ZN(n14389) );
  INV_X1 U17578 ( .A(n14393), .ZN(n14378) );
  NAND2_X1 U17579 ( .A1(n14378), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14379) );
  OAI22_X1 U17580 ( .A1(n14389), .A2(n15923), .B1(n14601), .B2(n14379), .ZN(
        n14380) );
  XNOR2_X1 U17581 ( .A(n14380), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14581) );
  NAND2_X1 U17582 ( .A1(n14381), .A2(n20117), .ZN(n14386) );
  NOR2_X1 U17583 ( .A1(n19990), .A2(n14043), .ZN(n14574) );
  NOR2_X1 U17584 ( .A1(n14416), .A2(n14382), .ZN(n14383) );
  AOI211_X1 U17585 ( .C1(n15932), .C2(n14384), .A(n14574), .B(n14383), .ZN(
        n14385) );
  OAI211_X1 U17586 ( .C1(n14581), .C2(n19955), .A(n14386), .B(n14385), .ZN(
        P1_U2978) );
  INV_X1 U17587 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n14387) );
  NOR2_X1 U17588 ( .A1(n19990), .A2(n14387), .ZN(n14586) );
  NOR2_X1 U17589 ( .A1(n20122), .A2(n15859), .ZN(n14388) );
  AOI211_X1 U17590 ( .C1(n20111), .C2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n14586), .B(n14388), .ZN(n14392) );
  OAI21_X1 U17591 ( .B1(n14390), .B2(n10038), .A(n14389), .ZN(n14582) );
  NAND2_X1 U17592 ( .A1(n14582), .A2(n20118), .ZN(n14391) );
  OAI211_X1 U17593 ( .C1(n15854), .C2(n20161), .A(n14392), .B(n14391), .ZN(
        P1_U2979) );
  NAND2_X1 U17594 ( .A1(n14394), .A2(n14393), .ZN(n14395) );
  XNOR2_X1 U17595 ( .A(n14396), .B(n14395), .ZN(n14600) );
  NAND2_X1 U17596 ( .A1(n15932), .A2(n14397), .ZN(n14398) );
  NAND2_X1 U17597 ( .A1(n20123), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n14593) );
  OAI211_X1 U17598 ( .C1(n14416), .C2(n14399), .A(n14398), .B(n14593), .ZN(
        n14400) );
  AOI21_X1 U17599 ( .B1(n14401), .B2(n20117), .A(n14400), .ZN(n14402) );
  OAI21_X1 U17600 ( .B1(n19955), .B2(n14600), .A(n14402), .ZN(P1_U2980) );
  AND2_X1 U17601 ( .A1(n20123), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n14608) );
  NOR2_X1 U17602 ( .A1(n20122), .A2(n15868), .ZN(n14403) );
  AOI211_X1 U17603 ( .C1(n20111), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n14608), .B(n14403), .ZN(n14407) );
  OR2_X1 U17604 ( .A1(n14405), .A2(n14404), .ZN(n14602) );
  NAND3_X1 U17605 ( .A1(n14602), .A2(n14601), .A3(n20118), .ZN(n14406) );
  OAI211_X1 U17606 ( .C1(n14408), .C2(n20161), .A(n14407), .B(n14406), .ZN(
        P1_U2981) );
  AOI21_X1 U17607 ( .B1(n15936), .B2(n15909), .A(n14410), .ZN(n14413) );
  NOR2_X1 U17608 ( .A1(n14413), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14412) );
  MUX2_X1 U17609 ( .A(n14413), .B(n14412), .S(n14411), .Z(n14414) );
  XNOR2_X1 U17610 ( .A(n14414), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15958) );
  OAI22_X1 U17611 ( .A1(n14416), .A2(n14415), .B1(n19990), .B2(n20814), .ZN(
        n14419) );
  NOR2_X1 U17612 ( .A1(n14417), .A2(n20161), .ZN(n14418) );
  AOI211_X1 U17613 ( .C1(n15932), .C2(n14420), .A(n14419), .B(n14418), .ZN(
        n14421) );
  OAI21_X1 U17614 ( .B1(n19955), .B2(n15958), .A(n14421), .ZN(P1_U2982) );
  NOR2_X1 U17615 ( .A1(n15936), .A2(n14422), .ZN(n15912) );
  NOR3_X1 U17616 ( .A1(n15912), .A2(n15920), .A3(n14423), .ZN(n14425) );
  INV_X1 U17617 ( .A(n15910), .ZN(n14424) );
  XNOR2_X1 U17618 ( .A(n14425), .B(n9814), .ZN(n15979) );
  INV_X1 U17619 ( .A(n15979), .ZN(n14431) );
  AOI22_X1 U17620 ( .A1(n20111), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20123), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n14426) );
  OAI21_X1 U17621 ( .B1(n20122), .B2(n14427), .A(n14426), .ZN(n14428) );
  AOI21_X1 U17622 ( .B1(n14429), .B2(n20117), .A(n14428), .ZN(n14430) );
  OAI21_X1 U17623 ( .B1(n14431), .B2(n19955), .A(n14430), .ZN(P1_U2984) );
  INV_X1 U17624 ( .A(n14432), .ZN(n14433) );
  AOI21_X1 U17625 ( .B1(n10122), .B2(n14434), .A(n14433), .ZN(n14622) );
  AND2_X1 U17626 ( .A1(n14435), .A2(n14436), .ZN(n14621) );
  NAND2_X1 U17627 ( .A1(n14622), .A2(n14621), .ZN(n14620) );
  NAND2_X1 U17628 ( .A1(n14620), .A2(n14436), .ZN(n14438) );
  XNOR2_X1 U17629 ( .A(n14438), .B(n14437), .ZN(n15994) );
  AOI22_X1 U17630 ( .A1(n20111), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n20123), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14439) );
  OAI21_X1 U17631 ( .B1(n20122), .B2(n14440), .A(n14439), .ZN(n14441) );
  AOI21_X1 U17632 ( .B1(n14442), .B2(n20117), .A(n14441), .ZN(n14443) );
  OAI21_X1 U17633 ( .B1(n15994), .B2(n19955), .A(n14443), .ZN(P1_U2986) );
  MUX2_X1 U17634 ( .A(n14444), .B(n15936), .S(n15937), .Z(n14445) );
  XOR2_X1 U17635 ( .A(n12514), .B(n14445), .Z(n16010) );
  NAND2_X1 U17636 ( .A1(n16010), .A2(n20118), .ZN(n14449) );
  NOR2_X1 U17637 ( .A1(n19990), .A2(n20805), .ZN(n16008) );
  NOR2_X1 U17638 ( .A1(n20122), .A2(n14446), .ZN(n14447) );
  AOI211_X1 U17639 ( .C1(n20111), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16008), .B(n14447), .ZN(n14448) );
  OAI211_X1 U17640 ( .C1(n20161), .C2(n14450), .A(n14449), .B(n14448), .ZN(
        P1_U2989) );
  OR2_X1 U17641 ( .A1(n20141), .A2(n16017), .ZN(n14461) );
  INV_X1 U17642 ( .A(n14461), .ZN(n14452) );
  NOR2_X1 U17643 ( .A1(n14452), .A2(n10115), .ZN(n14471) );
  AND2_X1 U17644 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14511) );
  NAND2_X1 U17645 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16007) );
  NOR3_X1 U17646 ( .A1(n14454), .A2(n14453), .A3(n16007), .ZN(n14615) );
  NAND3_X1 U17647 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n14615), .ZN(n14562) );
  NOR2_X1 U17648 ( .A1(n15999), .A2(n14562), .ZN(n14605) );
  INV_X1 U17649 ( .A(n16007), .ZN(n14456) );
  NAND3_X1 U17650 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14456), .A3(
        n14455), .ZN(n14626) );
  NOR2_X1 U17651 ( .A1(n15984), .A2(n14626), .ZN(n14558) );
  NAND2_X1 U17652 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14558), .ZN(
        n14464) );
  NAND2_X1 U17653 ( .A1(n14618), .A2(n14464), .ZN(n14457) );
  NAND4_X1 U17654 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14603) );
  NOR2_X1 U17655 ( .A1(n14603), .A2(n14609), .ZN(n14563) );
  INV_X1 U17656 ( .A(n14563), .ZN(n14458) );
  NAND2_X1 U17657 ( .A1(n16017), .A2(n14458), .ZN(n14459) );
  OAI211_X1 U17658 ( .C1(n14616), .C2(n14605), .A(n14604), .B(n14459), .ZN(
        n14598) );
  OR2_X1 U17659 ( .A1(n14598), .A2(n14564), .ZN(n14460) );
  NAND2_X1 U17660 ( .A1(n14460), .A2(n14461), .ZN(n14577) );
  NAND2_X1 U17661 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14554) );
  NAND2_X1 U17662 ( .A1(n14461), .A2(n14554), .ZN(n14462) );
  AND2_X1 U17663 ( .A1(n14577), .A2(n14462), .ZN(n14533) );
  NAND2_X1 U17664 ( .A1(n16017), .A2(n14530), .ZN(n14463) );
  OAI21_X1 U17665 ( .B1(n14511), .B2(n15969), .A(n14522), .ZN(n14500) );
  AOI21_X1 U17666 ( .B1(n10053), .B2(n16017), .A(n14500), .ZN(n14483) );
  OAI211_X1 U17667 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15969), .A(
        n14483), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14480) );
  NAND2_X1 U17668 ( .A1(n20140), .A2(n14605), .ZN(n14532) );
  OR2_X1 U17669 ( .A1(n20147), .A2(n14464), .ZN(n14465) );
  NAND2_X1 U17670 ( .A1(n14532), .A2(n14465), .ZN(n15970) );
  NOR2_X1 U17671 ( .A1(n14564), .A2(n14554), .ZN(n14466) );
  AND2_X1 U17672 ( .A1(n14563), .A2(n14466), .ZN(n14467) );
  NAND2_X1 U17673 ( .A1(n15970), .A2(n14467), .ZN(n14543) );
  NOR2_X1 U17674 ( .A1(n14543), .A2(n14530), .ZN(n14526) );
  AND2_X1 U17675 ( .A1(n14526), .A2(n14511), .ZN(n14506) );
  NAND2_X1 U17676 ( .A1(n14506), .A2(n14468), .ZN(n14484) );
  INV_X1 U17677 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14475) );
  NOR4_X1 U17678 ( .A1(n14484), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14476), .A4(n14475), .ZN(n14469) );
  AOI211_X1 U17679 ( .C1(n14471), .C2(n14480), .A(n14470), .B(n14469), .ZN(
        n14474) );
  NAND2_X1 U17680 ( .A1(n14472), .A2(n20133), .ZN(n14473) );
  OAI21_X1 U17681 ( .B1(n14484), .B2(n14476), .A(n14475), .ZN(n14479) );
  NAND2_X1 U17682 ( .A1(n14482), .A2(n20152), .ZN(n14489) );
  INV_X1 U17683 ( .A(n14483), .ZN(n14487) );
  NOR2_X1 U17684 ( .A1(n14484), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14485) );
  AOI211_X1 U17685 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n14487), .A(
        n14486), .B(n14485), .ZN(n14488) );
  OAI211_X1 U17686 ( .C1(n20149), .C2(n14490), .A(n14489), .B(n14488), .ZN(
        P1_U3002) );
  INV_X1 U17687 ( .A(n14491), .ZN(n14497) );
  INV_X1 U17688 ( .A(n14506), .ZN(n14495) );
  XNOR2_X1 U17689 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14494) );
  AOI21_X1 U17690 ( .B1(n14500), .B2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14492), .ZN(n14493) );
  OAI21_X1 U17691 ( .B1(n14495), .B2(n14494), .A(n14493), .ZN(n14496) );
  AOI21_X1 U17692 ( .B1(n14497), .B2(n20133), .A(n14496), .ZN(n14498) );
  OAI21_X1 U17693 ( .B1(n14499), .B2(n15986), .A(n14498), .ZN(P1_U3003) );
  INV_X1 U17694 ( .A(n14500), .ZN(n14502) );
  OAI21_X1 U17695 ( .B1(n14502), .B2(n10056), .A(n14501), .ZN(n14505) );
  NOR2_X1 U17696 ( .A1(n14503), .A2(n20149), .ZN(n14504) );
  AOI211_X1 U17697 ( .C1(n14506), .C2(n10056), .A(n14505), .B(n14504), .ZN(
        n14507) );
  OAI21_X1 U17698 ( .B1(n14508), .B2(n15986), .A(n14507), .ZN(P1_U3004) );
  INV_X1 U17699 ( .A(n14522), .ZN(n14510) );
  AOI21_X1 U17700 ( .B1(n14510), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n14509), .ZN(n14516) );
  INV_X1 U17701 ( .A(n14511), .ZN(n14514) );
  NAND2_X1 U17702 ( .A1(n14525), .A2(n14512), .ZN(n14513) );
  NAND3_X1 U17703 ( .A1(n14526), .A2(n14514), .A3(n14513), .ZN(n14515) );
  OAI211_X1 U17704 ( .C1(n14517), .C2(n20149), .A(n14516), .B(n14515), .ZN(
        n14518) );
  INV_X1 U17705 ( .A(n14518), .ZN(n14519) );
  OAI21_X1 U17706 ( .B1(n14520), .B2(n15986), .A(n14519), .ZN(P1_U3005) );
  OAI21_X1 U17707 ( .B1(n14522), .B2(n14525), .A(n14521), .ZN(n14523) );
  AOI21_X1 U17708 ( .B1(n14524), .B2(n20133), .A(n14523), .ZN(n14528) );
  NAND2_X1 U17709 ( .A1(n14526), .A2(n14525), .ZN(n14527) );
  OAI211_X1 U17710 ( .C1(n14529), .C2(n15986), .A(n14528), .B(n14527), .ZN(
        P1_U3006) );
  INV_X1 U17711 ( .A(n14530), .ZN(n14531) );
  AOI21_X1 U17712 ( .B1(n14532), .B2(n20147), .A(n14531), .ZN(n14536) );
  INV_X1 U17713 ( .A(n14533), .ZN(n14544) );
  INV_X1 U17714 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14549) );
  OAI21_X1 U17715 ( .B1(n14543), .B2(n14549), .A(n14534), .ZN(n14535) );
  OAI21_X1 U17716 ( .B1(n14536), .B2(n14544), .A(n14535), .ZN(n14537) );
  OAI211_X1 U17717 ( .C1(n14539), .C2(n20149), .A(n14538), .B(n14537), .ZN(
        n14540) );
  INV_X1 U17718 ( .A(n14540), .ZN(n14541) );
  OAI21_X1 U17719 ( .B1(n14542), .B2(n15986), .A(n14541), .ZN(P1_U3007) );
  INV_X1 U17720 ( .A(n14543), .ZN(n14550) );
  NAND2_X1 U17721 ( .A1(n14544), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14545) );
  OAI211_X1 U17722 ( .C1(n14547), .C2(n20149), .A(n14546), .B(n14545), .ZN(
        n14548) );
  AOI21_X1 U17723 ( .B1(n14550), .B2(n14549), .A(n14548), .ZN(n14551) );
  OAI21_X1 U17724 ( .B1(n14552), .B2(n15986), .A(n14551), .ZN(P1_U3008) );
  NAND2_X1 U17725 ( .A1(n14553), .A2(n20152), .ZN(n14572) );
  INV_X1 U17726 ( .A(n14577), .ZN(n14570) );
  INV_X1 U17727 ( .A(n14554), .ZN(n14566) );
  INV_X1 U17728 ( .A(n14555), .ZN(n14583) );
  INV_X1 U17729 ( .A(n14562), .ZN(n14556) );
  NAND3_X1 U17730 ( .A1(n14557), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n14556), .ZN(n14561) );
  INV_X1 U17731 ( .A(n14558), .ZN(n14559) );
  OR2_X1 U17732 ( .A1(n20147), .A2(n14559), .ZN(n14560) );
  AND2_X1 U17733 ( .A1(n14561), .A2(n14560), .ZN(n14584) );
  OAI21_X1 U17734 ( .B1(n14583), .B2(n14562), .A(n14584), .ZN(n15993) );
  NAND3_X1 U17735 ( .A1(n15993), .A2(n14563), .A3(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14594) );
  NOR2_X1 U17736 ( .A1(n14594), .A2(n14564), .ZN(n14575) );
  INV_X1 U17737 ( .A(n14575), .ZN(n14565) );
  AOI211_X1 U17738 ( .C1(n10039), .C2(n14567), .A(n14566), .B(n14565), .ZN(
        n14568) );
  AOI211_X1 U17739 ( .C1(n14570), .C2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n14569), .B(n14568), .ZN(n14571) );
  OAI211_X1 U17740 ( .C1(n20149), .C2(n14573), .A(n14572), .B(n14571), .ZN(
        P1_U3009) );
  AOI21_X1 U17741 ( .B1(n14575), .B2(n10039), .A(n14574), .ZN(n14576) );
  OAI21_X1 U17742 ( .B1(n10039), .B2(n14577), .A(n14576), .ZN(n14578) );
  AOI21_X1 U17743 ( .B1(n14579), .B2(n20133), .A(n14578), .ZN(n14580) );
  OAI21_X1 U17744 ( .B1(n14581), .B2(n15986), .A(n14580), .ZN(P1_U3010) );
  INV_X1 U17745 ( .A(n14582), .ZN(n14592) );
  NAND2_X1 U17746 ( .A1(n10038), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14589) );
  AOI21_X1 U17747 ( .B1(n14584), .B2(n14583), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14585) );
  OAI21_X1 U17748 ( .B1(n14598), .B2(n14585), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14588) );
  INV_X1 U17749 ( .A(n14586), .ZN(n14587) );
  OAI211_X1 U17750 ( .C1(n14594), .C2(n14589), .A(n14588), .B(n14587), .ZN(
        n14590) );
  AOI21_X1 U17751 ( .B1(n15856), .B2(n20133), .A(n14590), .ZN(n14591) );
  OAI21_X1 U17752 ( .B1(n14592), .B2(n15986), .A(n14591), .ZN(P1_U3011) );
  OAI21_X1 U17753 ( .B1(n14594), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n14593), .ZN(n14597) );
  NOR2_X1 U17754 ( .A1(n14595), .A2(n20149), .ZN(n14596) );
  AOI211_X1 U17755 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n14598), .A(
        n14597), .B(n14596), .ZN(n14599) );
  OAI21_X1 U17756 ( .B1(n14600), .B2(n15986), .A(n14599), .ZN(P1_U3012) );
  NAND3_X1 U17757 ( .A1(n14602), .A2(n14601), .A3(n20152), .ZN(n14613) );
  INV_X1 U17758 ( .A(n14603), .ZN(n14610) );
  OAI21_X1 U17759 ( .B1(n14616), .B2(n14605), .A(n14604), .ZN(n14606) );
  INV_X1 U17760 ( .A(n14606), .ZN(n16000) );
  OAI21_X1 U17761 ( .B1(n14610), .B2(n15969), .A(n16000), .ZN(n15962) );
  NOR2_X1 U17762 ( .A1(n15864), .A2(n20149), .ZN(n14607) );
  AOI211_X1 U17763 ( .C1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n15962), .A(
        n14608), .B(n14607), .ZN(n14612) );
  NAND3_X1 U17764 ( .A1(n15970), .A2(n14610), .A3(n14609), .ZN(n14611) );
  NAND3_X1 U17765 ( .A1(n14613), .A2(n14612), .A3(n14611), .ZN(P1_U3013) );
  OAI21_X1 U17766 ( .B1(n14616), .B2(n14615), .A(n14614), .ZN(n14617) );
  AOI21_X1 U17767 ( .B1(n14618), .B2(n14626), .A(n14617), .ZN(n16006) );
  OAI21_X1 U17768 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n14619), .A(
        n16006), .ZN(n14628) );
  OAI21_X1 U17769 ( .B1(n14622), .B2(n14621), .A(n14620), .ZN(n14623) );
  INV_X1 U17770 ( .A(n14623), .ZN(n15935) );
  NAND2_X1 U17771 ( .A1(n15984), .A2(n14624), .ZN(n14625) );
  OAI22_X1 U17772 ( .A1(n15935), .A2(n15986), .B1(n14626), .B2(n14625), .ZN(
        n14627) );
  AOI21_X1 U17773 ( .B1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n14628), .A(
        n14627), .ZN(n14630) );
  NAND2_X1 U17774 ( .A1(n20123), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n14629) );
  OAI211_X1 U17775 ( .C1(n20149), .C2(n15882), .A(n14630), .B(n14629), .ZN(
        P1_U3019) );
  OR3_X1 U17776 ( .A1(n15969), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n14631), .ZN(n14640) );
  NAND3_X1 U17777 ( .A1(n14632), .A2(n13057), .A3(n20152), .ZN(n14639) );
  INV_X1 U17778 ( .A(n14633), .ZN(n14637) );
  NOR2_X1 U17779 ( .A1(n20973), .A2(n14634), .ZN(n14635) );
  AOI211_X1 U17780 ( .C1(n20133), .C2(n14637), .A(n14636), .B(n14635), .ZN(
        n14638) );
  NAND3_X1 U17781 ( .A1(n14640), .A2(n14639), .A3(n14638), .ZN(P1_U3030) );
  NAND3_X1 U17782 ( .A1(n14642), .A2(n16047), .A3(n14641), .ZN(n15818) );
  NAND2_X1 U17783 ( .A1(n20284), .A2(n14643), .ZN(n14644) );
  OAI211_X1 U17784 ( .C1(n20711), .C2(n12437), .A(n15818), .B(n14644), .ZN(
        n14645) );
  MUX2_X1 U17785 ( .A(n14645), .B(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .S(
        n20158), .Z(P1_U3478) );
  NOR2_X1 U17786 ( .A1(n11044), .A2(n14646), .ZN(n14648) );
  INV_X1 U17787 ( .A(n14648), .ZN(n14652) );
  AOI22_X1 U17788 ( .A1(n15787), .A2(n11027), .B1(n14648), .B2(n9743), .ZN(
        n14649) );
  OAI21_X1 U17789 ( .B1(n9741), .B2(n14650), .A(n14649), .ZN(n15791) );
  NOR2_X1 U17790 ( .A1(n20772), .A2(n20143), .ZN(n14656) );
  OAI22_X1 U17791 ( .A1(n10115), .A2(n20973), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14654) );
  AOI22_X1 U17792 ( .A1(n15791), .A2(n14657), .B1(n14656), .B2(n14654), .ZN(
        n14651) );
  OAI21_X1 U17793 ( .B1(n14661), .B2(n14652), .A(n14651), .ZN(n14653) );
  MUX2_X1 U17794 ( .A(n14653), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n14662), .Z(P1_U3473) );
  INV_X1 U17795 ( .A(n14654), .ZN(n14655) );
  AOI22_X1 U17796 ( .A1(n14658), .A2(n14657), .B1(n14656), .B2(n14655), .ZN(
        n14659) );
  OAI21_X1 U17797 ( .B1(n14661), .B2(n14660), .A(n14659), .ZN(n14663) );
  MUX2_X1 U17798 ( .A(n14663), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n14662), .Z(P1_U3472) );
  AOI21_X1 U17799 ( .B1(n14666), .B2(n14665), .A(n14664), .ZN(n14667) );
  NAND2_X1 U17800 ( .A1(n14667), .A2(n19021), .ZN(n14674) );
  OAI22_X1 U17801 ( .A1(n19010), .A2(n19882), .B1(n19037), .B2(n14668), .ZN(
        n14669) );
  AOI21_X1 U17802 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n19026), .A(n14669), .ZN(
        n14670) );
  OAI21_X1 U17803 ( .B1(n14822), .B2(n19029), .A(n14670), .ZN(n14671) );
  AOI21_X1 U17804 ( .B1(n14672), .B2(n19032), .A(n14671), .ZN(n14673) );
  OAI211_X1 U17805 ( .C1(n19034), .C2(n14723), .A(n14674), .B(n14673), .ZN(
        P2_U2827) );
  AOI211_X1 U17806 ( .C1(n14930), .C2(n14676), .A(n14675), .B(n19820), .ZN(
        n14677) );
  INV_X1 U17807 ( .A(n14677), .ZN(n14688) );
  NAND2_X1 U17808 ( .A1(n14756), .A2(n14678), .ZN(n14679) );
  NAND2_X1 U17809 ( .A1(n14738), .A2(n14679), .ZN(n15113) );
  INV_X1 U17810 ( .A(n15113), .ZN(n14686) );
  INV_X1 U17811 ( .A(n14854), .ZN(n14682) );
  INV_X1 U17812 ( .A(n14680), .ZN(n14681) );
  OAI21_X1 U17813 ( .B1(n14682), .B2(n14681), .A(n14837), .ZN(n15112) );
  AOI22_X1 U17814 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n18996), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19025), .ZN(n14684) );
  NAND2_X1 U17815 ( .A1(n19026), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n14683) );
  OAI211_X1 U17816 ( .C1(n15112), .C2(n19029), .A(n14684), .B(n14683), .ZN(
        n14685) );
  AOI21_X1 U17817 ( .B1(n14686), .B2(n19020), .A(n14685), .ZN(n14687) );
  OAI211_X1 U17818 ( .C1(n19018), .C2(n14689), .A(n14688), .B(n14687), .ZN(
        P2_U2830) );
  INV_X1 U17819 ( .A(n14973), .ZN(n14692) );
  INV_X1 U17820 ( .A(n14690), .ZN(n14691) );
  OAI221_X1 U17821 ( .B1(n14692), .B2(n14691), .C1(n14973), .C2(n14690), .A(
        n19021), .ZN(n14703) );
  OR2_X1 U17822 ( .A1(n14790), .A2(n14693), .ZN(n14694) );
  NAND2_X1 U17823 ( .A1(n9807), .A2(n14694), .ZN(n15183) );
  INV_X1 U17824 ( .A(n15183), .ZN(n14701) );
  INV_X1 U17825 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14695) );
  OAI22_X1 U17826 ( .A1(n14695), .A2(n19037), .B1(n14972), .B2(n19010), .ZN(
        n14700) );
  NOR2_X1 U17827 ( .A1(n14871), .A2(n14696), .ZN(n14697) );
  NOR2_X1 U17828 ( .A1(n12569), .A2(n14697), .ZN(n16127) );
  INV_X1 U17829 ( .A(n16127), .ZN(n14698) );
  OAI22_X1 U17830 ( .A1(n14698), .A2(n19029), .B1(n10930), .B2(n19012), .ZN(
        n14699) );
  AOI211_X1 U17831 ( .C1(n14701), .C2(n19020), .A(n14700), .B(n14699), .ZN(
        n14702) );
  OAI211_X1 U17832 ( .C1(n14704), .C2(n19018), .A(n14703), .B(n14702), .ZN(
        P2_U2835) );
  NOR2_X1 U17833 ( .A1(n9753), .A2(n14705), .ZN(n18939) );
  AOI21_X1 U17834 ( .B1(n16167), .B2(n14706), .A(n19820), .ZN(n14707) );
  AOI22_X1 U17835 ( .A1(n16167), .A2(n18931), .B1(n18939), .B2(n14707), .ZN(
        n14716) );
  INV_X1 U17836 ( .A(n18983), .ZN(n19000) );
  OAI22_X1 U17837 ( .A1(n16174), .A2(n19037), .B1(n12187), .B2(n19010), .ZN(
        n14708) );
  AOI211_X1 U17838 ( .C1(P2_EBX_REG_11__SCAN_IN), .C2(n19026), .A(n19000), .B(
        n14708), .ZN(n14715) );
  INV_X1 U17839 ( .A(n14709), .ZN(n14711) );
  AOI211_X1 U17840 ( .C1(P2_EBX_REG_11__SCAN_IN), .C2(n14711), .A(n19018), .B(
        n14710), .ZN(n14713) );
  OAI22_X1 U17841 ( .A1(n15314), .A2(n19034), .B1(n19029), .B2(n15313), .ZN(
        n14712) );
  NOR2_X1 U17842 ( .A1(n14713), .A2(n14712), .ZN(n14714) );
  NAND3_X1 U17843 ( .A1(n14716), .A2(n14715), .A3(n14714), .ZN(P2_U2844) );
  NAND2_X1 U17844 ( .A1(n16057), .A2(n14808), .ZN(n14717) );
  OAI21_X1 U17845 ( .B1(n14808), .B2(n14718), .A(n14717), .ZN(P2_U2856) );
  NOR2_X1 U17846 ( .A1(n14719), .A2(n14720), .ZN(n14722) );
  XNOR2_X1 U17847 ( .A(n14722), .B(n14721), .ZN(n14827) );
  NOR2_X1 U17848 ( .A1(n14723), .A2(n14791), .ZN(n14724) );
  AOI21_X1 U17849 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n14791), .A(n14724), .ZN(
        n14725) );
  OAI21_X1 U17850 ( .B1(n14827), .B2(n14811), .A(n14725), .ZN(P2_U2859) );
  OAI21_X1 U17851 ( .B1(n9799), .B2(n14727), .A(n14726), .ZN(n14835) );
  OR2_X1 U17852 ( .A1(n14740), .A2(n14728), .ZN(n14729) );
  NAND2_X1 U17853 ( .A1(n14730), .A2(n14729), .ZN(n16085) );
  NOR2_X1 U17854 ( .A1(n16085), .A2(n14791), .ZN(n14731) );
  AOI21_X1 U17855 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n14791), .A(n14731), .ZN(
        n14732) );
  OAI21_X1 U17856 ( .B1(n14835), .B2(n14811), .A(n14732), .ZN(P2_U2860) );
  OAI21_X1 U17857 ( .B1(n14734), .B2(n14736), .A(n14735), .ZN(n14845) );
  NAND2_X1 U17858 ( .A1(n14804), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14742) );
  AND2_X1 U17859 ( .A1(n14738), .A2(n14737), .ZN(n14739) );
  NOR2_X1 U17860 ( .A1(n14740), .A2(n14739), .ZN(n16093) );
  NAND2_X1 U17861 ( .A1(n16093), .A2(n14808), .ZN(n14741) );
  OAI211_X1 U17862 ( .C1(n14845), .C2(n14811), .A(n14742), .B(n14741), .ZN(
        P2_U2861) );
  OAI21_X1 U17863 ( .B1(n14744), .B2(n14746), .A(n14745), .ZN(n14850) );
  MUX2_X1 U17864 ( .A(n15113), .B(n14747), .S(n14791), .Z(n14748) );
  OAI21_X1 U17865 ( .B1(n14850), .B2(n14811), .A(n14748), .ZN(P2_U2862) );
  AOI21_X1 U17866 ( .B1(n14749), .B2(n14750), .A(n9790), .ZN(n14751) );
  XOR2_X1 U17867 ( .A(n14752), .B(n14751), .Z(n14860) );
  NAND2_X1 U17868 ( .A1(n14754), .A2(n14753), .ZN(n14755) );
  NAND2_X1 U17869 ( .A1(n14756), .A2(n14755), .ZN(n16110) );
  NOR2_X1 U17870 ( .A1(n16110), .A2(n14791), .ZN(n14757) );
  AOI21_X1 U17871 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n14791), .A(n14757), .ZN(
        n14758) );
  OAI21_X1 U17872 ( .B1(n14860), .B2(n14811), .A(n14758), .ZN(P2_U2863) );
  AOI21_X1 U17873 ( .B1(n14759), .B2(n14762), .A(n14761), .ZN(n14763) );
  INV_X1 U17874 ( .A(n14763), .ZN(n14865) );
  NOR2_X1 U17875 ( .A1(n14808), .A2(n10984), .ZN(n14764) );
  AOI21_X1 U17876 ( .B1(n16142), .B2(n14808), .A(n14764), .ZN(n14765) );
  OAI21_X1 U17877 ( .B1(n14865), .B2(n14811), .A(n14765), .ZN(P2_U2864) );
  AND2_X1 U17878 ( .A1(n9778), .A2(n14766), .ZN(n14768) );
  OR2_X1 U17879 ( .A1(n14768), .A2(n14767), .ZN(n16148) );
  INV_X1 U17880 ( .A(n14770), .ZN(n14771) );
  AOI21_X1 U17881 ( .B1(n14773), .B2(n14771), .A(n14772), .ZN(n16123) );
  NAND2_X1 U17882 ( .A1(n16123), .A2(n14783), .ZN(n14775) );
  NAND2_X1 U17883 ( .A1(n14804), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n14774) );
  OAI211_X1 U17884 ( .C1(n16148), .C2(n14804), .A(n14775), .B(n14774), .ZN(
        P2_U2865) );
  AOI21_X1 U17885 ( .B1(n14777), .B2(n14776), .A(n14770), .ZN(n14869) );
  NAND2_X1 U17886 ( .A1(n14869), .A2(n14783), .ZN(n14779) );
  NAND2_X1 U17887 ( .A1(n14804), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n14778) );
  OAI211_X1 U17888 ( .C1(n15163), .C2(n14804), .A(n14779), .B(n14778), .ZN(
        P2_U2866) );
  OR2_X1 U17889 ( .A1(n14780), .A2(n14781), .ZN(n14782) );
  AND2_X1 U17890 ( .A1(n14782), .A2(n14776), .ZN(n16128) );
  NAND2_X1 U17891 ( .A1(n16128), .A2(n14783), .ZN(n14785) );
  NAND2_X1 U17892 ( .A1(n14804), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n14784) );
  OAI211_X1 U17893 ( .C1(n15183), .C2(n14804), .A(n14785), .B(n14784), .ZN(
        P2_U2867) );
  AOI21_X1 U17894 ( .B1(n14786), .B2(n9768), .A(n14780), .ZN(n14787) );
  INV_X1 U17895 ( .A(n14787), .ZN(n14879) );
  NOR2_X1 U17896 ( .A1(n14799), .A2(n14788), .ZN(n14789) );
  OR2_X1 U17897 ( .A1(n14790), .A2(n14789), .ZN(n15190) );
  NOR2_X1 U17898 ( .A1(n15190), .A2(n14791), .ZN(n14792) );
  AOI21_X1 U17899 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n14791), .A(n14792), .ZN(
        n14793) );
  OAI21_X1 U17900 ( .B1(n14879), .B2(n14811), .A(n14793), .ZN(P2_U2868) );
  NAND2_X1 U17901 ( .A1(n14794), .A2(n14795), .ZN(n14796) );
  NAND2_X1 U17902 ( .A1(n9768), .A2(n14796), .ZN(n16134) );
  AND2_X1 U17903 ( .A1(n14805), .A2(n14797), .ZN(n14798) );
  NOR2_X1 U17904 ( .A1(n14799), .A2(n14798), .ZN(n18897) );
  NOR2_X1 U17905 ( .A1(n14808), .A2(n14800), .ZN(n14801) );
  AOI21_X1 U17906 ( .B1(n18897), .B2(n14808), .A(n14801), .ZN(n14802) );
  OAI21_X1 U17907 ( .B1(n16134), .B2(n14811), .A(n14802), .ZN(P2_U2869) );
  OAI21_X1 U17908 ( .B1(n14803), .B2(n10267), .A(n14794), .ZN(n14886) );
  NAND2_X1 U17909 ( .A1(n14804), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n14810) );
  AOI21_X1 U17910 ( .B1(n14807), .B2(n14806), .A(n10794), .ZN(n18907) );
  NAND2_X1 U17911 ( .A1(n18907), .A2(n14808), .ZN(n14809) );
  OAI211_X1 U17912 ( .C1(n14886), .C2(n14811), .A(n14810), .B(n14809), .ZN(
        P2_U2870) );
  NAND3_X1 U17913 ( .A1(n14812), .A2(n13871), .A3(n19064), .ZN(n14820) );
  OAI21_X1 U17914 ( .B1(n14815), .B2(n14814), .A(n14813), .ZN(n16074) );
  INV_X1 U17915 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n19083) );
  OAI22_X1 U17916 ( .A1(n16074), .A2(n16132), .B1(n19060), .B2(n19083), .ZN(
        n14816) );
  AOI21_X1 U17917 ( .B1(n14883), .B2(n14817), .A(n14816), .ZN(n14819) );
  AOI22_X1 U17918 ( .A1(n19044), .A2(BUF1_REG_29__SCAN_IN), .B1(n19046), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n14818) );
  NAND3_X1 U17919 ( .A1(n14820), .A2(n14819), .A3(n14818), .ZN(P2_U2890) );
  INV_X1 U17920 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n14821) );
  OAI22_X1 U17921 ( .A1(n14822), .A2(n16132), .B1(n19060), .B2(n14821), .ZN(
        n14824) );
  INV_X1 U17922 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n19230) );
  OAI22_X1 U17923 ( .A1(n19051), .A2(n19230), .B1(n19059), .B2(n19231), .ZN(
        n14823) );
  AOI211_X1 U17924 ( .C1(n14883), .C2(n14825), .A(n14824), .B(n14823), .ZN(
        n14826) );
  OAI21_X1 U17925 ( .B1(n14827), .B2(n16133), .A(n14826), .ZN(P2_U2891) );
  AOI21_X1 U17926 ( .B1(n14829), .B2(n14839), .A(n14828), .ZN(n14830) );
  INV_X1 U17927 ( .A(n14830), .ZN(n16089) );
  OAI22_X1 U17928 ( .A1(n16089), .A2(n16132), .B1(n19060), .B2(n19086), .ZN(
        n14831) );
  AOI21_X1 U17929 ( .B1(n14883), .B2(n14832), .A(n14831), .ZN(n14834) );
  AOI22_X1 U17930 ( .A1(n19044), .A2(BUF1_REG_27__SCAN_IN), .B1(n19046), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n14833) );
  OAI211_X1 U17931 ( .C1(n14835), .C2(n16133), .A(n14834), .B(n14833), .ZN(
        P2_U2892) );
  NAND2_X1 U17932 ( .A1(n14837), .A2(n14836), .ZN(n14838) );
  AND2_X1 U17933 ( .A1(n14839), .A2(n14838), .ZN(n16104) );
  INV_X1 U17934 ( .A(n16104), .ZN(n14840) );
  OAI22_X1 U17935 ( .A1(n14840), .A2(n16132), .B1(n19060), .B2(n20996), .ZN(
        n14841) );
  AOI21_X1 U17936 ( .B1(n14883), .B2(n14842), .A(n14841), .ZN(n14844) );
  AOI22_X1 U17937 ( .A1(n19044), .A2(BUF1_REG_26__SCAN_IN), .B1(n19046), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n14843) );
  OAI211_X1 U17938 ( .C1(n14845), .C2(n16133), .A(n14844), .B(n14843), .ZN(
        P2_U2893) );
  OAI22_X1 U17939 ( .A1(n15112), .A2(n16132), .B1(n19060), .B2(n19089), .ZN(
        n14846) );
  AOI21_X1 U17940 ( .B1(n14883), .B2(n14847), .A(n14846), .ZN(n14849) );
  AOI22_X1 U17941 ( .A1(n19044), .A2(BUF1_REG_25__SCAN_IN), .B1(n19046), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n14848) );
  OAI211_X1 U17942 ( .C1(n14850), .C2(n16133), .A(n14849), .B(n14848), .ZN(
        P2_U2894) );
  OR2_X1 U17943 ( .A1(n14852), .A2(n14851), .ZN(n14853) );
  NAND2_X1 U17944 ( .A1(n14854), .A2(n14853), .ZN(n16109) );
  INV_X1 U17945 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n14855) );
  OAI22_X1 U17946 ( .A1(n16109), .A2(n16132), .B1(n19060), .B2(n14855), .ZN(
        n14857) );
  INV_X1 U17947 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n19206) );
  OAI22_X1 U17948 ( .A1(n19051), .A2(n19206), .B1(n19059), .B2(n19207), .ZN(
        n14856) );
  AOI211_X1 U17949 ( .C1(n14883), .C2(n14858), .A(n14857), .B(n14856), .ZN(
        n14859) );
  OAI21_X1 U17950 ( .B1(n14860), .B2(n16133), .A(n14859), .ZN(P2_U2895) );
  INV_X1 U17951 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n19092) );
  OAI22_X1 U17952 ( .A1(n15135), .A2(n16132), .B1(n19060), .B2(n19092), .ZN(
        n14861) );
  AOI21_X1 U17953 ( .B1(n14883), .B2(n14862), .A(n14861), .ZN(n14864) );
  AOI22_X1 U17954 ( .A1(n19044), .A2(BUF1_REG_23__SCAN_IN), .B1(n19046), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n14863) );
  OAI211_X1 U17955 ( .C1(n14865), .C2(n16133), .A(n14864), .B(n14863), .ZN(
        P2_U2896) );
  INV_X1 U17956 ( .A(n14883), .ZN(n19049) );
  AOI22_X1 U17957 ( .A1(n19044), .A2(BUF1_REG_21__SCAN_IN), .B1(n19046), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n14867) );
  AOI22_X1 U17958 ( .A1(n15166), .A2(n19055), .B1(P2_EAX_REG_21__SCAN_IN), 
        .B2(n19053), .ZN(n14866) );
  OAI211_X1 U17959 ( .C1(n19237), .C2(n19049), .A(n14867), .B(n14866), .ZN(
        n14868) );
  AOI21_X1 U17960 ( .B1(n14869), .B2(n19064), .A(n14868), .ZN(n14870) );
  INV_X1 U17961 ( .A(n14870), .ZN(P2_U2898) );
  INV_X1 U17962 ( .A(n14871), .ZN(n14872) );
  OAI21_X1 U17963 ( .B1(n15203), .B2(n14873), .A(n14872), .ZN(n18888) );
  INV_X1 U17964 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14874) );
  OAI22_X1 U17965 ( .A1(n18888), .A2(n16132), .B1(n19060), .B2(n14874), .ZN(
        n14875) );
  AOI21_X1 U17966 ( .B1(n14883), .B2(n14876), .A(n14875), .ZN(n14878) );
  AOI22_X1 U17967 ( .A1(n19044), .A2(BUF1_REG_19__SCAN_IN), .B1(n19046), .B2(
        BUF2_REG_19__SCAN_IN), .ZN(n14877) );
  OAI211_X1 U17968 ( .C1(n14879), .C2(n16133), .A(n14878), .B(n14877), .ZN(
        P2_U2900) );
  OAI21_X1 U17969 ( .B1(n12246), .B2(n14880), .A(n15202), .ZN(n18911) );
  INV_X1 U17970 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n19103) );
  OAI22_X1 U17971 ( .A1(n18911), .A2(n16132), .B1(n19060), .B2(n19103), .ZN(
        n14881) );
  AOI21_X1 U17972 ( .B1(n14883), .B2(n14882), .A(n14881), .ZN(n14885) );
  AOI22_X1 U17973 ( .A1(n19044), .A2(BUF1_REG_17__SCAN_IN), .B1(n19046), .B2(
        BUF2_REG_17__SCAN_IN), .ZN(n14884) );
  OAI211_X1 U17974 ( .C1(n14886), .C2(n16133), .A(n14885), .B(n14884), .ZN(
        P2_U2902) );
  XNOR2_X1 U17975 ( .A(n9780), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15073) );
  NAND2_X1 U17976 ( .A1(n10151), .A2(n14888), .ZN(n14889) );
  XNOR2_X1 U17977 ( .A(n14890), .B(n14889), .ZN(n15063) );
  NAND2_X1 U17978 ( .A1(n15063), .A2(n19162), .ZN(n14895) );
  INV_X1 U17979 ( .A(n14891), .ZN(n15070) );
  NAND2_X1 U17980 ( .A1(n19000), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15066) );
  NAND2_X1 U17981 ( .A1(n19154), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14892) );
  OAI211_X1 U17982 ( .C1(n19152), .C2(n16058), .A(n15066), .B(n14892), .ZN(
        n14893) );
  AOI21_X1 U17983 ( .B1(n15070), .B2(n19156), .A(n14893), .ZN(n14894) );
  OAI211_X1 U17984 ( .C1(n15073), .C2(n19159), .A(n14895), .B(n14894), .ZN(
        P2_U2984) );
  NAND2_X1 U17985 ( .A1(n14897), .A2(n14896), .ZN(n14898) );
  XOR2_X1 U17986 ( .A(n14899), .B(n14898), .Z(n15086) );
  AOI21_X1 U17987 ( .B1(n15076), .B2(n14900), .A(n9780), .ZN(n15084) );
  NOR2_X1 U17988 ( .A1(n16226), .A2(n19884), .ZN(n15079) );
  AOI21_X1 U17989 ( .B1(n19154), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15079), .ZN(n14902) );
  NAND2_X1 U17990 ( .A1(n16217), .A2(n16064), .ZN(n14901) );
  OAI211_X1 U17991 ( .C1(n16070), .C2(n16211), .A(n14902), .B(n14901), .ZN(
        n14903) );
  AOI21_X1 U17992 ( .B1(n15084), .B2(n16186), .A(n14903), .ZN(n14904) );
  OAI21_X1 U17993 ( .B1(n15086), .B2(n16219), .A(n14904), .ZN(P2_U2985) );
  INV_X1 U17994 ( .A(n14905), .ZN(n14906) );
  OAI21_X1 U17995 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14919), .A(
        n14906), .ZN(n15097) );
  NAND3_X1 U17996 ( .A1(n14907), .A2(n19162), .A3(n15087), .ZN(n14912) );
  INV_X1 U17997 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19881) );
  OR2_X1 U17998 ( .A1(n18983), .A2(n19881), .ZN(n15091) );
  OAI21_X1 U17999 ( .B1(n16225), .B2(n16078), .A(n15091), .ZN(n14910) );
  NOR2_X1 U18000 ( .A1(n16085), .A2(n16211), .ZN(n14909) );
  AOI211_X1 U18001 ( .C1(n16217), .C2(n16076), .A(n14910), .B(n14909), .ZN(
        n14911) );
  OAI211_X1 U18002 ( .C1(n19159), .C2(n15097), .A(n14912), .B(n14911), .ZN(
        P2_U2987) );
  NAND2_X1 U18003 ( .A1(n14913), .A2(n14923), .ZN(n14914) );
  XOR2_X1 U18004 ( .A(n14915), .B(n14914), .Z(n15109) );
  NAND2_X1 U18005 ( .A1(n16243), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15098) );
  NAND2_X1 U18006 ( .A1(n19154), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14916) );
  OAI211_X1 U18007 ( .C1(n19152), .C2(n14917), .A(n15098), .B(n14916), .ZN(
        n14921) );
  NOR2_X1 U18008 ( .A1(n9788), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14918) );
  OR2_X1 U18009 ( .A1(n14919), .A2(n14918), .ZN(n15105) );
  NOR2_X1 U18010 ( .A1(n15105), .A2(n19159), .ZN(n14920) );
  AOI211_X1 U18011 ( .C1(n19156), .C2(n16093), .A(n14921), .B(n14920), .ZN(
        n14922) );
  OAI21_X1 U18012 ( .B1(n15109), .B2(n16219), .A(n14922), .ZN(P2_U2988) );
  NAND2_X1 U18013 ( .A1(n14924), .A2(n14923), .ZN(n14926) );
  XOR2_X1 U18014 ( .A(n14926), .B(n14925), .Z(n15121) );
  INV_X1 U18015 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n21077) );
  OAI22_X1 U18016 ( .A1(n16225), .A2(n14927), .B1(n21077), .B2(n18983), .ZN(
        n14929) );
  NOR2_X1 U18017 ( .A1(n15113), .A2(n16211), .ZN(n14928) );
  AOI211_X1 U18018 ( .C1(n16217), .C2(n14930), .A(n14929), .B(n14928), .ZN(
        n14932) );
  INV_X1 U18019 ( .A(n9788), .ZN(n15118) );
  NAND2_X1 U18020 ( .A1(n14936), .A2(n21137), .ZN(n15117) );
  NAND3_X1 U18021 ( .A1(n15118), .A2(n16186), .A3(n15117), .ZN(n14931) );
  OAI211_X1 U18022 ( .C1(n15121), .C2(n16219), .A(n14932), .B(n14931), .ZN(
        P2_U2989) );
  XNOR2_X1 U18023 ( .A(n14933), .B(n15124), .ZN(n14934) );
  XNOR2_X1 U18024 ( .A(n14935), .B(n14934), .ZN(n15130) );
  INV_X1 U18025 ( .A(n14936), .ZN(n14937) );
  AOI21_X1 U18026 ( .B1(n15124), .B2(n15142), .A(n14937), .ZN(n15128) );
  NOR2_X1 U18027 ( .A1(n16110), .A2(n16211), .ZN(n14941) );
  AOI22_X1 U18028 ( .A1(n19154), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19000), .ZN(n14938) );
  OAI21_X1 U18029 ( .B1(n19152), .B2(n14939), .A(n14938), .ZN(n14940) );
  AOI211_X1 U18030 ( .C1(n15128), .C2(n16186), .A(n14941), .B(n14940), .ZN(
        n14942) );
  OAI21_X1 U18031 ( .B1(n15130), .B2(n16219), .A(n14942), .ZN(P2_U2990) );
  NAND2_X1 U18032 ( .A1(n14943), .A2(n15276), .ZN(n15029) );
  INV_X1 U18033 ( .A(n15026), .ZN(n14944) );
  AOI21_X1 U18034 ( .B1(n15029), .B2(n15027), .A(n14944), .ZN(n15018) );
  INV_X1 U18035 ( .A(n15016), .ZN(n14945) );
  INV_X1 U18036 ( .A(n14946), .ZN(n14947) );
  INV_X1 U18037 ( .A(n14948), .ZN(n14949) );
  AND2_X1 U18038 ( .A1(n14949), .A2(n14950), .ZN(n15000) );
  INV_X1 U18039 ( .A(n14950), .ZN(n14951) );
  INV_X1 U18040 ( .A(n14952), .ZN(n14953) );
  OAI211_X1 U18041 ( .C1(n14991), .C2(n14953), .A(n14990), .B(n14979), .ZN(
        n14967) );
  NAND2_X1 U18042 ( .A1(n14967), .A2(n14968), .ZN(n14966) );
  NAND2_X1 U18043 ( .A1(n14966), .A2(n14970), .ZN(n14957) );
  NAND2_X1 U18044 ( .A1(n14955), .A2(n14954), .ZN(n14956) );
  XNOR2_X1 U18045 ( .A(n14957), .B(n14956), .ZN(n15174) );
  NAND2_X1 U18046 ( .A1(n15320), .A2(n15207), .ZN(n15002) );
  AOI21_X1 U18047 ( .B1(n14983), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14959) );
  INV_X1 U18048 ( .A(n15159), .ZN(n14958) );
  NOR2_X1 U18049 ( .A1(n14959), .A2(n14958), .ZN(n15172) );
  NOR2_X1 U18050 ( .A1(n16226), .A2(n19874), .ZN(n15165) );
  NOR2_X1 U18051 ( .A1(n16225), .A2(n14960), .ZN(n14961) );
  AOI211_X1 U18052 ( .C1(n14962), .C2(n16217), .A(n15165), .B(n14961), .ZN(
        n14963) );
  OAI21_X1 U18053 ( .B1(n15163), .B2(n16211), .A(n14963), .ZN(n14964) );
  AOI21_X1 U18054 ( .B1(n15172), .B2(n16186), .A(n14964), .ZN(n14965) );
  OAI21_X1 U18055 ( .B1(n15174), .B2(n16219), .A(n14965), .ZN(P2_U2993) );
  INV_X1 U18056 ( .A(n14966), .ZN(n14971) );
  AOI21_X1 U18057 ( .B1(n14970), .B2(n14968), .A(n14967), .ZN(n14969) );
  AOI21_X1 U18058 ( .B1(n14971), .B2(n14970), .A(n14969), .ZN(n15189) );
  XNOR2_X1 U18059 ( .A(n14983), .B(n15179), .ZN(n15186) );
  NOR2_X1 U18060 ( .A1(n16226), .A2(n14972), .ZN(n15178) );
  NOR2_X1 U18061 ( .A1(n19152), .A2(n14973), .ZN(n14974) );
  AOI211_X1 U18062 ( .C1(n19154), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15178), .B(n14974), .ZN(n14975) );
  OAI21_X1 U18063 ( .B1(n15183), .B2(n16211), .A(n14975), .ZN(n14976) );
  AOI21_X1 U18064 ( .B1(n15186), .B2(n16186), .A(n14976), .ZN(n14977) );
  OAI21_X1 U18065 ( .B1(n15189), .B2(n16219), .A(n14977), .ZN(P2_U2994) );
  INV_X1 U18066 ( .A(n14989), .ZN(n14978) );
  OAI21_X1 U18067 ( .B1(n14991), .B2(n14978), .A(n14990), .ZN(n14982) );
  NAND2_X1 U18068 ( .A1(n14980), .A2(n14979), .ZN(n14981) );
  XNOR2_X1 U18069 ( .A(n14982), .B(n14981), .ZN(n15200) );
  AOI21_X1 U18070 ( .B1(n15195), .B2(n14993), .A(n14983), .ZN(n15198) );
  NAND2_X1 U18071 ( .A1(n19000), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15191) );
  OAI21_X1 U18072 ( .B1(n16225), .B2(n14984), .A(n15191), .ZN(n14985) );
  AOI21_X1 U18073 ( .B1(n16217), .B2(n18881), .A(n14985), .ZN(n14986) );
  OAI21_X1 U18074 ( .B1(n15190), .B2(n16211), .A(n14986), .ZN(n14987) );
  AOI21_X1 U18075 ( .B1(n15198), .B2(n16186), .A(n14987), .ZN(n14988) );
  OAI21_X1 U18076 ( .B1(n15200), .B2(n16219), .A(n14988), .ZN(P2_U2995) );
  NAND2_X1 U18077 ( .A1(n14990), .A2(n14989), .ZN(n14992) );
  XOR2_X1 U18078 ( .A(n14992), .B(n14991), .Z(n15214) );
  INV_X1 U18079 ( .A(n14993), .ZN(n14994) );
  AOI21_X1 U18080 ( .B1(n20943), .B2(n15002), .A(n14994), .ZN(n15212) );
  NAND2_X1 U18081 ( .A1(n18897), .A2(n19156), .ZN(n14996) );
  NOR2_X1 U18082 ( .A1(n16226), .A2(n19869), .ZN(n15206) );
  AOI21_X1 U18083 ( .B1(n19154), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15206), .ZN(n14995) );
  OAI211_X1 U18084 ( .C1(n19152), .C2(n18890), .A(n14996), .B(n14995), .ZN(
        n14997) );
  AOI21_X1 U18085 ( .B1(n15212), .B2(n16186), .A(n14997), .ZN(n14998) );
  OAI21_X1 U18086 ( .B1(n15214), .B2(n16219), .A(n14998), .ZN(P2_U2996) );
  XOR2_X1 U18087 ( .A(n15000), .B(n14999), .Z(n15230) );
  NAND2_X1 U18088 ( .A1(n16217), .A2(n18905), .ZN(n15001) );
  NAND2_X1 U18089 ( .A1(n19000), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15215) );
  OAI211_X1 U18090 ( .C1(n16225), .C2(n9987), .A(n15001), .B(n15215), .ZN(
        n15006) );
  NOR2_X2 U18091 ( .A1(n15303), .A2(n15259), .ZN(n15273) );
  INV_X1 U18092 ( .A(n15002), .ZN(n15003) );
  AOI211_X1 U18093 ( .C1(n15221), .C2(n15004), .A(n15003), .B(n19159), .ZN(
        n15005) );
  AOI211_X1 U18094 ( .C1(n19156), .C2(n18907), .A(n15006), .B(n15005), .ZN(
        n15007) );
  OAI21_X1 U18095 ( .B1(n15230), .B2(n16219), .A(n15007), .ZN(P2_U2997) );
  XNOR2_X1 U18096 ( .A(n15009), .B(n15008), .ZN(n15243) );
  XOR2_X1 U18097 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n15217), .Z(
        n15010) );
  NAND2_X1 U18098 ( .A1(n15010), .A2(n16186), .ZN(n15014) );
  INV_X1 U18099 ( .A(n15236), .ZN(n18919) );
  NOR2_X1 U18100 ( .A1(n15235), .A2(n16226), .ZN(n15012) );
  OAI22_X1 U18101 ( .A1(n16225), .A2(n9986), .B1(n19152), .B2(n18913), .ZN(
        n15011) );
  AOI211_X1 U18102 ( .C1(n19156), .C2(n18919), .A(n15012), .B(n15011), .ZN(
        n15013) );
  OAI211_X1 U18103 ( .C1(n16219), .C2(n15243), .A(n15014), .B(n15013), .ZN(
        P2_U2998) );
  NAND2_X1 U18104 ( .A1(n15016), .A2(n15015), .ZN(n15017) );
  XNOR2_X1 U18105 ( .A(n15018), .B(n15017), .ZN(n15256) );
  AOI21_X1 U18106 ( .B1(n15252), .B2(n15025), .A(n15217), .ZN(n15244) );
  NAND2_X1 U18107 ( .A1(n15244), .A2(n16186), .ZN(n15024) );
  OAI22_X1 U18108 ( .A1(n16225), .A2(n15019), .B1(n21120), .B2(n16226), .ZN(
        n15021) );
  NOR2_X1 U18109 ( .A1(n15248), .A2(n16211), .ZN(n15020) );
  AOI211_X1 U18110 ( .C1(n16217), .C2(n15022), .A(n15021), .B(n15020), .ZN(
        n15023) );
  OAI211_X1 U18111 ( .C1(n15256), .C2(n16219), .A(n15024), .B(n15023), .ZN(
        P2_U2999) );
  OAI21_X1 U18112 ( .B1(n15273), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15025), .ZN(n15272) );
  NAND2_X1 U18113 ( .A1(n15027), .A2(n15026), .ZN(n15028) );
  XNOR2_X1 U18114 ( .A(n15029), .B(n15028), .ZN(n15270) );
  NOR2_X1 U18115 ( .A1(n18983), .A2(n19864), .ZN(n15263) );
  NOR2_X1 U18116 ( .A1(n19152), .A2(n15030), .ZN(n15031) );
  AOI211_X1 U18117 ( .C1(n19154), .C2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n15263), .B(n15031), .ZN(n15032) );
  OAI21_X1 U18118 ( .B1(n16211), .B2(n15262), .A(n15032), .ZN(n15033) );
  AOI21_X1 U18119 ( .B1(n15270), .B2(n19162), .A(n15033), .ZN(n15034) );
  OAI21_X1 U18120 ( .B1(n15272), .B2(n19159), .A(n15034), .ZN(P2_U3000) );
  AND2_X1 U18121 ( .A1(n15035), .A2(n15036), .ZN(n16197) );
  INV_X1 U18122 ( .A(n16197), .ZN(n15039) );
  INV_X1 U18123 ( .A(n15036), .ZN(n15037) );
  NOR2_X1 U18124 ( .A1(n15037), .A2(n16196), .ZN(n15038) );
  OAI22_X1 U18125 ( .A1(n15039), .A2(n16196), .B1(n15038), .B2(n15035), .ZN(
        n15344) );
  OR2_X1 U18126 ( .A1(n15040), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15336) );
  NAND3_X1 U18127 ( .A1(n15336), .A2(n15335), .A3(n16186), .ZN(n15046) );
  OAI22_X1 U18128 ( .A1(n16225), .A2(n15041), .B1(n19853), .B2(n18983), .ZN(
        n15044) );
  INV_X1 U18129 ( .A(n18972), .ZN(n15042) );
  NOR2_X1 U18130 ( .A1(n19152), .A2(n15042), .ZN(n15043) );
  AOI211_X1 U18131 ( .C1(n19156), .C2(n18976), .A(n15044), .B(n15043), .ZN(
        n15045) );
  OAI211_X1 U18132 ( .C1(n16219), .C2(n15344), .A(n15046), .B(n15045), .ZN(
        P2_U3007) );
  NAND2_X1 U18133 ( .A1(n15047), .A2(n19182), .ZN(n15061) );
  INV_X1 U18134 ( .A(n16057), .ZN(n15058) );
  INV_X1 U18135 ( .A(n19192), .ZN(n15050) );
  NOR2_X1 U18136 ( .A1(n15076), .A2(n15077), .ZN(n15075) );
  INV_X1 U18137 ( .A(n15075), .ZN(n15049) );
  AOI211_X1 U18138 ( .C1(n15050), .C2(n15049), .A(n15048), .B(n15094), .ZN(
        n15065) );
  AOI222_X1 U18139 ( .A1(n12095), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n12253), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C1(n12264), .C2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n15051) );
  INV_X1 U18140 ( .A(n15053), .ZN(n15055) );
  NAND4_X1 U18141 ( .A1(n15089), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15075), .A4(n10698), .ZN(n15054) );
  OAI211_X1 U18142 ( .C1(n16056), .C2(n16251), .A(n15055), .B(n15054), .ZN(
        n15056) );
  INV_X1 U18143 ( .A(n15056), .ZN(n15057) );
  INV_X1 U18144 ( .A(n15059), .ZN(n15060) );
  OAI211_X1 U18145 ( .C1(n15062), .C2(n19202), .A(n15061), .B(n15060), .ZN(
        P2_U3015) );
  NAND2_X1 U18146 ( .A1(n15063), .A2(n19182), .ZN(n15072) );
  AOI21_X1 U18147 ( .B1(n15089), .B2(n15075), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15064) );
  NOR2_X1 U18148 ( .A1(n15065), .A2(n15064), .ZN(n15069) );
  OAI21_X1 U18149 ( .B1(n15067), .B2(n16251), .A(n15066), .ZN(n15068) );
  AOI211_X1 U18150 ( .C1(n15070), .C2(n19199), .A(n15069), .B(n15068), .ZN(
        n15071) );
  OAI211_X1 U18151 ( .C1(n19202), .C2(n15073), .A(n15072), .B(n15071), .ZN(
        P2_U3016) );
  INV_X1 U18152 ( .A(n16074), .ZN(n15080) );
  INV_X1 U18153 ( .A(n15089), .ZN(n15074) );
  AOI211_X1 U18154 ( .C1(n15077), .C2(n15076), .A(n15075), .B(n15074), .ZN(
        n15078) );
  AOI211_X1 U18155 ( .C1(n15080), .C2(n19187), .A(n15079), .B(n15078), .ZN(
        n15082) );
  NAND2_X1 U18156 ( .A1(n15094), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15081) );
  OAI211_X1 U18157 ( .C1(n16070), .C2(n16266), .A(n15082), .B(n15081), .ZN(
        n15083) );
  AOI21_X1 U18158 ( .B1(n15084), .B2(n16231), .A(n15083), .ZN(n15085) );
  OAI21_X1 U18159 ( .B1(n15086), .B2(n19190), .A(n15085), .ZN(P2_U3017) );
  NAND3_X1 U18160 ( .A1(n14907), .A2(n19182), .A3(n15087), .ZN(n15096) );
  NAND2_X1 U18161 ( .A1(n15089), .A2(n15088), .ZN(n15090) );
  OAI211_X1 U18162 ( .C1(n16251), .C2(n16089), .A(n15091), .B(n15090), .ZN(
        n15093) );
  NOR2_X1 U18163 ( .A1(n16085), .A2(n16266), .ZN(n15092) );
  AOI211_X1 U18164 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15094), .A(
        n15093), .B(n15092), .ZN(n15095) );
  OAI211_X1 U18165 ( .C1(n15097), .C2(n19202), .A(n15096), .B(n15095), .ZN(
        P2_U3019) );
  INV_X1 U18166 ( .A(n15110), .ZN(n15100) );
  XNOR2_X1 U18167 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15099) );
  OAI21_X1 U18168 ( .B1(n15100), .B2(n15099), .A(n15098), .ZN(n15101) );
  AOI21_X1 U18169 ( .B1(n19187), .B2(n16104), .A(n15101), .ZN(n15102) );
  OAI21_X1 U18170 ( .B1(n15104), .B2(n15103), .A(n15102), .ZN(n15107) );
  NOR2_X1 U18171 ( .A1(n15105), .A2(n19202), .ZN(n15106) );
  AOI211_X1 U18172 ( .C1(n16093), .C2(n19199), .A(n15107), .B(n15106), .ZN(
        n15108) );
  OAI21_X1 U18173 ( .B1(n15109), .B2(n19190), .A(n15108), .ZN(P2_U3020) );
  AOI22_X1 U18174 ( .A1(n15110), .A2(n21137), .B1(n19000), .B2(
        P2_REIP_REG_25__SCAN_IN), .ZN(n15111) );
  OAI21_X1 U18175 ( .B1(n16251), .B2(n15112), .A(n15111), .ZN(n15115) );
  NOR2_X1 U18176 ( .A1(n15113), .A2(n16266), .ZN(n15114) );
  AOI211_X1 U18177 ( .C1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n15116), .A(
        n15115), .B(n15114), .ZN(n15120) );
  NAND3_X1 U18178 ( .A1(n15118), .A2(n16231), .A3(n15117), .ZN(n15119) );
  OAI211_X1 U18179 ( .C1(n15121), .C2(n19190), .A(n15120), .B(n15119), .ZN(
        P2_U3021) );
  INV_X1 U18180 ( .A(n18983), .ZN(n16243) );
  NAND2_X1 U18181 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n16243), .ZN(n15122) );
  OAI221_X1 U18182 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15125), 
        .C1(n15124), .C2(n15123), .A(n15122), .ZN(n15127) );
  OAI22_X1 U18183 ( .A1(n16110), .A2(n16266), .B1(n16251), .B2(n16109), .ZN(
        n15126) );
  AOI211_X1 U18184 ( .C1(n15128), .C2(n16231), .A(n15127), .B(n15126), .ZN(
        n15129) );
  OAI21_X1 U18185 ( .B1(n15130), .B2(n19190), .A(n15129), .ZN(P2_U3022) );
  XNOR2_X1 U18186 ( .A(n15131), .B(n15132), .ZN(n16140) );
  OR2_X1 U18187 ( .A1(n15307), .A2(n15133), .ZN(n15170) );
  INV_X1 U18188 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15141) );
  AOI21_X1 U18189 ( .B1(n15141), .B2(n10980), .A(n15134), .ZN(n15139) );
  NOR2_X1 U18190 ( .A1(n21110), .A2(n16226), .ZN(n15137) );
  NOR2_X1 U18191 ( .A1(n16251), .A2(n15135), .ZN(n15136) );
  AOI211_X1 U18192 ( .C1(n15139), .C2(n15138), .A(n15137), .B(n15136), .ZN(
        n15140) );
  OAI21_X1 U18193 ( .B1(n15170), .B2(n15141), .A(n15140), .ZN(n15145) );
  OR2_X1 U18194 ( .A1(n15159), .A2(n10980), .ZN(n16146) );
  NAND2_X1 U18195 ( .A1(n16146), .A2(n15141), .ZN(n15143) );
  NAND2_X1 U18196 ( .A1(n15143), .A2(n15142), .ZN(n16139) );
  NOR2_X1 U18197 ( .A1(n16139), .A2(n19202), .ZN(n15144) );
  AOI211_X1 U18198 ( .C1(n19199), .C2(n16142), .A(n15145), .B(n15144), .ZN(
        n15146) );
  OAI21_X1 U18199 ( .B1(n16140), .B2(n19190), .A(n15146), .ZN(P2_U3023) );
  NAND2_X1 U18200 ( .A1(n15149), .A2(n15148), .ZN(n15150) );
  XNOR2_X1 U18201 ( .A(n15147), .B(n15150), .ZN(n16150) );
  INV_X1 U18202 ( .A(n16150), .ZN(n15162) );
  NAND2_X1 U18203 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n16243), .ZN(n15151) );
  OAI221_X1 U18204 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15152), 
        .C1(n10980), .C2(n15170), .A(n15151), .ZN(n15158) );
  NOR2_X1 U18205 ( .A1(n15154), .A2(n15153), .ZN(n15155) );
  OR2_X1 U18206 ( .A1(n15156), .A2(n15155), .ZN(n16121) );
  OAI22_X1 U18207 ( .A1(n16148), .A2(n16266), .B1(n16251), .B2(n16121), .ZN(
        n15157) );
  NOR2_X1 U18208 ( .A1(n15158), .A2(n15157), .ZN(n15161) );
  NAND2_X1 U18209 ( .A1(n15159), .A2(n10980), .ZN(n16145) );
  NAND3_X1 U18210 ( .A1(n16146), .A2(n16145), .A3(n16231), .ZN(n15160) );
  OAI211_X1 U18211 ( .C1(n15162), .C2(n19190), .A(n15161), .B(n15160), .ZN(
        P2_U3024) );
  NOR2_X1 U18212 ( .A1(n15163), .A2(n16266), .ZN(n15164) );
  AOI211_X1 U18213 ( .C1(n19187), .C2(n15166), .A(n15165), .B(n15164), .ZN(
        n15168) );
  NAND4_X1 U18214 ( .A1(n15329), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n15180), .A4(n15169), .ZN(n15167) );
  OAI211_X1 U18215 ( .C1(n15170), .C2(n15169), .A(n15168), .B(n15167), .ZN(
        n15171) );
  AOI21_X1 U18216 ( .B1(n15172), .B2(n16231), .A(n15171), .ZN(n15173) );
  OAI21_X1 U18217 ( .B1(n15174), .B2(n19190), .A(n15173), .ZN(P2_U3025) );
  NOR2_X1 U18218 ( .A1(n19192), .A2(n15207), .ZN(n15175) );
  NOR2_X1 U18219 ( .A1(n15330), .A2(n15175), .ZN(n15210) );
  OR2_X1 U18220 ( .A1(n19192), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15176) );
  AND2_X1 U18221 ( .A1(n15210), .A2(n15176), .ZN(n15196) );
  AND3_X1 U18222 ( .A1(n15207), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15195), .ZN(n15177) );
  NAND2_X1 U18223 ( .A1(n15329), .A2(n15177), .ZN(n15193) );
  AOI21_X1 U18224 ( .B1(n15196), .B2(n15193), .A(n15179), .ZN(n15185) );
  AOI21_X1 U18225 ( .B1(n19187), .B2(n16127), .A(n15178), .ZN(n15182) );
  NAND3_X1 U18226 ( .A1(n15329), .A2(n15180), .A3(n15179), .ZN(n15181) );
  OAI211_X1 U18227 ( .C1(n15183), .C2(n16266), .A(n15182), .B(n15181), .ZN(
        n15184) );
  NOR2_X1 U18228 ( .A1(n15185), .A2(n15184), .ZN(n15188) );
  NAND2_X1 U18229 ( .A1(n15186), .A2(n16231), .ZN(n15187) );
  OAI211_X1 U18230 ( .C1(n15189), .C2(n19190), .A(n15188), .B(n15187), .ZN(
        P2_U3026) );
  INV_X1 U18231 ( .A(n15190), .ZN(n18883) );
  OAI21_X1 U18232 ( .B1(n16251), .B2(n18888), .A(n15191), .ZN(n15192) );
  AOI21_X1 U18233 ( .B1(n18883), .B2(n19199), .A(n15192), .ZN(n15194) );
  OAI211_X1 U18234 ( .C1(n15196), .C2(n15195), .A(n15194), .B(n15193), .ZN(
        n15197) );
  AOI21_X1 U18235 ( .B1(n15198), .B2(n16231), .A(n15197), .ZN(n15199) );
  OAI21_X1 U18236 ( .B1(n15200), .B2(n19190), .A(n15199), .ZN(P2_U3027) );
  AND2_X1 U18237 ( .A1(n15202), .A2(n15201), .ZN(n15204) );
  OR2_X1 U18238 ( .A1(n15204), .A2(n15203), .ZN(n18895) );
  NOR2_X1 U18239 ( .A1(n16251), .A2(n18895), .ZN(n15205) );
  AOI211_X1 U18240 ( .C1(n18897), .C2(n19199), .A(n15206), .B(n15205), .ZN(
        n15209) );
  NAND3_X1 U18241 ( .A1(n15329), .A2(n15207), .A3(n20943), .ZN(n15208) );
  OAI211_X1 U18242 ( .C1(n15210), .C2(n20943), .A(n15209), .B(n15208), .ZN(
        n15211) );
  AOI21_X1 U18243 ( .B1(n15212), .B2(n16231), .A(n15211), .ZN(n15213) );
  OAI21_X1 U18244 ( .B1(n15214), .B2(n19190), .A(n15213), .ZN(P2_U3028) );
  OAI21_X1 U18245 ( .B1(n16251), .B2(n18911), .A(n15215), .ZN(n15220) );
  NAND2_X1 U18246 ( .A1(n15329), .A2(n15258), .ZN(n15257) );
  OR2_X1 U18247 ( .A1(n15257), .A2(n15216), .ZN(n15281) );
  NOR3_X1 U18248 ( .A1(n15281), .A2(n15260), .A3(n15282), .ZN(n15253) );
  AOI22_X1 U18249 ( .A1(n15217), .A2(n16231), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15253), .ZN(n15237) );
  NOR3_X1 U18250 ( .A1(n15237), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15218), .ZN(n15219) );
  AOI211_X1 U18251 ( .C1(n18907), .C2(n19199), .A(n15220), .B(n15219), .ZN(
        n15229) );
  INV_X1 U18252 ( .A(n15307), .ZN(n15223) );
  OAI21_X1 U18253 ( .B1(n15330), .B2(n15224), .A(n15223), .ZN(n15249) );
  OAI211_X1 U18254 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15226), .A(
        n15225), .B(n15249), .ZN(n15240) );
  NOR2_X1 U18255 ( .A1(n19192), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15227) );
  OAI21_X1 U18256 ( .B1(n15240), .B2(n15227), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15228) );
  OAI211_X1 U18257 ( .C1(n15230), .C2(n19190), .A(n15229), .B(n15228), .ZN(
        P2_U3029) );
  OR2_X1 U18258 ( .A1(n15232), .A2(n15231), .ZN(n15233) );
  AND2_X1 U18259 ( .A1(n15234), .A2(n15233), .ZN(n19054) );
  OAI22_X1 U18260 ( .A1(n15236), .A2(n16266), .B1(n15235), .B2(n16226), .ZN(
        n15239) );
  NOR2_X1 U18261 ( .A1(n15237), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15238) );
  AOI211_X1 U18262 ( .C1(n19187), .C2(n19054), .A(n15239), .B(n15238), .ZN(
        n15242) );
  NAND2_X1 U18263 ( .A1(n15240), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15241) );
  OAI211_X1 U18264 ( .C1(n15243), .C2(n19190), .A(n15242), .B(n15241), .ZN(
        P2_U3030) );
  NAND2_X1 U18265 ( .A1(n15244), .A2(n16231), .ZN(n15255) );
  NAND2_X1 U18266 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n16243), .ZN(n15247) );
  OR2_X1 U18267 ( .A1(n16251), .A2(n15245), .ZN(n15246) );
  OAI211_X1 U18268 ( .C1(n15248), .C2(n16266), .A(n15247), .B(n15246), .ZN(
        n15251) );
  NOR2_X1 U18269 ( .A1(n15249), .A2(n15252), .ZN(n15250) );
  AOI211_X1 U18270 ( .C1(n15253), .C2(n15252), .A(n15251), .B(n15250), .ZN(
        n15254) );
  OAI211_X1 U18271 ( .C1(n15256), .C2(n19190), .A(n15255), .B(n15254), .ZN(
        P2_U3031) );
  INV_X1 U18272 ( .A(n15257), .ZN(n15299) );
  OAI21_X1 U18273 ( .B1(n15258), .B2(n19192), .A(n15308), .ZN(n15296) );
  AOI21_X1 U18274 ( .B1(n15299), .B2(n15259), .A(n15296), .ZN(n15280) );
  NOR2_X1 U18275 ( .A1(n15280), .A2(n15260), .ZN(n15269) );
  INV_X1 U18276 ( .A(n15281), .ZN(n15261) );
  NAND3_X1 U18277 ( .A1(n15261), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n15260), .ZN(n15266) );
  INV_X1 U18278 ( .A(n15262), .ZN(n15264) );
  AOI21_X1 U18279 ( .B1(n19199), .B2(n15264), .A(n15263), .ZN(n15265) );
  OAI211_X1 U18280 ( .C1(n16251), .C2(n15267), .A(n15266), .B(n15265), .ZN(
        n15268) );
  AOI211_X1 U18281 ( .C1(n15270), .C2(n19182), .A(n15269), .B(n15268), .ZN(
        n15271) );
  OAI21_X1 U18282 ( .B1(n15272), .B2(n19202), .A(n15271), .ZN(P2_U3032) );
  NOR2_X1 U18283 ( .A1(n15303), .A2(n15216), .ZN(n16161) );
  INV_X1 U18284 ( .A(n15273), .ZN(n15274) );
  OAI21_X1 U18285 ( .B1(n16161), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15274), .ZN(n16155) );
  NAND2_X1 U18286 ( .A1(n15275), .A2(n15291), .ZN(n15279) );
  NAND2_X1 U18287 ( .A1(n15277), .A2(n15276), .ZN(n15278) );
  XNOR2_X1 U18288 ( .A(n15279), .B(n15278), .ZN(n16154) );
  INV_X1 U18289 ( .A(n16154), .ZN(n15288) );
  AOI21_X1 U18290 ( .B1(n15282), .B2(n15281), .A(n15280), .ZN(n15285) );
  NOR2_X1 U18291 ( .A1(n16226), .A2(n15283), .ZN(n15284) );
  AOI211_X1 U18292 ( .C1(n19199), .C2(n18933), .A(n15285), .B(n15284), .ZN(
        n15286) );
  OAI21_X1 U18293 ( .B1(n16251), .B2(n18936), .A(n15286), .ZN(n15287) );
  AOI21_X1 U18294 ( .B1(n15288), .B2(n19182), .A(n15287), .ZN(n15289) );
  OAI21_X1 U18295 ( .B1(n16155), .B2(n19202), .A(n15289), .ZN(P2_U3033) );
  NAND2_X1 U18296 ( .A1(n15291), .A2(n15290), .ZN(n15292) );
  XNOR2_X1 U18297 ( .A(n15293), .B(n15292), .ZN(n16162) );
  AND2_X1 U18298 ( .A1(n15303), .A2(n15216), .ZN(n16160) );
  OR3_X1 U18299 ( .A1(n16160), .A2(n16161), .A3(n19202), .ZN(n15301) );
  INV_X1 U18300 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19861) );
  NOR2_X1 U18301 ( .A1(n19861), .A2(n16226), .ZN(n15295) );
  NOR2_X1 U18302 ( .A1(n16266), .A2(n18942), .ZN(n15294) );
  AOI211_X1 U18303 ( .C1(n15296), .C2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15295), .B(n15294), .ZN(n15297) );
  OAI21_X1 U18304 ( .B1(n16251), .B2(n18941), .A(n15297), .ZN(n15298) );
  AOI21_X1 U18305 ( .B1(n15299), .B2(n15216), .A(n15298), .ZN(n15300) );
  OAI211_X1 U18306 ( .C1(n16162), .C2(n19190), .A(n15301), .B(n15300), .ZN(
        P2_U3034) );
  INV_X1 U18307 ( .A(n15302), .ZN(n16175) );
  OAI21_X1 U18308 ( .B1(n16175), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15303), .ZN(n16169) );
  XNOR2_X1 U18309 ( .A(n15305), .B(n15310), .ZN(n15306) );
  XNOR2_X1 U18310 ( .A(n15304), .B(n15306), .ZN(n16168) );
  AOI21_X1 U18311 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15308), .A(
        n15307), .ZN(n16230) );
  NOR2_X1 U18312 ( .A1(n12187), .A2(n16226), .ZN(n15312) );
  NAND2_X1 U18313 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15329), .ZN(
        n16227) );
  AOI211_X1 U18314 ( .C1(n16177), .C2(n15310), .A(n15309), .B(n16227), .ZN(
        n15311) );
  AOI211_X1 U18315 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n16230), .A(
        n15312), .B(n15311), .ZN(n15317) );
  OAI22_X1 U18316 ( .A1(n16266), .A2(n15314), .B1(n16251), .B2(n15313), .ZN(
        n15315) );
  INV_X1 U18317 ( .A(n15315), .ZN(n15316) );
  OAI211_X1 U18318 ( .C1(n16168), .C2(n19190), .A(n15317), .B(n15316), .ZN(
        n15318) );
  INV_X1 U18319 ( .A(n15318), .ZN(n15319) );
  OAI21_X1 U18320 ( .B1(n16169), .B2(n19202), .A(n15319), .ZN(P2_U3035) );
  OAI21_X1 U18321 ( .B1(n15320), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16176), .ZN(n16190) );
  INV_X1 U18322 ( .A(n15321), .ZN(n16178) );
  OR2_X1 U18323 ( .A1(n16178), .A2(n15322), .ZN(n15323) );
  XNOR2_X1 U18324 ( .A(n15324), .B(n15323), .ZN(n16189) );
  INV_X1 U18325 ( .A(n16192), .ZN(n18966) );
  OR2_X1 U18326 ( .A1(n16251), .A2(n18965), .ZN(n15326) );
  OR2_X1 U18327 ( .A1(n12161), .A2(n18983), .ZN(n15325) );
  OAI211_X1 U18328 ( .C1(n16266), .C2(n18966), .A(n15326), .B(n15325), .ZN(
        n15327) );
  AOI21_X1 U18329 ( .B1(n15329), .B2(n15328), .A(n15327), .ZN(n15332) );
  NAND2_X1 U18330 ( .A1(n15330), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15331) );
  OAI211_X1 U18331 ( .C1(n16189), .C2(n19190), .A(n15332), .B(n15331), .ZN(
        n15333) );
  INV_X1 U18332 ( .A(n15333), .ZN(n15334) );
  OAI21_X1 U18333 ( .B1(n16190), .B2(n19202), .A(n15334), .ZN(P2_U3037) );
  NAND3_X1 U18334 ( .A1(n15336), .A2(n15335), .A3(n16231), .ZN(n15343) );
  OAI21_X1 U18335 ( .B1(n19192), .B2(n15338), .A(n16261), .ZN(n16238) );
  NAND2_X1 U18336 ( .A1(n19199), .A2(n18976), .ZN(n15340) );
  AND2_X1 U18337 ( .A1(n15338), .A2(n15337), .ZN(n16244) );
  AOI22_X1 U18338 ( .A1(n19000), .A2(P2_REIP_REG_7__SCAN_IN), .B1(n16244), 
        .B2(n16245), .ZN(n15339) );
  OAI211_X1 U18339 ( .C1(n16251), .C2(n18977), .A(n15340), .B(n15339), .ZN(
        n15341) );
  AOI21_X1 U18340 ( .B1(n16238), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n15341), .ZN(n15342) );
  OAI211_X1 U18341 ( .C1(n15344), .C2(n19190), .A(n15343), .B(n15342), .ZN(
        P2_U3039) );
  OAI21_X1 U18342 ( .B1(n15346), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15345), .ZN(n16212) );
  XOR2_X1 U18343 ( .A(n15348), .B(n15347), .Z(n16214) );
  NAND2_X1 U18344 ( .A1(n16214), .A2(n19182), .ZN(n15357) );
  NOR2_X1 U18345 ( .A1(n15350), .A2(n15349), .ZN(n15355) );
  NAND2_X1 U18346 ( .A1(n16238), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15352) );
  AOI22_X1 U18347 ( .A1(n19199), .A2(n18991), .B1(n19000), .B2(
        P2_REIP_REG_6__SCAN_IN), .ZN(n15351) );
  OAI211_X1 U18348 ( .C1(n16251), .C2(n18995), .A(n15352), .B(n15351), .ZN(
        n15353) );
  AOI21_X1 U18349 ( .B1(n15355), .B2(n15354), .A(n15353), .ZN(n15356) );
  OAI211_X1 U18350 ( .C1(n16212), .C2(n19202), .A(n15357), .B(n15356), .ZN(
        P2_U3040) );
  NAND2_X1 U18351 ( .A1(n19169), .A2(n15358), .ZN(n15369) );
  NAND2_X1 U18352 ( .A1(n15360), .A2(n15359), .ZN(n15366) );
  NOR2_X1 U18353 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15363) );
  INV_X1 U18354 ( .A(n15361), .ZN(n15362) );
  OAI22_X1 U18355 ( .A1(n15364), .A2(n15363), .B1(n15362), .B2(n15366), .ZN(
        n15365) );
  AOI21_X1 U18356 ( .B1(n15367), .B2(n15366), .A(n15365), .ZN(n15368) );
  NAND2_X1 U18357 ( .A1(n15369), .A2(n15368), .ZN(n16281) );
  INV_X1 U18358 ( .A(n15370), .ZN(n15372) );
  NOR2_X1 U18359 ( .A1(n15372), .A2(n15371), .ZN(n15373) );
  AOI21_X1 U18360 ( .B1(n16281), .B2(n19817), .A(n15373), .ZN(n15374) );
  OAI21_X1 U18361 ( .B1(n19909), .B2(n15375), .A(n15374), .ZN(n15377) );
  MUX2_X1 U18362 ( .A(n15377), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15376), .Z(P2_U3599) );
  INV_X2 U18363 ( .A(n9783), .ZN(n17124) );
  NOR2_X2 U18364 ( .A1(n15386), .A2(n16885), .ZN(n15672) );
  INV_X4 U18365 ( .A(n15682), .ZN(n17155) );
  AOI22_X1 U18366 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15383) );
  NOR2_X1 U18367 ( .A1(n15386), .A2(n16884), .ZN(n15378) );
  INV_X2 U18368 ( .A(n16981), .ZN(n17147) );
  AOI22_X1 U18369 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15382) );
  AOI22_X1 U18370 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15381) );
  NAND3_X1 U18371 ( .A1(n18818), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n18635), .ZN(n17008) );
  AOI22_X1 U18372 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17167), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15380) );
  NAND4_X1 U18373 ( .A1(n15383), .A2(n15382), .A3(n15381), .A4(n15380), .ZN(
        n15395) );
  NOR2_X2 U18374 ( .A1(n15385), .A2(n15388), .ZN(n15484) );
  CLKBUF_X3 U18375 ( .A(n15484), .Z(n17154) );
  AOI22_X1 U18376 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15393) );
  INV_X2 U18377 ( .A(n15458), .ZN(n17156) );
  NOR2_X2 U18378 ( .A1(n15384), .A2(n15387), .ZN(n15670) );
  BUF_X4 U18379 ( .A(n15670), .Z(n17165) );
  AOI22_X1 U18380 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15392) );
  AOI22_X1 U18381 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9735), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15391) );
  INV_X2 U18382 ( .A(n9776), .ZN(n17148) );
  AOI22_X1 U18383 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15390) );
  NAND4_X1 U18384 ( .A1(n15393), .A2(n15392), .A3(n15391), .A4(n15390), .ZN(
        n15394) );
  AOI22_X1 U18385 ( .A1(n9735), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(n9734), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15400) );
  AOI22_X1 U18386 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15399) );
  INV_X2 U18387 ( .A(n15669), .ZN(n17123) );
  AOI22_X1 U18388 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15398) );
  AOI22_X1 U18389 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15397) );
  NAND4_X1 U18390 ( .A1(n15400), .A2(n15399), .A3(n15398), .A4(n15397), .ZN(
        n15407) );
  AOI22_X1 U18391 ( .A1(n17170), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15405) );
  INV_X2 U18392 ( .A(n17169), .ZN(n17089) );
  AOI22_X1 U18393 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15404) );
  AOI22_X1 U18394 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15403) );
  AOI22_X1 U18395 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15402) );
  NAND4_X1 U18396 ( .A1(n15405), .A2(n15404), .A3(n15403), .A4(n15402), .ZN(
        n15406) );
  AOI22_X1 U18397 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17123), .ZN(n15417) );
  AOI22_X1 U18398 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15416) );
  INV_X1 U18399 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17184) );
  AOI22_X1 U18400 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17154), .B1(
        n9735), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15408) );
  OAI21_X1 U18401 ( .B1(n9776), .B2(n17184), .A(n15408), .ZN(n15414) );
  AOI22_X1 U18402 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n17165), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n9734), .ZN(n15412) );
  AOI22_X1 U18403 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n17166), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15411) );
  AOI22_X1 U18404 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17089), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15410) );
  AOI22_X1 U18405 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n17155), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n17049), .ZN(n15409) );
  NAND4_X1 U18406 ( .A1(n15412), .A2(n15411), .A3(n15410), .A4(n15409), .ZN(
        n15413) );
  AOI22_X1 U18407 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15484), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15427) );
  INV_X2 U18408 ( .A(n17169), .ZN(n17075) );
  AOI22_X1 U18409 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15426) );
  AOI22_X1 U18410 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15418) );
  OAI21_X1 U18411 ( .B1(n15694), .B2(n21030), .A(n15418), .ZN(n15424) );
  AOI22_X1 U18412 ( .A1(n9735), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15422) );
  AOI22_X1 U18413 ( .A1(n17080), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15421) );
  AOI22_X1 U18414 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15420) );
  AOI22_X1 U18415 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15419) );
  NAND4_X1 U18416 ( .A1(n15422), .A2(n15421), .A3(n15420), .A4(n15419), .ZN(
        n15423) );
  AOI211_X1 U18417 ( .C1(n17148), .C2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A(
        n15424), .B(n15423), .ZN(n15425) );
  INV_X1 U18418 ( .A(n15601), .ZN(n15468) );
  AOI22_X1 U18419 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15436) );
  AOI22_X1 U18420 ( .A1(n15645), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15435) );
  AOI22_X1 U18421 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9735), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15428) );
  OAI21_X1 U18422 ( .B1(n17169), .B2(n20976), .A(n15428), .ZN(n15434) );
  AOI22_X1 U18423 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15432) );
  AOI22_X1 U18424 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15431) );
  AOI22_X1 U18425 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15430) );
  AOI22_X1 U18426 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15670), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15429) );
  NAND4_X1 U18427 ( .A1(n15432), .A2(n15431), .A3(n15430), .A4(n15429), .ZN(
        n15433) );
  AOI22_X1 U18428 ( .A1(n17170), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15440) );
  AOI22_X1 U18429 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9735), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15439) );
  AOI22_X1 U18430 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15438) );
  AOI22_X1 U18431 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15437) );
  NAND4_X1 U18432 ( .A1(n15440), .A2(n15439), .A3(n15438), .A4(n15437), .ZN(
        n15446) );
  BUF_X1 U18433 ( .A(n15533), .Z(n17047) );
  AOI22_X1 U18434 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17047), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15444) );
  AOI22_X1 U18435 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15443) );
  AOI22_X1 U18436 ( .A1(n17080), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15484), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15442) );
  AOI22_X1 U18437 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15672), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15441) );
  NAND4_X1 U18438 ( .A1(n15444), .A2(n15443), .A3(n15442), .A4(n15441), .ZN(
        n15445) );
  AOI22_X1 U18439 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15456) );
  AOI22_X1 U18440 ( .A1(n9735), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n15672), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n15455) );
  INV_X1 U18441 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17191) );
  AOI22_X1 U18442 ( .A1(n17080), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15447) );
  OAI21_X1 U18443 ( .B1(n9776), .B2(n17191), .A(n15447), .ZN(n15453) );
  AOI22_X1 U18444 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15451) );
  AOI22_X1 U18445 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15450) );
  AOI22_X1 U18446 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n15484), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15449) );
  AOI22_X1 U18447 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15448) );
  NAND4_X1 U18448 ( .A1(n15451), .A2(n15450), .A3(n15449), .A4(n15448), .ZN(
        n15452) );
  AOI211_X1 U18449 ( .C1(n15645), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n15453), .B(n15452), .ZN(n15454) );
  NAND3_X1 U18450 ( .A1(n15456), .A2(n15455), .A3(n15454), .ZN(n17222) );
  AOI22_X1 U18451 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15467) );
  AOI22_X1 U18452 ( .A1(n17080), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n15672), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15466) );
  INV_X1 U18453 ( .A(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n21112) );
  AOI22_X1 U18454 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15457) );
  OAI21_X1 U18455 ( .B1(n15458), .B2(n21112), .A(n15457), .ZN(n15464) );
  AOI22_X1 U18456 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9735), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15462) );
  AOI22_X1 U18457 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15461) );
  AOI22_X1 U18458 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15460) );
  AOI22_X1 U18459 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15459) );
  NAND4_X1 U18460 ( .A1(n15462), .A2(n15461), .A3(n15460), .A4(n15459), .ZN(
        n15463) );
  AOI211_X1 U18461 ( .C1(n17146), .C2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n15464), .B(n15463), .ZN(n15465) );
  NAND3_X1 U18462 ( .A1(n15467), .A2(n15466), .A3(n15465), .ZN(n15561) );
  NAND2_X1 U18463 ( .A1(n18215), .A2(n15561), .ZN(n18621) );
  AOI22_X1 U18464 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n18646), .B2(n18811), .ZN(
        n15577) );
  AOI22_X1 U18465 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21113), .B1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18803), .ZN(n15476) );
  NAND2_X1 U18466 ( .A1(n18477), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15578) );
  OR2_X1 U18467 ( .A1(n15577), .A2(n15578), .ZN(n15469) );
  NAND2_X1 U18468 ( .A1(n15476), .A2(n15477), .ZN(n15470) );
  OAI21_X1 U18469 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18803), .A(
        n15470), .ZN(n15471) );
  OAI22_X1 U18470 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18665), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n15471), .ZN(n15473) );
  NOR2_X1 U18471 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18665), .ZN(
        n15472) );
  NAND2_X1 U18472 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n15471), .ZN(
        n15474) );
  AOI22_X1 U18473 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15473), .B1(
        n15472), .B2(n15474), .ZN(n15478) );
  OAI211_X1 U18474 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18477), .A(
        n15478), .B(n15578), .ZN(n15605) );
  AOI21_X1 U18475 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15474), .A(
        n15473), .ZN(n15475) );
  XOR2_X1 U18476 ( .A(n15477), .B(n15476), .Z(n15607) );
  NAND2_X1 U18477 ( .A1(n15478), .A2(n15607), .ZN(n15580) );
  OAI211_X1 U18478 ( .C1(n15577), .C2(n15605), .A(n15579), .B(n15580), .ZN(
        n16340) );
  INV_X1 U18479 ( .A(n16340), .ZN(n18660) );
  NOR2_X1 U18480 ( .A1(n15574), .A2(n15608), .ZN(n18623) );
  NAND3_X1 U18481 ( .A1(n18210), .A2(n18623), .A3(n17222), .ZN(n15559) );
  NOR3_X1 U18482 ( .A1(n17263), .A2(n15561), .A3(n15559), .ZN(n15479) );
  AOI22_X1 U18483 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n15672), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15483) );
  AOI22_X1 U18484 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15482) );
  AOI22_X1 U18485 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15481) );
  AOI22_X1 U18486 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15480) );
  NAND4_X1 U18487 ( .A1(n15483), .A2(n15482), .A3(n15481), .A4(n15480), .ZN(
        n15490) );
  AOI22_X1 U18488 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15488) );
  AOI22_X1 U18489 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9735), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15487) );
  AOI22_X1 U18490 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15484), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15486) );
  AOI22_X1 U18491 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17047), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15485) );
  NAND4_X1 U18492 ( .A1(n15488), .A2(n15487), .A3(n15486), .A4(n15485), .ZN(
        n15489) );
  NOR2_X1 U18493 ( .A1(n15490), .A2(n15489), .ZN(n16942) );
  AOI22_X1 U18494 ( .A1(n15645), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15495) );
  AOI22_X1 U18495 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15494) );
  AOI22_X1 U18496 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15493) );
  AOI22_X1 U18497 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15672), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15492) );
  NAND4_X1 U18498 ( .A1(n15495), .A2(n15494), .A3(n15493), .A4(n15492), .ZN(
        n15501) );
  AOI22_X1 U18499 ( .A1(n9735), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15499) );
  AOI22_X1 U18500 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15498) );
  AOI22_X1 U18501 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15497) );
  AOI22_X1 U18502 ( .A1(n17170), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15496) );
  NAND4_X1 U18503 ( .A1(n15499), .A2(n15498), .A3(n15497), .A4(n15496), .ZN(
        n15500) );
  NOR2_X1 U18504 ( .A1(n15501), .A2(n15500), .ZN(n16953) );
  AOI22_X1 U18505 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15505) );
  AOI22_X1 U18506 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15670), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15504) );
  AOI22_X1 U18507 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15503) );
  AOI22_X1 U18508 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15502) );
  NAND4_X1 U18509 ( .A1(n15505), .A2(n15504), .A3(n15503), .A4(n15502), .ZN(
        n15511) );
  AOI22_X1 U18510 ( .A1(n17170), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15672), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15509) );
  AOI22_X1 U18511 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9735), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15508) );
  AOI22_X1 U18512 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15507) );
  AOI22_X1 U18513 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15506) );
  NAND4_X1 U18514 ( .A1(n15509), .A2(n15508), .A3(n15507), .A4(n15506), .ZN(
        n15510) );
  NOR2_X1 U18515 ( .A1(n15511), .A2(n15510), .ZN(n16964) );
  AOI22_X1 U18516 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17154), .ZN(n15515) );
  AOI22_X1 U18517 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n9735), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n17124), .ZN(n15514) );
  AOI22_X1 U18518 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n17165), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n9734), .ZN(n15513) );
  AOI22_X1 U18519 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n17049), .ZN(n15512) );
  NAND4_X1 U18520 ( .A1(n15515), .A2(n15514), .A3(n15513), .A4(n15512), .ZN(
        n15521) );
  AOI22_X1 U18521 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15519) );
  AOI22_X1 U18522 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17166), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n17155), .ZN(n15518) );
  AOI22_X1 U18523 ( .A1(n15645), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15517) );
  AOI22_X1 U18524 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n17107), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17147), .ZN(n15516) );
  NAND4_X1 U18525 ( .A1(n15519), .A2(n15518), .A3(n15517), .A4(n15516), .ZN(
        n15520) );
  NOR2_X1 U18526 ( .A1(n15521), .A2(n15520), .ZN(n16963) );
  NOR2_X1 U18527 ( .A1(n16964), .A2(n16963), .ZN(n16959) );
  AOI22_X1 U18528 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15531) );
  AOI22_X1 U18529 ( .A1(n17170), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9735), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15530) );
  INV_X1 U18530 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n21063) );
  AOI22_X1 U18531 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15522) );
  OAI21_X1 U18532 ( .B1(n15682), .B2(n21063), .A(n15522), .ZN(n15528) );
  AOI22_X1 U18533 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15526) );
  AOI22_X1 U18534 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15525) );
  AOI22_X1 U18535 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15524) );
  AOI22_X1 U18536 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15523) );
  NAND4_X1 U18537 ( .A1(n15526), .A2(n15525), .A3(n15524), .A4(n15523), .ZN(
        n15527) );
  AOI211_X1 U18538 ( .C1(n17075), .C2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n15528), .B(n15527), .ZN(n15529) );
  NAND3_X1 U18539 ( .A1(n15531), .A2(n15530), .A3(n15529), .ZN(n16958) );
  NAND2_X1 U18540 ( .A1(n16959), .A2(n16958), .ZN(n16957) );
  NOR2_X1 U18541 ( .A1(n16953), .A2(n16957), .ZN(n16949) );
  AOI22_X1 U18542 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15542) );
  AOI22_X1 U18543 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15541) );
  INV_X1 U18544 ( .A(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n20993) );
  AOI22_X1 U18545 ( .A1(n9735), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15532) );
  OAI21_X1 U18546 ( .B1(n9783), .B2(n20993), .A(n15532), .ZN(n15539) );
  AOI22_X1 U18547 ( .A1(n15645), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15537) );
  AOI22_X1 U18548 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15670), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15536) );
  AOI22_X1 U18549 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15535) );
  AOI22_X1 U18550 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15534) );
  NAND4_X1 U18551 ( .A1(n15537), .A2(n15536), .A3(n15535), .A4(n15534), .ZN(
        n15538) );
  AOI211_X1 U18552 ( .C1(n17146), .C2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n15539), .B(n15538), .ZN(n15540) );
  NAND3_X1 U18553 ( .A1(n15542), .A2(n15541), .A3(n15540), .ZN(n16948) );
  NAND2_X1 U18554 ( .A1(n16949), .A2(n16948), .ZN(n16947) );
  NOR2_X1 U18555 ( .A1(n16942), .A2(n16947), .ZN(n16941) );
  AOI22_X1 U18556 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15552) );
  AOI22_X1 U18557 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15672), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15551) );
  INV_X1 U18558 ( .A(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n20949) );
  AOI22_X1 U18559 ( .A1(n9735), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n9734), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15543) );
  OAI21_X1 U18560 ( .B1(n9776), .B2(n20949), .A(n15543), .ZN(n15549) );
  AOI22_X1 U18561 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15547) );
  AOI22_X1 U18562 ( .A1(n15645), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15484), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15546) );
  AOI22_X1 U18563 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15545) );
  AOI22_X1 U18564 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15670), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15544) );
  NAND4_X1 U18565 ( .A1(n15547), .A2(n15546), .A3(n15545), .A4(n15544), .ZN(
        n15548) );
  AOI211_X1 U18566 ( .C1(n17075), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n15549), .B(n15548), .ZN(n15550) );
  NAND3_X1 U18567 ( .A1(n15552), .A2(n15551), .A3(n15550), .ZN(n16933) );
  XNOR2_X1 U18568 ( .A(n16941), .B(n16933), .ZN(n17237) );
  INV_X1 U18569 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16945) );
  INV_X1 U18570 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16901) );
  INV_X1 U18571 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17115) );
  INV_X1 U18572 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16796) );
  INV_X1 U18573 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17188) );
  NAND4_X1 U18574 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .A4(P3_EBX_REG_2__SCAN_IN), .ZN(n17202) );
  NAND4_X1 U18575 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(P3_EBX_REG_17__SCAN_IN), 
        .A3(P3_EBX_REG_16__SCAN_IN), .A4(n17059), .ZN(n17019) );
  INV_X1 U18576 ( .A(n17019), .ZN(n16993) );
  AND4_X1 U18577 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n16903)
         );
  NAND2_X1 U18578 ( .A1(n16991), .A2(n16903), .ZN(n16952) );
  INV_X1 U18579 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n21075) );
  OAI21_X1 U18580 ( .B1(n16945), .B2(n16946), .A(n21075), .ZN(n15553) );
  NOR2_X1 U18581 ( .A1(n21075), .A2(n16945), .ZN(n16937) );
  NAND2_X1 U18582 ( .A1(n18222), .A2(n17212), .ZN(n17218) );
  NAND2_X1 U18583 ( .A1(n15553), .A2(n16938), .ZN(n15554) );
  OAI21_X1 U18584 ( .B1(n17197), .B2(n17237), .A(n15554), .ZN(P3_U2675) );
  NOR2_X1 U18585 ( .A1(n21113), .A2(n18646), .ZN(n18356) );
  INV_X1 U18586 ( .A(n18356), .ZN(n18185) );
  AOI221_X1 U18587 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18185), .C1(n15556), 
        .C2(n18185), .A(n15555), .ZN(n18179) );
  NOR2_X1 U18588 ( .A1(n15557), .A2(n18646), .ZN(n15558) );
  OAI21_X1 U18589 ( .B1(n15558), .B2(n18267), .A(n18180), .ZN(n18177) );
  AOI22_X1 U18590 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18179), .B1(
        n18177), .B2(n21113), .ZN(P3_U2865) );
  NAND2_X1 U18591 ( .A1(n17416), .A2(n16523), .ZN(n15582) );
  NAND2_X1 U18592 ( .A1(n18183), .A2(n17263), .ZN(n15571) );
  NOR2_X1 U18593 ( .A1(n15571), .A2(n15559), .ZN(n15562) );
  NAND2_X1 U18594 ( .A1(n15560), .A2(n17222), .ZN(n15568) );
  NOR4_X1 U18595 ( .A1(n15574), .A2(n15561), .A3(n15571), .A4(n15568), .ZN(
        n15575) );
  AND2_X1 U18596 ( .A1(n15575), .A2(n15608), .ZN(n15587) );
  NOR2_X1 U18597 ( .A1(n18210), .A2(n17222), .ZN(n18642) );
  OAI211_X1 U18598 ( .C1(n18222), .C2(n18642), .A(n18835), .B(n17377), .ZN(
        n15590) );
  NAND2_X1 U18599 ( .A1(n18210), .A2(n15564), .ZN(n15583) );
  NAND3_X1 U18600 ( .A1(n18197), .A2(n15590), .A3(n15583), .ZN(n15573) );
  NAND2_X1 U18601 ( .A1(n18183), .A2(n16523), .ZN(n15584) );
  NAND2_X1 U18602 ( .A1(n18197), .A2(n15584), .ZN(n15566) );
  AOI21_X1 U18603 ( .B1(n18197), .B2(n18183), .A(n18642), .ZN(n15563) );
  AOI21_X1 U18604 ( .B1(n15564), .B2(n15568), .A(n15563), .ZN(n15565) );
  AOI21_X1 U18605 ( .B1(n15568), .B2(n15566), .A(n15565), .ZN(n15567) );
  INV_X1 U18606 ( .A(n15567), .ZN(n15570) );
  AOI21_X1 U18607 ( .B1(n17263), .B2(n15568), .A(n18206), .ZN(n15569) );
  AOI211_X2 U18608 ( .C1(n15571), .C2(n18200), .A(n15570), .B(n15569), .ZN(
        n15588) );
  INV_X1 U18609 ( .A(n15588), .ZN(n15572) );
  NAND2_X1 U18610 ( .A1(n15575), .A2(n15599), .ZN(n15603) );
  INV_X1 U18611 ( .A(n15603), .ZN(n15576) );
  NAND2_X1 U18612 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18836) );
  XNOR2_X1 U18613 ( .A(n15578), .B(n15577), .ZN(n15581) );
  AND2_X1 U18614 ( .A1(n18660), .A2(n15602), .ZN(n15593) );
  NOR2_X2 U18615 ( .A1(n18700), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18773) );
  NOR2_X1 U18616 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18698) );
  NOR4_X1 U18617 ( .A1(n18707), .A2(n18654), .A3(n17376), .A4(n18833), .ZN(
        n15592) );
  OAI211_X1 U18618 ( .C1(n18206), .C2(n18215), .A(n15584), .B(n15583), .ZN(
        n15585) );
  NOR2_X1 U18619 ( .A1(n15586), .A2(n15585), .ZN(n15752) );
  AOI21_X1 U18620 ( .B1(n15752), .B2(n15588), .A(n15587), .ZN(n15589) );
  INV_X1 U18621 ( .A(n15589), .ZN(n15591) );
  NAND2_X1 U18622 ( .A1(n15591), .A2(n15590), .ZN(n15614) );
  NOR4_X2 U18623 ( .A1(n9725), .A2(n15593), .A3(n15592), .A4(n15614), .ZN(
        n18668) );
  INV_X1 U18624 ( .A(n18668), .ZN(n18640) );
  NOR2_X1 U18625 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18787), .ZN(n18182) );
  INV_X1 U18626 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18175) );
  NOR2_X1 U18627 ( .A1(n18175), .A2(n18785), .ZN(n15594) );
  INV_X1 U18628 ( .A(n18819), .ZN(n18816) );
  INV_X1 U18629 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15597) );
  INV_X1 U18630 ( .A(n18845), .ZN(n18808) );
  NOR2_X1 U18631 ( .A1(n15595), .A2(n16515), .ZN(n18667) );
  NAND3_X1 U18632 ( .A1(n18816), .A2(n18808), .A3(n18667), .ZN(n15596) );
  OAI21_X1 U18633 ( .B1(n18816), .B2(n15597), .A(n15596), .ZN(P3_U3284) );
  INV_X1 U18634 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17871) );
  INV_X1 U18635 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17490) );
  NOR2_X1 U18636 ( .A1(n17871), .A2(n17490), .ZN(n16367) );
  NAND2_X1 U18637 ( .A1(n16523), .A2(n16514), .ZN(n15600) );
  OAI21_X1 U18638 ( .B1(n15601), .B2(n15600), .A(n15599), .ZN(n18622) );
  AOI21_X2 U18639 ( .B1(n18623), .B2(n15604), .A(n18622), .ZN(n18057) );
  NAND2_X1 U18640 ( .A1(n18197), .A2(n16523), .ZN(n15609) );
  NOR2_X1 U18641 ( .A1(n18215), .A2(n15609), .ZN(n15753) );
  INV_X1 U18642 ( .A(n15605), .ZN(n15606) );
  NAND2_X1 U18643 ( .A1(n15607), .A2(n15606), .ZN(n16337) );
  AOI21_X1 U18644 ( .B1(n18835), .B2(n15608), .A(n16518), .ZN(n15610) );
  AOI21_X1 U18645 ( .B1(n15610), .B2(n15609), .A(n18707), .ZN(n16496) );
  AOI22_X1 U18646 ( .A1(n15753), .A2(n16337), .B1(n16496), .B2(n15611), .ZN(
        n15612) );
  OAI22_X1 U18647 ( .A1(n15612), .A2(n18654), .B1(n16340), .B2(n15611), .ZN(
        n15613) );
  NAND2_X1 U18648 ( .A1(n18001), .A2(n18154), .ZN(n18130) );
  NAND2_X1 U18649 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18055) );
  INV_X1 U18650 ( .A(n18055), .ZN(n17730) );
  NAND2_X1 U18651 ( .A1(n17730), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18035) );
  INV_X1 U18652 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18048) );
  NOR2_X1 U18653 ( .A1(n18035), .A2(n18048), .ZN(n18032) );
  INV_X1 U18654 ( .A(n18032), .ZN(n18014) );
  NAND2_X1 U18655 ( .A1(n18015), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17990) );
  INV_X1 U18656 ( .A(n17990), .ZN(n17662) );
  AOI22_X1 U18657 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17089), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15624) );
  AOI22_X1 U18658 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15623) );
  AOI22_X1 U18659 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15615) );
  OAI21_X1 U18660 ( .B1(n15694), .B2(n17184), .A(n15615), .ZN(n15621) );
  AOI22_X1 U18661 ( .A1(n17080), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15619) );
  AOI22_X1 U18662 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9735), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15618) );
  AOI22_X1 U18663 ( .A1(n17165), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15617) );
  AOI22_X1 U18664 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n15672), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15616) );
  NAND4_X1 U18665 ( .A1(n15619), .A2(n15618), .A3(n15617), .A4(n15616), .ZN(
        n15620) );
  AOI211_X1 U18666 ( .C1(n17148), .C2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n15621), .B(n15620), .ZN(n15622) );
  NAND3_X1 U18667 ( .A1(n15624), .A2(n15623), .A3(n15622), .ZN(n16403) );
  AOI22_X1 U18668 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15628) );
  AOI22_X1 U18669 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15627) );
  AOI22_X1 U18670 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15626) );
  AOI22_X1 U18671 ( .A1(n9735), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15625) );
  NAND4_X1 U18672 ( .A1(n15628), .A2(n15627), .A3(n15626), .A4(n15625), .ZN(
        n15634) );
  AOI22_X1 U18673 ( .A1(n17170), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15632) );
  AOI22_X1 U18674 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15672), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15631) );
  AOI22_X1 U18675 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15630) );
  AOI22_X1 U18676 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15629) );
  NAND4_X1 U18677 ( .A1(n15632), .A2(n15631), .A3(n15630), .A4(n15629), .ZN(
        n15633) );
  AOI22_X1 U18678 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15638) );
  AOI22_X1 U18679 ( .A1(n17170), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n15672), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15637) );
  AOI22_X1 U18680 ( .A1(n15645), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15636) );
  AOI22_X1 U18681 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15635) );
  NAND4_X1 U18682 ( .A1(n15638), .A2(n15637), .A3(n15636), .A4(n15635), .ZN(
        n15644) );
  AOI22_X1 U18683 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9735), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15642) );
  AOI22_X1 U18684 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15641) );
  AOI22_X1 U18685 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15640) );
  AOI22_X1 U18686 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15639) );
  NAND4_X1 U18687 ( .A1(n15642), .A2(n15641), .A3(n15640), .A4(n15639), .ZN(
        n15643) );
  AOI22_X1 U18688 ( .A1(n15484), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n15670), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15657) );
  AOI22_X1 U18689 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n15672), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15656) );
  AOI22_X1 U18690 ( .A1(n15378), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15645), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15646) );
  OAI21_X1 U18691 ( .B1(n17008), .B2(n21063), .A(n15646), .ZN(n15654) );
  AOI22_X1 U18692 ( .A1(n17170), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15652) );
  AOI22_X1 U18693 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n15379), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15651) );
  AOI22_X1 U18694 ( .A1(n15533), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n15647), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15650) );
  AOI22_X1 U18695 ( .A1(n9735), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n15648), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15649) );
  NAND4_X1 U18696 ( .A1(n15652), .A2(n15651), .A3(n15650), .A4(n15649), .ZN(
        n15653) );
  NAND3_X1 U18697 ( .A1(n15657), .A2(n15656), .A3(n15655), .ZN(n15736) );
  AOI22_X1 U18698 ( .A1(n17170), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15661) );
  AOI22_X1 U18699 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15660) );
  AOI22_X1 U18700 ( .A1(n15645), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15659) );
  AOI22_X1 U18701 ( .A1(n9735), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15658) );
  NAND4_X1 U18702 ( .A1(n15661), .A2(n15660), .A3(n15659), .A4(n15658), .ZN(
        n15667) );
  AOI22_X1 U18703 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15665) );
  AOI22_X1 U18704 ( .A1(n17080), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15664) );
  AOI22_X1 U18705 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15663) );
  AOI22_X1 U18706 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15662) );
  NAND4_X1 U18707 ( .A1(n15665), .A2(n15664), .A3(n15663), .A4(n15662), .ZN(
        n15666) );
  NOR2_X1 U18708 ( .A1(n15667), .A2(n15666), .ZN(n17855) );
  AOI22_X1 U18709 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15681) );
  AOI22_X1 U18710 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15680) );
  INV_X1 U18711 ( .A(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n20967) );
  AOI22_X1 U18712 ( .A1(n17080), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15668) );
  OAI21_X1 U18713 ( .B1(n15669), .B2(n20967), .A(n15668), .ZN(n15678) );
  AOI22_X1 U18714 ( .A1(n15647), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15670), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15676) );
  AOI22_X1 U18715 ( .A1(n15671), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15533), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15675) );
  AOI22_X1 U18716 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9735), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15674) );
  AOI22_X1 U18717 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15672), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15673) );
  NAND4_X1 U18718 ( .A1(n15676), .A2(n15675), .A3(n15674), .A4(n15673), .ZN(
        n15677) );
  AOI211_X1 U18719 ( .C1(n17148), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n15678), .B(n15677), .ZN(n15679) );
  NAND3_X1 U18720 ( .A1(n15681), .A2(n15680), .A3(n15679), .ZN(n17363) );
  NOR2_X1 U18721 ( .A1(n15710), .A2(n17363), .ZN(n15708) );
  NOR2_X1 U18722 ( .A1(n17358), .A2(n15708), .ZN(n15706) );
  AOI22_X1 U18723 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15692) );
  AOI22_X1 U18724 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15691) );
  INV_X1 U18725 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n21166) );
  AOI22_X1 U18726 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15683) );
  OAI21_X1 U18727 ( .B1(n17169), .B2(n21166), .A(n15683), .ZN(n15689) );
  AOI22_X1 U18728 ( .A1(n15645), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9735), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15687) );
  AOI22_X1 U18729 ( .A1(n17170), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15686) );
  AOI22_X1 U18730 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15685) );
  AOI22_X1 U18731 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15684) );
  NAND4_X1 U18732 ( .A1(n15687), .A2(n15686), .A3(n15685), .A4(n15684), .ZN(
        n15688) );
  AOI211_X1 U18733 ( .C1(n17146), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n15689), .B(n15688), .ZN(n15690) );
  NAND3_X1 U18734 ( .A1(n15692), .A2(n15691), .A3(n15690), .ZN(n17353) );
  NAND2_X1 U18735 ( .A1(n15706), .A2(n17353), .ZN(n15705) );
  NOR2_X1 U18736 ( .A1(n17350), .A2(n15705), .ZN(n15718) );
  AOI22_X1 U18737 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15703) );
  AOI22_X1 U18738 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n15702) );
  AOI22_X1 U18739 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n15693) );
  OAI21_X1 U18740 ( .B1(n15694), .B2(n17191), .A(n15693), .ZN(n15700) );
  AOI22_X1 U18741 ( .A1(n9735), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n15698) );
  AOI22_X1 U18742 ( .A1(n17170), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n15697) );
  AOI22_X1 U18743 ( .A1(n17080), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15696) );
  AOI22_X1 U18744 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15695) );
  NAND4_X1 U18745 ( .A1(n15698), .A2(n15697), .A3(n15696), .A4(n15695), .ZN(
        n15699) );
  AOI211_X1 U18746 ( .C1(n17156), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n15700), .B(n15699), .ZN(n15701) );
  NAND3_X1 U18747 ( .A1(n15703), .A2(n15702), .A3(n15701), .ZN(n17345) );
  NAND2_X1 U18748 ( .A1(n15718), .A2(n17345), .ZN(n15704) );
  NOR2_X1 U18749 ( .A1(n17342), .A2(n15704), .ZN(n15726) );
  XOR2_X1 U18750 ( .A(n17342), .B(n15704), .Z(n17779) );
  INV_X1 U18751 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18113) );
  XOR2_X1 U18752 ( .A(n17350), .B(n15705), .Z(n17798) );
  XOR2_X1 U18753 ( .A(n17353), .B(n15706), .Z(n15707) );
  NAND2_X1 U18754 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15707), .ZN(
        n15716) );
  XOR2_X1 U18755 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n15707), .Z(
        n17813) );
  XOR2_X1 U18756 ( .A(n17358), .B(n15708), .Z(n15709) );
  NAND2_X1 U18757 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15709), .ZN(
        n15715) );
  XOR2_X1 U18758 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n15709), .Z(
        n17827) );
  INV_X1 U18759 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21167) );
  XOR2_X1 U18760 ( .A(n17363), .B(n15710), .Z(n15713) );
  OR2_X1 U18761 ( .A1(n21167), .A2(n15713), .ZN(n15714) );
  INV_X1 U18762 ( .A(n17855), .ZN(n15848) );
  AOI21_X1 U18763 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n9724), .A(
        n15848), .ZN(n15712) );
  INV_X1 U18764 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18796) );
  NOR2_X1 U18765 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n9724), .ZN(
        n15711) );
  AOI221_X1 U18766 ( .B1(n15848), .B2(n9724), .C1(n15712), .C2(n18796), .A(
        n15711), .ZN(n17835) );
  XOR2_X1 U18767 ( .A(n21167), .B(n15713), .Z(n17834) );
  NAND2_X1 U18768 ( .A1(n17835), .A2(n17834), .ZN(n17833) );
  NAND2_X1 U18769 ( .A1(n15714), .A2(n17833), .ZN(n17826) );
  NAND2_X1 U18770 ( .A1(n17827), .A2(n17826), .ZN(n17825) );
  NAND2_X1 U18771 ( .A1(n15715), .A2(n17825), .ZN(n17812) );
  NAND2_X1 U18772 ( .A1(n17813), .A2(n17812), .ZN(n17811) );
  NAND2_X1 U18773 ( .A1(n15716), .A2(n17811), .ZN(n17799) );
  NAND2_X1 U18774 ( .A1(n17798), .A2(n17799), .ZN(n17797) );
  NOR2_X1 U18775 ( .A1(n17798), .A2(n17799), .ZN(n15717) );
  AOI21_X1 U18776 ( .B1(n18113), .B2(n17797), .A(n15717), .ZN(n15719) );
  XOR2_X1 U18777 ( .A(n17345), .B(n15718), .Z(n15720) );
  NAND2_X1 U18778 ( .A1(n15719), .A2(n15720), .ZN(n15721) );
  XOR2_X1 U18779 ( .A(n15720), .B(n15719), .Z(n17792) );
  NAND2_X1 U18780 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17792), .ZN(
        n17791) );
  NAND2_X1 U18781 ( .A1(n15721), .A2(n17791), .ZN(n17778) );
  INV_X1 U18782 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18094) );
  NAND2_X1 U18783 ( .A1(n15726), .A2(n15722), .ZN(n15727) );
  INV_X1 U18784 ( .A(n15722), .ZN(n15725) );
  NAND2_X1 U18785 ( .A1(n17779), .A2(n17778), .ZN(n15724) );
  NAND2_X1 U18786 ( .A1(n15726), .A2(n15725), .ZN(n15723) );
  OAI211_X1 U18787 ( .C1(n15726), .C2(n15725), .A(n15724), .B(n15723), .ZN(
        n17763) );
  NAND2_X1 U18788 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17763), .ZN(
        n17762) );
  NOR2_X1 U18789 ( .A1(n17992), .A2(n17970), .ZN(n17628) );
  NAND2_X1 U18790 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17628), .ZN(
        n17941) );
  INV_X1 U18791 ( .A(n17941), .ZN(n17919) );
  INV_X1 U18792 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17926) );
  NOR2_X1 U18793 ( .A1(n17964), .A2(n17926), .ZN(n17938) );
  NAND2_X1 U18794 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17938), .ZN(
        n17921) );
  INV_X1 U18795 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17920) );
  NOR2_X1 U18796 ( .A1(n17921), .A2(n17920), .ZN(n15769) );
  NAND2_X1 U18797 ( .A1(n17919), .A2(n15769), .ZN(n17911) );
  INV_X1 U18798 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17901) );
  INV_X1 U18799 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17904) );
  NOR3_X1 U18800 ( .A1(n17911), .A2(n17901), .A3(n17904), .ZN(n17885) );
  NAND2_X1 U18801 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17885), .ZN(
        n17517) );
  NOR2_X1 U18802 ( .A1(n18000), .A2(n17517), .ZN(n17540) );
  NAND2_X1 U18803 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17540), .ZN(
        n17868) );
  INV_X1 U18804 ( .A(n17517), .ZN(n16399) );
  NAND2_X1 U18805 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18154), .ZN(
        n17878) );
  INV_X1 U18806 ( .A(n17878), .ZN(n15730) );
  AOI21_X1 U18807 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18144) );
  INV_X1 U18808 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18136) );
  NAND2_X1 U18809 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18087) );
  NOR2_X1 U18810 ( .A1(n18136), .A2(n18087), .ZN(n17971) );
  INV_X1 U18811 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18104) );
  NOR2_X1 U18812 ( .A1(n18104), .A2(n18094), .ZN(n18088) );
  NAND2_X1 U18813 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18088), .ZN(
        n17972) );
  INV_X1 U18814 ( .A(n17972), .ZN(n15728) );
  NAND2_X1 U18815 ( .A1(n17971), .A2(n15728), .ZN(n15729) );
  NOR2_X1 U18816 ( .A1(n18144), .A2(n15729), .ZN(n17987) );
  NAND2_X1 U18817 ( .A1(n15760), .A2(n17987), .ZN(n17966) );
  NAND2_X1 U18818 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18083) );
  NOR2_X1 U18819 ( .A1(n15729), .A2(n18083), .ZN(n18013) );
  NAND2_X1 U18820 ( .A1(n15760), .A2(n18013), .ZN(n17965) );
  AOI21_X1 U18821 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18641), .A(
        n18628), .ZN(n18137) );
  OAI22_X1 U18822 ( .A1(n18659), .A2(n17966), .B1(n17965), .B2(n18137), .ZN(
        n17884) );
  NAND3_X1 U18823 ( .A1(n16399), .A2(n15730), .A3(n17884), .ZN(n16387) );
  INV_X1 U18824 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17896) );
  NAND2_X1 U18825 ( .A1(n9724), .A2(n17363), .ZN(n15739) );
  NAND2_X1 U18826 ( .A1(n15734), .A2(n17353), .ZN(n15733) );
  XOR2_X1 U18827 ( .A(n15731), .B(n17345), .Z(n15732) );
  NAND2_X1 U18828 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15732), .ZN(
        n15747) );
  XOR2_X1 U18829 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n15732), .Z(
        n17786) );
  XOR2_X1 U18830 ( .A(n15733), .B(n17350), .Z(n15743) );
  XOR2_X1 U18831 ( .A(n15734), .B(n17353), .Z(n15741) );
  XOR2_X1 U18832 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n15741), .Z(
        n17815) );
  NAND2_X1 U18833 ( .A1(n17375), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15735) );
  NOR2_X1 U18834 ( .A1(n17855), .A2(n18796), .ZN(n17854) );
  XNOR2_X1 U18835 ( .A(n9724), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17846) );
  NAND2_X1 U18836 ( .A1(n17854), .A2(n17846), .ZN(n17845) );
  NAND2_X1 U18837 ( .A1(n15735), .A2(n17845), .ZN(n17837) );
  XNOR2_X1 U18838 ( .A(n17363), .B(n9724), .ZN(n15737) );
  NAND2_X1 U18839 ( .A1(n17837), .A2(n17838), .ZN(n17836) );
  OR2_X1 U18840 ( .A1(n21167), .A2(n15737), .ZN(n15738) );
  XOR2_X1 U18841 ( .A(n15739), .B(n17358), .Z(n17823) );
  NAND2_X1 U18842 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15741), .ZN(
        n15742) );
  NAND2_X1 U18843 ( .A1(n15743), .A2(n15745), .ZN(n15746) );
  AOI21_X1 U18844 ( .B1(n17342), .B2(n15748), .A(n17761), .ZN(n15750) );
  NAND2_X1 U18845 ( .A1(n15750), .A2(n15749), .ZN(n15751) );
  INV_X1 U18846 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21143) );
  NOR2_X1 U18847 ( .A1(n17911), .A2(n17901), .ZN(n15764) );
  INV_X1 U18848 ( .A(n15764), .ZN(n17552) );
  NAND2_X1 U18849 ( .A1(n17898), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17539) );
  NOR2_X1 U18850 ( .A1(n17896), .A2(n17539), .ZN(n17538) );
  NAND2_X1 U18851 ( .A1(n17538), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17488) );
  INV_X1 U18852 ( .A(n17488), .ZN(n17870) );
  NAND2_X1 U18853 ( .A1(n15753), .A2(n15752), .ZN(n16339) );
  NOR2_X1 U18854 ( .A1(n16403), .A2(n16339), .ZN(n17999) );
  NAND2_X1 U18855 ( .A1(n18154), .A2(n17999), .ZN(n15757) );
  INV_X1 U18856 ( .A(n15757), .ZN(n18082) );
  NAND2_X1 U18857 ( .A1(n17870), .A2(n18082), .ZN(n15754) );
  OAI211_X1 U18858 ( .C1(n18130), .C2(n17868), .A(n16387), .B(n15754), .ZN(
        n15833) );
  NAND2_X1 U18859 ( .A1(n16367), .A2(n15833), .ZN(n15775) );
  INV_X1 U18860 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16369) );
  NOR2_X1 U18861 ( .A1(n18170), .A2(n9908), .ZN(n18117) );
  INV_X1 U18862 ( .A(n16367), .ZN(n16380) );
  NAND2_X1 U18863 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17866) );
  NOR2_X1 U18864 ( .A1(n17552), .A2(n17966), .ZN(n17903) );
  AOI21_X1 U18865 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17903), .A(
        n18659), .ZN(n17864) );
  NAND2_X1 U18866 ( .A1(n18057), .A2(n18643), .ZN(n18084) );
  INV_X1 U18867 ( .A(n18084), .ZN(n18139) );
  INV_X1 U18868 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17525) );
  NOR3_X1 U18869 ( .A1(n17525), .A2(n17517), .A3(n17965), .ZN(n15755) );
  NOR2_X1 U18870 ( .A1(n18057), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18141) );
  INV_X1 U18871 ( .A(n18141), .ZN(n18085) );
  OAI21_X1 U18872 ( .B1(n18139), .B2(n15755), .A(n18085), .ZN(n15756) );
  AOI211_X1 U18873 ( .C1(n18639), .C2(n17866), .A(n17864), .B(n15756), .ZN(
        n16405) );
  NOR2_X1 U18874 ( .A1(n16405), .A2(n18170), .ZN(n15830) );
  OR3_X2 U18875 ( .A1(n18845), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18169) );
  NAND2_X1 U18876 ( .A1(n16367), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16388) );
  NOR2_X1 U18877 ( .A1(n16388), .A2(n17868), .ZN(n16381) );
  NOR2_X1 U18878 ( .A1(n17488), .A2(n16388), .ZN(n16368) );
  OAI22_X1 U18879 ( .A1(n16381), .A2(n18130), .B1(n16368), .B2(n15757), .ZN(
        n15758) );
  NOR2_X1 U18880 ( .A1(n18149), .A2(n15758), .ZN(n15831) );
  INV_X1 U18881 ( .A(n15831), .ZN(n15759) );
  AOI211_X1 U18882 ( .C1(n18117), .C2(n16380), .A(n15830), .B(n15759), .ZN(
        n15774) );
  INV_X1 U18883 ( .A(n16339), .ZN(n18656) );
  NOR4_X1 U18884 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15763) );
  INV_X1 U18885 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18069) );
  INV_X1 U18886 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18062) );
  NAND2_X1 U18887 ( .A1(n18069), .A2(n18062), .ZN(n17739) );
  INV_X1 U18888 ( .A(n17739), .ZN(n15762) );
  INV_X1 U18889 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18026) );
  NAND2_X1 U18890 ( .A1(n17598), .A2(n17665), .ZN(n17694) );
  NOR2_X1 U18891 ( .A1(n17761), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17634) );
  NAND2_X1 U18892 ( .A1(n17634), .A2(n17964), .ZN(n15765) );
  NOR2_X1 U18893 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15765), .ZN(
        n17600) );
  INV_X1 U18894 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17927) );
  NAND2_X1 U18895 ( .A1(n17600), .A2(n17927), .ZN(n17575) );
  NAND2_X1 U18896 ( .A1(n17628), .A2(n15768), .ZN(n17597) );
  NAND2_X1 U18897 ( .A1(n17605), .A2(n17597), .ZN(n17599) );
  NAND3_X1 U18898 ( .A1(n15769), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17599), .ZN(n17558) );
  NAND2_X1 U18899 ( .A1(n17504), .A2(n17490), .ZN(n15827) );
  NOR2_X1 U18900 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17598), .ZN(
        n16400) );
  AOI21_X1 U18901 ( .B1(n15828), .B2(n15827), .A(n16400), .ZN(n15771) );
  XNOR2_X1 U18902 ( .A(n15771), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16385) );
  INV_X1 U18903 ( .A(n16385), .ZN(n15772) );
  AOI22_X1 U18904 ( .A1(n9736), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n18073), 
        .B2(n15772), .ZN(n15773) );
  OAI221_X1 U18905 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15775), 
        .C1(n16369), .C2(n15774), .A(n15773), .ZN(P3_U2833) );
  OAI22_X1 U18906 ( .A1(n16148), .A2(n19034), .B1(n19029), .B2(n16121), .ZN(
        n15776) );
  INV_X1 U18907 ( .A(n15776), .ZN(n15785) );
  AOI211_X1 U18908 ( .C1(n15779), .C2(n15778), .A(n15777), .B(n19820), .ZN(
        n15783) );
  AOI22_X1 U18909 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18996), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19025), .ZN(n15780) );
  OAI21_X1 U18910 ( .B1(n15781), .B2(n19018), .A(n15780), .ZN(n15782) );
  AOI211_X1 U18911 ( .C1(n19026), .C2(P2_EBX_REG_22__SCAN_IN), .A(n15783), .B(
        n15782), .ZN(n15784) );
  NAND2_X1 U18912 ( .A1(n15785), .A2(n15784), .ZN(P2_U2833) );
  INV_X1 U18913 ( .A(n15786), .ZN(n15798) );
  AOI21_X1 U18914 ( .B1(n15787), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n20602), .ZN(n15788) );
  AND2_X1 U18915 ( .A1(n15789), .A2(n15788), .ZN(n15794) );
  INV_X1 U18916 ( .A(n15794), .ZN(n15796) );
  INV_X1 U18917 ( .A(n15790), .ZN(n15793) );
  INV_X1 U18918 ( .A(n15791), .ZN(n15792) );
  OAI22_X1 U18919 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n15794), .B1(
        n15793), .B2(n15792), .ZN(n15795) );
  OAI21_X1 U18920 ( .B1(n15796), .B2(n20492), .A(n15795), .ZN(n15797) );
  AOI222_X1 U18921 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n15798), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15797), .C1(n15798), 
        .C2(n15797), .ZN(n15799) );
  OR2_X1 U18922 ( .A1(n15800), .A2(n15799), .ZN(n15801) );
  AOI22_X1 U18923 ( .A1(n15801), .A2(n20565), .B1(n15800), .B2(n15799), .ZN(
        n15808) );
  INV_X1 U18924 ( .A(n15802), .ZN(n15803) );
  NOR2_X1 U18925 ( .A1(n15804), .A2(n15803), .ZN(n15807) );
  OAI21_X1 U18926 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15805), .ZN(n15806) );
  OAI211_X1 U18927 ( .C1(n15808), .C2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n15807), .B(n15806), .ZN(n15809) );
  NOR3_X1 U18928 ( .A1(n15811), .A2(n15810), .A3(n15809), .ZN(n15821) );
  INV_X1 U18929 ( .A(n15821), .ZN(n15816) );
  NOR3_X1 U18930 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n11307), .A3(n20856), 
        .ZN(n15814) );
  OAI22_X1 U18931 ( .A1(n15815), .A2(n15814), .B1(n15813), .B2(n15812), .ZN(
        n16046) );
  AOI221_X1 U18932 ( .B1(n20773), .B2(n20772), .C1(n15816), .C2(n20772), .A(
        n16046), .ZN(n16051) );
  AOI21_X1 U18933 ( .B1(n20783), .B2(n11307), .A(n15817), .ZN(n15819) );
  OAI211_X1 U18934 ( .C1(n15821), .C2(n15820), .A(n15819), .B(n15818), .ZN(
        n15822) );
  NOR2_X1 U18935 ( .A1(n16051), .A2(n15822), .ZN(n15826) );
  NAND2_X1 U18936 ( .A1(n20859), .A2(n15823), .ZN(n15824) );
  NAND2_X1 U18937 ( .A1(n20773), .A2(n15824), .ZN(n15825) );
  OAI22_X1 U18938 ( .A1(n15826), .A2(n20773), .B1(n16051), .B2(n15825), .ZN(
        P1_U3161) );
  OAI21_X1 U18939 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15829), .A(
        n16342), .ZN(n16366) );
  NOR2_X1 U18940 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16388), .ZN(
        n16362) );
  AOI21_X1 U18941 ( .B1(n18117), .B2(n16388), .A(n15830), .ZN(n16386) );
  INV_X1 U18942 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16389) );
  AOI21_X1 U18943 ( .B1(n16386), .B2(n15831), .A(n16389), .ZN(n15832) );
  AOI21_X1 U18944 ( .B1(n16362), .B2(n15833), .A(n15832), .ZN(n15834) );
  NAND2_X1 U18945 ( .A1(n9736), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16358) );
  OAI211_X1 U18946 ( .C1(n18078), .C2(n16366), .A(n15834), .B(n16358), .ZN(
        P3_U2832) );
  INV_X1 U18947 ( .A(HOLD), .ZN(n20778) );
  NAND2_X1 U18948 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20794), .ZN(n20782) );
  AOI21_X1 U18949 ( .B1(n20783), .B2(P1_STATE_REG_1__SCAN_IN), .A(n15835), 
        .ZN(n15837) );
  OAI211_X1 U18950 ( .C1(n20794), .C2(n20778), .A(P1_STATE_REG_0__SCAN_IN), 
        .B(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n15836) );
  OAI211_X1 U18951 ( .C1(n20778), .C2(n20782), .A(n15837), .B(n15836), .ZN(
        P1_U3195) );
  AND2_X1 U18952 ( .A1(n20074), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR2_X1 U18953 ( .A1(n19834), .A2(n16324), .ZN(n19816) );
  NAND2_X1 U18954 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19816), .ZN(n15839) );
  AOI21_X1 U18955 ( .B1(n19916), .B2(n16324), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15838) );
  AOI21_X1 U18956 ( .B1(n15839), .B2(n15838), .A(n15843), .ZN(P2_U3178) );
  INV_X1 U18957 ( .A(n15840), .ZN(n19939) );
  AOI221_X1 U18958 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n15843), .C1(n19939), .C2(
        n15843), .A(n19753), .ZN(n19931) );
  INV_X1 U18959 ( .A(n19931), .ZN(n19932) );
  NOR2_X1 U18960 ( .A1(n15844), .A2(n19932), .ZN(P2_U3047) );
  NOR3_X1 U18961 ( .A1(n15845), .A2(n17377), .A3(n16523), .ZN(n15846) );
  NOR2_X1 U18962 ( .A1(n17263), .A2(n17368), .ZN(n17371) );
  INV_X1 U18963 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17448) );
  INV_X1 U18964 ( .A(n17368), .ZN(n15850) );
  AOI22_X1 U18965 ( .A1(n17369), .A2(BUF2_REG_0__SCAN_IN), .B1(n17335), .B2(
        n15848), .ZN(n15849) );
  OAI221_X1 U18966 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17340), .C1(n17448), 
        .C2(n15850), .A(n15849), .ZN(P3_U2735) );
  AOI22_X1 U18967 ( .A1(n20021), .A2(P1_EBX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20024), .ZN(n15858) );
  AOI21_X1 U18968 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(n15851), .A(
        P1_REIP_REG_20__SCAN_IN), .ZN(n15853) );
  OAI22_X1 U18969 ( .A1(n15854), .A2(n19996), .B1(n15853), .B2(n15852), .ZN(
        n15855) );
  AOI21_X1 U18970 ( .B1(n20025), .B2(n15856), .A(n15855), .ZN(n15857) );
  OAI211_X1 U18971 ( .C1(n15859), .C2(n20016), .A(n15858), .B(n15857), .ZN(
        P1_U2820) );
  AOI211_X1 U18972 ( .C1(n20024), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15860), .B(n20123), .ZN(n15863) );
  AOI22_X1 U18973 ( .A1(n15861), .A2(P1_REIP_REG_18__SCAN_IN), .B1(n20021), 
        .B2(P1_EBX_REG_18__SCAN_IN), .ZN(n15862) );
  OAI211_X1 U18974 ( .C1(n19978), .C2(n15864), .A(n15863), .B(n15862), .ZN(
        n15865) );
  AOI21_X1 U18975 ( .B1(n15866), .B2(n19980), .A(n15865), .ZN(n15867) );
  OAI21_X1 U18976 ( .B1(n15868), .B2(n20016), .A(n15867), .ZN(P1_U2822) );
  OAI22_X1 U18977 ( .A1(n20009), .A2(n21002), .B1(n20016), .B2(n15918), .ZN(
        n15869) );
  AOI211_X1 U18978 ( .C1(n20024), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n20123), .B(n15869), .ZN(n15879) );
  XNOR2_X1 U18979 ( .A(n15872), .B(n15871), .ZN(n15966) );
  AOI22_X1 U18980 ( .A1(n15915), .A2(n19980), .B1(n20025), .B2(n15966), .ZN(
        n15878) );
  OAI21_X1 U18981 ( .B1(n15874), .B2(n15873), .A(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n15877) );
  INV_X1 U18982 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20815) );
  NAND3_X1 U18983 ( .A1(n20005), .A2(n15875), .A3(n20815), .ZN(n15876) );
  NAND4_X1 U18984 ( .A1(n15879), .A2(n15878), .A3(n15877), .A4(n15876), .ZN(
        P1_U2824) );
  INV_X1 U18985 ( .A(n15880), .ZN(n15896) );
  AOI21_X1 U18986 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15896), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15888) );
  OAI21_X1 U18987 ( .B1(n20006), .B2(n15881), .A(n19990), .ZN(n15884) );
  NOR2_X1 U18988 ( .A1(n19978), .A2(n15882), .ZN(n15883) );
  AOI211_X1 U18989 ( .C1(P1_EBX_REG_12__SCAN_IN), .C2(n20021), .A(n15884), .B(
        n15883), .ZN(n15887) );
  INV_X1 U18990 ( .A(n15885), .ZN(n15930) );
  AOI22_X1 U18991 ( .A1(n15931), .A2(n20027), .B1(n19980), .B2(n15930), .ZN(
        n15886) );
  OAI211_X1 U18992 ( .C1(n15889), .C2(n15888), .A(n15887), .B(n15886), .ZN(
        P1_U2828) );
  INV_X1 U18993 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20808) );
  NAND2_X1 U18994 ( .A1(n15891), .A2(n15890), .ZN(n15892) );
  AND2_X1 U18995 ( .A1(n15893), .A2(n15892), .ZN(n16001) );
  AOI22_X1 U18996 ( .A1(n20025), .A2(n16001), .B1(n20021), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n15894) );
  OAI211_X1 U18997 ( .C1(n20006), .C2(n11444), .A(n15894), .B(n19990), .ZN(
        n15895) );
  AOI221_X1 U18998 ( .B1(n15897), .B2(P1_REIP_REG_11__SCAN_IN), .C1(n15896), 
        .C2(n20808), .A(n15895), .ZN(n15901) );
  XOR2_X1 U18999 ( .A(n15899), .B(n15898), .Z(n15942) );
  NAND2_X1 U19000 ( .A1(n19980), .A2(n15942), .ZN(n15900) );
  OAI211_X1 U19001 ( .C1(n20016), .C2(n15945), .A(n15901), .B(n15900), .ZN(
        P1_U2829) );
  AOI22_X1 U19002 ( .A1(n15915), .A2(n20037), .B1(n20036), .B2(n15966), .ZN(
        n15902) );
  OAI21_X1 U19003 ( .B1(n20040), .B2(n21002), .A(n15902), .ZN(P1_U2856) );
  AOI22_X1 U19004 ( .A1(n15942), .A2(n20037), .B1(n20036), .B2(n16001), .ZN(
        n15903) );
  OAI21_X1 U19005 ( .B1(n20040), .B2(n15904), .A(n15903), .ZN(P1_U2861) );
  INV_X1 U19006 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n21141) );
  AOI22_X1 U19007 ( .A1(n15942), .A2(n15906), .B1(n20086), .B2(n15905), .ZN(
        n15907) );
  OAI21_X1 U19008 ( .B1(n21141), .B2(n15908), .A(n15907), .ZN(P1_U2893) );
  AOI22_X1 U19009 ( .A1(n20111), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20123), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15917) );
  INV_X1 U19010 ( .A(n15909), .ZN(n15911) );
  OAI21_X1 U19011 ( .B1(n15912), .B2(n15911), .A(n15910), .ZN(n15914) );
  XNOR2_X1 U19012 ( .A(n15914), .B(n15913), .ZN(n15967) );
  AOI22_X1 U19013 ( .A1(n15967), .A2(n20118), .B1(n15915), .B2(n20117), .ZN(
        n15916) );
  OAI211_X1 U19014 ( .C1(n20122), .C2(n15918), .A(n15917), .B(n15916), .ZN(
        P1_U2983) );
  OAI21_X1 U19015 ( .B1(n10122), .B2(n15920), .A(n15919), .ZN(n15922) );
  NAND2_X1 U19016 ( .A1(n15922), .A2(n15921), .ZN(n15925) );
  XNOR2_X1 U19017 ( .A(n15923), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15924) );
  XNOR2_X1 U19018 ( .A(n15925), .B(n15924), .ZN(n15987) );
  AOI22_X1 U19019 ( .A1(n20111), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20123), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15929) );
  AOI22_X1 U19020 ( .A1(n15927), .A2(n20117), .B1(n15932), .B2(n15926), .ZN(
        n15928) );
  OAI211_X1 U19021 ( .C1(n15987), .C2(n19955), .A(n15929), .B(n15928), .ZN(
        P1_U2985) );
  AOI22_X1 U19022 ( .A1(n20111), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20123), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15934) );
  AOI22_X1 U19023 ( .A1(n15932), .A2(n15931), .B1(n20117), .B2(n15930), .ZN(
        n15933) );
  OAI211_X1 U19024 ( .C1(n15935), .C2(n19955), .A(n15934), .B(n15933), .ZN(
        P1_U2987) );
  AOI22_X1 U19025 ( .A1(n20111), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20123), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15944) );
  NOR2_X1 U19026 ( .A1(n14444), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15939) );
  NOR2_X1 U19027 ( .A1(n15936), .A2(n12514), .ZN(n15938) );
  MUX2_X1 U19028 ( .A(n15939), .B(n15938), .S(n15937), .Z(n15941) );
  XNOR2_X1 U19029 ( .A(n15941), .B(n15940), .ZN(n16003) );
  AOI22_X1 U19030 ( .A1(n20118), .A2(n16003), .B1(n20117), .B2(n15942), .ZN(
        n15943) );
  OAI211_X1 U19031 ( .C1(n20122), .C2(n15945), .A(n15944), .B(n15943), .ZN(
        P1_U2988) );
  AOI22_X1 U19032 ( .A1(n20111), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20123), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15951) );
  NAND2_X1 U19033 ( .A1(n15948), .A2(n15947), .ZN(n15949) );
  XNOR2_X1 U19034 ( .A(n15946), .B(n15949), .ZN(n16027) );
  AOI22_X1 U19035 ( .A1(n16027), .A2(n20118), .B1(n20117), .B2(n19981), .ZN(
        n15950) );
  OAI211_X1 U19036 ( .C1(n20122), .C2(n19986), .A(n15951), .B(n15950), .ZN(
        P1_U2992) );
  AOI22_X1 U19037 ( .A1(n20111), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20123), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15957) );
  OAI21_X1 U19038 ( .B1(n15954), .B2(n15953), .A(n15952), .ZN(n15955) );
  INV_X1 U19039 ( .A(n15955), .ZN(n16039) );
  AOI22_X1 U19040 ( .A1(n16039), .A2(n20118), .B1(n20117), .B2(n20038), .ZN(
        n15956) );
  OAI211_X1 U19041 ( .C1(n20122), .C2(n20017), .A(n15957), .B(n15956), .ZN(
        P1_U2994) );
  INV_X1 U19042 ( .A(n15958), .ZN(n15961) );
  INV_X1 U19043 ( .A(n15959), .ZN(n15960) );
  AOI22_X1 U19044 ( .A1(n15961), .A2(n20152), .B1(n20133), .B2(n15960), .ZN(
        n15965) );
  NOR3_X1 U19045 ( .A1(n21157), .A2(n15992), .A3(n15971), .ZN(n15963) );
  OAI221_X1 U19046 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n15963), 
        .C1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n15970), .A(n15962), .ZN(
        n15964) );
  OAI211_X1 U19047 ( .C1(n20814), .C2(n19990), .A(n15965), .B(n15964), .ZN(
        P1_U3014) );
  AOI22_X1 U19048 ( .A1(n15967), .A2(n20152), .B1(n20133), .B2(n15966), .ZN(
        n15975) );
  NAND2_X1 U19049 ( .A1(n20123), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n15974) );
  NAND2_X1 U19050 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15970), .ZN(
        n15968) );
  NOR2_X1 U19051 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n15968), .ZN(
        n15978) );
  OAI21_X1 U19052 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15969), .A(
        n16000), .ZN(n15980) );
  OAI21_X1 U19053 ( .B1(n15978), .B2(n15980), .A(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15973) );
  NAND4_X1 U19054 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n15971), .A4(n15970), .ZN(
        n15972) );
  NAND4_X1 U19055 ( .A1(n15975), .A2(n15974), .A3(n15973), .A4(n15972), .ZN(
        P1_U3015) );
  NOR2_X1 U19056 ( .A1(n19990), .A2(n15976), .ZN(n15977) );
  AOI211_X1 U19057 ( .C1(n20152), .C2(n15979), .A(n15978), .B(n15977), .ZN(
        n15983) );
  AOI22_X1 U19058 ( .A1(n15981), .A2(n20133), .B1(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15980), .ZN(n15982) );
  NAND2_X1 U19059 ( .A1(n15983), .A2(n15982), .ZN(P1_U3016) );
  NOR2_X1 U19060 ( .A1(n16007), .A2(n16015), .ZN(n16002) );
  NOR4_X1 U19061 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15940), .A3(
        n15984), .A4(n15999), .ZN(n15989) );
  OAI22_X1 U19062 ( .A1(n15987), .A2(n15986), .B1(n20149), .B2(n15985), .ZN(
        n15988) );
  AOI21_X1 U19063 ( .B1(n16002), .B2(n15989), .A(n15988), .ZN(n15991) );
  NAND2_X1 U19064 ( .A1(n20123), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n15990) );
  OAI211_X1 U19065 ( .C1(n16000), .C2(n15992), .A(n15991), .B(n15990), .ZN(
        P1_U3017) );
  AOI22_X1 U19066 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n20123), .B1(n15999), 
        .B2(n15993), .ZN(n15998) );
  INV_X1 U19067 ( .A(n15994), .ZN(n15996) );
  AOI22_X1 U19068 ( .A1(n15996), .A2(n20152), .B1(n20133), .B2(n15995), .ZN(
        n15997) );
  OAI211_X1 U19069 ( .C1(n16000), .C2(n15999), .A(n15998), .B(n15997), .ZN(
        P1_U3018) );
  AOI22_X1 U19070 ( .A1(n16001), .A2(n20133), .B1(n20123), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16005) );
  AOI22_X1 U19071 ( .A1(n16003), .A2(n20152), .B1(n16002), .B2(n15940), .ZN(
        n16004) );
  OAI211_X1 U19072 ( .C1(n16006), .C2(n15940), .A(n16005), .B(n16004), .ZN(
        P1_U3020) );
  OAI21_X1 U19073 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n16007), .ZN(n16014) );
  AOI21_X1 U19074 ( .B1(n16009), .B2(n20133), .A(n16008), .ZN(n16013) );
  AOI22_X1 U19075 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n16011), .B1(
        n20152), .B2(n16010), .ZN(n16012) );
  OAI211_X1 U19076 ( .C1(n16015), .C2(n16014), .A(n16013), .B(n16012), .ZN(
        P1_U3021) );
  AOI21_X1 U19077 ( .B1(n12481), .B2(n16017), .A(n16016), .ZN(n16029) );
  INV_X1 U19078 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16025) );
  INV_X1 U19079 ( .A(n16018), .ZN(n16023) );
  INV_X1 U19080 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16030) );
  NAND3_X1 U19081 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16019), .A3(
        n20127), .ZN(n16031) );
  AOI221_X1 U19082 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16025), .C2(n16030), .A(
        n16031), .ZN(n16022) );
  OAI22_X1 U19083 ( .A1(n16020), .A2(n20149), .B1(n20803), .B2(n19990), .ZN(
        n16021) );
  AOI211_X1 U19084 ( .C1(n16023), .C2(n20152), .A(n16022), .B(n16021), .ZN(
        n16024) );
  OAI21_X1 U19085 ( .B1(n16029), .B2(n16025), .A(n16024), .ZN(P1_U3023) );
  AOI222_X1 U19086 ( .A1(n16027), .A2(n20152), .B1(n20133), .B2(n16026), .C1(
        P1_REIP_REG_7__SCAN_IN), .C2(n20123), .ZN(n16028) );
  OAI221_X1 U19087 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16031), .C1(
        n16030), .C2(n16029), .A(n16028), .ZN(P1_U3024) );
  INV_X1 U19088 ( .A(n16032), .ZN(n16035) );
  AOI21_X1 U19089 ( .B1(n16035), .B2(n16034), .A(n16033), .ZN(n16037) );
  AOI22_X1 U19090 ( .A1(n20133), .A2(n9819), .B1(n20123), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n16041) );
  AOI22_X1 U19091 ( .A1(n16039), .A2(n20152), .B1(n20127), .B2(n16038), .ZN(
        n16040) );
  OAI211_X1 U19092 ( .C1(n16043), .C2(n16042), .A(n16041), .B(n16040), .ZN(
        P1_U3026) );
  NAND4_X1 U19093 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n11307), .A4(n20856), .ZN(n16044) );
  NAND2_X1 U19094 ( .A1(n16045), .A2(n16044), .ZN(n20774) );
  OAI21_X1 U19095 ( .B1(n16047), .B2(n20774), .A(n16046), .ZN(n16048) );
  OAI221_X1 U19096 ( .B1(n16049), .B2(n20573), .C1(n16049), .C2(n20856), .A(
        n16048), .ZN(n16050) );
  AOI221_X1 U19097 ( .B1(n16051), .B2(n20772), .C1(n20773), .C2(n20772), .A(
        n16050), .ZN(P1_U3162) );
  NOR2_X1 U19098 ( .A1(n16051), .A2(n20773), .ZN(n16053) );
  OAI21_X1 U19099 ( .B1(n16053), .B2(n20573), .A(n16052), .ZN(P1_U3466) );
  INV_X1 U19100 ( .A(n16054), .ZN(n16055) );
  AOI22_X1 U19101 ( .A1(n16055), .A2(n19032), .B1(P2_REIP_REG_31__SCAN_IN), 
        .B2(n19025), .ZN(n16062) );
  AOI22_X1 U19102 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n18996), .B1(
        P2_EBX_REG_31__SCAN_IN), .B2(n19026), .ZN(n16061) );
  INV_X1 U19103 ( .A(n16056), .ZN(n19045) );
  AOI22_X1 U19104 ( .A1(n16057), .A2(n19020), .B1(n19015), .B2(n19045), .ZN(
        n16060) );
  NAND4_X1 U19105 ( .A1(n19021), .A2(n16063), .A3(n16058), .A4(n19002), .ZN(
        n16059) );
  NAND4_X1 U19106 ( .A1(n16062), .A2(n16061), .A3(n16060), .A4(n16059), .ZN(
        P2_U2824) );
  AOI21_X1 U19107 ( .B1(n16065), .B2(n16064), .A(n16063), .ZN(n16072) );
  OAI22_X1 U19108 ( .A1(n19010), .A2(n19884), .B1(n19037), .B2(n10002), .ZN(
        n16068) );
  NOR2_X1 U19109 ( .A1(n16066), .A2(n19018), .ZN(n16067) );
  AOI211_X1 U19110 ( .C1(n19026), .C2(P2_EBX_REG_29__SCAN_IN), .A(n16068), .B(
        n16067), .ZN(n16069) );
  OAI21_X1 U19111 ( .B1(n16070), .B2(n19034), .A(n16069), .ZN(n16071) );
  AOI21_X1 U19112 ( .B1(n19021), .B2(n16072), .A(n16071), .ZN(n16073) );
  OAI21_X1 U19113 ( .B1(n16074), .B2(n19029), .A(n16073), .ZN(P2_U2826) );
  AOI21_X1 U19114 ( .B1(n16077), .B2(n16076), .A(n16075), .ZN(n16087) );
  OAI22_X1 U19115 ( .A1(n19010), .A2(n19881), .B1(n19037), .B2(n16078), .ZN(
        n16079) );
  AOI21_X1 U19116 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n19026), .A(n16079), .ZN(
        n16084) );
  OAI211_X1 U19117 ( .C1(n16082), .C2(n16081), .A(n16080), .B(n19032), .ZN(
        n16083) );
  OAI211_X1 U19118 ( .C1(n16085), .C2(n19034), .A(n16084), .B(n16083), .ZN(
        n16086) );
  AOI21_X1 U19119 ( .B1(n19021), .B2(n16087), .A(n16086), .ZN(n16088) );
  OAI21_X1 U19120 ( .B1(n16089), .B2(n19029), .A(n16088), .ZN(P2_U2828) );
  AOI211_X1 U19121 ( .C1(n16092), .C2(n16091), .A(n16090), .B(n19820), .ZN(
        n16103) );
  INV_X1 U19122 ( .A(n16093), .ZN(n16101) );
  INV_X1 U19123 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n16095) );
  INV_X1 U19124 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16094) );
  OAI22_X1 U19125 ( .A1(n19010), .A2(n16095), .B1(n19037), .B2(n16094), .ZN(
        n16099) );
  AOI211_X1 U19126 ( .C1(P2_EBX_REG_26__SCAN_IN), .C2(n16097), .A(n19018), .B(
        n16096), .ZN(n16098) );
  AOI211_X1 U19127 ( .C1(n19026), .C2(P2_EBX_REG_26__SCAN_IN), .A(n16099), .B(
        n16098), .ZN(n16100) );
  OAI21_X1 U19128 ( .B1(n16101), .B2(n19034), .A(n16100), .ZN(n16102) );
  AOI211_X1 U19129 ( .C1(n19015), .C2(n16104), .A(n16103), .B(n16102), .ZN(
        n16105) );
  INV_X1 U19130 ( .A(n16105), .ZN(P2_U2829) );
  OAI22_X1 U19131 ( .A1(n16107), .A2(n19018), .B1(n16106), .B2(n19010), .ZN(
        n16108) );
  INV_X1 U19132 ( .A(n16108), .ZN(n16119) );
  AOI22_X1 U19133 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n19026), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n18996), .ZN(n16118) );
  OAI22_X1 U19134 ( .A1(n16110), .A2(n19034), .B1(n19029), .B2(n16109), .ZN(
        n16111) );
  INV_X1 U19135 ( .A(n16111), .ZN(n16117) );
  AOI21_X1 U19136 ( .B1(n16114), .B2(n16113), .A(n16112), .ZN(n16115) );
  NAND2_X1 U19137 ( .A1(n19021), .A2(n16115), .ZN(n16116) );
  NAND4_X1 U19138 ( .A1(n16119), .A2(n16118), .A3(n16117), .A4(n16116), .ZN(
        P2_U2831) );
  INV_X1 U19139 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n18213) );
  OAI22_X1 U19140 ( .A1(n19049), .A2(n19242), .B1(n14246), .B2(n19059), .ZN(
        n16120) );
  AOI21_X1 U19141 ( .B1(P2_EAX_REG_22__SCAN_IN), .B2(n19053), .A(n16120), .ZN(
        n16125) );
  INV_X1 U19142 ( .A(n16121), .ZN(n16122) );
  AOI22_X1 U19143 ( .A1(n16123), .A2(n19064), .B1(n19055), .B2(n16122), .ZN(
        n16124) );
  OAI211_X1 U19144 ( .C1(n19051), .C2(n18213), .A(n16125), .B(n16124), .ZN(
        P2_U2897) );
  INV_X1 U19145 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n17276) );
  OAI22_X1 U19146 ( .A1(n19051), .A2(n17276), .B1(n19049), .B2(n19232), .ZN(
        n16126) );
  AOI21_X1 U19147 ( .B1(P2_EAX_REG_20__SCAN_IN), .B2(n19053), .A(n16126), .ZN(
        n16130) );
  AOI22_X1 U19148 ( .A1(n16128), .A2(n19064), .B1(n19055), .B2(n16127), .ZN(
        n16129) );
  OAI211_X1 U19149 ( .C1(n19059), .C2(n14255), .A(n16130), .B(n16129), .ZN(
        P2_U2899) );
  INV_X1 U19150 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n18195) );
  OAI22_X1 U19151 ( .A1(n19051), .A2(n18195), .B1(n19049), .B2(n19222), .ZN(
        n16131) );
  AOI21_X1 U19152 ( .B1(P2_EAX_REG_18__SCAN_IN), .B2(n19053), .A(n16131), .ZN(
        n16137) );
  OAI22_X1 U19153 ( .A1(n16134), .A2(n16133), .B1(n16132), .B2(n18895), .ZN(
        n16135) );
  INV_X1 U19154 ( .A(n16135), .ZN(n16136) );
  OAI211_X1 U19155 ( .C1(n19059), .C2(n14264), .A(n16137), .B(n16136), .ZN(
        P2_U2901) );
  AOI22_X1 U19156 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19000), .B1(n16217), 
        .B2(n16138), .ZN(n16144) );
  OAI22_X1 U19157 ( .A1(n16140), .A2(n16219), .B1(n19159), .B2(n16139), .ZN(
        n16141) );
  AOI21_X1 U19158 ( .B1(n19156), .B2(n16142), .A(n16141), .ZN(n16143) );
  OAI211_X1 U19159 ( .C1(n16225), .C2(n9983), .A(n16144), .B(n16143), .ZN(
        P2_U2991) );
  AOI22_X1 U19160 ( .A1(n19154), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19000), .ZN(n16152) );
  NAND3_X1 U19161 ( .A1(n16146), .A2(n16145), .A3(n16186), .ZN(n16147) );
  OAI21_X1 U19162 ( .B1(n16211), .B2(n16148), .A(n16147), .ZN(n16149) );
  AOI21_X1 U19163 ( .B1(n16150), .B2(n19162), .A(n16149), .ZN(n16151) );
  OAI211_X1 U19164 ( .C1(n19152), .C2(n16153), .A(n16152), .B(n16151), .ZN(
        P2_U2992) );
  AOI22_X1 U19165 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n16243), .B1(n16217), 
        .B2(n18932), .ZN(n16158) );
  OAI22_X1 U19166 ( .A1(n16155), .A2(n19159), .B1(n16219), .B2(n16154), .ZN(
        n16156) );
  AOI21_X1 U19167 ( .B1(n19156), .B2(n18933), .A(n16156), .ZN(n16157) );
  OAI211_X1 U19168 ( .C1(n16225), .C2(n16159), .A(n16158), .B(n16157), .ZN(
        P2_U3001) );
  AOI22_X1 U19169 ( .A1(n19154), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19000), .ZN(n16166) );
  NOR3_X1 U19170 ( .A1(n16161), .A2(n16160), .A3(n19159), .ZN(n16164) );
  OAI22_X1 U19171 ( .A1(n16162), .A2(n16219), .B1(n16211), .B2(n18942), .ZN(
        n16163) );
  NOR2_X1 U19172 ( .A1(n16164), .A2(n16163), .ZN(n16165) );
  OAI211_X1 U19173 ( .C1(n19152), .C2(n18940), .A(n16166), .B(n16165), .ZN(
        P2_U3002) );
  AOI22_X1 U19174 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n16243), .B1(n16217), 
        .B2(n16167), .ZN(n16173) );
  OAI22_X1 U19175 ( .A1(n16169), .A2(n19159), .B1(n16168), .B2(n16219), .ZN(
        n16170) );
  AOI21_X1 U19176 ( .B1(n19156), .B2(n16171), .A(n16170), .ZN(n16172) );
  OAI211_X1 U19177 ( .C1(n16225), .C2(n16174), .A(n16173), .B(n16172), .ZN(
        P2_U3003) );
  AOI22_X1 U19178 ( .A1(n19154), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19000), .ZN(n16188) );
  AOI21_X1 U19179 ( .B1(n16177), .B2(n16176), .A(n16175), .ZN(n16232) );
  NOR2_X1 U19180 ( .A1(n16179), .A2(n16178), .ZN(n16183) );
  NAND2_X1 U19181 ( .A1(n16181), .A2(n16180), .ZN(n16182) );
  XNOR2_X1 U19182 ( .A(n16183), .B(n16182), .ZN(n16235) );
  OAI22_X1 U19183 ( .A1(n16235), .A2(n16219), .B1(n16211), .B2(n16184), .ZN(
        n16185) );
  AOI21_X1 U19184 ( .B1(n16232), .B2(n16186), .A(n16185), .ZN(n16187) );
  OAI211_X1 U19185 ( .C1(n19152), .C2(n18953), .A(n16188), .B(n16187), .ZN(
        P2_U3004) );
  AOI22_X1 U19186 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19000), .B1(n16217), 
        .B2(n18961), .ZN(n16194) );
  OAI22_X1 U19187 ( .A1(n16190), .A2(n19159), .B1(n16219), .B2(n16189), .ZN(
        n16191) );
  AOI21_X1 U19188 ( .B1(n19156), .B2(n16192), .A(n16191), .ZN(n16193) );
  OAI211_X1 U19189 ( .C1(n16225), .C2(n16195), .A(n16194), .B(n16193), .ZN(
        P2_U3005) );
  AOI22_X1 U19190 ( .A1(n19154), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19000), .ZN(n16208) );
  NOR2_X1 U19191 ( .A1(n16197), .A2(n16196), .ZN(n16202) );
  INV_X1 U19192 ( .A(n16198), .ZN(n16200) );
  NAND2_X1 U19193 ( .A1(n16200), .A2(n16199), .ZN(n16201) );
  XNOR2_X1 U19194 ( .A(n16202), .B(n16201), .ZN(n16240) );
  OAI21_X1 U19195 ( .B1(n16205), .B2(n16204), .A(n16203), .ZN(n16239) );
  OAI222_X1 U19196 ( .A1(n16241), .A2(n16211), .B1(n16219), .B2(n16240), .C1(
        n19159), .C2(n16239), .ZN(n16206) );
  INV_X1 U19197 ( .A(n16206), .ZN(n16207) );
  OAI211_X1 U19198 ( .C1(n19152), .C2(n16209), .A(n16208), .B(n16207), .ZN(
        P2_U3006) );
  AOI22_X1 U19199 ( .A1(n19154), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n19000), .ZN(n16216) );
  OAI22_X1 U19200 ( .A1(n16212), .A2(n19159), .B1(n16211), .B2(n16210), .ZN(
        n16213) );
  AOI21_X1 U19201 ( .B1(n19162), .B2(n16214), .A(n16213), .ZN(n16215) );
  OAI211_X1 U19202 ( .C1(n19152), .C2(n18989), .A(n16216), .B(n16215), .ZN(
        P2_U3008) );
  AOI22_X1 U19203 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19000), .B1(n16217), 
        .B2(n19004), .ZN(n16223) );
  OAI22_X1 U19204 ( .A1(n16220), .A2(n16219), .B1(n16218), .B2(n19159), .ZN(
        n16221) );
  AOI21_X1 U19205 ( .B1(n19156), .B2(n19005), .A(n16221), .ZN(n16222) );
  OAI211_X1 U19206 ( .C1(n16225), .C2(n16224), .A(n16223), .B(n16222), .ZN(
        P2_U3009) );
  INV_X1 U19207 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19858) );
  NOR2_X1 U19208 ( .A1(n19858), .A2(n16226), .ZN(n16229) );
  OAI22_X1 U19209 ( .A1(n16251), .A2(n18959), .B1(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16227), .ZN(n16228) );
  AOI211_X1 U19210 ( .C1(n16230), .C2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16229), .B(n16228), .ZN(n16234) );
  AOI22_X1 U19211 ( .A1(n16232), .A2(n16231), .B1(n19199), .B2(n18955), .ZN(
        n16233) );
  OAI211_X1 U19212 ( .C1(n16235), .C2(n19190), .A(n16234), .B(n16233), .ZN(
        P2_U3036) );
  INV_X1 U19213 ( .A(n16236), .ZN(n16237) );
  AOI22_X1 U19214 ( .A1(n16238), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19187), .B2(n16237), .ZN(n16250) );
  OAI222_X1 U19215 ( .A1(n16241), .A2(n16266), .B1(n19190), .B2(n16240), .C1(
        n19202), .C2(n16239), .ZN(n16242) );
  INV_X1 U19216 ( .A(n16242), .ZN(n16249) );
  NAND2_X1 U19217 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n16243), .ZN(n16248) );
  OAI221_X1 U19218 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16246), .C2(n16245), .A(
        n16244), .ZN(n16247) );
  NAND4_X1 U19219 ( .A1(n16250), .A2(n16249), .A3(n16248), .A4(n16247), .ZN(
        P2_U3038) );
  OAI22_X1 U19220 ( .A1(n16251), .A2(n19905), .B1(n13258), .B2(n18983), .ZN(
        n16254) );
  AOI211_X1 U19221 ( .C1(n19172), .C2(n16252), .A(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n19192), .ZN(n16253) );
  AOI211_X1 U19222 ( .C1(n19199), .C2(n16255), .A(n16254), .B(n16253), .ZN(
        n16256) );
  OAI21_X1 U19223 ( .B1(n16257), .B2(n19202), .A(n16256), .ZN(n16258) );
  AOI21_X1 U19224 ( .B1(n16259), .B2(n19182), .A(n16258), .ZN(n16260) );
  OAI21_X1 U19225 ( .B1(n16261), .B2(n21153), .A(n16260), .ZN(P2_U3043) );
  INV_X1 U19226 ( .A(n16262), .ZN(n19188) );
  AOI22_X1 U19227 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n19188), .B1(
        n19187), .B2(n16263), .ZN(n16274) );
  OAI21_X1 U19228 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19031), .A(
        n16264), .ZN(n16265) );
  INV_X1 U19229 ( .A(n16265), .ZN(n19161) );
  NAND2_X1 U19230 ( .A1(n19182), .A2(n19161), .ZN(n16272) );
  OR2_X1 U19231 ( .A1(n16266), .A2(n19035), .ZN(n16271) );
  OR2_X1 U19232 ( .A1(n18983), .A2(n18870), .ZN(n19157) );
  OR2_X1 U19233 ( .A1(n16267), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16268) );
  NAND2_X1 U19234 ( .A1(n16269), .A2(n16268), .ZN(n19158) );
  OR2_X1 U19235 ( .A1(n19202), .A2(n19158), .ZN(n16270) );
  AND4_X1 U19236 ( .A1(n16272), .A2(n16271), .A3(n19157), .A4(n16270), .ZN(
        n16273) );
  OAI211_X1 U19237 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n19192), .A(
        n16274), .B(n16273), .ZN(P2_U3046) );
  INV_X1 U19238 ( .A(n16308), .ZN(n16284) );
  NAND2_X1 U19239 ( .A1(n16277), .A2(n19924), .ZN(n16279) );
  INV_X1 U19240 ( .A(n16275), .ZN(n16276) );
  OAI22_X1 U19241 ( .A1(n16277), .A2(n19924), .B1(n19933), .B2(n16276), .ZN(
        n16278) );
  NAND2_X1 U19242 ( .A1(n16279), .A2(n16278), .ZN(n16280) );
  OAI211_X1 U19243 ( .C1(n19908), .C2(n16285), .A(n16284), .B(n16280), .ZN(
        n16283) );
  NAND2_X1 U19244 ( .A1(n16283), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n16282) );
  MUX2_X1 U19245 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n16281), .S(
        n16284), .Z(n16290) );
  NAND3_X1 U19246 ( .A1(n16282), .A2(n16290), .A3(n19908), .ZN(n16288) );
  OR2_X1 U19247 ( .A1(n16283), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n16287) );
  MUX2_X1 U19248 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16285), .S(
        n16284), .Z(n16289) );
  NAND2_X1 U19249 ( .A1(n16289), .A2(n19908), .ZN(n16286) );
  NAND3_X1 U19250 ( .A1(n16288), .A2(n16287), .A3(n16286), .ZN(n16313) );
  INV_X1 U19251 ( .A(n16289), .ZN(n16311) );
  INV_X1 U19252 ( .A(n16290), .ZN(n16310) );
  AOI22_X1 U19253 ( .A1(n16294), .A2(n16293), .B1(n16292), .B2(n16291), .ZN(
        n16298) );
  NAND2_X1 U19254 ( .A1(n16296), .A2(n16295), .ZN(n16297) );
  AND2_X1 U19255 ( .A1(n16298), .A2(n16297), .ZN(n19941) );
  NAND2_X1 U19256 ( .A1(n16316), .A2(n16299), .ZN(n16301) );
  OAI22_X1 U19257 ( .A1(n16302), .A2(n16301), .B1(n10721), .B2(n16300), .ZN(
        n16303) );
  INV_X1 U19258 ( .A(n16303), .ZN(n16306) );
  OAI21_X1 U19259 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n16304), .ZN(n16305) );
  NAND3_X1 U19260 ( .A1(n19941), .A2(n16306), .A3(n16305), .ZN(n16307) );
  AOI21_X1 U19261 ( .B1(n16308), .B2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n16307), .ZN(n16309) );
  OAI21_X1 U19262 ( .B1(n16311), .B2(n16310), .A(n16309), .ZN(n16312) );
  AOI21_X1 U19263 ( .B1(n16313), .B2(n15844), .A(n16312), .ZN(n16334) );
  NOR2_X1 U19264 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n16324), .ZN(n19818) );
  NAND2_X1 U19265 ( .A1(n16334), .A2(n21119), .ZN(n16314) );
  NAND2_X1 U19266 ( .A1(n16314), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n16322) );
  NAND2_X1 U19267 ( .A1(n10412), .A2(n16315), .ZN(n16318) );
  OAI21_X1 U19268 ( .B1(n16319), .B2(n16318), .A(n16317), .ZN(n16320) );
  INV_X1 U19269 ( .A(n16320), .ZN(n16321) );
  AND2_X1 U19270 ( .A1(n16322), .A2(n16321), .ZN(n19822) );
  NAND2_X1 U19271 ( .A1(n16323), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19926) );
  AOI21_X1 U19272 ( .B1(n16336), .B2(n19926), .A(n16324), .ZN(n16326) );
  AOI211_X1 U19273 ( .C1(n19834), .C2(n19818), .A(n16326), .B(n16325), .ZN(
        n16332) );
  NOR2_X1 U19274 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16327), .ZN(n16329) );
  OAI22_X1 U19275 ( .A1(n16330), .A2(n16329), .B1(n16328), .B2(n16336), .ZN(
        n16331) );
  OAI211_X1 U19276 ( .C1(n16334), .C2(n16333), .A(n16332), .B(n16331), .ZN(
        P2_U3176) );
  OAI221_X1 U19277 ( .B1(n19576), .B2(P2_STATE2_REG_0__SCAN_IN), .C1(n19576), 
        .C2(n16336), .A(n16335), .ZN(P2_U3593) );
  INV_X1 U19278 ( .A(n18654), .ZN(n16338) );
  NAND2_X1 U19279 ( .A1(n16338), .A2(n16337), .ZN(n18655) );
  NOR2_X1 U19280 ( .A1(n17761), .A2(n16341), .ZN(n16348) );
  NAND2_X1 U19281 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17761), .ZN(
        n16344) );
  OAI21_X1 U19282 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16389), .A(
        n16343), .ZN(n16346) );
  OAI22_X1 U19283 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17761), .B1(
        n16344), .B2(n16389), .ZN(n16345) );
  OAI21_X1 U19284 ( .B1(n16348), .B2(n16346), .A(n16345), .ZN(n16347) );
  INV_X1 U19285 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16544) );
  NAND2_X1 U19286 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17809) );
  NAND2_X1 U19287 ( .A1(n17806), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17787) );
  NAND2_X1 U19288 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17767) );
  INV_X1 U19289 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16774) );
  NAND2_X1 U19290 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17703) );
  NAND2_X1 U19291 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17656) );
  NAND2_X1 U19292 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17618) );
  NAND2_X1 U19293 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17584) );
  NAND2_X1 U19294 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17533) );
  INV_X1 U19295 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16370) );
  INV_X1 U19296 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18772) );
  NOR2_X1 U19297 ( .A1(n18772), .A2(n18169), .ZN(n16391) );
  INV_X1 U19298 ( .A(n17498), .ZN(n17485) );
  NAND3_X1 U19299 ( .A1(n17485), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16375) );
  NOR2_X1 U19300 ( .A1(n16370), .A2(n16375), .ZN(n16350) );
  NAND2_X1 U19301 ( .A1(n16516), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17856) );
  NAND2_X1 U19302 ( .A1(n16350), .A2(n17654), .ZN(n16360) );
  XNOR2_X1 U19303 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16351) );
  NOR2_X1 U19304 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17640), .ZN(
        n16372) );
  INV_X1 U19305 ( .A(n16371), .ZN(n16526) );
  OR2_X1 U19306 ( .A1(n18219), .A2(n16350), .ZN(n16376) );
  OAI211_X1 U19307 ( .C1(n16526), .C2(n17856), .A(n17857), .B(n16376), .ZN(
        n16379) );
  NOR2_X1 U19308 ( .A1(n16372), .A2(n16379), .ZN(n16359) );
  OAI22_X1 U19309 ( .A1(n16360), .A2(n16351), .B1(n16359), .B2(n16544), .ZN(
        n16352) );
  AOI211_X1 U19310 ( .C1(n17692), .C2(n16815), .A(n16391), .B(n16352), .ZN(
        n16357) );
  NAND2_X1 U19311 ( .A1(n17342), .A2(n16353), .ZN(n17579) );
  INV_X1 U19312 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18797) );
  NAND2_X1 U19313 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16368), .ZN(
        n16354) );
  XOR2_X1 U19314 ( .A(n18797), .B(n16354), .Z(n16394) );
  NOR2_X2 U19315 ( .A1(n16523), .A2(n16498), .ZN(n17848) );
  NAND2_X1 U19316 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16381), .ZN(
        n16355) );
  XOR2_X1 U19317 ( .A(n18797), .B(n16355), .Z(n16393) );
  AOI22_X1 U19318 ( .A1(n17766), .A2(n16394), .B1(n17848), .B2(n16393), .ZN(
        n16356) );
  OAI211_X1 U19319 ( .C1(n17764), .C2(n16397), .A(n16357), .B(n16356), .ZN(
        P3_U2799) );
  XNOR2_X1 U19320 ( .A(n9841), .B(n10020), .ZN(n16547) );
  OAI221_X1 U19321 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16360), .C1(
        n10020), .C2(n16359), .A(n16358), .ZN(n16361) );
  AOI21_X1 U19322 ( .B1(n17692), .B2(n16547), .A(n16361), .ZN(n16365) );
  OAI22_X1 U19323 ( .A1(n16368), .A2(n17579), .B1(n16381), .B2(n17861), .ZN(
        n16363) );
  INV_X1 U19324 ( .A(n17661), .ZN(n17590) );
  NOR3_X1 U19325 ( .A1(n17525), .A2(n17517), .A3(n17590), .ZN(n17512) );
  AOI22_X1 U19326 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16363), .B1(
        n16362), .B2(n17512), .ZN(n16364) );
  OAI211_X1 U19327 ( .C1(n17764), .C2(n16366), .A(n16365), .B(n16364), .ZN(
        P3_U2800) );
  NAND2_X1 U19328 ( .A1(n17870), .A2(n16367), .ZN(n16402) );
  AOI211_X1 U19329 ( .C1(n16369), .C2(n16402), .A(n16368), .B(n17579), .ZN(
        n16378) );
  NAND2_X1 U19330 ( .A1(n9736), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16374) );
  AOI21_X1 U19331 ( .B1(n16371), .B2(n16370), .A(n9841), .ZN(n16556) );
  OAI21_X1 U19332 ( .B1(n17692), .B2(n16372), .A(n16556), .ZN(n16373) );
  OAI211_X1 U19333 ( .C1(n16376), .C2(n16375), .A(n16374), .B(n16373), .ZN(
        n16377) );
  AOI211_X1 U19334 ( .C1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n16379), .A(
        n16378), .B(n16377), .ZN(n16384) );
  NOR2_X1 U19335 ( .A1(n16380), .A2(n17868), .ZN(n16407) );
  NOR2_X1 U19336 ( .A1(n16381), .A2(n17861), .ZN(n16382) );
  OAI21_X1 U19337 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16407), .A(
        n16382), .ZN(n16383) );
  OAI211_X1 U19338 ( .C1(n16385), .C2(n17764), .A(n16384), .B(n16383), .ZN(
        P3_U2801) );
  INV_X1 U19339 ( .A(n18117), .ZN(n18156) );
  OAI211_X1 U19340 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n18156), .A(
        n16386), .B(n18155), .ZN(n16392) );
  NOR4_X1 U19341 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16389), .A3(
        n16388), .A4(n16387), .ZN(n16390) );
  AOI211_X1 U19342 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16392), .A(
        n16391), .B(n16390), .ZN(n16396) );
  AOI22_X1 U19343 ( .A1(n16394), .A2(n18082), .B1(n16393), .B2(n18166), .ZN(
        n16395) );
  OAI211_X1 U19344 ( .C1(n16397), .C2(n18078), .A(n16396), .B(n16395), .ZN(
        P3_U2831) );
  INV_X1 U19345 ( .A(n17999), .ZN(n18028) );
  OAI22_X1 U19346 ( .A1(n18658), .A2(n18000), .B1(n17998), .B2(n18028), .ZN(
        n16398) );
  NOR2_X1 U19347 ( .A1(n17884), .A2(n16398), .ZN(n17912) );
  NOR2_X1 U19348 ( .A1(n17912), .A2(n18170), .ZN(n17918) );
  NAND2_X1 U19349 ( .A1(n16399), .A2(n17918), .ZN(n17877) );
  NOR2_X1 U19350 ( .A1(n17525), .A2(n17877), .ZN(n17873) );
  NOR2_X1 U19351 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17871), .ZN(
        n17497) );
  AOI22_X1 U19352 ( .A1(n9736), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n17873), 
        .B2(n17497), .ZN(n16416) );
  INV_X1 U19353 ( .A(n18162), .ZN(n18168) );
  AOI21_X1 U19354 ( .B1(n17761), .B2(n17505), .A(n17504), .ZN(n17494) );
  NAND3_X1 U19355 ( .A1(n18168), .A2(n16400), .A3(n17494), .ZN(n16415) );
  AOI22_X1 U19356 ( .A1(n17761), .A2(n17490), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17598), .ZN(n17493) );
  NAND3_X1 U19357 ( .A1(n17504), .A2(n18073), .A3(n17493), .ZN(n16414) );
  NOR2_X1 U19358 ( .A1(n16401), .A2(n17492), .ZN(n16404) );
  OAI221_X1 U19359 ( .B1(n17342), .B2(n16404), .C1(n16403), .C2(n16402), .A(
        n18656), .ZN(n16410) );
  OAI211_X1 U19360 ( .C1(n9908), .C2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16405), .B(n18155), .ZN(n16406) );
  OR2_X1 U19361 ( .A1(n16407), .A2(n18658), .ZN(n16408) );
  NAND3_X1 U19362 ( .A1(n16410), .A2(n16409), .A3(n16408), .ZN(n16412) );
  NAND4_X1 U19363 ( .A1(n16416), .A2(n16415), .A3(n16414), .A4(n16413), .ZN(
        P3_U2834) );
  NOR3_X1 U19364 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16418) );
  NOR4_X1 U19365 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16417) );
  NAND4_X1 U19366 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16418), .A3(n16417), .A4(
        U215), .ZN(U213) );
  INV_X2 U19367 ( .A(U214), .ZN(n16453) );
  NOR2_X1 U19368 ( .A1(n16453), .A2(n16419), .ZN(n16454) );
  AOI222_X1 U19369 ( .A1(n16453), .A2(P1_DATAO_REG_31__SCAN_IN), .B1(n16454), 
        .B2(BUF1_REG_31__SCAN_IN), .C1(n16449), .C2(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n16420) );
  INV_X1 U19370 ( .A(n16420), .ZN(U216) );
  INV_X1 U19371 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19080) );
  INV_X1 U19372 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n20043) );
  OAI222_X1 U19373 ( .A1(U212), .A2(n19080), .B1(n16451), .B2(n19241), .C1(
        U214), .C2(n20043), .ZN(U217) );
  AOI22_X1 U19374 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n16453), .ZN(n16421) );
  OAI21_X1 U19375 ( .B1(n14210), .B2(n16451), .A(n16421), .ZN(U218) );
  AOI22_X1 U19376 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n16453), .ZN(n16422) );
  OAI21_X1 U19377 ( .B1(n19231), .B2(n16451), .A(n16422), .ZN(U219) );
  AOI22_X1 U19378 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16453), .ZN(n16423) );
  OAI21_X1 U19379 ( .B1(n14225), .B2(n16451), .A(n16423), .ZN(U220) );
  AOI22_X1 U19380 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16453), .ZN(n16424) );
  OAI21_X1 U19381 ( .B1(n16425), .B2(n16451), .A(n16424), .ZN(U221) );
  AOI22_X1 U19382 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n16453), .ZN(n16426) );
  OAI21_X1 U19383 ( .B1(n14233), .B2(n16451), .A(n16426), .ZN(U222) );
  AOI22_X1 U19384 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n16453), .ZN(n16427) );
  OAI21_X1 U19385 ( .B1(n19207), .B2(n16451), .A(n16427), .ZN(U223) );
  AOI22_X1 U19386 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n16453), .ZN(n16428) );
  OAI21_X1 U19387 ( .B1(n14241), .B2(n16451), .A(n16428), .ZN(U224) );
  AOI22_X1 U19388 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n16453), .ZN(n16429) );
  OAI21_X1 U19389 ( .B1(n14246), .B2(n16451), .A(n16429), .ZN(U225) );
  AOI22_X1 U19390 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n16453), .ZN(n16430) );
  OAI21_X1 U19391 ( .B1(n14250), .B2(n16451), .A(n16430), .ZN(U226) );
  AOI22_X1 U19392 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16453), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16449), .ZN(n16431) );
  OAI21_X1 U19393 ( .B1(n14255), .B2(n16451), .A(n16431), .ZN(U227) );
  AOI22_X1 U19394 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n16453), .ZN(n16432) );
  OAI21_X1 U19395 ( .B1(n14259), .B2(n16451), .A(n16432), .ZN(U228) );
  AOI22_X1 U19396 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n16453), .ZN(n16433) );
  OAI21_X1 U19397 ( .B1(n14264), .B2(n16451), .A(n16433), .ZN(U229) );
  AOI22_X1 U19398 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n16453), .ZN(n16434) );
  OAI21_X1 U19399 ( .B1(n14268), .B2(n16451), .A(n16434), .ZN(U230) );
  AOI22_X1 U19400 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n16453), .ZN(n16435) );
  OAI21_X1 U19401 ( .B1(n14275), .B2(n16451), .A(n16435), .ZN(U231) );
  AOI22_X1 U19402 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16453), .ZN(n16436) );
  OAI21_X1 U19403 ( .B1(n12876), .B2(n16451), .A(n16436), .ZN(U232) );
  AOI22_X1 U19404 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16453), .ZN(n16437) );
  OAI21_X1 U19405 ( .B1(n14199), .B2(n16451), .A(n16437), .ZN(U233) );
  AOI22_X1 U19406 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16453), .ZN(n16438) );
  OAI21_X1 U19407 ( .B1(n14206), .B2(n16451), .A(n16438), .ZN(U234) );
  AOI22_X1 U19408 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16453), .ZN(n16439) );
  OAI21_X1 U19409 ( .B1(n14213), .B2(n16451), .A(n16439), .ZN(U235) );
  AOI22_X1 U19410 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16453), .ZN(n16440) );
  OAI21_X1 U19411 ( .B1(n14220), .B2(n16451), .A(n16440), .ZN(U236) );
  AOI22_X1 U19412 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16453), .ZN(n16441) );
  OAI21_X1 U19413 ( .B1(n13532), .B2(n16451), .A(n16441), .ZN(U237) );
  AOI22_X1 U19414 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16453), .ZN(n16442) );
  OAI21_X1 U19415 ( .B1(n13513), .B2(n16451), .A(n16442), .ZN(U238) );
  AOI22_X1 U19416 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16453), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16449), .ZN(n16443) );
  OAI21_X1 U19417 ( .B1(n13479), .B2(n16451), .A(n16443), .ZN(U239) );
  AOI22_X1 U19418 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16453), .ZN(n16444) );
  OAI21_X1 U19419 ( .B1(n13101), .B2(n16451), .A(n16444), .ZN(U240) );
  AOI22_X1 U19420 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16453), .ZN(n16445) );
  OAI21_X1 U19421 ( .B1(n13092), .B2(n16451), .A(n16445), .ZN(U241) );
  AOI22_X1 U19422 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16453), .ZN(n16446) );
  OAI21_X1 U19423 ( .B1(n13105), .B2(n16451), .A(n16446), .ZN(U242) );
  INV_X1 U19424 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16459) );
  AOI22_X1 U19425 ( .A1(BUF1_REG_4__SCAN_IN), .A2(n16454), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16453), .ZN(n16447) );
  OAI21_X1 U19426 ( .B1(n16459), .B2(U212), .A(n16447), .ZN(U243) );
  INV_X1 U19427 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n21089) );
  AOI22_X1 U19428 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16454), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16453), .ZN(n16448) );
  OAI21_X1 U19429 ( .B1(n21089), .B2(U212), .A(n16448), .ZN(U244) );
  AOI22_X1 U19430 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16453), .ZN(n16450) );
  OAI21_X1 U19431 ( .B1(n13131), .B2(n16451), .A(n16450), .ZN(U245) );
  INV_X1 U19432 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16457) );
  AOI22_X1 U19433 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16454), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16453), .ZN(n16452) );
  OAI21_X1 U19434 ( .B1(n16457), .B2(U212), .A(n16452), .ZN(U246) );
  INV_X1 U19435 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16456) );
  AOI22_X1 U19436 ( .A1(BUF1_REG_0__SCAN_IN), .A2(n16454), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16453), .ZN(n16455) );
  OAI21_X1 U19437 ( .B1(n16456), .B2(U212), .A(n16455), .ZN(U247) );
  INV_X1 U19438 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18184) );
  AOI22_X1 U19439 ( .A1(n16487), .A2(n16456), .B1(n18184), .B2(U215), .ZN(U251) );
  INV_X1 U19440 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18191) );
  AOI22_X1 U19441 ( .A1(n16487), .A2(n16457), .B1(n18191), .B2(U215), .ZN(U252) );
  OAI22_X1 U19442 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16484), .ZN(n16458) );
  INV_X1 U19443 ( .A(n16458), .ZN(U253) );
  INV_X1 U19444 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18201) );
  AOI22_X1 U19445 ( .A1(n16487), .A2(n21089), .B1(n18201), .B2(U215), .ZN(U254) );
  INV_X1 U19446 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18205) );
  AOI22_X1 U19447 ( .A1(n16487), .A2(n16459), .B1(n18205), .B2(U215), .ZN(U255) );
  OAI22_X1 U19448 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16487), .ZN(n16460) );
  INV_X1 U19449 ( .A(n16460), .ZN(U256) );
  OAI22_X1 U19450 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16487), .ZN(n16461) );
  INV_X1 U19451 ( .A(n16461), .ZN(U257) );
  OAI22_X1 U19452 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16484), .ZN(n16462) );
  INV_X1 U19453 ( .A(n16462), .ZN(U258) );
  OAI22_X1 U19454 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16487), .ZN(n16463) );
  INV_X1 U19455 ( .A(n16463), .ZN(U259) );
  OAI22_X1 U19456 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16487), .ZN(n16464) );
  INV_X1 U19457 ( .A(n16464), .ZN(U260) );
  OAI22_X1 U19458 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16487), .ZN(n16465) );
  INV_X1 U19459 ( .A(n16465), .ZN(U261) );
  OAI22_X1 U19460 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16487), .ZN(n16466) );
  INV_X1 U19461 ( .A(n16466), .ZN(U262) );
  OAI22_X1 U19462 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16487), .ZN(n16467) );
  INV_X1 U19463 ( .A(n16467), .ZN(U263) );
  OAI22_X1 U19464 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16487), .ZN(n16468) );
  INV_X1 U19465 ( .A(n16468), .ZN(U264) );
  OAI22_X1 U19466 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16487), .ZN(n16469) );
  INV_X1 U19467 ( .A(n16469), .ZN(U265) );
  OAI22_X1 U19468 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16487), .ZN(n16470) );
  INV_X1 U19469 ( .A(n16470), .ZN(U266) );
  OAI22_X1 U19470 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16487), .ZN(n16471) );
  INV_X1 U19471 ( .A(n16471), .ZN(U267) );
  OAI22_X1 U19472 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16484), .ZN(n16472) );
  INV_X1 U19473 ( .A(n16472), .ZN(U268) );
  OAI22_X1 U19474 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16487), .ZN(n16473) );
  INV_X1 U19475 ( .A(n16473), .ZN(U269) );
  OAI22_X1 U19476 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16484), .ZN(n16474) );
  INV_X1 U19477 ( .A(n16474), .ZN(U270) );
  OAI22_X1 U19478 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16487), .ZN(n16475) );
  INV_X1 U19479 ( .A(n16475), .ZN(U271) );
  OAI22_X1 U19480 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16484), .ZN(n16476) );
  INV_X1 U19481 ( .A(n16476), .ZN(U272) );
  OAI22_X1 U19482 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16487), .ZN(n16477) );
  INV_X1 U19483 ( .A(n16477), .ZN(U273) );
  INV_X1 U19484 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n16478) );
  INV_X1 U19485 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n19254) );
  AOI22_X1 U19486 ( .A1(n16487), .A2(n16478), .B1(n19254), .B2(U215), .ZN(U274) );
  OAI22_X1 U19487 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16487), .ZN(n16479) );
  INV_X1 U19488 ( .A(n16479), .ZN(U275) );
  OAI22_X1 U19489 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16484), .ZN(n16480) );
  INV_X1 U19490 ( .A(n16480), .ZN(U276) );
  OAI22_X1 U19491 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16484), .ZN(n16481) );
  INV_X1 U19492 ( .A(n16481), .ZN(U277) );
  OAI22_X1 U19493 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16484), .ZN(n16482) );
  INV_X1 U19494 ( .A(n16482), .ZN(U278) );
  OAI22_X1 U19495 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16484), .ZN(n16483) );
  INV_X1 U19496 ( .A(n16483), .ZN(U279) );
  OAI22_X1 U19497 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16484), .ZN(n16485) );
  INV_X1 U19498 ( .A(n16485), .ZN(U280) );
  AOI22_X1 U19499 ( .A1(n16487), .A2(n19080), .B1(n19240), .B2(U215), .ZN(U281) );
  INV_X1 U19500 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n21034) );
  INV_X1 U19501 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n16486) );
  AOI22_X1 U19502 ( .A1(n16487), .A2(n21034), .B1(n16486), .B2(U215), .ZN(U282) );
  INV_X1 U19503 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n16488) );
  OAI222_X1 U19504 ( .A1(P3_DATAO_REG_31__SCAN_IN), .A2(n16488), .B1(
        P1_DATAO_REG_31__SCAN_IN), .B2(n20043), .C1(P2_DATAO_REG_31__SCAN_IN), 
        .C2(n19080), .ZN(n16490) );
  INV_X2 U19505 ( .A(n16491), .ZN(n16489) );
  INV_X1 U19506 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18733) );
  INV_X1 U19507 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19859) );
  AOI22_X1 U19508 ( .A1(n16489), .A2(n18733), .B1(n19859), .B2(n16491), .ZN(
        U347) );
  INV_X1 U19509 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18731) );
  INV_X1 U19510 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19857) );
  AOI22_X1 U19511 ( .A1(n16489), .A2(n18731), .B1(n19857), .B2(n16491), .ZN(
        U348) );
  INV_X1 U19512 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18728) );
  INV_X1 U19513 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19856) );
  AOI22_X1 U19514 ( .A1(n16489), .A2(n18728), .B1(n19856), .B2(n16491), .ZN(
        U349) );
  INV_X1 U19515 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18727) );
  INV_X1 U19516 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19854) );
  AOI22_X1 U19517 ( .A1(n16489), .A2(n18727), .B1(n19854), .B2(n16491), .ZN(
        U350) );
  INV_X1 U19518 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18725) );
  INV_X1 U19519 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19852) );
  AOI22_X1 U19520 ( .A1(n16489), .A2(n18725), .B1(n19852), .B2(n16491), .ZN(
        U351) );
  INV_X1 U19521 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18723) );
  INV_X1 U19522 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19850) );
  AOI22_X1 U19523 ( .A1(n16489), .A2(n18723), .B1(n19850), .B2(n16491), .ZN(
        U352) );
  INV_X1 U19524 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18721) );
  INV_X1 U19525 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19849) );
  AOI22_X1 U19526 ( .A1(n16489), .A2(n18721), .B1(n19849), .B2(n16491), .ZN(
        U353) );
  INV_X1 U19527 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18720) );
  AOI22_X1 U19528 ( .A1(n16489), .A2(n18720), .B1(n19847), .B2(n16491), .ZN(
        U354) );
  INV_X1 U19529 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18774) );
  INV_X1 U19530 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19887) );
  AOI22_X1 U19531 ( .A1(n16489), .A2(n18774), .B1(n19887), .B2(n16490), .ZN(
        U355) );
  INV_X1 U19532 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18771) );
  INV_X1 U19533 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19885) );
  AOI22_X1 U19534 ( .A1(n16489), .A2(n18771), .B1(n19885), .B2(n16491), .ZN(
        U356) );
  INV_X1 U19535 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18767) );
  INV_X1 U19536 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19883) );
  AOI22_X1 U19537 ( .A1(n16489), .A2(n18767), .B1(n19883), .B2(n16491), .ZN(
        U357) );
  INV_X1 U19538 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18766) );
  INV_X1 U19539 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19880) );
  AOI22_X1 U19540 ( .A1(n16489), .A2(n18766), .B1(n19880), .B2(n16490), .ZN(
        U358) );
  INV_X1 U19541 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18764) );
  INV_X1 U19542 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19879) );
  AOI22_X1 U19543 ( .A1(n16489), .A2(n18764), .B1(n19879), .B2(n16490), .ZN(
        U359) );
  INV_X1 U19544 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18762) );
  INV_X1 U19545 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19878) );
  AOI22_X1 U19546 ( .A1(n16489), .A2(n18762), .B1(n19878), .B2(n16490), .ZN(
        U360) );
  INV_X1 U19547 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18759) );
  INV_X1 U19548 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19877) );
  AOI22_X1 U19549 ( .A1(n16489), .A2(n18759), .B1(n19877), .B2(n16490), .ZN(
        U361) );
  INV_X1 U19550 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18757) );
  INV_X1 U19551 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19876) );
  AOI22_X1 U19552 ( .A1(n16489), .A2(n18757), .B1(n19876), .B2(n16490), .ZN(
        U362) );
  INV_X1 U19553 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18755) );
  INV_X1 U19554 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n21079) );
  AOI22_X1 U19555 ( .A1(n16489), .A2(n18755), .B1(n21079), .B2(n16490), .ZN(
        U363) );
  INV_X1 U19556 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18753) );
  INV_X1 U19557 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19875) );
  AOI22_X1 U19558 ( .A1(n16489), .A2(n18753), .B1(n19875), .B2(n16491), .ZN(
        U364) );
  INV_X1 U19559 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18718) );
  INV_X1 U19560 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19846) );
  AOI22_X1 U19561 ( .A1(n16489), .A2(n18718), .B1(n19846), .B2(n16491), .ZN(
        U365) );
  INV_X1 U19562 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18751) );
  INV_X1 U19563 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19873) );
  AOI22_X1 U19564 ( .A1(n16489), .A2(n18751), .B1(n19873), .B2(n16491), .ZN(
        U366) );
  INV_X1 U19565 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18749) );
  INV_X1 U19566 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19872) );
  AOI22_X1 U19567 ( .A1(n16489), .A2(n18749), .B1(n19872), .B2(n16491), .ZN(
        U367) );
  INV_X1 U19568 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18747) );
  INV_X1 U19569 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19870) );
  AOI22_X1 U19570 ( .A1(n16489), .A2(n18747), .B1(n19870), .B2(n16491), .ZN(
        U368) );
  INV_X1 U19571 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18745) );
  INV_X1 U19572 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19868) );
  AOI22_X1 U19573 ( .A1(n16489), .A2(n18745), .B1(n19868), .B2(n16491), .ZN(
        U369) );
  INV_X1 U19574 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18743) );
  INV_X1 U19575 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19867) );
  AOI22_X1 U19576 ( .A1(n16489), .A2(n18743), .B1(n19867), .B2(n16491), .ZN(
        U370) );
  INV_X1 U19577 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18741) );
  INV_X1 U19578 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19866) );
  AOI22_X1 U19579 ( .A1(n16489), .A2(n18741), .B1(n19866), .B2(n16491), .ZN(
        U371) );
  INV_X1 U19580 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18740) );
  INV_X1 U19581 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19865) );
  AOI22_X1 U19582 ( .A1(n16489), .A2(n18740), .B1(n19865), .B2(n16491), .ZN(
        U372) );
  INV_X1 U19583 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18739) );
  INV_X1 U19584 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19863) );
  AOI22_X1 U19585 ( .A1(n16489), .A2(n18739), .B1(n19863), .B2(n16491), .ZN(
        U373) );
  INV_X1 U19586 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18737) );
  INV_X1 U19587 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19862) );
  AOI22_X1 U19588 ( .A1(n16489), .A2(n18737), .B1(n19862), .B2(n16491), .ZN(
        U374) );
  INV_X1 U19589 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18735) );
  INV_X1 U19590 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19860) );
  AOI22_X1 U19591 ( .A1(n16489), .A2(n18735), .B1(n19860), .B2(n16490), .ZN(
        U375) );
  INV_X1 U19592 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18715) );
  INV_X1 U19593 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19844) );
  AOI22_X1 U19594 ( .A1(n16489), .A2(n18715), .B1(n19844), .B2(n16491), .ZN(
        U376) );
  INV_X1 U19595 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18714) );
  NAND2_X1 U19596 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18714), .ZN(n18702) );
  INV_X1 U19597 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18712) );
  AOI22_X1 U19598 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18702), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18712), .ZN(n18784) );
  AOI21_X1 U19599 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18784), .ZN(n16492) );
  INV_X1 U19600 ( .A(n16492), .ZN(P3_U2633) );
  INV_X1 U19601 ( .A(n16517), .ZN(n18689) );
  INV_X1 U19602 ( .A(n17415), .ZN(n17414) );
  OAI21_X1 U19603 ( .B1(n16497), .B2(n17414), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16493) );
  OAI21_X1 U19604 ( .B1(n16494), .B2(n18689), .A(n16493), .ZN(P3_U2634) );
  AOI21_X1 U19605 ( .B1(n18712), .B2(n18714), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16495) );
  AOI22_X1 U19606 ( .A1(n18779), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16495), 
        .B2(n18843), .ZN(P3_U2635) );
  OAI21_X1 U19607 ( .B1(n18698), .B2(BS16), .A(n18784), .ZN(n18782) );
  OAI21_X1 U19608 ( .B1(n18784), .B2(n18834), .A(n18782), .ZN(P3_U2636) );
  NOR3_X1 U19609 ( .A1(n16497), .A2(n16496), .A3(n18654), .ZN(n18669) );
  NOR2_X1 U19610 ( .A1(n18669), .A2(n18685), .ZN(n18827) );
  OAI21_X1 U19611 ( .B1(n18827), .B2(n18175), .A(n16498), .ZN(P3_U2637) );
  NOR4_X1 U19612 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16502) );
  NOR4_X1 U19613 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_15__SCAN_IN), .A3(P3_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16501) );
  NOR4_X1 U19614 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16500) );
  NOR4_X1 U19615 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16499) );
  NAND4_X1 U19616 ( .A1(n16502), .A2(n16501), .A3(n16500), .A4(n16499), .ZN(
        n16508) );
  NOR4_X1 U19617 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16506) );
  AOI211_X1 U19618 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_4__SCAN_IN), .B(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16505) );
  NOR4_X1 U19619 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_10__SCAN_IN), .A3(P3_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_13__SCAN_IN), .ZN(n16504) );
  NOR4_X1 U19620 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_8__SCAN_IN), .ZN(n16503) );
  NAND4_X1 U19621 ( .A1(n16506), .A2(n16505), .A3(n16504), .A4(n16503), .ZN(
        n16507) );
  NOR2_X1 U19622 ( .A1(n16508), .A2(n16507), .ZN(n18826) );
  INV_X1 U19623 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16510) );
  NOR3_X1 U19624 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16511) );
  OAI21_X1 U19625 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16511), .A(n18826), .ZN(
        n16509) );
  OAI21_X1 U19626 ( .B1(n18826), .B2(n16510), .A(n16509), .ZN(P3_U2638) );
  INV_X1 U19627 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18716) );
  INV_X1 U19628 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18783) );
  AOI21_X1 U19629 ( .B1(n18716), .B2(n18783), .A(n16511), .ZN(n16513) );
  INV_X1 U19630 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16512) );
  INV_X1 U19631 ( .A(n18826), .ZN(n18823) );
  AOI22_X1 U19632 ( .A1(n18826), .A2(n16513), .B1(n16512), .B2(n18823), .ZN(
        P3_U2639) );
  NAND2_X1 U19633 ( .A1(n16515), .A2(n16514), .ZN(n18653) );
  NAND3_X1 U19634 ( .A1(n16516), .A2(n18687), .A3(n18834), .ZN(n18695) );
  NAND2_X1 U19635 ( .A1(n16517), .A2(n9722), .ZN(n18683) );
  OAI211_X1 U19636 ( .C1(n16523), .C2(n16518), .A(n18836), .B(n18834), .ZN(
        n18679) );
  INV_X1 U19637 ( .A(n18679), .ZN(n16519) );
  AOI211_X1 U19638 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n16523), .A(n16519), .B(
        n16525), .ZN(n16520) );
  INV_X1 U19639 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18775) );
  INV_X1 U19640 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18768) );
  INV_X1 U19641 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18761) );
  INV_X1 U19642 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18756) );
  INV_X1 U19643 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18752) );
  INV_X1 U19644 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18748) );
  INV_X1 U19645 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18746) );
  INV_X1 U19646 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n21154) );
  INV_X1 U19647 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18738) );
  INV_X1 U19648 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18736) );
  INV_X1 U19649 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18726) );
  INV_X1 U19650 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18722) );
  INV_X1 U19651 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n20931) );
  NAND2_X1 U19652 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16850) );
  NOR2_X1 U19653 ( .A1(n20931), .A2(n16850), .ZN(n16843) );
  NAND2_X1 U19654 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16843), .ZN(n16825) );
  NOR2_X1 U19655 ( .A1(n18722), .A2(n16825), .ZN(n16819) );
  NAND2_X1 U19656 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16819), .ZN(n16800) );
  NOR2_X1 U19657 ( .A1(n18726), .A2(n16800), .ZN(n16786) );
  NAND2_X1 U19658 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16786), .ZN(n16769) );
  INV_X1 U19659 ( .A(n16769), .ZN(n16521) );
  INV_X1 U19660 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18732) );
  INV_X1 U19661 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18730) );
  NOR2_X1 U19662 ( .A1(n18732), .A2(n18730), .ZN(n16750) );
  NAND3_X1 U19663 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16521), .A3(n16750), 
        .ZN(n16744) );
  OR2_X1 U19664 ( .A1(n18736), .A2(n16744), .ZN(n16729) );
  NOR2_X1 U19665 ( .A1(n18738), .A2(n16729), .ZN(n16715) );
  NAND2_X1 U19666 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16715), .ZN(n16694) );
  NOR2_X1 U19667 ( .A1(n21154), .A2(n16694), .ZN(n16680) );
  NAND3_X1 U19668 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(n16680), .ZN(n16660) );
  NOR3_X1 U19669 ( .A1(n18748), .A2(n18746), .A3(n16660), .ZN(n16654) );
  NAND2_X1 U19670 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16654), .ZN(n16646) );
  NOR2_X1 U19671 ( .A1(n18752), .A2(n16646), .ZN(n16628) );
  NAND2_X1 U19672 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16628), .ZN(n16620) );
  NAND2_X1 U19673 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16618), .ZN(n16600) );
  NOR2_X1 U19674 ( .A1(n18761), .A2(n16600), .ZN(n16587) );
  NAND2_X1 U19675 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16587), .ZN(n16538) );
  NOR2_X1 U19676 ( .A1(n16894), .A2(n16538), .ZN(n16578) );
  NAND2_X1 U19677 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16578), .ZN(n16566) );
  NOR2_X1 U19678 ( .A1(n18768), .A2(n16566), .ZN(n16560) );
  NAND2_X1 U19679 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16560), .ZN(n16540) );
  NOR3_X1 U19680 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18775), .A3(n16540), 
        .ZN(n16522) );
  AOI21_X1 U19681 ( .B1(n16888), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16522), .ZN(
        n16543) );
  NAND2_X1 U19682 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n16523), .ZN(n16524) );
  AOI211_X4 U19683 ( .C1(n18834), .C2(n18836), .A(n16525), .B(n16524), .ZN(
        n16862) );
  NOR3_X1 U19684 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16867) );
  INV_X1 U19685 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17201) );
  NAND2_X1 U19686 ( .A1(n16867), .A2(n17201), .ZN(n16861) );
  NOR2_X1 U19687 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16861), .ZN(n16841) );
  INV_X1 U19688 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16837) );
  NAND2_X1 U19689 ( .A1(n16841), .A2(n16837), .ZN(n16829) );
  NAND2_X1 U19690 ( .A1(n16811), .A2(n16796), .ZN(n16798) );
  INV_X1 U19691 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16784) );
  NAND2_X1 U19692 ( .A1(n16785), .A2(n16784), .ZN(n16763) );
  INV_X1 U19693 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16760) );
  NAND2_X1 U19694 ( .A1(n16762), .A2(n16760), .ZN(n16757) );
  INV_X1 U19695 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16735) );
  NAND2_X1 U19696 ( .A1(n16742), .A2(n16735), .ZN(n16734) );
  INV_X1 U19697 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16707) );
  NAND2_X1 U19698 ( .A1(n16719), .A2(n16707), .ZN(n16705) );
  INV_X1 U19699 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16690) );
  NAND2_X1 U19700 ( .A1(n16691), .A2(n16690), .ZN(n16687) );
  INV_X1 U19701 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16665) );
  NAND2_X1 U19702 ( .A1(n16673), .A2(n16665), .ZN(n16664) );
  INV_X1 U19703 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n21016) );
  NAND2_X1 U19704 ( .A1(n16648), .A2(n21016), .ZN(n16643) );
  INV_X1 U19705 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16956) );
  NAND2_X1 U19706 ( .A1(n16629), .A2(n16956), .ZN(n16623) );
  NAND2_X1 U19707 ( .A1(n16608), .A2(n16901), .ZN(n16603) );
  NAND2_X1 U19708 ( .A1(n16596), .A2(n16945), .ZN(n16579) );
  INV_X1 U19709 ( .A(n16579), .ZN(n16570) );
  NAND2_X1 U19710 ( .A1(n21075), .A2(n16570), .ZN(n16569) );
  NOR2_X1 U19711 ( .A1(n16892), .A2(n16545), .ZN(n16551) );
  INV_X1 U19712 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16907) );
  INV_X1 U19713 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16565) );
  NAND2_X1 U19714 ( .A1(n16528), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16527) );
  AOI21_X1 U19715 ( .B1(n16565), .B2(n16527), .A(n16526), .ZN(n17487) );
  OAI21_X1 U19716 ( .B1(n16528), .B2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16527), .ZN(n17507) );
  INV_X1 U19717 ( .A(n17507), .ZN(n16576) );
  INV_X1 U19718 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16590) );
  NOR2_X1 U19719 ( .A1(n17849), .A2(n17532), .ZN(n16531) );
  INV_X1 U19720 ( .A(n16531), .ZN(n16532) );
  NOR2_X1 U19721 ( .A1(n17533), .A2(n16532), .ZN(n17484) );
  INV_X1 U19722 ( .A(n17484), .ZN(n16529) );
  AOI21_X1 U19723 ( .B1(n16590), .B2(n16529), .A(n16528), .ZN(n17519) );
  INV_X1 U19724 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17535) );
  NAND2_X1 U19725 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16531), .ZN(
        n16530) );
  AOI21_X1 U19726 ( .B1(n17535), .B2(n16530), .A(n17484), .ZN(n17537) );
  INV_X1 U19727 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17547) );
  AOI22_X1 U19728 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16531), .B1(
        n16532), .B2(n17547), .ZN(n17550) );
  NAND2_X1 U19729 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9802), .ZN(
        n16658) );
  NAND2_X1 U19730 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17580), .ZN(
        n16535) );
  NOR2_X1 U19731 ( .A1(n17584), .A2(n16535), .ZN(n17531) );
  OAI21_X1 U19732 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17531), .A(
        n16532), .ZN(n16533) );
  INV_X1 U19733 ( .A(n16533), .ZN(n17562) );
  INV_X1 U19734 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16637) );
  INV_X1 U19735 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17595) );
  OR2_X1 U19736 ( .A1(n17595), .A2(n16535), .ZN(n16534) );
  AOI21_X1 U19737 ( .B1(n16637), .B2(n16534), .A(n17531), .ZN(n17582) );
  XOR2_X1 U19738 ( .A(n17595), .B(n16535), .Z(n17591) );
  OAI21_X1 U19739 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17580), .A(
        n16535), .ZN(n16536) );
  INV_X1 U19740 ( .A(n16536), .ZN(n17610) );
  INV_X1 U19741 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n21128) );
  INV_X1 U19742 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17664) );
  INV_X1 U19743 ( .A(n16537), .ZN(n17655) );
  NAND2_X1 U19744 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17655), .ZN(
        n17653) );
  NOR2_X1 U19745 ( .A1(n17664), .A2(n17653), .ZN(n16710) );
  AOI21_X1 U19746 ( .B1(n21128), .B2(n16710), .A(n16852), .ZN(n16700) );
  INV_X1 U19747 ( .A(n16700), .ZN(n16699) );
  OAI21_X1 U19748 ( .B1(n17580), .B2(n16852), .A(n16699), .ZN(n16650) );
  NOR2_X1 U19749 ( .A1(n17610), .A2(n16650), .ZN(n16649) );
  NOR2_X1 U19750 ( .A1(n16649), .A2(n16852), .ZN(n16639) );
  NOR2_X1 U19751 ( .A1(n17591), .A2(n16639), .ZN(n16638) );
  NOR2_X1 U19752 ( .A1(n16638), .A2(n16852), .ZN(n16631) );
  NOR2_X1 U19753 ( .A1(n17582), .A2(n16631), .ZN(n16630) );
  NOR2_X1 U19754 ( .A1(n16630), .A2(n16852), .ZN(n16617) );
  NOR2_X1 U19755 ( .A1(n17562), .A2(n16617), .ZN(n16616) );
  NOR2_X1 U19756 ( .A1(n16616), .A2(n16852), .ZN(n16610) );
  NOR2_X1 U19757 ( .A1(n17519), .A2(n16586), .ZN(n16585) );
  NOR2_X1 U19758 ( .A1(n16564), .A2(n16852), .ZN(n16555) );
  NOR2_X1 U19759 ( .A1(n16556), .A2(n16555), .ZN(n16554) );
  NOR2_X1 U19760 ( .A1(n16852), .A2(n18693), .ZN(n16881) );
  INV_X1 U19761 ( .A(n16881), .ZN(n16728) );
  NAND3_X1 U19762 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16539) );
  NAND2_X1 U19763 ( .A1(n16876), .A2(n16538), .ZN(n16588) );
  NAND2_X1 U19764 ( .A1(n16897), .A2(n16588), .ZN(n16593) );
  AOI21_X1 U19765 ( .B1(n16876), .B2(n16539), .A(n16593), .ZN(n16563) );
  NOR2_X1 U19766 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16540), .ZN(n16549) );
  INV_X1 U19767 ( .A(n16549), .ZN(n16541) );
  AOI21_X1 U19768 ( .B1(n16563), .B2(n16541), .A(n18772), .ZN(n16542) );
  NAND2_X1 U19769 ( .A1(n16862), .A2(n16545), .ZN(n16557) );
  XOR2_X1 U19770 ( .A(n16547), .B(n16546), .Z(n16550) );
  OAI22_X1 U19771 ( .A1(n16563), .A2(n18775), .B1(n10020), .B2(n16868), .ZN(
        n16548) );
  AOI211_X1 U19772 ( .C1(n16550), .C2(n16853), .A(n16549), .B(n16548), .ZN(
        n16553) );
  OAI21_X1 U19773 ( .B1(n16888), .B2(n16551), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16552) );
  OAI211_X1 U19774 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16557), .A(n16553), .B(
        n16552), .ZN(P3_U2641) );
  INV_X1 U19775 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18770) );
  AOI22_X1 U19776 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16880), .B1(
        n16888), .B2(P3_EBX_REG_29__SCAN_IN), .ZN(n16562) );
  AOI211_X1 U19777 ( .C1(n16556), .C2(n16555), .A(n16554), .B(n18693), .ZN(
        n16559) );
  AOI21_X1 U19778 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16569), .A(n16557), .ZN(
        n16558) );
  AOI211_X1 U19779 ( .C1(n16560), .C2(n18770), .A(n16559), .B(n16558), .ZN(
        n16561) );
  OAI211_X1 U19780 ( .C1(n16563), .C2(n18770), .A(n16562), .B(n16561), .ZN(
        P3_U2642) );
  INV_X1 U19781 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18765) );
  AOI21_X1 U19782 ( .B1(n16578), .B2(n18765), .A(n16593), .ZN(n16573) );
  AOI211_X1 U19783 ( .C1(n17487), .C2(n10009), .A(n16564), .B(n18693), .ZN(
        n16568) );
  OAI22_X1 U19784 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n16566), .B1(n16565), 
        .B2(n16868), .ZN(n16567) );
  AOI211_X1 U19785 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16888), .A(n16568), .B(
        n16567), .ZN(n16572) );
  OAI211_X1 U19786 ( .C1(n16570), .C2(n21075), .A(n16862), .B(n16569), .ZN(
        n16571) );
  OAI211_X1 U19787 ( .C1(n16573), .C2(n18768), .A(n16572), .B(n16571), .ZN(
        P3_U2643) );
  AOI22_X1 U19788 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16880), .B1(
        n16888), .B2(P3_EBX_REG_27__SCAN_IN), .ZN(n16583) );
  AOI211_X1 U19789 ( .C1(n16576), .C2(n16575), .A(n16574), .B(n18693), .ZN(
        n16577) );
  AOI21_X1 U19790 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n16593), .A(n16577), 
        .ZN(n16582) );
  NAND2_X1 U19791 ( .A1(n16578), .A2(n18765), .ZN(n16581) );
  OAI211_X1 U19792 ( .C1(n16596), .C2(n16945), .A(n16862), .B(n16579), .ZN(
        n16580) );
  NAND4_X1 U19793 ( .A1(n16583), .A2(n16582), .A3(n16581), .A4(n16580), .ZN(
        P3_U2644) );
  AOI21_X1 U19794 ( .B1(n16603), .B2(P3_EBX_REG_26__SCAN_IN), .A(n16892), .ZN(
        n16584) );
  AOI21_X1 U19795 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n16888), .A(n16584), .ZN(
        n16595) );
  AOI211_X1 U19796 ( .C1(n17519), .C2(n16586), .A(n16585), .B(n18693), .ZN(
        n16592) );
  INV_X1 U19797 ( .A(n16587), .ZN(n16589) );
  OAI22_X1 U19798 ( .A1(n16590), .A2(n16868), .B1(n16589), .B2(n16588), .ZN(
        n16591) );
  AOI211_X1 U19799 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16593), .A(n16592), 
        .B(n16591), .ZN(n16594) );
  OAI21_X1 U19800 ( .B1(n16596), .B2(n16595), .A(n16594), .ZN(P3_U2645) );
  INV_X1 U19801 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18758) );
  OAI21_X1 U19802 ( .B1(n16618), .B2(n16894), .A(n16897), .ZN(n16615) );
  AOI21_X1 U19803 ( .B1(n16876), .B2(n18758), .A(n16615), .ZN(n16606) );
  AOI211_X1 U19804 ( .C1(n17537), .C2(n16598), .A(n16597), .B(n18693), .ZN(
        n16602) );
  NAND2_X1 U19805 ( .A1(n16876), .A2(n18761), .ZN(n16599) );
  OAI22_X1 U19806 ( .A1(n17535), .A2(n16868), .B1(n16600), .B2(n16599), .ZN(
        n16601) );
  AOI211_X1 U19807 ( .C1(P3_EBX_REG_25__SCAN_IN), .C2(n16888), .A(n16602), .B(
        n16601), .ZN(n16605) );
  OAI211_X1 U19808 ( .C1(n16608), .C2(n16901), .A(n16862), .B(n16603), .ZN(
        n16604) );
  OAI211_X1 U19809 ( .C1(n16606), .C2(n18761), .A(n16605), .B(n16604), .ZN(
        P3_U2646) );
  NOR2_X1 U19810 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16894), .ZN(n16607) );
  AOI22_X1 U19811 ( .A1(n16888), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16618), 
        .B2(n16607), .ZN(n16614) );
  AOI211_X1 U19812 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16623), .A(n16608), .B(
        n16892), .ZN(n16612) );
  AOI211_X1 U19813 ( .C1(n17550), .C2(n16610), .A(n16609), .B(n18693), .ZN(
        n16611) );
  AOI211_X1 U19814 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16615), .A(n16612), 
        .B(n16611), .ZN(n16613) );
  OAI211_X1 U19815 ( .C1(n17547), .C2(n16868), .A(n16614), .B(n16613), .ZN(
        P3_U2647) );
  INV_X1 U19816 ( .A(n16615), .ZN(n16626) );
  AOI211_X1 U19817 ( .C1(n17562), .C2(n16617), .A(n16616), .B(n18693), .ZN(
        n16622) );
  INV_X1 U19818 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n21169) );
  OR2_X1 U19819 ( .A1(n16894), .A2(n16618), .ZN(n16619) );
  OAI22_X1 U19820 ( .A1(n21169), .A2(n16868), .B1(n16620), .B2(n16619), .ZN(
        n16621) );
  AOI211_X1 U19821 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n16888), .A(n16622), .B(
        n16621), .ZN(n16625) );
  OAI211_X1 U19822 ( .C1(n16629), .C2(n16956), .A(n16862), .B(n16623), .ZN(
        n16624) );
  OAI211_X1 U19823 ( .C1(n16626), .C2(n18756), .A(n16625), .B(n16624), .ZN(
        P3_U2648) );
  NOR2_X1 U19824 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16894), .ZN(n16627) );
  AOI22_X1 U19825 ( .A1(n16888), .A2(P3_EBX_REG_22__SCAN_IN), .B1(n16628), 
        .B2(n16627), .ZN(n16636) );
  AOI21_X1 U19826 ( .B1(n16876), .B2(n16646), .A(n16768), .ZN(n16657) );
  OAI21_X1 U19827 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n16894), .A(n16657), 
        .ZN(n16634) );
  AOI211_X1 U19828 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16643), .A(n16629), .B(
        n16892), .ZN(n16633) );
  AOI211_X1 U19829 ( .C1(n17582), .C2(n16631), .A(n16630), .B(n18693), .ZN(
        n16632) );
  AOI211_X1 U19830 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16634), .A(n16633), 
        .B(n16632), .ZN(n16635) );
  OAI211_X1 U19831 ( .C1(n16637), .C2(n16868), .A(n16636), .B(n16635), .ZN(
        P3_U2649) );
  NAND2_X1 U19832 ( .A1(n16876), .A2(n18752), .ZN(n16647) );
  INV_X1 U19833 ( .A(n16657), .ZN(n16642) );
  AOI211_X1 U19834 ( .C1(n17591), .C2(n16639), .A(n16638), .B(n18693), .ZN(
        n16641) );
  OAI22_X1 U19835 ( .A1(n17595), .A2(n16868), .B1(n16893), .B2(n21016), .ZN(
        n16640) );
  AOI211_X1 U19836 ( .C1(n16642), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16641), 
        .B(n16640), .ZN(n16645) );
  OAI211_X1 U19837 ( .C1(n16648), .C2(n21016), .A(n16862), .B(n16643), .ZN(
        n16644) );
  OAI211_X1 U19838 ( .C1(n16647), .C2(n16646), .A(n16645), .B(n16644), .ZN(
        P3_U2650) );
  INV_X1 U19839 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18750) );
  AOI22_X1 U19840 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n16880), .B1(
        n16888), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n16656) );
  NOR2_X1 U19841 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16894), .ZN(n16653) );
  AOI211_X1 U19842 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16664), .A(n16648), .B(
        n16892), .ZN(n16652) );
  AOI211_X1 U19843 ( .C1(n17610), .C2(n16650), .A(n16649), .B(n18693), .ZN(
        n16651) );
  AOI211_X1 U19844 ( .C1(n16654), .C2(n16653), .A(n16652), .B(n16651), .ZN(
        n16655) );
  OAI211_X1 U19845 ( .C1(n18750), .C2(n16657), .A(n16656), .B(n16655), .ZN(
        P3_U2651) );
  AOI22_X1 U19846 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n16880), .B1(
        n16888), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n16668) );
  NOR2_X1 U19847 ( .A1(n17849), .A2(n17617), .ZN(n17616) );
  NAND2_X1 U19848 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17616), .ZN(
        n16669) );
  INV_X1 U19849 ( .A(n16669), .ZN(n16659) );
  OAI21_X1 U19850 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16659), .A(
        n16658), .ZN(n17620) );
  AOI21_X1 U19851 ( .B1(n16669), .B2(n16815), .A(n16700), .ZN(n16672) );
  XOR2_X1 U19852 ( .A(n17620), .B(n16672), .Z(n16663) );
  NAND4_X1 U19853 ( .A1(n16876), .A2(P3_REIP_REG_17__SCAN_IN), .A3(
        P3_REIP_REG_16__SCAN_IN), .A4(n16680), .ZN(n16679) );
  XOR2_X1 U19854 ( .A(P3_REIP_REG_19__SCAN_IN), .B(n18746), .Z(n16661) );
  AOI21_X1 U19855 ( .B1(n16876), .B2(n16660), .A(n16768), .ZN(n16684) );
  OAI22_X1 U19856 ( .A1(n16679), .A2(n16661), .B1(n18748), .B2(n16684), .ZN(
        n16662) );
  AOI21_X1 U19857 ( .B1(n16663), .B2(n16853), .A(n16662), .ZN(n16667) );
  OAI211_X1 U19858 ( .C1(n16673), .C2(n16665), .A(n16862), .B(n16664), .ZN(
        n16666) );
  NAND4_X1 U19859 ( .A1(n16668), .A2(n16667), .A3(n18169), .A4(n16666), .ZN(
        P3_U2652) );
  OAI21_X1 U19860 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17616), .A(
        n16669), .ZN(n17629) );
  NOR2_X1 U19861 ( .A1(n18693), .A2(n16815), .ZN(n16805) );
  INV_X1 U19862 ( .A(n16805), .ZN(n16879) );
  NOR2_X1 U19863 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16670) );
  OAI21_X1 U19864 ( .B1(n16670), .B2(n17629), .A(n16853), .ZN(n16671) );
  AOI22_X1 U19865 ( .A1(n16672), .A2(n17629), .B1(n16879), .B2(n16671), .ZN(
        n16677) );
  AOI211_X1 U19866 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16687), .A(n16673), .B(
        n16892), .ZN(n16676) );
  AOI22_X1 U19867 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16880), .B1(
        n16888), .B2(P3_EBX_REG_18__SCAN_IN), .ZN(n16674) );
  INV_X1 U19868 ( .A(n16674), .ZN(n16675) );
  NOR4_X1 U19869 ( .A1(n9736), .A2(n16677), .A3(n16676), .A4(n16675), .ZN(
        n16678) );
  OAI221_X1 U19870 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16679), .C1(n18746), 
        .C2(n16684), .A(n16678), .ZN(P3_U2653) );
  AND2_X1 U19871 ( .A1(n16876), .A2(n16680), .ZN(n16693) );
  AOI21_X1 U19872 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(n16693), .A(
        P3_REIP_REG_17__SCAN_IN), .ZN(n16685) );
  NOR2_X1 U19873 ( .A1(n17656), .A2(n17653), .ZN(n16696) );
  AOI21_X1 U19874 ( .B1(n16696), .B2(n21128), .A(n16852), .ZN(n16682) );
  INV_X1 U19875 ( .A(n17616), .ZN(n16681) );
  OAI21_X1 U19876 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16696), .A(
        n16681), .ZN(n17641) );
  XOR2_X1 U19877 ( .A(n16682), .B(n17641), .Z(n16683) );
  OAI22_X1 U19878 ( .A1(n16685), .A2(n16684), .B1(n18693), .B2(n16683), .ZN(
        n16686) );
  AOI211_X1 U19879 ( .C1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(n16880), .A(
        n9736), .B(n16686), .ZN(n16689) );
  OAI211_X1 U19880 ( .C1(n16691), .C2(n16690), .A(n16862), .B(n16687), .ZN(
        n16688) );
  OAI211_X1 U19881 ( .C1(n16690), .C2(n16893), .A(n16689), .B(n16688), .ZN(
        P3_U2654) );
  AOI22_X1 U19882 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16880), .B1(
        n16888), .B2(P3_EBX_REG_16__SCAN_IN), .ZN(n16704) );
  INV_X1 U19883 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18742) );
  AOI211_X1 U19884 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16705), .A(n16691), .B(
        n16892), .ZN(n16692) );
  AOI211_X1 U19885 ( .C1(n16693), .C2(n18742), .A(n9736), .B(n16692), .ZN(
        n16703) );
  AOI21_X1 U19886 ( .B1(n16876), .B2(n16694), .A(n16768), .ZN(n16724) );
  INV_X1 U19887 ( .A(n16724), .ZN(n16695) );
  NOR3_X1 U19888 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16894), .A3(n16694), 
        .ZN(n16709) );
  OAI21_X1 U19889 ( .B1(n16695), .B2(n16709), .A(P3_REIP_REG_16__SCAN_IN), 
        .ZN(n16702) );
  INV_X1 U19890 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17659) );
  INV_X1 U19891 ( .A(n16710), .ZN(n16697) );
  AOI21_X1 U19892 ( .B1(n17659), .B2(n16697), .A(n16696), .ZN(n17658) );
  INV_X1 U19893 ( .A(n17658), .ZN(n16698) );
  OAI221_X1 U19894 ( .B1(n16700), .B2(n17658), .C1(n16699), .C2(n16698), .A(
        n16853), .ZN(n16701) );
  NAND4_X1 U19895 ( .A1(n16704), .A2(n16703), .A3(n16702), .A4(n16701), .ZN(
        P3_U2655) );
  OAI211_X1 U19896 ( .C1(n16719), .C2(n16707), .A(n16862), .B(n16705), .ZN(
        n16706) );
  OAI211_X1 U19897 ( .C1(n16893), .C2(n16707), .A(n18169), .B(n16706), .ZN(
        n16708) );
  AOI211_X1 U19898 ( .C1(n16880), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16709), .B(n16708), .ZN(n16714) );
  AOI21_X1 U19899 ( .B1(n17664), .B2(n17653), .A(n16710), .ZN(n17672) );
  NOR2_X1 U19900 ( .A1(n17849), .A2(n17701), .ZN(n17690) );
  INV_X1 U19901 ( .A(n17690), .ZN(n16751) );
  NOR2_X1 U19902 ( .A1(n17703), .A2(n16751), .ZN(n16725) );
  OAI21_X1 U19903 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16725), .A(
        n17653), .ZN(n17680) );
  INV_X1 U19904 ( .A(n17680), .ZN(n16718) );
  NOR2_X1 U19905 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17849), .ZN(
        n16869) );
  AOI21_X1 U19906 ( .B1(n17678), .B2(n16869), .A(n16852), .ZN(n16717) );
  NOR2_X1 U19907 ( .A1(n16718), .A2(n16717), .ZN(n16716) );
  NOR2_X1 U19908 ( .A1(n16716), .A2(n16852), .ZN(n16712) );
  AOI21_X1 U19909 ( .B1(n17672), .B2(n16712), .A(n18693), .ZN(n16711) );
  OAI21_X1 U19910 ( .B1(n17672), .B2(n16712), .A(n16711), .ZN(n16713) );
  OAI211_X1 U19911 ( .C1(n16724), .C2(n21154), .A(n16714), .B(n16713), .ZN(
        P3_U2656) );
  INV_X1 U19912 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n20962) );
  AOI211_X1 U19913 ( .C1(n16888), .C2(P3_EBX_REG_14__SCAN_IN), .A(n9736), .B(
        n10264), .ZN(n16723) );
  AOI211_X1 U19914 ( .C1(n16718), .C2(n16717), .A(n16716), .B(n18693), .ZN(
        n16721) );
  AOI211_X1 U19915 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16734), .A(n16719), .B(
        n16892), .ZN(n16720) );
  AOI211_X1 U19916 ( .C1(n16880), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16721), .B(n16720), .ZN(n16722) );
  OAI211_X1 U19917 ( .C1(n20962), .C2(n16724), .A(n16723), .B(n16722), .ZN(
        P3_U2657) );
  AOI22_X1 U19918 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n16880), .B1(
        n16888), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n16738) );
  NAND2_X1 U19919 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17690), .ZN(
        n16740) );
  OAI21_X1 U19920 ( .B1(n16852), .B2(n21128), .A(n16853), .ZN(n16891) );
  INV_X1 U19921 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16726) );
  AOI21_X1 U19922 ( .B1(n16726), .B2(n16740), .A(n16725), .ZN(n17691) );
  INV_X1 U19923 ( .A(n17691), .ZN(n16727) );
  AOI211_X1 U19924 ( .C1(n16815), .C2(n16740), .A(n16891), .B(n16727), .ZN(
        n16733) );
  AOI21_X1 U19925 ( .B1(n16876), .B2(n16744), .A(n16768), .ZN(n16754) );
  NAND2_X1 U19926 ( .A1(n16876), .A2(n18736), .ZN(n16743) );
  AOI21_X1 U19927 ( .B1(n16754), .B2(n16743), .A(n18738), .ZN(n16732) );
  AOI211_X1 U19928 ( .C1(n17678), .C2(n16869), .A(n17691), .B(n16728), .ZN(
        n16731) );
  NOR3_X1 U19929 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16894), .A3(n16729), 
        .ZN(n16730) );
  NOR4_X1 U19930 ( .A1(n16733), .A2(n16732), .A3(n16731), .A4(n16730), .ZN(
        n16737) );
  OAI211_X1 U19931 ( .C1(n16742), .C2(n16735), .A(n16862), .B(n16734), .ZN(
        n16736) );
  NAND4_X1 U19932 ( .A1(n16738), .A2(n16737), .A3(n18169), .A4(n16736), .ZN(
        P3_U2658) );
  AOI22_X1 U19933 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16880), .B1(
        n16888), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n16749) );
  INV_X1 U19934 ( .A(n17701), .ZN(n16739) );
  AOI21_X1 U19935 ( .B1(n16739), .B2(n16869), .A(n16852), .ZN(n16741) );
  OAI21_X1 U19936 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17690), .A(
        n16740), .ZN(n17708) );
  XNOR2_X1 U19937 ( .A(n16741), .B(n17708), .ZN(n16747) );
  AOI211_X1 U19938 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16757), .A(n16742), .B(
        n16892), .ZN(n16746) );
  OAI21_X1 U19939 ( .B1(n16744), .B2(n16743), .A(n18169), .ZN(n16745) );
  AOI211_X1 U19940 ( .C1(n16747), .C2(n16853), .A(n16746), .B(n16745), .ZN(
        n16748) );
  OAI211_X1 U19941 ( .C1(n18736), .C2(n16754), .A(n16749), .B(n16748), .ZN(
        P3_U2659) );
  NOR2_X1 U19942 ( .A1(n16894), .A2(n16769), .ZN(n16764) );
  AOI21_X1 U19943 ( .B1(n16750), .B2(n16764), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16755) );
  INV_X1 U19944 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16788) );
  NAND3_X1 U19945 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17757), .A3(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16802) );
  NOR2_X1 U19946 ( .A1(n16788), .A2(n16802), .ZN(n16787) );
  NAND2_X1 U19947 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16787), .ZN(
        n16773) );
  NOR2_X1 U19948 ( .A1(n17735), .A2(n16773), .ZN(n16761) );
  AOI21_X1 U19949 ( .B1(n16761), .B2(n21128), .A(n16852), .ZN(n16752) );
  OAI21_X1 U19950 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16761), .A(
        n16751), .ZN(n17727) );
  XOR2_X1 U19951 ( .A(n16752), .B(n17727), .Z(n16753) );
  OAI22_X1 U19952 ( .A1(n16755), .A2(n16754), .B1(n18693), .B2(n16753), .ZN(
        n16756) );
  AOI211_X1 U19953 ( .C1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n16880), .A(
        n9736), .B(n16756), .ZN(n16759) );
  OAI211_X1 U19954 ( .C1(n16762), .C2(n16760), .A(n16862), .B(n16757), .ZN(
        n16758) );
  OAI211_X1 U19955 ( .C1(n16760), .C2(n16893), .A(n16759), .B(n16758), .ZN(
        P3_U2660) );
  AOI21_X1 U19956 ( .B1(n17735), .B2(n16773), .A(n16761), .ZN(n17738) );
  OAI21_X1 U19957 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16773), .A(
        n16815), .ZN(n16775) );
  XOR2_X1 U19958 ( .A(n17738), .B(n16775), .Z(n16772) );
  AOI211_X1 U19959 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16763), .A(n16762), .B(
        n16892), .ZN(n16767) );
  NAND3_X1 U19960 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16764), .A3(n18732), 
        .ZN(n16765) );
  OAI211_X1 U19961 ( .C1(n17735), .C2(n16868), .A(n18169), .B(n16765), .ZN(
        n16766) );
  AOI211_X1 U19962 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16888), .A(n16767), .B(
        n16766), .ZN(n16771) );
  AOI21_X1 U19963 ( .B1(n16769), .B2(n16876), .A(n16768), .ZN(n16790) );
  INV_X1 U19964 ( .A(n16790), .ZN(n16780) );
  NOR3_X1 U19965 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16769), .A3(n16894), .ZN(
        n16779) );
  OAI21_X1 U19966 ( .B1(n16780), .B2(n16779), .A(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n16770) );
  OAI211_X1 U19967 ( .C1(n16772), .C2(n18693), .A(n16771), .B(n16770), .ZN(
        P3_U2661) );
  AOI21_X1 U19968 ( .B1(n16862), .B2(n16785), .A(n16888), .ZN(n16783) );
  OAI21_X1 U19969 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16787), .A(
        n16773), .ZN(n17750) );
  OAI221_X1 U19970 ( .B1(n17750), .B2(n16774), .C1(n17750), .C2(n21128), .A(
        n16853), .ZN(n16776) );
  AOI22_X1 U19971 ( .A1(n16776), .A2(n16879), .B1(n17750), .B2(n16775), .ZN(
        n16777) );
  AOI211_X1 U19972 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n16880), .A(
        n9736), .B(n16777), .ZN(n16782) );
  NOR3_X1 U19973 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n16785), .A3(n16892), .ZN(
        n16778) );
  AOI211_X1 U19974 ( .C1(n16780), .C2(P3_REIP_REG_9__SCAN_IN), .A(n16779), .B(
        n16778), .ZN(n16781) );
  OAI211_X1 U19975 ( .C1(n16784), .C2(n16783), .A(n16782), .B(n16781), .ZN(
        P3_U2662) );
  INV_X1 U19976 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n16795) );
  AOI211_X1 U19977 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16798), .A(n16785), .B(
        n16892), .ZN(n16793) );
  AOI21_X1 U19978 ( .B1(n16876), .B2(n16786), .A(P3_REIP_REG_8__SCAN_IN), .ZN(
        n16791) );
  AOI21_X1 U19979 ( .B1(n16788), .B2(n16802), .A(n16787), .ZN(n17758) );
  AND2_X1 U19980 ( .A1(n17757), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17768) );
  AOI21_X1 U19981 ( .B1(n17768), .B2(n16869), .A(n16852), .ZN(n16806) );
  XNOR2_X1 U19982 ( .A(n17758), .B(n16806), .ZN(n16789) );
  OAI22_X1 U19983 ( .A1(n16791), .A2(n16790), .B1(n18693), .B2(n16789), .ZN(
        n16792) );
  AOI211_X1 U19984 ( .C1(n16880), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16793), .B(n16792), .ZN(n16794) );
  OAI211_X1 U19985 ( .C1(n16893), .C2(n16795), .A(n16794), .B(n18169), .ZN(
        P3_U2663) );
  OAI21_X1 U19986 ( .B1(n16796), .B2(n16811), .A(n16862), .ZN(n16797) );
  INV_X1 U19987 ( .A(n16797), .ZN(n16799) );
  AOI22_X1 U19988 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n16880), .B1(
        n16799), .B2(n16798), .ZN(n16810) );
  NOR3_X1 U19989 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n16894), .A3(n16800), .ZN(
        n16801) );
  AOI211_X1 U19990 ( .C1(n16888), .C2(P3_EBX_REG_7__SCAN_IN), .A(n9736), .B(
        n16801), .ZN(n16809) );
  OAI21_X1 U19991 ( .B1(n16819), .B2(n16894), .A(n16897), .ZN(n16835) );
  NOR2_X1 U19992 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16894), .ZN(n16818) );
  OAI21_X1 U19993 ( .B1(n16835), .B2(n16818), .A(P3_REIP_REG_7__SCAN_IN), .ZN(
        n16808) );
  INV_X1 U19994 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17775) );
  NOR2_X1 U19995 ( .A1(n17849), .A2(n17787), .ZN(n16826) );
  NAND2_X1 U19996 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16826), .ZN(
        n16813) );
  INV_X1 U19997 ( .A(n16802), .ZN(n16803) );
  AOI21_X1 U19998 ( .B1(n17775), .B2(n16813), .A(n16803), .ZN(n17781) );
  NAND2_X1 U19999 ( .A1(n17757), .A2(n16869), .ZN(n16816) );
  AOI21_X1 U20000 ( .B1(n17781), .B2(n16816), .A(n18693), .ZN(n16804) );
  OAI22_X1 U20001 ( .A1(n17781), .A2(n16806), .B1(n16805), .B2(n16804), .ZN(
        n16807) );
  NAND4_X1 U20002 ( .A1(n16810), .A2(n16809), .A3(n16808), .A4(n16807), .ZN(
        P3_U2664) );
  AOI211_X1 U20003 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16829), .A(n16811), .B(
        n16892), .ZN(n16812) );
  AOI211_X1 U20004 ( .C1(n16888), .C2(P3_EBX_REG_6__SCAN_IN), .A(n9736), .B(
        n16812), .ZN(n16824) );
  INV_X1 U20005 ( .A(n16826), .ZN(n16814) );
  OAI21_X1 U20006 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16826), .A(
        n16813), .ZN(n17793) );
  AOI211_X1 U20007 ( .C1(n16815), .C2(n16814), .A(n16891), .B(n17793), .ZN(
        n16822) );
  AND2_X1 U20008 ( .A1(n17793), .A2(n16816), .ZN(n16817) );
  AOI22_X1 U20009 ( .A1(n16819), .A2(n16818), .B1(n16881), .B2(n16817), .ZN(
        n16820) );
  INV_X1 U20010 ( .A(n16820), .ZN(n16821) );
  AOI211_X1 U20011 ( .C1(n16835), .C2(P3_REIP_REG_6__SCAN_IN), .A(n16822), .B(
        n16821), .ZN(n16823) );
  OAI211_X1 U20012 ( .C1(n17788), .C2(n16868), .A(n16824), .B(n16823), .ZN(
        P3_U2665) );
  OAI21_X1 U20013 ( .B1(n16894), .B2(n16825), .A(n18722), .ZN(n16834) );
  INV_X1 U20014 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16832) );
  NAND2_X1 U20015 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17806), .ZN(
        n16838) );
  AOI21_X1 U20016 ( .B1(n16832), .B2(n16838), .A(n16826), .ZN(n17804) );
  AOI21_X1 U20017 ( .B1(n17806), .B2(n16869), .A(n16852), .ZN(n16839) );
  INV_X1 U20018 ( .A(n17804), .ZN(n16828) );
  INV_X1 U20019 ( .A(n16839), .ZN(n16827) );
  OAI221_X1 U20020 ( .B1(n17804), .B2(n16839), .C1(n16828), .C2(n16827), .A(
        n16853), .ZN(n16831) );
  OAI211_X1 U20021 ( .C1(n16841), .C2(n16837), .A(n16862), .B(n16829), .ZN(
        n16830) );
  OAI211_X1 U20022 ( .C1(n16868), .C2(n16832), .A(n16831), .B(n16830), .ZN(
        n16833) );
  AOI21_X1 U20023 ( .B1(n16835), .B2(n16834), .A(n16833), .ZN(n16836) );
  OAI211_X1 U20024 ( .C1(n16893), .C2(n16837), .A(n16836), .B(n18169), .ZN(
        P3_U2666) );
  NOR2_X1 U20025 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17809), .ZN(
        n17819) );
  NOR2_X1 U20026 ( .A1(n17849), .A2(n17809), .ZN(n16851) );
  OAI21_X1 U20027 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16851), .A(
        n16838), .ZN(n17816) );
  AOI22_X1 U20028 ( .A1(n16869), .A2(n17819), .B1(n16839), .B2(n17816), .ZN(
        n16849) );
  OAI21_X1 U20029 ( .B1(n16843), .B2(n16894), .A(n16897), .ZN(n16860) );
  NOR2_X1 U20030 ( .A1(n17377), .A2(n18846), .ZN(n16856) );
  OAI21_X1 U20031 ( .B1(n17118), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n16856), .ZN(n16840) );
  OAI211_X1 U20032 ( .C1(n17816), .C2(n16879), .A(n18169), .B(n16840), .ZN(
        n16847) );
  AOI211_X1 U20033 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16861), .A(n16841), .B(
        n16892), .ZN(n16842) );
  AOI21_X1 U20034 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n16888), .A(n16842), .ZN(
        n16845) );
  INV_X1 U20035 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20983) );
  NAND3_X1 U20036 ( .A1(n16876), .A2(n16843), .A3(n20983), .ZN(n16844) );
  OAI211_X1 U20037 ( .C1(n16868), .C2(n17821), .A(n16845), .B(n16844), .ZN(
        n16846) );
  AOI211_X1 U20038 ( .C1(P3_REIP_REG_4__SCAN_IN), .C2(n16860), .A(n16847), .B(
        n16846), .ZN(n16848) );
  OAI21_X1 U20039 ( .B1(n16849), .B2(n18693), .A(n16848), .ZN(P3_U2667) );
  INV_X1 U20040 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16865) );
  OAI21_X1 U20041 ( .B1(n16894), .B2(n16850), .A(n20931), .ZN(n16859) );
  NAND2_X1 U20042 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16866) );
  AOI21_X1 U20043 ( .B1(n16865), .B2(n16866), .A(n16851), .ZN(n17831) );
  NOR2_X1 U20044 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16866), .ZN(
        n16871) );
  NOR2_X1 U20045 ( .A1(n16871), .A2(n16852), .ZN(n16855) );
  OAI21_X1 U20046 ( .B1(n17831), .B2(n16855), .A(n16853), .ZN(n16854) );
  AOI21_X1 U20047 ( .B1(n17831), .B2(n16855), .A(n16854), .ZN(n16858) );
  NAND2_X1 U20048 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18635), .ZN(
        n18626) );
  AOI21_X1 U20049 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18626), .A(
        n17107), .ZN(n18788) );
  INV_X1 U20050 ( .A(n16856), .ZN(n18849) );
  OAI22_X1 U20051 ( .A1(n18788), .A2(n18849), .B1(n16893), .B2(n17201), .ZN(
        n16857) );
  AOI211_X1 U20052 ( .C1(n16860), .C2(n16859), .A(n16858), .B(n16857), .ZN(
        n16864) );
  OAI211_X1 U20053 ( .C1(n16867), .C2(n17201), .A(n16862), .B(n16861), .ZN(
        n16863) );
  OAI211_X1 U20054 ( .C1(n16868), .C2(n16865), .A(n16864), .B(n16863), .ZN(
        P3_U2668) );
  OAI21_X1 U20055 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16866), .ZN(n17839) );
  NAND2_X1 U20056 ( .A1(n16876), .A2(n18716), .ZN(n16883) );
  INV_X1 U20057 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18717) );
  AOI21_X1 U20058 ( .B1(n16897), .B2(n16883), .A(n18717), .ZN(n16875) );
  OR2_X1 U20059 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), .ZN(
        n16882) );
  AOI211_X1 U20060 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16882), .A(n16867), .B(
        n16892), .ZN(n16874) );
  INV_X1 U20061 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17842) );
  INV_X1 U20062 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17200) );
  OAI22_X1 U20063 ( .A1(n17842), .A2(n16868), .B1(n16893), .B2(n17200), .ZN(
        n16873) );
  OAI21_X1 U20064 ( .B1(n16869), .B2(n17839), .A(n16881), .ZN(n16870) );
  NOR2_X1 U20065 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18634), .ZN(
        n18629) );
  AOI21_X1 U20066 ( .B1(n18635), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n18629), .ZN(n18801) );
  INV_X1 U20067 ( .A(n18801), .ZN(n18638) );
  OAI22_X1 U20068 ( .A1(n16871), .A2(n16870), .B1(n18638), .B2(n18849), .ZN(
        n16872) );
  NOR4_X1 U20069 ( .A1(n16875), .A2(n16874), .A3(n16873), .A4(n16872), .ZN(
        n16878) );
  NAND3_X1 U20070 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16876), .A3(n18717), 
        .ZN(n16877) );
  OAI211_X1 U20071 ( .C1(n16879), .C2(n17839), .A(n16878), .B(n16877), .ZN(
        P3_U2669) );
  AOI21_X1 U20072 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16881), .A(
        n16880), .ZN(n16890) );
  NAND2_X1 U20073 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17206) );
  NAND2_X1 U20074 ( .A1(n16882), .A2(n17206), .ZN(n17214) );
  OAI21_X1 U20075 ( .B1(n16892), .B2(n17214), .A(n16883), .ZN(n16887) );
  NAND2_X1 U20076 ( .A1(n16885), .A2(n16884), .ZN(n18804) );
  OAI22_X1 U20077 ( .A1(n18716), .A2(n16897), .B1(n18804), .B2(n18849), .ZN(
        n16886) );
  AOI211_X1 U20078 ( .C1(n16888), .C2(P3_EBX_REG_1__SCAN_IN), .A(n16887), .B(
        n16886), .ZN(n16889) );
  OAI221_X1 U20079 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16891), .C1(
        n17849), .C2(n16890), .A(n16889), .ZN(P3_U2670) );
  NAND2_X1 U20080 ( .A1(n16893), .A2(n16892), .ZN(n16896) );
  NAND2_X1 U20081 ( .A1(n16894), .A2(n16897), .ZN(n16895) );
  AOI22_X1 U20082 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n16896), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n16895), .ZN(n16899) );
  NAND3_X1 U20083 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18845), .A3(
        n16897), .ZN(n16898) );
  OAI211_X1 U20084 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18849), .A(
        n16899), .B(n16898), .ZN(P3_U2671) );
  INV_X1 U20085 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16936) );
  NAND3_X1 U20086 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(P3_EBX_REG_17__SCAN_IN), 
        .A3(P3_EBX_REG_16__SCAN_IN), .ZN(n16900) );
  NOR2_X1 U20087 ( .A1(n17046), .A2(n16900), .ZN(n17006) );
  NAND3_X1 U20088 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(P3_EBX_REG_19__SCAN_IN), 
        .A3(n17006), .ZN(n16979) );
  NOR3_X1 U20089 ( .A1(n16936), .A2(n16901), .A3(n16979), .ZN(n16902) );
  NAND4_X1 U20090 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16903), .A3(n16937), 
        .A4(n16902), .ZN(n16906) );
  NOR2_X1 U20091 ( .A1(n16907), .A2(n16906), .ZN(n16932) );
  NAND2_X1 U20092 ( .A1(n17197), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16905) );
  NAND2_X1 U20093 ( .A1(n16932), .A2(n18222), .ZN(n16904) );
  OAI22_X1 U20094 ( .A1(n16932), .A2(n16905), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16904), .ZN(P3_U2672) );
  NAND2_X1 U20095 ( .A1(n16907), .A2(n16906), .ZN(n16908) );
  NAND2_X1 U20096 ( .A1(n16908), .A2(n17197), .ZN(n16931) );
  AOI22_X1 U20097 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16912) );
  AOI22_X1 U20098 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n15484), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16911) );
  AOI22_X1 U20099 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16910) );
  AOI22_X1 U20100 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16909) );
  NAND4_X1 U20101 ( .A1(n16912), .A2(n16911), .A3(n16910), .A4(n16909), .ZN(
        n16918) );
  AOI22_X1 U20102 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16916) );
  AOI22_X1 U20103 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16915) );
  AOI22_X1 U20104 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16914) );
  AOI22_X1 U20105 ( .A1(n9735), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16913) );
  NAND4_X1 U20106 ( .A1(n16916), .A2(n16915), .A3(n16914), .A4(n16913), .ZN(
        n16917) );
  OR2_X1 U20107 ( .A1(n16918), .A2(n16917), .ZN(n16934) );
  NAND3_X1 U20108 ( .A1(n16933), .A2(n16941), .A3(n16934), .ZN(n16930) );
  AOI22_X1 U20109 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n17154), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17166), .ZN(n16922) );
  AOI22_X1 U20110 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n17155), .ZN(n16921) );
  AOI22_X1 U20111 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n17165), .B1(
        P3_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n17171), .ZN(n16920) );
  AOI22_X1 U20112 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n17167), .ZN(n16919) );
  NAND4_X1 U20113 ( .A1(n16922), .A2(n16921), .A3(n16920), .A4(n16919), .ZN(
        n16928) );
  AOI22_X1 U20114 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16926) );
  AOI22_X1 U20115 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n9735), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16925) );
  AOI22_X1 U20116 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n9734), .ZN(n16924) );
  AOI22_X1 U20117 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n17080), .ZN(n16923) );
  NAND4_X1 U20118 ( .A1(n16926), .A2(n16925), .A3(n16924), .A4(n16923), .ZN(
        n16927) );
  NOR2_X1 U20119 ( .A1(n16928), .A2(n16927), .ZN(n16929) );
  XNOR2_X1 U20120 ( .A(n16930), .B(n16929), .ZN(n17228) );
  OAI22_X1 U20121 ( .A1(n16932), .A2(n16931), .B1(n17228), .B2(n17197), .ZN(
        P3_U2673) );
  NAND2_X1 U20122 ( .A1(n16933), .A2(n16941), .ZN(n16935) );
  XOR2_X1 U20123 ( .A(n16935), .B(n16934), .Z(n17233) );
  NAND4_X1 U20124 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16955), .A3(n16937), 
        .A4(n16936), .ZN(n16940) );
  NAND2_X1 U20125 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16938), .ZN(n16939) );
  OAI211_X1 U20126 ( .C1(n17197), .C2(n17233), .A(n16940), .B(n16939), .ZN(
        P3_U2674) );
  AOI21_X1 U20127 ( .B1(n16942), .B2(n16947), .A(n16941), .ZN(n17241) );
  NAND2_X1 U20128 ( .A1(n17216), .A2(n17241), .ZN(n16943) );
  OAI221_X1 U20129 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n16946), .C1(n16945), 
        .C2(n16944), .A(n16943), .ZN(P3_U2676) );
  INV_X1 U20130 ( .A(n16946), .ZN(n16951) );
  AOI21_X1 U20131 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17197), .A(n16955), .ZN(
        n16950) );
  OAI21_X1 U20132 ( .B1(n16949), .B2(n16948), .A(n16947), .ZN(n17247) );
  OAI22_X1 U20133 ( .A1(n16951), .A2(n16950), .B1(n17197), .B2(n17247), .ZN(
        P3_U2677) );
  INV_X1 U20134 ( .A(n16952), .ZN(n16961) );
  AOI21_X1 U20135 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17197), .A(n16961), .ZN(
        n16954) );
  XNOR2_X1 U20136 ( .A(n16953), .B(n16957), .ZN(n17252) );
  OAI22_X1 U20137 ( .A1(n16955), .A2(n16954), .B1(n17197), .B2(n17252), .ZN(
        P3_U2678) );
  NAND3_X1 U20138 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n16991), .ZN(n16962) );
  NOR2_X1 U20139 ( .A1(n16956), .A2(n16962), .ZN(n16966) );
  AOI21_X1 U20140 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17197), .A(n16966), .ZN(
        n16960) );
  OAI21_X1 U20141 ( .B1(n16959), .B2(n16958), .A(n16957), .ZN(n17257) );
  OAI22_X1 U20142 ( .A1(n16961), .A2(n16960), .B1(n17197), .B2(n17257), .ZN(
        P3_U2679) );
  INV_X1 U20143 ( .A(n16962), .ZN(n16978) );
  AOI21_X1 U20144 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17197), .A(n16978), .ZN(
        n16965) );
  XNOR2_X1 U20145 ( .A(n16964), .B(n16963), .ZN(n17262) );
  OAI22_X1 U20146 ( .A1(n16966), .A2(n16965), .B1(n17197), .B2(n17262), .ZN(
        P3_U2680) );
  AOI22_X1 U20147 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17197), .B1(
        P3_EBX_REG_21__SCAN_IN), .B2(n16991), .ZN(n16977) );
  AOI22_X1 U20148 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16970) );
  AOI22_X1 U20149 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16969) );
  AOI22_X1 U20150 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16968) );
  AOI22_X1 U20151 ( .A1(n17080), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16967) );
  NAND4_X1 U20152 ( .A1(n16970), .A2(n16969), .A3(n16968), .A4(n16967), .ZN(
        n16976) );
  AOI22_X1 U20153 ( .A1(n17107), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16974) );
  AOI22_X1 U20154 ( .A1(n17165), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16973) );
  AOI22_X1 U20155 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9735), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16972) );
  AOI22_X1 U20156 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16971) );
  NAND4_X1 U20157 ( .A1(n16974), .A2(n16973), .A3(n16972), .A4(n16971), .ZN(
        n16975) );
  NOR2_X1 U20158 ( .A1(n16976), .A2(n16975), .ZN(n17266) );
  OAI22_X1 U20159 ( .A1(n16978), .A2(n16977), .B1(n17266), .B2(n17197), .ZN(
        P3_U2681) );
  NAND2_X1 U20160 ( .A1(n17197), .A2(n16979), .ZN(n17004) );
  AOI22_X1 U20161 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16990) );
  AOI22_X1 U20162 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16989) );
  INV_X1 U20163 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20946) );
  AOI22_X1 U20164 ( .A1(n9735), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16980) );
  OAI21_X1 U20165 ( .B1(n16981), .B2(n20946), .A(n16980), .ZN(n16987) );
  AOI22_X1 U20166 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16985) );
  AOI22_X1 U20167 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16984) );
  AOI22_X1 U20168 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16983) );
  AOI22_X1 U20169 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16982) );
  NAND4_X1 U20170 ( .A1(n16985), .A2(n16984), .A3(n16983), .A4(n16982), .ZN(
        n16986) );
  AOI211_X1 U20171 ( .C1(n17124), .C2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        n16987), .B(n16986), .ZN(n16988) );
  NAND3_X1 U20172 ( .A1(n16990), .A2(n16989), .A3(n16988), .ZN(n17272) );
  AOI22_X1 U20173 ( .A1(n17216), .A2(n17272), .B1(n16991), .B2(n21016), .ZN(
        n16992) );
  OAI21_X1 U20174 ( .B1(n21016), .B2(n17004), .A(n16992), .ZN(P3_U2682) );
  AOI21_X1 U20175 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n16993), .A(
        P3_EBX_REG_20__SCAN_IN), .ZN(n17005) );
  AOI22_X1 U20176 ( .A1(n9735), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16997) );
  AOI22_X1 U20177 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16996) );
  AOI22_X1 U20178 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16995) );
  AOI22_X1 U20179 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16994) );
  NAND4_X1 U20180 ( .A1(n16997), .A2(n16996), .A3(n16995), .A4(n16994), .ZN(
        n17003) );
  AOI22_X1 U20181 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17001) );
  AOI22_X1 U20182 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17000) );
  AOI22_X1 U20183 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16999) );
  AOI22_X1 U20184 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16998) );
  NAND4_X1 U20185 ( .A1(n17001), .A2(n17000), .A3(n16999), .A4(n16998), .ZN(
        n17002) );
  NOR2_X1 U20186 ( .A1(n17003), .A2(n17002), .ZN(n17277) );
  OAI22_X1 U20187 ( .A1(n17005), .A2(n17004), .B1(n17277), .B2(n17197), .ZN(
        P3_U2683) );
  NOR2_X1 U20188 ( .A1(n17216), .A2(n17006), .ZN(n17030) );
  AOI22_X1 U20189 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17017) );
  AOI22_X1 U20190 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17016) );
  INV_X1 U20191 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n20952) );
  AOI22_X1 U20192 ( .A1(n9735), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17007) );
  OAI21_X1 U20193 ( .B1(n17008), .B2(n20952), .A(n17007), .ZN(n17014) );
  AOI22_X1 U20194 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17012) );
  AOI22_X1 U20195 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17011) );
  AOI22_X1 U20196 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17010) );
  AOI22_X1 U20197 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17009) );
  NAND4_X1 U20198 ( .A1(n17012), .A2(n17011), .A3(n17010), .A4(n17009), .ZN(
        n17013) );
  AOI211_X1 U20199 ( .C1(n17166), .C2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A(
        n17014), .B(n17013), .ZN(n17015) );
  NAND3_X1 U20200 ( .A1(n17017), .A2(n17016), .A3(n17015), .ZN(n17281) );
  AOI22_X1 U20201 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17030), .B1(n17216), 
        .B2(n17281), .ZN(n17018) );
  OAI21_X1 U20202 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17019), .A(n17018), .ZN(
        P3_U2684) );
  NAND3_X1 U20203 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(P3_EBX_REG_16__SCAN_IN), 
        .A3(n17059), .ZN(n17032) );
  AOI22_X1 U20204 ( .A1(n9735), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17029) );
  AOI22_X1 U20205 ( .A1(n17080), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17028) );
  AOI22_X1 U20206 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17020) );
  OAI21_X1 U20207 ( .B1(n17169), .B2(n20967), .A(n17020), .ZN(n17026) );
  AOI22_X1 U20208 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17024) );
  AOI22_X1 U20209 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17023) );
  AOI22_X1 U20210 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17022) );
  AOI22_X1 U20211 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17021) );
  NAND4_X1 U20212 ( .A1(n17024), .A2(n17023), .A3(n17022), .A4(n17021), .ZN(
        n17025) );
  AOI211_X1 U20213 ( .C1(n17047), .C2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A(
        n17026), .B(n17025), .ZN(n17027) );
  NAND3_X1 U20214 ( .A1(n17029), .A2(n17028), .A3(n17027), .ZN(n17285) );
  AOI22_X1 U20215 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17030), .B1(n17216), 
        .B2(n17285), .ZN(n17031) );
  OAI21_X1 U20216 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17032), .A(n17031), .ZN(
        P3_U2685) );
  INV_X1 U20217 ( .A(n17032), .ZN(n17045) );
  AOI22_X1 U20218 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17197), .B1(
        P3_EBX_REG_16__SCAN_IN), .B2(n17059), .ZN(n17044) );
  AOI22_X1 U20219 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9735), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17036) );
  AOI22_X1 U20220 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17035) );
  AOI22_X1 U20221 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17034) );
  AOI22_X1 U20222 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17033) );
  NAND4_X1 U20223 ( .A1(n17036), .A2(n17035), .A3(n17034), .A4(n17033), .ZN(
        n17043) );
  AOI22_X1 U20224 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17041) );
  AOI22_X1 U20225 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17040) );
  AOI22_X1 U20226 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17039) );
  AOI22_X1 U20227 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17038) );
  NAND4_X1 U20228 ( .A1(n17041), .A2(n17040), .A3(n17039), .A4(n17038), .ZN(
        n17042) );
  NOR2_X1 U20229 ( .A1(n17043), .A2(n17042), .ZN(n17295) );
  OAI22_X1 U20230 ( .A1(n17045), .A2(n17044), .B1(n17295), .B2(n17197), .ZN(
        P3_U2686) );
  INV_X1 U20231 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17061) );
  NAND2_X1 U20232 ( .A1(n17197), .A2(n17046), .ZN(n17072) );
  AOI22_X1 U20233 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17047), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17058) );
  AOI22_X1 U20234 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17057) );
  INV_X1 U20235 ( .A(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n20966) );
  AOI22_X1 U20236 ( .A1(n9735), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17048) );
  OAI21_X1 U20237 ( .B1(n9783), .B2(n20966), .A(n17048), .ZN(n17055) );
  AOI22_X1 U20238 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17053) );
  AOI22_X1 U20239 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17052) );
  AOI22_X1 U20240 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17051) );
  AOI22_X1 U20241 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17050) );
  NAND4_X1 U20242 ( .A1(n17053), .A2(n17052), .A3(n17051), .A4(n17050), .ZN(
        n17054) );
  AOI211_X1 U20243 ( .C1(n17075), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n17055), .B(n17054), .ZN(n17056) );
  NAND3_X1 U20244 ( .A1(n17058), .A2(n17057), .A3(n17056), .ZN(n17296) );
  AOI22_X1 U20245 ( .A1(n17216), .A2(n17296), .B1(n17059), .B2(n17061), .ZN(
        n17060) );
  OAI21_X1 U20246 ( .B1(n17061), .B2(n17072), .A(n17060), .ZN(P3_U2687) );
  NOR2_X1 U20247 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17088), .ZN(n17073) );
  AOI22_X1 U20248 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17154), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17065) );
  AOI22_X1 U20249 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17064) );
  AOI22_X1 U20250 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17118), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17063) );
  AOI22_X1 U20251 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n17089), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17049), .ZN(n17062) );
  NAND4_X1 U20252 ( .A1(n17065), .A2(n17064), .A3(n17063), .A4(n17062), .ZN(
        n17071) );
  AOI22_X1 U20253 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n17124), .ZN(n17069) );
  AOI22_X1 U20254 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17165), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17068) );
  AOI22_X1 U20255 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n9735), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n9734), .ZN(n17067) );
  AOI22_X1 U20256 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17066) );
  NAND4_X1 U20257 ( .A1(n17069), .A2(n17068), .A3(n17067), .A4(n17066), .ZN(
        n17070) );
  NOR2_X1 U20258 ( .A1(n17071), .A2(n17070), .ZN(n17305) );
  OAI22_X1 U20259 ( .A1(n17073), .A2(n17072), .B1(n17305), .B2(n17197), .ZN(
        P3_U2688) );
  OAI21_X1 U20260 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17074), .A(n17197), .ZN(
        n17087) );
  AOI22_X1 U20261 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17079) );
  AOI22_X1 U20262 ( .A1(n9735), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17078) );
  AOI22_X1 U20263 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17077) );
  AOI22_X1 U20264 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17076) );
  NAND4_X1 U20265 ( .A1(n17079), .A2(n17078), .A3(n17077), .A4(n17076), .ZN(
        n17086) );
  AOI22_X1 U20266 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17084) );
  AOI22_X1 U20267 ( .A1(n17080), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17083) );
  AOI22_X1 U20268 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17082) );
  AOI22_X1 U20269 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17081) );
  NAND4_X1 U20270 ( .A1(n17084), .A2(n17083), .A3(n17082), .A4(n17081), .ZN(
        n17085) );
  NOR2_X1 U20271 ( .A1(n17086), .A2(n17085), .ZN(n17310) );
  OAI22_X1 U20272 ( .A1(n17088), .A2(n17087), .B1(n17310), .B2(n17197), .ZN(
        P3_U2689) );
  AOI22_X1 U20273 ( .A1(n17047), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17093) );
  AOI22_X1 U20274 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17092) );
  AOI22_X1 U20275 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17091) );
  AOI22_X1 U20276 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17090) );
  NAND4_X1 U20277 ( .A1(n17093), .A2(n17092), .A3(n17091), .A4(n17090), .ZN(
        n17099) );
  AOI22_X1 U20278 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17097) );
  AOI22_X1 U20279 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17096) );
  AOI22_X1 U20280 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17095) );
  AOI22_X1 U20281 ( .A1(n9735), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17094) );
  NAND4_X1 U20282 ( .A1(n17097), .A2(n17096), .A3(n17095), .A4(n17094), .ZN(
        n17098) );
  NOR2_X1 U20283 ( .A1(n17099), .A2(n17098), .ZN(n17311) );
  OAI21_X1 U20284 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17101), .A(n17100), .ZN(
        n17102) );
  AOI22_X1 U20285 ( .A1(n17216), .A2(n17311), .B1(n17102), .B2(n17197), .ZN(
        P3_U2690) );
  AOI22_X1 U20286 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17106) );
  AOI22_X1 U20287 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17105) );
  AOI22_X1 U20288 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17104) );
  AOI22_X1 U20289 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17103) );
  NAND4_X1 U20290 ( .A1(n17106), .A2(n17105), .A3(n17104), .A4(n17103), .ZN(
        n17113) );
  AOI22_X1 U20291 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17107), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17111) );
  AOI22_X1 U20292 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17110) );
  AOI22_X1 U20293 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17109) );
  AOI22_X1 U20294 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9735), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17108) );
  NAND4_X1 U20295 ( .A1(n17111), .A2(n17110), .A3(n17109), .A4(n17108), .ZN(
        n17112) );
  NOR2_X1 U20296 ( .A1(n17113), .A2(n17112), .ZN(n17315) );
  INV_X1 U20297 ( .A(n17131), .ZN(n17114) );
  OAI33_X1 U20298 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17263), .A3(n17131), 
        .B1(n17115), .B2(n17216), .B3(n17114), .ZN(n17116) );
  INV_X1 U20299 ( .A(n17116), .ZN(n17117) );
  OAI21_X1 U20300 ( .B1(n17315), .B2(n17197), .A(n17117), .ZN(P3_U2691) );
  AOI22_X1 U20301 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17122) );
  AOI22_X1 U20302 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17121) );
  AOI22_X1 U20303 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17120) );
  AOI22_X1 U20304 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17119) );
  NAND4_X1 U20305 ( .A1(n17122), .A2(n17121), .A3(n17120), .A4(n17119), .ZN(
        n17130) );
  AOI22_X1 U20306 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9735), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17128) );
  AOI22_X1 U20307 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17127) );
  AOI22_X1 U20308 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17126) );
  AOI22_X1 U20309 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17123), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17125) );
  NAND4_X1 U20310 ( .A1(n17128), .A2(n17127), .A3(n17126), .A4(n17125), .ZN(
        n17129) );
  NOR2_X1 U20311 ( .A1(n17130), .A2(n17129), .ZN(n17320) );
  OAI211_X1 U20312 ( .C1(P3_EBX_REG_11__SCAN_IN), .C2(n17145), .A(n17131), .B(
        n17197), .ZN(n17132) );
  OAI21_X1 U20313 ( .B1(n17320), .B2(n17197), .A(n17132), .ZN(P3_U2692) );
  OAI21_X1 U20314 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17133), .A(n17197), .ZN(
        n17144) );
  AOI22_X1 U20315 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17137) );
  AOI22_X1 U20316 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17136) );
  AOI22_X1 U20317 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17135) );
  AOI22_X1 U20318 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17134) );
  NAND4_X1 U20319 ( .A1(n17137), .A2(n17136), .A3(n17135), .A4(n17134), .ZN(
        n17143) );
  AOI22_X1 U20320 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17141) );
  AOI22_X1 U20321 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17140) );
  AOI22_X1 U20322 ( .A1(n9735), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17139) );
  AOI22_X1 U20323 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17138) );
  NAND4_X1 U20324 ( .A1(n17141), .A2(n17140), .A3(n17139), .A4(n17138), .ZN(
        n17142) );
  NOR2_X1 U20325 ( .A1(n17143), .A2(n17142), .ZN(n17329) );
  OAI22_X1 U20326 ( .A1(n17145), .A2(n17144), .B1(n17329), .B2(n17197), .ZN(
        P3_U2693) );
  AOI22_X1 U20327 ( .A1(n17146), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17152) );
  AOI22_X1 U20328 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17151) );
  AOI22_X1 U20329 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17150) );
  AOI22_X1 U20330 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17167), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17149) );
  NAND4_X1 U20331 ( .A1(n17152), .A2(n17151), .A3(n17150), .A4(n17149), .ZN(
        n17162) );
  AOI22_X1 U20332 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17160) );
  AOI22_X1 U20333 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9735), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17159) );
  AOI22_X1 U20334 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17158) );
  AOI22_X1 U20335 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17157) );
  NAND4_X1 U20336 ( .A1(n17160), .A2(n17159), .A3(n17158), .A4(n17157), .ZN(
        n17161) );
  NOR2_X1 U20337 ( .A1(n17162), .A2(n17161), .ZN(n17330) );
  OAI21_X1 U20338 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17183), .A(n17163), .ZN(
        n17164) );
  AOI22_X1 U20339 ( .A1(n17216), .A2(n17330), .B1(n17164), .B2(n17197), .ZN(
        P3_U2694) );
  OAI21_X1 U20340 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17186), .A(n17197), .ZN(
        n17182) );
  AOI22_X1 U20341 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17180) );
  AOI22_X1 U20342 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17179) );
  INV_X1 U20343 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n21014) );
  AOI22_X1 U20344 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17168) );
  OAI21_X1 U20345 ( .B1(n17169), .B2(n21014), .A(n17168), .ZN(n17177) );
  AOI22_X1 U20346 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9735), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17175) );
  AOI22_X1 U20347 ( .A1(n17170), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17174) );
  AOI22_X1 U20348 ( .A1(n17123), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n15484), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17173) );
  AOI22_X1 U20349 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17172) );
  NAND4_X1 U20350 ( .A1(n17175), .A2(n17174), .A3(n17173), .A4(n17172), .ZN(
        n17176) );
  AOI211_X1 U20351 ( .C1(n17124), .C2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n17177), .B(n17176), .ZN(n17178) );
  NAND3_X1 U20352 ( .A1(n17180), .A2(n17179), .A3(n17178), .ZN(n17334) );
  INV_X1 U20353 ( .A(n17334), .ZN(n17181) );
  OAI22_X1 U20354 ( .A1(n17183), .A2(n17182), .B1(n17181), .B2(n17197), .ZN(
        P3_U2695) );
  NOR2_X1 U20355 ( .A1(n17263), .A2(n17187), .ZN(n17189) );
  AOI22_X1 U20356 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17197), .B1(
        P3_EBX_REG_6__SCAN_IN), .B2(n17189), .ZN(n17185) );
  OAI22_X1 U20357 ( .A1(n17186), .A2(n17185), .B1(n17184), .B2(n17197), .ZN(
        P3_U2696) );
  AND2_X1 U20358 ( .A1(n17197), .A2(n17187), .ZN(n17192) );
  AOI22_X1 U20359 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17192), .B1(n17189), .B2(
        n17188), .ZN(n17190) );
  OAI21_X1 U20360 ( .B1(n17191), .B2(n17197), .A(n17190), .ZN(P3_U2697) );
  OAI21_X1 U20361 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17193), .A(n17192), .ZN(
        n17194) );
  OAI21_X1 U20362 ( .B1(n17197), .B2(n20946), .A(n17194), .ZN(P3_U2698) );
  INV_X1 U20363 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17199) );
  OAI21_X1 U20364 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17196), .A(n17195), .ZN(
        n17198) );
  AOI22_X1 U20365 ( .A1(n17216), .A2(n17199), .B1(n17198), .B2(n17197), .ZN(
        P3_U2699) );
  INV_X1 U20366 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17205) );
  NOR3_X1 U20367 ( .A1(n17200), .A2(n17206), .A3(n17218), .ZN(n17208) );
  NOR2_X1 U20368 ( .A1(n17216), .A2(n17201), .ZN(n17203) );
  OAI22_X1 U20369 ( .A1(n17208), .A2(n17203), .B1(n17202), .B2(n17218), .ZN(
        n17204) );
  OAI21_X1 U20370 ( .B1(n17197), .B2(n17205), .A(n17204), .ZN(P3_U2700) );
  INV_X1 U20371 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17210) );
  INV_X1 U20372 ( .A(n17206), .ZN(n17207) );
  AOI221_X1 U20373 ( .B1(n17207), .B2(n17212), .C1(n17263), .C2(n17212), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17209) );
  AOI211_X1 U20374 ( .C1(n17216), .C2(n17210), .A(n17209), .B(n17208), .ZN(
        P3_U2701) );
  INV_X1 U20375 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17213) );
  INV_X1 U20376 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17211) );
  OAI222_X1 U20377 ( .A1(n17214), .A2(n17218), .B1(n17213), .B2(n17212), .C1(
        n17211), .C2(n17197), .ZN(P3_U2702) );
  AOI22_X1 U20378 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17216), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17215), .ZN(n17217) );
  OAI21_X1 U20379 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17218), .A(n17217), .ZN(
        P3_U2703) );
  INV_X1 U20380 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17444) );
  INV_X1 U20381 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17440) );
  INV_X1 U20382 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17436) );
  INV_X1 U20383 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17483) );
  NAND2_X1 U20384 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n17370) );
  NAND3_X1 U20385 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .ZN(n17341) );
  NOR2_X1 U20386 ( .A1(n17370), .A2(n17341), .ZN(n17219) );
  NAND4_X1 U20387 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(P3_EAX_REG_7__SCAN_IN), 
        .A3(P3_EAX_REG_6__SCAN_IN), .A4(n17219), .ZN(n17339) );
  NOR2_X1 U20388 ( .A1(n17368), .A2(n17339), .ZN(n17333) );
  INV_X1 U20389 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17468) );
  INV_X1 U20390 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17466) );
  INV_X1 U20391 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17464) );
  NAND2_X1 U20392 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .ZN(n17306) );
  NOR4_X1 U20393 ( .A1(n17468), .A2(n17466), .A3(n17464), .A4(n17306), .ZN(
        n17220) );
  NAND4_X1 U20394 ( .A1(n17333), .A2(P3_EAX_REG_14__SCAN_IN), .A3(
        P3_EAX_REG_13__SCAN_IN), .A4(n17220), .ZN(n17307) );
  NAND2_X1 U20395 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17302), .ZN(n17298) );
  NAND2_X1 U20396 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .ZN(n17264) );
  NAND4_X1 U20397 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_21__SCAN_IN), 
        .A3(P3_EAX_REG_20__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n17221)
         );
  NAND2_X1 U20398 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17259), .ZN(n17258) );
  NOR2_X1 U20399 ( .A1(n17263), .A2(n17258), .ZN(n17254) );
  NAND2_X1 U20400 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17254), .ZN(n17253) );
  NAND2_X1 U20401 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17248), .ZN(n17244) );
  NAND2_X1 U20402 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17238), .ZN(n17234) );
  NOR2_X2 U20403 ( .A1(n17444), .A2(n17234), .ZN(n17229) );
  NAND2_X1 U20404 ( .A1(n17229), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17225) );
  NAND2_X1 U20405 ( .A1(n17222), .A2(n17325), .ZN(n17301) );
  OAI22_X1 U20406 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17340), .B1(n17325), 
        .B2(n17229), .ZN(n17223) );
  AOI22_X1 U20407 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17290), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17223), .ZN(n17224) );
  OAI21_X1 U20408 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17225), .A(n17224), .ZN(
        P3_U2704) );
  NAND2_X1 U20409 ( .A1(n18210), .A2(n17325), .ZN(n17271) );
  AOI22_X1 U20410 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n17290), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n17297), .ZN(n17227) );
  OAI211_X1 U20411 ( .C1(n17229), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17362), .B(
        n17225), .ZN(n17226) );
  OAI211_X1 U20412 ( .C1(n17228), .C2(n17374), .A(n17227), .B(n17226), .ZN(
        P3_U2705) );
  AOI22_X1 U20413 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n17290), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n17297), .ZN(n17232) );
  AOI211_X1 U20414 ( .C1(n17444), .C2(n17234), .A(n17229), .B(n17325), .ZN(
        n17230) );
  INV_X1 U20415 ( .A(n17230), .ZN(n17231) );
  OAI211_X1 U20416 ( .C1(n17374), .C2(n17233), .A(n17232), .B(n17231), .ZN(
        P3_U2706) );
  AOI22_X1 U20417 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n17290), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n17297), .ZN(n17236) );
  OAI211_X1 U20418 ( .C1(n17238), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17362), .B(
        n17234), .ZN(n17235) );
  OAI211_X1 U20419 ( .C1(n17374), .C2(n17237), .A(n17236), .B(n17235), .ZN(
        P3_U2707) );
  INV_X1 U20420 ( .A(n17238), .ZN(n17240) );
  OAI21_X1 U20421 ( .B1(n17325), .B2(n17440), .A(n17244), .ZN(n17239) );
  AOI22_X1 U20422 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n17290), .B1(n17240), .B2(
        n17239), .ZN(n17243) );
  AOI22_X1 U20423 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17297), .B1(n17241), .B2(
        n17335), .ZN(n17242) );
  NAND2_X1 U20424 ( .A1(n17243), .A2(n17242), .ZN(P3_U2708) );
  AOI22_X1 U20425 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n17290), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n17297), .ZN(n17246) );
  OAI211_X1 U20426 ( .C1(n17248), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17362), .B(
        n17244), .ZN(n17245) );
  OAI211_X1 U20427 ( .C1(n17247), .C2(n17374), .A(n17246), .B(n17245), .ZN(
        P3_U2709) );
  AOI22_X1 U20428 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n17290), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n17297), .ZN(n17251) );
  AOI211_X1 U20429 ( .C1(n17436), .C2(n17253), .A(n17248), .B(n17325), .ZN(
        n17249) );
  INV_X1 U20430 ( .A(n17249), .ZN(n17250) );
  OAI211_X1 U20431 ( .C1(n17252), .C2(n17374), .A(n17251), .B(n17250), .ZN(
        P3_U2710) );
  AOI22_X1 U20432 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n17290), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n17297), .ZN(n17256) );
  OAI211_X1 U20433 ( .C1(n17254), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17362), .B(
        n17253), .ZN(n17255) );
  OAI211_X1 U20434 ( .C1(n17374), .C2(n17257), .A(n17256), .B(n17255), .ZN(
        P3_U2711) );
  AOI22_X1 U20435 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n17290), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n17297), .ZN(n17261) );
  OAI211_X1 U20436 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17259), .A(n17362), .B(
        n17258), .ZN(n17260) );
  OAI211_X1 U20437 ( .C1(n17262), .C2(n17374), .A(n17261), .B(n17260), .ZN(
        P3_U2712) );
  INV_X1 U20438 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18214) );
  INV_X1 U20439 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17426) );
  NOR2_X1 U20440 ( .A1(n17263), .A2(n17298), .ZN(n17292) );
  NAND2_X1 U20441 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17292), .ZN(n17291) );
  NOR2_X1 U20442 ( .A1(n17426), .A2(n17282), .ZN(n17273) );
  INV_X1 U20443 ( .A(n17273), .ZN(n17265) );
  NAND2_X1 U20444 ( .A1(n17362), .A2(n17265), .ZN(n17280) );
  OAI21_X1 U20445 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17340), .A(n17280), .ZN(
        n17269) );
  INV_X1 U20446 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17428) );
  NOR3_X1 U20447 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17428), .A3(n17265), .ZN(
        n17268) );
  OAI22_X1 U20448 ( .A1(n17266), .A2(n17374), .B1(n18213), .B2(n17301), .ZN(
        n17267) );
  AOI211_X1 U20449 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n17269), .A(n17268), .B(
        n17267), .ZN(n17270) );
  OAI21_X1 U20450 ( .B1(n18214), .B2(n17271), .A(n17270), .ZN(P3_U2713) );
  AOI22_X1 U20451 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n17290), .B1(n17335), .B2(
        n17272), .ZN(n17275) );
  AOI22_X1 U20452 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17297), .B1(n17273), .B2(
        n17428), .ZN(n17274) );
  OAI211_X1 U20453 ( .C1(n17428), .C2(n17280), .A(n17275), .B(n17274), .ZN(
        P3_U2714) );
  OAI22_X1 U20454 ( .A1(n17277), .A2(n17374), .B1(n17276), .B2(n17301), .ZN(
        n17278) );
  AOI21_X1 U20455 ( .B1(BUF2_REG_4__SCAN_IN), .B2(n17297), .A(n17278), .ZN(
        n17279) );
  OAI221_X1 U20456 ( .B1(P3_EAX_REG_20__SCAN_IN), .B2(n17282), .C1(n17426), 
        .C2(n17280), .A(n17279), .ZN(P3_U2715) );
  INV_X1 U20457 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n18202) );
  AOI22_X1 U20458 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17297), .B1(n17335), .B2(
        n17281), .ZN(n17284) );
  INV_X1 U20459 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17422) );
  NOR2_X1 U20460 ( .A1(n17422), .A2(n17291), .ZN(n17286) );
  OAI211_X1 U20461 ( .C1(n17286), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17362), .B(
        n17282), .ZN(n17283) );
  OAI211_X1 U20462 ( .C1(n17301), .C2(n18202), .A(n17284), .B(n17283), .ZN(
        P3_U2716) );
  AOI22_X1 U20463 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17297), .B1(n17335), .B2(
        n17285), .ZN(n17289) );
  AOI211_X1 U20464 ( .C1(n17422), .C2(n17291), .A(n17286), .B(n17325), .ZN(
        n17287) );
  INV_X1 U20465 ( .A(n17287), .ZN(n17288) );
  OAI211_X1 U20466 ( .C1(n17301), .C2(n18195), .A(n17289), .B(n17288), .ZN(
        P3_U2717) );
  AOI22_X1 U20467 ( .A1(BUF2_REG_17__SCAN_IN), .A2(n17290), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n17297), .ZN(n17294) );
  OAI211_X1 U20468 ( .C1(n17292), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17362), .B(
        n17291), .ZN(n17293) );
  OAI211_X1 U20469 ( .C1(n17295), .C2(n17374), .A(n17294), .B(n17293), .ZN(
        P3_U2718) );
  INV_X1 U20470 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n19050) );
  AOI22_X1 U20471 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17297), .B1(n17335), .B2(
        n17296), .ZN(n17300) );
  OAI211_X1 U20472 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17302), .A(n17362), .B(
        n17298), .ZN(n17299) );
  OAI211_X1 U20473 ( .C1(n17301), .C2(n19050), .A(n17300), .B(n17299), .ZN(
        P3_U2719) );
  AOI211_X1 U20474 ( .C1(n17483), .C2(n17307), .A(n17325), .B(n17302), .ZN(
        n17303) );
  AOI21_X1 U20475 ( .B1(n17369), .B2(BUF2_REG_15__SCAN_IN), .A(n17303), .ZN(
        n17304) );
  OAI21_X1 U20476 ( .B1(n17305), .B2(n17374), .A(n17304), .ZN(P3_U2720) );
  NAND2_X1 U20477 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17338), .ZN(n17326) );
  INV_X1 U20478 ( .A(n17326), .ZN(n17332) );
  NAND2_X1 U20479 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17332), .ZN(n17319) );
  NOR2_X1 U20480 ( .A1(n17306), .A2(n17319), .ZN(n17317) );
  AND2_X1 U20481 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17317), .ZN(n17313) );
  INV_X1 U20482 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17478) );
  AOI22_X1 U20483 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17369), .B1(n17313), .B2(
        n17478), .ZN(n17309) );
  NAND3_X1 U20484 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17362), .A3(n17307), 
        .ZN(n17308) );
  OAI211_X1 U20485 ( .C1(n17310), .C2(n17374), .A(n17309), .B(n17308), .ZN(
        P3_U2721) );
  INV_X1 U20486 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17314) );
  AOI21_X1 U20487 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17362), .A(n17317), .ZN(
        n17312) );
  OAI222_X1 U20488 ( .A1(n17367), .A2(n17314), .B1(n17313), .B2(n17312), .C1(
        n17374), .C2(n17311), .ZN(P3_U2722) );
  INV_X1 U20489 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17318) );
  INV_X1 U20490 ( .A(n17319), .ZN(n17324) );
  AOI22_X1 U20491 ( .A1(n17324), .A2(P3_EAX_REG_11__SCAN_IN), .B1(
        P3_EAX_REG_12__SCAN_IN), .B2(n17362), .ZN(n17316) );
  OAI222_X1 U20492 ( .A1(n17367), .A2(n17318), .B1(n17317), .B2(n17316), .C1(
        n17374), .C2(n17315), .ZN(P3_U2723) );
  INV_X1 U20493 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17323) );
  INV_X1 U20494 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17471) );
  NOR2_X1 U20495 ( .A1(n17471), .A2(n17319), .ZN(n17322) );
  AOI21_X1 U20496 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17362), .A(n17324), .ZN(
        n17321) );
  OAI222_X1 U20497 ( .A1(n17367), .A2(n17323), .B1(n17322), .B2(n17321), .C1(
        n17374), .C2(n17320), .ZN(P3_U2724) );
  AOI211_X1 U20498 ( .C1(n17468), .C2(n17326), .A(n17325), .B(n17324), .ZN(
        n17327) );
  AOI21_X1 U20499 ( .B1(n17369), .B2(BUF2_REG_10__SCAN_IN), .A(n17327), .ZN(
        n17328) );
  OAI21_X1 U20500 ( .B1(n17329), .B2(n17374), .A(n17328), .ZN(P3_U2725) );
  INV_X1 U20501 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n20999) );
  AOI21_X1 U20502 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17362), .A(n17338), .ZN(
        n17331) );
  OAI222_X1 U20503 ( .A1(n17367), .A2(n20999), .B1(n17332), .B2(n17331), .C1(
        n17374), .C2(n17330), .ZN(P3_U2726) );
  OAI21_X1 U20504 ( .B1(n17333), .B2(P3_EAX_REG_8__SCAN_IN), .A(n17362), .ZN(
        n17337) );
  AOI22_X1 U20505 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17369), .B1(n17335), .B2(
        n17334), .ZN(n17336) );
  OAI21_X1 U20506 ( .B1(n17338), .B2(n17337), .A(n17336), .ZN(P3_U2727) );
  INV_X1 U20507 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18218) );
  NOR2_X1 U20508 ( .A1(n17339), .A2(n17340), .ZN(n17344) );
  NOR2_X1 U20509 ( .A1(n17370), .A2(n17340), .ZN(n17361) );
  NAND2_X1 U20510 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17361), .ZN(n17357) );
  NOR2_X1 U20511 ( .A1(n17341), .A2(n17357), .ZN(n17352) );
  AOI22_X1 U20512 ( .A1(n17352), .A2(P3_EAX_REG_6__SCAN_IN), .B1(
        P3_EAX_REG_7__SCAN_IN), .B2(n17362), .ZN(n17343) );
  OAI222_X1 U20513 ( .A1(n17367), .A2(n18218), .B1(n17344), .B2(n17343), .C1(
        n17374), .C2(n17342), .ZN(P3_U2728) );
  AOI21_X1 U20514 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17362), .A(n17352), .ZN(
        n17348) );
  AND2_X1 U20515 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17352), .ZN(n17347) );
  INV_X1 U20516 ( .A(n17345), .ZN(n17346) );
  OAI222_X1 U20517 ( .A1(n17367), .A2(n18214), .B1(n17348), .B2(n17347), .C1(
        n17374), .C2(n17346), .ZN(P3_U2729) );
  INV_X1 U20518 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18209) );
  NAND2_X1 U20519 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .ZN(n17349) );
  NOR2_X1 U20520 ( .A1(n17349), .A2(n17357), .ZN(n17356) );
  AOI21_X1 U20521 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17362), .A(n17356), .ZN(
        n17351) );
  OAI222_X1 U20522 ( .A1(n18209), .A2(n17367), .B1(n17352), .B2(n17351), .C1(
        n17374), .C2(n17350), .ZN(P3_U2730) );
  INV_X1 U20523 ( .A(n17357), .ZN(n17366) );
  AOI22_X1 U20524 ( .A1(n17366), .A2(P3_EAX_REG_3__SCAN_IN), .B1(
        P3_EAX_REG_4__SCAN_IN), .B2(n17362), .ZN(n17355) );
  INV_X1 U20525 ( .A(n17353), .ZN(n17354) );
  OAI222_X1 U20526 ( .A1(n18205), .A2(n17367), .B1(n17356), .B2(n17355), .C1(
        n17374), .C2(n17354), .ZN(P3_U2731) );
  INV_X1 U20527 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17454) );
  NOR2_X1 U20528 ( .A1(n17454), .A2(n17357), .ZN(n17360) );
  AOI21_X1 U20529 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17362), .A(n17366), .ZN(
        n17359) );
  OAI222_X1 U20530 ( .A1(n18201), .A2(n17367), .B1(n17360), .B2(n17359), .C1(
        n17374), .C2(n17358), .ZN(P3_U2732) );
  INV_X1 U20531 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18196) );
  AOI21_X1 U20532 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17362), .A(n17361), .ZN(
        n17365) );
  INV_X1 U20533 ( .A(n17363), .ZN(n17364) );
  OAI222_X1 U20534 ( .A1(n18196), .A2(n17367), .B1(n17366), .B2(n17365), .C1(
        n17374), .C2(n17364), .ZN(P3_U2733) );
  AOI22_X1 U20535 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17369), .B1(
        P3_EAX_REG_1__SCAN_IN), .B2(n17368), .ZN(n17373) );
  OAI211_X1 U20536 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(P3_EAX_REG_0__SCAN_IN), 
        .A(n17371), .B(n17370), .ZN(n17372) );
  OAI211_X1 U20537 ( .C1(n17375), .C2(n17374), .A(n17373), .B(n17372), .ZN(
        P3_U2734) );
  NOR2_X2 U20538 ( .A1(n20974), .A2(n17856), .ZN(n18832) );
  NOR2_X4 U20539 ( .A1(n18832), .A2(n17394), .ZN(n17409) );
  AND2_X1 U20540 ( .A1(n17409), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20541 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17446) );
  CLKBUF_X1 U20542 ( .A(n18832), .Z(n17410) );
  AOI22_X1 U20543 ( .A1(n17410), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17378) );
  OAI21_X1 U20544 ( .B1(n17446), .B2(n17393), .A(n17378), .ZN(P3_U2737) );
  AOI22_X1 U20545 ( .A1(n17410), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17379) );
  OAI21_X1 U20546 ( .B1(n17444), .B2(n17393), .A(n17379), .ZN(P3_U2738) );
  INV_X1 U20547 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17442) );
  AOI22_X1 U20548 ( .A1(P3_DATAO_REG_28__SCAN_IN), .A2(n17409), .B1(n18832), 
        .B2(P3_UWORD_REG_12__SCAN_IN), .ZN(n17380) );
  OAI21_X1 U20549 ( .B1(n17442), .B2(n17393), .A(n17380), .ZN(P3_U2739) );
  AOI22_X1 U20550 ( .A1(P3_DATAO_REG_27__SCAN_IN), .A2(n17409), .B1(n18832), 
        .B2(P3_UWORD_REG_11__SCAN_IN), .ZN(n17381) );
  OAI21_X1 U20551 ( .B1(n17440), .B2(n17393), .A(n17381), .ZN(P3_U2740) );
  INV_X1 U20552 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17438) );
  AOI22_X1 U20553 ( .A1(n17410), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17382) );
  OAI21_X1 U20554 ( .B1(n17438), .B2(n17393), .A(n17382), .ZN(P3_U2741) );
  AOI22_X1 U20555 ( .A1(n17410), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17383) );
  OAI21_X1 U20556 ( .B1(n17436), .B2(n17393), .A(n17383), .ZN(P3_U2742) );
  INV_X1 U20557 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17434) );
  AOI22_X1 U20558 ( .A1(P3_DATAO_REG_24__SCAN_IN), .A2(n17409), .B1(n18832), 
        .B2(P3_UWORD_REG_8__SCAN_IN), .ZN(n17384) );
  OAI21_X1 U20559 ( .B1(n17434), .B2(n17393), .A(n17384), .ZN(P3_U2743) );
  INV_X1 U20560 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17432) );
  AOI22_X1 U20561 ( .A1(P3_UWORD_REG_7__SCAN_IN), .A2(n18832), .B1(n17409), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17385) );
  OAI21_X1 U20562 ( .B1(n17432), .B2(n17393), .A(n17385), .ZN(P3_U2744) );
  INV_X1 U20563 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17430) );
  AOI22_X1 U20564 ( .A1(n17410), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17386) );
  OAI21_X1 U20565 ( .B1(n17430), .B2(n17393), .A(n17386), .ZN(P3_U2745) );
  AOI22_X1 U20566 ( .A1(P3_UWORD_REG_5__SCAN_IN), .A2(n17410), .B1(n17409), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17387) );
  OAI21_X1 U20567 ( .B1(n17428), .B2(n17393), .A(n17387), .ZN(P3_U2746) );
  AOI22_X1 U20568 ( .A1(n17410), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17388) );
  OAI21_X1 U20569 ( .B1(n17426), .B2(n17393), .A(n17388), .ZN(P3_U2747) );
  INV_X1 U20570 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17424) );
  AOI22_X1 U20571 ( .A1(n17410), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17389) );
  OAI21_X1 U20572 ( .B1(n17424), .B2(n17393), .A(n17389), .ZN(P3_U2748) );
  AOI22_X1 U20573 ( .A1(n17410), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17390) );
  OAI21_X1 U20574 ( .B1(n17422), .B2(n17393), .A(n17390), .ZN(P3_U2749) );
  INV_X1 U20575 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17420) );
  AOI22_X1 U20576 ( .A1(n17410), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17391) );
  OAI21_X1 U20577 ( .B1(n17420), .B2(n17393), .A(n17391), .ZN(P3_U2750) );
  INV_X1 U20578 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17418) );
  AOI22_X1 U20579 ( .A1(n17410), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17392) );
  OAI21_X1 U20580 ( .B1(n17418), .B2(n17393), .A(n17392), .ZN(P3_U2751) );
  AOI22_X1 U20581 ( .A1(n17410), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17395) );
  OAI21_X1 U20582 ( .B1(n17483), .B2(n17413), .A(n17395), .ZN(P3_U2752) );
  AOI22_X1 U20583 ( .A1(n17410), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17396) );
  OAI21_X1 U20584 ( .B1(n17478), .B2(n17413), .A(n17396), .ZN(P3_U2753) );
  INV_X1 U20585 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17475) );
  AOI22_X1 U20586 ( .A1(n17410), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17397) );
  OAI21_X1 U20587 ( .B1(n17475), .B2(n17413), .A(n17397), .ZN(P3_U2754) );
  INV_X1 U20588 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17473) );
  AOI22_X1 U20589 ( .A1(n17410), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17398) );
  OAI21_X1 U20590 ( .B1(n17473), .B2(n17413), .A(n17398), .ZN(P3_U2755) );
  AOI22_X1 U20591 ( .A1(n17410), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17399) );
  OAI21_X1 U20592 ( .B1(n17471), .B2(n17413), .A(n17399), .ZN(P3_U2756) );
  AOI22_X1 U20593 ( .A1(n17410), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17400) );
  OAI21_X1 U20594 ( .B1(n17468), .B2(n17413), .A(n17400), .ZN(P3_U2757) );
  AOI22_X1 U20595 ( .A1(n17410), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17401) );
  OAI21_X1 U20596 ( .B1(n17466), .B2(n17413), .A(n17401), .ZN(P3_U2758) );
  AOI22_X1 U20597 ( .A1(n17410), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17402) );
  OAI21_X1 U20598 ( .B1(n17464), .B2(n17413), .A(n17402), .ZN(P3_U2759) );
  INV_X1 U20599 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17462) );
  AOI22_X1 U20600 ( .A1(P3_LWORD_REG_7__SCAN_IN), .A2(n18832), .B1(n17409), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17403) );
  OAI21_X1 U20601 ( .B1(n17462), .B2(n17413), .A(n17403), .ZN(P3_U2760) );
  INV_X1 U20602 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17460) );
  AOI22_X1 U20603 ( .A1(P3_LWORD_REG_6__SCAN_IN), .A2(n18832), .B1(n17409), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17404) );
  OAI21_X1 U20604 ( .B1(n17460), .B2(n17413), .A(n17404), .ZN(P3_U2761) );
  INV_X1 U20605 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17458) );
  AOI22_X1 U20606 ( .A1(n17410), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17405) );
  OAI21_X1 U20607 ( .B1(n17458), .B2(n17413), .A(n17405), .ZN(P3_U2762) );
  INV_X1 U20608 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17456) );
  AOI22_X1 U20609 ( .A1(n17410), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17406) );
  OAI21_X1 U20610 ( .B1(n17456), .B2(n17413), .A(n17406), .ZN(P3_U2763) );
  AOI22_X1 U20611 ( .A1(n17410), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17407) );
  OAI21_X1 U20612 ( .B1(n17454), .B2(n17413), .A(n17407), .ZN(P3_U2764) );
  INV_X1 U20613 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17452) );
  AOI22_X1 U20614 ( .A1(n17410), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17408) );
  OAI21_X1 U20615 ( .B1(n17452), .B2(n17413), .A(n17408), .ZN(P3_U2765) );
  INV_X1 U20616 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17450) );
  AOI22_X1 U20617 ( .A1(n17410), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17411) );
  OAI21_X1 U20618 ( .B1(n17450), .B2(n17413), .A(n17411), .ZN(P3_U2766) );
  AOI22_X1 U20619 ( .A1(P3_DATAO_REG_0__SCAN_IN), .A2(n17409), .B1(n18832), 
        .B2(P3_LWORD_REG_0__SCAN_IN), .ZN(n17412) );
  OAI21_X1 U20620 ( .B1(n17448), .B2(n17413), .A(n17412), .ZN(P3_U2767) );
  NAND2_X1 U20621 ( .A1(n18835), .A2(n17416), .ZN(n18678) );
  AOI22_X1 U20622 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17480), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17479), .ZN(n17417) );
  OAI21_X1 U20623 ( .B1(n17418), .B2(n17482), .A(n17417), .ZN(P3_U2768) );
  AOI22_X1 U20624 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17480), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17479), .ZN(n17419) );
  OAI21_X1 U20625 ( .B1(n17420), .B2(n17482), .A(n17419), .ZN(P3_U2769) );
  AOI22_X1 U20626 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17480), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17479), .ZN(n17421) );
  OAI21_X1 U20627 ( .B1(n17422), .B2(n17482), .A(n17421), .ZN(P3_U2770) );
  AOI22_X1 U20628 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17480), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17479), .ZN(n17423) );
  OAI21_X1 U20629 ( .B1(n17424), .B2(n17482), .A(n17423), .ZN(P3_U2771) );
  AOI22_X1 U20630 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17476), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17479), .ZN(n17425) );
  OAI21_X1 U20631 ( .B1(n17426), .B2(n17482), .A(n17425), .ZN(P3_U2772) );
  AOI22_X1 U20632 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17476), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17479), .ZN(n17427) );
  OAI21_X1 U20633 ( .B1(n17428), .B2(n17482), .A(n17427), .ZN(P3_U2773) );
  AOI22_X1 U20634 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17476), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17479), .ZN(n17429) );
  OAI21_X1 U20635 ( .B1(n17430), .B2(n17482), .A(n17429), .ZN(P3_U2774) );
  AOI22_X1 U20636 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17476), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17479), .ZN(n17431) );
  OAI21_X1 U20637 ( .B1(n17432), .B2(n17482), .A(n17431), .ZN(P3_U2775) );
  AOI22_X1 U20638 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17476), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17479), .ZN(n17433) );
  OAI21_X1 U20639 ( .B1(n17434), .B2(n17482), .A(n17433), .ZN(P3_U2776) );
  AOI22_X1 U20640 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17476), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17479), .ZN(n17435) );
  OAI21_X1 U20641 ( .B1(n17436), .B2(n17482), .A(n17435), .ZN(P3_U2777) );
  AOI22_X1 U20642 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17476), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17479), .ZN(n17437) );
  OAI21_X1 U20643 ( .B1(n17438), .B2(n17482), .A(n17437), .ZN(P3_U2778) );
  AOI22_X1 U20644 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17476), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17479), .ZN(n17439) );
  OAI21_X1 U20645 ( .B1(n17440), .B2(n17482), .A(n17439), .ZN(P3_U2779) );
  AOI22_X1 U20646 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17480), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17479), .ZN(n17441) );
  OAI21_X1 U20647 ( .B1(n17442), .B2(n17482), .A(n17441), .ZN(P3_U2780) );
  AOI22_X1 U20648 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17480), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17479), .ZN(n17443) );
  OAI21_X1 U20649 ( .B1(n17444), .B2(n17482), .A(n17443), .ZN(P3_U2781) );
  AOI22_X1 U20650 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17480), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17479), .ZN(n17445) );
  OAI21_X1 U20651 ( .B1(n17446), .B2(n17482), .A(n17445), .ZN(P3_U2782) );
  AOI22_X1 U20652 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17480), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17479), .ZN(n17447) );
  OAI21_X1 U20653 ( .B1(n17448), .B2(n17482), .A(n17447), .ZN(P3_U2783) );
  AOI22_X1 U20654 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17480), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17479), .ZN(n17449) );
  OAI21_X1 U20655 ( .B1(n17450), .B2(n17482), .A(n17449), .ZN(P3_U2784) );
  AOI22_X1 U20656 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17480), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17469), .ZN(n17451) );
  OAI21_X1 U20657 ( .B1(n17452), .B2(n17482), .A(n17451), .ZN(P3_U2785) );
  AOI22_X1 U20658 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17480), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17469), .ZN(n17453) );
  OAI21_X1 U20659 ( .B1(n17454), .B2(n17482), .A(n17453), .ZN(P3_U2786) );
  AOI22_X1 U20660 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17480), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17469), .ZN(n17455) );
  OAI21_X1 U20661 ( .B1(n17456), .B2(n17482), .A(n17455), .ZN(P3_U2787) );
  AOI22_X1 U20662 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17480), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17469), .ZN(n17457) );
  OAI21_X1 U20663 ( .B1(n17458), .B2(n17482), .A(n17457), .ZN(P3_U2788) );
  AOI22_X1 U20664 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17480), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17469), .ZN(n17459) );
  OAI21_X1 U20665 ( .B1(n17460), .B2(n17482), .A(n17459), .ZN(P3_U2789) );
  AOI22_X1 U20666 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17480), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17469), .ZN(n17461) );
  OAI21_X1 U20667 ( .B1(n17462), .B2(n17482), .A(n17461), .ZN(P3_U2790) );
  AOI22_X1 U20668 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17480), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17469), .ZN(n17463) );
  OAI21_X1 U20669 ( .B1(n17464), .B2(n17482), .A(n17463), .ZN(P3_U2791) );
  AOI22_X1 U20670 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17476), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17469), .ZN(n17465) );
  OAI21_X1 U20671 ( .B1(n17466), .B2(n17482), .A(n17465), .ZN(P3_U2792) );
  AOI22_X1 U20672 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17480), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17469), .ZN(n17467) );
  OAI21_X1 U20673 ( .B1(n17468), .B2(n17482), .A(n17467), .ZN(P3_U2793) );
  AOI22_X1 U20674 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17480), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17469), .ZN(n17470) );
  OAI21_X1 U20675 ( .B1(n17471), .B2(n17482), .A(n17470), .ZN(P3_U2794) );
  AOI22_X1 U20676 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17476), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17479), .ZN(n17472) );
  OAI21_X1 U20677 ( .B1(n17473), .B2(n17482), .A(n17472), .ZN(P3_U2795) );
  AOI22_X1 U20678 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17480), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17479), .ZN(n17474) );
  OAI21_X1 U20679 ( .B1(n17475), .B2(n17482), .A(n17474), .ZN(P3_U2796) );
  AOI22_X1 U20680 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17476), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17479), .ZN(n17477) );
  OAI21_X1 U20681 ( .B1(n17478), .B2(n17482), .A(n17477), .ZN(P3_U2797) );
  AOI22_X1 U20682 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17480), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17479), .ZN(n17481) );
  OAI21_X1 U20683 ( .B1(n17483), .B2(n17482), .A(n17481), .ZN(P3_U2798) );
  INV_X1 U20684 ( .A(n17810), .ZN(n17756) );
  OAI22_X1 U20685 ( .A1(n17485), .A2(n17756), .B1(n17484), .B2(n17856), .ZN(
        n17486) );
  NOR2_X1 U20686 ( .A1(n17843), .A2(n17486), .ZN(n17522) );
  OAI21_X1 U20687 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17640), .A(
        n17522), .ZN(n17509) );
  AOI22_X1 U20688 ( .A1(n17692), .A2(n17487), .B1(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n17509), .ZN(n17503) );
  NOR2_X1 U20689 ( .A1(n17766), .A2(n17848), .ZN(n17612) );
  AOI22_X1 U20690 ( .A1(n17488), .A2(n17766), .B1(n17868), .B2(n17848), .ZN(
        n17489) );
  INV_X1 U20691 ( .A(n17489), .ZN(n17524) );
  NOR2_X1 U20692 ( .A1(n17871), .A2(n17524), .ZN(n17491) );
  NOR3_X1 U20693 ( .A1(n17612), .A2(n17491), .A3(n17490), .ZN(n17496) );
  AOI211_X1 U20694 ( .C1(n17494), .C2(n17493), .A(n17492), .B(n17764), .ZN(
        n17495) );
  AOI211_X1 U20695 ( .C1(n17497), .C2(n17512), .A(n17496), .B(n17495), .ZN(
        n17502) );
  NAND2_X1 U20696 ( .A1(n9736), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17501) );
  NOR2_X1 U20697 ( .A1(n17702), .A2(n17498), .ZN(n17511) );
  NAND2_X1 U20698 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17499) );
  OAI211_X1 U20699 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17511), .B(n17499), .ZN(n17500) );
  NAND4_X1 U20700 ( .A1(n17503), .A2(n17502), .A3(n17501), .A4(n17500), .ZN(
        P3_U2802) );
  NAND2_X1 U20701 ( .A1(n17505), .A2(n9933), .ZN(n17506) );
  XOR2_X1 U20702 ( .A(n17506), .B(n17598), .Z(n17876) );
  INV_X1 U20703 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17510) );
  OAI22_X1 U20704 ( .A1(n18169), .A2(n18765), .B1(n17709), .B2(n17507), .ZN(
        n17508) );
  AOI221_X1 U20705 ( .B1(n17511), .B2(n17510), .C1(n17509), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17508), .ZN(n17514) );
  AOI22_X1 U20706 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17524), .B1(
        n17512), .B2(n17871), .ZN(n17513) );
  OAI211_X1 U20707 ( .C1(n17876), .C2(n17764), .A(n17514), .B(n17513), .ZN(
        P3_U2803) );
  AOI21_X1 U20708 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17516), .A(
        n17515), .ZN(n17883) );
  NOR2_X1 U20709 ( .A1(n17517), .A2(n17590), .ZN(n17526) );
  AOI21_X1 U20710 ( .B1(n17518), .B2(n18566), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17521) );
  OAI21_X1 U20711 ( .B1(n17692), .B2(n17563), .A(n17519), .ZN(n17520) );
  NAND2_X1 U20712 ( .A1(n9736), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17881) );
  OAI211_X1 U20713 ( .C1(n17522), .C2(n17521), .A(n17520), .B(n17881), .ZN(
        n17523) );
  AOI221_X1 U20714 ( .B1(n17526), .B2(n17525), .C1(n17524), .C2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n17523), .ZN(n17527) );
  OAI21_X1 U20715 ( .B1(n17883), .B2(n17764), .A(n17527), .ZN(P3_U2804) );
  OAI21_X1 U20716 ( .B1(n17598), .B2(n17529), .A(n17528), .ZN(n17530) );
  XOR2_X1 U20717 ( .A(n17530), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17890) );
  NAND2_X1 U20718 ( .A1(n18566), .A2(n17532), .ZN(n17564) );
  OAI211_X1 U20719 ( .C1(n17531), .C2(n17856), .A(n17857), .B(n17564), .ZN(
        n17561) );
  AOI21_X1 U20720 ( .B1(n17563), .B2(n21169), .A(n17561), .ZN(n17546) );
  NOR2_X1 U20721 ( .A1(n17702), .A2(n17532), .ZN(n17545) );
  OAI211_X1 U20722 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17545), .B(n17533), .ZN(n17534) );
  NAND2_X1 U20723 ( .A1(n9736), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17894) );
  OAI211_X1 U20724 ( .C1(n17546), .C2(n17535), .A(n17534), .B(n17894), .ZN(
        n17536) );
  AOI21_X1 U20725 ( .B1(n17692), .B2(n17537), .A(n17536), .ZN(n17542) );
  AOI21_X1 U20726 ( .B1(n17896), .B2(n17539), .A(n17538), .ZN(n17889) );
  NOR2_X1 U20727 ( .A1(n17552), .A2(n18000), .ZN(n17897) );
  INV_X1 U20728 ( .A(n17897), .ZN(n17551) );
  AOI221_X1 U20729 ( .B1(n17904), .B2(n17896), .C1(n17551), .C2(n17896), .A(
        n17540), .ZN(n17893) );
  AOI22_X1 U20730 ( .A1(n17766), .A2(n17889), .B1(n17848), .B2(n17893), .ZN(
        n17541) );
  OAI211_X1 U20731 ( .C1(n17764), .C2(n17890), .A(n17542), .B(n17541), .ZN(
        P3_U2805) );
  AOI21_X1 U20732 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17544), .A(
        n17543), .ZN(n17910) );
  INV_X1 U20733 ( .A(n17545), .ZN(n17548) );
  NAND2_X1 U20734 ( .A1(n9736), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n17908) );
  OAI221_X1 U20735 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n17548), .C1(
        n17547), .C2(n17546), .A(n17908), .ZN(n17549) );
  AOI21_X1 U20736 ( .B1(n17692), .B2(n17550), .A(n17549), .ZN(n17554) );
  NAND2_X1 U20737 ( .A1(n17551), .A2(n17848), .ZN(n17555) );
  OAI21_X1 U20738 ( .B1(n17898), .B2(n17579), .A(n17555), .ZN(n17571) );
  NOR2_X1 U20739 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17552), .ZN(
        n17907) );
  AOI22_X1 U20740 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17571), .B1(
        n17661), .B2(n17907), .ZN(n17553) );
  OAI211_X1 U20741 ( .C1(n17910), .C2(n17764), .A(n17554), .B(n17553), .ZN(
        P3_U2806) );
  NOR2_X1 U20742 ( .A1(n17898), .A2(n17579), .ZN(n17557) );
  INV_X1 U20743 ( .A(n17555), .ZN(n17556) );
  AOI22_X1 U20744 ( .A1(n17578), .A2(n17557), .B1(n17577), .B2(n17556), .ZN(
        n17573) );
  AOI22_X1 U20745 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17598), .B1(
        n17558), .B2(n17575), .ZN(n17559) );
  NAND2_X1 U20746 ( .A1(n17605), .A2(n17559), .ZN(n17560) );
  XOR2_X1 U20747 ( .A(n17560), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(
        n17917) );
  AOI22_X1 U20748 ( .A1(n17692), .A2(n17562), .B1(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17561), .ZN(n17569) );
  NAND2_X1 U20749 ( .A1(n17563), .A2(n21169), .ZN(n17565) );
  OAI21_X1 U20750 ( .B1(n17565), .B2(n17849), .A(n17564), .ZN(n17566) );
  AOI22_X1 U20751 ( .A1(n9736), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n17567), 
        .B2(n17566), .ZN(n17568) );
  OAI211_X1 U20752 ( .C1(n17764), .C2(n17917), .A(n17569), .B(n17568), .ZN(
        n17570) );
  AOI21_X1 U20753 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17571), .A(
        n17570), .ZN(n17572) );
  OAI21_X1 U20754 ( .B1(n17573), .B2(n17911), .A(n17572), .ZN(P3_U2807) );
  NOR2_X1 U20755 ( .A1(n17941), .A2(n17921), .ZN(n17924) );
  INV_X1 U20756 ( .A(n17924), .ZN(n17862) );
  INV_X1 U20757 ( .A(n17605), .ZN(n17574) );
  AOI221_X1 U20758 ( .B1(n17651), .B2(n17575), .C1(n17862), .C2(n17575), .A(
        n17574), .ZN(n17576) );
  XOR2_X1 U20759 ( .A(n17920), .B(n17576), .Z(n17935) );
  OAI22_X1 U20760 ( .A1(n17579), .A2(n17578), .B1(n17861), .B2(n17577), .ZN(
        n17660) );
  INV_X1 U20761 ( .A(n17660), .ZN(n17611) );
  OAI21_X1 U20762 ( .B1(n17612), .B2(n17924), .A(n17611), .ZN(n17602) );
  OAI21_X1 U20763 ( .B1(n17580), .B2(n17856), .A(n17857), .ZN(n17581) );
  AOI21_X1 U20764 ( .B1(n17810), .B2(n17583), .A(n17581), .ZN(n17608) );
  OAI21_X1 U20765 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17640), .A(
        n17608), .ZN(n17594) );
  AOI22_X1 U20766 ( .A1(n17692), .A2(n17582), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17594), .ZN(n17587) );
  NAND2_X1 U20767 ( .A1(n9736), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17933) );
  NAND3_X1 U20768 ( .A1(n17661), .A2(n17924), .A3(n17920), .ZN(n17586) );
  NOR2_X1 U20769 ( .A1(n17702), .A2(n17583), .ZN(n17596) );
  OAI211_X1 U20770 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17596), .B(n17584), .ZN(n17585) );
  NAND4_X1 U20771 ( .A1(n17587), .A2(n17933), .A3(n17586), .A4(n17585), .ZN(
        n17588) );
  AOI21_X1 U20772 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17602), .A(
        n17588), .ZN(n17589) );
  OAI21_X1 U20773 ( .B1(n17764), .B2(n17935), .A(n17589), .ZN(P3_U2808) );
  NAND2_X1 U20774 ( .A1(n17938), .A2(n17927), .ZN(n17946) );
  NOR2_X1 U20775 ( .A1(n17941), .A2(n17590), .ZN(n17613) );
  INV_X1 U20776 ( .A(n17613), .ZN(n17627) );
  AOI22_X1 U20777 ( .A1(n9736), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n17692), 
        .B2(n17591), .ZN(n17592) );
  INV_X1 U20778 ( .A(n17592), .ZN(n17593) );
  AOI221_X1 U20779 ( .B1(n17596), .B2(n17595), .C1(n17594), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17593), .ZN(n17604) );
  INV_X1 U20780 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21138) );
  NOR3_X1 U20781 ( .A1(n17598), .A2(n21138), .A3(n17597), .ZN(n17622) );
  INV_X1 U20782 ( .A(n17599), .ZN(n17635) );
  AOI22_X1 U20783 ( .A1(n17938), .A2(n17622), .B1(n17635), .B2(n17600), .ZN(
        n17601) );
  XOR2_X1 U20784 ( .A(n17927), .B(n17601), .Z(n17936) );
  AOI22_X1 U20785 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17602), .B1(
        n17752), .B2(n17936), .ZN(n17603) );
  OAI211_X1 U20786 ( .C1(n17946), .C2(n17627), .A(n17604), .B(n17603), .ZN(
        P3_U2809) );
  OAI221_X1 U20787 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17634), 
        .C1(n17964), .C2(n17622), .A(n17605), .ZN(n17606) );
  XOR2_X1 U20788 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17606), .Z(
        n17958) );
  AOI21_X1 U20789 ( .B1(n9802), .B2(n18566), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17607) );
  NAND2_X1 U20790 ( .A1(n9736), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17956) );
  OAI21_X1 U20791 ( .B1(n17608), .B2(n17607), .A(n17956), .ZN(n17609) );
  AOI221_X1 U20792 ( .B1(n17692), .B2(n17610), .C1(n17563), .C2(n17610), .A(
        n17609), .ZN(n17615) );
  NOR2_X1 U20793 ( .A1(n17941), .A2(n17964), .ZN(n17949) );
  OAI21_X1 U20794 ( .B1(n17612), .B2(n17949), .A(n17611), .ZN(n17624) );
  NOR2_X1 U20795 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17964), .ZN(
        n17954) );
  AOI22_X1 U20796 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17624), .B1(
        n17613), .B2(n17954), .ZN(n17614) );
  OAI211_X1 U20797 ( .C1(n17764), .C2(n17958), .A(n17615), .B(n17614), .ZN(
        P3_U2810) );
  AOI21_X1 U20798 ( .B1(n17810), .B2(n17617), .A(n17843), .ZN(n17642) );
  OAI21_X1 U20799 ( .B1(n17616), .B2(n17856), .A(n17642), .ZN(n17631) );
  NOR2_X1 U20800 ( .A1(n17702), .A2(n17617), .ZN(n17633) );
  OAI211_X1 U20801 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17633), .B(n17618), .ZN(n17619) );
  NAND2_X1 U20802 ( .A1(n9736), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17961) );
  OAI211_X1 U20803 ( .C1(n17709), .C2(n17620), .A(n17619), .B(n17961), .ZN(
        n17621) );
  AOI21_X1 U20804 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17631), .A(
        n17621), .ZN(n17626) );
  AOI21_X1 U20805 ( .B1(n17634), .B2(n17635), .A(n17622), .ZN(n17623) );
  XOR2_X1 U20806 ( .A(n17964), .B(n17623), .Z(n17960) );
  AOI22_X1 U20807 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17624), .B1(
        n17752), .B2(n17960), .ZN(n17625) );
  OAI211_X1 U20808 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17627), .A(
        n17626), .B(n17625), .ZN(P3_U2811) );
  INV_X1 U20809 ( .A(n17628), .ZN(n17967) );
  AOI21_X1 U20810 ( .B1(n17661), .B2(n17967), .A(n17660), .ZN(n17649) );
  INV_X1 U20811 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17632) );
  OAI22_X1 U20812 ( .A1(n18169), .A2(n18746), .B1(n17709), .B2(n17629), .ZN(
        n17630) );
  AOI221_X1 U20813 ( .B1(n17633), .B2(n17632), .C1(n17631), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17630), .ZN(n17638) );
  AOI21_X1 U20814 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17761), .A(
        n17634), .ZN(n17636) );
  XOR2_X1 U20815 ( .A(n17636), .B(n17635), .Z(n17978) );
  NOR2_X1 U20816 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17967), .ZN(
        n17977) );
  AOI22_X1 U20817 ( .A1(n17752), .A2(n17978), .B1(n17661), .B2(n17977), .ZN(
        n17637) );
  OAI211_X1 U20818 ( .C1(n17649), .C2(n21138), .A(n17638), .B(n17637), .ZN(
        P3_U2812) );
  AOI21_X1 U20819 ( .B1(n17639), .B2(n18566), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17643) );
  OAI22_X1 U20820 ( .A1(n17643), .A2(n17642), .B1(n17840), .B2(n17641), .ZN(
        n17644) );
  AOI21_X1 U20821 ( .B1(n9736), .B2(P3_REIP_REG_17__SCAN_IN), .A(n17644), .ZN(
        n17648) );
  OAI21_X1 U20822 ( .B1(n17646), .B2(n17970), .A(n17645), .ZN(n17983) );
  NOR2_X1 U20823 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17992), .ZN(
        n17982) );
  AOI22_X1 U20824 ( .A1(n17752), .A2(n17983), .B1(n17661), .B2(n17982), .ZN(
        n17647) );
  OAI211_X1 U20825 ( .C1(n17649), .C2(n17970), .A(n17648), .B(n17647), .ZN(
        P3_U2813) );
  AOI21_X1 U20826 ( .B1(n17761), .B2(n17651), .A(n17650), .ZN(n17652) );
  XOR2_X1 U20827 ( .A(n17992), .B(n17652), .Z(n17997) );
  INV_X1 U20828 ( .A(n17856), .ZN(n17688) );
  OAI21_X1 U20829 ( .B1(n17655), .B2(n17756), .A(n17857), .ZN(n17677) );
  AOI21_X1 U20830 ( .B1(n17688), .B2(n17653), .A(n17677), .ZN(n17663) );
  AOI21_X1 U20831 ( .B1(n17664), .B2(n17659), .A(n9761), .ZN(n17657) );
  NAND2_X1 U20832 ( .A1(n9736), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n17995) );
  AOI21_X1 U20833 ( .B1(n17662), .B2(n18029), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18007) );
  NAND2_X1 U20834 ( .A1(n17766), .A2(n17998), .ZN(n17674) );
  NAND2_X1 U20835 ( .A1(n9736), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18010) );
  OAI221_X1 U20836 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n9761), .C1(
        n17664), .C2(n17663), .A(n18010), .ZN(n17671) );
  INV_X1 U20837 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18019) );
  INV_X1 U20838 ( .A(n18015), .ZN(n17683) );
  NOR3_X1 U20839 ( .A1(n17974), .A2(n18019), .A3(n17683), .ZN(n17684) );
  NOR2_X1 U20840 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17684), .ZN(
        n18005) );
  NAND2_X1 U20841 ( .A1(n17848), .A2(n18000), .ZN(n17669) );
  NAND2_X1 U20842 ( .A1(n17699), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17698) );
  INV_X1 U20843 ( .A(n17698), .ZN(n18036) );
  NAND2_X1 U20844 ( .A1(n17761), .A2(n17759), .ZN(n17744) );
  NOR3_X1 U20845 ( .A1(n18035), .A2(n18048), .A3(n17744), .ZN(n17675) );
  NOR2_X1 U20846 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17666) );
  NOR2_X1 U20847 ( .A1(n17761), .A2(n17665), .ZN(n17714) );
  AOI22_X1 U20848 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17675), .B1(
        n17666), .B2(n17714), .ZN(n17667) );
  NOR2_X1 U20849 ( .A1(n18036), .A2(n17667), .ZN(n17668) );
  XNOR2_X1 U20850 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17668), .ZN(
        n18012) );
  OAI22_X1 U20851 ( .A1(n18005), .A2(n17669), .B1(n17764), .B2(n18012), .ZN(
        n17670) );
  AOI211_X1 U20852 ( .C1(n17692), .C2(n17672), .A(n17671), .B(n17670), .ZN(
        n17673) );
  OAI21_X1 U20853 ( .B1(n18007), .B2(n17674), .A(n17673), .ZN(P3_U2815) );
  OAI221_X1 U20854 ( .B1(n17675), .B2(n17714), .C1(n17675), .C2(n17699), .A(
        n17698), .ZN(n17676) );
  XOR2_X1 U20855 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17676), .Z(
        n18025) );
  OAI221_X1 U20856 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n17678), .C1(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n18566), .A(n17677), .ZN(
        n17679) );
  OAI21_X1 U20857 ( .B1(n17840), .B2(n17680), .A(n17679), .ZN(n17681) );
  AOI21_X1 U20858 ( .B1(n9736), .B2(P3_REIP_REG_14__SCAN_IN), .A(n17681), .ZN(
        n17687) );
  NOR2_X1 U20859 ( .A1(n17973), .A2(n17990), .ZN(n17682) );
  AOI221_X1 U20860 ( .B1(n17683), .B2(n18019), .C1(n17973), .C2(n18019), .A(
        n17682), .ZN(n18022) );
  NAND2_X1 U20861 ( .A1(n18015), .A2(n18027), .ZN(n17685) );
  AOI21_X1 U20862 ( .B1(n18019), .B2(n17685), .A(n17684), .ZN(n18021) );
  AOI22_X1 U20863 ( .A1(n17766), .A2(n18022), .B1(n17848), .B2(n18021), .ZN(
        n17686) );
  OAI211_X1 U20864 ( .C1(n17764), .C2(n18025), .A(n17687), .B(n17686), .ZN(
        P3_U2816) );
  AOI21_X1 U20865 ( .B1(n17810), .B2(n17701), .A(n17688), .ZN(n17689) );
  OAI21_X1 U20866 ( .B1(n17690), .B2(n17689), .A(n17857), .ZN(n17711) );
  AOI22_X1 U20867 ( .A1(n17692), .A2(n17691), .B1(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17711), .ZN(n17707) );
  OAI22_X1 U20868 ( .A1(n17761), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n17693), .B2(n18014), .ZN(n17695) );
  NAND2_X1 U20869 ( .A1(n17695), .A2(n17694), .ZN(n17696) );
  XOR2_X1 U20870 ( .A(n17696), .B(n17699), .Z(n18037) );
  INV_X1 U20871 ( .A(n17755), .ZN(n17697) );
  AOI22_X1 U20872 ( .A1(n17973), .A2(n17766), .B1(n17848), .B2(n17974), .ZN(
        n17754) );
  INV_X1 U20873 ( .A(n17754), .ZN(n17740) );
  AOI21_X1 U20874 ( .B1(n18014), .B2(n17697), .A(n17740), .ZN(n17717) );
  OR2_X1 U20875 ( .A1(n18035), .A2(n17755), .ZN(n17718) );
  OAI22_X1 U20876 ( .A1(n17717), .A2(n17699), .B1(n17698), .B2(n17718), .ZN(
        n17700) );
  AOI21_X1 U20877 ( .B1(n17752), .B2(n18037), .A(n17700), .ZN(n17706) );
  NAND2_X1 U20878 ( .A1(n9736), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17705) );
  NOR2_X1 U20879 ( .A1(n17702), .A2(n17701), .ZN(n17713) );
  OAI211_X1 U20880 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17713), .B(n17703), .ZN(n17704) );
  NAND4_X1 U20881 ( .A1(n17707), .A2(n17706), .A3(n17705), .A4(n17704), .ZN(
        P3_U2817) );
  INV_X1 U20882 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17712) );
  NAND2_X1 U20883 ( .A1(n9736), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18046) );
  OAI21_X1 U20884 ( .B1(n17709), .B2(n17708), .A(n18046), .ZN(n17710) );
  AOI221_X1 U20885 ( .B1(n17713), .B2(n17712), .C1(n17711), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17710), .ZN(n17721) );
  INV_X1 U20886 ( .A(n17714), .ZN(n17715) );
  OAI21_X1 U20887 ( .B1(n17744), .B2(n18035), .A(n17715), .ZN(n17716) );
  XOR2_X1 U20888 ( .A(n17716), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n18045) );
  AOI21_X1 U20889 ( .B1(n18048), .B2(n17718), .A(n17717), .ZN(n17719) );
  AOI21_X1 U20890 ( .B1(n18045), .B2(n17752), .A(n17719), .ZN(n17720) );
  NAND2_X1 U20891 ( .A1(n17721), .A2(n17720), .ZN(P3_U2818) );
  NAND2_X1 U20892 ( .A1(n17730), .A2(n18026), .ZN(n18061) );
  NAND2_X1 U20893 ( .A1(n17722), .A2(n21143), .ZN(n17745) );
  OAI22_X1 U20894 ( .A1(n18055), .A2(n17744), .B1(n17739), .B2(n17745), .ZN(
        n17723) );
  XOR2_X1 U20895 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17723), .Z(
        n18049) );
  NOR3_X1 U20896 ( .A1(n17787), .A2(n17788), .A3(n18219), .ZN(n17776) );
  INV_X1 U20897 ( .A(n17790), .ZN(n17851) );
  INV_X1 U20898 ( .A(n17776), .ZN(n17724) );
  NOR2_X1 U20899 ( .A1(n17767), .A2(n17724), .ZN(n17748) );
  NAND2_X1 U20900 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17748), .ZN(
        n17747) );
  NOR2_X1 U20901 ( .A1(n17735), .A2(n17747), .ZN(n17734) );
  AOI21_X1 U20902 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17851), .A(
        n17734), .ZN(n17725) );
  AOI21_X1 U20903 ( .B1(n17776), .B2(n17726), .A(n17725), .ZN(n17729) );
  INV_X1 U20904 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18734) );
  OAI22_X1 U20905 ( .A1(n17840), .A2(n17727), .B1(n18169), .B2(n18734), .ZN(
        n17728) );
  AOI211_X1 U20906 ( .C1(n17752), .C2(n18049), .A(n17729), .B(n17728), .ZN(
        n17732) );
  NOR2_X1 U20907 ( .A1(n17730), .A2(n17755), .ZN(n17741) );
  OAI21_X1 U20908 ( .B1(n17741), .B2(n17740), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17731) );
  OAI211_X1 U20909 ( .C1(n17755), .C2(n18061), .A(n17732), .B(n17731), .ZN(
        P3_U2819) );
  AOI22_X1 U20910 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17744), .B1(
        n17745), .B2(n18069), .ZN(n17733) );
  XOR2_X1 U20911 ( .A(n18062), .B(n17733), .Z(n18068) );
  AOI211_X1 U20912 ( .C1(n17747), .C2(n17735), .A(n17790), .B(n17734), .ZN(
        n17737) );
  NOR2_X1 U20913 ( .A1(n18169), .A2(n18732), .ZN(n17736) );
  AOI211_X1 U20914 ( .C1(n17738), .C2(n17850), .A(n17737), .B(n17736), .ZN(
        n17743) );
  OAI221_X1 U20915 ( .B1(n17741), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), 
        .C1(n17741), .C2(n17740), .A(n17739), .ZN(n17742) );
  OAI211_X1 U20916 ( .C1(n18068), .C2(n17764), .A(n17743), .B(n17742), .ZN(
        P3_U2820) );
  NAND2_X1 U20917 ( .A1(n17745), .A2(n17744), .ZN(n17746) );
  XOR2_X1 U20918 ( .A(n17746), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n18072) );
  OAI211_X1 U20919 ( .C1(n17748), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n17851), .B(n17747), .ZN(n17749) );
  NAND2_X1 U20920 ( .A1(n9736), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n18074) );
  OAI211_X1 U20921 ( .C1(n17840), .C2(n17750), .A(n17749), .B(n18074), .ZN(
        n17751) );
  AOI21_X1 U20922 ( .B1(n17752), .B2(n18072), .A(n17751), .ZN(n17753) );
  OAI221_X1 U20923 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17755), .C1(
        n18069), .C2(n17754), .A(n17753), .ZN(P3_U2821) );
  OAI21_X1 U20924 ( .B1(n17757), .B2(n17756), .A(n17857), .ZN(n17774) );
  AOI22_X1 U20925 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17774), .B1(
        n17758), .B2(n17850), .ZN(n17771) );
  NOR2_X1 U20926 ( .A1(n17760), .A2(n17759), .ZN(n18081) );
  XOR2_X1 U20927 ( .A(n18081), .B(n17761), .Z(n18079) );
  OAI21_X1 U20928 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17763), .A(
        n17762), .ZN(n18077) );
  OAI22_X1 U20929 ( .A1(n18079), .A2(n17764), .B1(n17861), .B2(n18077), .ZN(
        n17765) );
  AOI21_X1 U20930 ( .B1(n17766), .B2(n18081), .A(n17765), .ZN(n17770) );
  NAND2_X1 U20931 ( .A1(n9736), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18091) );
  OAI211_X1 U20932 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17768), .A(
        n18566), .B(n17767), .ZN(n17769) );
  NAND4_X1 U20933 ( .A1(n17771), .A2(n17770), .A3(n18091), .A4(n17769), .ZN(
        P3_U2822) );
  OAI21_X1 U20934 ( .B1(n17773), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n17772), .ZN(n18101) );
  NOR2_X1 U20935 ( .A1(n18169), .A2(n18726), .ZN(n18093) );
  AOI221_X1 U20936 ( .B1(n17776), .B2(n17775), .C1(n17774), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18093), .ZN(n17783) );
  AOI21_X1 U20937 ( .B1(n17779), .B2(n17778), .A(n17777), .ZN(n17780) );
  XOR2_X1 U20938 ( .A(n17780), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18098) );
  AOI22_X1 U20939 ( .A1(n17848), .A2(n18098), .B1(n17781), .B2(n17850), .ZN(
        n17782) );
  OAI211_X1 U20940 ( .C1(n17860), .C2(n18101), .A(n17783), .B(n17782), .ZN(
        P3_U2823) );
  OAI21_X1 U20941 ( .B1(n17786), .B2(n17785), .A(n17784), .ZN(n18103) );
  NOR2_X1 U20942 ( .A1(n17787), .A2(n18219), .ZN(n17789) );
  AOI22_X1 U20943 ( .A1(n9736), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n17789), .B2(
        n17788), .ZN(n17796) );
  NOR2_X1 U20944 ( .A1(n17790), .A2(n17789), .ZN(n17805) );
  OAI21_X1 U20945 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17792), .A(
        n17791), .ZN(n18109) );
  OAI22_X1 U20946 ( .A1(n17840), .A2(n17793), .B1(n17861), .B2(n18109), .ZN(
        n17794) );
  AOI21_X1 U20947 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17805), .A(
        n17794), .ZN(n17795) );
  OAI211_X1 U20948 ( .C1(n17860), .C2(n18103), .A(n17796), .B(n17795), .ZN(
        P3_U2824) );
  OAI21_X1 U20949 ( .B1(n17799), .B2(n17798), .A(n17797), .ZN(n17800) );
  XOR2_X1 U20950 ( .A(n17800), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(
        n18110) );
  OAI21_X1 U20951 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17802), .A(
        n17801), .ZN(n18116) );
  OAI22_X1 U20952 ( .A1(n17860), .A2(n18116), .B1(n18169), .B2(n18722), .ZN(
        n17803) );
  AOI21_X1 U20953 ( .B1(n17804), .B2(n17850), .A(n17803), .ZN(n17808) );
  OAI221_X1 U20954 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17806), .C1(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n17857), .A(n17805), .ZN(n17807) );
  OAI211_X1 U20955 ( .C1(n18110), .C2(n17861), .A(n17808), .B(n17807), .ZN(
        P3_U2825) );
  AOI21_X1 U20956 ( .B1(n17810), .B2(n17809), .A(n17843), .ZN(n17829) );
  OAI21_X1 U20957 ( .B1(n17813), .B2(n17812), .A(n17811), .ZN(n18118) );
  OAI22_X1 U20958 ( .A1(n17861), .A2(n18118), .B1(n18169), .B2(n20983), .ZN(
        n17818) );
  OAI22_X1 U20959 ( .A1(n17840), .A2(n17816), .B1(n17860), .B2(n18119), .ZN(
        n17817) );
  AOI211_X1 U20960 ( .C1(n18566), .C2(n17819), .A(n17818), .B(n17817), .ZN(
        n17820) );
  OAI21_X1 U20961 ( .B1(n17829), .B2(n17821), .A(n17820), .ZN(P3_U2826) );
  XOR2_X1 U20962 ( .A(n17824), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(
        n18128) );
  AOI21_X1 U20963 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17857), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17828) );
  OAI21_X1 U20964 ( .B1(n17827), .B2(n17826), .A(n17825), .ZN(n18129) );
  OAI22_X1 U20965 ( .A1(n17829), .A2(n17828), .B1(n17861), .B2(n18129), .ZN(
        n17830) );
  AOI21_X1 U20966 ( .B1(n17831), .B2(n17850), .A(n17830), .ZN(n17832) );
  NAND2_X1 U20967 ( .A1(n9736), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18134) );
  OAI211_X1 U20968 ( .C1(n17860), .C2(n18128), .A(n17832), .B(n18134), .ZN(
        P3_U2827) );
  OAI21_X1 U20969 ( .B1(n17835), .B2(n17834), .A(n17833), .ZN(n18147) );
  OAI21_X1 U20970 ( .B1(n17838), .B2(n17837), .A(n17836), .ZN(n18152) );
  OAI22_X1 U20971 ( .A1(n17840), .A2(n17839), .B1(n17860), .B2(n18152), .ZN(
        n17841) );
  AOI221_X1 U20972 ( .B1(n17843), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18566), .C2(n17842), .A(n17841), .ZN(n17844) );
  NAND2_X1 U20973 ( .A1(n9736), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18150) );
  OAI211_X1 U20974 ( .C1(n17861), .C2(n18147), .A(n17844), .B(n18150), .ZN(
        P3_U2828) );
  OAI21_X1 U20975 ( .B1(n17854), .B2(n17846), .A(n17845), .ZN(n18163) );
  NAND2_X1 U20976 ( .A1(n18796), .A2(n17855), .ZN(n17847) );
  XNOR2_X1 U20977 ( .A(n17847), .B(n17846), .ZN(n18159) );
  AOI22_X1 U20978 ( .A1(n17848), .A2(n18159), .B1(n9736), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17853) );
  AOI22_X1 U20979 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17851), .B1(
        n17850), .B2(n17849), .ZN(n17852) );
  OAI211_X1 U20980 ( .C1(n17860), .C2(n18163), .A(n17853), .B(n17852), .ZN(
        P3_U2829) );
  AOI21_X1 U20981 ( .B1(n17855), .B2(n18796), .A(n17854), .ZN(n18167) );
  INV_X1 U20982 ( .A(n18167), .ZN(n18165) );
  NAND3_X1 U20983 ( .A1(n20974), .A2(n17857), .A3(n17856), .ZN(n17858) );
  AOI22_X1 U20984 ( .A1(n9736), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17858), .ZN(n17859) );
  OAI221_X1 U20985 ( .B1(n18167), .B2(n17861), .C1(n18165), .C2(n17860), .A(
        n17859), .ZN(P3_U2830) );
  AOI22_X1 U20986 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18149), .B1(
        n9736), .B2(P3_REIP_REG_27__SCAN_IN), .ZN(n17875) );
  NOR2_X1 U20987 ( .A1(n18170), .A2(n17871), .ZN(n17872) );
  NAND2_X1 U20988 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17865) );
  NOR2_X1 U20989 ( .A1(n17965), .A2(n17862), .ZN(n17863) );
  NOR2_X1 U20990 ( .A1(n18796), .A2(n17965), .ZN(n17986) );
  INV_X1 U20991 ( .A(n17986), .ZN(n17940) );
  OAI22_X1 U20992 ( .A1(n18641), .A2(n17920), .B1(n17911), .B2(n17940), .ZN(
        n17929) );
  AOI21_X1 U20993 ( .B1(n17863), .B2(n17929), .A(n18139), .ZN(n17900) );
  AOI211_X1 U20994 ( .C1(n17865), .C2(n18084), .A(n17900), .B(n17864), .ZN(
        n17887) );
  AOI22_X1 U20995 ( .A1(n18001), .A2(n17868), .B1(n17867), .B2(n17866), .ZN(
        n17869) );
  OAI211_X1 U20996 ( .C1(n17870), .C2(n18028), .A(n17887), .B(n17869), .ZN(
        n17880) );
  OAI22_X1 U20997 ( .A1(n17873), .A2(n17872), .B1(n17880), .B2(n17871), .ZN(
        n17874) );
  OAI211_X1 U20998 ( .C1(n17876), .C2(n18078), .A(n17875), .B(n17874), .ZN(
        P3_U2835) );
  NAND2_X1 U20999 ( .A1(n17878), .A2(n17877), .ZN(n17879) );
  AOI22_X1 U21000 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18149), .B1(
        n17880), .B2(n17879), .ZN(n17882) );
  OAI211_X1 U21001 ( .C1(n17883), .C2(n18078), .A(n17882), .B(n17881), .ZN(
        P3_U2836) );
  NAND3_X1 U21002 ( .A1(n17885), .A2(n17884), .A3(n17896), .ZN(n17886) );
  OAI21_X1 U21003 ( .B1(n17887), .B2(n17896), .A(n17886), .ZN(n17888) );
  AOI21_X1 U21004 ( .B1(n17999), .B2(n17889), .A(n17888), .ZN(n17891) );
  OAI22_X1 U21005 ( .A1(n17891), .A2(n18170), .B1(n18078), .B2(n17890), .ZN(
        n17892) );
  AOI21_X1 U21006 ( .B1(n18166), .B2(n17893), .A(n17892), .ZN(n17895) );
  OAI211_X1 U21007 ( .C1(n18155), .C2(n17896), .A(n17895), .B(n17894), .ZN(
        P3_U2837) );
  OAI22_X1 U21008 ( .A1(n17898), .A2(n18028), .B1(n17897), .B2(n18658), .ZN(
        n17899) );
  NOR3_X1 U21009 ( .A1(n18149), .A2(n17900), .A3(n17899), .ZN(n17905) );
  NOR2_X1 U21010 ( .A1(n18639), .A2(n17901), .ZN(n17902) );
  AOI221_X1 U21011 ( .B1(n17903), .B2(n17905), .C1(n17902), .C2(n17905), .A(
        n9736), .ZN(n17913) );
  AOI21_X1 U21012 ( .B1(n9908), .B2(n17905), .A(n17904), .ZN(n17906) );
  AOI22_X1 U21013 ( .A1(n17918), .A2(n17907), .B1(n17913), .B2(n17906), .ZN(
        n17909) );
  OAI211_X1 U21014 ( .C1(n17910), .C2(n18078), .A(n17909), .B(n17908), .ZN(
        P3_U2838) );
  NAND2_X1 U21015 ( .A1(n9736), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17916) );
  NOR3_X1 U21016 ( .A1(n18149), .A2(n17912), .A3(n17911), .ZN(n17914) );
  OAI21_X1 U21017 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17914), .A(
        n17913), .ZN(n17915) );
  OAI211_X1 U21018 ( .C1(n17917), .C2(n18078), .A(n17916), .B(n17915), .ZN(
        P3_U2839) );
  NAND2_X1 U21019 ( .A1(n17919), .A2(n17918), .ZN(n17953) );
  OAI22_X1 U21020 ( .A1(n17921), .A2(n17953), .B1(n17920), .B2(n18170), .ZN(
        n17932) );
  AOI22_X1 U21021 ( .A1(n17998), .A2(n17999), .B1(n18000), .B2(n18001), .ZN(
        n17939) );
  NAND2_X1 U21022 ( .A1(n18658), .A2(n18028), .ZN(n18054) );
  INV_X1 U21023 ( .A(n18054), .ZN(n18031) );
  INV_X1 U21024 ( .A(n17965), .ZN(n17922) );
  AOI21_X1 U21025 ( .B1(n17922), .B2(n17949), .A(n18643), .ZN(n17923) );
  AOI221_X1 U21026 ( .B1(n17941), .B2(n18639), .C1(n17966), .C2(n18639), .A(
        n17923), .ZN(n17948) );
  OAI21_X1 U21027 ( .B1(n17924), .B2(n18031), .A(n17948), .ZN(n17925) );
  AOI21_X1 U21028 ( .B1(n18628), .B2(n17926), .A(n17925), .ZN(n17937) );
  INV_X1 U21029 ( .A(n17938), .ZN(n17928) );
  NOR2_X1 U21030 ( .A1(n18628), .A2(n18639), .ZN(n18063) );
  INV_X1 U21031 ( .A(n18063), .ZN(n17989) );
  AOI22_X1 U21032 ( .A1(n18639), .A2(n17928), .B1(n17927), .B2(n17989), .ZN(
        n17930) );
  NAND4_X1 U21033 ( .A1(n17939), .A2(n17937), .A3(n17930), .A4(n17929), .ZN(
        n17931) );
  AOI22_X1 U21034 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18149), .B1(
        n17932), .B2(n17931), .ZN(n17934) );
  OAI211_X1 U21035 ( .C1(n17935), .C2(n18078), .A(n17934), .B(n17933), .ZN(
        P3_U2840) );
  AOI22_X1 U21036 ( .A1(n9736), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18073), 
        .B2(n17936), .ZN(n17945) );
  OAI21_X1 U21037 ( .B1(n17947), .B2(n17938), .A(n17937), .ZN(n17943) );
  OAI21_X1 U21038 ( .B1(n17941), .B2(n17940), .A(n18641), .ZN(n17942) );
  NAND2_X1 U21039 ( .A1(n17991), .A2(n17942), .ZN(n17951) );
  OAI211_X1 U21040 ( .C1(n17943), .C2(n17951), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18169), .ZN(n17944) );
  OAI211_X1 U21041 ( .C1(n17946), .C2(n17953), .A(n17945), .B(n17944), .ZN(
        P3_U2841) );
  INV_X1 U21042 ( .A(n17947), .ZN(n18153) );
  NAND2_X1 U21043 ( .A1(n18153), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17952) );
  OAI21_X1 U21044 ( .B1(n17949), .B2(n18031), .A(n17948), .ZN(n17950) );
  OAI21_X1 U21045 ( .B1(n17951), .B2(n17950), .A(n18169), .ZN(n17963) );
  OAI21_X1 U21046 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17952), .A(
        n17963), .ZN(n17955) );
  INV_X1 U21047 ( .A(n17953), .ZN(n17959) );
  AOI22_X1 U21048 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17955), .B1(
        n17959), .B2(n17954), .ZN(n17957) );
  OAI211_X1 U21049 ( .C1(n17958), .C2(n18078), .A(n17957), .B(n17956), .ZN(
        P3_U2842) );
  AOI22_X1 U21050 ( .A1(n18073), .A2(n17960), .B1(n17959), .B2(n17964), .ZN(
        n17962) );
  OAI211_X1 U21051 ( .C1(n17964), .C2(n17963), .A(n17962), .B(n17961), .ZN(
        P3_U2843) );
  NOR3_X1 U21052 ( .A1(n18141), .A2(n17992), .A3(n17965), .ZN(n17969) );
  AOI222_X1 U21053 ( .A1(n18639), .A2(n17967), .B1(n18639), .B2(n17966), .C1(
        n17967), .C2(n18054), .ZN(n17968) );
  OAI211_X1 U21054 ( .C1(n18139), .C2(n17969), .A(n17991), .B(n17968), .ZN(
        n17981) );
  OAI221_X1 U21055 ( .B1(n17981), .B2(n17970), .C1(n17981), .C2(n18084), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17980) );
  OAI22_X1 U21056 ( .A1(n18144), .A2(n18659), .B1(n18083), .B2(n18137), .ZN(
        n18126) );
  NAND2_X1 U21057 ( .A1(n17971), .A2(n18126), .ZN(n18095) );
  NOR2_X1 U21058 ( .A1(n17972), .A2(n18095), .ZN(n18002) );
  OAI22_X1 U21059 ( .A1(n17974), .A2(n18658), .B1(n17973), .B2(n18028), .ZN(
        n17975) );
  NOR2_X1 U21060 ( .A1(n17976), .A2(n18076), .ZN(n17993) );
  AOI22_X1 U21061 ( .A1(n18073), .A2(n17978), .B1(n17993), .B2(n17977), .ZN(
        n17979) );
  OAI221_X1 U21062 ( .B1(n9736), .B2(n17980), .C1(n18169), .C2(n18746), .A(
        n17979), .ZN(P3_U2844) );
  NAND2_X1 U21063 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17981), .ZN(
        n17985) );
  INV_X1 U21064 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18744) );
  AOI22_X1 U21065 ( .A1(n18073), .A2(n17983), .B1(n17993), .B2(n17982), .ZN(
        n17984) );
  OAI221_X1 U21066 ( .B1(n9736), .B2(n17985), .C1(n18169), .C2(n18744), .A(
        n17984), .ZN(P3_U2845) );
  AOI21_X1 U21067 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18057), .A(
        n17986), .ZN(n17988) );
  OAI22_X1 U21068 ( .A1(n18643), .A2(n18013), .B1(n17987), .B2(n18659), .ZN(
        n18051) );
  AOI211_X1 U21069 ( .C1(n17990), .C2(n17989), .A(n17988), .B(n18051), .ZN(
        n18003) );
  AOI221_X1 U21070 ( .B1(n9908), .B2(n17991), .C1(n18003), .C2(n17991), .A(
        n9736), .ZN(n17994) );
  AOI22_X1 U21071 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17994), .B1(
        n17993), .B2(n17992), .ZN(n17996) );
  OAI211_X1 U21072 ( .C1(n17997), .C2(n18078), .A(n17996), .B(n17995), .ZN(
        P3_U2846) );
  NAND2_X1 U21073 ( .A1(n17999), .A2(n17998), .ZN(n18008) );
  NAND2_X1 U21074 ( .A1(n18001), .A2(n18000), .ZN(n18006) );
  AND2_X1 U21075 ( .A1(n18015), .A2(n18002), .ZN(n18017) );
  AOI21_X1 U21076 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18017), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18004) );
  OAI222_X1 U21077 ( .A1(n18008), .A2(n18007), .B1(n18006), .B2(n18005), .C1(
        n18004), .C2(n18003), .ZN(n18009) );
  AOI22_X1 U21078 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18149), .B1(
        n18154), .B2(n18009), .ZN(n18011) );
  OAI211_X1 U21079 ( .C1(n18078), .C2(n18012), .A(n18011), .B(n18010), .ZN(
        P3_U2847) );
  NAND2_X1 U21080 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18013), .ZN(
        n18052) );
  AOI221_X1 U21081 ( .B1(n18014), .B2(n18641), .C1(n18052), .C2(n18641), .A(
        n18051), .ZN(n18030) );
  OAI21_X1 U21082 ( .B1(n9908), .B2(n18015), .A(n18030), .ZN(n18016) );
  OAI221_X1 U21083 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18017), 
        .C1(n18019), .C2(n18016), .A(n18154), .ZN(n18018) );
  OAI21_X1 U21084 ( .B1(n18155), .B2(n18019), .A(n18018), .ZN(n18020) );
  AOI21_X1 U21085 ( .B1(n9736), .B2(P3_REIP_REG_14__SCAN_IN), .A(n18020), .ZN(
        n18024) );
  AOI22_X1 U21086 ( .A1(n18082), .A2(n18022), .B1(n18166), .B2(n18021), .ZN(
        n18023) );
  OAI211_X1 U21087 ( .C1(n18078), .C2(n18025), .A(n18024), .B(n18023), .ZN(
        P3_U2848) );
  AOI21_X1 U21088 ( .B1(n18628), .B2(n18026), .A(n18048), .ZN(n18043) );
  OAI22_X1 U21089 ( .A1(n18029), .A2(n18028), .B1(n18658), .B2(n18027), .ZN(
        n18050) );
  AOI22_X1 U21090 ( .A1(n18639), .A2(n18035), .B1(n18628), .B2(n18055), .ZN(
        n18056) );
  OAI211_X1 U21091 ( .C1(n18032), .C2(n18031), .A(n18056), .B(n18030), .ZN(
        n18033) );
  NOR2_X1 U21092 ( .A1(n18050), .A2(n18033), .ZN(n18042) );
  OAI211_X1 U21093 ( .C1(n18063), .C2(n18043), .A(n18154), .B(n18042), .ZN(
        n18034) );
  NAND2_X1 U21094 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18034), .ZN(
        n18039) );
  NOR2_X1 U21095 ( .A1(n18035), .A2(n18076), .ZN(n18040) );
  AOI22_X1 U21096 ( .A1(n18073), .A2(n18037), .B1(n18036), .B2(n18040), .ZN(
        n18038) );
  OAI221_X1 U21097 ( .B1(n9736), .B2(n18039), .C1(n18169), .C2(n18738), .A(
        n18038), .ZN(P3_U2849) );
  AOI21_X1 U21098 ( .B1(n18154), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18040), .ZN(n18041) );
  AOI21_X1 U21099 ( .B1(n18043), .B2(n18042), .A(n18041), .ZN(n18044) );
  AOI21_X1 U21100 ( .B1(n18073), .B2(n18045), .A(n18044), .ZN(n18047) );
  OAI211_X1 U21101 ( .C1(n18155), .C2(n18048), .A(n18047), .B(n18046), .ZN(
        P3_U2850) );
  AOI22_X1 U21102 ( .A1(n9736), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18073), 
        .B2(n18049), .ZN(n18060) );
  AOI211_X1 U21103 ( .C1(n18641), .C2(n18052), .A(n18051), .B(n18050), .ZN(
        n18070) );
  OAI211_X1 U21104 ( .C1(n18057), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18070), .B(n18155), .ZN(n18053) );
  AOI21_X1 U21105 ( .B1(n18055), .B2(n18054), .A(n18053), .ZN(n18064) );
  OAI211_X1 U21106 ( .C1(n18057), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18056), .B(n18064), .ZN(n18058) );
  NAND3_X1 U21107 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18169), .A3(
        n18058), .ZN(n18059) );
  OAI211_X1 U21108 ( .C1(n18061), .C2(n18076), .A(n18060), .B(n18059), .ZN(
        P3_U2851) );
  AOI221_X1 U21109 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18064), .C1(
        n18063), .C2(n18064), .A(n18062), .ZN(n18066) );
  NOR3_X1 U21110 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18069), .A3(
        n18076), .ZN(n18065) );
  AOI221_X1 U21111 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n9736), .C1(n18066), 
        .C2(n18169), .A(n18065), .ZN(n18067) );
  OAI21_X1 U21112 ( .B1(n18068), .B2(n18078), .A(n18067), .ZN(P3_U2852) );
  AOI211_X1 U21113 ( .C1(n18154), .C2(n18070), .A(n9736), .B(n18069), .ZN(
        n18071) );
  AOI21_X1 U21114 ( .B1(n18073), .B2(n18072), .A(n18071), .ZN(n18075) );
  OAI211_X1 U21115 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18076), .A(
        n18075), .B(n18074), .ZN(P3_U2853) );
  OAI22_X1 U21116 ( .A1(n18079), .A2(n18078), .B1(n18130), .B2(n18077), .ZN(
        n18080) );
  AOI21_X1 U21117 ( .B1(n18082), .B2(n18081), .A(n18080), .ZN(n18092) );
  AOI22_X1 U21118 ( .A1(n18639), .A2(n18144), .B1(n18084), .B2(n18083), .ZN(
        n18086) );
  NAND3_X1 U21119 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18086), .A3(
        n18085), .ZN(n18132) );
  NOR2_X1 U21120 ( .A1(n18087), .A2(n18132), .ZN(n18102) );
  AOI21_X1 U21121 ( .B1(n18088), .B2(n18102), .A(n18156), .ZN(n18097) );
  OAI21_X1 U21122 ( .B1(n18149), .B2(n18097), .A(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18090) );
  NAND3_X1 U21123 ( .A1(n18154), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18126), .ZN(n18125) );
  NOR2_X1 U21124 ( .A1(n18087), .A2(n18125), .ZN(n18105) );
  NAND3_X1 U21125 ( .A1(n18088), .A2(n18105), .A3(n21143), .ZN(n18089) );
  NAND4_X1 U21126 ( .A1(n18092), .A2(n18091), .A3(n18090), .A4(n18089), .ZN(
        P3_U2854) );
  AOI21_X1 U21127 ( .B1(n18149), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18093), .ZN(n18100) );
  OAI21_X1 U21128 ( .B1(n18104), .B2(n18095), .A(n18094), .ZN(n18096) );
  AOI22_X1 U21129 ( .A1(n18166), .A2(n18098), .B1(n18097), .B2(n18096), .ZN(
        n18099) );
  OAI211_X1 U21130 ( .C1(n18162), .C2(n18101), .A(n18100), .B(n18099), .ZN(
        P3_U2855) );
  OAI21_X1 U21131 ( .B1(n18102), .B2(n18156), .A(n18155), .ZN(n18112) );
  AOI22_X1 U21132 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18112), .B1(
        n9736), .B2(P3_REIP_REG_6__SCAN_IN), .ZN(n18108) );
  INV_X1 U21133 ( .A(n18103), .ZN(n18106) );
  AOI22_X1 U21134 ( .A1(n18106), .A2(n18168), .B1(n18105), .B2(n18104), .ZN(
        n18107) );
  OAI211_X1 U21135 ( .C1(n18130), .C2(n18109), .A(n18108), .B(n18107), .ZN(
        P3_U2856) );
  INV_X1 U21136 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18124) );
  NOR2_X1 U21137 ( .A1(n18124), .A2(n18125), .ZN(n18114) );
  OAI22_X1 U21138 ( .A1(n18169), .A2(n18722), .B1(n18130), .B2(n18110), .ZN(
        n18111) );
  AOI221_X1 U21139 ( .B1(n18114), .B2(n18113), .C1(n18112), .C2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n18111), .ZN(n18115) );
  OAI21_X1 U21140 ( .B1(n18162), .B2(n18116), .A(n18115), .ZN(P3_U2857) );
  AOI21_X1 U21141 ( .B1(n18117), .B2(n18132), .A(n18149), .ZN(n18123) );
  INV_X1 U21142 ( .A(n18118), .ZN(n18121) );
  OAI22_X1 U21143 ( .A1(n18169), .A2(n20983), .B1(n18162), .B2(n18119), .ZN(
        n18120) );
  AOI21_X1 U21144 ( .B1(n18166), .B2(n18121), .A(n18120), .ZN(n18122) );
  OAI221_X1 U21145 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18125), .C1(
        n18124), .C2(n18123), .A(n18122), .ZN(P3_U2858) );
  OAI21_X1 U21146 ( .B1(n18126), .B2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n18154), .ZN(n18127) );
  INV_X1 U21147 ( .A(n18127), .ZN(n18133) );
  OAI22_X1 U21148 ( .A1(n18130), .A2(n18129), .B1(n18162), .B2(n18128), .ZN(
        n18131) );
  AOI21_X1 U21149 ( .B1(n18133), .B2(n18132), .A(n18131), .ZN(n18135) );
  OAI211_X1 U21150 ( .C1(n18155), .C2(n18136), .A(n18135), .B(n18134), .ZN(
        P3_U2859) );
  INV_X1 U21151 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18798) );
  OR2_X1 U21152 ( .A1(n18798), .A2(n18137), .ZN(n18143) );
  NAND2_X1 U21153 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18138) );
  OAI22_X1 U21154 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18139), .B1(
        n18659), .B2(n18138), .ZN(n18140) );
  NOR2_X1 U21155 ( .A1(n18141), .A2(n18140), .ZN(n18142) );
  MUX2_X1 U21156 ( .A(n18143), .B(n18142), .S(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n18146) );
  NAND2_X1 U21157 ( .A1(n18639), .A2(n18144), .ZN(n18145) );
  OAI211_X1 U21158 ( .C1(n18658), .C2(n18147), .A(n18146), .B(n18145), .ZN(
        n18148) );
  AOI22_X1 U21159 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18149), .B1(
        n18154), .B2(n18148), .ZN(n18151) );
  OAI211_X1 U21160 ( .C1(n18152), .C2(n18162), .A(n18151), .B(n18150), .ZN(
        P3_U2860) );
  NAND3_X1 U21161 ( .A1(n18154), .A2(n18153), .A3(n18796), .ZN(n18172) );
  AOI21_X1 U21162 ( .B1(n18155), .B2(n18172), .A(n18798), .ZN(n18158) );
  AOI211_X1 U21163 ( .C1(n18643), .C2(n18796), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18156), .ZN(n18157) );
  AOI211_X1 U21164 ( .C1(n18166), .C2(n18159), .A(n18158), .B(n18157), .ZN(
        n18161) );
  NAND2_X1 U21165 ( .A1(n9736), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18160) );
  OAI211_X1 U21166 ( .C1(n18163), .C2(n18162), .A(n18161), .B(n18160), .ZN(
        P3_U2861) );
  AND2_X1 U21167 ( .A1(n9736), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18164) );
  AOI221_X1 U21168 ( .B1(n18168), .B2(n18167), .C1(n18166), .C2(n18165), .A(
        n18164), .ZN(n18173) );
  OAI211_X1 U21169 ( .C1(n18628), .C2(n18170), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n18169), .ZN(n18171) );
  NAND3_X1 U21170 ( .A1(n18173), .A2(n18172), .A3(n18171), .ZN(P3_U2862) );
  AOI211_X1 U21171 ( .C1(n18175), .C2(n18174), .A(n18687), .B(n20974), .ZN(
        n18680) );
  OAI21_X1 U21172 ( .B1(n18680), .B2(n18226), .A(n18180), .ZN(n18176) );
  OAI221_X1 U21173 ( .B1(n18477), .B2(n18829), .C1(n18477), .C2(n18180), .A(
        n18176), .ZN(P3_U2863) );
  INV_X1 U21174 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18664) );
  NAND2_X1 U21175 ( .A1(n18664), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18332) );
  NAND2_X1 U21176 ( .A1(n21113), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18452) );
  INV_X1 U21177 ( .A(n18452), .ZN(n18454) );
  NAND2_X1 U21178 ( .A1(n18267), .A2(n18454), .ZN(n18478) );
  AND2_X1 U21179 ( .A1(n18332), .A2(n18478), .ZN(n18178) );
  OAI22_X1 U21180 ( .A1(n18179), .A2(n18664), .B1(n18178), .B2(n18177), .ZN(
        P3_U2866) );
  NOR2_X1 U21181 ( .A1(n18665), .A2(n18180), .ZN(P3_U2867) );
  NAND2_X1 U21182 ( .A1(n18182), .A2(n18181), .ZN(n18221) );
  NOR2_X1 U21183 ( .A1(n18183), .A2(n18221), .ZN(n18428) );
  INV_X1 U21184 ( .A(n18428), .ZN(n18570) );
  NAND2_X1 U21185 ( .A1(n18646), .A2(n18477), .ZN(n18647) );
  NAND2_X1 U21186 ( .A1(n21113), .A2(n18664), .ZN(n18245) );
  NOR2_X2 U21187 ( .A1(n18647), .A2(n18245), .ZN(n18280) );
  INV_X1 U21188 ( .A(n18280), .ZN(n18287) );
  NOR2_X2 U21189 ( .A1(n18219), .A2(n19050), .ZN(n18567) );
  NOR2_X1 U21190 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18646), .ZN(
        n18186) );
  NAND2_X1 U21191 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18526) );
  NOR2_X2 U21192 ( .A1(n18425), .A2(n18526), .ZN(n18554) );
  NOR2_X2 U21193 ( .A1(n18334), .A2(n18184), .ZN(n18562) );
  NOR2_X1 U21194 ( .A1(n18664), .A2(n18185), .ZN(n18564) );
  NAND2_X1 U21195 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18564), .ZN(
        n18588) );
  INV_X1 U21196 ( .A(n18588), .ZN(n18614) );
  NOR2_X1 U21197 ( .A1(n18614), .A2(n18280), .ZN(n18246) );
  NOR2_X1 U21198 ( .A1(n9722), .A2(n18246), .ZN(n18220) );
  AOI22_X1 U21199 ( .A1(n18567), .A2(n18554), .B1(n18562), .B2(n18220), .ZN(
        n18190) );
  NOR2_X1 U21200 ( .A1(n18477), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18401) );
  NOR2_X1 U21201 ( .A1(n18186), .A2(n18401), .ZN(n18527) );
  NOR2_X1 U21202 ( .A1(n18527), .A2(n18526), .ZN(n18188) );
  AOI211_X1 U21203 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18246), .B(n18334), .ZN(
        n18187) );
  AOI21_X1 U21204 ( .B1(n18188), .B2(n18566), .A(n18187), .ZN(n18223) );
  NOR2_X2 U21205 ( .A1(n19206), .A2(n18219), .ZN(n18561) );
  NOR2_X1 U21206 ( .A1(n18526), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18565) );
  INV_X1 U21207 ( .A(n18565), .ZN(n18502) );
  NOR2_X2 U21208 ( .A1(n18477), .A2(n18502), .ZN(n18596) );
  AOI22_X1 U21209 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18223), .B1(
        n18561), .B2(n18596), .ZN(n18189) );
  OAI211_X1 U21210 ( .C1(n18570), .C2(n18287), .A(n18190), .B(n18189), .ZN(
        P3_U2868) );
  NAND2_X1 U21211 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18566), .ZN(n18509) );
  INV_X1 U21212 ( .A(n18596), .ZN(n18619) );
  NOR2_X2 U21213 ( .A1(n18334), .A2(n18191), .ZN(n18571) );
  INV_X1 U21214 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n18192) );
  NOR2_X2 U21215 ( .A1(n18219), .A2(n18192), .ZN(n18573) );
  AOI22_X1 U21216 ( .A1(n18571), .A2(n18220), .B1(n18573), .B2(n18554), .ZN(
        n18194) );
  NOR2_X1 U21217 ( .A1(n18835), .A2(n18221), .ZN(n18506) );
  AOI22_X1 U21218 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18223), .B1(
        n18506), .B2(n18280), .ZN(n18193) );
  OAI211_X1 U21219 ( .C1(n18509), .C2(n18619), .A(n18194), .B(n18193), .ZN(
        P3_U2869) );
  NOR2_X1 U21220 ( .A1(n18219), .A2(n18195), .ZN(n18536) );
  INV_X1 U21221 ( .A(n18536), .ZN(n18582) );
  NOR2_X2 U21222 ( .A1(n18334), .A2(n18196), .ZN(n18578) );
  AND2_X1 U21223 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18566), .ZN(n18577) );
  AOI22_X1 U21224 ( .A1(n18578), .A2(n18220), .B1(n18577), .B2(n18596), .ZN(
        n18199) );
  NOR2_X1 U21225 ( .A1(n18197), .A2(n18221), .ZN(n18579) );
  AOI22_X1 U21226 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18223), .B1(
        n18579), .B2(n18280), .ZN(n18198) );
  OAI211_X1 U21227 ( .C1(n18582), .C2(n18543), .A(n18199), .B(n18198), .ZN(
        P3_U2870) );
  NOR2_X1 U21228 ( .A1(n18200), .A2(n18221), .ZN(n18436) );
  INV_X1 U21229 ( .A(n18436), .ZN(n18589) );
  NAND2_X1 U21230 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18566), .ZN(n18439) );
  NOR2_X2 U21231 ( .A1(n18334), .A2(n18201), .ZN(n18583) );
  AOI22_X1 U21232 ( .A1(n18584), .A2(n18596), .B1(n18583), .B2(n18220), .ZN(
        n18204) );
  NOR2_X2 U21233 ( .A1(n18219), .A2(n18202), .ZN(n18585) );
  AOI22_X1 U21234 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18223), .B1(
        n18585), .B2(n18554), .ZN(n18203) );
  OAI211_X1 U21235 ( .C1(n18589), .C2(n18287), .A(n18204), .B(n18203), .ZN(
        P3_U2871) );
  NOR2_X1 U21236 ( .A1(n19230), .A2(n18219), .ZN(n18488) );
  INV_X1 U21237 ( .A(n18488), .ZN(n18595) );
  NOR2_X2 U21238 ( .A1(n18334), .A2(n18205), .ZN(n18591) );
  NAND2_X1 U21239 ( .A1(n18566), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18491) );
  INV_X1 U21240 ( .A(n18491), .ZN(n18590) );
  AOI22_X1 U21241 ( .A1(n18591), .A2(n18220), .B1(n18590), .B2(n18554), .ZN(
        n18208) );
  NOR2_X2 U21242 ( .A1(n18206), .A2(n18221), .ZN(n18592) );
  AOI22_X1 U21243 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18223), .B1(
        n18592), .B2(n18280), .ZN(n18207) );
  OAI211_X1 U21244 ( .C1(n18595), .C2(n18619), .A(n18208), .B(n18207), .ZN(
        P3_U2872) );
  NAND2_X1 U21245 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18566), .ZN(n18603) );
  NOR2_X2 U21246 ( .A1(n18334), .A2(n18209), .ZN(n18598) );
  NAND2_X1 U21247 ( .A1(n18566), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18468) );
  INV_X1 U21248 ( .A(n18468), .ZN(n18597) );
  AOI22_X1 U21249 ( .A1(n18598), .A2(n18220), .B1(n18597), .B2(n18554), .ZN(
        n18212) );
  NOR2_X2 U21250 ( .A1(n18210), .A2(n18221), .ZN(n18599) );
  AOI22_X1 U21251 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18223), .B1(
        n18599), .B2(n18280), .ZN(n18211) );
  OAI211_X1 U21252 ( .C1(n18603), .C2(n18619), .A(n18212), .B(n18211), .ZN(
        P3_U2873) );
  NOR2_X1 U21253 ( .A1(n18213), .A2(n18219), .ZN(n18548) );
  NAND2_X1 U21254 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18566), .ZN(n18551) );
  INV_X1 U21255 ( .A(n18551), .ZN(n18605) );
  NOR2_X2 U21256 ( .A1(n18214), .A2(n18334), .ZN(n18604) );
  AOI22_X1 U21257 ( .A1(n18605), .A2(n18596), .B1(n18604), .B2(n18220), .ZN(
        n18217) );
  NOR2_X2 U21258 ( .A1(n18215), .A2(n18221), .ZN(n18606) );
  AOI22_X1 U21259 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18223), .B1(
        n18606), .B2(n18280), .ZN(n18216) );
  OAI211_X1 U21260 ( .C1(n18609), .C2(n18543), .A(n18217), .B(n18216), .ZN(
        P3_U2874) );
  NAND2_X1 U21261 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18566), .ZN(n18559) );
  NOR2_X2 U21262 ( .A1(n18218), .A2(n18334), .ZN(n18611) );
  NOR2_X2 U21263 ( .A1(n19254), .A2(n18219), .ZN(n18552) );
  AOI22_X1 U21264 ( .A1(n18611), .A2(n18220), .B1(n18552), .B2(n18554), .ZN(
        n18225) );
  NOR2_X2 U21265 ( .A1(n18222), .A2(n18221), .ZN(n18615) );
  AOI22_X1 U21266 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18223), .B1(
        n18615), .B2(n18280), .ZN(n18224) );
  OAI211_X1 U21267 ( .C1(n18559), .C2(n18619), .A(n18225), .B(n18224), .ZN(
        P3_U2875) );
  INV_X1 U21268 ( .A(n18245), .ZN(n18266) );
  NAND2_X1 U21269 ( .A1(n18401), .A2(n18266), .ZN(n18309) );
  AOI22_X1 U21270 ( .A1(n18562), .A2(n18241), .B1(n18561), .B2(n18554), .ZN(
        n18228) );
  NOR2_X1 U21271 ( .A1(n18334), .A2(n18226), .ZN(n18563) );
  AND2_X1 U21272 ( .A1(n18646), .A2(n18563), .ZN(n18403) );
  AOI22_X1 U21273 ( .A1(n18566), .A2(n18564), .B1(n18266), .B2(n18403), .ZN(
        n18242) );
  AOI22_X1 U21274 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18242), .B1(
        n18567), .B2(n18614), .ZN(n18227) );
  OAI211_X1 U21275 ( .C1(n18570), .C2(n18309), .A(n18228), .B(n18227), .ZN(
        P3_U2876) );
  AOI22_X1 U21276 ( .A1(n18571), .A2(n18241), .B1(n18573), .B2(n18614), .ZN(
        n18230) );
  INV_X1 U21277 ( .A(n18509), .ZN(n18572) );
  AOI22_X1 U21278 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18242), .B1(
        n18572), .B2(n18554), .ZN(n18229) );
  OAI211_X1 U21279 ( .C1(n18576), .C2(n18309), .A(n18230), .B(n18229), .ZN(
        P3_U2877) );
  AOI22_X1 U21280 ( .A1(n18536), .A2(n18614), .B1(n18578), .B2(n18241), .ZN(
        n18232) );
  AOI22_X1 U21281 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18242), .B1(
        n18577), .B2(n18554), .ZN(n18231) );
  OAI211_X1 U21282 ( .C1(n18539), .C2(n18309), .A(n18232), .B(n18231), .ZN(
        P3_U2878) );
  AOI22_X1 U21283 ( .A1(n18584), .A2(n18554), .B1(n18583), .B2(n18241), .ZN(
        n18234) );
  AOI22_X1 U21284 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18242), .B1(
        n18585), .B2(n18614), .ZN(n18233) );
  OAI211_X1 U21285 ( .C1(n18589), .C2(n18309), .A(n18234), .B(n18233), .ZN(
        P3_U2879) );
  AOI22_X1 U21286 ( .A1(n18591), .A2(n18241), .B1(n18590), .B2(n18614), .ZN(
        n18236) );
  INV_X1 U21287 ( .A(n18309), .ZN(n18298) );
  AOI22_X1 U21288 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18242), .B1(
        n18592), .B2(n18298), .ZN(n18235) );
  OAI211_X1 U21289 ( .C1(n18595), .C2(n18543), .A(n18236), .B(n18235), .ZN(
        P3_U2880) );
  AOI22_X1 U21290 ( .A1(n18598), .A2(n18241), .B1(n18597), .B2(n18614), .ZN(
        n18238) );
  AOI22_X1 U21291 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18242), .B1(
        n18599), .B2(n18298), .ZN(n18237) );
  OAI211_X1 U21292 ( .C1(n18603), .C2(n18543), .A(n18238), .B(n18237), .ZN(
        P3_U2881) );
  AOI22_X1 U21293 ( .A1(n18605), .A2(n18554), .B1(n18604), .B2(n18241), .ZN(
        n18240) );
  AOI22_X1 U21294 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18242), .B1(
        n18606), .B2(n18298), .ZN(n18239) );
  OAI211_X1 U21295 ( .C1(n18609), .C2(n18588), .A(n18240), .B(n18239), .ZN(
        P3_U2882) );
  AOI22_X1 U21296 ( .A1(n18611), .A2(n18241), .B1(n18552), .B2(n18614), .ZN(
        n18244) );
  AOI22_X1 U21297 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18242), .B1(
        n18615), .B2(n18298), .ZN(n18243) );
  OAI211_X1 U21298 ( .C1(n18559), .C2(n18543), .A(n18244), .B(n18243), .ZN(
        P3_U2883) );
  NOR2_X2 U21299 ( .A1(n18425), .A2(n18245), .ZN(n18328) );
  INV_X1 U21300 ( .A(n18328), .ZN(n18324) );
  NOR2_X1 U21301 ( .A1(n18298), .A2(n18328), .ZN(n18288) );
  NOR2_X1 U21302 ( .A1(n9722), .A2(n18288), .ZN(n18262) );
  AOI22_X1 U21303 ( .A1(n18567), .A2(n18280), .B1(n18562), .B2(n18262), .ZN(
        n18249) );
  INV_X1 U21304 ( .A(n18334), .ZN(n18530) );
  OAI21_X1 U21305 ( .B1(n18246), .B2(n18528), .A(n18288), .ZN(n18247) );
  OAI211_X1 U21306 ( .C1(n18328), .C2(n18787), .A(n18530), .B(n18247), .ZN(
        n18263) );
  AOI22_X1 U21307 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18263), .B1(
        n18561), .B2(n18614), .ZN(n18248) );
  OAI211_X1 U21308 ( .C1(n18570), .C2(n18324), .A(n18249), .B(n18248), .ZN(
        P3_U2884) );
  AOI22_X1 U21309 ( .A1(n18572), .A2(n18614), .B1(n18571), .B2(n18262), .ZN(
        n18251) );
  AOI22_X1 U21310 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18263), .B1(
        n18573), .B2(n18280), .ZN(n18250) );
  OAI211_X1 U21311 ( .C1(n18576), .C2(n18324), .A(n18251), .B(n18250), .ZN(
        P3_U2885) );
  AOI22_X1 U21312 ( .A1(n18578), .A2(n18262), .B1(n18577), .B2(n18614), .ZN(
        n18253) );
  AOI22_X1 U21313 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18263), .B1(
        n18579), .B2(n18328), .ZN(n18252) );
  OAI211_X1 U21314 ( .C1(n18582), .C2(n18287), .A(n18253), .B(n18252), .ZN(
        P3_U2886) );
  AOI22_X1 U21315 ( .A1(n18584), .A2(n18614), .B1(n18583), .B2(n18262), .ZN(
        n18255) );
  AOI22_X1 U21316 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18263), .B1(
        n18585), .B2(n18280), .ZN(n18254) );
  OAI211_X1 U21317 ( .C1(n18589), .C2(n18324), .A(n18255), .B(n18254), .ZN(
        P3_U2887) );
  AOI22_X1 U21318 ( .A1(n18591), .A2(n18262), .B1(n18590), .B2(n18280), .ZN(
        n18257) );
  AOI22_X1 U21319 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18263), .B1(
        n18592), .B2(n18328), .ZN(n18256) );
  OAI211_X1 U21320 ( .C1(n18595), .C2(n18588), .A(n18257), .B(n18256), .ZN(
        P3_U2888) );
  INV_X1 U21321 ( .A(n18603), .ZN(n18465) );
  AOI22_X1 U21322 ( .A1(n18465), .A2(n18614), .B1(n18598), .B2(n18262), .ZN(
        n18259) );
  AOI22_X1 U21323 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18263), .B1(
        n18599), .B2(n18328), .ZN(n18258) );
  OAI211_X1 U21324 ( .C1(n18468), .C2(n18287), .A(n18259), .B(n18258), .ZN(
        P3_U2889) );
  AOI22_X1 U21325 ( .A1(n18605), .A2(n18614), .B1(n18604), .B2(n18262), .ZN(
        n18261) );
  AOI22_X1 U21326 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18263), .B1(
        n18606), .B2(n18328), .ZN(n18260) );
  OAI211_X1 U21327 ( .C1(n18609), .C2(n18287), .A(n18261), .B(n18260), .ZN(
        P3_U2890) );
  AOI22_X1 U21328 ( .A1(n18611), .A2(n18262), .B1(n18552), .B2(n18280), .ZN(
        n18265) );
  AOI22_X1 U21329 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18263), .B1(
        n18615), .B2(n18328), .ZN(n18264) );
  OAI211_X1 U21330 ( .C1(n18559), .C2(n18588), .A(n18265), .B(n18264), .ZN(
        P3_U2891) );
  NAND2_X1 U21331 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18266), .ZN(
        n18310) );
  NOR2_X2 U21332 ( .A1(n18477), .A2(n18310), .ZN(n18346) );
  NOR2_X1 U21333 ( .A1(n9722), .A2(n18310), .ZN(n18283) );
  AOI22_X1 U21334 ( .A1(n18567), .A2(n18298), .B1(n18562), .B2(n18283), .ZN(
        n18269) );
  OAI211_X1 U21335 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18267), .A(
        n18266), .B(n18563), .ZN(n18284) );
  AOI22_X1 U21336 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18284), .B1(
        n18561), .B2(n18280), .ZN(n18268) );
  OAI211_X1 U21337 ( .C1(n18570), .C2(n18355), .A(n18269), .B(n18268), .ZN(
        P3_U2892) );
  AOI22_X1 U21338 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18284), .B1(
        n18571), .B2(n18283), .ZN(n18271) );
  AOI22_X1 U21339 ( .A1(n18572), .A2(n18280), .B1(n18573), .B2(n18298), .ZN(
        n18270) );
  OAI211_X1 U21340 ( .C1(n18576), .C2(n18355), .A(n18271), .B(n18270), .ZN(
        P3_U2893) );
  AOI22_X1 U21341 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18284), .B1(
        n18578), .B2(n18283), .ZN(n18273) );
  AOI22_X1 U21342 ( .A1(n18536), .A2(n18298), .B1(n18577), .B2(n18280), .ZN(
        n18272) );
  OAI211_X1 U21343 ( .C1(n18539), .C2(n18355), .A(n18273), .B(n18272), .ZN(
        P3_U2894) );
  AOI22_X1 U21344 ( .A1(n18585), .A2(n18298), .B1(n18583), .B2(n18283), .ZN(
        n18275) );
  AOI22_X1 U21345 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18284), .B1(
        n18584), .B2(n18280), .ZN(n18274) );
  OAI211_X1 U21346 ( .C1(n18589), .C2(n18355), .A(n18275), .B(n18274), .ZN(
        P3_U2895) );
  AOI22_X1 U21347 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18284), .B1(
        n18591), .B2(n18283), .ZN(n18277) );
  AOI22_X1 U21348 ( .A1(n18592), .A2(n18346), .B1(n18590), .B2(n18298), .ZN(
        n18276) );
  OAI211_X1 U21349 ( .C1(n18595), .C2(n18287), .A(n18277), .B(n18276), .ZN(
        P3_U2896) );
  AOI22_X1 U21350 ( .A1(n18598), .A2(n18283), .B1(n18597), .B2(n18298), .ZN(
        n18279) );
  AOI22_X1 U21351 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18284), .B1(
        n18599), .B2(n18346), .ZN(n18278) );
  OAI211_X1 U21352 ( .C1(n18603), .C2(n18287), .A(n18279), .B(n18278), .ZN(
        P3_U2897) );
  AOI22_X1 U21353 ( .A1(n18605), .A2(n18280), .B1(n18604), .B2(n18283), .ZN(
        n18282) );
  AOI22_X1 U21354 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18284), .B1(
        n18606), .B2(n18346), .ZN(n18281) );
  OAI211_X1 U21355 ( .C1(n18609), .C2(n18309), .A(n18282), .B(n18281), .ZN(
        P3_U2898) );
  AOI22_X1 U21356 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18284), .B1(
        n18611), .B2(n18283), .ZN(n18286) );
  AOI22_X1 U21357 ( .A1(n18615), .A2(n18346), .B1(n18552), .B2(n18298), .ZN(
        n18285) );
  OAI211_X1 U21358 ( .C1(n18559), .C2(n18287), .A(n18286), .B(n18285), .ZN(
        P3_U2899) );
  NOR2_X2 U21359 ( .A1(n18647), .A2(n18332), .ZN(n18369) );
  AOI21_X1 U21360 ( .B1(n18355), .B2(n18378), .A(n9722), .ZN(n18305) );
  AOI22_X1 U21361 ( .A1(n18567), .A2(n18328), .B1(n18562), .B2(n18305), .ZN(
        n18291) );
  OAI21_X1 U21362 ( .B1(n18346), .B2(n18369), .A(n18530), .ZN(n18333) );
  OAI21_X1 U21363 ( .B1(n18288), .B2(n18219), .A(n18333), .ZN(n18289) );
  OAI21_X1 U21364 ( .B1(n18369), .B2(n18787), .A(n18289), .ZN(n18306) );
  AOI22_X1 U21365 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18306), .B1(
        n18561), .B2(n18298), .ZN(n18290) );
  OAI211_X1 U21366 ( .C1(n18570), .C2(n18378), .A(n18291), .B(n18290), .ZN(
        P3_U2900) );
  AOI22_X1 U21367 ( .A1(n18572), .A2(n18298), .B1(n18571), .B2(n18305), .ZN(
        n18293) );
  AOI22_X1 U21368 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18306), .B1(
        n18573), .B2(n18328), .ZN(n18292) );
  OAI211_X1 U21369 ( .C1(n18576), .C2(n18378), .A(n18293), .B(n18292), .ZN(
        P3_U2901) );
  AOI22_X1 U21370 ( .A1(n18578), .A2(n18305), .B1(n18577), .B2(n18298), .ZN(
        n18295) );
  AOI22_X1 U21371 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18306), .B1(
        n18579), .B2(n18369), .ZN(n18294) );
  OAI211_X1 U21372 ( .C1(n18582), .C2(n18324), .A(n18295), .B(n18294), .ZN(
        P3_U2902) );
  AOI22_X1 U21373 ( .A1(n18585), .A2(n18328), .B1(n18583), .B2(n18305), .ZN(
        n18297) );
  AOI22_X1 U21374 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18306), .B1(
        n18436), .B2(n18369), .ZN(n18296) );
  OAI211_X1 U21375 ( .C1(n18439), .C2(n18309), .A(n18297), .B(n18296), .ZN(
        P3_U2903) );
  AOI22_X1 U21376 ( .A1(n18488), .A2(n18298), .B1(n18591), .B2(n18305), .ZN(
        n18300) );
  AOI22_X1 U21377 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18306), .B1(
        n18592), .B2(n18369), .ZN(n18299) );
  OAI211_X1 U21378 ( .C1(n18491), .C2(n18324), .A(n18300), .B(n18299), .ZN(
        P3_U2904) );
  AOI22_X1 U21379 ( .A1(n18598), .A2(n18305), .B1(n18597), .B2(n18328), .ZN(
        n18302) );
  AOI22_X1 U21380 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18306), .B1(
        n18599), .B2(n18369), .ZN(n18301) );
  OAI211_X1 U21381 ( .C1(n18603), .C2(n18309), .A(n18302), .B(n18301), .ZN(
        P3_U2905) );
  AOI22_X1 U21382 ( .A1(n18548), .A2(n18328), .B1(n18604), .B2(n18305), .ZN(
        n18304) );
  AOI22_X1 U21383 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18306), .B1(
        n18606), .B2(n18369), .ZN(n18303) );
  OAI211_X1 U21384 ( .C1(n18551), .C2(n18309), .A(n18304), .B(n18303), .ZN(
        P3_U2906) );
  AOI22_X1 U21385 ( .A1(n18611), .A2(n18305), .B1(n18552), .B2(n18328), .ZN(
        n18308) );
  AOI22_X1 U21386 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18306), .B1(
        n18615), .B2(n18369), .ZN(n18307) );
  OAI211_X1 U21387 ( .C1(n18559), .C2(n18309), .A(n18308), .B(n18307), .ZN(
        P3_U2907) );
  INV_X1 U21388 ( .A(n18332), .ZN(n18358) );
  NAND2_X1 U21389 ( .A1(n18401), .A2(n18358), .ZN(n18400) );
  AOI22_X1 U21390 ( .A1(n18567), .A2(n18346), .B1(n18562), .B2(n18327), .ZN(
        n18313) );
  INV_X1 U21391 ( .A(n18310), .ZN(n18311) );
  AOI22_X1 U21392 ( .A1(n18566), .A2(n18311), .B1(n18403), .B2(n18358), .ZN(
        n18329) );
  AOI22_X1 U21393 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18329), .B1(
        n18561), .B2(n18328), .ZN(n18312) );
  OAI211_X1 U21394 ( .C1(n18570), .C2(n18400), .A(n18313), .B(n18312), .ZN(
        P3_U2908) );
  AOI22_X1 U21395 ( .A1(n18572), .A2(n18328), .B1(n18571), .B2(n18327), .ZN(
        n18315) );
  AOI22_X1 U21396 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18329), .B1(
        n18573), .B2(n18346), .ZN(n18314) );
  OAI211_X1 U21397 ( .C1(n18576), .C2(n18400), .A(n18315), .B(n18314), .ZN(
        P3_U2909) );
  AOI22_X1 U21398 ( .A1(n18578), .A2(n18327), .B1(n18577), .B2(n18328), .ZN(
        n18317) );
  AOI22_X1 U21399 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18329), .B1(
        n18536), .B2(n18346), .ZN(n18316) );
  OAI211_X1 U21400 ( .C1(n18539), .C2(n18400), .A(n18317), .B(n18316), .ZN(
        P3_U2910) );
  AOI22_X1 U21401 ( .A1(n18584), .A2(n18328), .B1(n18583), .B2(n18327), .ZN(
        n18319) );
  AOI22_X1 U21402 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18329), .B1(
        n18585), .B2(n18346), .ZN(n18318) );
  OAI211_X1 U21403 ( .C1(n18589), .C2(n18400), .A(n18319), .B(n18318), .ZN(
        P3_U2911) );
  AOI22_X1 U21404 ( .A1(n18591), .A2(n18327), .B1(n18590), .B2(n18346), .ZN(
        n18321) );
  INV_X1 U21405 ( .A(n18400), .ZN(n18393) );
  AOI22_X1 U21406 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18329), .B1(
        n18592), .B2(n18393), .ZN(n18320) );
  OAI211_X1 U21407 ( .C1(n18595), .C2(n18324), .A(n18321), .B(n18320), .ZN(
        P3_U2912) );
  AOI22_X1 U21408 ( .A1(n18598), .A2(n18327), .B1(n18597), .B2(n18346), .ZN(
        n18323) );
  AOI22_X1 U21409 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18329), .B1(
        n18599), .B2(n18393), .ZN(n18322) );
  OAI211_X1 U21410 ( .C1(n18603), .C2(n18324), .A(n18323), .B(n18322), .ZN(
        P3_U2913) );
  AOI22_X1 U21411 ( .A1(n18605), .A2(n18328), .B1(n18604), .B2(n18327), .ZN(
        n18326) );
  AOI22_X1 U21412 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18329), .B1(
        n18606), .B2(n18393), .ZN(n18325) );
  OAI211_X1 U21413 ( .C1(n18609), .C2(n18355), .A(n18326), .B(n18325), .ZN(
        P3_U2914) );
  INV_X1 U21414 ( .A(n18552), .ZN(n18620) );
  INV_X1 U21415 ( .A(n18559), .ZN(n18613) );
  AOI22_X1 U21416 ( .A1(n18613), .A2(n18328), .B1(n18611), .B2(n18327), .ZN(
        n18331) );
  AOI22_X1 U21417 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18329), .B1(
        n18615), .B2(n18393), .ZN(n18330) );
  OAI211_X1 U21418 ( .C1(n18620), .C2(n18355), .A(n18331), .B(n18330), .ZN(
        P3_U2915) );
  NOR2_X2 U21419 ( .A1(n18425), .A2(n18332), .ZN(n18417) );
  NOR2_X1 U21420 ( .A1(n18393), .A2(n18417), .ZN(n18379) );
  NOR2_X1 U21421 ( .A1(n9722), .A2(n18379), .ZN(n18351) );
  AOI22_X1 U21422 ( .A1(n18567), .A2(n18369), .B1(n18562), .B2(n18351), .ZN(
        n18337) );
  OAI22_X1 U21423 ( .A1(n18379), .A2(n18334), .B1(n18528), .B2(n18333), .ZN(
        n18335) );
  OAI21_X1 U21424 ( .B1(n18417), .B2(n18787), .A(n18335), .ZN(n18352) );
  AOI22_X1 U21425 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18352), .B1(
        n18561), .B2(n18346), .ZN(n18336) );
  OAI211_X1 U21426 ( .C1(n18570), .C2(n18424), .A(n18337), .B(n18336), .ZN(
        P3_U2916) );
  AOI22_X1 U21427 ( .A1(n18572), .A2(n18346), .B1(n18571), .B2(n18351), .ZN(
        n18339) );
  AOI22_X1 U21428 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18352), .B1(
        n18573), .B2(n18369), .ZN(n18338) );
  OAI211_X1 U21429 ( .C1(n18576), .C2(n18424), .A(n18339), .B(n18338), .ZN(
        P3_U2917) );
  AOI22_X1 U21430 ( .A1(n18578), .A2(n18351), .B1(n18577), .B2(n18346), .ZN(
        n18341) );
  AOI22_X1 U21431 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18352), .B1(
        n18579), .B2(n18417), .ZN(n18340) );
  OAI211_X1 U21432 ( .C1(n18582), .C2(n18378), .A(n18341), .B(n18340), .ZN(
        P3_U2918) );
  AOI22_X1 U21433 ( .A1(n18584), .A2(n18346), .B1(n18583), .B2(n18351), .ZN(
        n18343) );
  AOI22_X1 U21434 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18352), .B1(
        n18585), .B2(n18369), .ZN(n18342) );
  OAI211_X1 U21435 ( .C1(n18589), .C2(n18424), .A(n18343), .B(n18342), .ZN(
        P3_U2919) );
  AOI22_X1 U21436 ( .A1(n18488), .A2(n18346), .B1(n18591), .B2(n18351), .ZN(
        n18345) );
  AOI22_X1 U21437 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18352), .B1(
        n18592), .B2(n18417), .ZN(n18344) );
  OAI211_X1 U21438 ( .C1(n18491), .C2(n18378), .A(n18345), .B(n18344), .ZN(
        P3_U2920) );
  AOI22_X1 U21439 ( .A1(n18465), .A2(n18346), .B1(n18598), .B2(n18351), .ZN(
        n18348) );
  AOI22_X1 U21440 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18352), .B1(
        n18599), .B2(n18417), .ZN(n18347) );
  OAI211_X1 U21441 ( .C1(n18468), .C2(n18378), .A(n18348), .B(n18347), .ZN(
        P3_U2921) );
  AOI22_X1 U21442 ( .A1(n18548), .A2(n18369), .B1(n18604), .B2(n18351), .ZN(
        n18350) );
  AOI22_X1 U21443 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18352), .B1(
        n18606), .B2(n18417), .ZN(n18349) );
  OAI211_X1 U21444 ( .C1(n18551), .C2(n18355), .A(n18350), .B(n18349), .ZN(
        P3_U2922) );
  AOI22_X1 U21445 ( .A1(n18611), .A2(n18351), .B1(n18552), .B2(n18369), .ZN(
        n18354) );
  AOI22_X1 U21446 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18352), .B1(
        n18615), .B2(n18417), .ZN(n18353) );
  OAI211_X1 U21447 ( .C1(n18559), .C2(n18355), .A(n18354), .B(n18353), .ZN(
        P3_U2923) );
  NAND2_X1 U21448 ( .A1(n18664), .A2(n18356), .ZN(n18402) );
  NOR2_X2 U21449 ( .A1(n18477), .A2(n18402), .ZN(n18444) );
  NOR2_X1 U21450 ( .A1(n9722), .A2(n18402), .ZN(n18374) );
  AOI22_X1 U21451 ( .A1(n18562), .A2(n18374), .B1(n18561), .B2(n18369), .ZN(
        n18360) );
  AOI22_X1 U21452 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18451), .B1(n18646), 
        .B2(n18528), .ZN(n18357) );
  NAND3_X1 U21453 ( .A1(n18530), .A2(n18358), .A3(n18357), .ZN(n18375) );
  AOI22_X1 U21454 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18375), .B1(
        n18567), .B2(n18393), .ZN(n18359) );
  OAI211_X1 U21455 ( .C1(n18451), .C2(n18570), .A(n18360), .B(n18359), .ZN(
        P3_U2924) );
  AOI22_X1 U21456 ( .A1(n18572), .A2(n18369), .B1(n18571), .B2(n18374), .ZN(
        n18362) );
  AOI22_X1 U21457 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18375), .B1(
        n18573), .B2(n18393), .ZN(n18361) );
  OAI211_X1 U21458 ( .C1(n18451), .C2(n18576), .A(n18362), .B(n18361), .ZN(
        P3_U2925) );
  AOI22_X1 U21459 ( .A1(n18578), .A2(n18374), .B1(n18577), .B2(n18369), .ZN(
        n18364) );
  AOI22_X1 U21460 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18375), .B1(
        n18444), .B2(n18579), .ZN(n18363) );
  OAI211_X1 U21461 ( .C1(n18582), .C2(n18400), .A(n18364), .B(n18363), .ZN(
        P3_U2926) );
  AOI22_X1 U21462 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18375), .B1(
        n18583), .B2(n18374), .ZN(n18366) );
  AOI22_X1 U21463 ( .A1(n18444), .A2(n18436), .B1(n18585), .B2(n18393), .ZN(
        n18365) );
  OAI211_X1 U21464 ( .C1(n18439), .C2(n18378), .A(n18366), .B(n18365), .ZN(
        P3_U2927) );
  AOI22_X1 U21465 ( .A1(n18591), .A2(n18374), .B1(n18590), .B2(n18393), .ZN(
        n18368) );
  AOI22_X1 U21466 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18375), .B1(
        n18444), .B2(n18592), .ZN(n18367) );
  OAI211_X1 U21467 ( .C1(n18595), .C2(n18378), .A(n18368), .B(n18367), .ZN(
        P3_U2928) );
  AOI22_X1 U21468 ( .A1(n18465), .A2(n18369), .B1(n18598), .B2(n18374), .ZN(
        n18371) );
  AOI22_X1 U21469 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18375), .B1(
        n18444), .B2(n18599), .ZN(n18370) );
  OAI211_X1 U21470 ( .C1(n18468), .C2(n18400), .A(n18371), .B(n18370), .ZN(
        P3_U2929) );
  AOI22_X1 U21471 ( .A1(n18548), .A2(n18393), .B1(n18604), .B2(n18374), .ZN(
        n18373) );
  AOI22_X1 U21472 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18375), .B1(
        n18444), .B2(n18606), .ZN(n18372) );
  OAI211_X1 U21473 ( .C1(n18551), .C2(n18378), .A(n18373), .B(n18372), .ZN(
        P3_U2930) );
  AOI22_X1 U21474 ( .A1(n18611), .A2(n18374), .B1(n18552), .B2(n18393), .ZN(
        n18377) );
  AOI22_X1 U21475 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18375), .B1(
        n18444), .B2(n18615), .ZN(n18376) );
  OAI211_X1 U21476 ( .C1(n18559), .C2(n18378), .A(n18377), .B(n18376), .ZN(
        P3_U2931) );
  NOR2_X2 U21477 ( .A1(n18647), .A2(n18452), .ZN(n18473) );
  INV_X1 U21478 ( .A(n18473), .ZN(n18471) );
  NOR2_X1 U21479 ( .A1(n18473), .A2(n18444), .ZN(n18426) );
  NOR2_X1 U21480 ( .A1(n9722), .A2(n18426), .ZN(n18396) );
  AOI22_X1 U21481 ( .A1(n18562), .A2(n18396), .B1(n18561), .B2(n18393), .ZN(
        n18382) );
  AOI221_X1 U21482 ( .B1(n18379), .B2(n18451), .C1(n18528), .C2(n18451), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18380) );
  OAI21_X1 U21483 ( .B1(n18473), .B2(n18380), .A(n18530), .ZN(n18397) );
  AOI22_X1 U21484 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18397), .B1(
        n18567), .B2(n18417), .ZN(n18381) );
  OAI211_X1 U21485 ( .C1(n18471), .C2(n18570), .A(n18382), .B(n18381), .ZN(
        P3_U2932) );
  AOI22_X1 U21486 ( .A1(n18571), .A2(n18396), .B1(n18573), .B2(n18417), .ZN(
        n18384) );
  AOI22_X1 U21487 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18397), .B1(
        n18473), .B2(n18506), .ZN(n18383) );
  OAI211_X1 U21488 ( .C1(n18509), .C2(n18400), .A(n18384), .B(n18383), .ZN(
        P3_U2933) );
  AOI22_X1 U21489 ( .A1(n18536), .A2(n18417), .B1(n18578), .B2(n18396), .ZN(
        n18386) );
  AOI22_X1 U21490 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18397), .B1(
        n18577), .B2(n18393), .ZN(n18385) );
  OAI211_X1 U21491 ( .C1(n18471), .C2(n18539), .A(n18386), .B(n18385), .ZN(
        P3_U2934) );
  AOI22_X1 U21492 ( .A1(n18584), .A2(n18393), .B1(n18583), .B2(n18396), .ZN(
        n18388) );
  AOI22_X1 U21493 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18397), .B1(
        n18585), .B2(n18417), .ZN(n18387) );
  OAI211_X1 U21494 ( .C1(n18471), .C2(n18589), .A(n18388), .B(n18387), .ZN(
        P3_U2935) );
  AOI22_X1 U21495 ( .A1(n18488), .A2(n18393), .B1(n18591), .B2(n18396), .ZN(
        n18390) );
  AOI22_X1 U21496 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18397), .B1(
        n18473), .B2(n18592), .ZN(n18389) );
  OAI211_X1 U21497 ( .C1(n18491), .C2(n18424), .A(n18390), .B(n18389), .ZN(
        P3_U2936) );
  AOI22_X1 U21498 ( .A1(n18465), .A2(n18393), .B1(n18598), .B2(n18396), .ZN(
        n18392) );
  AOI22_X1 U21499 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18397), .B1(
        n18473), .B2(n18599), .ZN(n18391) );
  OAI211_X1 U21500 ( .C1(n18468), .C2(n18424), .A(n18392), .B(n18391), .ZN(
        P3_U2937) );
  AOI22_X1 U21501 ( .A1(n18605), .A2(n18393), .B1(n18604), .B2(n18396), .ZN(
        n18395) );
  AOI22_X1 U21502 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18397), .B1(
        n18473), .B2(n18606), .ZN(n18394) );
  OAI211_X1 U21503 ( .C1(n18609), .C2(n18424), .A(n18395), .B(n18394), .ZN(
        P3_U2938) );
  AOI22_X1 U21504 ( .A1(n18611), .A2(n18396), .B1(n18552), .B2(n18417), .ZN(
        n18399) );
  AOI22_X1 U21505 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18397), .B1(
        n18473), .B2(n18615), .ZN(n18398) );
  OAI211_X1 U21506 ( .C1(n18559), .C2(n18400), .A(n18399), .B(n18398), .ZN(
        P3_U2939) );
  NAND2_X1 U21507 ( .A1(n18454), .A2(n18401), .ZN(n18501) );
  AOI22_X1 U21508 ( .A1(n18562), .A2(n18420), .B1(n18561), .B2(n18417), .ZN(
        n18406) );
  INV_X1 U21509 ( .A(n18402), .ZN(n18404) );
  AOI22_X1 U21510 ( .A1(n18566), .A2(n18404), .B1(n18454), .B2(n18403), .ZN(
        n18421) );
  AOI22_X1 U21511 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18421), .B1(
        n18567), .B2(n18444), .ZN(n18405) );
  OAI211_X1 U21512 ( .C1(n18501), .C2(n18570), .A(n18406), .B(n18405), .ZN(
        P3_U2940) );
  AOI22_X1 U21513 ( .A1(n18444), .A2(n18573), .B1(n18571), .B2(n18420), .ZN(
        n18408) );
  INV_X1 U21514 ( .A(n18501), .ZN(n18494) );
  AOI22_X1 U21515 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18421), .B1(
        n18494), .B2(n18506), .ZN(n18407) );
  OAI211_X1 U21516 ( .C1(n18509), .C2(n18424), .A(n18408), .B(n18407), .ZN(
        P3_U2941) );
  AOI22_X1 U21517 ( .A1(n18444), .A2(n18536), .B1(n18578), .B2(n18420), .ZN(
        n18410) );
  AOI22_X1 U21518 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18421), .B1(
        n18577), .B2(n18417), .ZN(n18409) );
  OAI211_X1 U21519 ( .C1(n18501), .C2(n18539), .A(n18410), .B(n18409), .ZN(
        P3_U2942) );
  AOI22_X1 U21520 ( .A1(n18444), .A2(n18585), .B1(n18583), .B2(n18420), .ZN(
        n18412) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18421), .B1(
        n18494), .B2(n18436), .ZN(n18411) );
  OAI211_X1 U21522 ( .C1(n18439), .C2(n18424), .A(n18412), .B(n18411), .ZN(
        P3_U2943) );
  AOI22_X1 U21523 ( .A1(n18444), .A2(n18590), .B1(n18591), .B2(n18420), .ZN(
        n18414) );
  AOI22_X1 U21524 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18421), .B1(
        n18494), .B2(n18592), .ZN(n18413) );
  OAI211_X1 U21525 ( .C1(n18595), .C2(n18424), .A(n18414), .B(n18413), .ZN(
        P3_U2944) );
  AOI22_X1 U21526 ( .A1(n18444), .A2(n18597), .B1(n18598), .B2(n18420), .ZN(
        n18416) );
  AOI22_X1 U21527 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18421), .B1(
        n18494), .B2(n18599), .ZN(n18415) );
  OAI211_X1 U21528 ( .C1(n18603), .C2(n18424), .A(n18416), .B(n18415), .ZN(
        P3_U2945) );
  AOI22_X1 U21529 ( .A1(n18605), .A2(n18417), .B1(n18604), .B2(n18420), .ZN(
        n18419) );
  AOI22_X1 U21530 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18421), .B1(
        n18494), .B2(n18606), .ZN(n18418) );
  OAI211_X1 U21531 ( .C1(n18451), .C2(n18609), .A(n18419), .B(n18418), .ZN(
        P3_U2946) );
  AOI22_X1 U21532 ( .A1(n18444), .A2(n18552), .B1(n18611), .B2(n18420), .ZN(
        n18423) );
  AOI22_X1 U21533 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18421), .B1(
        n18494), .B2(n18615), .ZN(n18422) );
  OAI211_X1 U21534 ( .C1(n18559), .C2(n18424), .A(n18423), .B(n18422), .ZN(
        P3_U2947) );
  NOR2_X2 U21535 ( .A1(n18452), .A2(n18425), .ZN(n18522) );
  AOI221_X1 U21536 ( .B1(n18501), .B2(n18528), .C1(n18501), .C2(n18426), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18427) );
  OAI21_X1 U21537 ( .B1(n18522), .B2(n18427), .A(n18530), .ZN(n18448) );
  INV_X1 U21538 ( .A(n18448), .ZN(n18431) );
  AOI22_X1 U21539 ( .A1(n18444), .A2(n18561), .B1(n18562), .B2(n18447), .ZN(
        n18430) );
  AOI22_X1 U21540 ( .A1(n18567), .A2(n18473), .B1(n18522), .B2(n18428), .ZN(
        n18429) );
  OAI211_X1 U21541 ( .C1(n18431), .C2(n21014), .A(n18430), .B(n18429), .ZN(
        P3_U2948) );
  AOI22_X1 U21542 ( .A1(n18473), .A2(n18573), .B1(n18447), .B2(n18571), .ZN(
        n18433) );
  AOI22_X1 U21543 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18448), .B1(
        n18522), .B2(n18506), .ZN(n18432) );
  OAI211_X1 U21544 ( .C1(n18451), .C2(n18509), .A(n18433), .B(n18432), .ZN(
        P3_U2949) );
  AOI22_X1 U21545 ( .A1(n18444), .A2(n18577), .B1(n18447), .B2(n18578), .ZN(
        n18435) );
  AOI22_X1 U21546 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18448), .B1(
        n18522), .B2(n18579), .ZN(n18434) );
  OAI211_X1 U21547 ( .C1(n18471), .C2(n18582), .A(n18435), .B(n18434), .ZN(
        P3_U2950) );
  AOI22_X1 U21548 ( .A1(n18473), .A2(n18585), .B1(n18447), .B2(n18583), .ZN(
        n18438) );
  AOI22_X1 U21549 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18448), .B1(
        n18522), .B2(n18436), .ZN(n18437) );
  OAI211_X1 U21550 ( .C1(n18451), .C2(n18439), .A(n18438), .B(n18437), .ZN(
        P3_U2951) );
  AOI22_X1 U21551 ( .A1(n18473), .A2(n18590), .B1(n18447), .B2(n18591), .ZN(
        n18441) );
  AOI22_X1 U21552 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18448), .B1(
        n18522), .B2(n18592), .ZN(n18440) );
  OAI211_X1 U21553 ( .C1(n18451), .C2(n18595), .A(n18441), .B(n18440), .ZN(
        P3_U2952) );
  AOI22_X1 U21554 ( .A1(n18473), .A2(n18597), .B1(n18447), .B2(n18598), .ZN(
        n18443) );
  AOI22_X1 U21555 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18448), .B1(
        n18522), .B2(n18599), .ZN(n18442) );
  OAI211_X1 U21556 ( .C1(n18451), .C2(n18603), .A(n18443), .B(n18442), .ZN(
        P3_U2953) );
  AOI22_X1 U21557 ( .A1(n18444), .A2(n18605), .B1(n18447), .B2(n18604), .ZN(
        n18446) );
  AOI22_X1 U21558 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18448), .B1(
        n18522), .B2(n18606), .ZN(n18445) );
  OAI211_X1 U21559 ( .C1(n18471), .C2(n18609), .A(n18446), .B(n18445), .ZN(
        P3_U2954) );
  AOI22_X1 U21560 ( .A1(n18473), .A2(n18552), .B1(n18447), .B2(n18611), .ZN(
        n18450) );
  AOI22_X1 U21561 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18448), .B1(
        n18522), .B2(n18615), .ZN(n18449) );
  OAI211_X1 U21562 ( .C1(n18451), .C2(n18559), .A(n18450), .B(n18449), .ZN(
        P3_U2955) );
  NOR2_X1 U21563 ( .A1(n18646), .A2(n18452), .ZN(n18503) );
  NAND2_X1 U21564 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18503), .ZN(
        n18558) );
  INV_X1 U21565 ( .A(n18503), .ZN(n18453) );
  NOR2_X1 U21566 ( .A1(n9722), .A2(n18453), .ZN(n18472) );
  AOI22_X1 U21567 ( .A1(n18473), .A2(n18561), .B1(n18562), .B2(n18472), .ZN(
        n18456) );
  AOI22_X1 U21568 ( .A1(n18566), .A2(n18454), .B1(n18503), .B2(n18563), .ZN(
        n18474) );
  AOI22_X1 U21569 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18474), .B1(
        n18567), .B2(n18494), .ZN(n18455) );
  OAI211_X1 U21570 ( .C1(n18570), .C2(n18558), .A(n18456), .B(n18455), .ZN(
        P3_U2956) );
  AOI22_X1 U21571 ( .A1(n18494), .A2(n18573), .B1(n18571), .B2(n18472), .ZN(
        n18458) );
  AOI22_X1 U21572 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18474), .B1(
        n18506), .B2(n18540), .ZN(n18457) );
  OAI211_X1 U21573 ( .C1(n18471), .C2(n18509), .A(n18458), .B(n18457), .ZN(
        P3_U2957) );
  AOI22_X1 U21574 ( .A1(n18494), .A2(n18536), .B1(n18578), .B2(n18472), .ZN(
        n18460) );
  AOI22_X1 U21575 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18474), .B1(
        n18473), .B2(n18577), .ZN(n18459) );
  OAI211_X1 U21576 ( .C1(n18539), .C2(n18558), .A(n18460), .B(n18459), .ZN(
        P3_U2958) );
  AOI22_X1 U21577 ( .A1(n18473), .A2(n18584), .B1(n18583), .B2(n18472), .ZN(
        n18462) );
  AOI22_X1 U21578 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18474), .B1(
        n18494), .B2(n18585), .ZN(n18461) );
  OAI211_X1 U21579 ( .C1(n18589), .C2(n18558), .A(n18462), .B(n18461), .ZN(
        P3_U2959) );
  AOI22_X1 U21580 ( .A1(n18473), .A2(n18488), .B1(n18591), .B2(n18472), .ZN(
        n18464) );
  AOI22_X1 U21581 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18474), .B1(
        n18592), .B2(n18540), .ZN(n18463) );
  OAI211_X1 U21582 ( .C1(n18501), .C2(n18491), .A(n18464), .B(n18463), .ZN(
        P3_U2960) );
  AOI22_X1 U21583 ( .A1(n18473), .A2(n18465), .B1(n18598), .B2(n18472), .ZN(
        n18467) );
  AOI22_X1 U21584 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18474), .B1(
        n18599), .B2(n18540), .ZN(n18466) );
  OAI211_X1 U21585 ( .C1(n18501), .C2(n18468), .A(n18467), .B(n18466), .ZN(
        P3_U2961) );
  AOI22_X1 U21586 ( .A1(n18494), .A2(n18548), .B1(n18604), .B2(n18472), .ZN(
        n18470) );
  AOI22_X1 U21587 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18474), .B1(
        n18606), .B2(n18540), .ZN(n18469) );
  OAI211_X1 U21588 ( .C1(n18471), .C2(n18551), .A(n18470), .B(n18469), .ZN(
        P3_U2962) );
  AOI22_X1 U21589 ( .A1(n18473), .A2(n18613), .B1(n18611), .B2(n18472), .ZN(
        n18476) );
  AOI22_X1 U21590 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18474), .B1(
        n18615), .B2(n18540), .ZN(n18475) );
  OAI211_X1 U21591 ( .C1(n18501), .C2(n18620), .A(n18476), .B(n18475), .ZN(
        P3_U2963) );
  NAND2_X1 U21592 ( .A1(n18477), .A2(n18565), .ZN(n18602) );
  INV_X1 U21593 ( .A(n18602), .ZN(n18612) );
  NOR2_X1 U21594 ( .A1(n18540), .A2(n18612), .ZN(n18529) );
  NOR2_X1 U21595 ( .A1(n9722), .A2(n18529), .ZN(n18497) );
  AOI22_X1 U21596 ( .A1(n18567), .A2(n18522), .B1(n18562), .B2(n18497), .ZN(
        n18481) );
  OAI21_X1 U21597 ( .B1(n18527), .B2(n18478), .A(n18529), .ZN(n18479) );
  OAI211_X1 U21598 ( .C1(n18612), .C2(n18787), .A(n18530), .B(n18479), .ZN(
        n18498) );
  AOI22_X1 U21599 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18498), .B1(
        n18494), .B2(n18561), .ZN(n18480) );
  OAI211_X1 U21600 ( .C1(n18570), .C2(n18602), .A(n18481), .B(n18480), .ZN(
        P3_U2964) );
  AOI22_X1 U21601 ( .A1(n18522), .A2(n18573), .B1(n18571), .B2(n18497), .ZN(
        n18483) );
  AOI22_X1 U21602 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18498), .B1(
        n18506), .B2(n18612), .ZN(n18482) );
  OAI211_X1 U21603 ( .C1(n18501), .C2(n18509), .A(n18483), .B(n18482), .ZN(
        P3_U2965) );
  AOI22_X1 U21604 ( .A1(n18522), .A2(n18536), .B1(n18578), .B2(n18497), .ZN(
        n18485) );
  AOI22_X1 U21605 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18498), .B1(
        n18494), .B2(n18577), .ZN(n18484) );
  OAI211_X1 U21606 ( .C1(n18539), .C2(n18602), .A(n18485), .B(n18484), .ZN(
        P3_U2966) );
  AOI22_X1 U21607 ( .A1(n18494), .A2(n18584), .B1(n18583), .B2(n18497), .ZN(
        n18487) );
  AOI22_X1 U21608 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18498), .B1(
        n18522), .B2(n18585), .ZN(n18486) );
  OAI211_X1 U21609 ( .C1(n18589), .C2(n18602), .A(n18487), .B(n18486), .ZN(
        P3_U2967) );
  INV_X1 U21610 ( .A(n18522), .ZN(n18520) );
  AOI22_X1 U21611 ( .A1(n18494), .A2(n18488), .B1(n18591), .B2(n18497), .ZN(
        n18490) );
  AOI22_X1 U21612 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18498), .B1(
        n18592), .B2(n18612), .ZN(n18489) );
  OAI211_X1 U21613 ( .C1(n18520), .C2(n18491), .A(n18490), .B(n18489), .ZN(
        P3_U2968) );
  AOI22_X1 U21614 ( .A1(n18522), .A2(n18597), .B1(n18598), .B2(n18497), .ZN(
        n18493) );
  AOI22_X1 U21615 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18498), .B1(
        n18599), .B2(n18612), .ZN(n18492) );
  OAI211_X1 U21616 ( .C1(n18501), .C2(n18603), .A(n18493), .B(n18492), .ZN(
        P3_U2969) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18498), .B1(
        n18604), .B2(n18497), .ZN(n18496) );
  AOI22_X1 U21618 ( .A1(n18494), .A2(n18605), .B1(n18606), .B2(n18612), .ZN(
        n18495) );
  OAI211_X1 U21619 ( .C1(n18520), .C2(n18609), .A(n18496), .B(n18495), .ZN(
        P3_U2970) );
  AOI22_X1 U21620 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18498), .B1(
        n18611), .B2(n18497), .ZN(n18500) );
  AOI22_X1 U21621 ( .A1(n18522), .A2(n18552), .B1(n18615), .B2(n18612), .ZN(
        n18499) );
  OAI211_X1 U21622 ( .C1(n18501), .C2(n18559), .A(n18500), .B(n18499), .ZN(
        P3_U2971) );
  NOR2_X1 U21623 ( .A1(n9722), .A2(n18502), .ZN(n18521) );
  AOI22_X1 U21624 ( .A1(n18522), .A2(n18561), .B1(n18562), .B2(n18521), .ZN(
        n18505) );
  AOI22_X1 U21625 ( .A1(n18566), .A2(n18503), .B1(n18565), .B2(n18563), .ZN(
        n18523) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18523), .B1(
        n18567), .B2(n18540), .ZN(n18504) );
  OAI211_X1 U21627 ( .C1(n18570), .C2(n18619), .A(n18505), .B(n18504), .ZN(
        P3_U2972) );
  AOI22_X1 U21628 ( .A1(n18571), .A2(n18521), .B1(n18573), .B2(n18540), .ZN(
        n18508) );
  AOI22_X1 U21629 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18523), .B1(
        n18506), .B2(n18596), .ZN(n18507) );
  OAI211_X1 U21630 ( .C1(n18520), .C2(n18509), .A(n18508), .B(n18507), .ZN(
        P3_U2973) );
  AOI22_X1 U21631 ( .A1(n18536), .A2(n18540), .B1(n18578), .B2(n18521), .ZN(
        n18511) );
  AOI22_X1 U21632 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18523), .B1(
        n18522), .B2(n18577), .ZN(n18510) );
  OAI211_X1 U21633 ( .C1(n18539), .C2(n18619), .A(n18511), .B(n18510), .ZN(
        P3_U2974) );
  AOI22_X1 U21634 ( .A1(n18522), .A2(n18584), .B1(n18583), .B2(n18521), .ZN(
        n18513) );
  AOI22_X1 U21635 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18523), .B1(
        n18585), .B2(n18540), .ZN(n18512) );
  OAI211_X1 U21636 ( .C1(n18589), .C2(n18619), .A(n18513), .B(n18512), .ZN(
        P3_U2975) );
  AOI22_X1 U21637 ( .A1(n18591), .A2(n18521), .B1(n18590), .B2(n18540), .ZN(
        n18515) );
  AOI22_X1 U21638 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18523), .B1(
        n18592), .B2(n18596), .ZN(n18514) );
  OAI211_X1 U21639 ( .C1(n18520), .C2(n18595), .A(n18515), .B(n18514), .ZN(
        P3_U2976) );
  AOI22_X1 U21640 ( .A1(n18598), .A2(n18521), .B1(n18597), .B2(n18540), .ZN(
        n18517) );
  AOI22_X1 U21641 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18523), .B1(
        n18599), .B2(n18596), .ZN(n18516) );
  OAI211_X1 U21642 ( .C1(n18520), .C2(n18603), .A(n18517), .B(n18516), .ZN(
        P3_U2977) );
  AOI22_X1 U21643 ( .A1(n18548), .A2(n18540), .B1(n18604), .B2(n18521), .ZN(
        n18519) );
  AOI22_X1 U21644 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18523), .B1(
        n18606), .B2(n18596), .ZN(n18518) );
  OAI211_X1 U21645 ( .C1(n18520), .C2(n18551), .A(n18519), .B(n18518), .ZN(
        P3_U2978) );
  AOI22_X1 U21646 ( .A1(n18522), .A2(n18613), .B1(n18611), .B2(n18521), .ZN(
        n18525) );
  AOI22_X1 U21647 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18523), .B1(
        n18615), .B2(n18596), .ZN(n18524) );
  OAI211_X1 U21648 ( .C1(n18620), .C2(n18558), .A(n18525), .B(n18524), .ZN(
        P3_U2979) );
  AOI22_X1 U21649 ( .A1(n18567), .A2(n18612), .B1(n18562), .B2(n18553), .ZN(
        n18533) );
  AOI221_X1 U21650 ( .B1(n18529), .B2(n18619), .C1(n18528), .C2(n18619), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18531) );
  OAI21_X1 U21651 ( .B1(n18554), .B2(n18531), .A(n18530), .ZN(n18555) );
  AOI22_X1 U21652 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18555), .B1(
        n18561), .B2(n18540), .ZN(n18532) );
  OAI211_X1 U21653 ( .C1(n18570), .C2(n18543), .A(n18533), .B(n18532), .ZN(
        P3_U2980) );
  AOI22_X1 U21654 ( .A1(n18572), .A2(n18540), .B1(n18571), .B2(n18553), .ZN(
        n18535) );
  AOI22_X1 U21655 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18555), .B1(
        n18573), .B2(n18612), .ZN(n18534) );
  OAI211_X1 U21656 ( .C1(n18576), .C2(n18543), .A(n18535), .B(n18534), .ZN(
        P3_U2981) );
  AOI22_X1 U21657 ( .A1(n18536), .A2(n18612), .B1(n18578), .B2(n18553), .ZN(
        n18538) );
  AOI22_X1 U21658 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18555), .B1(
        n18577), .B2(n18540), .ZN(n18537) );
  OAI211_X1 U21659 ( .C1(n18539), .C2(n18543), .A(n18538), .B(n18537), .ZN(
        P3_U2982) );
  AOI22_X1 U21660 ( .A1(n18584), .A2(n18540), .B1(n18583), .B2(n18553), .ZN(
        n18542) );
  AOI22_X1 U21661 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18555), .B1(
        n18585), .B2(n18612), .ZN(n18541) );
  OAI211_X1 U21662 ( .C1(n18589), .C2(n18543), .A(n18542), .B(n18541), .ZN(
        P3_U2983) );
  AOI22_X1 U21663 ( .A1(n18591), .A2(n18553), .B1(n18590), .B2(n18612), .ZN(
        n18545) );
  AOI22_X1 U21664 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18555), .B1(
        n18592), .B2(n18554), .ZN(n18544) );
  OAI211_X1 U21665 ( .C1(n18595), .C2(n18558), .A(n18545), .B(n18544), .ZN(
        P3_U2984) );
  AOI22_X1 U21666 ( .A1(n18598), .A2(n18553), .B1(n18597), .B2(n18612), .ZN(
        n18547) );
  AOI22_X1 U21667 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18555), .B1(
        n18599), .B2(n18554), .ZN(n18546) );
  OAI211_X1 U21668 ( .C1(n18603), .C2(n18558), .A(n18547), .B(n18546), .ZN(
        P3_U2985) );
  AOI22_X1 U21669 ( .A1(n18548), .A2(n18612), .B1(n18604), .B2(n18553), .ZN(
        n18550) );
  AOI22_X1 U21670 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18555), .B1(
        n18606), .B2(n18554), .ZN(n18549) );
  OAI211_X1 U21671 ( .C1(n18551), .C2(n18558), .A(n18550), .B(n18549), .ZN(
        P3_U2986) );
  AOI22_X1 U21672 ( .A1(n18611), .A2(n18553), .B1(n18552), .B2(n18612), .ZN(
        n18557) );
  AOI22_X1 U21673 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18555), .B1(
        n18615), .B2(n18554), .ZN(n18556) );
  OAI211_X1 U21674 ( .C1(n18559), .C2(n18558), .A(n18557), .B(n18556), .ZN(
        P3_U2987) );
  INV_X1 U21675 ( .A(n18564), .ZN(n18560) );
  NOR2_X1 U21676 ( .A1(n9722), .A2(n18560), .ZN(n18610) );
  AOI22_X1 U21677 ( .A1(n18562), .A2(n18610), .B1(n18561), .B2(n18612), .ZN(
        n18569) );
  AOI22_X1 U21678 ( .A1(n18566), .A2(n18565), .B1(n18564), .B2(n18563), .ZN(
        n18616) );
  AOI22_X1 U21679 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18616), .B1(
        n18567), .B2(n18596), .ZN(n18568) );
  OAI211_X1 U21680 ( .C1(n18570), .C2(n18588), .A(n18569), .B(n18568), .ZN(
        P3_U2988) );
  AOI22_X1 U21681 ( .A1(n18572), .A2(n18612), .B1(n18571), .B2(n18610), .ZN(
        n18575) );
  AOI22_X1 U21682 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18616), .B1(
        n18573), .B2(n18596), .ZN(n18574) );
  OAI211_X1 U21683 ( .C1(n18576), .C2(n18588), .A(n18575), .B(n18574), .ZN(
        P3_U2989) );
  AOI22_X1 U21684 ( .A1(n18578), .A2(n18610), .B1(n18577), .B2(n18612), .ZN(
        n18581) );
  AOI22_X1 U21685 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18616), .B1(
        n18579), .B2(n18614), .ZN(n18580) );
  OAI211_X1 U21686 ( .C1(n18582), .C2(n18619), .A(n18581), .B(n18580), .ZN(
        P3_U2990) );
  AOI22_X1 U21687 ( .A1(n18584), .A2(n18612), .B1(n18583), .B2(n18610), .ZN(
        n18587) );
  AOI22_X1 U21688 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18616), .B1(
        n18585), .B2(n18596), .ZN(n18586) );
  OAI211_X1 U21689 ( .C1(n18589), .C2(n18588), .A(n18587), .B(n18586), .ZN(
        P3_U2991) );
  AOI22_X1 U21690 ( .A1(n18591), .A2(n18610), .B1(n18590), .B2(n18596), .ZN(
        n18594) );
  AOI22_X1 U21691 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18616), .B1(
        n18592), .B2(n18614), .ZN(n18593) );
  OAI211_X1 U21692 ( .C1(n18595), .C2(n18602), .A(n18594), .B(n18593), .ZN(
        P3_U2992) );
  AOI22_X1 U21693 ( .A1(n18598), .A2(n18610), .B1(n18597), .B2(n18596), .ZN(
        n18601) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18616), .B1(
        n18599), .B2(n18614), .ZN(n18600) );
  OAI211_X1 U21695 ( .C1(n18603), .C2(n18602), .A(n18601), .B(n18600), .ZN(
        P3_U2993) );
  AOI22_X1 U21696 ( .A1(n18605), .A2(n18612), .B1(n18604), .B2(n18610), .ZN(
        n18608) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18616), .B1(
        n18606), .B2(n18614), .ZN(n18607) );
  OAI211_X1 U21698 ( .C1(n18609), .C2(n18619), .A(n18608), .B(n18607), .ZN(
        P3_U2994) );
  AOI22_X1 U21699 ( .A1(n18613), .A2(n18612), .B1(n18611), .B2(n18610), .ZN(
        n18618) );
  AOI22_X1 U21700 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18616), .B1(
        n18615), .B2(n18614), .ZN(n18617) );
  OAI211_X1 U21701 ( .C1(n18620), .C2(n18619), .A(n18618), .B(n18617), .ZN(
        P3_U2995) );
  INV_X1 U21702 ( .A(n18621), .ZN(n18624) );
  AOI21_X1 U21703 ( .B1(n18624), .B2(n18623), .A(n18622), .ZN(n18633) );
  OAI21_X1 U21704 ( .B1(n18635), .B2(n18643), .A(n18633), .ZN(n18625) );
  AOI21_X1 U21705 ( .B1(n18626), .B2(n18625), .A(n18629), .ZN(n18627) );
  INV_X1 U21706 ( .A(n18627), .ZN(n18792) );
  NOR2_X1 U21707 ( .A1(n18668), .A2(n18792), .ZN(n18632) );
  AOI21_X1 U21708 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18641), .A(
        n18628), .ZN(n18644) );
  INV_X1 U21709 ( .A(n18635), .ZN(n18630) );
  OAI22_X1 U21710 ( .A1(n18644), .A2(n18630), .B1(n18629), .B2(n18659), .ZN(
        n18789) );
  NAND2_X1 U21711 ( .A1(n18793), .A2(n18789), .ZN(n18631) );
  OAI22_X1 U21712 ( .A1(n18632), .A2(n18793), .B1(n18668), .B2(n18631), .ZN(
        n18676) );
  NOR3_X1 U21713 ( .A1(n18634), .A2(n18633), .A3(n18803), .ZN(n18637) );
  AOI211_X1 U21714 ( .C1(n18803), .C2(n18811), .A(n18644), .B(n18635), .ZN(
        n18636) );
  AOI211_X1 U21715 ( .C1(n18639), .C2(n18638), .A(n18637), .B(n18636), .ZN(
        n18799) );
  AOI22_X1 U21716 ( .A1(n18668), .A2(n18803), .B1(n18799), .B2(n18640), .ZN(
        n18663) );
  NOR2_X1 U21717 ( .A1(n18642), .A2(n18641), .ZN(n18645) );
  AOI22_X1 U21718 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18643), .B1(
        n18645), .B2(n18818), .ZN(n18649) );
  OAI22_X1 U21719 ( .A1(n18645), .A2(n18804), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18644), .ZN(n18809) );
  AOI21_X1 U21720 ( .B1(n18649), .B2(n18646), .A(n18809), .ZN(n18648) );
  OAI21_X1 U21721 ( .B1(n18668), .B2(n18648), .A(n18647), .ZN(n18651) );
  INV_X1 U21722 ( .A(n18649), .ZN(n18812) );
  NAND3_X1 U21723 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n18812), .ZN(n18650) );
  OAI211_X1 U21724 ( .C1(n21113), .C2(n18663), .A(n18651), .B(n18650), .ZN(
        n18661) );
  INV_X1 U21725 ( .A(n18663), .ZN(n18652) );
  OAI221_X1 U21726 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n18661), .A(n18652), .ZN(
        n18675) );
  AOI22_X1 U21727 ( .A1(n18656), .A2(n18655), .B1(n18654), .B2(n18653), .ZN(
        n18657) );
  OAI221_X1 U21728 ( .B1(n18660), .B2(n18659), .C1(n18660), .C2(n18658), .A(
        n18657), .ZN(n18828) );
  INV_X1 U21729 ( .A(n18661), .ZN(n18662) );
  AOI21_X1 U21730 ( .B1(n21113), .B2(n18663), .A(n18662), .ZN(n18673) );
  NAND2_X1 U21731 ( .A1(n18665), .A2(n18664), .ZN(n18672) );
  AOI211_X1 U21732 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18668), .A(
        n18667), .B(n18666), .ZN(n18671) );
  OAI21_X1 U21733 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18669), .ZN(n18670) );
  OAI211_X1 U21734 ( .C1(n18673), .C2(n18672), .A(n18671), .B(n18670), .ZN(
        n18674) );
  AOI211_X1 U21735 ( .C1(n18676), .C2(n18675), .A(n18828), .B(n18674), .ZN(
        n18686) );
  NAND2_X1 U21736 ( .A1(n20974), .A2(n18687), .ZN(n18696) );
  INV_X1 U21737 ( .A(n18696), .ZN(n18838) );
  AOI22_X1 U21738 ( .A1(n18815), .A2(n18838), .B1(n18707), .B2(n18832), .ZN(
        n18677) );
  INV_X1 U21739 ( .A(n18677), .ZN(n18682) );
  OAI211_X1 U21740 ( .C1(n18679), .C2(n18678), .A(n18830), .B(n18686), .ZN(
        n18786) );
  OAI21_X1 U21741 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18836), .A(n18786), 
        .ZN(n18688) );
  NOR2_X1 U21742 ( .A1(n18680), .A2(n18688), .ZN(n18681) );
  MUX2_X1 U21743 ( .A(n18682), .B(n18681), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18684) );
  OAI211_X1 U21744 ( .C1(n18686), .C2(n18685), .A(n18684), .B(n18683), .ZN(
        P3_U2996) );
  NAND2_X1 U21745 ( .A1(n18707), .A2(n18832), .ZN(n18692) );
  NAND4_X1 U21746 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n18707), .A4(n18687), .ZN(n18694) );
  OR3_X1 U21747 ( .A1(n9722), .A2(n18689), .A3(n18688), .ZN(n18691) );
  NAND4_X1 U21748 ( .A1(n18693), .A2(n18692), .A3(n18694), .A4(n18691), .ZN(
        P3_U2997) );
  AND4_X1 U21749 ( .A1(n18696), .A2(n18695), .A3(n18694), .A4(n18785), .ZN(
        P3_U2998) );
  AND2_X1 U21750 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18697), .ZN(
        P3_U2999) );
  AND2_X1 U21751 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18697), .ZN(
        P3_U3000) );
  AND2_X1 U21752 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18697), .ZN(
        P3_U3001) );
  AND2_X1 U21753 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18697), .ZN(
        P3_U3002) );
  AND2_X1 U21754 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18697), .ZN(
        P3_U3003) );
  AND2_X1 U21755 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18697), .ZN(
        P3_U3004) );
  AND2_X1 U21756 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18697), .ZN(
        P3_U3005) );
  AND2_X1 U21757 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18697), .ZN(
        P3_U3006) );
  AND2_X1 U21758 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18697), .ZN(
        P3_U3007) );
  AND2_X1 U21759 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18697), .ZN(
        P3_U3008) );
  AND2_X1 U21760 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18697), .ZN(
        P3_U3009) );
  AND2_X1 U21761 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18697), .ZN(
        P3_U3010) );
  AND2_X1 U21762 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18697), .ZN(
        P3_U3011) );
  AND2_X1 U21763 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18697), .ZN(
        P3_U3012) );
  AND2_X1 U21764 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18697), .ZN(
        P3_U3013) );
  AND2_X1 U21765 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18697), .ZN(
        P3_U3014) );
  AND2_X1 U21766 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18697), .ZN(
        P3_U3015) );
  AND2_X1 U21767 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18697), .ZN(
        P3_U3016) );
  AND2_X1 U21768 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18697), .ZN(
        P3_U3017) );
  AND2_X1 U21769 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18697), .ZN(
        P3_U3018) );
  AND2_X1 U21770 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18697), .ZN(
        P3_U3019) );
  AND2_X1 U21771 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18697), .ZN(
        P3_U3020) );
  AND2_X1 U21772 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18697), .ZN(P3_U3021) );
  AND2_X1 U21773 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18697), .ZN(P3_U3022) );
  INV_X1 U21774 ( .A(P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n21045) );
  NOR2_X1 U21775 ( .A1(n21045), .A2(n18784), .ZN(P3_U3023) );
  AND2_X1 U21776 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18697), .ZN(P3_U3024) );
  AND2_X1 U21777 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18697), .ZN(P3_U3025) );
  AND2_X1 U21778 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18697), .ZN(P3_U3026) );
  AND2_X1 U21779 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18697), .ZN(P3_U3027) );
  AND2_X1 U21780 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18697), .ZN(P3_U3028) );
  OAI21_X1 U21781 ( .B1(n18698), .B2(n20778), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18699) );
  AOI22_X1 U21782 ( .A1(n18712), .A2(n18714), .B1(n18843), .B2(n18699), .ZN(
        n18701) );
  NAND3_X1 U21783 ( .A1(NA), .A2(n18712), .A3(n18700), .ZN(n18706) );
  OAI211_X1 U21784 ( .C1(n18836), .C2(n18702), .A(n18701), .B(n18706), .ZN(
        P3_U3029) );
  NOR2_X1 U21785 ( .A1(n18714), .A2(n20778), .ZN(n18710) );
  INV_X1 U21786 ( .A(n18710), .ZN(n18704) );
  INV_X1 U21787 ( .A(n18702), .ZN(n18703) );
  AOI22_X1 U21788 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(n18704), .B1(HOLD), 
        .B2(n18703), .ZN(n18705) );
  NAND2_X1 U21789 ( .A1(n18707), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18708) );
  OAI211_X1 U21790 ( .C1(n18705), .C2(n18712), .A(n18708), .B(n18833), .ZN(
        P3_U3030) );
  AOI22_X1 U21791 ( .A1(n18707), .A2(P3_STATE_REG_1__SCAN_IN), .B1(n18712), 
        .B2(n18706), .ZN(n18713) );
  OAI22_X1 U21792 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18708), .ZN(n18709) );
  OAI22_X1 U21793 ( .A1(n18710), .A2(n18709), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18711) );
  OAI22_X1 U21794 ( .A1(n18713), .A2(n18714), .B1(n18712), .B2(n18711), .ZN(
        P3_U3031) );
  INV_X2 U21795 ( .A(n18719), .ZN(n18769) );
  OAI222_X1 U21796 ( .A1(n18716), .A2(n18769), .B1(n18715), .B2(n18773), .C1(
        n18717), .C2(n18760), .ZN(P3_U3032) );
  OAI222_X1 U21797 ( .A1(n18760), .A2(n20931), .B1(n18718), .B2(n18773), .C1(
        n18717), .C2(n18769), .ZN(P3_U3033) );
  OAI222_X1 U21798 ( .A1(n18760), .A2(n20983), .B1(n18720), .B2(n18773), .C1(
        n20931), .C2(n18769), .ZN(P3_U3034) );
  OAI222_X1 U21799 ( .A1(n18760), .A2(n18722), .B1(n18721), .B2(n18773), .C1(
        n20983), .C2(n18769), .ZN(P3_U3035) );
  INV_X1 U21800 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18724) );
  OAI222_X1 U21801 ( .A1(n18760), .A2(n18724), .B1(n18723), .B2(n18773), .C1(
        n18722), .C2(n18769), .ZN(P3_U3036) );
  OAI222_X1 U21802 ( .A1(n18760), .A2(n18726), .B1(n18725), .B2(n18773), .C1(
        n18724), .C2(n18769), .ZN(P3_U3037) );
  INV_X1 U21803 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18729) );
  OAI222_X1 U21804 ( .A1(n18760), .A2(n18729), .B1(n18727), .B2(n18779), .C1(
        n18726), .C2(n18769), .ZN(P3_U3038) );
  OAI222_X1 U21805 ( .A1(n18729), .A2(n18769), .B1(n18728), .B2(n18773), .C1(
        n18730), .C2(n18760), .ZN(P3_U3039) );
  OAI222_X1 U21806 ( .A1(n18760), .A2(n18732), .B1(n18731), .B2(n18773), .C1(
        n18730), .C2(n18769), .ZN(P3_U3040) );
  OAI222_X1 U21807 ( .A1(n18760), .A2(n18734), .B1(n18733), .B2(n18779), .C1(
        n18732), .C2(n18769), .ZN(P3_U3041) );
  OAI222_X1 U21808 ( .A1(n18760), .A2(n18736), .B1(n18735), .B2(n18779), .C1(
        n18734), .C2(n18769), .ZN(P3_U3042) );
  OAI222_X1 U21809 ( .A1(n18760), .A2(n18738), .B1(n18737), .B2(n18779), .C1(
        n18736), .C2(n18769), .ZN(P3_U3043) );
  OAI222_X1 U21810 ( .A1(n18760), .A2(n20962), .B1(n18739), .B2(n18779), .C1(
        n18738), .C2(n18769), .ZN(P3_U3044) );
  OAI222_X1 U21811 ( .A1(n18760), .A2(n21154), .B1(n18740), .B2(n18779), .C1(
        n20962), .C2(n18769), .ZN(P3_U3045) );
  OAI222_X1 U21812 ( .A1(n18760), .A2(n18742), .B1(n18741), .B2(n18779), .C1(
        n21154), .C2(n18769), .ZN(P3_U3046) );
  OAI222_X1 U21813 ( .A1(n18760), .A2(n18744), .B1(n18743), .B2(n18779), .C1(
        n18742), .C2(n18769), .ZN(P3_U3047) );
  OAI222_X1 U21814 ( .A1(n18760), .A2(n18746), .B1(n18745), .B2(n18779), .C1(
        n18744), .C2(n18769), .ZN(P3_U3048) );
  OAI222_X1 U21815 ( .A1(n18760), .A2(n18748), .B1(n18747), .B2(n18779), .C1(
        n18746), .C2(n18769), .ZN(P3_U3049) );
  OAI222_X1 U21816 ( .A1(n18760), .A2(n18750), .B1(n18749), .B2(n18779), .C1(
        n18748), .C2(n18769), .ZN(P3_U3050) );
  OAI222_X1 U21817 ( .A1(n18760), .A2(n18752), .B1(n18751), .B2(n18779), .C1(
        n18750), .C2(n18769), .ZN(P3_U3051) );
  INV_X1 U21818 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18754) );
  OAI222_X1 U21819 ( .A1(n18760), .A2(n18754), .B1(n18753), .B2(n18779), .C1(
        n18752), .C2(n18769), .ZN(P3_U3052) );
  OAI222_X1 U21820 ( .A1(n18760), .A2(n18756), .B1(n18755), .B2(n18779), .C1(
        n18754), .C2(n18769), .ZN(P3_U3053) );
  OAI222_X1 U21821 ( .A1(n18760), .A2(n18758), .B1(n18757), .B2(n18773), .C1(
        n18756), .C2(n18769), .ZN(P3_U3054) );
  OAI222_X1 U21822 ( .A1(n18760), .A2(n18761), .B1(n18759), .B2(n18773), .C1(
        n18758), .C2(n18769), .ZN(P3_U3055) );
  INV_X1 U21823 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18763) );
  OAI222_X1 U21824 ( .A1(n18760), .A2(n18763), .B1(n18762), .B2(n18773), .C1(
        n18761), .C2(n18769), .ZN(P3_U3056) );
  OAI222_X1 U21825 ( .A1(n18760), .A2(n18765), .B1(n18764), .B2(n18773), .C1(
        n18763), .C2(n18769), .ZN(P3_U3057) );
  OAI222_X1 U21826 ( .A1(n18760), .A2(n18768), .B1(n18766), .B2(n18773), .C1(
        n18765), .C2(n18769), .ZN(P3_U3058) );
  OAI222_X1 U21827 ( .A1(n18768), .A2(n18769), .B1(n18767), .B2(n18773), .C1(
        n18770), .C2(n18760), .ZN(P3_U3059) );
  OAI222_X1 U21828 ( .A1(n18760), .A2(n18775), .B1(n18771), .B2(n18773), .C1(
        n18770), .C2(n18769), .ZN(P3_U3060) );
  OAI222_X1 U21829 ( .A1(n18769), .A2(n18775), .B1(n18774), .B2(n18773), .C1(
        n18772), .C2(n18760), .ZN(P3_U3061) );
  OAI22_X1 U21830 ( .A1(n18843), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18779), .ZN(n18776) );
  INV_X1 U21831 ( .A(n18776), .ZN(P3_U3274) );
  OAI22_X1 U21832 ( .A1(n18843), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18773), .ZN(n18777) );
  INV_X1 U21833 ( .A(n18777), .ZN(P3_U3275) );
  OAI22_X1 U21834 ( .A1(n18843), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18773), .ZN(n18778) );
  INV_X1 U21835 ( .A(n18778), .ZN(P3_U3276) );
  OAI22_X1 U21836 ( .A1(n18843), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18779), .ZN(n18780) );
  INV_X1 U21837 ( .A(n18780), .ZN(P3_U3277) );
  OAI21_X1 U21838 ( .B1(n18784), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18782), 
        .ZN(n18781) );
  INV_X1 U21839 ( .A(n18781), .ZN(P3_U3280) );
  OAI21_X1 U21840 ( .B1(n18784), .B2(n18783), .A(n18782), .ZN(P3_U3281) );
  OAI221_X1 U21841 ( .B1(n18787), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18787), 
        .C2(n18786), .A(n18785), .ZN(P3_U3282) );
  INV_X1 U21842 ( .A(n18788), .ZN(n18791) );
  NOR2_X1 U21843 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18845), .ZN(
        n18790) );
  AOI22_X1 U21844 ( .A1(n18815), .A2(n18791), .B1(n18790), .B2(n18789), .ZN(
        n18795) );
  AOI21_X1 U21845 ( .B1(n18808), .B2(n18792), .A(n18819), .ZN(n18794) );
  OAI22_X1 U21846 ( .A1(n18819), .A2(n18795), .B1(n18794), .B2(n18793), .ZN(
        P3_U3285) );
  NOR2_X1 U21847 ( .A1(n20974), .A2(n18796), .ZN(n18805) );
  INV_X1 U21848 ( .A(n18805), .ZN(n18814) );
  AOI22_X1 U21849 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n18798), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18797), .ZN(n18806) );
  OAI22_X1 U21850 ( .A1(n18799), .A2(n18845), .B1(n18814), .B2(n18806), .ZN(
        n18800) );
  AOI21_X1 U21851 ( .B1(n18815), .B2(n18801), .A(n18800), .ZN(n18802) );
  AOI22_X1 U21852 ( .A1(n18819), .A2(n18803), .B1(n18802), .B2(n18816), .ZN(
        P3_U3288) );
  INV_X1 U21853 ( .A(n18804), .ZN(n18807) );
  AOI222_X1 U21854 ( .A1(n18809), .A2(n18808), .B1(n18815), .B2(n18807), .C1(
        n18806), .C2(n18805), .ZN(n18810) );
  AOI22_X1 U21855 ( .A1(n18819), .A2(n18811), .B1(n18810), .B2(n18816), .ZN(
        P3_U3289) );
  OAI21_X1 U21856 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18812), .A(n20974), 
        .ZN(n18813) );
  AOI22_X1 U21857 ( .A1(n18815), .A2(n18818), .B1(n18814), .B2(n18813), .ZN(
        n18817) );
  AOI22_X1 U21858 ( .A1(n18819), .A2(n18818), .B1(n18817), .B2(n18816), .ZN(
        P3_U3290) );
  AOI211_X1 U21859 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_REIP_REG_1__SCAN_IN), .B(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18820) );
  AOI21_X1 U21860 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18820), .ZN(n18822) );
  INV_X1 U21861 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18821) );
  AOI22_X1 U21862 ( .A1(n18826), .A2(n18822), .B1(n18821), .B2(n18823), .ZN(
        P3_U3292) );
  NOR2_X1 U21863 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n18825) );
  INV_X1 U21864 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18824) );
  AOI22_X1 U21865 ( .A1(n18826), .A2(n18825), .B1(n18824), .B2(n18823), .ZN(
        P3_U3293) );
  INV_X1 U21866 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n21072) );
  AOI22_X1 U21867 ( .A1(n18779), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n21072), 
        .B2(n18843), .ZN(P3_U3294) );
  MUX2_X1 U21868 ( .A(P3_MORE_REG_SCAN_IN), .B(n18828), .S(n18827), .Z(
        P3_U3295) );
  OAI21_X1 U21869 ( .B1(n18830), .B2(n18829), .A(n18846), .ZN(n18831) );
  AOI21_X1 U21870 ( .B1(n18832), .B2(n18836), .A(n18831), .ZN(n18842) );
  AOI21_X1 U21871 ( .B1(n18835), .B2(n18834), .A(n18833), .ZN(n18837) );
  OAI211_X1 U21872 ( .C1(n18837), .C2(n18847), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18836), .ZN(n18839) );
  AOI21_X1 U21873 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18839), .A(n18838), 
        .ZN(n18841) );
  NAND2_X1 U21874 ( .A1(n18842), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18840) );
  OAI21_X1 U21875 ( .B1(n18842), .B2(n18841), .A(n18840), .ZN(P3_U3296) );
  OAI22_X1 U21876 ( .A1(n18843), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18773), .ZN(n18844) );
  INV_X1 U21877 ( .A(n18844), .ZN(P3_U3297) );
  OAI21_X1 U21878 ( .B1(n18845), .B2(P3_STATE2_REG_2__SCAN_IN), .A(n18846), 
        .ZN(n18850) );
  OAI22_X1 U21879 ( .A1(n18847), .A2(n18846), .B1(n18850), .B2(
        P3_READREQUEST_REG_SCAN_IN), .ZN(n18848) );
  INV_X1 U21880 ( .A(n18848), .ZN(P3_U3298) );
  OAI21_X1 U21881 ( .B1(n18850), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n18849), 
        .ZN(n18851) );
  INV_X1 U21882 ( .A(n18851), .ZN(P3_U3299) );
  NAND2_X1 U21883 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19842), .ZN(n19831) );
  AOI22_X1 U21884 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19831), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n18855), .ZN(n19896) );
  AOI21_X1 U21885 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19896), .ZN(n18852) );
  INV_X1 U21886 ( .A(n18852), .ZN(P2_U2815) );
  AOI22_X1 U21887 ( .A1(n18853), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n19817), 
        .B2(n19818), .ZN(n18854) );
  INV_X1 U21888 ( .A(n18854), .ZN(P2_U2816) );
  NAND2_X1 U21889 ( .A1(n18855), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19945) );
  INV_X2 U21890 ( .A(n19945), .ZN(n19944) );
  AOI21_X1 U21891 ( .B1(n18855), .B2(n19842), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18856) );
  AOI22_X1 U21892 ( .A1(n19944), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18856), 
        .B2(n19945), .ZN(P2_U2817) );
  OAI21_X1 U21893 ( .B1(n19824), .B2(BS16), .A(n19896), .ZN(n19894) );
  OAI21_X1 U21894 ( .B1(n19896), .B2(n19898), .A(n19894), .ZN(P2_U2818) );
  NOR4_X1 U21895 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18860) );
  NOR4_X1 U21896 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18859) );
  NOR4_X1 U21897 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18858) );
  NOR4_X1 U21898 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18857) );
  NAND4_X1 U21899 ( .A1(n18860), .A2(n18859), .A3(n18858), .A4(n18857), .ZN(
        n18866) );
  NOR4_X1 U21900 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18864) );
  AOI211_X1 U21901 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_12__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18863) );
  NOR4_X1 U21902 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n18862) );
  NOR4_X1 U21903 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18861) );
  NAND4_X1 U21904 ( .A1(n18864), .A2(n18863), .A3(n18862), .A4(n18861), .ZN(
        n18865) );
  NOR2_X1 U21905 ( .A1(n18866), .A2(n18865), .ZN(n18877) );
  INV_X1 U21906 ( .A(n18877), .ZN(n18875) );
  NOR2_X1 U21907 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18875), .ZN(n18869) );
  INV_X1 U21908 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18867) );
  AOI22_X1 U21909 ( .A1(n18869), .A2(n18870), .B1(n18875), .B2(n18867), .ZN(
        P2_U2820) );
  OR3_X1 U21910 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18874) );
  INV_X1 U21911 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18868) );
  AOI22_X1 U21912 ( .A1(n18869), .A2(n18874), .B1(n18875), .B2(n18868), .ZN(
        P2_U2821) );
  INV_X1 U21913 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19895) );
  NAND2_X1 U21914 ( .A1(n18869), .A2(n19895), .ZN(n18873) );
  OAI21_X1 U21915 ( .B1(n19843), .B2(n18870), .A(n18877), .ZN(n18871) );
  OAI21_X1 U21916 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18877), .A(n18871), 
        .ZN(n18872) );
  OAI221_X1 U21917 ( .B1(n18873), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18873), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18872), .ZN(P2_U2822) );
  INV_X1 U21918 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18876) );
  OAI221_X1 U21919 ( .B1(n18877), .B2(n18876), .C1(n18875), .C2(n18874), .A(
        n18873), .ZN(P2_U2823) );
  AOI22_X1 U21920 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18996), .B1(
        P2_REIP_REG_19__SCAN_IN), .B2(n19025), .ZN(n18878) );
  OAI21_X1 U21921 ( .B1(n18879), .B2(n19018), .A(n18878), .ZN(n18880) );
  AOI211_X1 U21922 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19026), .A(n19000), .B(
        n18880), .ZN(n18887) );
  AOI21_X1 U21923 ( .B1(n18882), .B2(n18881), .A(n19820), .ZN(n18885) );
  AOI22_X1 U21924 ( .A1(n18885), .A2(n18884), .B1(n18883), .B2(n19020), .ZN(
        n18886) );
  OAI211_X1 U21925 ( .C1(n18888), .C2(n19029), .A(n18887), .B(n18886), .ZN(
        P2_U2836) );
  NOR2_X1 U21926 ( .A1(n9753), .A2(n18889), .ZN(n18891) );
  XOR2_X1 U21927 ( .A(n18891), .B(n18890), .Z(n18900) );
  AOI22_X1 U21928 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18996), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19025), .ZN(n18892) );
  OAI21_X1 U21929 ( .B1(n18893), .B2(n19018), .A(n18892), .ZN(n18894) );
  AOI211_X1 U21930 ( .C1(P2_EBX_REG_18__SCAN_IN), .C2(n19026), .A(n19000), .B(
        n18894), .ZN(n18899) );
  NOR2_X1 U21931 ( .A1(n18895), .A2(n19029), .ZN(n18896) );
  AOI21_X1 U21932 ( .B1(n18897), .B2(n19020), .A(n18896), .ZN(n18898) );
  OAI211_X1 U21933 ( .C1(n19820), .C2(n18900), .A(n18899), .B(n18898), .ZN(
        P2_U2837) );
  OAI21_X1 U21934 ( .B1(n21170), .B2(n19010), .A(n18983), .ZN(n18903) );
  OAI22_X1 U21935 ( .A1(n18901), .A2(n19018), .B1(n19037), .B2(n9987), .ZN(
        n18902) );
  AOI211_X1 U21936 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n19026), .A(n18903), .B(
        n18902), .ZN(n18910) );
  NAND2_X1 U21937 ( .A1(n19002), .A2(n18904), .ZN(n18906) );
  XNOR2_X1 U21938 ( .A(n18906), .B(n18905), .ZN(n18908) );
  AOI22_X1 U21939 ( .A1(n18908), .A2(n19021), .B1(n19020), .B2(n18907), .ZN(
        n18909) );
  OAI211_X1 U21940 ( .C1(n18911), .C2(n19029), .A(n18910), .B(n18909), .ZN(
        P2_U2838) );
  NOR2_X1 U21941 ( .A1(n9753), .A2(n18912), .ZN(n18914) );
  XOR2_X1 U21942 ( .A(n18914), .B(n18913), .Z(n18922) );
  OAI21_X1 U21943 ( .B1(n15235), .B2(n19010), .A(n18983), .ZN(n18918) );
  INV_X1 U21944 ( .A(n18915), .ZN(n18916) );
  OAI22_X1 U21945 ( .A1(n18916), .A2(n19018), .B1(n19037), .B2(n9986), .ZN(
        n18917) );
  AOI211_X1 U21946 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n19026), .A(n18918), .B(
        n18917), .ZN(n18921) );
  AOI22_X1 U21947 ( .A1(n18919), .A2(n19020), .B1(n19015), .B2(n19054), .ZN(
        n18920) );
  OAI211_X1 U21948 ( .C1(n19820), .C2(n18922), .A(n18921), .B(n18920), .ZN(
        P2_U2839) );
  AOI211_X1 U21949 ( .C1(n18932), .C2(n18924), .A(n18923), .B(n19042), .ZN(
        n18930) );
  NAND2_X1 U21950 ( .A1(n18925), .A2(n19032), .ZN(n18928) );
  AOI22_X1 U21951 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n18996), .B1(
        P2_EBX_REG_13__SCAN_IN), .B2(n19026), .ZN(n18927) );
  NAND2_X1 U21952 ( .A1(n19025), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n18926) );
  NAND4_X1 U21953 ( .A1(n18928), .A2(n18927), .A3(n18983), .A4(n18926), .ZN(
        n18929) );
  NOR2_X1 U21954 ( .A1(n18930), .A2(n18929), .ZN(n18935) );
  AOI22_X1 U21955 ( .A1(n18933), .A2(n19020), .B1(n18932), .B2(n18931), .ZN(
        n18934) );
  OAI211_X1 U21956 ( .C1(n18936), .C2(n19029), .A(n18935), .B(n18934), .ZN(
        P2_U2842) );
  INV_X1 U21957 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18947) );
  OAI22_X1 U21958 ( .A1(n18937), .A2(n19018), .B1(n19861), .B2(n19010), .ZN(
        n18938) );
  AOI211_X1 U21959 ( .C1(P2_EBX_REG_12__SCAN_IN), .C2(n19026), .A(n19000), .B(
        n18938), .ZN(n18946) );
  XNOR2_X1 U21960 ( .A(n18940), .B(n18939), .ZN(n18944) );
  OAI22_X1 U21961 ( .A1(n18942), .A2(n19034), .B1(n19029), .B2(n18941), .ZN(
        n18943) );
  AOI21_X1 U21962 ( .B1(n18944), .B2(n19021), .A(n18943), .ZN(n18945) );
  OAI211_X1 U21963 ( .C1(n18947), .C2(n19037), .A(n18946), .B(n18945), .ZN(
        P2_U2843) );
  OAI21_X1 U21964 ( .B1(n19858), .B2(n19010), .A(n18983), .ZN(n18951) );
  OAI22_X1 U21965 ( .A1(n18949), .A2(n19018), .B1(n18948), .B2(n19012), .ZN(
        n18950) );
  AOI211_X1 U21966 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n18996), .A(
        n18951), .B(n18950), .ZN(n18958) );
  NOR2_X1 U21967 ( .A1(n9753), .A2(n18952), .ZN(n18954) );
  XNOR2_X1 U21968 ( .A(n18954), .B(n18953), .ZN(n18956) );
  AOI22_X1 U21969 ( .A1(n18956), .A2(n19021), .B1(n19020), .B2(n18955), .ZN(
        n18957) );
  OAI211_X1 U21970 ( .C1(n18959), .C2(n19029), .A(n18958), .B(n18957), .ZN(
        P2_U2845) );
  NAND2_X1 U21971 ( .A1(n19002), .A2(n18960), .ZN(n18962) );
  XOR2_X1 U21972 ( .A(n18962), .B(n18961), .Z(n18970) );
  AOI22_X1 U21973 ( .A1(n18963), .A2(n19032), .B1(P2_REIP_REG_9__SCAN_IN), 
        .B2(n19025), .ZN(n18964) );
  OAI211_X1 U21974 ( .C1(n10906), .C2(n19012), .A(n18964), .B(n18983), .ZN(
        n18968) );
  OAI22_X1 U21975 ( .A1(n18966), .A2(n19034), .B1(n19029), .B2(n18965), .ZN(
        n18967) );
  AOI211_X1 U21976 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n18996), .A(
        n18968), .B(n18967), .ZN(n18969) );
  OAI21_X1 U21977 ( .B1(n18970), .B2(n19820), .A(n18969), .ZN(P2_U2846) );
  NAND2_X1 U21978 ( .A1(n19002), .A2(n18971), .ZN(n18973) );
  XOR2_X1 U21979 ( .A(n18973), .B(n18972), .Z(n18982) );
  AOI22_X1 U21980 ( .A1(n18974), .A2(n19032), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n19026), .ZN(n18975) );
  OAI211_X1 U21981 ( .C1(n19853), .C2(n19010), .A(n18975), .B(n18983), .ZN(
        n18980) );
  INV_X1 U21982 ( .A(n18976), .ZN(n18978) );
  OAI22_X1 U21983 ( .A1(n19034), .A2(n18978), .B1(n18977), .B2(n19029), .ZN(
        n18979) );
  AOI211_X1 U21984 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n18996), .A(
        n18980), .B(n18979), .ZN(n18981) );
  OAI21_X1 U21985 ( .B1(n18982), .B2(n19820), .A(n18981), .ZN(P2_U2848) );
  INV_X1 U21986 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19851) );
  OAI21_X1 U21987 ( .B1(n19851), .B2(n19010), .A(n18983), .ZN(n18987) );
  OAI22_X1 U21988 ( .A1(n18985), .A2(n19018), .B1(n19012), .B2(n18984), .ZN(
        n18986) );
  AOI211_X1 U21989 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n18996), .A(
        n18987), .B(n18986), .ZN(n18994) );
  NOR2_X1 U21990 ( .A1(n9753), .A2(n18988), .ZN(n18990) );
  XNOR2_X1 U21991 ( .A(n18990), .B(n18989), .ZN(n18992) );
  AOI22_X1 U21992 ( .A1(n18992), .A2(n19021), .B1(n19020), .B2(n18991), .ZN(
        n18993) );
  OAI211_X1 U21993 ( .C1(n19029), .C2(n18995), .A(n18994), .B(n18993), .ZN(
        P2_U2849) );
  AOI22_X1 U21994 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n18996), .B1(
        P2_REIP_REG_5__SCAN_IN), .B2(n19025), .ZN(n18997) );
  OAI21_X1 U21995 ( .B1(n18998), .B2(n19018), .A(n18997), .ZN(n18999) );
  AOI211_X1 U21996 ( .C1(P2_EBX_REG_5__SCAN_IN), .C2(n19026), .A(n19000), .B(
        n18999), .ZN(n19008) );
  NAND2_X1 U21997 ( .A1(n19002), .A2(n19001), .ZN(n19003) );
  XNOR2_X1 U21998 ( .A(n19004), .B(n19003), .ZN(n19006) );
  AOI22_X1 U21999 ( .A1(n19006), .A2(n19021), .B1(n19020), .B2(n19005), .ZN(
        n19007) );
  OAI211_X1 U22000 ( .C1(n19029), .C2(n19069), .A(n19008), .B(n19007), .ZN(
        P2_U2850) );
  OAI22_X1 U22001 ( .A1(n19010), .A2(n19843), .B1(n19037), .B2(n19009), .ZN(
        n19014) );
  INV_X1 U22002 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n19011) );
  NOR2_X1 U22003 ( .A1(n19012), .A2(n19011), .ZN(n19013) );
  AOI211_X1 U22004 ( .C1(n19015), .C2(n19922), .A(n19014), .B(n19013), .ZN(
        n19016) );
  OAI21_X1 U22005 ( .B1(n19018), .B2(n19017), .A(n19016), .ZN(n19019) );
  AOI21_X1 U22006 ( .B1(n19198), .B2(n19020), .A(n19019), .ZN(n19024) );
  AOI22_X1 U22007 ( .A1(n19022), .A2(n19021), .B1(n19920), .B2(n19040), .ZN(
        n19023) );
  OAI211_X1 U22008 ( .C1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n19036), .A(
        n19024), .B(n19023), .ZN(P2_U2854) );
  AOI22_X1 U22009 ( .A1(n19026), .A2(P2_EBX_REG_0__SCAN_IN), .B1(
        P2_REIP_REG_0__SCAN_IN), .B2(n19025), .ZN(n19027) );
  OAI21_X1 U22010 ( .B1(n19029), .B2(n19028), .A(n19027), .ZN(n19030) );
  AOI21_X1 U22011 ( .B1(n19032), .B2(n19031), .A(n19030), .ZN(n19033) );
  OAI21_X1 U22012 ( .B1(n19035), .B2(n19034), .A(n19033), .ZN(n19039) );
  INV_X1 U22013 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19167) );
  AOI21_X1 U22014 ( .B1(n19037), .B2(n19036), .A(n19167), .ZN(n19038) );
  AOI211_X1 U22015 ( .C1(n19265), .C2(n19040), .A(n19039), .B(n19038), .ZN(
        n19041) );
  OAI21_X1 U22016 ( .B1(n19043), .B2(n19042), .A(n19041), .ZN(P2_U2855) );
  AOI22_X1 U22017 ( .A1(n19045), .A2(n19055), .B1(n19044), .B2(
        BUF1_REG_31__SCAN_IN), .ZN(n19048) );
  AOI22_X1 U22018 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19053), .B1(n19046), 
        .B2(BUF2_REG_31__SCAN_IN), .ZN(n19047) );
  NAND2_X1 U22019 ( .A1(n19048), .A2(n19047), .ZN(P2_U2888) );
  OAI22_X1 U22020 ( .A1(n19051), .A2(n19050), .B1(n19049), .B2(n19211), .ZN(
        n19052) );
  AOI21_X1 U22021 ( .B1(P2_EAX_REG_16__SCAN_IN), .B2(n19053), .A(n19052), .ZN(
        n19058) );
  AOI22_X1 U22022 ( .A1(n19056), .A2(n19064), .B1(n19055), .B2(n19054), .ZN(
        n19057) );
  OAI211_X1 U22023 ( .C1(n19059), .C2(n14275), .A(n19058), .B(n19057), .ZN(
        P2_U2903) );
  INV_X1 U22024 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19127) );
  OAI22_X1 U22025 ( .A1(n19061), .A2(n19237), .B1(n19060), .B2(n19127), .ZN(
        n19062) );
  INV_X1 U22026 ( .A(n19062), .ZN(n19068) );
  INV_X1 U22027 ( .A(n19063), .ZN(n19065) );
  NAND3_X1 U22028 ( .A1(n19066), .A2(n19065), .A3(n19064), .ZN(n19067) );
  OAI211_X1 U22029 ( .C1(n19070), .C2(n19069), .A(n19068), .B(n19067), .ZN(
        P2_U2914) );
  NAND3_X1 U22030 ( .A1(n19072), .A2(n19071), .A3(n19815), .ZN(n19074) );
  NAND2_X1 U22031 ( .A1(n19074), .A2(n19073), .ZN(n19075) );
  INV_X1 U22032 ( .A(n19076), .ZN(n19139) );
  NOR2_X1 U22033 ( .A1(n21034), .A2(n19133), .ZN(P2_U2920) );
  INV_X1 U22034 ( .A(n19077), .ZN(n19078) );
  AND2_X1 U22035 ( .A1(n19131), .A2(n19078), .ZN(n19081) );
  AOI22_X1 U22036 ( .A1(P2_EAX_REG_30__SCAN_IN), .A2(n19081), .B1(n19139), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19079) );
  OAI21_X1 U22037 ( .B1(n19133), .B2(n19080), .A(n19079), .ZN(P2_U2921) );
  INV_X2 U22038 ( .A(n19133), .ZN(n19136) );
  AOI22_X1 U22039 ( .A1(n19130), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19136), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n19082) );
  OAI21_X1 U22040 ( .B1(n19083), .B2(n19105), .A(n19082), .ZN(P2_U2922) );
  AOI22_X1 U22041 ( .A1(n19139), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19136), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n19084) );
  OAI21_X1 U22042 ( .B1(n14821), .B2(n19105), .A(n19084), .ZN(P2_U2923) );
  AOI22_X1 U22043 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n19136), .B1(n19130), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n19085) );
  OAI21_X1 U22044 ( .B1(n19086), .B2(n19105), .A(n19085), .ZN(P2_U2924) );
  AOI22_X1 U22045 ( .A1(n19139), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19136), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n19087) );
  OAI21_X1 U22046 ( .B1(n20996), .B2(n19105), .A(n19087), .ZN(P2_U2925) );
  AOI22_X1 U22047 ( .A1(n19139), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19136), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n19088) );
  OAI21_X1 U22048 ( .B1(n19089), .B2(n19105), .A(n19088), .ZN(P2_U2926) );
  AOI22_X1 U22049 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n19136), .B1(n19130), 
        .B2(P2_UWORD_REG_8__SCAN_IN), .ZN(n19090) );
  OAI21_X1 U22050 ( .B1(n14855), .B2(n19105), .A(n19090), .ZN(P2_U2927) );
  AOI22_X1 U22051 ( .A1(n19139), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19136), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n19091) );
  OAI21_X1 U22052 ( .B1(n19092), .B2(n19105), .A(n19091), .ZN(P2_U2928) );
  INV_X1 U22053 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n19094) );
  AOI22_X1 U22054 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n19136), .B1(n19130), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n19093) );
  OAI21_X1 U22055 ( .B1(n19094), .B2(n19105), .A(n19093), .ZN(P2_U2929) );
  INV_X1 U22056 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n19096) );
  AOI22_X1 U22057 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n19136), .B1(n19130), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n19095) );
  OAI21_X1 U22058 ( .B1(n19096), .B2(n19105), .A(n19095), .ZN(P2_U2930) );
  INV_X1 U22059 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n19098) );
  AOI22_X1 U22060 ( .A1(n19139), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19136), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n19097) );
  OAI21_X1 U22061 ( .B1(n19098), .B2(n19105), .A(n19097), .ZN(P2_U2931) );
  AOI22_X1 U22062 ( .A1(P2_UWORD_REG_3__SCAN_IN), .A2(n19130), .B1(n19136), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n19099) );
  OAI21_X1 U22063 ( .B1(n14874), .B2(n19105), .A(n19099), .ZN(P2_U2932) );
  INV_X1 U22064 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n19101) );
  AOI22_X1 U22065 ( .A1(n19139), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19136), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n19100) );
  OAI21_X1 U22066 ( .B1(n19101), .B2(n19105), .A(n19100), .ZN(P2_U2933) );
  AOI22_X1 U22067 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n19136), .B1(n19130), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n19102) );
  OAI21_X1 U22068 ( .B1(n19103), .B2(n19105), .A(n19102), .ZN(P2_U2934) );
  INV_X1 U22069 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n19106) );
  AOI22_X1 U22070 ( .A1(n19139), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19136), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n19104) );
  OAI21_X1 U22071 ( .B1(n19106), .B2(n19105), .A(n19104), .ZN(P2_U2935) );
  AOI22_X1 U22072 ( .A1(n19139), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19136), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19107) );
  OAI21_X1 U22073 ( .B1(n19108), .B2(n19141), .A(n19107), .ZN(P2_U2936) );
  AOI22_X1 U22074 ( .A1(n19139), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19136), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19109) );
  OAI21_X1 U22075 ( .B1(n19110), .B2(n19141), .A(n19109), .ZN(P2_U2937) );
  AOI22_X1 U22076 ( .A1(P2_LWORD_REG_13__SCAN_IN), .A2(n19130), .B1(n19136), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19111) );
  OAI21_X1 U22077 ( .B1(n19112), .B2(n19141), .A(n19111), .ZN(P2_U2938) );
  AOI22_X1 U22078 ( .A1(n19139), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19136), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19113) );
  OAI21_X1 U22079 ( .B1(n19114), .B2(n19141), .A(n19113), .ZN(P2_U2939) );
  AOI22_X1 U22080 ( .A1(n19139), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19136), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19115) );
  OAI21_X1 U22081 ( .B1(n19116), .B2(n19141), .A(n19115), .ZN(P2_U2940) );
  AOI22_X1 U22082 ( .A1(n19139), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19136), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19117) );
  OAI21_X1 U22083 ( .B1(n21013), .B2(n19141), .A(n19117), .ZN(P2_U2941) );
  AOI22_X1 U22084 ( .A1(n19139), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19136), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19118) );
  OAI21_X1 U22085 ( .B1(n19119), .B2(n19141), .A(n19118), .ZN(P2_U2942) );
  AOI22_X1 U22086 ( .A1(n19139), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19136), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19120) );
  OAI21_X1 U22087 ( .B1(n19121), .B2(n19141), .A(n19120), .ZN(P2_U2943) );
  AOI22_X1 U22088 ( .A1(n19139), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19136), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19122) );
  OAI21_X1 U22089 ( .B1(n19123), .B2(n19141), .A(n19122), .ZN(P2_U2944) );
  AOI22_X1 U22090 ( .A1(n19139), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19136), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19124) );
  OAI21_X1 U22091 ( .B1(n19125), .B2(n19141), .A(n19124), .ZN(P2_U2945) );
  AOI22_X1 U22092 ( .A1(n19139), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19136), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19126) );
  OAI21_X1 U22093 ( .B1(n19127), .B2(n19141), .A(n19126), .ZN(P2_U2946) );
  INV_X1 U22094 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19129) );
  AOI22_X1 U22095 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n19136), .B1(n19130), 
        .B2(P2_LWORD_REG_4__SCAN_IN), .ZN(n19128) );
  OAI21_X1 U22096 ( .B1(n19129), .B2(n19141), .A(n19128), .ZN(P2_U2947) );
  AOI22_X1 U22097 ( .A1(P2_EAX_REG_3__SCAN_IN), .A2(n19131), .B1(n19130), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n19132) );
  OAI21_X1 U22098 ( .B1(n21089), .B2(n19133), .A(n19132), .ZN(P2_U2948) );
  INV_X1 U22099 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19135) );
  AOI22_X1 U22100 ( .A1(n19139), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19136), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19134) );
  OAI21_X1 U22101 ( .B1(n19135), .B2(n19141), .A(n19134), .ZN(P2_U2949) );
  AOI22_X1 U22102 ( .A1(n19139), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19136), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19137) );
  OAI21_X1 U22103 ( .B1(n19138), .B2(n19141), .A(n19137), .ZN(P2_U2950) );
  INV_X1 U22104 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19142) );
  AOI22_X1 U22105 ( .A1(n19139), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19136), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19140) );
  OAI21_X1 U22106 ( .B1(n19142), .B2(n19141), .A(n19140), .ZN(P2_U2951) );
  AOI22_X1 U22107 ( .A1(n19154), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19000), .ZN(n19150) );
  NAND2_X1 U22108 ( .A1(n19143), .A2(n19162), .ZN(n19146) );
  NAND2_X1 U22109 ( .A1(n19144), .A2(n19156), .ZN(n19145) );
  OAI211_X1 U22110 ( .C1(n19147), .C2(n19159), .A(n19146), .B(n19145), .ZN(
        n19148) );
  INV_X1 U22111 ( .A(n19148), .ZN(n19149) );
  OAI211_X1 U22112 ( .C1(n19152), .C2(n19151), .A(n19150), .B(n19149), .ZN(
        P2_U3010) );
  NOR2_X1 U22113 ( .A1(n19154), .A2(n19153), .ZN(n19168) );
  NAND2_X1 U22114 ( .A1(n19156), .A2(n19155), .ZN(n19165) );
  OAI21_X1 U22115 ( .B1(n19159), .B2(n19158), .A(n19157), .ZN(n19160) );
  INV_X1 U22116 ( .A(n19160), .ZN(n19164) );
  NAND2_X1 U22117 ( .A1(n19162), .A2(n19161), .ZN(n19163) );
  AND3_X1 U22118 ( .A1(n19165), .A2(n19164), .A3(n19163), .ZN(n19166) );
  OAI21_X1 U22119 ( .B1(n19168), .B2(n19167), .A(n19166), .ZN(P2_U3014) );
  NAND2_X1 U22120 ( .A1(n19199), .A2(n19169), .ZN(n19171) );
  OAI211_X1 U22121 ( .C1(n19172), .C2(n19175), .A(n19171), .B(n19170), .ZN(
        n19173) );
  AOI21_X1 U22122 ( .B1(n19913), .B2(n19187), .A(n19173), .ZN(n19184) );
  NOR2_X1 U22123 ( .A1(n19175), .A2(n19174), .ZN(n19180) );
  OAI22_X1 U22124 ( .A1(n19202), .A2(n19178), .B1(n19177), .B2(n19176), .ZN(
        n19179) );
  AOI211_X1 U22125 ( .C1(n19182), .C2(n19181), .A(n19180), .B(n19179), .ZN(
        n19183) );
  OAI211_X1 U22126 ( .C1(n19186), .C2(n19185), .A(n19184), .B(n19183), .ZN(
        P2_U3044) );
  AOI22_X1 U22127 ( .A1(n19188), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19187), .B2(n19922), .ZN(n19189) );
  OAI21_X1 U22128 ( .B1(n19191), .B2(n19190), .A(n19189), .ZN(n19197) );
  AOI211_X1 U22129 ( .C1(n19195), .C2(n19194), .A(n19193), .B(n19192), .ZN(
        n19196) );
  AOI211_X1 U22130 ( .C1(n19199), .C2(n19198), .A(n19197), .B(n19196), .ZN(
        n19201) );
  OAI211_X1 U22131 ( .C1(n19203), .C2(n19202), .A(n19201), .B(n19200), .ZN(
        P2_U3045) );
  NOR2_X1 U22132 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19318) );
  NAND2_X1 U22133 ( .A1(n19924), .A2(n19318), .ZN(n19264) );
  NOR2_X1 U22134 ( .A1(n19264), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19251) );
  INV_X1 U22135 ( .A(n19251), .ZN(n19208) );
  AND2_X1 U22136 ( .A1(n19804), .A2(n19208), .ZN(n19210) );
  OAI21_X1 U22137 ( .B1(n10590), .B2(n19251), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19209) );
  OAI21_X1 U22138 ( .B1(n19210), .B2(n19679), .A(n19209), .ZN(n19252) );
  NOR2_X2 U22139 ( .A1(n19211), .A2(n19682), .ZN(n19694) );
  NAND2_X1 U22140 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19753), .ZN(n19233) );
  AND2_X1 U22141 ( .A1(n19212), .A2(n19249), .ZN(n19687) );
  AOI22_X1 U22142 ( .A1(n19252), .A2(n19694), .B1(n19687), .B2(n19251), .ZN(
        n19218) );
  INV_X1 U22143 ( .A(n10590), .ZN(n19215) );
  NOR2_X2 U22144 ( .A1(n19506), .A2(n19413), .ZN(n19286) );
  INV_X1 U22145 ( .A(n19804), .ZN(n19213) );
  AOI221_X1 U22146 ( .B1(n19809), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19286), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19213), .ZN(n19214) );
  AOI211_X1 U22147 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19215), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19214), .ZN(n19216) );
  OAI21_X1 U22148 ( .B1(n19216), .B2(n19251), .A(n19753), .ZN(n19256) );
  AOI22_X1 U22149 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19247), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19246), .ZN(n19648) );
  AOI22_X1 U22150 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19256), .B1(
        n19286), .B2(n19755), .ZN(n19217) );
  OAI211_X1 U22151 ( .C1(n19758), .C2(n19801), .A(n19218), .B(n19217), .ZN(
        P2_U3048) );
  AOI22_X2 U22152 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19247), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19246), .ZN(n19765) );
  NOR2_X2 U22153 ( .A1(n19219), .A2(n19682), .ZN(n19699) );
  NAND2_X1 U22154 ( .A1(n9740), .A2(n19249), .ZN(n19759) );
  AOI22_X1 U22155 ( .A1(n19252), .A2(n19699), .B1(n19609), .B2(n19251), .ZN(
        n19221) );
  AOI22_X1 U22156 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19247), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19246), .ZN(n19653) );
  AOI22_X1 U22157 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19256), .B1(
        n19286), .B2(n19762), .ZN(n19220) );
  OAI211_X1 U22158 ( .C1(n19765), .C2(n19801), .A(n19221), .B(n19220), .ZN(
        P2_U3049) );
  AOI22_X1 U22159 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19247), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19246), .ZN(n19709) );
  NOR2_X2 U22160 ( .A1(n19222), .A2(n19682), .ZN(n19706) );
  AOI22_X1 U22161 ( .A1(n19252), .A2(n19706), .B1(n19703), .B2(n19251), .ZN(
        n19225) );
  AOI22_X1 U22162 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19247), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19246), .ZN(n19772) );
  AOI22_X1 U22163 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19256), .B1(
        n19286), .B2(n19704), .ZN(n19224) );
  OAI211_X1 U22164 ( .C1(n19709), .C2(n19801), .A(n19225), .B(n19224), .ZN(
        P2_U3050) );
  AOI22_X1 U22165 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19246), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19247), .ZN(n19710) );
  NOR2_X2 U22166 ( .A1(n19226), .A2(n19682), .ZN(n19712) );
  NAND2_X1 U22167 ( .A1(n19227), .A2(n19249), .ZN(n19773) );
  AOI22_X1 U22168 ( .A1(n19252), .A2(n19712), .B1(n19614), .B2(n19251), .ZN(
        n19229) );
  AOI22_X1 U22169 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19247), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19246), .ZN(n19779) );
  INV_X1 U22170 ( .A(n19779), .ZN(n19615) );
  AOI22_X1 U22171 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19256), .B1(
        n19286), .B2(n19615), .ZN(n19228) );
  OAI211_X1 U22172 ( .C1(n19710), .C2(n19801), .A(n19229), .B(n19228), .ZN(
        P2_U3051) );
  NOR2_X2 U22173 ( .A1(n19232), .A2(n19682), .ZN(n19717) );
  NOR2_X2 U22174 ( .A1(n19234), .A2(n19233), .ZN(n19715) );
  AOI22_X1 U22175 ( .A1(n19252), .A2(n19717), .B1(n19715), .B2(n19251), .ZN(
        n19236) );
  AOI22_X1 U22176 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19247), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19246), .ZN(n19720) );
  INV_X1 U22177 ( .A(n19720), .ZN(n19783) );
  AOI22_X1 U22178 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19256), .B1(
        n19286), .B2(n19783), .ZN(n19235) );
  OAI211_X1 U22179 ( .C1(n19786), .C2(n19801), .A(n19236), .B(n19235), .ZN(
        P2_U3052) );
  AOI22_X2 U22180 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19247), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19246), .ZN(n19793) );
  NOR2_X2 U22181 ( .A1(n19237), .A2(n19682), .ZN(n19723) );
  NAND2_X1 U22182 ( .A1(n10102), .A2(n19249), .ZN(n19787) );
  AOI22_X1 U22183 ( .A1(n19252), .A2(n19723), .B1(n19620), .B2(n19251), .ZN(
        n19239) );
  AOI22_X1 U22184 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19247), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19246), .ZN(n19726) );
  AOI22_X1 U22185 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19256), .B1(
        n19286), .B2(n19790), .ZN(n19238) );
  OAI211_X1 U22186 ( .C1(n19793), .C2(n19801), .A(n19239), .B(n19238), .ZN(
        P2_U3053) );
  NOR2_X2 U22187 ( .A1(n19242), .A2(n19682), .ZN(n19729) );
  AOI22_X1 U22188 ( .A1(n19252), .A2(n19729), .B1(n19727), .B2(n19251), .ZN(
        n19245) );
  AOI22_X1 U22189 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19247), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19246), .ZN(n19802) );
  INV_X1 U22190 ( .A(n19802), .ZN(n19623) );
  AOI22_X1 U22191 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19256), .B1(
        n19286), .B2(n19623), .ZN(n19244) );
  OAI211_X1 U22192 ( .C1(n19626), .C2(n19801), .A(n19245), .B(n19244), .ZN(
        P2_U3054) );
  AOI22_X2 U22193 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19247), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19246), .ZN(n19814) );
  NOR2_X2 U22194 ( .A1(n19248), .A2(n19682), .ZN(n19735) );
  AOI22_X1 U22195 ( .A1(n19252), .A2(n19735), .B1(n19733), .B2(n19251), .ZN(
        n19258) );
  OAI22_X2 U22196 ( .A1(n14241), .A2(n19255), .B1(n19254), .B2(n19253), .ZN(
        n19808) );
  AOI22_X1 U22197 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19256), .B1(
        n19286), .B2(n19808), .ZN(n19257) );
  OAI211_X1 U22198 ( .C1(n19814), .C2(n19801), .A(n19258), .B(n19257), .ZN(
        P2_U3055) );
  NAND2_X1 U22199 ( .A1(n19266), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19445) );
  OAI21_X1 U22200 ( .B1(n19445), .B2(n19506), .A(n19264), .ZN(n19262) );
  NAND2_X1 U22201 ( .A1(n10589), .A2(n19576), .ZN(n19260) );
  INV_X1 U22202 ( .A(n19318), .ZN(n19320) );
  NOR2_X1 U22203 ( .A1(n19505), .A2(n19320), .ZN(n19284) );
  NOR2_X1 U22204 ( .A1(n12882), .A2(n19284), .ZN(n19259) );
  AOI21_X1 U22205 ( .B1(n19260), .B2(n19259), .A(n19682), .ZN(n19261) );
  OAI21_X1 U22206 ( .B1(n10589), .B2(n19284), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19263) );
  OAI21_X1 U22207 ( .B1(n19264), .B2(n19679), .A(n19263), .ZN(n19285) );
  AOI22_X1 U22208 ( .A1(n19285), .A2(n19694), .B1(n19687), .B2(n19284), .ZN(
        n19268) );
  AOI22_X1 U22209 ( .A1(n19293), .A2(n19755), .B1(n19286), .B2(n19688), .ZN(
        n19267) );
  OAI211_X1 U22210 ( .C1(n19289), .C2(n19269), .A(n19268), .B(n19267), .ZN(
        P2_U3056) );
  AOI22_X1 U22211 ( .A1(n19285), .A2(n19699), .B1(n19609), .B2(n19284), .ZN(
        n19271) );
  INV_X1 U22212 ( .A(n19765), .ZN(n19650) );
  AOI22_X1 U22213 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19281), .B1(
        n19286), .B2(n19650), .ZN(n19270) );
  OAI211_X1 U22214 ( .C1(n19653), .C2(n19317), .A(n19271), .B(n19270), .ZN(
        P2_U3057) );
  AOI22_X1 U22215 ( .A1(n19285), .A2(n19706), .B1(n19703), .B2(n19284), .ZN(
        n19273) );
  INV_X1 U22216 ( .A(n19709), .ZN(n19769) );
  AOI22_X1 U22217 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19281), .B1(
        n19286), .B2(n19769), .ZN(n19272) );
  OAI211_X1 U22218 ( .C1(n19772), .C2(n19317), .A(n19273), .B(n19272), .ZN(
        P2_U3058) );
  INV_X1 U22219 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n19276) );
  AOI22_X1 U22220 ( .A1(n19285), .A2(n19712), .B1(n19614), .B2(n19284), .ZN(
        n19275) );
  INV_X1 U22221 ( .A(n19710), .ZN(n19776) );
  AOI22_X1 U22222 ( .A1(n19293), .A2(n19615), .B1(n19286), .B2(n19776), .ZN(
        n19274) );
  OAI211_X1 U22223 ( .C1(n19289), .C2(n19276), .A(n19275), .B(n19274), .ZN(
        P2_U3059) );
  AOI22_X1 U22224 ( .A1(n19285), .A2(n19717), .B1(n19715), .B2(n19284), .ZN(
        n19278) );
  AOI22_X1 U22225 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19281), .B1(
        n19286), .B2(n19716), .ZN(n19277) );
  OAI211_X1 U22226 ( .C1(n19720), .C2(n19317), .A(n19278), .B(n19277), .ZN(
        P2_U3060) );
  AOI22_X1 U22227 ( .A1(n19285), .A2(n19723), .B1(n19620), .B2(n19284), .ZN(
        n19280) );
  INV_X1 U22228 ( .A(n19793), .ZN(n19664) );
  AOI22_X1 U22229 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19281), .B1(
        n19286), .B2(n19664), .ZN(n19279) );
  OAI211_X1 U22230 ( .C1(n19726), .C2(n19317), .A(n19280), .B(n19279), .ZN(
        P2_U3061) );
  AOI22_X1 U22231 ( .A1(n19285), .A2(n19729), .B1(n19727), .B2(n19284), .ZN(
        n19283) );
  AOI22_X1 U22232 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19281), .B1(
        n19286), .B2(n19797), .ZN(n19282) );
  OAI211_X1 U22233 ( .C1(n19802), .C2(n19317), .A(n19283), .B(n19282), .ZN(
        P2_U3062) );
  INV_X1 U22234 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n20977) );
  AOI22_X1 U22235 ( .A1(n19285), .A2(n19735), .B1(n19733), .B2(n19284), .ZN(
        n19288) );
  INV_X1 U22236 ( .A(n19814), .ZN(n19348) );
  AOI22_X1 U22237 ( .A1(n19293), .A2(n19808), .B1(n19286), .B2(n19348), .ZN(
        n19287) );
  OAI211_X1 U22238 ( .C1(n19289), .C2(n20977), .A(n19288), .B(n19287), .ZN(
        P2_U3063) );
  NOR2_X1 U22239 ( .A1(n19538), .A2(n19320), .ZN(n19312) );
  OAI21_X1 U22240 ( .B1(n19291), .B2(n19312), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19290) );
  OR2_X1 U22241 ( .A1(n19320), .A2(n19540), .ZN(n19294) );
  NAND2_X1 U22242 ( .A1(n19290), .A2(n19294), .ZN(n19313) );
  AOI22_X1 U22243 ( .A1(n19313), .A2(n19694), .B1(n19687), .B2(n19312), .ZN(
        n19299) );
  INV_X1 U22244 ( .A(n19291), .ZN(n19292) );
  AOI21_X1 U22245 ( .B1(n19292), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19297) );
  NOR2_X2 U22246 ( .A1(n19413), .A2(n19572), .ZN(n19347) );
  OAI21_X1 U22247 ( .B1(n19293), .B2(n19347), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19295) );
  NAND3_X1 U22248 ( .A1(n19295), .A2(n12682), .A3(n19294), .ZN(n19296) );
  OAI211_X1 U22249 ( .C1(n19312), .C2(n19297), .A(n19296), .B(n19753), .ZN(
        n19314) );
  AOI22_X1 U22250 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19314), .B1(
        n19347), .B2(n19755), .ZN(n19298) );
  OAI211_X1 U22251 ( .C1(n19758), .C2(n19317), .A(n19299), .B(n19298), .ZN(
        P2_U3064) );
  AOI22_X1 U22252 ( .A1(n19313), .A2(n19699), .B1(n19609), .B2(n19312), .ZN(
        n19301) );
  AOI22_X1 U22253 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19314), .B1(
        n19347), .B2(n19762), .ZN(n19300) );
  OAI211_X1 U22254 ( .C1(n19765), .C2(n19317), .A(n19301), .B(n19300), .ZN(
        P2_U3065) );
  AOI22_X1 U22255 ( .A1(n19313), .A2(n19706), .B1(n19703), .B2(n19312), .ZN(
        n19303) );
  AOI22_X1 U22256 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19314), .B1(
        n19347), .B2(n19704), .ZN(n19302) );
  OAI211_X1 U22257 ( .C1(n19709), .C2(n19317), .A(n19303), .B(n19302), .ZN(
        P2_U3066) );
  AOI22_X1 U22258 ( .A1(n19313), .A2(n19712), .B1(n19614), .B2(n19312), .ZN(
        n19305) );
  AOI22_X1 U22259 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19314), .B1(
        n19347), .B2(n19615), .ZN(n19304) );
  OAI211_X1 U22260 ( .C1(n19710), .C2(n19317), .A(n19305), .B(n19304), .ZN(
        P2_U3067) );
  AOI22_X1 U22261 ( .A1(n19313), .A2(n19717), .B1(n19715), .B2(n19312), .ZN(
        n19307) );
  AOI22_X1 U22262 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19314), .B1(
        n19347), .B2(n19783), .ZN(n19306) );
  OAI211_X1 U22263 ( .C1(n19786), .C2(n19317), .A(n19307), .B(n19306), .ZN(
        P2_U3068) );
  AOI22_X1 U22264 ( .A1(n19313), .A2(n19723), .B1(n19620), .B2(n19312), .ZN(
        n19309) );
  AOI22_X1 U22265 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19314), .B1(
        n19347), .B2(n19790), .ZN(n19308) );
  OAI211_X1 U22266 ( .C1(n19793), .C2(n19317), .A(n19309), .B(n19308), .ZN(
        P2_U3069) );
  AOI22_X1 U22267 ( .A1(n19313), .A2(n19729), .B1(n19727), .B2(n19312), .ZN(
        n19311) );
  AOI22_X1 U22268 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19314), .B1(
        n19347), .B2(n19623), .ZN(n19310) );
  OAI211_X1 U22269 ( .C1(n19626), .C2(n19317), .A(n19311), .B(n19310), .ZN(
        P2_U3070) );
  AOI22_X1 U22270 ( .A1(n19313), .A2(n19735), .B1(n19733), .B2(n19312), .ZN(
        n19316) );
  AOI22_X1 U22271 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19314), .B1(
        n19347), .B2(n19808), .ZN(n19315) );
  OAI211_X1 U22272 ( .C1(n19814), .C2(n19317), .A(n19316), .B(n19315), .ZN(
        P2_U3071) );
  OAI21_X1 U22273 ( .B1(n19445), .B2(n19572), .A(n12682), .ZN(n19328) );
  NAND2_X1 U22274 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19318), .ZN(
        n19327) );
  INV_X1 U22275 ( .A(n19327), .ZN(n19319) );
  OR2_X1 U22276 ( .A1(n19328), .A2(n19319), .ZN(n19324) );
  NAND2_X1 U22277 ( .A1(n19325), .A2(n19576), .ZN(n19322) );
  NOR2_X1 U22278 ( .A1(n19320), .A2(n19566), .ZN(n19346) );
  NOR2_X1 U22279 ( .A1(n19346), .A2(n12682), .ZN(n19321) );
  AOI21_X1 U22280 ( .B1(n19322), .B2(n19321), .A(n19682), .ZN(n19323) );
  AOI22_X1 U22281 ( .A1(n19347), .A2(n19688), .B1(n19346), .B2(n19687), .ZN(
        n19330) );
  OAI21_X1 U22282 ( .B1(n19325), .B2(n19346), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19326) );
  OAI21_X1 U22283 ( .B1(n19328), .B2(n19327), .A(n19326), .ZN(n19349) );
  AOI22_X1 U22284 ( .A1(n19694), .A2(n19349), .B1(n19375), .B2(n19755), .ZN(
        n19329) );
  OAI211_X1 U22285 ( .C1(n19352), .C2(n19331), .A(n19330), .B(n19329), .ZN(
        P2_U3072) );
  AOI22_X1 U22286 ( .A1(n19375), .A2(n19762), .B1(n19346), .B2(n19609), .ZN(
        n19333) );
  AOI22_X1 U22287 ( .A1(n19699), .A2(n19349), .B1(n19347), .B2(n19650), .ZN(
        n19332) );
  OAI211_X1 U22288 ( .C1(n19352), .C2(n13684), .A(n19333), .B(n19332), .ZN(
        P2_U3073) );
  INV_X1 U22289 ( .A(n19347), .ZN(n19345) );
  AOI22_X1 U22290 ( .A1(n19704), .A2(n19375), .B1(n19346), .B2(n19703), .ZN(
        n19335) );
  INV_X1 U22291 ( .A(n19352), .ZN(n19342) );
  AOI22_X1 U22292 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19342), .B1(
        n19706), .B2(n19349), .ZN(n19334) );
  OAI211_X1 U22293 ( .C1(n19709), .C2(n19345), .A(n19335), .B(n19334), .ZN(
        P2_U3074) );
  AOI22_X1 U22294 ( .A1(n19375), .A2(n19615), .B1(n19346), .B2(n19614), .ZN(
        n19337) );
  AOI22_X1 U22295 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19342), .B1(
        n19712), .B2(n19349), .ZN(n19336) );
  OAI211_X1 U22296 ( .C1(n19710), .C2(n19345), .A(n19337), .B(n19336), .ZN(
        P2_U3075) );
  AOI22_X1 U22297 ( .A1(n19783), .A2(n19375), .B1(n19346), .B2(n19715), .ZN(
        n19339) );
  AOI22_X1 U22298 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19342), .B1(
        n19717), .B2(n19349), .ZN(n19338) );
  OAI211_X1 U22299 ( .C1(n19786), .C2(n19345), .A(n19339), .B(n19338), .ZN(
        P2_U3076) );
  AOI22_X1 U22300 ( .A1(n19347), .A2(n19664), .B1(n19346), .B2(n19620), .ZN(
        n19341) );
  AOI22_X1 U22301 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19342), .B1(
        n19723), .B2(n19349), .ZN(n19340) );
  OAI211_X1 U22302 ( .C1(n19726), .C2(n19383), .A(n19341), .B(n19340), .ZN(
        P2_U3077) );
  AOI22_X1 U22303 ( .A1(n19623), .A2(n19375), .B1(n19346), .B2(n19727), .ZN(
        n19344) );
  AOI22_X1 U22304 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19342), .B1(
        n19729), .B2(n19349), .ZN(n19343) );
  OAI211_X1 U22305 ( .C1(n19626), .C2(n19345), .A(n19344), .B(n19343), .ZN(
        P2_U3078) );
  INV_X1 U22306 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n21095) );
  AOI22_X1 U22307 ( .A1(n19348), .A2(n19347), .B1(n19346), .B2(n19733), .ZN(
        n19351) );
  AOI22_X1 U22308 ( .A1(n19735), .A2(n19349), .B1(n19375), .B2(n19808), .ZN(
        n19350) );
  OAI211_X1 U22309 ( .C1(n19352), .C2(n21095), .A(n19351), .B(n19350), .ZN(
        P2_U3079) );
  INV_X1 U22310 ( .A(n19414), .ZN(n19353) );
  NAND2_X1 U22311 ( .A1(n19354), .A2(n19353), .ZN(n19604) );
  NOR2_X1 U22312 ( .A1(n19604), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19362) );
  INV_X1 U22313 ( .A(n19362), .ZN(n19356) );
  NAND2_X1 U22314 ( .A1(n19908), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19440) );
  INV_X1 U22315 ( .A(n19440), .ZN(n19415) );
  NAND2_X1 U22316 ( .A1(n19415), .A2(n19924), .ZN(n19388) );
  NOR2_X1 U22317 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19388), .ZN(
        n19378) );
  OAI21_X1 U22318 ( .B1(n19357), .B2(n19378), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19355) );
  OAI21_X1 U22319 ( .B1(n19679), .B2(n19356), .A(n19355), .ZN(n19379) );
  AOI22_X1 U22320 ( .A1(n19379), .A2(n19694), .B1(n19687), .B2(n19378), .ZN(
        n19364) );
  AOI21_X1 U22321 ( .B1(n19383), .B2(n19410), .A(n19898), .ZN(n19361) );
  OAI21_X1 U22322 ( .B1(n19357), .B2(n19441), .A(n19576), .ZN(n19359) );
  INV_X1 U22323 ( .A(n19378), .ZN(n19358) );
  NAND2_X1 U22324 ( .A1(n19359), .A2(n19358), .ZN(n19360) );
  OAI211_X1 U22325 ( .C1(n19362), .C2(n19361), .A(n19360), .B(n19753), .ZN(
        n19380) );
  AOI22_X1 U22326 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19380), .B1(
        n19398), .B2(n19755), .ZN(n19363) );
  OAI211_X1 U22327 ( .C1(n19758), .C2(n19383), .A(n19364), .B(n19363), .ZN(
        P2_U3080) );
  AOI22_X1 U22328 ( .A1(n19379), .A2(n19699), .B1(n19609), .B2(n19378), .ZN(
        n19366) );
  AOI22_X1 U22329 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19380), .B1(
        n19398), .B2(n19762), .ZN(n19365) );
  OAI211_X1 U22330 ( .C1(n19765), .C2(n19383), .A(n19366), .B(n19365), .ZN(
        P2_U3081) );
  AOI22_X1 U22331 ( .A1(n19379), .A2(n19706), .B1(n19703), .B2(n19378), .ZN(
        n19368) );
  AOI22_X1 U22332 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19380), .B1(
        n19398), .B2(n19704), .ZN(n19367) );
  OAI211_X1 U22333 ( .C1(n19709), .C2(n19383), .A(n19368), .B(n19367), .ZN(
        P2_U3082) );
  AOI22_X1 U22334 ( .A1(n19379), .A2(n19712), .B1(n19614), .B2(n19378), .ZN(
        n19370) );
  AOI22_X1 U22335 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19380), .B1(
        n19375), .B2(n19776), .ZN(n19369) );
  OAI211_X1 U22336 ( .C1(n19779), .C2(n19410), .A(n19370), .B(n19369), .ZN(
        P2_U3083) );
  AOI22_X1 U22337 ( .A1(n19379), .A2(n19717), .B1(n19715), .B2(n19378), .ZN(
        n19372) );
  AOI22_X1 U22338 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19380), .B1(
        n19398), .B2(n19783), .ZN(n19371) );
  OAI211_X1 U22339 ( .C1(n19786), .C2(n19383), .A(n19372), .B(n19371), .ZN(
        P2_U3084) );
  AOI22_X1 U22340 ( .A1(n19379), .A2(n19723), .B1(n19620), .B2(n19378), .ZN(
        n19374) );
  AOI22_X1 U22341 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19380), .B1(
        n19398), .B2(n19790), .ZN(n19373) );
  OAI211_X1 U22342 ( .C1(n19793), .C2(n19383), .A(n19374), .B(n19373), .ZN(
        P2_U3085) );
  AOI22_X1 U22343 ( .A1(n19379), .A2(n19729), .B1(n19727), .B2(n19378), .ZN(
        n19377) );
  AOI22_X1 U22344 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19380), .B1(
        n19375), .B2(n19797), .ZN(n19376) );
  OAI211_X1 U22345 ( .C1(n19802), .C2(n19410), .A(n19377), .B(n19376), .ZN(
        P2_U3086) );
  AOI22_X1 U22346 ( .A1(n19379), .A2(n19735), .B1(n19733), .B2(n19378), .ZN(
        n19382) );
  AOI22_X1 U22347 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19380), .B1(
        n19398), .B2(n19808), .ZN(n19381) );
  OAI211_X1 U22348 ( .C1(n19814), .C2(n19383), .A(n19382), .B(n19381), .ZN(
        P2_U3087) );
  NOR2_X1 U22349 ( .A1(n19505), .A2(n19440), .ZN(n19405) );
  AOI22_X1 U22350 ( .A1(n19755), .A2(n19431), .B1(n19687), .B2(n19405), .ZN(
        n19391) );
  OAI21_X1 U22351 ( .B1(n19445), .B2(n19640), .A(n12682), .ZN(n19389) );
  INV_X1 U22352 ( .A(n19389), .ZN(n19385) );
  NOR2_X1 U22353 ( .A1(n19384), .A2(n19405), .ZN(n19387) );
  AOI22_X1 U22354 ( .A1(n19385), .A2(n19388), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n19387), .ZN(n19386) );
  OAI211_X1 U22355 ( .C1(n19405), .C2(n19576), .A(n19386), .B(n19753), .ZN(
        n19407) );
  OAI22_X1 U22356 ( .A1(n19389), .A2(n19388), .B1(n19387), .B2(n19441), .ZN(
        n19406) );
  AOI22_X1 U22357 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19407), .B1(
        n19694), .B2(n19406), .ZN(n19390) );
  OAI211_X1 U22358 ( .C1(n19758), .C2(n19410), .A(n19391), .B(n19390), .ZN(
        P2_U3088) );
  AOI22_X1 U22359 ( .A1(n19431), .A2(n19762), .B1(n19609), .B2(n19405), .ZN(
        n19393) );
  AOI22_X1 U22360 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19407), .B1(
        n19699), .B2(n19406), .ZN(n19392) );
  OAI211_X1 U22361 ( .C1(n19765), .C2(n19410), .A(n19393), .B(n19392), .ZN(
        P2_U3089) );
  AOI22_X1 U22362 ( .A1(n19398), .A2(n19769), .B1(n19703), .B2(n19405), .ZN(
        n19395) );
  AOI22_X1 U22363 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19407), .B1(
        n19706), .B2(n19406), .ZN(n19394) );
  OAI211_X1 U22364 ( .C1(n19772), .C2(n19439), .A(n19395), .B(n19394), .ZN(
        P2_U3090) );
  AOI22_X1 U22365 ( .A1(n19398), .A2(n19776), .B1(n19614), .B2(n19405), .ZN(
        n19397) );
  AOI22_X1 U22366 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19407), .B1(
        n19712), .B2(n19406), .ZN(n19396) );
  OAI211_X1 U22367 ( .C1(n19779), .C2(n19439), .A(n19397), .B(n19396), .ZN(
        P2_U3091) );
  AOI22_X1 U22368 ( .A1(n19398), .A2(n19716), .B1(n19715), .B2(n19405), .ZN(
        n19400) );
  AOI22_X1 U22369 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19407), .B1(
        n19717), .B2(n19406), .ZN(n19399) );
  OAI211_X1 U22370 ( .C1(n19720), .C2(n19439), .A(n19400), .B(n19399), .ZN(
        P2_U3092) );
  AOI22_X1 U22371 ( .A1(n19431), .A2(n19790), .B1(n19620), .B2(n19405), .ZN(
        n19402) );
  AOI22_X1 U22372 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19407), .B1(
        n19723), .B2(n19406), .ZN(n19401) );
  OAI211_X1 U22373 ( .C1(n19793), .C2(n19410), .A(n19402), .B(n19401), .ZN(
        P2_U3093) );
  AOI22_X1 U22374 ( .A1(n19623), .A2(n19431), .B1(n19727), .B2(n19405), .ZN(
        n19404) );
  AOI22_X1 U22375 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19407), .B1(
        n19729), .B2(n19406), .ZN(n19403) );
  OAI211_X1 U22376 ( .C1(n19626), .C2(n19410), .A(n19404), .B(n19403), .ZN(
        P2_U3094) );
  AOI22_X1 U22377 ( .A1(n19808), .A2(n19431), .B1(n19733), .B2(n19405), .ZN(
        n19409) );
  AOI22_X1 U22378 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19407), .B1(
        n19735), .B2(n19406), .ZN(n19408) );
  OAI211_X1 U22379 ( .C1(n19814), .C2(n19410), .A(n19409), .B(n19408), .ZN(
        P2_U3095) );
  NOR2_X1 U22380 ( .A1(n19538), .A2(n19440), .ZN(n19434) );
  OAI21_X1 U22381 ( .B1(n10595), .B2(n19434), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19411) );
  OAI21_X1 U22382 ( .B1(n19540), .B2(n19440), .A(n19411), .ZN(n19435) );
  AOI22_X1 U22383 ( .A1(n19435), .A2(n19694), .B1(n19687), .B2(n19434), .ZN(
        n19420) );
  INV_X1 U22384 ( .A(n10595), .ZN(n19412) );
  AOI21_X1 U22385 ( .B1(n19412), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19418) );
  NAND2_X1 U22386 ( .A1(n19415), .A2(n19414), .ZN(n19416) );
  OAI221_X1 U22387 ( .B1(n19898), .B2(n19439), .C1(n19898), .C2(n19470), .A(
        n19416), .ZN(n19417) );
  OAI211_X1 U22388 ( .C1(n19418), .C2(n19434), .A(n19417), .B(n19753), .ZN(
        n19436) );
  AOI22_X1 U22389 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19436), .B1(
        n19459), .B2(n19755), .ZN(n19419) );
  OAI211_X1 U22390 ( .C1(n19758), .C2(n19439), .A(n19420), .B(n19419), .ZN(
        P2_U3096) );
  AOI22_X1 U22391 ( .A1(n19435), .A2(n19699), .B1(n19609), .B2(n19434), .ZN(
        n19422) );
  AOI22_X1 U22392 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19436), .B1(
        n19459), .B2(n19762), .ZN(n19421) );
  OAI211_X1 U22393 ( .C1(n19765), .C2(n19439), .A(n19422), .B(n19421), .ZN(
        P2_U3097) );
  AOI22_X1 U22394 ( .A1(n19435), .A2(n19706), .B1(n19703), .B2(n19434), .ZN(
        n19424) );
  AOI22_X1 U22395 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19436), .B1(
        n19431), .B2(n19769), .ZN(n19423) );
  OAI211_X1 U22396 ( .C1(n19772), .C2(n19470), .A(n19424), .B(n19423), .ZN(
        P2_U3098) );
  AOI22_X1 U22397 ( .A1(n19435), .A2(n19712), .B1(n19614), .B2(n19434), .ZN(
        n19426) );
  AOI22_X1 U22398 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19436), .B1(
        n19431), .B2(n19776), .ZN(n19425) );
  OAI211_X1 U22399 ( .C1(n19779), .C2(n19470), .A(n19426), .B(n19425), .ZN(
        P2_U3099) );
  AOI22_X1 U22400 ( .A1(n19435), .A2(n19717), .B1(n19715), .B2(n19434), .ZN(
        n19428) );
  AOI22_X1 U22401 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19436), .B1(
        n19431), .B2(n19716), .ZN(n19427) );
  OAI211_X1 U22402 ( .C1(n19720), .C2(n19470), .A(n19428), .B(n19427), .ZN(
        P2_U3100) );
  AOI22_X1 U22403 ( .A1(n19435), .A2(n19723), .B1(n19620), .B2(n19434), .ZN(
        n19430) );
  AOI22_X1 U22404 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19436), .B1(
        n19459), .B2(n19790), .ZN(n19429) );
  OAI211_X1 U22405 ( .C1(n19793), .C2(n19439), .A(n19430), .B(n19429), .ZN(
        P2_U3101) );
  AOI22_X1 U22406 ( .A1(n19435), .A2(n19729), .B1(n19727), .B2(n19434), .ZN(
        n19433) );
  AOI22_X1 U22407 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19436), .B1(
        n19431), .B2(n19797), .ZN(n19432) );
  OAI211_X1 U22408 ( .C1(n19802), .C2(n19470), .A(n19433), .B(n19432), .ZN(
        P2_U3102) );
  AOI22_X1 U22409 ( .A1(n19435), .A2(n19735), .B1(n19733), .B2(n19434), .ZN(
        n19438) );
  AOI22_X1 U22410 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19436), .B1(
        n19459), .B2(n19808), .ZN(n19437) );
  OAI211_X1 U22411 ( .C1(n19814), .C2(n19439), .A(n19438), .B(n19437), .ZN(
        P2_U3103) );
  NOR2_X1 U22412 ( .A1(n19566), .A2(n19440), .ZN(n19476) );
  NOR2_X1 U22413 ( .A1(n19742), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19449) );
  INV_X1 U22414 ( .A(n19449), .ZN(n19443) );
  OAI21_X1 U22415 ( .B1(n19443), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19441), 
        .ZN(n19444) );
  AOI22_X1 U22416 ( .A1(n19466), .A2(n19694), .B1(n19476), .B2(n19687), .ZN(
        n19452) );
  NOR2_X1 U22417 ( .A1(n19445), .A2(n19899), .ZN(n19897) );
  OAI211_X1 U22418 ( .C1(n19476), .C2(n19576), .A(n19446), .B(n19753), .ZN(
        n19447) );
  INV_X1 U22419 ( .A(n19447), .ZN(n19448) );
  OAI21_X1 U22420 ( .B1(n19897), .B2(n19449), .A(n19448), .ZN(n19467) );
  AOI22_X1 U22421 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19467), .B1(
        n19471), .B2(n19755), .ZN(n19451) );
  OAI211_X1 U22422 ( .C1(n19758), .C2(n19470), .A(n19452), .B(n19451), .ZN(
        P2_U3104) );
  AOI22_X1 U22423 ( .A1(n19466), .A2(n19699), .B1(n19476), .B2(n19609), .ZN(
        n19454) );
  AOI22_X1 U22424 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19467), .B1(
        n19459), .B2(n19650), .ZN(n19453) );
  OAI211_X1 U22425 ( .C1(n19653), .C2(n19504), .A(n19454), .B(n19453), .ZN(
        P2_U3105) );
  AOI22_X1 U22426 ( .A1(n19466), .A2(n19706), .B1(n19476), .B2(n19703), .ZN(
        n19456) );
  AOI22_X1 U22427 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19467), .B1(
        n19459), .B2(n19769), .ZN(n19455) );
  OAI211_X1 U22428 ( .C1(n19772), .C2(n19504), .A(n19456), .B(n19455), .ZN(
        P2_U3106) );
  AOI22_X1 U22429 ( .A1(n19466), .A2(n19712), .B1(n19476), .B2(n19614), .ZN(
        n19458) );
  AOI22_X1 U22430 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19467), .B1(
        n19471), .B2(n19615), .ZN(n19457) );
  OAI211_X1 U22431 ( .C1(n19710), .C2(n19470), .A(n19458), .B(n19457), .ZN(
        P2_U3107) );
  AOI22_X1 U22432 ( .A1(n19466), .A2(n19717), .B1(n19476), .B2(n19715), .ZN(
        n19461) );
  AOI22_X1 U22433 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19467), .B1(
        n19459), .B2(n19716), .ZN(n19460) );
  OAI211_X1 U22434 ( .C1(n19720), .C2(n19504), .A(n19461), .B(n19460), .ZN(
        P2_U3108) );
  AOI22_X1 U22435 ( .A1(n19466), .A2(n19723), .B1(n19476), .B2(n19620), .ZN(
        n19463) );
  AOI22_X1 U22436 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19467), .B1(
        n19471), .B2(n19790), .ZN(n19462) );
  OAI211_X1 U22437 ( .C1(n19793), .C2(n19470), .A(n19463), .B(n19462), .ZN(
        P2_U3109) );
  AOI22_X1 U22438 ( .A1(n19466), .A2(n19729), .B1(n19476), .B2(n19727), .ZN(
        n19465) );
  AOI22_X1 U22439 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19467), .B1(
        n19471), .B2(n19623), .ZN(n19464) );
  OAI211_X1 U22440 ( .C1(n19626), .C2(n19470), .A(n19465), .B(n19464), .ZN(
        P2_U3110) );
  AOI22_X1 U22441 ( .A1(n19466), .A2(n19735), .B1(n19476), .B2(n19733), .ZN(
        n19469) );
  AOI22_X1 U22442 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19467), .B1(
        n19471), .B2(n19808), .ZN(n19468) );
  OAI211_X1 U22443 ( .C1(n19814), .C2(n19470), .A(n19469), .B(n19468), .ZN(
        P2_U3111) );
  NAND2_X1 U22444 ( .A1(n19915), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19569) );
  NOR2_X1 U22445 ( .A1(n19569), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19509) );
  INV_X1 U22446 ( .A(n19509), .ZN(n19512) );
  NOR2_X1 U22447 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19512), .ZN(
        n19499) );
  AOI22_X1 U22448 ( .A1(n19755), .A2(n19530), .B1(n19687), .B2(n19499), .ZN(
        n19482) );
  OAI21_X1 U22449 ( .B1(n19530), .B2(n19471), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19472) );
  NAND2_X1 U22450 ( .A1(n19472), .A2(n12682), .ZN(n19480) );
  NOR2_X1 U22451 ( .A1(n19480), .A2(n19476), .ZN(n19473) );
  AOI211_X1 U22452 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19474), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19473), .ZN(n19475) );
  OAI21_X1 U22453 ( .B1(n19499), .B2(n19475), .A(n19753), .ZN(n19501) );
  NOR2_X1 U22454 ( .A1(n19476), .A2(n19499), .ZN(n19479) );
  OAI21_X1 U22455 ( .B1(n19477), .B2(n19499), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19478) );
  AOI22_X1 U22456 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19501), .B1(
        n19694), .B2(n19500), .ZN(n19481) );
  OAI211_X1 U22457 ( .C1(n19758), .C2(n19504), .A(n19482), .B(n19481), .ZN(
        P2_U3112) );
  INV_X1 U22458 ( .A(n19499), .ZN(n19493) );
  OAI22_X1 U22459 ( .A1(n19537), .A2(n19653), .B1(n19759), .B2(n19493), .ZN(
        n19483) );
  INV_X1 U22460 ( .A(n19483), .ZN(n19485) );
  AOI22_X1 U22461 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19501), .B1(
        n19500), .B2(n19699), .ZN(n19484) );
  OAI211_X1 U22462 ( .C1(n19765), .C2(n19504), .A(n19485), .B(n19484), .ZN(
        P2_U3113) );
  AOI22_X1 U22463 ( .A1(n19704), .A2(n19530), .B1(n19703), .B2(n19499), .ZN(
        n19487) );
  AOI22_X1 U22464 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19501), .B1(
        n19500), .B2(n19706), .ZN(n19486) );
  OAI211_X1 U22465 ( .C1(n19709), .C2(n19504), .A(n19487), .B(n19486), .ZN(
        P2_U3114) );
  OAI22_X1 U22466 ( .A1(n19537), .A2(n19779), .B1(n19773), .B2(n19493), .ZN(
        n19488) );
  INV_X1 U22467 ( .A(n19488), .ZN(n19490) );
  AOI22_X1 U22468 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19501), .B1(
        n19500), .B2(n19712), .ZN(n19489) );
  OAI211_X1 U22469 ( .C1(n19710), .C2(n19504), .A(n19490), .B(n19489), .ZN(
        P2_U3115) );
  AOI22_X1 U22470 ( .A1(n19783), .A2(n19530), .B1(n19715), .B2(n19499), .ZN(
        n19492) );
  AOI22_X1 U22471 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19501), .B1(
        n19500), .B2(n19717), .ZN(n19491) );
  OAI211_X1 U22472 ( .C1(n19786), .C2(n19504), .A(n19492), .B(n19491), .ZN(
        P2_U3116) );
  OAI22_X1 U22473 ( .A1(n19537), .A2(n19726), .B1(n19787), .B2(n19493), .ZN(
        n19494) );
  INV_X1 U22474 ( .A(n19494), .ZN(n19496) );
  AOI22_X1 U22475 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19501), .B1(
        n19500), .B2(n19723), .ZN(n19495) );
  OAI211_X1 U22476 ( .C1(n19793), .C2(n19504), .A(n19496), .B(n19495), .ZN(
        P2_U3117) );
  AOI22_X1 U22477 ( .A1(n19623), .A2(n19530), .B1(n19727), .B2(n19499), .ZN(
        n19498) );
  AOI22_X1 U22478 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19501), .B1(
        n19500), .B2(n19729), .ZN(n19497) );
  OAI211_X1 U22479 ( .C1(n19626), .C2(n19504), .A(n19498), .B(n19497), .ZN(
        P2_U3118) );
  AOI22_X1 U22480 ( .A1(n19808), .A2(n19530), .B1(n19733), .B2(n19499), .ZN(
        n19503) );
  AOI22_X1 U22481 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19501), .B1(
        n19500), .B2(n19735), .ZN(n19502) );
  OAI211_X1 U22482 ( .C1(n19814), .C2(n19504), .A(n19503), .B(n19502), .ZN(
        P2_U3119) );
  NOR2_X1 U22483 ( .A1(n19505), .A2(n19569), .ZN(n19541) );
  AOI22_X1 U22484 ( .A1(n19530), .A2(n19688), .B1(n19687), .B2(n19541), .ZN(
        n19515) );
  NAND2_X1 U22485 ( .A1(n19902), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19639) );
  OAI21_X1 U22486 ( .B1(n19639), .B2(n19506), .A(n12682), .ZN(n19513) );
  INV_X1 U22487 ( .A(n19510), .ZN(n19507) );
  INV_X1 U22488 ( .A(n19541), .ZN(n19526) );
  OAI211_X1 U22489 ( .C1(n19507), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19526), 
        .B(n19679), .ZN(n19508) );
  OAI211_X1 U22490 ( .C1(n19513), .C2(n19509), .A(n19753), .B(n19508), .ZN(
        n19534) );
  OAI21_X1 U22491 ( .B1(n19510), .B2(n19541), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19511) );
  OAI21_X1 U22492 ( .B1(n19513), .B2(n19512), .A(n19511), .ZN(n19533) );
  AOI22_X1 U22493 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19534), .B1(
        n19694), .B2(n19533), .ZN(n19514) );
  OAI211_X1 U22494 ( .C1(n19648), .C2(n19565), .A(n19515), .B(n19514), .ZN(
        P2_U3120) );
  OAI22_X1 U22495 ( .A1(n19537), .A2(n19765), .B1(n19759), .B2(n19526), .ZN(
        n19516) );
  INV_X1 U22496 ( .A(n19516), .ZN(n19518) );
  AOI22_X1 U22497 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19534), .B1(
        n19699), .B2(n19533), .ZN(n19517) );
  OAI211_X1 U22498 ( .C1(n19653), .C2(n19565), .A(n19518), .B(n19517), .ZN(
        P2_U3121) );
  AOI22_X1 U22499 ( .A1(n19704), .A2(n19542), .B1(n19703), .B2(n19541), .ZN(
        n19520) );
  AOI22_X1 U22500 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19534), .B1(
        n19706), .B2(n19533), .ZN(n19519) );
  OAI211_X1 U22501 ( .C1(n19709), .C2(n19537), .A(n19520), .B(n19519), .ZN(
        P2_U3122) );
  OAI22_X1 U22502 ( .A1(n19537), .A2(n19710), .B1(n19773), .B2(n19526), .ZN(
        n19521) );
  INV_X1 U22503 ( .A(n19521), .ZN(n19523) );
  AOI22_X1 U22504 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19534), .B1(
        n19712), .B2(n19533), .ZN(n19522) );
  OAI211_X1 U22505 ( .C1(n19779), .C2(n19565), .A(n19523), .B(n19522), .ZN(
        P2_U3123) );
  AOI22_X1 U22506 ( .A1(n19783), .A2(n19542), .B1(n19715), .B2(n19541), .ZN(
        n19525) );
  AOI22_X1 U22507 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19534), .B1(
        n19717), .B2(n19533), .ZN(n19524) );
  OAI211_X1 U22508 ( .C1(n19786), .C2(n19537), .A(n19525), .B(n19524), .ZN(
        P2_U3124) );
  OAI22_X1 U22509 ( .A1(n19537), .A2(n19793), .B1(n19787), .B2(n19526), .ZN(
        n19527) );
  INV_X1 U22510 ( .A(n19527), .ZN(n19529) );
  AOI22_X1 U22511 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19534), .B1(
        n19723), .B2(n19533), .ZN(n19528) );
  OAI211_X1 U22512 ( .C1(n19726), .C2(n19565), .A(n19529), .B(n19528), .ZN(
        P2_U3125) );
  AOI22_X1 U22513 ( .A1(n19530), .A2(n19797), .B1(n19727), .B2(n19541), .ZN(
        n19532) );
  AOI22_X1 U22514 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19534), .B1(
        n19729), .B2(n19533), .ZN(n19531) );
  OAI211_X1 U22515 ( .C1(n19802), .C2(n19565), .A(n19532), .B(n19531), .ZN(
        P2_U3126) );
  AOI22_X1 U22516 ( .A1(n19808), .A2(n19542), .B1(n19733), .B2(n19541), .ZN(
        n19536) );
  AOI22_X1 U22517 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19534), .B1(
        n19735), .B2(n19533), .ZN(n19535) );
  OAI211_X1 U22518 ( .C1(n19814), .C2(n19537), .A(n19536), .B(n19535), .ZN(
        P2_U3127) );
  NOR2_X1 U22519 ( .A1(n19538), .A2(n19569), .ZN(n19560) );
  OAI21_X1 U22520 ( .B1(n9730), .B2(n19560), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19539) );
  OAI21_X1 U22521 ( .B1(n19569), .B2(n19540), .A(n19539), .ZN(n19561) );
  AOI22_X1 U22522 ( .A1(n19561), .A2(n19694), .B1(n19687), .B2(n19560), .ZN(
        n19547) );
  NOR2_X2 U22523 ( .A1(n19678), .A2(n19572), .ZN(n19591) );
  AOI221_X1 U22524 ( .B1(n19591), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19542), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19541), .ZN(n19543) );
  AOI211_X1 U22525 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19544), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19543), .ZN(n19545) );
  OAI21_X1 U22526 ( .B1(n19545), .B2(n19560), .A(n19753), .ZN(n19562) );
  AOI22_X1 U22527 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19562), .B1(
        n19591), .B2(n19755), .ZN(n19546) );
  OAI211_X1 U22528 ( .C1(n19758), .C2(n19565), .A(n19547), .B(n19546), .ZN(
        P2_U3128) );
  AOI22_X1 U22529 ( .A1(n19561), .A2(n19699), .B1(n19609), .B2(n19560), .ZN(
        n19549) );
  AOI22_X1 U22530 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19562), .B1(
        n19591), .B2(n19762), .ZN(n19548) );
  OAI211_X1 U22531 ( .C1(n19765), .C2(n19565), .A(n19549), .B(n19548), .ZN(
        P2_U3129) );
  AOI22_X1 U22532 ( .A1(n19561), .A2(n19706), .B1(n19703), .B2(n19560), .ZN(
        n19551) );
  AOI22_X1 U22533 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19562), .B1(
        n19591), .B2(n19704), .ZN(n19550) );
  OAI211_X1 U22534 ( .C1(n19709), .C2(n19565), .A(n19551), .B(n19550), .ZN(
        P2_U3130) );
  AOI22_X1 U22535 ( .A1(n19561), .A2(n19712), .B1(n19614), .B2(n19560), .ZN(
        n19553) );
  AOI22_X1 U22536 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19562), .B1(
        n19591), .B2(n19615), .ZN(n19552) );
  OAI211_X1 U22537 ( .C1(n19710), .C2(n19565), .A(n19553), .B(n19552), .ZN(
        P2_U3131) );
  AOI22_X1 U22538 ( .A1(n19561), .A2(n19717), .B1(n19715), .B2(n19560), .ZN(
        n19555) );
  AOI22_X1 U22539 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19562), .B1(
        n19591), .B2(n19783), .ZN(n19554) );
  OAI211_X1 U22540 ( .C1(n19786), .C2(n19565), .A(n19555), .B(n19554), .ZN(
        P2_U3132) );
  AOI22_X1 U22541 ( .A1(n19561), .A2(n19723), .B1(n19620), .B2(n19560), .ZN(
        n19557) );
  AOI22_X1 U22542 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19562), .B1(
        n19591), .B2(n19790), .ZN(n19556) );
  OAI211_X1 U22543 ( .C1(n19793), .C2(n19565), .A(n19557), .B(n19556), .ZN(
        P2_U3133) );
  AOI22_X1 U22544 ( .A1(n19561), .A2(n19729), .B1(n19727), .B2(n19560), .ZN(
        n19559) );
  AOI22_X1 U22545 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19562), .B1(
        n19591), .B2(n19623), .ZN(n19558) );
  OAI211_X1 U22546 ( .C1(n19626), .C2(n19565), .A(n19559), .B(n19558), .ZN(
        P2_U3134) );
  AOI22_X1 U22547 ( .A1(n19561), .A2(n19735), .B1(n19733), .B2(n19560), .ZN(
        n19564) );
  AOI22_X1 U22548 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19562), .B1(
        n19591), .B2(n19808), .ZN(n19563) );
  OAI211_X1 U22549 ( .C1(n19814), .C2(n19565), .A(n19564), .B(n19563), .ZN(
        P2_U3135) );
  NOR2_X1 U22550 ( .A1(n19566), .A2(n19569), .ZN(n19592) );
  NOR2_X1 U22551 ( .A1(n19592), .A2(n19441), .ZN(n19567) );
  NAND2_X1 U22552 ( .A1(n19568), .A2(n19567), .ZN(n19573) );
  OR2_X1 U22553 ( .A1(n19924), .A2(n19569), .ZN(n19571) );
  OAI21_X1 U22554 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19571), .A(n19441), 
        .ZN(n19570) );
  AND2_X1 U22555 ( .A1(n19573), .A2(n19570), .ZN(n19593) );
  AOI22_X1 U22556 ( .A1(n19593), .A2(n19694), .B1(n19687), .B2(n19592), .ZN(
        n19578) );
  OAI21_X1 U22557 ( .B1(n19639), .B2(n19572), .A(n19571), .ZN(n19574) );
  AND2_X1 U22558 ( .A1(n19574), .A2(n19573), .ZN(n19575) );
  OAI211_X1 U22559 ( .C1(n19592), .C2(n19576), .A(n19575), .B(n19753), .ZN(
        n19594) );
  AOI22_X1 U22560 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19594), .B1(
        n19591), .B2(n19688), .ZN(n19577) );
  OAI211_X1 U22561 ( .C1(n19648), .C2(n19632), .A(n19578), .B(n19577), .ZN(
        P2_U3136) );
  AOI22_X1 U22562 ( .A1(n19593), .A2(n19699), .B1(n19609), .B2(n19592), .ZN(
        n19580) );
  AOI22_X1 U22563 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19594), .B1(
        n19591), .B2(n19650), .ZN(n19579) );
  OAI211_X1 U22564 ( .C1(n19653), .C2(n19632), .A(n19580), .B(n19579), .ZN(
        P2_U3137) );
  AOI22_X1 U22565 ( .A1(n19593), .A2(n19706), .B1(n19703), .B2(n19592), .ZN(
        n19582) );
  AOI22_X1 U22566 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19594), .B1(
        n19591), .B2(n19769), .ZN(n19581) );
  OAI211_X1 U22567 ( .C1(n19772), .C2(n19632), .A(n19582), .B(n19581), .ZN(
        P2_U3138) );
  AOI22_X1 U22568 ( .A1(n19593), .A2(n19712), .B1(n19614), .B2(n19592), .ZN(
        n19584) );
  AOI22_X1 U22569 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19594), .B1(
        n19591), .B2(n19776), .ZN(n19583) );
  OAI211_X1 U22570 ( .C1(n19779), .C2(n19632), .A(n19584), .B(n19583), .ZN(
        P2_U3139) );
  AOI22_X1 U22571 ( .A1(n19593), .A2(n19717), .B1(n19715), .B2(n19592), .ZN(
        n19586) );
  AOI22_X1 U22572 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19594), .B1(
        n19591), .B2(n19716), .ZN(n19585) );
  OAI211_X1 U22573 ( .C1(n19720), .C2(n19632), .A(n19586), .B(n19585), .ZN(
        P2_U3140) );
  AOI22_X1 U22574 ( .A1(n19593), .A2(n19723), .B1(n19620), .B2(n19592), .ZN(
        n19588) );
  AOI22_X1 U22575 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19594), .B1(
        n19591), .B2(n19664), .ZN(n19587) );
  OAI211_X1 U22576 ( .C1(n19726), .C2(n19632), .A(n19588), .B(n19587), .ZN(
        P2_U3141) );
  AOI22_X1 U22577 ( .A1(n19593), .A2(n19729), .B1(n19727), .B2(n19592), .ZN(
        n19590) );
  AOI22_X1 U22578 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19594), .B1(
        n19591), .B2(n19797), .ZN(n19589) );
  OAI211_X1 U22579 ( .C1(n19802), .C2(n19632), .A(n19590), .B(n19589), .ZN(
        P2_U3142) );
  INV_X1 U22580 ( .A(n19591), .ZN(n19597) );
  AOI22_X1 U22581 ( .A1(n19593), .A2(n19735), .B1(n19733), .B2(n19592), .ZN(
        n19596) );
  AOI22_X1 U22582 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19594), .B1(
        n19602), .B2(n19808), .ZN(n19595) );
  OAI211_X1 U22583 ( .C1(n19814), .C2(n19597), .A(n19596), .B(n19595), .ZN(
        P2_U3143) );
  NAND3_X1 U22584 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19924), .ZN(n19643) );
  NOR2_X1 U22585 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19643), .ZN(
        n19627) );
  OAI21_X1 U22586 ( .B1(n19600), .B2(n19627), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19598) );
  OAI21_X1 U22587 ( .B1(n19599), .B2(n19604), .A(n19598), .ZN(n19628) );
  AOI22_X1 U22588 ( .A1(n19628), .A2(n19694), .B1(n19687), .B2(n19627), .ZN(
        n19608) );
  INV_X1 U22589 ( .A(n19600), .ZN(n19601) );
  AOI21_X1 U22590 ( .B1(n19601), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19606) );
  NOR2_X2 U22591 ( .A1(n19678), .A2(n19640), .ZN(n19670) );
  OAI21_X1 U22592 ( .B1(n19670), .B2(n19602), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19603) );
  OAI21_X1 U22593 ( .B1(n19604), .B2(n19908), .A(n19603), .ZN(n19605) );
  OAI211_X1 U22594 ( .C1(n19627), .C2(n19606), .A(n19605), .B(n19753), .ZN(
        n19629) );
  AOI22_X1 U22595 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19629), .B1(
        n19670), .B2(n19755), .ZN(n19607) );
  OAI211_X1 U22596 ( .C1(n19758), .C2(n19632), .A(n19608), .B(n19607), .ZN(
        P2_U3144) );
  AOI22_X1 U22597 ( .A1(n19628), .A2(n19699), .B1(n19609), .B2(n19627), .ZN(
        n19611) );
  AOI22_X1 U22598 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19629), .B1(
        n19670), .B2(n19762), .ZN(n19610) );
  OAI211_X1 U22599 ( .C1(n19765), .C2(n19632), .A(n19611), .B(n19610), .ZN(
        P2_U3145) );
  AOI22_X1 U22600 ( .A1(n19628), .A2(n19706), .B1(n19703), .B2(n19627), .ZN(
        n19613) );
  AOI22_X1 U22601 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19629), .B1(
        n19670), .B2(n19704), .ZN(n19612) );
  OAI211_X1 U22602 ( .C1(n19709), .C2(n19632), .A(n19613), .B(n19612), .ZN(
        P2_U3146) );
  AOI22_X1 U22603 ( .A1(n19628), .A2(n19712), .B1(n19614), .B2(n19627), .ZN(
        n19617) );
  AOI22_X1 U22604 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19629), .B1(
        n19670), .B2(n19615), .ZN(n19616) );
  OAI211_X1 U22605 ( .C1(n19710), .C2(n19632), .A(n19617), .B(n19616), .ZN(
        P2_U3147) );
  AOI22_X1 U22606 ( .A1(n19628), .A2(n19717), .B1(n19715), .B2(n19627), .ZN(
        n19619) );
  AOI22_X1 U22607 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19629), .B1(
        n19670), .B2(n19783), .ZN(n19618) );
  OAI211_X1 U22608 ( .C1(n19786), .C2(n19632), .A(n19619), .B(n19618), .ZN(
        P2_U3148) );
  AOI22_X1 U22609 ( .A1(n19628), .A2(n19723), .B1(n19620), .B2(n19627), .ZN(
        n19622) );
  AOI22_X1 U22610 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19629), .B1(
        n19670), .B2(n19790), .ZN(n19621) );
  OAI211_X1 U22611 ( .C1(n19793), .C2(n19632), .A(n19622), .B(n19621), .ZN(
        P2_U3149) );
  AOI22_X1 U22612 ( .A1(n19628), .A2(n19729), .B1(n19727), .B2(n19627), .ZN(
        n19625) );
  AOI22_X1 U22613 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19629), .B1(
        n19670), .B2(n19623), .ZN(n19624) );
  OAI211_X1 U22614 ( .C1(n19626), .C2(n19632), .A(n19625), .B(n19624), .ZN(
        P2_U3150) );
  AOI22_X1 U22615 ( .A1(n19628), .A2(n19735), .B1(n19733), .B2(n19627), .ZN(
        n19631) );
  AOI22_X1 U22616 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19629), .B1(
        n19670), .B2(n19808), .ZN(n19630) );
  OAI211_X1 U22617 ( .C1(n19814), .C2(n19632), .A(n19631), .B(n19630), .ZN(
        P2_U3151) );
  NOR2_X1 U22618 ( .A1(n19933), .A2(n19643), .ZN(n19681) );
  INV_X1 U22619 ( .A(n19681), .ZN(n19671) );
  NAND2_X1 U22620 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19671), .ZN(n19634) );
  NOR2_X1 U22621 ( .A1(n19635), .A2(n19634), .ZN(n19642) );
  INV_X1 U22622 ( .A(n19643), .ZN(n19636) );
  AOI21_X1 U22623 ( .B1(n19576), .B2(n19636), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19637) );
  OR2_X1 U22624 ( .A1(n19642), .A2(n19637), .ZN(n19672) );
  INV_X1 U22625 ( .A(n19694), .ZN(n19746) );
  INV_X1 U22626 ( .A(n19687), .ZN(n19745) );
  OAI22_X1 U22627 ( .A1(n19672), .A2(n19746), .B1(n19745), .B2(n19671), .ZN(
        n19638) );
  INV_X1 U22628 ( .A(n19638), .ZN(n19647) );
  INV_X1 U22629 ( .A(n19639), .ZN(n19749) );
  INV_X1 U22630 ( .A(n19640), .ZN(n19641) );
  NAND2_X1 U22631 ( .A1(n19749), .A2(n19641), .ZN(n19644) );
  AOI21_X1 U22632 ( .B1(n19644), .B2(n19643), .A(n19642), .ZN(n19645) );
  OAI211_X1 U22633 ( .C1(n19681), .C2(n19576), .A(n19645), .B(n19753), .ZN(
        n19674) );
  AOI22_X1 U22634 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19674), .B1(
        n19670), .B2(n19688), .ZN(n19646) );
  OAI211_X1 U22635 ( .C1(n19648), .C2(n19739), .A(n19647), .B(n19646), .ZN(
        P2_U3152) );
  INV_X1 U22636 ( .A(n19699), .ZN(n19760) );
  OAI22_X1 U22637 ( .A1(n19672), .A2(n19760), .B1(n19759), .B2(n19671), .ZN(
        n19649) );
  INV_X1 U22638 ( .A(n19649), .ZN(n19652) );
  AOI22_X1 U22639 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19674), .B1(
        n19670), .B2(n19650), .ZN(n19651) );
  OAI211_X1 U22640 ( .C1(n19653), .C2(n19739), .A(n19652), .B(n19651), .ZN(
        P2_U3153) );
  INV_X1 U22641 ( .A(n19706), .ZN(n19767) );
  INV_X1 U22642 ( .A(n19703), .ZN(n19766) );
  OAI22_X1 U22643 ( .A1(n19672), .A2(n19767), .B1(n19766), .B2(n19671), .ZN(
        n19654) );
  INV_X1 U22644 ( .A(n19654), .ZN(n19656) );
  AOI22_X1 U22645 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19674), .B1(
        n19670), .B2(n19769), .ZN(n19655) );
  OAI211_X1 U22646 ( .C1(n19772), .C2(n19739), .A(n19656), .B(n19655), .ZN(
        P2_U3154) );
  INV_X1 U22647 ( .A(n19712), .ZN(n19774) );
  OAI22_X1 U22648 ( .A1(n19672), .A2(n19774), .B1(n19773), .B2(n19671), .ZN(
        n19657) );
  INV_X1 U22649 ( .A(n19657), .ZN(n19659) );
  AOI22_X1 U22650 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19674), .B1(
        n19670), .B2(n19776), .ZN(n19658) );
  OAI211_X1 U22651 ( .C1(n19779), .C2(n19739), .A(n19659), .B(n19658), .ZN(
        P2_U3155) );
  INV_X1 U22652 ( .A(n19717), .ZN(n19781) );
  INV_X1 U22653 ( .A(n19715), .ZN(n19780) );
  OAI22_X1 U22654 ( .A1(n19672), .A2(n19781), .B1(n19780), .B2(n19671), .ZN(
        n19660) );
  INV_X1 U22655 ( .A(n19660), .ZN(n19662) );
  AOI22_X1 U22656 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19674), .B1(
        n19670), .B2(n19716), .ZN(n19661) );
  OAI211_X1 U22657 ( .C1(n19720), .C2(n19739), .A(n19662), .B(n19661), .ZN(
        P2_U3156) );
  INV_X1 U22658 ( .A(n19723), .ZN(n19788) );
  OAI22_X1 U22659 ( .A1(n19672), .A2(n19788), .B1(n19787), .B2(n19671), .ZN(
        n19663) );
  INV_X1 U22660 ( .A(n19663), .ZN(n19666) );
  AOI22_X1 U22661 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19674), .B1(
        n19670), .B2(n19664), .ZN(n19665) );
  OAI211_X1 U22662 ( .C1(n19726), .C2(n19739), .A(n19666), .B(n19665), .ZN(
        P2_U3157) );
  INV_X1 U22663 ( .A(n19729), .ZN(n19795) );
  INV_X1 U22664 ( .A(n19727), .ZN(n19794) );
  OAI22_X1 U22665 ( .A1(n19672), .A2(n19795), .B1(n19794), .B2(n19671), .ZN(
        n19667) );
  INV_X1 U22666 ( .A(n19667), .ZN(n19669) );
  AOI22_X1 U22667 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19674), .B1(
        n19670), .B2(n19797), .ZN(n19668) );
  OAI211_X1 U22668 ( .C1(n19802), .C2(n19739), .A(n19669), .B(n19668), .ZN(
        P2_U3158) );
  INV_X1 U22669 ( .A(n19670), .ZN(n19677) );
  INV_X1 U22670 ( .A(n19735), .ZN(n19805) );
  INV_X1 U22671 ( .A(n19733), .ZN(n19803) );
  OAI22_X1 U22672 ( .A1(n19672), .A2(n19805), .B1(n19803), .B2(n19671), .ZN(
        n19673) );
  INV_X1 U22673 ( .A(n19673), .ZN(n19676) );
  INV_X1 U22674 ( .A(n19739), .ZN(n19728) );
  AOI22_X1 U22675 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19674), .B1(
        n19728), .B2(n19808), .ZN(n19675) );
  OAI211_X1 U22676 ( .C1(n19814), .C2(n19677), .A(n19676), .B(n19675), .ZN(
        P2_U3159) );
  NAND2_X1 U22677 ( .A1(n19813), .A2(n19739), .ZN(n19680) );
  AOI21_X1 U22678 ( .B1(n19680), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19679), 
        .ZN(n19689) );
  NOR3_X2 U22679 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19908), .A3(
        n19742), .ZN(n19732) );
  NOR2_X1 U22680 ( .A1(n19732), .A2(n19681), .ZN(n19692) );
  NAND2_X1 U22681 ( .A1(n19689), .A2(n19692), .ZN(n19686) );
  NAND2_X1 U22682 ( .A1(n19690), .A2(n19576), .ZN(n19684) );
  NOR2_X1 U22683 ( .A1(n12882), .A2(n19732), .ZN(n19683) );
  AOI21_X1 U22684 ( .B1(n19684), .B2(n19683), .A(n19682), .ZN(n19685) );
  INV_X1 U22685 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n19697) );
  AOI22_X1 U22686 ( .A1(n19728), .A2(n19688), .B1(n19687), .B2(n19732), .ZN(
        n19696) );
  INV_X1 U22687 ( .A(n19689), .ZN(n19693) );
  OAI21_X1 U22688 ( .B1(n19690), .B2(n19732), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19691) );
  AOI22_X1 U22689 ( .A1(n19694), .A2(n19734), .B1(n19798), .B2(n19755), .ZN(
        n19695) );
  OAI211_X1 U22690 ( .C1(n19705), .C2(n19697), .A(n19696), .B(n19695), .ZN(
        P2_U3160) );
  INV_X1 U22691 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n19702) );
  INV_X1 U22692 ( .A(n19732), .ZN(n19721) );
  OAI22_X1 U22693 ( .A1(n19739), .A2(n19765), .B1(n19759), .B2(n19721), .ZN(
        n19698) );
  INV_X1 U22694 ( .A(n19698), .ZN(n19701) );
  AOI22_X1 U22695 ( .A1(n19699), .A2(n19734), .B1(n19798), .B2(n19762), .ZN(
        n19700) );
  OAI211_X1 U22696 ( .C1(n19705), .C2(n19702), .A(n19701), .B(n19700), .ZN(
        P2_U3161) );
  AOI22_X1 U22697 ( .A1(n19704), .A2(n19798), .B1(n19703), .B2(n19732), .ZN(
        n19708) );
  AOI22_X1 U22698 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19736), .B1(
        n19706), .B2(n19734), .ZN(n19707) );
  OAI211_X1 U22699 ( .C1(n19709), .C2(n19739), .A(n19708), .B(n19707), .ZN(
        P2_U3162) );
  OAI22_X1 U22700 ( .A1(n19739), .A2(n19710), .B1(n19773), .B2(n19721), .ZN(
        n19711) );
  INV_X1 U22701 ( .A(n19711), .ZN(n19714) );
  AOI22_X1 U22702 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19736), .B1(
        n19712), .B2(n19734), .ZN(n19713) );
  OAI211_X1 U22703 ( .C1(n19779), .C2(n19813), .A(n19714), .B(n19713), .ZN(
        P2_U3163) );
  AOI22_X1 U22704 ( .A1(n19728), .A2(n19716), .B1(n19715), .B2(n19732), .ZN(
        n19719) );
  AOI22_X1 U22705 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19736), .B1(
        n19717), .B2(n19734), .ZN(n19718) );
  OAI211_X1 U22706 ( .C1(n19720), .C2(n19813), .A(n19719), .B(n19718), .ZN(
        P2_U3164) );
  OAI22_X1 U22707 ( .A1(n19739), .A2(n19793), .B1(n19787), .B2(n19721), .ZN(
        n19722) );
  INV_X1 U22708 ( .A(n19722), .ZN(n19725) );
  AOI22_X1 U22709 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19736), .B1(
        n19723), .B2(n19734), .ZN(n19724) );
  OAI211_X1 U22710 ( .C1(n19726), .C2(n19813), .A(n19725), .B(n19724), .ZN(
        P2_U3165) );
  AOI22_X1 U22711 ( .A1(n19728), .A2(n19797), .B1(n19727), .B2(n19732), .ZN(
        n19731) );
  AOI22_X1 U22712 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19736), .B1(
        n19729), .B2(n19734), .ZN(n19730) );
  OAI211_X1 U22713 ( .C1(n19802), .C2(n19813), .A(n19731), .B(n19730), .ZN(
        P2_U3166) );
  AOI22_X1 U22714 ( .A1(n19808), .A2(n19798), .B1(n19733), .B2(n19732), .ZN(
        n19738) );
  AOI22_X1 U22715 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19736), .B1(
        n19735), .B2(n19734), .ZN(n19737) );
  OAI211_X1 U22716 ( .C1(n19814), .C2(n19739), .A(n19738), .B(n19737), .ZN(
        P2_U3167) );
  NAND2_X1 U22717 ( .A1(n19804), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19740) );
  NOR2_X1 U22718 ( .A1(n19741), .A2(n19740), .ZN(n19750) );
  OR2_X1 U22719 ( .A1(n19908), .A2(n19742), .ZN(n19751) );
  INV_X1 U22720 ( .A(n19751), .ZN(n19743) );
  AOI21_X1 U22721 ( .B1(n19576), .B2(n19743), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19744) );
  OAI22_X1 U22722 ( .A1(n19806), .A2(n19746), .B1(n19804), .B2(n19745), .ZN(
        n19747) );
  INV_X1 U22723 ( .A(n19747), .ZN(n19757) );
  INV_X1 U22724 ( .A(n19899), .ZN(n19748) );
  NAND2_X1 U22725 ( .A1(n19749), .A2(n19748), .ZN(n19752) );
  AOI21_X1 U22726 ( .B1(n19752), .B2(n19751), .A(n19750), .ZN(n19754) );
  OAI211_X1 U22727 ( .C1(n19213), .C2(n19576), .A(n19754), .B(n19753), .ZN(
        n19810) );
  AOI22_X1 U22728 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19810), .B1(
        n19809), .B2(n19755), .ZN(n19756) );
  OAI211_X1 U22729 ( .C1(n19758), .C2(n19813), .A(n19757), .B(n19756), .ZN(
        P2_U3168) );
  OAI22_X1 U22730 ( .A1(n19806), .A2(n19760), .B1(n19804), .B2(n19759), .ZN(
        n19761) );
  INV_X1 U22731 ( .A(n19761), .ZN(n19764) );
  AOI22_X1 U22732 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19810), .B1(
        n19809), .B2(n19762), .ZN(n19763) );
  OAI211_X1 U22733 ( .C1(n19765), .C2(n19813), .A(n19764), .B(n19763), .ZN(
        P2_U3169) );
  OAI22_X1 U22734 ( .A1(n19806), .A2(n19767), .B1(n19804), .B2(n19766), .ZN(
        n19768) );
  INV_X1 U22735 ( .A(n19768), .ZN(n19771) );
  AOI22_X1 U22736 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19810), .B1(
        n19798), .B2(n19769), .ZN(n19770) );
  OAI211_X1 U22737 ( .C1(n19772), .C2(n19801), .A(n19771), .B(n19770), .ZN(
        P2_U3170) );
  OAI22_X1 U22738 ( .A1(n19806), .A2(n19774), .B1(n19804), .B2(n19773), .ZN(
        n19775) );
  INV_X1 U22739 ( .A(n19775), .ZN(n19778) );
  AOI22_X1 U22740 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19810), .B1(
        n19798), .B2(n19776), .ZN(n19777) );
  OAI211_X1 U22741 ( .C1(n19779), .C2(n19801), .A(n19778), .B(n19777), .ZN(
        P2_U3171) );
  OAI22_X1 U22742 ( .A1(n19806), .A2(n19781), .B1(n19804), .B2(n19780), .ZN(
        n19782) );
  INV_X1 U22743 ( .A(n19782), .ZN(n19785) );
  AOI22_X1 U22744 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19810), .B1(
        n19809), .B2(n19783), .ZN(n19784) );
  OAI211_X1 U22745 ( .C1(n19786), .C2(n19813), .A(n19785), .B(n19784), .ZN(
        P2_U3172) );
  OAI22_X1 U22746 ( .A1(n19806), .A2(n19788), .B1(n19804), .B2(n19787), .ZN(
        n19789) );
  INV_X1 U22747 ( .A(n19789), .ZN(n19792) );
  AOI22_X1 U22748 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19810), .B1(
        n19809), .B2(n19790), .ZN(n19791) );
  OAI211_X1 U22749 ( .C1(n19793), .C2(n19813), .A(n19792), .B(n19791), .ZN(
        P2_U3173) );
  OAI22_X1 U22750 ( .A1(n19806), .A2(n19795), .B1(n19804), .B2(n19794), .ZN(
        n19796) );
  INV_X1 U22751 ( .A(n19796), .ZN(n19800) );
  AOI22_X1 U22752 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19810), .B1(
        n19798), .B2(n19797), .ZN(n19799) );
  OAI211_X1 U22753 ( .C1(n19802), .C2(n19801), .A(n19800), .B(n19799), .ZN(
        P2_U3174) );
  OAI22_X1 U22754 ( .A1(n19806), .A2(n19805), .B1(n19804), .B2(n19803), .ZN(
        n19807) );
  INV_X1 U22755 ( .A(n19807), .ZN(n19812) );
  AOI22_X1 U22756 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19810), .B1(
        n19809), .B2(n19808), .ZN(n19811) );
  OAI211_X1 U22757 ( .C1(n19814), .C2(n19813), .A(n19812), .B(n19811), .ZN(
        P2_U3175) );
  AOI21_X1 U22758 ( .B1(n19817), .B2(n19816), .A(n19815), .ZN(n19821) );
  OAI211_X1 U22759 ( .C1(n19822), .C2(n19818), .A(n19834), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19819) );
  OAI211_X1 U22760 ( .C1(n19822), .C2(n19821), .A(n19820), .B(n19819), .ZN(
        P2_U3177) );
  AND2_X1 U22761 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19823), .ZN(
        P2_U3179) );
  AND2_X1 U22762 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19823), .ZN(
        P2_U3180) );
  AND2_X1 U22763 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19823), .ZN(
        P2_U3181) );
  AND2_X1 U22764 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19823), .ZN(
        P2_U3182) );
  AND2_X1 U22765 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19823), .ZN(
        P2_U3183) );
  AND2_X1 U22766 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19823), .ZN(
        P2_U3184) );
  AND2_X1 U22767 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19823), .ZN(
        P2_U3185) );
  AND2_X1 U22768 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19823), .ZN(
        P2_U3186) );
  AND2_X1 U22769 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19823), .ZN(
        P2_U3187) );
  AND2_X1 U22770 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19823), .ZN(
        P2_U3188) );
  AND2_X1 U22771 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19823), .ZN(
        P2_U3189) );
  AND2_X1 U22772 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19823), .ZN(
        P2_U3190) );
  AND2_X1 U22773 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19823), .ZN(
        P2_U3191) );
  AND2_X1 U22774 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19823), .ZN(
        P2_U3192) );
  AND2_X1 U22775 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19823), .ZN(
        P2_U3193) );
  AND2_X1 U22776 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19823), .ZN(
        P2_U3194) );
  AND2_X1 U22777 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19823), .ZN(
        P2_U3195) );
  AND2_X1 U22778 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19823), .ZN(
        P2_U3196) );
  AND2_X1 U22779 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19823), .ZN(
        P2_U3197) );
  AND2_X1 U22780 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19823), .ZN(
        P2_U3198) );
  AND2_X1 U22781 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19823), .ZN(
        P2_U3199) );
  AND2_X1 U22782 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19823), .ZN(
        P2_U3200) );
  AND2_X1 U22783 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19823), .ZN(P2_U3201) );
  AND2_X1 U22784 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19823), .ZN(P2_U3202) );
  AND2_X1 U22785 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19823), .ZN(P2_U3203) );
  AND2_X1 U22786 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19823), .ZN(P2_U3204) );
  AND2_X1 U22787 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19823), .ZN(P2_U3205) );
  AND2_X1 U22788 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19823), .ZN(P2_U3206) );
  AND2_X1 U22789 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19823), .ZN(P2_U3207) );
  AND2_X1 U22790 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19823), .ZN(P2_U3208) );
  NAND2_X1 U22791 ( .A1(n19834), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19836) );
  NAND3_X1 U22792 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n19836), .ZN(n19826) );
  AOI211_X1 U22793 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n20778), .A(
        n19824), .B(n19944), .ZN(n19825) );
  INV_X1 U22794 ( .A(NA), .ZN(n20788) );
  NOR3_X1 U22795 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n20788), .ZN(n19841) );
  AOI211_X1 U22796 ( .C1(n19842), .C2(n19826), .A(n19825), .B(n19841), .ZN(
        n19827) );
  INV_X1 U22797 ( .A(n19827), .ZN(P2_U3209) );
  AOI21_X1 U22798 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20778), .A(n19842), 
        .ZN(n19833) );
  NOR2_X1 U22799 ( .A1(n18855), .A2(n19833), .ZN(n19829) );
  AOI21_X1 U22800 ( .B1(n19829), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .A(n19828), .ZN(n19830) );
  OAI211_X1 U22801 ( .C1(n20778), .C2(n19831), .A(n19830), .B(n19836), .ZN(
        P2_U3210) );
  NOR2_X1 U22802 ( .A1(n19832), .A2(n19842), .ZN(n19835) );
  AOI21_X1 U22803 ( .B1(n19835), .B2(n19834), .A(n19833), .ZN(n19840) );
  OAI22_X1 U22804 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19837), .B1(NA), 
        .B2(n19836), .ZN(n19838) );
  OAI211_X1 U22805 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19838), .ZN(n19839) );
  OAI21_X1 U22806 ( .B1(n19841), .B2(n19840), .A(n19839), .ZN(P2_U3211) );
  NAND2_X2 U22807 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19944), .ZN(n19886) );
  OAI222_X1 U22808 ( .A1(n19889), .A2(n19845), .B1(n19844), .B2(n19944), .C1(
        n19843), .C2(n19886), .ZN(P2_U3212) );
  OAI222_X1 U22809 ( .A1(n19889), .A2(n13258), .B1(n19846), .B2(n19944), .C1(
        n19845), .C2(n19886), .ZN(P2_U3213) );
  OAI222_X1 U22810 ( .A1(n19889), .A2(n19848), .B1(n19847), .B2(n19944), .C1(
        n13258), .C2(n19886), .ZN(P2_U3214) );
  OAI222_X1 U22811 ( .A1(n19889), .A2(n12101), .B1(n19849), .B2(n19944), .C1(
        n19848), .C2(n19886), .ZN(P2_U3215) );
  OAI222_X1 U22812 ( .A1(n19889), .A2(n19851), .B1(n19850), .B2(n19944), .C1(
        n12101), .C2(n19886), .ZN(P2_U3216) );
  OAI222_X1 U22813 ( .A1(n19889), .A2(n19853), .B1(n19852), .B2(n19944), .C1(
        n19851), .C2(n19886), .ZN(P2_U3217) );
  INV_X1 U22814 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19855) );
  OAI222_X1 U22815 ( .A1(n19889), .A2(n19855), .B1(n19854), .B2(n19944), .C1(
        n19853), .C2(n19886), .ZN(P2_U3218) );
  OAI222_X1 U22816 ( .A1(n19889), .A2(n12161), .B1(n19856), .B2(n19944), .C1(
        n19855), .C2(n19886), .ZN(P2_U3219) );
  OAI222_X1 U22817 ( .A1(n19889), .A2(n19858), .B1(n19857), .B2(n19944), .C1(
        n12161), .C2(n19886), .ZN(P2_U3220) );
  OAI222_X1 U22818 ( .A1(n19889), .A2(n12187), .B1(n19859), .B2(n19944), .C1(
        n19858), .C2(n19886), .ZN(P2_U3221) );
  OAI222_X1 U22819 ( .A1(n19889), .A2(n19861), .B1(n19860), .B2(n19944), .C1(
        n12187), .C2(n19886), .ZN(P2_U3222) );
  OAI222_X1 U22820 ( .A1(n19889), .A2(n15283), .B1(n19862), .B2(n19944), .C1(
        n19861), .C2(n19886), .ZN(P2_U3223) );
  OAI222_X1 U22821 ( .A1(n19889), .A2(n19864), .B1(n19863), .B2(n19944), .C1(
        n15283), .C2(n19886), .ZN(P2_U3224) );
  OAI222_X1 U22822 ( .A1(n19889), .A2(n21120), .B1(n19865), .B2(n19944), .C1(
        n19864), .C2(n19886), .ZN(P2_U3225) );
  OAI222_X1 U22823 ( .A1(n19889), .A2(n15235), .B1(n19866), .B2(n19944), .C1(
        n21120), .C2(n19886), .ZN(P2_U3226) );
  OAI222_X1 U22824 ( .A1(n19889), .A2(n21170), .B1(n19867), .B2(n19944), .C1(
        n15235), .C2(n19886), .ZN(P2_U3227) );
  OAI222_X1 U22825 ( .A1(n19889), .A2(n19869), .B1(n19868), .B2(n19944), .C1(
        n21170), .C2(n19886), .ZN(P2_U3228) );
  OAI222_X1 U22826 ( .A1(n19889), .A2(n19871), .B1(n19870), .B2(n19944), .C1(
        n19869), .C2(n19886), .ZN(P2_U3229) );
  OAI222_X1 U22827 ( .A1(n19889), .A2(n14972), .B1(n19872), .B2(n19944), .C1(
        n19871), .C2(n19886), .ZN(P2_U3230) );
  OAI222_X1 U22828 ( .A1(n19889), .A2(n19874), .B1(n19873), .B2(n19944), .C1(
        n14972), .C2(n19886), .ZN(P2_U3231) );
  OAI222_X1 U22829 ( .A1(n19889), .A2(n12255), .B1(n19875), .B2(n19944), .C1(
        n19874), .C2(n19886), .ZN(P2_U3232) );
  OAI222_X1 U22830 ( .A1(n19889), .A2(n21110), .B1(n21079), .B2(n19944), .C1(
        n12255), .C2(n19886), .ZN(P2_U3233) );
  OAI222_X1 U22831 ( .A1(n19889), .A2(n16106), .B1(n19876), .B2(n19944), .C1(
        n21110), .C2(n19886), .ZN(P2_U3234) );
  OAI222_X1 U22832 ( .A1(n19889), .A2(n21077), .B1(n19877), .B2(n19944), .C1(
        n16106), .C2(n19886), .ZN(P2_U3235) );
  OAI222_X1 U22833 ( .A1(n19889), .A2(n16095), .B1(n19878), .B2(n19944), .C1(
        n21077), .C2(n19886), .ZN(P2_U3236) );
  OAI222_X1 U22834 ( .A1(n19889), .A2(n19881), .B1(n19879), .B2(n19944), .C1(
        n16095), .C2(n19886), .ZN(P2_U3237) );
  OAI222_X1 U22835 ( .A1(n19886), .A2(n19881), .B1(n19880), .B2(n19944), .C1(
        n19882), .C2(n19889), .ZN(P2_U3238) );
  OAI222_X1 U22836 ( .A1(n19889), .A2(n19884), .B1(n19883), .B2(n19944), .C1(
        n19882), .C2(n19886), .ZN(P2_U3239) );
  OAI222_X1 U22837 ( .A1(n19889), .A2(n12266), .B1(n19885), .B2(n19944), .C1(
        n19884), .C2(n19886), .ZN(P2_U3240) );
  OAI222_X1 U22838 ( .A1(n19889), .A2(n19888), .B1(n19887), .B2(n19944), .C1(
        n12266), .C2(n19886), .ZN(P2_U3241) );
  OAI22_X1 U22839 ( .A1(n19945), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19944), .ZN(n19890) );
  INV_X1 U22840 ( .A(n19890), .ZN(P2_U3585) );
  MUX2_X1 U22841 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n19945), .Z(P2_U3586) );
  OAI22_X1 U22842 ( .A1(n19945), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19944), .ZN(n19891) );
  INV_X1 U22843 ( .A(n19891), .ZN(P2_U3587) );
  OAI22_X1 U22844 ( .A1(n19945), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19944), .ZN(n19892) );
  INV_X1 U22845 ( .A(n19892), .ZN(P2_U3588) );
  OAI21_X1 U22846 ( .B1(n19896), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19894), 
        .ZN(n19893) );
  INV_X1 U22847 ( .A(n19893), .ZN(P2_U3591) );
  OAI21_X1 U22848 ( .B1(n19896), .B2(n19895), .A(n19894), .ZN(P2_U3592) );
  NAND2_X1 U22849 ( .A1(n19897), .A2(n12682), .ZN(n19904) );
  OAI21_X1 U22850 ( .B1(n19899), .B2(n19898), .A(n12682), .ZN(n19901) );
  NAND2_X1 U22851 ( .A1(n19901), .A2(n19900), .ZN(n19912) );
  NAND2_X1 U22852 ( .A1(n19912), .A2(n19902), .ZN(n19903) );
  OAI211_X1 U22853 ( .C1(n19905), .C2(n19576), .A(n19904), .B(n19903), .ZN(
        n19906) );
  INV_X1 U22854 ( .A(n19906), .ZN(n19907) );
  AOI22_X1 U22855 ( .A1(n19931), .A2(n19908), .B1(n19907), .B2(n19932), .ZN(
        P2_U3602) );
  NAND2_X1 U22856 ( .A1(n12882), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19919) );
  OAI21_X1 U22857 ( .B1(n19910), .B2(n19919), .A(n19909), .ZN(n19911) );
  AOI22_X1 U22858 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19913), .B1(n19912), 
        .B2(n19911), .ZN(n19914) );
  AOI22_X1 U22859 ( .A1(n19931), .A2(n19915), .B1(n19914), .B2(n19932), .ZN(
        P2_U3603) );
  INV_X1 U22860 ( .A(n19916), .ZN(n19917) );
  NAND3_X1 U22861 ( .A1(n19920), .A2(n19925), .A3(n19917), .ZN(n19918) );
  OAI21_X1 U22862 ( .B1(n19920), .B2(n19919), .A(n19918), .ZN(n19921) );
  AOI21_X1 U22863 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19922), .A(n19921), 
        .ZN(n19923) );
  AOI22_X1 U22864 ( .A1(n19931), .A2(n19924), .B1(n19923), .B2(n19932), .ZN(
        P2_U3604) );
  INV_X1 U22865 ( .A(n19925), .ZN(n19927) );
  OAI21_X1 U22866 ( .B1(n19928), .B2(n19927), .A(n19926), .ZN(n19929) );
  AOI21_X1 U22867 ( .B1(n19933), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19929), 
        .ZN(n19930) );
  OAI22_X1 U22868 ( .A1(n19933), .A2(n19932), .B1(n19931), .B2(n19930), .ZN(
        P2_U3605) );
  INV_X1 U22869 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19934) );
  AOI22_X1 U22870 ( .A1(n19944), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19934), 
        .B2(n19945), .ZN(P2_U3608) );
  INV_X1 U22871 ( .A(n19935), .ZN(n19936) );
  AOI22_X1 U22872 ( .A1(n19939), .A2(n19938), .B1(n19937), .B2(n19936), .ZN(
        n19940) );
  NAND2_X1 U22873 ( .A1(n19941), .A2(n19940), .ZN(n19943) );
  MUX2_X1 U22874 ( .A(P2_MORE_REG_SCAN_IN), .B(n19943), .S(n19942), .Z(
        P2_U3609) );
  OAI22_X1 U22875 ( .A1(n19945), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19944), .ZN(n19946) );
  INV_X1 U22876 ( .A(n19946), .ZN(P2_U3611) );
  AND2_X1 U22877 ( .A1(n20782), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n19948) );
  INV_X1 U22878 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19947) );
  AOI21_X1 U22879 ( .B1(n19948), .B2(n19947), .A(n20853), .ZN(P1_U2802) );
  OAI21_X1 U22880 ( .B1(n19950), .B2(n19949), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19951) );
  OAI21_X1 U22881 ( .B1(n19952), .B2(n20773), .A(n19951), .ZN(P1_U2803) );
  INV_X2 U22882 ( .A(n20853), .ZN(n20864) );
  NOR2_X1 U22883 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19954) );
  OAI21_X1 U22884 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(n19954), .A(n20864), .ZN(
        n19953) );
  OAI21_X1 U22885 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20864), .A(n19953), 
        .ZN(P1_U2804) );
  AOI21_X1 U22886 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20782), .A(n20853), 
        .ZN(n20844) );
  OAI21_X1 U22887 ( .B1(BS16), .B2(n19954), .A(n20844), .ZN(n20842) );
  OAI21_X1 U22888 ( .B1(n20844), .B2(n20649), .A(n20842), .ZN(P1_U2805) );
  OAI21_X1 U22889 ( .B1(n19957), .B2(n19956), .A(n19955), .ZN(P1_U2806) );
  NOR4_X1 U22890 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19961) );
  NOR4_X1 U22891 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19960) );
  NOR4_X1 U22892 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19959) );
  NOR4_X1 U22893 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19958) );
  NAND4_X1 U22894 ( .A1(n19961), .A2(n19960), .A3(n19959), .A4(n19958), .ZN(
        n19967) );
  NOR4_X1 U22895 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_3__SCAN_IN), .A3(P1_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n19965) );
  AOI211_X1 U22896 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_11__SCAN_IN), .B(
        P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(n19964) );
  NOR4_X1 U22897 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19963) );
  NOR4_X1 U22898 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_7__SCAN_IN), .A3(P1_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n19962) );
  NAND4_X1 U22899 ( .A1(n19965), .A2(n19964), .A3(n19963), .A4(n19962), .ZN(
        n19966) );
  NOR2_X1 U22900 ( .A1(n19967), .A2(n19966), .ZN(n20851) );
  INV_X1 U22901 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19969) );
  NOR3_X1 U22902 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19970) );
  OAI21_X1 U22903 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19970), .A(n20851), .ZN(
        n19968) );
  OAI21_X1 U22904 ( .B1(n20851), .B2(n19969), .A(n19968), .ZN(P1_U2807) );
  INV_X1 U22905 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20843) );
  AOI21_X1 U22906 ( .B1(n14140), .B2(n20843), .A(n19970), .ZN(n19972) );
  INV_X1 U22907 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19971) );
  INV_X1 U22908 ( .A(n20851), .ZN(n20848) );
  AOI22_X1 U22909 ( .A1(n20851), .A2(n19972), .B1(n19971), .B2(n20848), .ZN(
        P1_U2808) );
  INV_X1 U22910 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20801) );
  NAND3_X1 U22911 ( .A1(n20005), .A2(n19983), .A3(n20801), .ZN(n19976) );
  INV_X1 U22912 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19973) );
  OAI21_X1 U22913 ( .B1(n20006), .B2(n19973), .A(n19990), .ZN(n19974) );
  AOI21_X1 U22914 ( .B1(n20021), .B2(P1_EBX_REG_7__SCAN_IN), .A(n19974), .ZN(
        n19975) );
  OAI211_X1 U22915 ( .C1(n19978), .C2(n19977), .A(n19976), .B(n19975), .ZN(
        n19979) );
  AOI21_X1 U22916 ( .B1(n19981), .B2(n19980), .A(n19979), .ZN(n19985) );
  OAI21_X1 U22917 ( .B1(n19983), .B2(n19994), .A(n19982), .ZN(n19999) );
  NAND2_X1 U22918 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19999), .ZN(n19984) );
  OAI211_X1 U22919 ( .C1(n20016), .C2(n19986), .A(n19985), .B(n19984), .ZN(
        P1_U2833) );
  INV_X1 U22920 ( .A(n19987), .ZN(n19988) );
  NAND2_X1 U22921 ( .A1(n20025), .A2(n19988), .ZN(n19992) );
  NAND2_X1 U22922 ( .A1(n20021), .A2(P1_EBX_REG_6__SCAN_IN), .ZN(n19991) );
  NAND2_X1 U22923 ( .A1(n20024), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n19989) );
  AND4_X1 U22924 ( .A1(n19992), .A2(n19991), .A3(n19990), .A4(n19989), .ZN(
        n20002) );
  NAND3_X1 U22925 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n19993) );
  NOR2_X1 U22926 ( .A1(n19994), .A2(n19993), .ZN(n20023) );
  NAND2_X1 U22927 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20023), .ZN(n20013) );
  NOR2_X1 U22928 ( .A1(n20012), .A2(n20013), .ZN(n20000) );
  OAI22_X1 U22929 ( .A1(n19997), .A2(n19996), .B1(n19995), .B2(n20016), .ZN(
        n19998) );
  AOI221_X1 U22930 ( .B1(n20000), .B2(n20928), .C1(n19999), .C2(
        P1_REIP_REG_6__SCAN_IN), .A(n19998), .ZN(n20001) );
  NAND2_X1 U22931 ( .A1(n20002), .A2(n20001), .ZN(P1_U2834) );
  AOI21_X1 U22932 ( .B1(n20005), .B2(n20004), .A(n20003), .ZN(n20034) );
  INV_X1 U22933 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20008) );
  INV_X1 U22934 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20007) );
  OAI22_X1 U22935 ( .A1(n20009), .A2(n20008), .B1(n20007), .B2(n20006), .ZN(
        n20010) );
  AOI211_X1 U22936 ( .C1(n20025), .C2(n9819), .A(n20123), .B(n20010), .ZN(
        n20011) );
  OAI221_X1 U22937 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(n20013), .C1(n20012), 
        .C2(n20034), .A(n20011), .ZN(n20014) );
  AOI21_X1 U22938 ( .B1(n20038), .B2(n20022), .A(n20014), .ZN(n20015) );
  OAI21_X1 U22939 ( .B1(n20017), .B2(n20016), .A(n20015), .ZN(P1_U2835) );
  INV_X1 U22940 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20035) );
  INV_X1 U22941 ( .A(n20018), .ZN(n20020) );
  AOI22_X1 U22942 ( .A1(n20021), .A2(P1_EBX_REG_4__SCAN_IN), .B1(n20020), .B2(
        n20019), .ZN(n20033) );
  NAND2_X1 U22943 ( .A1(n20116), .A2(n20022), .ZN(n20031) );
  AOI22_X1 U22944 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n20024), .B1(
        n20023), .B2(n20035), .ZN(n20030) );
  AOI21_X1 U22945 ( .B1(n20025), .B2(n20124), .A(n20123), .ZN(n20029) );
  INV_X1 U22946 ( .A(n20121), .ZN(n20026) );
  NAND2_X1 U22947 ( .A1(n20027), .A2(n20026), .ZN(n20028) );
  AND4_X1 U22948 ( .A1(n20031), .A2(n20030), .A3(n20029), .A4(n20028), .ZN(
        n20032) );
  OAI211_X1 U22949 ( .C1(n20035), .C2(n20034), .A(n20033), .B(n20032), .ZN(
        P1_U2836) );
  AOI22_X1 U22950 ( .A1(n20038), .A2(n20037), .B1(n20036), .B2(n9819), .ZN(
        n20039) );
  OAI21_X1 U22951 ( .B1(n20040), .B2(n20008), .A(n20039), .ZN(P1_U2867) );
  INV_X1 U22952 ( .A(n20044), .ZN(n20041) );
  AOI22_X1 U22953 ( .A1(n20041), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20075), .ZN(n20042) );
  OAI21_X1 U22954 ( .B1(n20043), .B2(n20047), .A(n20042), .ZN(P1_U2906) );
  INV_X1 U22955 ( .A(P1_UWORD_REG_2__SCAN_IN), .ZN(n21046) );
  INV_X1 U22956 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n20046) );
  INV_X1 U22957 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n20045) );
  OAI22_X1 U22958 ( .A1(n20047), .A2(n20046), .B1(n20045), .B2(n20044), .ZN(
        n20048) );
  INV_X1 U22959 ( .A(n20048), .ZN(n20049) );
  OAI21_X1 U22960 ( .B1(n21046), .B2(n20050), .A(n20049), .ZN(P1_U2918) );
  AOI22_X1 U22961 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20051) );
  OAI21_X1 U22962 ( .B1(n12857), .B2(n20077), .A(n20051), .ZN(P1_U2921) );
  INV_X1 U22963 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20053) );
  AOI22_X1 U22964 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20052) );
  OAI21_X1 U22965 ( .B1(n20053), .B2(n20077), .A(n20052), .ZN(P1_U2922) );
  AOI22_X1 U22966 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20054) );
  OAI21_X1 U22967 ( .B1(n14284), .B2(n20077), .A(n20054), .ZN(P1_U2923) );
  INV_X1 U22968 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20056) );
  AOI22_X1 U22969 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20055) );
  OAI21_X1 U22970 ( .B1(n20056), .B2(n20077), .A(n20055), .ZN(P1_U2924) );
  AOI22_X1 U22971 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20057) );
  OAI21_X1 U22972 ( .B1(n21141), .B2(n20077), .A(n20057), .ZN(P1_U2925) );
  INV_X1 U22973 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20059) );
  AOI22_X1 U22974 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20058) );
  OAI21_X1 U22975 ( .B1(n20059), .B2(n20077), .A(n20058), .ZN(P1_U2926) );
  INV_X1 U22976 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20061) );
  AOI22_X1 U22977 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20060) );
  OAI21_X1 U22978 ( .B1(n20061), .B2(n20077), .A(n20060), .ZN(P1_U2927) );
  INV_X1 U22979 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20964) );
  AOI22_X1 U22980 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n20074), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20075), .ZN(n20062) );
  OAI21_X1 U22981 ( .B1(n20964), .B2(n20077), .A(n20062), .ZN(P1_U2928) );
  AOI22_X1 U22982 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20063) );
  OAI21_X1 U22983 ( .B1(n11310), .B2(n20077), .A(n20063), .ZN(P1_U2929) );
  AOI22_X1 U22984 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20064) );
  OAI21_X1 U22985 ( .B1(n11382), .B2(n20077), .A(n20064), .ZN(P1_U2930) );
  AOI22_X1 U22986 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20065) );
  OAI21_X1 U22987 ( .B1(n13268), .B2(n20077), .A(n20065), .ZN(P1_U2931) );
  AOI22_X1 U22988 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20066) );
  OAI21_X1 U22989 ( .B1(n20067), .B2(n20077), .A(n20066), .ZN(P1_U2932) );
  AOI22_X1 U22990 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20068) );
  OAI21_X1 U22991 ( .B1(n20069), .B2(n20077), .A(n20068), .ZN(P1_U2933) );
  AOI22_X1 U22992 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20070) );
  OAI21_X1 U22993 ( .B1(n20071), .B2(n20077), .A(n20070), .ZN(P1_U2934) );
  AOI22_X1 U22994 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20072) );
  OAI21_X1 U22995 ( .B1(n20073), .B2(n20077), .A(n20072), .ZN(P1_U2935) );
  AOI22_X1 U22996 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20075), .B1(n20074), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20076) );
  OAI21_X1 U22997 ( .B1(n20078), .B2(n20077), .A(n20076), .ZN(P1_U2936) );
  AOI22_X1 U22998 ( .A1(n20104), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20083), .ZN(n20080) );
  NAND2_X1 U22999 ( .A1(n20093), .A2(n20079), .ZN(n20095) );
  NAND2_X1 U23000 ( .A1(n20080), .A2(n20095), .ZN(P1_U2945) );
  AOI22_X1 U23001 ( .A1(n20104), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20083), .ZN(n20082) );
  NAND2_X1 U23002 ( .A1(n20093), .A2(n20081), .ZN(n20097) );
  NAND2_X1 U23003 ( .A1(n20082), .A2(n20097), .ZN(P1_U2946) );
  AOI22_X1 U23004 ( .A1(n20104), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n20083), .ZN(n20085) );
  NAND2_X1 U23005 ( .A1(n20093), .A2(n20084), .ZN(n20099) );
  NAND2_X1 U23006 ( .A1(n20085), .A2(n20099), .ZN(P1_U2947) );
  AOI22_X1 U23007 ( .A1(n20104), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20101), .ZN(n20087) );
  NAND2_X1 U23008 ( .A1(n20093), .A2(n20086), .ZN(n20102) );
  NAND2_X1 U23009 ( .A1(n20087), .A2(n20102), .ZN(P1_U2948) );
  AOI22_X1 U23010 ( .A1(n20104), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20101), .ZN(n20089) );
  NAND2_X1 U23011 ( .A1(n20093), .A2(n20088), .ZN(n20105) );
  NAND2_X1 U23012 ( .A1(n20089), .A2(n20105), .ZN(P1_U2949) );
  AOI22_X1 U23013 ( .A1(n20104), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20101), .ZN(n20091) );
  NAND2_X1 U23014 ( .A1(n20093), .A2(n20090), .ZN(n20107) );
  NAND2_X1 U23015 ( .A1(n20091), .A2(n20107), .ZN(P1_U2950) );
  AOI22_X1 U23016 ( .A1(n20104), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20101), .ZN(n20094) );
  NAND2_X1 U23017 ( .A1(n20093), .A2(n20092), .ZN(n20109) );
  NAND2_X1 U23018 ( .A1(n20094), .A2(n20109), .ZN(P1_U2951) );
  AOI22_X1 U23019 ( .A1(n20104), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20101), .ZN(n20096) );
  NAND2_X1 U23020 ( .A1(n20096), .A2(n20095), .ZN(P1_U2960) );
  AOI22_X1 U23021 ( .A1(n20104), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20101), .ZN(n20098) );
  NAND2_X1 U23022 ( .A1(n20098), .A2(n20097), .ZN(P1_U2961) );
  AOI22_X1 U23023 ( .A1(n20104), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20101), .ZN(n20100) );
  NAND2_X1 U23024 ( .A1(n20100), .A2(n20099), .ZN(P1_U2962) );
  AOI22_X1 U23025 ( .A1(n20104), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20101), .ZN(n20103) );
  NAND2_X1 U23026 ( .A1(n20103), .A2(n20102), .ZN(P1_U2963) );
  AOI22_X1 U23027 ( .A1(n20104), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20101), .ZN(n20106) );
  NAND2_X1 U23028 ( .A1(n20106), .A2(n20105), .ZN(P1_U2964) );
  AOI22_X1 U23029 ( .A1(n20104), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20101), .ZN(n20108) );
  NAND2_X1 U23030 ( .A1(n20108), .A2(n20107), .ZN(P1_U2965) );
  AOI22_X1 U23031 ( .A1(n20104), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20101), .ZN(n20110) );
  NAND2_X1 U23032 ( .A1(n20110), .A2(n20109), .ZN(P1_U2966) );
  AOI22_X1 U23033 ( .A1(n20111), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20123), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20120) );
  OAI21_X1 U23034 ( .B1(n20114), .B2(n20113), .A(n20112), .ZN(n20115) );
  INV_X1 U23035 ( .A(n20115), .ZN(n20125) );
  AOI22_X1 U23036 ( .A1(n20125), .A2(n20118), .B1(n20117), .B2(n20116), .ZN(
        n20119) );
  OAI211_X1 U23037 ( .C1(n20122), .C2(n20121), .A(n20120), .B(n20119), .ZN(
        P1_U2995) );
  AOI22_X1 U23038 ( .A1(n20133), .A2(n20124), .B1(n20123), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n20130) );
  AOI22_X1 U23039 ( .A1(n20125), .A2(n20152), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n20135), .ZN(n20129) );
  OAI211_X1 U23040 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20127), .B(n20126), .ZN(n20128) );
  NAND3_X1 U23041 ( .A1(n20130), .A2(n20129), .A3(n20128), .ZN(P1_U3027) );
  AOI21_X1 U23042 ( .B1(n20133), .B2(n20132), .A(n20131), .ZN(n20138) );
  INV_X1 U23043 ( .A(n20134), .ZN(n20136) );
  AOI22_X1 U23044 ( .A1(n20136), .A2(n20152), .B1(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n20135), .ZN(n20137) );
  OAI211_X1 U23045 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n20139), .A(
        n20138), .B(n20137), .ZN(P1_U3028) );
  NAND2_X1 U23046 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20140), .ZN(
        n20157) );
  AOI21_X1 U23047 ( .B1(n20973), .B2(n20142), .A(n20141), .ZN(n20155) );
  NOR2_X1 U23048 ( .A1(n20143), .A2(n20973), .ZN(n20145) );
  AOI21_X1 U23049 ( .B1(n20145), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n20144), .ZN(n20146) );
  NOR2_X1 U23050 ( .A1(n20147), .A2(n20146), .ZN(n20151) );
  OAI22_X1 U23051 ( .A1(n20149), .A2(n20148), .B1(n13376), .B2(n19990), .ZN(
        n20150) );
  AOI211_X1 U23052 ( .C1(n20153), .C2(n20152), .A(n20151), .B(n20150), .ZN(
        n20154) );
  OAI221_X1 U23053 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20157), .C1(
        n20156), .C2(n20155), .A(n20154), .ZN(P1_U3029) );
  AND2_X1 U23054 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n20158), .ZN(
        P1_U3032) );
  AOI22_X2 U23055 ( .A1(DATAI_16_), .A2(n20207), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20208), .ZN(n20722) );
  INV_X1 U23056 ( .A(n12437), .ZN(n20164) );
  AOI22_X1 U23057 ( .A1(DATAI_24_), .A2(n20207), .B1(BUF1_REG_24__SCAN_IN), 
        .B2(n20208), .ZN(n21205) );
  NAND2_X1 U23058 ( .A1(n20210), .A2(n20166), .ZN(n20647) );
  NOR3_X1 U23059 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20224) );
  NAND2_X1 U23060 ( .A1(n20602), .A2(n20224), .ZN(n20211) );
  OAI22_X1 U23061 ( .A1(n20759), .A2(n21205), .B1(n20647), .B2(n20211), .ZN(
        n20167) );
  INV_X1 U23062 ( .A(n20167), .ZN(n20179) );
  INV_X1 U23063 ( .A(n20490), .ZN(n20168) );
  NOR2_X1 U23064 ( .A1(n20168), .A2(n20443), .ZN(n20175) );
  NAND2_X1 U23065 ( .A1(n20174), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20563) );
  NAND2_X1 U23066 ( .A1(n20230), .A2(n20759), .ZN(n20169) );
  AOI21_X1 U23067 ( .B1(n20169), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20711), 
        .ZN(n20173) );
  OR2_X1 U23068 ( .A1(n12753), .A2(n20170), .ZN(n20250) );
  NAND2_X1 U23069 ( .A1(n20287), .A2(n9741), .ZN(n20176) );
  AOI22_X1 U23070 ( .A1(n20173), .A2(n20176), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20211), .ZN(n20171) );
  NAND2_X1 U23071 ( .A1(n20172), .A2(n20213), .ZN(n20646) );
  INV_X1 U23072 ( .A(n20173), .ZN(n20177) );
  NOR2_X1 U23073 ( .A1(n20174), .A2(n11307), .ZN(n20491) );
  INV_X1 U23074 ( .A(n20491), .ZN(n20444) );
  INV_X1 U23075 ( .A(n20175), .ZN(n20324) );
  AOI22_X1 U23076 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20216), .B1(
        n21195), .B2(n20215), .ZN(n20178) );
  OAI211_X1 U23077 ( .C1(n20722), .C2(n20230), .A(n20179), .B(n20178), .ZN(
        P1_U3033) );
  AOI22_X1 U23078 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20208), .B1(DATAI_17_), 
        .B2(n20207), .ZN(n20728) );
  AOI22_X1 U23079 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20208), .B1(DATAI_25_), 
        .B2(n20207), .ZN(n20616) );
  NAND2_X1 U23080 ( .A1(n20210), .A2(n9729), .ZN(n20661) );
  OAI22_X1 U23081 ( .A1(n20759), .A2(n20616), .B1(n20211), .B2(n20661), .ZN(
        n20180) );
  INV_X1 U23082 ( .A(n20180), .ZN(n20183) );
  NAND2_X1 U23083 ( .A1(n20181), .A2(n20213), .ZN(n20660) );
  AOI22_X1 U23084 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20216), .B1(
        n20723), .B2(n20215), .ZN(n20182) );
  OAI211_X1 U23085 ( .C1(n20728), .C2(n20230), .A(n20183), .B(n20182), .ZN(
        P1_U3034) );
  AOI22_X1 U23086 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20208), .B1(DATAI_26_), 
        .B2(n20207), .ZN(n20734) );
  NAND2_X1 U23087 ( .A1(n20210), .A2(n20184), .ZN(n20666) );
  OAI22_X1 U23088 ( .A1(n20759), .A2(n20734), .B1(n20211), .B2(n20666), .ZN(
        n20185) );
  INV_X1 U23089 ( .A(n20185), .ZN(n20188) );
  NAND2_X1 U23090 ( .A1(n20186), .A2(n20213), .ZN(n20665) );
  AOI22_X1 U23091 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20216), .B1(
        n20729), .B2(n20215), .ZN(n20187) );
  OAI211_X1 U23092 ( .C1(n20671), .C2(n20230), .A(n20188), .B(n20187), .ZN(
        P1_U3035) );
  AOI22_X1 U23093 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20208), .B1(DATAI_27_), 
        .B2(n20207), .ZN(n20740) );
  NAND2_X1 U23094 ( .A1(n20210), .A2(n20189), .ZN(n20673) );
  OAI22_X1 U23095 ( .A1(n20759), .A2(n20740), .B1(n20211), .B2(n20673), .ZN(
        n20190) );
  INV_X1 U23096 ( .A(n20190), .ZN(n20193) );
  NAND2_X1 U23097 ( .A1(n20191), .A2(n20213), .ZN(n20672) );
  AOI22_X1 U23098 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20216), .B1(
        n20735), .B2(n20215), .ZN(n20192) );
  OAI211_X1 U23099 ( .C1(n20678), .C2(n20230), .A(n20193), .B(n20192), .ZN(
        P1_U3036) );
  AOI22_X2 U23100 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20208), .B1(DATAI_20_), 
        .B2(n20207), .ZN(n20746) );
  AOI22_X1 U23101 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20208), .B1(DATAI_28_), 
        .B2(n20207), .ZN(n20624) );
  NAND2_X1 U23102 ( .A1(n20210), .A2(n11204), .ZN(n20680) );
  OAI22_X1 U23103 ( .A1(n20759), .A2(n20624), .B1(n20211), .B2(n20680), .ZN(
        n20194) );
  INV_X1 U23104 ( .A(n20194), .ZN(n20197) );
  NAND2_X1 U23105 ( .A1(n20195), .A2(n20213), .ZN(n20679) );
  AOI22_X1 U23106 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20216), .B1(
        n20741), .B2(n20215), .ZN(n20196) );
  OAI211_X1 U23107 ( .C1(n20746), .C2(n20230), .A(n20197), .B(n20196), .ZN(
        P1_U3037) );
  AOI22_X1 U23108 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20208), .B1(DATAI_29_), 
        .B2(n20207), .ZN(n20752) );
  NAND2_X1 U23109 ( .A1(n20210), .A2(n20198), .ZN(n20685) );
  OAI22_X1 U23110 ( .A1(n20759), .A2(n20752), .B1(n20211), .B2(n20685), .ZN(
        n20199) );
  INV_X1 U23111 ( .A(n20199), .ZN(n20202) );
  NAND2_X1 U23112 ( .A1(n20200), .A2(n20213), .ZN(n20684) );
  AOI22_X1 U23113 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20216), .B1(
        n20747), .B2(n20215), .ZN(n20201) );
  OAI211_X1 U23114 ( .C1(n20690), .C2(n20230), .A(n20202), .B(n20201), .ZN(
        P1_U3038) );
  AOI22_X1 U23115 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20208), .B1(DATAI_30_), 
        .B2(n20207), .ZN(n20630) );
  NAND2_X1 U23116 ( .A1(n20210), .A2(n11155), .ZN(n20692) );
  OAI22_X1 U23117 ( .A1(n20759), .A2(n20630), .B1(n20211), .B2(n20692), .ZN(
        n20203) );
  INV_X1 U23118 ( .A(n20203), .ZN(n20206) );
  NAND2_X1 U23119 ( .A1(n20204), .A2(n20213), .ZN(n20691) );
  AOI22_X1 U23120 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20216), .B1(
        n20753), .B2(n20215), .ZN(n20205) );
  OAI211_X1 U23121 ( .C1(n20760), .C2(n20230), .A(n20206), .B(n20205), .ZN(
        P1_U3039) );
  AOI22_X1 U23122 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20208), .B1(DATAI_31_), 
        .B2(n20207), .ZN(n20771) );
  NAND2_X1 U23123 ( .A1(n20210), .A2(n20209), .ZN(n20699) );
  OAI22_X1 U23124 ( .A1(n20759), .A2(n20771), .B1(n20211), .B2(n20699), .ZN(
        n20212) );
  INV_X1 U23125 ( .A(n20212), .ZN(n20218) );
  NAND2_X1 U23126 ( .A1(n20214), .A2(n20213), .ZN(n20697) );
  AOI22_X1 U23127 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20216), .B1(
        n20762), .B2(n20215), .ZN(n20217) );
  OAI211_X1 U23128 ( .C1(n20706), .C2(n20230), .A(n20218), .B(n20217), .ZN(
        P1_U3040) );
  INV_X1 U23129 ( .A(n20219), .ZN(n20603) );
  INV_X1 U23130 ( .A(n20224), .ZN(n20220) );
  NOR2_X1 U23131 ( .A1(n20602), .A2(n20220), .ZN(n20241) );
  AOI21_X1 U23132 ( .B1(n20287), .B2(n20603), .A(n20241), .ZN(n20221) );
  OAI22_X1 U23133 ( .A1(n20221), .A2(n20711), .B1(n20220), .B2(n11307), .ZN(
        n20242) );
  INV_X1 U23134 ( .A(n20647), .ZN(n21198) );
  AOI22_X1 U23135 ( .A1(n21195), .A2(n20242), .B1(n21198), .B2(n20241), .ZN(
        n20226) );
  INV_X1 U23136 ( .A(n20289), .ZN(n20222) );
  OAI21_X1 U23137 ( .B1(n20222), .B2(n20471), .A(n20221), .ZN(n20223) );
  OAI221_X1 U23138 ( .B1(n20717), .B2(n20224), .C1(n20711), .C2(n20223), .A(
        n20716), .ZN(n20244) );
  INV_X1 U23139 ( .A(n21205), .ZN(n20719) );
  AOI22_X1 U23140 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20244), .B1(
        n20243), .B2(n20719), .ZN(n20225) );
  OAI211_X1 U23141 ( .C1(n20722), .C2(n20276), .A(n20226), .B(n20225), .ZN(
        P1_U3041) );
  INV_X1 U23142 ( .A(n20661), .ZN(n20724) );
  AOI22_X1 U23143 ( .A1(n20723), .A2(n20242), .B1(n20724), .B2(n20241), .ZN(
        n20229) );
  INV_X1 U23144 ( .A(n20276), .ZN(n20227) );
  INV_X1 U23145 ( .A(n20728), .ZN(n20613) );
  AOI22_X1 U23146 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20244), .B1(
        n20227), .B2(n20613), .ZN(n20228) );
  OAI211_X1 U23147 ( .C1(n20616), .C2(n20230), .A(n20229), .B(n20228), .ZN(
        P1_U3042) );
  INV_X1 U23148 ( .A(n20666), .ZN(n20730) );
  AOI22_X1 U23149 ( .A1(n20729), .A2(n20242), .B1(n20730), .B2(n20241), .ZN(
        n20232) );
  INV_X1 U23150 ( .A(n20734), .ZN(n20668) );
  AOI22_X1 U23151 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20244), .B1(
        n20243), .B2(n20668), .ZN(n20231) );
  OAI211_X1 U23152 ( .C1(n20671), .C2(n20276), .A(n20232), .B(n20231), .ZN(
        P1_U3043) );
  INV_X1 U23153 ( .A(n20673), .ZN(n20736) );
  AOI22_X1 U23154 ( .A1(n20735), .A2(n20242), .B1(n20736), .B2(n20241), .ZN(
        n20234) );
  INV_X1 U23155 ( .A(n20740), .ZN(n20675) );
  AOI22_X1 U23156 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20244), .B1(
        n20243), .B2(n20675), .ZN(n20233) );
  OAI211_X1 U23157 ( .C1(n20678), .C2(n20276), .A(n20234), .B(n20233), .ZN(
        P1_U3044) );
  INV_X1 U23158 ( .A(n20680), .ZN(n20742) );
  AOI22_X1 U23159 ( .A1(n20741), .A2(n20242), .B1(n20742), .B2(n20241), .ZN(
        n20236) );
  INV_X1 U23160 ( .A(n20624), .ZN(n20743) );
  AOI22_X1 U23161 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20244), .B1(
        n20243), .B2(n20743), .ZN(n20235) );
  OAI211_X1 U23162 ( .C1(n20746), .C2(n20276), .A(n20236), .B(n20235), .ZN(
        P1_U3045) );
  INV_X1 U23163 ( .A(n20685), .ZN(n20748) );
  AOI22_X1 U23164 ( .A1(n20747), .A2(n20242), .B1(n20748), .B2(n20241), .ZN(
        n20238) );
  INV_X1 U23165 ( .A(n20752), .ZN(n20687) );
  AOI22_X1 U23166 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20244), .B1(
        n20243), .B2(n20687), .ZN(n20237) );
  OAI211_X1 U23167 ( .C1(n20690), .C2(n20276), .A(n20238), .B(n20237), .ZN(
        P1_U3046) );
  INV_X1 U23168 ( .A(n20692), .ZN(n20754) );
  AOI22_X1 U23169 ( .A1(n20753), .A2(n20242), .B1(n20754), .B2(n20241), .ZN(
        n20240) );
  INV_X1 U23170 ( .A(n20630), .ZN(n20755) );
  AOI22_X1 U23171 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20244), .B1(
        n20243), .B2(n20755), .ZN(n20239) );
  OAI211_X1 U23172 ( .C1(n20760), .C2(n20276), .A(n20240), .B(n20239), .ZN(
        P1_U3047) );
  INV_X1 U23173 ( .A(n20699), .ZN(n20764) );
  AOI22_X1 U23174 ( .A1(n20762), .A2(n20242), .B1(n20764), .B2(n20241), .ZN(
        n20246) );
  INV_X1 U23175 ( .A(n20771), .ZN(n20701) );
  AOI22_X1 U23176 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20244), .B1(
        n20243), .B2(n20701), .ZN(n20245) );
  OAI211_X1 U23177 ( .C1(n20706), .C2(n20276), .A(n20246), .B(n20245), .ZN(
        P1_U3048) );
  NAND3_X1 U23178 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20565), .A3(
        n20566), .ZN(n20292) );
  OR2_X1 U23179 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20292), .ZN(
        n20275) );
  OAI22_X1 U23180 ( .A1(n20276), .A2(n21205), .B1(n20647), .B2(n20275), .ZN(
        n20248) );
  INV_X1 U23181 ( .A(n20248), .ZN(n20256) );
  NAND3_X1 U23182 ( .A1(n20316), .A2(n20276), .A3(n20717), .ZN(n20249) );
  NAND2_X1 U23183 ( .A1(n20717), .A2(n20649), .ZN(n20560) );
  NAND2_X1 U23184 ( .A1(n20249), .A2(n20560), .ZN(n20252) );
  OR2_X1 U23185 ( .A1(n20250), .A2(n9741), .ZN(n20253) );
  AOI22_X1 U23186 ( .A1(n20252), .A2(n20253), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20275), .ZN(n20251) );
  OR2_X1 U23187 ( .A1(n20490), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20383) );
  NAND2_X1 U23188 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20383), .ZN(n20380) );
  NAND3_X1 U23189 ( .A1(n20497), .A2(n20251), .A3(n20380), .ZN(n20279) );
  INV_X1 U23190 ( .A(n20252), .ZN(n20254) );
  AOI22_X1 U23191 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20279), .B1(
        n21195), .B2(n20278), .ZN(n20255) );
  OAI211_X1 U23192 ( .C1(n20722), .C2(n20316), .A(n20256), .B(n20255), .ZN(
        P1_U3049) );
  OAI22_X1 U23193 ( .A1(n20276), .A2(n20616), .B1(n20661), .B2(n20275), .ZN(
        n20257) );
  INV_X1 U23194 ( .A(n20257), .ZN(n20259) );
  AOI22_X1 U23195 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20279), .B1(
        n20723), .B2(n20278), .ZN(n20258) );
  OAI211_X1 U23196 ( .C1(n20728), .C2(n20316), .A(n20259), .B(n20258), .ZN(
        P1_U3050) );
  OAI22_X1 U23197 ( .A1(n20276), .A2(n20734), .B1(n20666), .B2(n20275), .ZN(
        n20260) );
  INV_X1 U23198 ( .A(n20260), .ZN(n20262) );
  AOI22_X1 U23199 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20279), .B1(
        n20729), .B2(n20278), .ZN(n20261) );
  OAI211_X1 U23200 ( .C1(n20671), .C2(n20316), .A(n20262), .B(n20261), .ZN(
        P1_U3051) );
  OAI22_X1 U23201 ( .A1(n20316), .A2(n20678), .B1(n20673), .B2(n20275), .ZN(
        n20263) );
  INV_X1 U23202 ( .A(n20263), .ZN(n20265) );
  AOI22_X1 U23203 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20279), .B1(
        n20735), .B2(n20278), .ZN(n20264) );
  OAI211_X1 U23204 ( .C1(n20740), .C2(n20276), .A(n20265), .B(n20264), .ZN(
        P1_U3052) );
  OAI22_X1 U23205 ( .A1(n20316), .A2(n20746), .B1(n20680), .B2(n20275), .ZN(
        n20266) );
  INV_X1 U23206 ( .A(n20266), .ZN(n20268) );
  AOI22_X1 U23207 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20279), .B1(
        n20741), .B2(n20278), .ZN(n20267) );
  OAI211_X1 U23208 ( .C1(n20624), .C2(n20276), .A(n20268), .B(n20267), .ZN(
        P1_U3053) );
  OAI22_X1 U23209 ( .A1(n20316), .A2(n20690), .B1(n20685), .B2(n20275), .ZN(
        n20269) );
  INV_X1 U23210 ( .A(n20269), .ZN(n20271) );
  AOI22_X1 U23211 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20279), .B1(
        n20747), .B2(n20278), .ZN(n20270) );
  OAI211_X1 U23212 ( .C1(n20752), .C2(n20276), .A(n20271), .B(n20270), .ZN(
        P1_U3054) );
  OAI22_X1 U23213 ( .A1(n20276), .A2(n20630), .B1(n20692), .B2(n20275), .ZN(
        n20272) );
  INV_X1 U23214 ( .A(n20272), .ZN(n20274) );
  AOI22_X1 U23215 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20279), .B1(
        n20753), .B2(n20278), .ZN(n20273) );
  OAI211_X1 U23216 ( .C1(n20760), .C2(n20316), .A(n20274), .B(n20273), .ZN(
        P1_U3055) );
  OAI22_X1 U23217 ( .A1(n20276), .A2(n20771), .B1(n20699), .B2(n20275), .ZN(
        n20277) );
  INV_X1 U23218 ( .A(n20277), .ZN(n20281) );
  AOI22_X1 U23219 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20279), .B1(
        n20762), .B2(n20278), .ZN(n20280) );
  OAI211_X1 U23220 ( .C1(n20706), .C2(n20316), .A(n20281), .B(n20280), .ZN(
        P1_U3056) );
  INV_X1 U23221 ( .A(n20528), .ZN(n20282) );
  NAND2_X1 U23222 ( .A1(n20282), .A2(n20565), .ZN(n20315) );
  OAI22_X1 U23223 ( .A1(n20316), .A2(n21205), .B1(n20647), .B2(n20315), .ZN(
        n20283) );
  INV_X1 U23224 ( .A(n20283), .ZN(n20296) );
  AND2_X1 U23225 ( .A1(n20285), .A2(n20284), .ZN(n20708) );
  INV_X1 U23226 ( .A(n20315), .ZN(n20286) );
  AOI21_X1 U23227 ( .B1(n20287), .B2(n20708), .A(n20286), .ZN(n20294) );
  AOI21_X1 U23228 ( .B1(n20289), .B2(n20288), .A(n20711), .ZN(n20291) );
  AOI22_X1 U23229 ( .A1(n20294), .A2(n20291), .B1(n20711), .B2(n20292), .ZN(
        n20290) );
  NAND2_X1 U23230 ( .A1(n20716), .A2(n20290), .ZN(n20319) );
  INV_X1 U23231 ( .A(n20291), .ZN(n20293) );
  OAI22_X1 U23232 ( .A1(n20294), .A2(n20293), .B1(n11307), .B2(n20292), .ZN(
        n20318) );
  AOI22_X1 U23233 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20319), .B1(
        n21195), .B2(n20318), .ZN(n20295) );
  OAI211_X1 U23234 ( .C1(n20722), .C2(n20329), .A(n20296), .B(n20295), .ZN(
        P1_U3057) );
  OAI22_X1 U23235 ( .A1(n20316), .A2(n20616), .B1(n20661), .B2(n20315), .ZN(
        n20297) );
  INV_X1 U23236 ( .A(n20297), .ZN(n20299) );
  AOI22_X1 U23237 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20319), .B1(
        n20723), .B2(n20318), .ZN(n20298) );
  OAI211_X1 U23238 ( .C1(n20728), .C2(n20329), .A(n20299), .B(n20298), .ZN(
        P1_U3058) );
  OAI22_X1 U23239 ( .A1(n20329), .A2(n20671), .B1(n20666), .B2(n20315), .ZN(
        n20300) );
  INV_X1 U23240 ( .A(n20300), .ZN(n20302) );
  AOI22_X1 U23241 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20319), .B1(
        n20729), .B2(n20318), .ZN(n20301) );
  OAI211_X1 U23242 ( .C1(n20734), .C2(n20316), .A(n20302), .B(n20301), .ZN(
        P1_U3059) );
  OAI22_X1 U23243 ( .A1(n20316), .A2(n20740), .B1(n20673), .B2(n20315), .ZN(
        n20303) );
  INV_X1 U23244 ( .A(n20303), .ZN(n20305) );
  AOI22_X1 U23245 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20319), .B1(
        n20735), .B2(n20318), .ZN(n20304) );
  OAI211_X1 U23246 ( .C1(n20678), .C2(n20329), .A(n20305), .B(n20304), .ZN(
        P1_U3060) );
  OAI22_X1 U23247 ( .A1(n20316), .A2(n20624), .B1(n20680), .B2(n20315), .ZN(
        n20306) );
  INV_X1 U23248 ( .A(n20306), .ZN(n20308) );
  AOI22_X1 U23249 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20319), .B1(
        n20741), .B2(n20318), .ZN(n20307) );
  OAI211_X1 U23250 ( .C1(n20746), .C2(n20329), .A(n20308), .B(n20307), .ZN(
        P1_U3061) );
  OAI22_X1 U23251 ( .A1(n20316), .A2(n20752), .B1(n20685), .B2(n20315), .ZN(
        n20309) );
  INV_X1 U23252 ( .A(n20309), .ZN(n20311) );
  AOI22_X1 U23253 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20319), .B1(
        n20747), .B2(n20318), .ZN(n20310) );
  OAI211_X1 U23254 ( .C1(n20690), .C2(n20329), .A(n20311), .B(n20310), .ZN(
        P1_U3062) );
  OAI22_X1 U23255 ( .A1(n20316), .A2(n20630), .B1(n20692), .B2(n20315), .ZN(
        n20312) );
  INV_X1 U23256 ( .A(n20312), .ZN(n20314) );
  AOI22_X1 U23257 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20319), .B1(
        n20753), .B2(n20318), .ZN(n20313) );
  OAI211_X1 U23258 ( .C1(n20760), .C2(n20329), .A(n20314), .B(n20313), .ZN(
        P1_U3063) );
  OAI22_X1 U23259 ( .A1(n20316), .A2(n20771), .B1(n20699), .B2(n20315), .ZN(
        n20317) );
  INV_X1 U23260 ( .A(n20317), .ZN(n20321) );
  AOI22_X1 U23261 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20319), .B1(
        n20762), .B2(n20318), .ZN(n20320) );
  OAI211_X1 U23262 ( .C1(n20706), .C2(n20329), .A(n20321), .B(n20320), .ZN(
        P1_U3064) );
  NOR3_X1 U23263 ( .A1(n20566), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20355) );
  INV_X1 U23264 ( .A(n20355), .ZN(n20351) );
  NOR2_X1 U23265 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20351), .ZN(
        n20345) );
  NOR2_X1 U23266 ( .A1(n13145), .A2(n20322), .ZN(n20414) );
  NAND3_X1 U23267 ( .A1(n20414), .A2(n20717), .A3(n9741), .ZN(n20323) );
  OAI21_X1 U23268 ( .B1(n20324), .B2(n20563), .A(n20323), .ZN(n20344) );
  AOI22_X1 U23269 ( .A1(n21198), .A2(n20345), .B1(n21195), .B2(n20344), .ZN(
        n20331) );
  AOI21_X1 U23270 ( .B1(n20329), .B2(n20377), .A(n20649), .ZN(n20325) );
  AOI21_X1 U23271 ( .B1(n20414), .B2(n9741), .A(n20325), .ZN(n20326) );
  NOR2_X1 U23272 ( .A1(n20326), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20328) );
  NOR2_X1 U23273 ( .A1(n20491), .A2(n20327), .ZN(n20655) );
  AOI22_X1 U23274 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20347), .B1(
        n20346), .B2(n20719), .ZN(n20330) );
  OAI211_X1 U23275 ( .C1(n20722), .C2(n20377), .A(n20331), .B(n20330), .ZN(
        P1_U3065) );
  AOI22_X1 U23276 ( .A1(n20724), .A2(n20345), .B1(n20723), .B2(n20344), .ZN(
        n20333) );
  INV_X1 U23277 ( .A(n20616), .ZN(n20725) );
  AOI22_X1 U23278 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20347), .B1(
        n20346), .B2(n20725), .ZN(n20332) );
  OAI211_X1 U23279 ( .C1(n20728), .C2(n20377), .A(n20333), .B(n20332), .ZN(
        P1_U3066) );
  AOI22_X1 U23280 ( .A1(n20730), .A2(n20345), .B1(n20729), .B2(n20344), .ZN(
        n20335) );
  AOI22_X1 U23281 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20347), .B1(
        n20346), .B2(n20668), .ZN(n20334) );
  OAI211_X1 U23282 ( .C1(n20671), .C2(n20377), .A(n20335), .B(n20334), .ZN(
        P1_U3067) );
  AOI22_X1 U23283 ( .A1(n20736), .A2(n20345), .B1(n20735), .B2(n20344), .ZN(
        n20337) );
  AOI22_X1 U23284 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20347), .B1(
        n20346), .B2(n20675), .ZN(n20336) );
  OAI211_X1 U23285 ( .C1(n20678), .C2(n20377), .A(n20337), .B(n20336), .ZN(
        P1_U3068) );
  AOI22_X1 U23286 ( .A1(n20742), .A2(n20345), .B1(n20741), .B2(n20344), .ZN(
        n20339) );
  AOI22_X1 U23287 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20347), .B1(
        n20346), .B2(n20743), .ZN(n20338) );
  OAI211_X1 U23288 ( .C1(n20746), .C2(n20377), .A(n20339), .B(n20338), .ZN(
        P1_U3069) );
  AOI22_X1 U23289 ( .A1(n20748), .A2(n20345), .B1(n20747), .B2(n20344), .ZN(
        n20341) );
  AOI22_X1 U23290 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20347), .B1(
        n20346), .B2(n20687), .ZN(n20340) );
  OAI211_X1 U23291 ( .C1(n20690), .C2(n20377), .A(n20341), .B(n20340), .ZN(
        P1_U3070) );
  AOI22_X1 U23292 ( .A1(n20754), .A2(n20345), .B1(n20753), .B2(n20344), .ZN(
        n20343) );
  AOI22_X1 U23293 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20347), .B1(
        n20346), .B2(n20755), .ZN(n20342) );
  OAI211_X1 U23294 ( .C1(n20760), .C2(n20377), .A(n20343), .B(n20342), .ZN(
        P1_U3071) );
  AOI22_X1 U23295 ( .A1(n20764), .A2(n20345), .B1(n20762), .B2(n20344), .ZN(
        n20349) );
  AOI22_X1 U23296 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20347), .B1(
        n20346), .B2(n20701), .ZN(n20348) );
  OAI211_X1 U23297 ( .C1(n20706), .C2(n20377), .A(n20349), .B(n20348), .ZN(
        P1_U3072) );
  NOR2_X1 U23298 ( .A1(n20602), .A2(n20351), .ZN(n20372) );
  AOI21_X1 U23299 ( .B1(n20414), .B2(n20603), .A(n20372), .ZN(n20352) );
  OAI22_X1 U23300 ( .A1(n20352), .A2(n20711), .B1(n20351), .B2(n11307), .ZN(
        n20371) );
  AOI22_X1 U23301 ( .A1(n21198), .A2(n20372), .B1(n21195), .B2(n20371), .ZN(
        n20358) );
  INV_X1 U23302 ( .A(n20420), .ZN(n20353) );
  OAI21_X1 U23303 ( .B1(n20353), .B2(n20471), .A(n20352), .ZN(n20354) );
  OAI221_X1 U23304 ( .B1(n20717), .B2(n20355), .C1(n20711), .C2(n20354), .A(
        n20716), .ZN(n20374) );
  INV_X1 U23305 ( .A(n20377), .ZN(n20356) );
  AOI22_X1 U23306 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20374), .B1(
        n20356), .B2(n20719), .ZN(n20357) );
  OAI211_X1 U23307 ( .C1(n20722), .C2(n20412), .A(n20358), .B(n20357), .ZN(
        P1_U3073) );
  AOI22_X1 U23308 ( .A1(n20724), .A2(n20372), .B1(n20723), .B2(n20371), .ZN(
        n20360) );
  AOI22_X1 U23309 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20374), .B1(
        n20373), .B2(n20613), .ZN(n20359) );
  OAI211_X1 U23310 ( .C1(n20616), .C2(n20377), .A(n20360), .B(n20359), .ZN(
        P1_U3074) );
  AOI22_X1 U23311 ( .A1(n20730), .A2(n20372), .B1(n20729), .B2(n20371), .ZN(
        n20362) );
  INV_X1 U23312 ( .A(n20671), .ZN(n20731) );
  AOI22_X1 U23313 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20374), .B1(
        n20373), .B2(n20731), .ZN(n20361) );
  OAI211_X1 U23314 ( .C1(n20734), .C2(n20377), .A(n20362), .B(n20361), .ZN(
        P1_U3075) );
  AOI22_X1 U23315 ( .A1(n20736), .A2(n20372), .B1(n20735), .B2(n20371), .ZN(
        n20364) );
  INV_X1 U23316 ( .A(n20678), .ZN(n20737) );
  AOI22_X1 U23317 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20374), .B1(
        n20373), .B2(n20737), .ZN(n20363) );
  OAI211_X1 U23318 ( .C1(n20740), .C2(n20377), .A(n20364), .B(n20363), .ZN(
        P1_U3076) );
  AOI22_X1 U23319 ( .A1(n20742), .A2(n20372), .B1(n20741), .B2(n20371), .ZN(
        n20366) );
  INV_X1 U23320 ( .A(n20746), .ZN(n20621) );
  AOI22_X1 U23321 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20374), .B1(
        n20373), .B2(n20621), .ZN(n20365) );
  OAI211_X1 U23322 ( .C1(n20624), .C2(n20377), .A(n20366), .B(n20365), .ZN(
        P1_U3077) );
  AOI22_X1 U23323 ( .A1(n20748), .A2(n20372), .B1(n20747), .B2(n20371), .ZN(
        n20368) );
  INV_X1 U23324 ( .A(n20690), .ZN(n20749) );
  AOI22_X1 U23325 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20374), .B1(
        n20373), .B2(n20749), .ZN(n20367) );
  OAI211_X1 U23326 ( .C1(n20752), .C2(n20377), .A(n20368), .B(n20367), .ZN(
        P1_U3078) );
  AOI22_X1 U23327 ( .A1(n20754), .A2(n20372), .B1(n20753), .B2(n20371), .ZN(
        n20370) );
  INV_X1 U23328 ( .A(n20760), .ZN(n20627) );
  AOI22_X1 U23329 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20374), .B1(
        n20373), .B2(n20627), .ZN(n20369) );
  OAI211_X1 U23330 ( .C1(n20630), .C2(n20377), .A(n20370), .B(n20369), .ZN(
        P1_U3079) );
  AOI22_X1 U23331 ( .A1(n20764), .A2(n20372), .B1(n20762), .B2(n20371), .ZN(
        n20376) );
  INV_X1 U23332 ( .A(n20706), .ZN(n20765) );
  AOI22_X1 U23333 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20374), .B1(
        n20373), .B2(n20765), .ZN(n20375) );
  OAI211_X1 U23334 ( .C1(n20771), .C2(n20377), .A(n20376), .B(n20375), .ZN(
        P1_U3080) );
  NAND2_X1 U23335 ( .A1(n20602), .A2(n11227), .ZN(n20406) );
  OAI22_X1 U23336 ( .A1(n20412), .A2(n21205), .B1(n20647), .B2(n20406), .ZN(
        n20378) );
  INV_X1 U23337 ( .A(n20378), .ZN(n20387) );
  NAND2_X1 U23338 ( .A1(n20435), .A2(n20412), .ZN(n20379) );
  AOI21_X1 U23339 ( .B1(n20379), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20711), 
        .ZN(n20382) );
  NAND2_X1 U23340 ( .A1(n20414), .A2(n20652), .ZN(n20384) );
  AOI22_X1 U23341 ( .A1(n20382), .A2(n20384), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20406), .ZN(n20381) );
  NAND3_X1 U23342 ( .A1(n20655), .A2(n20381), .A3(n20380), .ZN(n20409) );
  INV_X1 U23343 ( .A(n20382), .ZN(n20385) );
  AOI22_X1 U23344 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20409), .B1(
        n21195), .B2(n20408), .ZN(n20386) );
  OAI211_X1 U23345 ( .C1(n20722), .C2(n20435), .A(n20387), .B(n20386), .ZN(
        P1_U3081) );
  OAI22_X1 U23346 ( .A1(n20435), .A2(n20728), .B1(n20661), .B2(n20406), .ZN(
        n20388) );
  INV_X1 U23347 ( .A(n20388), .ZN(n20390) );
  AOI22_X1 U23348 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20409), .B1(
        n20723), .B2(n20408), .ZN(n20389) );
  OAI211_X1 U23349 ( .C1(n20616), .C2(n20412), .A(n20390), .B(n20389), .ZN(
        P1_U3082) );
  OAI22_X1 U23350 ( .A1(n20435), .A2(n20671), .B1(n20666), .B2(n20406), .ZN(
        n20391) );
  INV_X1 U23351 ( .A(n20391), .ZN(n20393) );
  AOI22_X1 U23352 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20409), .B1(
        n20729), .B2(n20408), .ZN(n20392) );
  OAI211_X1 U23353 ( .C1(n20734), .C2(n20412), .A(n20393), .B(n20392), .ZN(
        P1_U3083) );
  OAI22_X1 U23354 ( .A1(n20435), .A2(n20678), .B1(n20673), .B2(n20406), .ZN(
        n20394) );
  INV_X1 U23355 ( .A(n20394), .ZN(n20396) );
  AOI22_X1 U23356 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20409), .B1(
        n20735), .B2(n20408), .ZN(n20395) );
  OAI211_X1 U23357 ( .C1(n20740), .C2(n20412), .A(n20396), .B(n20395), .ZN(
        P1_U3084) );
  OAI22_X1 U23358 ( .A1(n20435), .A2(n20746), .B1(n20680), .B2(n20406), .ZN(
        n20397) );
  INV_X1 U23359 ( .A(n20397), .ZN(n20399) );
  AOI22_X1 U23360 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20409), .B1(
        n20741), .B2(n20408), .ZN(n20398) );
  OAI211_X1 U23361 ( .C1(n20624), .C2(n20412), .A(n20399), .B(n20398), .ZN(
        P1_U3085) );
  OAI22_X1 U23362 ( .A1(n20435), .A2(n20690), .B1(n20685), .B2(n20406), .ZN(
        n20400) );
  INV_X1 U23363 ( .A(n20400), .ZN(n20402) );
  AOI22_X1 U23364 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20409), .B1(
        n20747), .B2(n20408), .ZN(n20401) );
  OAI211_X1 U23365 ( .C1(n20752), .C2(n20412), .A(n20402), .B(n20401), .ZN(
        P1_U3086) );
  OAI22_X1 U23366 ( .A1(n20412), .A2(n20630), .B1(n20692), .B2(n20406), .ZN(
        n20403) );
  INV_X1 U23367 ( .A(n20403), .ZN(n20405) );
  AOI22_X1 U23368 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20409), .B1(
        n20753), .B2(n20408), .ZN(n20404) );
  OAI211_X1 U23369 ( .C1(n20760), .C2(n20435), .A(n20405), .B(n20404), .ZN(
        P1_U3087) );
  OAI22_X1 U23370 ( .A1(n20435), .A2(n20706), .B1(n20699), .B2(n20406), .ZN(
        n20407) );
  INV_X1 U23371 ( .A(n20407), .ZN(n20411) );
  AOI22_X1 U23372 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20409), .B1(
        n20762), .B2(n20408), .ZN(n20410) );
  OAI211_X1 U23373 ( .C1(n20771), .C2(n20412), .A(n20411), .B(n20410), .ZN(
        P1_U3088) );
  INV_X1 U23374 ( .A(n20413), .ZN(n20437) );
  AOI21_X1 U23375 ( .B1(n20414), .B2(n20708), .A(n20437), .ZN(n20416) );
  OAI22_X1 U23376 ( .A1(n20416), .A2(n20711), .B1(n20415), .B2(n11307), .ZN(
        n20436) );
  AOI22_X1 U23377 ( .A1(n21198), .A2(n20437), .B1(n21195), .B2(n20436), .ZN(
        n20422) );
  NAND2_X1 U23378 ( .A1(n20417), .A2(n20416), .ZN(n20418) );
  OAI221_X1 U23379 ( .B1(n20717), .B2(n11227), .C1(n20711), .C2(n20418), .A(
        n20716), .ZN(n20439) );
  INV_X1 U23380 ( .A(n20722), .ZN(n21199) );
  AOI22_X1 U23381 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20439), .B1(
        n20465), .B2(n21199), .ZN(n20421) );
  OAI211_X1 U23382 ( .C1(n21205), .C2(n20435), .A(n20422), .B(n20421), .ZN(
        P1_U3089) );
  AOI22_X1 U23383 ( .A1(n20724), .A2(n20437), .B1(n20723), .B2(n20436), .ZN(
        n20424) );
  INV_X1 U23384 ( .A(n20435), .ZN(n20438) );
  AOI22_X1 U23385 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20439), .B1(
        n20438), .B2(n20725), .ZN(n20423) );
  OAI211_X1 U23386 ( .C1(n20728), .C2(n20442), .A(n20424), .B(n20423), .ZN(
        P1_U3090) );
  AOI22_X1 U23387 ( .A1(n20730), .A2(n20437), .B1(n20729), .B2(n20436), .ZN(
        n20426) );
  AOI22_X1 U23388 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20439), .B1(
        n20438), .B2(n20668), .ZN(n20425) );
  OAI211_X1 U23389 ( .C1(n20671), .C2(n20442), .A(n20426), .B(n20425), .ZN(
        P1_U3091) );
  AOI22_X1 U23390 ( .A1(n20736), .A2(n20437), .B1(n20735), .B2(n20436), .ZN(
        n20428) );
  AOI22_X1 U23391 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20439), .B1(
        n20438), .B2(n20675), .ZN(n20427) );
  OAI211_X1 U23392 ( .C1(n20678), .C2(n20442), .A(n20428), .B(n20427), .ZN(
        P1_U3092) );
  AOI22_X1 U23393 ( .A1(n20742), .A2(n20437), .B1(n20741), .B2(n20436), .ZN(
        n20430) );
  AOI22_X1 U23394 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20439), .B1(
        n20438), .B2(n20743), .ZN(n20429) );
  OAI211_X1 U23395 ( .C1(n20746), .C2(n20442), .A(n20430), .B(n20429), .ZN(
        P1_U3093) );
  AOI22_X1 U23396 ( .A1(n20748), .A2(n20437), .B1(n20747), .B2(n20436), .ZN(
        n20432) );
  AOI22_X1 U23397 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20439), .B1(
        n20438), .B2(n20687), .ZN(n20431) );
  OAI211_X1 U23398 ( .C1(n20690), .C2(n20442), .A(n20432), .B(n20431), .ZN(
        P1_U3094) );
  AOI22_X1 U23399 ( .A1(n20754), .A2(n20437), .B1(n20753), .B2(n20436), .ZN(
        n20434) );
  AOI22_X1 U23400 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20439), .B1(
        n20465), .B2(n20627), .ZN(n20433) );
  OAI211_X1 U23401 ( .C1(n20630), .C2(n20435), .A(n20434), .B(n20433), .ZN(
        P1_U3095) );
  AOI22_X1 U23402 ( .A1(n20764), .A2(n20437), .B1(n20762), .B2(n20436), .ZN(
        n20441) );
  AOI22_X1 U23403 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20439), .B1(
        n20438), .B2(n20701), .ZN(n20440) );
  OAI211_X1 U23404 ( .C1(n20706), .C2(n20442), .A(n20441), .B(n20440), .ZN(
        P1_U3096) );
  NOR3_X1 U23405 ( .A1(n20565), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20473) );
  INV_X1 U23406 ( .A(n20473), .ZN(n20469) );
  NOR2_X1 U23407 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20469), .ZN(
        n20464) );
  AND2_X1 U23408 ( .A1(n12753), .A2(n13145), .ZN(n20529) );
  AOI21_X1 U23409 ( .B1(n20529), .B2(n9741), .A(n20464), .ZN(n20446) );
  AND2_X1 U23410 ( .A1(n20443), .A2(n20490), .ZN(n20564) );
  INV_X1 U23411 ( .A(n20564), .ZN(n20569) );
  OAI22_X1 U23412 ( .A1(n20446), .A2(n20711), .B1(n20569), .B2(n20444), .ZN(
        n20463) );
  AOI22_X1 U23413 ( .A1(n21198), .A2(n20464), .B1(n20463), .B2(n21195), .ZN(
        n20450) );
  INV_X1 U23414 ( .A(n21204), .ZN(n20445) );
  OAI21_X1 U23415 ( .B1(n20445), .B2(n20465), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20447) );
  NAND2_X1 U23416 ( .A1(n20447), .A2(n20446), .ZN(n20448) );
  AOI22_X1 U23417 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20466), .B1(
        n20465), .B2(n20719), .ZN(n20449) );
  OAI211_X1 U23418 ( .C1(n20722), .C2(n21204), .A(n20450), .B(n20449), .ZN(
        P1_U3097) );
  AOI22_X1 U23419 ( .A1(n20724), .A2(n20464), .B1(n20463), .B2(n20723), .ZN(
        n20452) );
  AOI22_X1 U23420 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20466), .B1(
        n20465), .B2(n20725), .ZN(n20451) );
  OAI211_X1 U23421 ( .C1(n20728), .C2(n21204), .A(n20452), .B(n20451), .ZN(
        P1_U3098) );
  AOI22_X1 U23422 ( .A1(n20730), .A2(n20464), .B1(n20463), .B2(n20729), .ZN(
        n20454) );
  AOI22_X1 U23423 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20466), .B1(
        n20465), .B2(n20668), .ZN(n20453) );
  OAI211_X1 U23424 ( .C1(n20671), .C2(n21204), .A(n20454), .B(n20453), .ZN(
        P1_U3099) );
  AOI22_X1 U23425 ( .A1(n20736), .A2(n20464), .B1(n20463), .B2(n20735), .ZN(
        n20456) );
  AOI22_X1 U23426 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20466), .B1(
        n20465), .B2(n20675), .ZN(n20455) );
  OAI211_X1 U23427 ( .C1(n20678), .C2(n21204), .A(n20456), .B(n20455), .ZN(
        P1_U3100) );
  AOI22_X1 U23428 ( .A1(n20742), .A2(n20464), .B1(n20463), .B2(n20741), .ZN(
        n20458) );
  AOI22_X1 U23429 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20466), .B1(
        n20465), .B2(n20743), .ZN(n20457) );
  OAI211_X1 U23430 ( .C1(n20746), .C2(n21204), .A(n20458), .B(n20457), .ZN(
        P1_U3101) );
  AOI22_X1 U23431 ( .A1(n20748), .A2(n20464), .B1(n20463), .B2(n20747), .ZN(
        n20460) );
  AOI22_X1 U23432 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20466), .B1(
        n20465), .B2(n20687), .ZN(n20459) );
  OAI211_X1 U23433 ( .C1(n20690), .C2(n21204), .A(n20460), .B(n20459), .ZN(
        P1_U3102) );
  AOI22_X1 U23434 ( .A1(n20754), .A2(n20464), .B1(n20463), .B2(n20753), .ZN(
        n20462) );
  AOI22_X1 U23435 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20466), .B1(
        n20465), .B2(n20755), .ZN(n20461) );
  OAI211_X1 U23436 ( .C1(n20760), .C2(n21204), .A(n20462), .B(n20461), .ZN(
        P1_U3103) );
  AOI22_X1 U23437 ( .A1(n20764), .A2(n20464), .B1(n20463), .B2(n20762), .ZN(
        n20468) );
  AOI22_X1 U23438 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20466), .B1(
        n20465), .B2(n20701), .ZN(n20467) );
  OAI211_X1 U23439 ( .C1(n20706), .C2(n21204), .A(n20468), .B(n20467), .ZN(
        P1_U3104) );
  NOR2_X1 U23440 ( .A1(n20602), .A2(n20469), .ZN(n21197) );
  AOI21_X1 U23441 ( .B1(n20529), .B2(n20603), .A(n21197), .ZN(n20470) );
  OAI22_X1 U23442 ( .A1(n20470), .A2(n20711), .B1(n20469), .B2(n11307), .ZN(
        n21196) );
  AOI22_X1 U23443 ( .A1(n20724), .A2(n21197), .B1(n21196), .B2(n20723), .ZN(
        n20475) );
  OAI21_X1 U23444 ( .B1(n20536), .B2(n20471), .A(n20470), .ZN(n20472) );
  OAI221_X1 U23445 ( .B1(n20717), .B2(n20473), .C1(n20711), .C2(n20472), .A(
        n20716), .ZN(n21201) );
  AOI22_X1 U23446 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n21201), .B1(
        n21200), .B2(n20613), .ZN(n20474) );
  OAI211_X1 U23447 ( .C1(n20616), .C2(n21204), .A(n20475), .B(n20474), .ZN(
        P1_U3106) );
  AOI22_X1 U23448 ( .A1(n20730), .A2(n21197), .B1(n21196), .B2(n20729), .ZN(
        n20477) );
  AOI22_X1 U23449 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n21201), .B1(
        n21200), .B2(n20731), .ZN(n20476) );
  OAI211_X1 U23450 ( .C1(n20734), .C2(n21204), .A(n20477), .B(n20476), .ZN(
        P1_U3107) );
  AOI22_X1 U23451 ( .A1(n20736), .A2(n21197), .B1(n21196), .B2(n20735), .ZN(
        n20479) );
  AOI22_X1 U23452 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n21201), .B1(
        n21200), .B2(n20737), .ZN(n20478) );
  OAI211_X1 U23453 ( .C1(n20740), .C2(n21204), .A(n20479), .B(n20478), .ZN(
        P1_U3108) );
  AOI22_X1 U23454 ( .A1(n20742), .A2(n21197), .B1(n21196), .B2(n20741), .ZN(
        n20481) );
  AOI22_X1 U23455 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n21201), .B1(
        n21200), .B2(n20621), .ZN(n20480) );
  OAI211_X1 U23456 ( .C1(n20624), .C2(n21204), .A(n20481), .B(n20480), .ZN(
        P1_U3109) );
  AOI22_X1 U23457 ( .A1(n20748), .A2(n21197), .B1(n21196), .B2(n20747), .ZN(
        n20483) );
  AOI22_X1 U23458 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n21201), .B1(
        n21200), .B2(n20749), .ZN(n20482) );
  OAI211_X1 U23459 ( .C1(n20752), .C2(n21204), .A(n20483), .B(n20482), .ZN(
        P1_U3110) );
  AOI22_X1 U23460 ( .A1(n20754), .A2(n21197), .B1(n21196), .B2(n20753), .ZN(
        n20485) );
  AOI22_X1 U23461 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n21201), .B1(
        n21200), .B2(n20627), .ZN(n20484) );
  OAI211_X1 U23462 ( .C1(n20630), .C2(n21204), .A(n20485), .B(n20484), .ZN(
        P1_U3111) );
  AOI22_X1 U23463 ( .A1(n20764), .A2(n21197), .B1(n21196), .B2(n20762), .ZN(
        n20487) );
  AOI22_X1 U23464 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n21201), .B1(
        n21200), .B2(n20765), .ZN(n20486) );
  OAI211_X1 U23465 ( .C1(n20771), .C2(n21204), .A(n20487), .B(n20486), .ZN(
        P1_U3112) );
  NAND2_X1 U23466 ( .A1(n20556), .A2(n20717), .ZN(n20489) );
  OAI21_X1 U23467 ( .B1(n20489), .B2(n21200), .A(n20560), .ZN(n20494) );
  AND2_X1 U23468 ( .A1(n20529), .A2(n20652), .ZN(n20499) );
  OR2_X1 U23469 ( .A1(n20490), .A2(n20565), .ZN(n20495) );
  INV_X1 U23470 ( .A(n20495), .ZN(n20642) );
  NOR3_X1 U23471 ( .A1(n20565), .A2(n20492), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20534) );
  INV_X1 U23472 ( .A(n20534), .ZN(n20530) );
  NOR2_X1 U23473 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20530), .ZN(
        n20503) );
  INV_X1 U23474 ( .A(n20503), .ZN(n20522) );
  OAI22_X1 U23475 ( .A1(n20556), .A2(n20722), .B1(n20647), .B2(n20522), .ZN(
        n20493) );
  INV_X1 U23476 ( .A(n20493), .ZN(n20502) );
  INV_X1 U23477 ( .A(n20494), .ZN(n20500) );
  NAND2_X1 U23478 ( .A1(n20495), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20654) );
  OAI21_X1 U23479 ( .B1(n20573), .B2(n20503), .A(n20654), .ZN(n20496) );
  INV_X1 U23480 ( .A(n20496), .ZN(n20498) );
  AOI22_X1 U23481 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20524), .B1(
        n21200), .B2(n20719), .ZN(n20501) );
  OAI211_X1 U23482 ( .C1(n20527), .C2(n20646), .A(n20502), .B(n20501), .ZN(
        P1_U3113) );
  AOI22_X1 U23483 ( .A1(n21200), .A2(n20725), .B1(n20724), .B2(n20503), .ZN(
        n20506) );
  INV_X1 U23484 ( .A(n20556), .ZN(n20504) );
  AOI22_X1 U23485 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20524), .B1(
        n20504), .B2(n20613), .ZN(n20505) );
  OAI211_X1 U23486 ( .C1(n20527), .C2(n20660), .A(n20506), .B(n20505), .ZN(
        P1_U3114) );
  OAI22_X1 U23487 ( .A1(n20556), .A2(n20671), .B1(n20666), .B2(n20522), .ZN(
        n20507) );
  INV_X1 U23488 ( .A(n20507), .ZN(n20509) );
  AOI22_X1 U23489 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20524), .B1(
        n21200), .B2(n20668), .ZN(n20508) );
  OAI211_X1 U23490 ( .C1(n20527), .C2(n20665), .A(n20509), .B(n20508), .ZN(
        P1_U3115) );
  OAI22_X1 U23491 ( .A1(n20556), .A2(n20678), .B1(n20673), .B2(n20522), .ZN(
        n20510) );
  INV_X1 U23492 ( .A(n20510), .ZN(n20512) );
  AOI22_X1 U23493 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20524), .B1(
        n21200), .B2(n20675), .ZN(n20511) );
  OAI211_X1 U23494 ( .C1(n20527), .C2(n20672), .A(n20512), .B(n20511), .ZN(
        P1_U3116) );
  OAI22_X1 U23495 ( .A1(n20556), .A2(n20746), .B1(n20680), .B2(n20522), .ZN(
        n20513) );
  INV_X1 U23496 ( .A(n20513), .ZN(n20515) );
  AOI22_X1 U23497 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20524), .B1(
        n21200), .B2(n20743), .ZN(n20514) );
  OAI211_X1 U23498 ( .C1(n20527), .C2(n20679), .A(n20515), .B(n20514), .ZN(
        P1_U3117) );
  OAI22_X1 U23499 ( .A1(n20556), .A2(n20690), .B1(n20685), .B2(n20522), .ZN(
        n20516) );
  INV_X1 U23500 ( .A(n20516), .ZN(n20518) );
  AOI22_X1 U23501 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20524), .B1(
        n21200), .B2(n20687), .ZN(n20517) );
  OAI211_X1 U23502 ( .C1(n20527), .C2(n20684), .A(n20518), .B(n20517), .ZN(
        P1_U3118) );
  OAI22_X1 U23503 ( .A1(n20556), .A2(n20760), .B1(n20692), .B2(n20522), .ZN(
        n20519) );
  INV_X1 U23504 ( .A(n20519), .ZN(n20521) );
  AOI22_X1 U23505 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20524), .B1(
        n21200), .B2(n20755), .ZN(n20520) );
  OAI211_X1 U23506 ( .C1(n20527), .C2(n20691), .A(n20521), .B(n20520), .ZN(
        P1_U3119) );
  OAI22_X1 U23507 ( .A1(n20556), .A2(n20706), .B1(n20699), .B2(n20522), .ZN(
        n20523) );
  INV_X1 U23508 ( .A(n20523), .ZN(n20526) );
  AOI22_X1 U23509 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20524), .B1(
        n21200), .B2(n20701), .ZN(n20525) );
  OAI211_X1 U23510 ( .C1(n20527), .C2(n20697), .A(n20526), .B(n20525), .ZN(
        P1_U3120) );
  NOR2_X1 U23511 ( .A1(n20528), .A2(n20565), .ZN(n20552) );
  AOI21_X1 U23512 ( .B1(n20529), .B2(n20708), .A(n20552), .ZN(n20531) );
  OAI22_X1 U23513 ( .A1(n20531), .A2(n20711), .B1(n20530), .B2(n11307), .ZN(
        n20551) );
  AOI22_X1 U23514 ( .A1(n21198), .A2(n20552), .B1(n20551), .B2(n21195), .ZN(
        n20538) );
  OAI21_X1 U23515 ( .B1(n20536), .B2(n20532), .A(n20531), .ZN(n20533) );
  OAI221_X1 U23516 ( .B1(n20717), .B2(n20534), .C1(n20711), .C2(n20533), .A(
        n20716), .ZN(n20553) );
  AOI22_X1 U23517 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20553), .B1(
        n20597), .B2(n21199), .ZN(n20537) );
  OAI211_X1 U23518 ( .C1(n21205), .C2(n20556), .A(n20538), .B(n20537), .ZN(
        P1_U3121) );
  AOI22_X1 U23519 ( .A1(n20724), .A2(n20552), .B1(n20551), .B2(n20723), .ZN(
        n20540) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20553), .B1(
        n20597), .B2(n20613), .ZN(n20539) );
  OAI211_X1 U23521 ( .C1(n20616), .C2(n20556), .A(n20540), .B(n20539), .ZN(
        P1_U3122) );
  AOI22_X1 U23522 ( .A1(n20730), .A2(n20552), .B1(n20551), .B2(n20729), .ZN(
        n20542) );
  AOI22_X1 U23523 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20553), .B1(
        n20597), .B2(n20731), .ZN(n20541) );
  OAI211_X1 U23524 ( .C1(n20734), .C2(n20556), .A(n20542), .B(n20541), .ZN(
        P1_U3123) );
  AOI22_X1 U23525 ( .A1(n20736), .A2(n20552), .B1(n20551), .B2(n20735), .ZN(
        n20544) );
  AOI22_X1 U23526 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20553), .B1(
        n20597), .B2(n20737), .ZN(n20543) );
  OAI211_X1 U23527 ( .C1(n20740), .C2(n20556), .A(n20544), .B(n20543), .ZN(
        P1_U3124) );
  AOI22_X1 U23528 ( .A1(n20742), .A2(n20552), .B1(n20551), .B2(n20741), .ZN(
        n20546) );
  AOI22_X1 U23529 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20553), .B1(
        n20597), .B2(n20621), .ZN(n20545) );
  OAI211_X1 U23530 ( .C1(n20624), .C2(n20556), .A(n20546), .B(n20545), .ZN(
        P1_U3125) );
  AOI22_X1 U23531 ( .A1(n20748), .A2(n20552), .B1(n20551), .B2(n20747), .ZN(
        n20548) );
  AOI22_X1 U23532 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20553), .B1(
        n20597), .B2(n20749), .ZN(n20547) );
  OAI211_X1 U23533 ( .C1(n20752), .C2(n20556), .A(n20548), .B(n20547), .ZN(
        P1_U3126) );
  AOI22_X1 U23534 ( .A1(n20754), .A2(n20552), .B1(n20551), .B2(n20753), .ZN(
        n20550) );
  AOI22_X1 U23535 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20553), .B1(
        n20597), .B2(n20627), .ZN(n20549) );
  OAI211_X1 U23536 ( .C1(n20630), .C2(n20556), .A(n20550), .B(n20549), .ZN(
        P1_U3127) );
  AOI22_X1 U23537 ( .A1(n20764), .A2(n20552), .B1(n20551), .B2(n20762), .ZN(
        n20555) );
  AOI22_X1 U23538 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20553), .B1(
        n20597), .B2(n20765), .ZN(n20554) );
  OAI211_X1 U23539 ( .C1(n20771), .C2(n20556), .A(n20555), .B(n20554), .ZN(
        P1_U3128) );
  INV_X1 U23540 ( .A(n20597), .ZN(n20559) );
  INV_X1 U23541 ( .A(n20557), .ZN(n20558) );
  NAND3_X1 U23542 ( .A1(n20559), .A2(n20717), .A3(n20636), .ZN(n20561) );
  NAND2_X1 U23543 ( .A1(n20561), .A2(n20560), .ZN(n20571) );
  OR2_X1 U23544 ( .A1(n13145), .A2(n20562), .ZN(n20641) );
  NOR2_X1 U23545 ( .A1(n20641), .A2(n20652), .ZN(n20568) );
  INV_X1 U23546 ( .A(n20563), .ZN(n20643) );
  NOR3_X1 U23547 ( .A1(n20566), .A2(n20565), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20609) );
  INV_X1 U23548 ( .A(n20609), .ZN(n20604) );
  NOR2_X1 U23549 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20604), .ZN(
        n20574) );
  INV_X1 U23550 ( .A(n20574), .ZN(n20595) );
  OAI22_X1 U23551 ( .A1(n20636), .A2(n20722), .B1(n20647), .B2(n20595), .ZN(
        n20567) );
  INV_X1 U23552 ( .A(n20567), .ZN(n20576) );
  INV_X1 U23553 ( .A(n20568), .ZN(n20570) );
  AOI22_X1 U23554 ( .A1(n20571), .A2(n20570), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20569), .ZN(n20572) );
  OAI211_X1 U23555 ( .C1(n20574), .C2(n20573), .A(n20655), .B(n20572), .ZN(
        n20598) );
  AOI22_X1 U23556 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20719), .ZN(n20575) );
  OAI211_X1 U23557 ( .C1(n20601), .C2(n20646), .A(n20576), .B(n20575), .ZN(
        P1_U3129) );
  OAI22_X1 U23558 ( .A1(n20636), .A2(n20728), .B1(n20661), .B2(n20595), .ZN(
        n20577) );
  INV_X1 U23559 ( .A(n20577), .ZN(n20579) );
  AOI22_X1 U23560 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20725), .ZN(n20578) );
  OAI211_X1 U23561 ( .C1(n20601), .C2(n20660), .A(n20579), .B(n20578), .ZN(
        P1_U3130) );
  OAI22_X1 U23562 ( .A1(n20636), .A2(n20671), .B1(n20666), .B2(n20595), .ZN(
        n20580) );
  INV_X1 U23563 ( .A(n20580), .ZN(n20582) );
  AOI22_X1 U23564 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20668), .ZN(n20581) );
  OAI211_X1 U23565 ( .C1(n20601), .C2(n20665), .A(n20582), .B(n20581), .ZN(
        P1_U3131) );
  OAI22_X1 U23566 ( .A1(n20636), .A2(n20678), .B1(n20673), .B2(n20595), .ZN(
        n20583) );
  INV_X1 U23567 ( .A(n20583), .ZN(n20585) );
  AOI22_X1 U23568 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20675), .ZN(n20584) );
  OAI211_X1 U23569 ( .C1(n20601), .C2(n20672), .A(n20585), .B(n20584), .ZN(
        P1_U3132) );
  OAI22_X1 U23570 ( .A1(n20636), .A2(n20746), .B1(n20680), .B2(n20595), .ZN(
        n20586) );
  INV_X1 U23571 ( .A(n20586), .ZN(n20588) );
  AOI22_X1 U23572 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20743), .ZN(n20587) );
  OAI211_X1 U23573 ( .C1(n20601), .C2(n20679), .A(n20588), .B(n20587), .ZN(
        P1_U3133) );
  OAI22_X1 U23574 ( .A1(n20636), .A2(n20690), .B1(n20685), .B2(n20595), .ZN(
        n20589) );
  INV_X1 U23575 ( .A(n20589), .ZN(n20591) );
  AOI22_X1 U23576 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20687), .ZN(n20590) );
  OAI211_X1 U23577 ( .C1(n20601), .C2(n20684), .A(n20591), .B(n20590), .ZN(
        P1_U3134) );
  OAI22_X1 U23578 ( .A1(n20636), .A2(n20760), .B1(n20692), .B2(n20595), .ZN(
        n20592) );
  INV_X1 U23579 ( .A(n20592), .ZN(n20594) );
  AOI22_X1 U23580 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20755), .ZN(n20593) );
  OAI211_X1 U23581 ( .C1(n20601), .C2(n20691), .A(n20594), .B(n20593), .ZN(
        P1_U3135) );
  OAI22_X1 U23582 ( .A1(n20636), .A2(n20706), .B1(n20699), .B2(n20595), .ZN(
        n20596) );
  INV_X1 U23583 ( .A(n20596), .ZN(n20600) );
  AOI22_X1 U23584 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20598), .B1(
        n20597), .B2(n20701), .ZN(n20599) );
  OAI211_X1 U23585 ( .C1(n20601), .C2(n20697), .A(n20600), .B(n20599), .ZN(
        P1_U3136) );
  NOR2_X1 U23586 ( .A1(n20602), .A2(n20604), .ZN(n20632) );
  INV_X1 U23587 ( .A(n20641), .ZN(n20709) );
  AOI21_X1 U23588 ( .B1(n20709), .B2(n20603), .A(n20632), .ZN(n20606) );
  OAI22_X1 U23589 ( .A1(n20606), .A2(n20711), .B1(n20604), .B2(n11307), .ZN(
        n20631) );
  AOI22_X1 U23590 ( .A1(n21198), .A2(n20632), .B1(n21195), .B2(n20631), .ZN(
        n20612) );
  INV_X1 U23591 ( .A(n20605), .ZN(n20607) );
  NAND2_X1 U23592 ( .A1(n20607), .A2(n20606), .ZN(n20608) );
  OAI221_X1 U23593 ( .B1(n20717), .B2(n20609), .C1(n20711), .C2(n20608), .A(
        n20716), .ZN(n20633) );
  AOI22_X1 U23594 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20633), .B1(
        n20702), .B2(n21199), .ZN(n20611) );
  OAI211_X1 U23595 ( .C1(n21205), .C2(n20636), .A(n20612), .B(n20611), .ZN(
        P1_U3137) );
  AOI22_X1 U23596 ( .A1(n20724), .A2(n20632), .B1(n20723), .B2(n20631), .ZN(
        n20615) );
  AOI22_X1 U23597 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20633), .B1(
        n20702), .B2(n20613), .ZN(n20614) );
  OAI211_X1 U23598 ( .C1(n20616), .C2(n20636), .A(n20615), .B(n20614), .ZN(
        P1_U3138) );
  AOI22_X1 U23599 ( .A1(n20730), .A2(n20632), .B1(n20729), .B2(n20631), .ZN(
        n20618) );
  AOI22_X1 U23600 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20633), .B1(
        n20702), .B2(n20731), .ZN(n20617) );
  OAI211_X1 U23601 ( .C1(n20734), .C2(n20636), .A(n20618), .B(n20617), .ZN(
        P1_U3139) );
  AOI22_X1 U23602 ( .A1(n20736), .A2(n20632), .B1(n20735), .B2(n20631), .ZN(
        n20620) );
  AOI22_X1 U23603 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20633), .B1(
        n20702), .B2(n20737), .ZN(n20619) );
  OAI211_X1 U23604 ( .C1(n20740), .C2(n20636), .A(n20620), .B(n20619), .ZN(
        P1_U3140) );
  AOI22_X1 U23605 ( .A1(n20742), .A2(n20632), .B1(n20741), .B2(n20631), .ZN(
        n20623) );
  AOI22_X1 U23606 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20633), .B1(
        n20702), .B2(n20621), .ZN(n20622) );
  OAI211_X1 U23607 ( .C1(n20624), .C2(n20636), .A(n20623), .B(n20622), .ZN(
        P1_U3141) );
  AOI22_X1 U23608 ( .A1(n20748), .A2(n20632), .B1(n20747), .B2(n20631), .ZN(
        n20626) );
  AOI22_X1 U23609 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20633), .B1(
        n20702), .B2(n20749), .ZN(n20625) );
  OAI211_X1 U23610 ( .C1(n20752), .C2(n20636), .A(n20626), .B(n20625), .ZN(
        P1_U3142) );
  AOI22_X1 U23611 ( .A1(n20754), .A2(n20632), .B1(n20753), .B2(n20631), .ZN(
        n20629) );
  AOI22_X1 U23612 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20633), .B1(
        n20702), .B2(n20627), .ZN(n20628) );
  OAI211_X1 U23613 ( .C1(n20630), .C2(n20636), .A(n20629), .B(n20628), .ZN(
        P1_U3143) );
  AOI22_X1 U23614 ( .A1(n20764), .A2(n20632), .B1(n20762), .B2(n20631), .ZN(
        n20635) );
  AOI22_X1 U23615 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20633), .B1(
        n20702), .B2(n20765), .ZN(n20634) );
  OAI211_X1 U23616 ( .C1(n20771), .C2(n20636), .A(n20635), .B(n20634), .ZN(
        P1_U3144) );
  INV_X1 U23617 ( .A(n20637), .ZN(n20638) );
  INV_X1 U23618 ( .A(n20718), .ZN(n20710) );
  NOR2_X1 U23619 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20710), .ZN(
        n20657) );
  INV_X1 U23620 ( .A(n20657), .ZN(n20698) );
  OR2_X1 U23621 ( .A1(n9741), .A2(n20711), .ZN(n20640) );
  OR2_X1 U23622 ( .A1(n20641), .A2(n20640), .ZN(n20645) );
  NAND2_X1 U23623 ( .A1(n20643), .A2(n20642), .ZN(n20644) );
  AND2_X1 U23624 ( .A1(n20645), .A2(n20644), .ZN(n20696) );
  OAI22_X1 U23625 ( .A1(n20647), .A2(n20698), .B1(n20646), .B2(n20696), .ZN(
        n20648) );
  INV_X1 U23626 ( .A(n20648), .ZN(n20659) );
  AOI21_X1 U23627 ( .B1(n20770), .B2(n20650), .A(n20649), .ZN(n20651) );
  AOI21_X1 U23628 ( .B1(n20709), .B2(n20652), .A(n20651), .ZN(n20653) );
  NOR2_X1 U23629 ( .A1(n20653), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20656) );
  AOI22_X1 U23630 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20703), .B1(
        n20702), .B2(n20719), .ZN(n20658) );
  OAI211_X1 U23631 ( .C1(n20722), .C2(n20770), .A(n20659), .B(n20658), .ZN(
        P1_U3145) );
  OAI22_X1 U23632 ( .A1(n20661), .A2(n20698), .B1(n20660), .B2(n20696), .ZN(
        n20662) );
  INV_X1 U23633 ( .A(n20662), .ZN(n20664) );
  AOI22_X1 U23634 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20703), .B1(
        n20702), .B2(n20725), .ZN(n20663) );
  OAI211_X1 U23635 ( .C1(n20728), .C2(n20770), .A(n20664), .B(n20663), .ZN(
        P1_U3146) );
  OAI22_X1 U23636 ( .A1(n20666), .A2(n20698), .B1(n20665), .B2(n20696), .ZN(
        n20667) );
  INV_X1 U23637 ( .A(n20667), .ZN(n20670) );
  AOI22_X1 U23638 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20703), .B1(
        n20702), .B2(n20668), .ZN(n20669) );
  OAI211_X1 U23639 ( .C1(n20671), .C2(n20770), .A(n20670), .B(n20669), .ZN(
        P1_U3147) );
  OAI22_X1 U23640 ( .A1(n20673), .A2(n20698), .B1(n20672), .B2(n20696), .ZN(
        n20674) );
  INV_X1 U23641 ( .A(n20674), .ZN(n20677) );
  AOI22_X1 U23642 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20703), .B1(
        n20702), .B2(n20675), .ZN(n20676) );
  OAI211_X1 U23643 ( .C1(n20678), .C2(n20770), .A(n20677), .B(n20676), .ZN(
        P1_U3148) );
  OAI22_X1 U23644 ( .A1(n20680), .A2(n20698), .B1(n20679), .B2(n20696), .ZN(
        n20681) );
  INV_X1 U23645 ( .A(n20681), .ZN(n20683) );
  AOI22_X1 U23646 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20703), .B1(
        n20702), .B2(n20743), .ZN(n20682) );
  OAI211_X1 U23647 ( .C1(n20746), .C2(n20770), .A(n20683), .B(n20682), .ZN(
        P1_U3149) );
  OAI22_X1 U23648 ( .A1(n20685), .A2(n20698), .B1(n20684), .B2(n20696), .ZN(
        n20686) );
  INV_X1 U23649 ( .A(n20686), .ZN(n20689) );
  AOI22_X1 U23650 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20703), .B1(
        n20702), .B2(n20687), .ZN(n20688) );
  OAI211_X1 U23651 ( .C1(n20690), .C2(n20770), .A(n20689), .B(n20688), .ZN(
        P1_U3150) );
  OAI22_X1 U23652 ( .A1(n20692), .A2(n20698), .B1(n20691), .B2(n20696), .ZN(
        n20693) );
  INV_X1 U23653 ( .A(n20693), .ZN(n20695) );
  AOI22_X1 U23654 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20703), .B1(
        n20702), .B2(n20755), .ZN(n20694) );
  OAI211_X1 U23655 ( .C1(n20760), .C2(n20770), .A(n20695), .B(n20694), .ZN(
        P1_U3151) );
  OAI22_X1 U23656 ( .A1(n20699), .A2(n20698), .B1(n20697), .B2(n20696), .ZN(
        n20700) );
  INV_X1 U23657 ( .A(n20700), .ZN(n20705) );
  AOI22_X1 U23658 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20703), .B1(
        n20702), .B2(n20701), .ZN(n20704) );
  OAI211_X1 U23659 ( .C1(n20706), .C2(n20770), .A(n20705), .B(n20704), .ZN(
        P1_U3152) );
  INV_X1 U23660 ( .A(n20707), .ZN(n20763) );
  AOI21_X1 U23661 ( .B1(n20709), .B2(n20708), .A(n20763), .ZN(n20712) );
  OAI22_X1 U23662 ( .A1(n20712), .A2(n20711), .B1(n11307), .B2(n20710), .ZN(
        n20761) );
  AOI22_X1 U23663 ( .A1(n21198), .A2(n20763), .B1(n21195), .B2(n20761), .ZN(
        n20721) );
  OAI21_X1 U23664 ( .B1(n20714), .B2(n20713), .A(n20712), .ZN(n20715) );
  INV_X1 U23665 ( .A(n20770), .ZN(n20756) );
  AOI22_X1 U23666 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20767), .B1(
        n20756), .B2(n20719), .ZN(n20720) );
  OAI211_X1 U23667 ( .C1(n20722), .C2(n20759), .A(n20721), .B(n20720), .ZN(
        P1_U3153) );
  AOI22_X1 U23668 ( .A1(n20724), .A2(n20763), .B1(n20723), .B2(n20761), .ZN(
        n20727) );
  AOI22_X1 U23669 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20767), .B1(
        n20756), .B2(n20725), .ZN(n20726) );
  OAI211_X1 U23670 ( .C1(n20728), .C2(n20759), .A(n20727), .B(n20726), .ZN(
        P1_U3154) );
  AOI22_X1 U23671 ( .A1(n20730), .A2(n20763), .B1(n20729), .B2(n20761), .ZN(
        n20733) );
  INV_X1 U23672 ( .A(n20759), .ZN(n20766) );
  AOI22_X1 U23673 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20767), .B1(
        n20766), .B2(n20731), .ZN(n20732) );
  OAI211_X1 U23674 ( .C1(n20734), .C2(n20770), .A(n20733), .B(n20732), .ZN(
        P1_U3155) );
  AOI22_X1 U23675 ( .A1(n20736), .A2(n20763), .B1(n20735), .B2(n20761), .ZN(
        n20739) );
  AOI22_X1 U23676 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20767), .B1(
        n20766), .B2(n20737), .ZN(n20738) );
  OAI211_X1 U23677 ( .C1(n20740), .C2(n20770), .A(n20739), .B(n20738), .ZN(
        P1_U3156) );
  AOI22_X1 U23678 ( .A1(n20742), .A2(n20763), .B1(n20741), .B2(n20761), .ZN(
        n20745) );
  AOI22_X1 U23679 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20767), .B1(
        n20756), .B2(n20743), .ZN(n20744) );
  OAI211_X1 U23680 ( .C1(n20746), .C2(n20759), .A(n20745), .B(n20744), .ZN(
        P1_U3157) );
  AOI22_X1 U23681 ( .A1(n20748), .A2(n20763), .B1(n20747), .B2(n20761), .ZN(
        n20751) );
  AOI22_X1 U23682 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20767), .B1(
        n20766), .B2(n20749), .ZN(n20750) );
  OAI211_X1 U23683 ( .C1(n20752), .C2(n20770), .A(n20751), .B(n20750), .ZN(
        P1_U3158) );
  AOI22_X1 U23684 ( .A1(n20754), .A2(n20763), .B1(n20753), .B2(n20761), .ZN(
        n20758) );
  AOI22_X1 U23685 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20767), .B1(
        n20756), .B2(n20755), .ZN(n20757) );
  OAI211_X1 U23686 ( .C1(n20760), .C2(n20759), .A(n20758), .B(n20757), .ZN(
        P1_U3159) );
  AOI22_X1 U23687 ( .A1(n20764), .A2(n20763), .B1(n20762), .B2(n20761), .ZN(
        n20769) );
  AOI22_X1 U23688 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20767), .B1(
        n20766), .B2(n20765), .ZN(n20768) );
  OAI211_X1 U23689 ( .C1(n20771), .C2(n20770), .A(n20769), .B(n20768), .ZN(
        P1_U3160) );
  NOR2_X1 U23690 ( .A1(n20773), .A2(n20772), .ZN(n20776) );
  INV_X1 U23691 ( .A(n20774), .ZN(n20775) );
  OAI21_X1 U23692 ( .B1(n20776), .B2(n11307), .A(n20775), .ZN(P1_U3163) );
  AND2_X1 U23693 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20777), .ZN(
        P1_U3164) );
  AND2_X1 U23694 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20777), .ZN(
        P1_U3165) );
  AND2_X1 U23695 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20777), .ZN(
        P1_U3166) );
  AND2_X1 U23696 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20777), .ZN(
        P1_U3167) );
  AND2_X1 U23697 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20777), .ZN(
        P1_U3168) );
  AND2_X1 U23698 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20777), .ZN(
        P1_U3169) );
  AND2_X1 U23699 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20777), .ZN(
        P1_U3170) );
  AND2_X1 U23700 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20777), .ZN(
        P1_U3171) );
  AND2_X1 U23701 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20777), .ZN(
        P1_U3172) );
  AND2_X1 U23702 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20777), .ZN(
        P1_U3173) );
  AND2_X1 U23703 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20777), .ZN(
        P1_U3174) );
  AND2_X1 U23704 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20777), .ZN(
        P1_U3175) );
  AND2_X1 U23705 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20777), .ZN(
        P1_U3176) );
  AND2_X1 U23706 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20777), .ZN(
        P1_U3177) );
  AND2_X1 U23707 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20777), .ZN(
        P1_U3178) );
  AND2_X1 U23708 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20777), .ZN(
        P1_U3179) );
  AND2_X1 U23709 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20777), .ZN(
        P1_U3180) );
  AND2_X1 U23710 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20777), .ZN(
        P1_U3181) );
  AND2_X1 U23711 ( .A1(n20777), .A2(P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(
        P1_U3182) );
  AND2_X1 U23712 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20777), .ZN(
        P1_U3183) );
  AND2_X1 U23713 ( .A1(n20777), .A2(P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(
        P1_U3184) );
  AND2_X1 U23714 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20777), .ZN(
        P1_U3185) );
  AND2_X1 U23715 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20777), .ZN(P1_U3186) );
  AND2_X1 U23716 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20777), .ZN(P1_U3187) );
  AND2_X1 U23717 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20777), .ZN(P1_U3188) );
  AND2_X1 U23718 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20777), .ZN(P1_U3189) );
  AND2_X1 U23719 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20777), .ZN(P1_U3190) );
  AND2_X1 U23720 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20777), .ZN(P1_U3191) );
  AND2_X1 U23721 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20777), .ZN(P1_U3192) );
  AND2_X1 U23722 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20777), .ZN(P1_U3193) );
  AOI21_X1 U23723 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20783), .A(n20786), 
        .ZN(n20791) );
  NOR2_X1 U23724 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20779) );
  OAI21_X1 U23725 ( .B1(n20779), .B2(n20778), .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20780) );
  AOI21_X1 U23726 ( .B1(NA), .B2(n20786), .A(n20780), .ZN(n20781) );
  OAI22_X1 U23727 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20791), .B1(n20853), 
        .B2(n20781), .ZN(P1_U3194) );
  AOI21_X1 U23728 ( .B1(n20783), .B2(n20788), .A(n20782), .ZN(n20793) );
  INV_X1 U23729 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20785) );
  OAI211_X1 U23730 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20785), .A(
        P1_STATE_REG_0__SCAN_IN), .B(HOLD), .ZN(n20792) );
  INV_X1 U23731 ( .A(n20784), .ZN(n20789) );
  NOR2_X1 U23732 ( .A1(n20786), .A2(n20785), .ZN(n20787) );
  OAI22_X1 U23733 ( .A1(n20789), .A2(n20788), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n20787), .ZN(n20790) );
  OAI22_X1 U23734 ( .A1(n20793), .A2(n20792), .B1(n20791), .B2(n20790), .ZN(
        P1_U3196) );
  OR2_X1 U23735 ( .A1(n20864), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20835) );
  NOR2_X1 U23736 ( .A1(n20794), .A2(n20864), .ZN(n20827) );
  OAI222_X1 U23737 ( .A1(n20835), .A2(n13376), .B1(n20795), .B2(n20853), .C1(
        n14140), .C2(n20831), .ZN(P1_U3197) );
  INV_X1 U23738 ( .A(n20831), .ZN(n20833) );
  AOI222_X1 U23739 ( .A1(n20833), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20864), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20829), .ZN(n20796) );
  INV_X1 U23740 ( .A(n20796), .ZN(P1_U3198) );
  AOI222_X1 U23741 ( .A1(n20833), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n20864), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20829), .ZN(n20797) );
  INV_X1 U23742 ( .A(n20797), .ZN(P1_U3199) );
  AOI222_X1 U23743 ( .A1(n20833), .A2(P1_REIP_REG_4__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20864), .C1(P1_REIP_REG_5__SCAN_IN), 
        .C2(n20829), .ZN(n20798) );
  INV_X1 U23744 ( .A(n20798), .ZN(P1_U3200) );
  AOI222_X1 U23745 ( .A1(n20833), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20864), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20829), .ZN(n20799) );
  INV_X1 U23746 ( .A(n20799), .ZN(P1_U3201) );
  AOI222_X1 U23747 ( .A1(n20833), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20864), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20829), .ZN(n20800) );
  INV_X1 U23748 ( .A(n20800), .ZN(P1_U3202) );
  INV_X1 U23749 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n21144) );
  OAI222_X1 U23750 ( .A1(n20831), .A2(n20801), .B1(n21144), .B2(n20853), .C1(
        n20803), .C2(n20835), .ZN(P1_U3203) );
  AOI22_X1 U23751 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n20864), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20829), .ZN(n20802) );
  OAI21_X1 U23752 ( .B1(n20803), .B2(n20831), .A(n20802), .ZN(P1_U3204) );
  AOI22_X1 U23753 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(n20864), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20833), .ZN(n20804) );
  OAI21_X1 U23754 ( .B1(n20805), .B2(n20835), .A(n20804), .ZN(P1_U3205) );
  AOI222_X1 U23755 ( .A1(n20829), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20864), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20833), .ZN(n20806) );
  INV_X1 U23756 ( .A(n20806), .ZN(P1_U3206) );
  AOI22_X1 U23757 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n20864), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20829), .ZN(n20807) );
  OAI21_X1 U23758 ( .B1(n20808), .B2(n20831), .A(n20807), .ZN(P1_U3207) );
  AOI22_X1 U23759 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n20864), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20833), .ZN(n20809) );
  OAI21_X1 U23760 ( .B1(n20810), .B2(n20835), .A(n20809), .ZN(P1_U3208) );
  AOI222_X1 U23761 ( .A1(n20833), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20864), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20829), .ZN(n20811) );
  INV_X1 U23762 ( .A(n20811), .ZN(P1_U3209) );
  AOI222_X1 U23763 ( .A1(n20833), .A2(P1_REIP_REG_14__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20864), .C1(P1_REIP_REG_15__SCAN_IN), 
        .C2(n20829), .ZN(n20812) );
  INV_X1 U23764 ( .A(n20812), .ZN(P1_U3210) );
  AOI222_X1 U23765 ( .A1(n20833), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20864), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20829), .ZN(n20813) );
  INV_X1 U23766 ( .A(n20813), .ZN(P1_U3211) );
  INV_X1 U23767 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n21125) );
  OAI222_X1 U23768 ( .A1(n20831), .A2(n20815), .B1(n21125), .B2(n20853), .C1(
        n20814), .C2(n20835), .ZN(P1_U3212) );
  AOI222_X1 U23769 ( .A1(n20833), .A2(P1_REIP_REG_17__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n20864), .C1(P1_REIP_REG_18__SCAN_IN), 
        .C2(n20829), .ZN(n20816) );
  INV_X1 U23770 ( .A(n20816), .ZN(P1_U3213) );
  AOI222_X1 U23771 ( .A1(n20827), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20864), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20829), .ZN(n20817) );
  INV_X1 U23772 ( .A(n20817), .ZN(P1_U3214) );
  AOI222_X1 U23773 ( .A1(n20827), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20864), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n20829), .ZN(n20818) );
  INV_X1 U23774 ( .A(n20818), .ZN(P1_U3215) );
  AOI222_X1 U23775 ( .A1(n20827), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20864), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20829), .ZN(n20819) );
  INV_X1 U23776 ( .A(n20819), .ZN(P1_U3216) );
  AOI222_X1 U23777 ( .A1(n20829), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20864), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20833), .ZN(n20820) );
  INV_X1 U23778 ( .A(n20820), .ZN(P1_U3217) );
  AOI222_X1 U23779 ( .A1(n20827), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20864), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20829), .ZN(n20821) );
  INV_X1 U23780 ( .A(n20821), .ZN(P1_U3218) );
  AOI222_X1 U23781 ( .A1(n20829), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20864), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20833), .ZN(n20822) );
  INV_X1 U23782 ( .A(n20822), .ZN(P1_U3219) );
  AOI222_X1 U23783 ( .A1(n20827), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20864), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20829), .ZN(n20823) );
  INV_X1 U23784 ( .A(n20823), .ZN(P1_U3220) );
  AOI222_X1 U23785 ( .A1(n20827), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20864), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20829), .ZN(n20824) );
  INV_X1 U23786 ( .A(n20824), .ZN(P1_U3221) );
  AOI222_X1 U23787 ( .A1(n20833), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20864), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20829), .ZN(n20825) );
  INV_X1 U23788 ( .A(n20825), .ZN(P1_U3222) );
  AOI222_X1 U23789 ( .A1(n20827), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20864), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20829), .ZN(n20826) );
  INV_X1 U23790 ( .A(n20826), .ZN(P1_U3223) );
  AOI222_X1 U23791 ( .A1(n20827), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20864), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20829), .ZN(n20828) );
  INV_X1 U23792 ( .A(n20828), .ZN(P1_U3224) );
  AOI22_X1 U23793 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20829), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20864), .ZN(n20830) );
  OAI21_X1 U23794 ( .B1(n20832), .B2(n20831), .A(n20830), .ZN(P1_U3225) );
  AOI22_X1 U23795 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20833), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20864), .ZN(n20834) );
  OAI21_X1 U23796 ( .B1(n20836), .B2(n20835), .A(n20834), .ZN(P1_U3226) );
  OAI22_X1 U23797 ( .A1(n20864), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20853), .ZN(n20837) );
  INV_X1 U23798 ( .A(n20837), .ZN(P1_U3458) );
  OAI22_X1 U23799 ( .A1(n20864), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20853), .ZN(n20838) );
  INV_X1 U23800 ( .A(n20838), .ZN(P1_U3459) );
  OAI22_X1 U23801 ( .A1(n20864), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20853), .ZN(n20839) );
  INV_X1 U23802 ( .A(n20839), .ZN(P1_U3460) );
  OAI22_X1 U23803 ( .A1(n20864), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20853), .ZN(n20840) );
  INV_X1 U23804 ( .A(n20840), .ZN(P1_U3461) );
  OAI21_X1 U23805 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20844), .A(n20842), 
        .ZN(n20841) );
  INV_X1 U23806 ( .A(n20841), .ZN(P1_U3464) );
  OAI21_X1 U23807 ( .B1(n20844), .B2(n20843), .A(n20842), .ZN(P1_U3465) );
  AOI211_X1 U23808 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_REIP_REG_1__SCAN_IN), .B(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20845) );
  AOI21_X1 U23809 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20845), .ZN(n20847) );
  INV_X1 U23810 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20846) );
  AOI22_X1 U23811 ( .A1(n20851), .A2(n20847), .B1(n20846), .B2(n20848), .ZN(
        P1_U3481) );
  NOR2_X1 U23812 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n20850) );
  INV_X1 U23813 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20849) );
  AOI22_X1 U23814 ( .A1(n20851), .A2(n20850), .B1(n20849), .B2(n20848), .ZN(
        P1_U3482) );
  AOI22_X1 U23815 ( .A1(n20853), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20852), 
        .B2(n20864), .ZN(P1_U3483) );
  AOI211_X1 U23816 ( .C1(n20075), .C2(n20856), .A(n20855), .B(n20854), .ZN(
        n20863) );
  OAI211_X1 U23817 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20858), .A(n20857), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20860) );
  AOI21_X1 U23818 ( .B1(n20860), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n20859), 
        .ZN(n20862) );
  NAND2_X1 U23819 ( .A1(n20863), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20861) );
  OAI21_X1 U23820 ( .B1(n20863), .B2(n20862), .A(n20861), .ZN(P1_U3485) );
  MUX2_X1 U23821 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n20864), .Z(P1_U3486) );
  INV_X1 U23822 ( .A(keyinput25), .ZN(n20865) );
  NAND4_X1 U23823 ( .A1(keyinput19), .A2(keyinput38), .A3(keyinput52), .A4(
        n20865), .ZN(n20866) );
  NOR3_X1 U23824 ( .A1(keyinput33), .A2(keyinput2), .A3(n20866), .ZN(n20878)
         );
  NAND2_X1 U23825 ( .A1(keyinput24), .A2(keyinput1), .ZN(n20867) );
  NOR3_X1 U23826 ( .A1(keyinput12), .A2(keyinput87), .A3(n20867), .ZN(n20868)
         );
  NAND3_X1 U23827 ( .A1(keyinput0), .A2(keyinput63), .A3(n20868), .ZN(n20876)
         );
  INV_X1 U23828 ( .A(keyinput55), .ZN(n20869) );
  NOR4_X1 U23829 ( .A1(keyinput18), .A2(keyinput66), .A3(keyinput67), .A4(
        n20869), .ZN(n20874) );
  NOR3_X1 U23830 ( .A1(keyinput79), .A2(keyinput3), .A3(keyinput96), .ZN(
        n20873) );
  NOR4_X1 U23831 ( .A1(keyinput49), .A2(keyinput68), .A3(keyinput20), .A4(
        keyinput58), .ZN(n20872) );
  NAND2_X1 U23832 ( .A1(keyinput98), .A2(keyinput57), .ZN(n20870) );
  NOR3_X1 U23833 ( .A1(keyinput15), .A2(keyinput102), .A3(n20870), .ZN(n20871)
         );
  NAND4_X1 U23834 ( .A1(n20874), .A2(n20873), .A3(n20872), .A4(n20871), .ZN(
        n20875) );
  NOR4_X1 U23835 ( .A1(keyinput108), .A2(keyinput27), .A3(n20876), .A4(n20875), 
        .ZN(n20877) );
  INV_X1 U23836 ( .A(keyinput74), .ZN(n21062) );
  NAND4_X1 U23837 ( .A1(keyinput6), .A2(n20878), .A3(n20877), .A4(n21062), 
        .ZN(n20925) );
  NOR4_X1 U23838 ( .A1(keyinput41), .A2(keyinput127), .A3(keyinput115), .A4(
        keyinput80), .ZN(n20923) );
  AND4_X1 U23839 ( .A1(keyinput43), .A2(keyinput29), .A3(keyinput22), .A4(
        keyinput60), .ZN(n20922) );
  NOR2_X1 U23840 ( .A1(keyinput39), .A2(keyinput125), .ZN(n20879) );
  NAND3_X1 U23841 ( .A1(keyinput61), .A2(keyinput76), .A3(n20879), .ZN(n20888)
         );
  INV_X1 U23842 ( .A(keyinput100), .ZN(n20880) );
  NAND4_X1 U23843 ( .A1(keyinput117), .A2(keyinput77), .A3(keyinput89), .A4(
        n20880), .ZN(n20887) );
  NOR4_X1 U23844 ( .A1(keyinput71), .A2(keyinput82), .A3(keyinput113), .A4(
        keyinput45), .ZN(n20885) );
  NAND2_X1 U23845 ( .A1(keyinput4), .A2(keyinput75), .ZN(n20881) );
  NOR3_X1 U23846 ( .A1(keyinput114), .A2(keyinput23), .A3(n20881), .ZN(n20884)
         );
  NOR4_X1 U23847 ( .A1(keyinput35), .A2(keyinput73), .A3(keyinput84), .A4(
        keyinput103), .ZN(n20883) );
  AND4_X1 U23848 ( .A1(keyinput118), .A2(keyinput11), .A3(keyinput53), .A4(
        keyinput109), .ZN(n20882) );
  NAND4_X1 U23849 ( .A1(n20885), .A2(n20884), .A3(n20883), .A4(n20882), .ZN(
        n20886) );
  NOR3_X1 U23850 ( .A1(n20888), .A2(n20887), .A3(n20886), .ZN(n20921) );
  INV_X1 U23851 ( .A(keyinput120), .ZN(n20891) );
  NOR4_X1 U23852 ( .A1(keyinput31), .A2(keyinput95), .A3(keyinput26), .A4(
        keyinput93), .ZN(n20889) );
  NAND3_X1 U23853 ( .A1(keyinput126), .A2(keyinput14), .A3(n20889), .ZN(n20890) );
  NOR3_X1 U23854 ( .A1(keyinput17), .A2(n20891), .A3(n20890), .ZN(n20903) );
  AND4_X1 U23855 ( .A1(keyinput50), .A2(keyinput86), .A3(keyinput44), .A4(
        keyinput8), .ZN(n20902) );
  NOR4_X1 U23856 ( .A1(keyinput62), .A2(keyinput78), .A3(keyinput105), .A4(
        keyinput13), .ZN(n20901) );
  INV_X1 U23857 ( .A(keyinput64), .ZN(n20892) );
  NAND4_X1 U23858 ( .A1(keyinput10), .A2(keyinput121), .A3(keyinput122), .A4(
        n20892), .ZN(n20899) );
  NOR2_X1 U23859 ( .A1(keyinput70), .A2(keyinput116), .ZN(n20893) );
  NAND3_X1 U23860 ( .A1(keyinput97), .A2(keyinput111), .A3(n20893), .ZN(n20898) );
  NOR2_X1 U23861 ( .A1(keyinput32), .A2(keyinput112), .ZN(n20894) );
  NAND3_X1 U23862 ( .A1(keyinput123), .A2(keyinput81), .A3(n20894), .ZN(n20897) );
  NOR2_X1 U23863 ( .A1(keyinput54), .A2(keyinput92), .ZN(n20895) );
  NAND3_X1 U23864 ( .A1(keyinput21), .A2(keyinput69), .A3(n20895), .ZN(n20896)
         );
  NOR4_X1 U23865 ( .A1(n20899), .A2(n20898), .A3(n20897), .A4(n20896), .ZN(
        n20900) );
  NAND4_X1 U23866 ( .A1(n20903), .A2(n20902), .A3(n20901), .A4(n20900), .ZN(
        n20919) );
  NAND4_X1 U23867 ( .A1(keyinput124), .A2(keyinput28), .A3(keyinput48), .A4(
        keyinput83), .ZN(n20918) );
  NOR2_X1 U23868 ( .A1(keyinput16), .A2(keyinput88), .ZN(n20904) );
  NAND3_X1 U23869 ( .A1(keyinput104), .A2(keyinput56), .A3(n20904), .ZN(n20917) );
  NOR2_X1 U23870 ( .A1(keyinput47), .A2(keyinput9), .ZN(n20905) );
  NAND3_X1 U23871 ( .A1(keyinput42), .A2(keyinput59), .A3(n20905), .ZN(n20906)
         );
  NOR3_X1 U23872 ( .A1(keyinput5), .A2(keyinput51), .A3(n20906), .ZN(n20915)
         );
  NOR2_X1 U23873 ( .A1(keyinput46), .A2(keyinput34), .ZN(n20907) );
  NAND3_X1 U23874 ( .A1(keyinput107), .A2(keyinput99), .A3(n20907), .ZN(n20913) );
  INV_X1 U23875 ( .A(keyinput106), .ZN(n20908) );
  NAND4_X1 U23876 ( .A1(keyinput72), .A2(keyinput65), .A3(keyinput7), .A4(
        n20908), .ZN(n20912) );
  INV_X1 U23877 ( .A(keyinput40), .ZN(n21027) );
  NAND4_X1 U23878 ( .A1(keyinput91), .A2(keyinput85), .A3(keyinput119), .A4(
        n21027), .ZN(n20911) );
  NOR2_X1 U23879 ( .A1(keyinput101), .A2(keyinput36), .ZN(n20909) );
  NAND3_X1 U23880 ( .A1(keyinput110), .A2(keyinput94), .A3(n20909), .ZN(n20910) );
  NOR4_X1 U23881 ( .A1(n20913), .A2(n20912), .A3(n20911), .A4(n20910), .ZN(
        n20914) );
  NAND4_X1 U23882 ( .A1(keyinput30), .A2(keyinput90), .A3(n20915), .A4(n20914), 
        .ZN(n20916) );
  NOR4_X1 U23883 ( .A1(n20919), .A2(n20918), .A3(n20917), .A4(n20916), .ZN(
        n20920) );
  NAND4_X1 U23884 ( .A1(n20923), .A2(n20922), .A3(n20921), .A4(n20920), .ZN(
        n20924) );
  OAI21_X1 U23885 ( .B1(n20925), .B2(n20924), .A(keyinput37), .ZN(n21194) );
  INV_X1 U23886 ( .A(keyinput80), .ZN(n20927) );
  AOI22_X1 U23887 ( .A1(n20928), .A2(keyinput117), .B1(
        P3_DATAO_REG_28__SCAN_IN), .B2(n20927), .ZN(n20926) );
  OAI221_X1 U23888 ( .B1(n20928), .B2(keyinput117), .C1(n20927), .C2(
        P3_DATAO_REG_28__SCAN_IN), .A(n20926), .ZN(n20940) );
  INV_X1 U23889 ( .A(keyinput127), .ZN(n20930) );
  AOI22_X1 U23890 ( .A1(n20931), .A2(keyinput115), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n20930), .ZN(n20929) );
  OAI221_X1 U23891 ( .B1(n20931), .B2(keyinput115), .C1(n20930), .C2(
        P1_DATAO_REG_20__SCAN_IN), .A(n20929), .ZN(n20939) );
  INV_X1 U23892 ( .A(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n20934) );
  INV_X1 U23893 ( .A(keyinput60), .ZN(n20933) );
  AOI22_X1 U23894 ( .A1(n20934), .A2(keyinput41), .B1(
        P3_DATAWIDTH_REG_4__SCAN_IN), .B2(n20933), .ZN(n20932) );
  OAI221_X1 U23895 ( .B1(n20934), .B2(keyinput41), .C1(n20933), .C2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A(n20932), .ZN(n20938) );
  XNOR2_X1 U23896 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B(keyinput22), 
        .ZN(n20936) );
  XNOR2_X1 U23897 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B(keyinput29), .ZN(
        n20935) );
  NAND2_X1 U23898 ( .A1(n20936), .A2(n20935), .ZN(n20937) );
  NOR4_X1 U23899 ( .A1(n20940), .A2(n20939), .A3(n20938), .A4(n20937), .ZN(
        n20991) );
  INV_X1 U23900 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n20942) );
  AOI22_X1 U23901 ( .A1(n20943), .A2(keyinput100), .B1(keyinput77), .B2(n20942), .ZN(n20941) );
  OAI221_X1 U23902 ( .B1(n20943), .B2(keyinput100), .C1(n20942), .C2(
        keyinput77), .A(n20941), .ZN(n20956) );
  INV_X1 U23903 ( .A(keyinput39), .ZN(n20945) );
  AOI22_X1 U23904 ( .A1(n20946), .A2(keyinput89), .B1(
        P1_DATAWIDTH_REG_11__SCAN_IN), .B2(n20945), .ZN(n20944) );
  OAI221_X1 U23905 ( .B1(n20946), .B2(keyinput89), .C1(n20945), .C2(
        P1_DATAWIDTH_REG_11__SCAN_IN), .A(n20944), .ZN(n20955) );
  INV_X1 U23906 ( .A(keyinput61), .ZN(n20948) );
  AOI22_X1 U23907 ( .A1(n20949), .A2(keyinput76), .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n20948), .ZN(n20947) );
  OAI221_X1 U23908 ( .B1(n20949), .B2(keyinput76), .C1(n20948), .C2(
        P3_CODEFETCH_REG_SCAN_IN), .A(n20947), .ZN(n20954) );
  INV_X1 U23909 ( .A(keyinput114), .ZN(n20951) );
  AOI22_X1 U23910 ( .A1(n20952), .A2(keyinput125), .B1(
        P2_DATAWIDTH_REG_12__SCAN_IN), .B2(n20951), .ZN(n20950) );
  OAI221_X1 U23911 ( .B1(n20952), .B2(keyinput125), .C1(n20951), .C2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A(n20950), .ZN(n20953) );
  NOR4_X1 U23912 ( .A1(n20956), .A2(n20955), .A3(n20954), .A4(n20953), .ZN(
        n20990) );
  INV_X1 U23913 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n20959) );
  AOI22_X1 U23914 ( .A1(n20959), .A2(keyinput75), .B1(keyinput23), .B2(n20958), 
        .ZN(n20957) );
  OAI221_X1 U23915 ( .B1(n20959), .B2(keyinput75), .C1(n20958), .C2(keyinput23), .A(n20957), .ZN(n20971) );
  INV_X1 U23916 ( .A(keyinput4), .ZN(n20961) );
  AOI22_X1 U23917 ( .A1(n20962), .A2(keyinput71), .B1(P1_LWORD_REG_5__SCAN_IN), 
        .B2(n20961), .ZN(n20960) );
  OAI221_X1 U23918 ( .B1(n20962), .B2(keyinput71), .C1(n20961), .C2(
        P1_LWORD_REG_5__SCAN_IN), .A(n20960), .ZN(n20970) );
  AOI22_X1 U23919 ( .A1(n20964), .A2(keyinput82), .B1(n13668), .B2(keyinput113), .ZN(n20963) );
  OAI221_X1 U23920 ( .B1(n20964), .B2(keyinput82), .C1(n13668), .C2(
        keyinput113), .A(n20963), .ZN(n20969) );
  AOI22_X1 U23921 ( .A1(n20967), .A2(keyinput45), .B1(n20966), .B2(keyinput118), .ZN(n20965) );
  OAI221_X1 U23922 ( .B1(n20967), .B2(keyinput45), .C1(n20966), .C2(
        keyinput118), .A(n20965), .ZN(n20968) );
  NOR4_X1 U23923 ( .A1(n20971), .A2(n20970), .A3(n20969), .A4(n20968), .ZN(
        n20989) );
  AOI22_X1 U23924 ( .A1(n20974), .A2(keyinput11), .B1(n20973), .B2(keyinput35), 
        .ZN(n20972) );
  OAI221_X1 U23925 ( .B1(n20974), .B2(keyinput11), .C1(n20973), .C2(keyinput35), .A(n20972), .ZN(n20987) );
  AOI22_X1 U23926 ( .A1(n20977), .A2(keyinput73), .B1(keyinput53), .B2(n20976), 
        .ZN(n20975) );
  OAI221_X1 U23927 ( .B1(n20977), .B2(keyinput73), .C1(n20976), .C2(keyinput53), .A(n20975), .ZN(n20986) );
  INV_X1 U23928 ( .A(DATAI_27_), .ZN(n20980) );
  INV_X1 U23929 ( .A(keyinput109), .ZN(n20979) );
  AOI22_X1 U23930 ( .A1(n20980), .A2(keyinput84), .B1(P3_UWORD_REG_5__SCAN_IN), 
        .B2(n20979), .ZN(n20978) );
  OAI221_X1 U23931 ( .B1(n20980), .B2(keyinput84), .C1(n20979), .C2(
        P3_UWORD_REG_5__SCAN_IN), .A(n20978), .ZN(n20985) );
  INV_X1 U23932 ( .A(keyinput16), .ZN(n20982) );
  AOI22_X1 U23933 ( .A1(n20983), .A2(keyinput103), .B1(
        P3_ADDRESS_REG_2__SCAN_IN), .B2(n20982), .ZN(n20981) );
  OAI221_X1 U23934 ( .B1(n20983), .B2(keyinput103), .C1(n20982), .C2(
        P3_ADDRESS_REG_2__SCAN_IN), .A(n20981), .ZN(n20984) );
  NOR4_X1 U23935 ( .A1(n20987), .A2(n20986), .A3(n20985), .A4(n20984), .ZN(
        n20988) );
  NAND4_X1 U23936 ( .A1(n20991), .A2(n20990), .A3(n20989), .A4(n20988), .ZN(
        n21193) );
  AOI22_X1 U23937 ( .A1(n20993), .A2(keyinput104), .B1(n9982), .B2(keyinput56), 
        .ZN(n20992) );
  OAI221_X1 U23938 ( .B1(n20993), .B2(keyinput104), .C1(n9982), .C2(keyinput56), .A(n20992), .ZN(n21006) );
  INV_X1 U23939 ( .A(keyinput124), .ZN(n20995) );
  AOI22_X1 U23940 ( .A1(n20996), .A2(keyinput88), .B1(P1_UWORD_REG_11__SCAN_IN), .B2(n20995), .ZN(n20994) );
  OAI221_X1 U23941 ( .B1(n20996), .B2(keyinput88), .C1(n20995), .C2(
        P1_UWORD_REG_11__SCAN_IN), .A(n20994), .ZN(n21005) );
  INV_X1 U23942 ( .A(keyinput48), .ZN(n20998) );
  AOI22_X1 U23943 ( .A1(n20999), .A2(keyinput28), .B1(P1_DATAO_REG_8__SCAN_IN), 
        .B2(n20998), .ZN(n20997) );
  OAI221_X1 U23944 ( .B1(n20999), .B2(keyinput28), .C1(n20998), .C2(
        P1_DATAO_REG_8__SCAN_IN), .A(n20997), .ZN(n21004) );
  INV_X1 U23945 ( .A(keyinput65), .ZN(n21001) );
  AOI22_X1 U23946 ( .A1(n21002), .A2(keyinput83), .B1(P2_LWORD_REG_13__SCAN_IN), .B2(n21001), .ZN(n21000) );
  OAI221_X1 U23947 ( .B1(n21002), .B2(keyinput83), .C1(n21001), .C2(
        P2_LWORD_REG_13__SCAN_IN), .A(n21000), .ZN(n21003) );
  NOR4_X1 U23948 ( .A1(n21006), .A2(n21005), .A3(n21004), .A4(n21003), .ZN(
        n21191) );
  AOI22_X1 U23949 ( .A1(n21008), .A2(keyinput72), .B1(n9983), .B2(keyinput106), 
        .ZN(n21007) );
  OAI221_X1 U23950 ( .B1(n21008), .B2(keyinput72), .C1(n9983), .C2(keyinput106), .A(n21007), .ZN(n21020) );
  INV_X1 U23951 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n21011) );
  INV_X1 U23952 ( .A(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n21010) );
  AOI22_X1 U23953 ( .A1(n21011), .A2(keyinput7), .B1(keyinput107), .B2(n21010), 
        .ZN(n21009) );
  OAI221_X1 U23954 ( .B1(n21011), .B2(keyinput7), .C1(n21010), .C2(keyinput107), .A(n21009), .ZN(n21019) );
  AOI22_X1 U23955 ( .A1(n21014), .A2(keyinput46), .B1(n21013), .B2(keyinput99), 
        .ZN(n21012) );
  OAI221_X1 U23956 ( .B1(n21014), .B2(keyinput46), .C1(n21013), .C2(keyinput99), .A(n21012), .ZN(n21018) );
  AOI22_X1 U23957 ( .A1(n21016), .A2(keyinput34), .B1(n10896), .B2(keyinput101), .ZN(n21015) );
  OAI221_X1 U23958 ( .B1(n21016), .B2(keyinput34), .C1(n10896), .C2(
        keyinput101), .A(n21015), .ZN(n21017) );
  NOR4_X1 U23959 ( .A1(n21020), .A2(n21019), .A3(n21018), .A4(n21017), .ZN(
        n21190) );
  INV_X1 U23960 ( .A(keyinput110), .ZN(n21023) );
  INV_X1 U23961 ( .A(keyinput94), .ZN(n21022) );
  AOI22_X1 U23962 ( .A1(n21023), .A2(P3_DATAO_REG_0__SCAN_IN), .B1(
        P3_ADDRESS_REG_7__SCAN_IN), .B2(n21022), .ZN(n21021) );
  OAI221_X1 U23963 ( .B1(n21023), .B2(P3_DATAO_REG_0__SCAN_IN), .C1(n21022), 
        .C2(P3_ADDRESS_REG_7__SCAN_IN), .A(n21021), .ZN(n21054) );
  INV_X1 U23964 ( .A(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n21026) );
  INV_X1 U23965 ( .A(keyinput85), .ZN(n21025) );
  AOI22_X1 U23966 ( .A1(n21026), .A2(keyinput36), .B1(P2_DATAO_REG_24__SCAN_IN), .B2(n21025), .ZN(n21024) );
  OAI221_X1 U23967 ( .B1(n21026), .B2(keyinput36), .C1(n21025), .C2(
        P2_DATAO_REG_24__SCAN_IN), .A(n21024), .ZN(n21053) );
  XNOR2_X1 U23968 ( .A(n21027), .B(P3_DATAWIDTH_REG_17__SCAN_IN), .ZN(n21032)
         );
  INV_X1 U23969 ( .A(keyinput91), .ZN(n21029) );
  AOI22_X1 U23970 ( .A1(n21030), .A2(keyinput119), .B1(
        P3_DATAWIDTH_REG_21__SCAN_IN), .B2(n21029), .ZN(n21028) );
  OAI221_X1 U23971 ( .B1(n21030), .B2(keyinput119), .C1(n21029), .C2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A(n21028), .ZN(n21031) );
  AOI211_X1 U23972 ( .C1(n21034), .C2(keyinput30), .A(n21032), .B(n21031), 
        .ZN(n21033) );
  OAI21_X1 U23973 ( .B1(n21034), .B2(keyinput30), .A(n21033), .ZN(n21052) );
  INV_X1 U23974 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n21037) );
  INV_X1 U23975 ( .A(keyinput90), .ZN(n21036) );
  OAI22_X1 U23976 ( .A1(n21037), .A2(keyinput5), .B1(n21036), .B2(
        P3_EAX_REG_18__SCAN_IN), .ZN(n21035) );
  AOI221_X1 U23977 ( .B1(n21037), .B2(keyinput5), .C1(P3_EAX_REG_18__SCAN_IN), 
        .C2(n21036), .A(n21035), .ZN(n21050) );
  INV_X1 U23978 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n21040) );
  INV_X1 U23979 ( .A(keyinput42), .ZN(n21039) );
  OAI22_X1 U23980 ( .A1(n21040), .A2(keyinput51), .B1(n21039), .B2(
        P2_UWORD_REG_3__SCAN_IN), .ZN(n21038) );
  AOI221_X1 U23981 ( .B1(n21040), .B2(keyinput51), .C1(P2_UWORD_REG_3__SCAN_IN), .C2(n21039), .A(n21038), .ZN(n21049) );
  INV_X1 U23982 ( .A(keyinput59), .ZN(n21042) );
  OAI22_X1 U23983 ( .A1(n21043), .A2(keyinput47), .B1(n21042), .B2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(n21041) );
  AOI221_X1 U23984 ( .B1(n21043), .B2(keyinput47), .C1(
        P1_DATAWIDTH_REG_13__SCAN_IN), .C2(n21042), .A(n21041), .ZN(n21048) );
  OAI22_X1 U23985 ( .A1(keyinput79), .A2(n21046), .B1(n21045), .B2(keyinput9), 
        .ZN(n21044) );
  AOI221_X1 U23986 ( .B1(n21046), .B2(keyinput79), .C1(n21045), .C2(keyinput9), 
        .A(n21044), .ZN(n21047) );
  NAND4_X1 U23987 ( .A1(n21050), .A2(n21049), .A3(n21048), .A4(n21047), .ZN(
        n21051) );
  NOR4_X1 U23988 ( .A1(n21054), .A2(n21053), .A3(n21052), .A4(n21051), .ZN(
        n21189) );
  INV_X1 U23989 ( .A(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n21056) );
  XNOR2_X1 U23990 ( .A(n11027), .B(keyinput3), .ZN(n21055) );
  AOI21_X1 U23991 ( .B1(keyinput37), .B2(n21056), .A(n21055), .ZN(n21059) );
  XNOR2_X1 U23992 ( .A(keyinput67), .B(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n21058) );
  XNOR2_X1 U23993 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(keyinput66), 
        .ZN(n21057) );
  NAND3_X1 U23994 ( .A1(n21059), .A2(n21058), .A3(n21057), .ZN(n21066) );
  INV_X1 U23995 ( .A(keyinput19), .ZN(n21061) );
  AOI22_X1 U23996 ( .A1(n21062), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n21061), .ZN(n21060) );
  OAI221_X1 U23997 ( .B1(n21062), .B2(P2_DATAO_REG_21__SCAN_IN), .C1(n21061), 
        .C2(P2_DATAO_REG_4__SCAN_IN), .A(n21060), .ZN(n21065) );
  XNOR2_X1 U23998 ( .A(n21063), .B(keyinput18), .ZN(n21064) );
  NOR3_X1 U23999 ( .A1(n21066), .A2(n21065), .A3(n21064), .ZN(n21086) );
  INV_X1 U24000 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21068) );
  OAI22_X1 U24001 ( .A1(n21069), .A2(keyinput25), .B1(n21068), .B2(keyinput38), 
        .ZN(n21067) );
  AOI221_X1 U24002 ( .B1(n21069), .B2(keyinput25), .C1(keyinput38), .C2(n21068), .A(n21067), .ZN(n21085) );
  INV_X1 U24003 ( .A(keyinput15), .ZN(n21071) );
  OAI22_X1 U24004 ( .A1(keyinput52), .A2(n21072), .B1(n21071), .B2(
        P3_DATAO_REG_27__SCAN_IN), .ZN(n21070) );
  AOI221_X1 U24005 ( .B1(n21072), .B2(keyinput52), .C1(n21071), .C2(
        P3_DATAO_REG_27__SCAN_IN), .A(n21070), .ZN(n21084) );
  AOI22_X1 U24006 ( .A1(n21075), .A2(keyinput55), .B1(n21074), .B2(keyinput33), 
        .ZN(n21073) );
  OAI221_X1 U24007 ( .B1(n21075), .B2(keyinput55), .C1(n21074), .C2(keyinput33), .A(n21073), .ZN(n21082) );
  INV_X1 U24008 ( .A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n21078) );
  AOI22_X1 U24009 ( .A1(n21078), .A2(keyinput2), .B1(n21077), .B2(keyinput6), 
        .ZN(n21076) );
  OAI221_X1 U24010 ( .B1(n21078), .B2(keyinput2), .C1(n21077), .C2(keyinput6), 
        .A(n21076), .ZN(n21081) );
  XNOR2_X1 U24011 ( .A(n21079), .B(keyinput96), .ZN(n21080) );
  NOR3_X1 U24012 ( .A1(n21082), .A2(n21081), .A3(n21080), .ZN(n21083) );
  NAND4_X1 U24013 ( .A1(n21086), .A2(n21085), .A3(n21084), .A4(n21083), .ZN(
        n21187) );
  INV_X1 U24014 ( .A(keyinput105), .ZN(n21088) );
  OAI22_X1 U24015 ( .A1(keyinput86), .A2(n21089), .B1(n21088), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n21087) );
  AOI221_X1 U24016 ( .B1(n21089), .B2(keyinput86), .C1(n21088), .C2(
        P2_DATAO_REG_17__SCAN_IN), .A(n21087), .ZN(n21102) );
  INV_X1 U24017 ( .A(keyinput78), .ZN(n21091) );
  OAI22_X1 U24018 ( .A1(n21092), .A2(keyinput50), .B1(n21091), .B2(
        P3_BE_N_REG_0__SCAN_IN), .ZN(n21090) );
  AOI221_X1 U24019 ( .B1(n21092), .B2(keyinput50), .C1(P3_BE_N_REG_0__SCAN_IN), 
        .C2(n21091), .A(n21090), .ZN(n21101) );
  INV_X1 U24020 ( .A(keyinput44), .ZN(n21094) );
  OAI22_X1 U24021 ( .A1(n21095), .A2(keyinput70), .B1(n21094), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n21093) );
  AOI221_X1 U24022 ( .B1(n21095), .B2(keyinput70), .C1(P1_EBX_REG_13__SCAN_IN), 
        .C2(n21094), .A(n21093), .ZN(n21100) );
  OAI22_X1 U24023 ( .A1(n21098), .A2(keyinput13), .B1(n21097), .B2(keyinput8), 
        .ZN(n21096) );
  AOI221_X1 U24024 ( .B1(n21098), .B2(keyinput13), .C1(keyinput8), .C2(n21097), 
        .A(n21096), .ZN(n21099) );
  NAND4_X1 U24025 ( .A1(n21102), .A2(n21101), .A3(n21100), .A4(n21099), .ZN(
        n21186) );
  INV_X1 U24026 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n21105) );
  INV_X1 U24027 ( .A(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n21104) );
  OAI22_X1 U24028 ( .A1(n21105), .A2(keyinput31), .B1(n21104), .B2(keyinput126), .ZN(n21103) );
  AOI221_X1 U24029 ( .B1(n21105), .B2(keyinput31), .C1(keyinput126), .C2(
        n21104), .A(n21103), .ZN(n21117) );
  INV_X1 U24030 ( .A(keyinput95), .ZN(n21107) );
  OAI22_X1 U24031 ( .A1(n9986), .A2(keyinput17), .B1(n21107), .B2(
        P2_DATAO_REG_22__SCAN_IN), .ZN(n21106) );
  AOI221_X1 U24032 ( .B1(n9986), .B2(keyinput17), .C1(P2_DATAO_REG_22__SCAN_IN), .C2(n21107), .A(n21106), .ZN(n21116) );
  INV_X1 U24033 ( .A(keyinput26), .ZN(n21109) );
  OAI22_X1 U24034 ( .A1(n21110), .A2(keyinput62), .B1(n21109), .B2(
        P3_LWORD_REG_6__SCAN_IN), .ZN(n21108) );
  AOI221_X1 U24035 ( .B1(n21110), .B2(keyinput62), .C1(P3_LWORD_REG_6__SCAN_IN), .C2(n21109), .A(n21108), .ZN(n21115) );
  OAI22_X1 U24036 ( .A1(n21113), .A2(keyinput14), .B1(n21112), .B2(keyinput93), 
        .ZN(n21111) );
  AOI221_X1 U24037 ( .B1(n21113), .B2(keyinput14), .C1(keyinput93), .C2(n21112), .A(n21111), .ZN(n21114) );
  NAND4_X1 U24038 ( .A1(n21117), .A2(n21116), .A3(n21115), .A4(n21114), .ZN(
        n21185) );
  AOI22_X1 U24039 ( .A1(n21120), .A2(keyinput63), .B1(n21119), .B2(keyinput108), .ZN(n21118) );
  OAI221_X1 U24040 ( .B1(n21120), .B2(keyinput63), .C1(n21119), .C2(
        keyinput108), .A(n21118), .ZN(n21132) );
  INV_X1 U24041 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n21123) );
  AOI22_X1 U24042 ( .A1(n21123), .A2(keyinput12), .B1(keyinput0), .B2(n21122), 
        .ZN(n21121) );
  OAI221_X1 U24043 ( .B1(n21123), .B2(keyinput12), .C1(n21122), .C2(keyinput0), 
        .A(n21121), .ZN(n21131) );
  AOI22_X1 U24044 ( .A1(n13776), .A2(keyinput87), .B1(keyinput120), .B2(n21125), .ZN(n21124) );
  OAI221_X1 U24045 ( .B1(n13776), .B2(keyinput87), .C1(n21125), .C2(
        keyinput120), .A(n21124), .ZN(n21130) );
  INV_X1 U24046 ( .A(keyinput24), .ZN(n21127) );
  AOI22_X1 U24047 ( .A1(n21128), .A2(keyinput27), .B1(P3_DATAO_REG_24__SCAN_IN), .B2(n21127), .ZN(n21126) );
  OAI221_X1 U24048 ( .B1(n21128), .B2(keyinput27), .C1(n21127), .C2(
        P3_DATAO_REG_24__SCAN_IN), .A(n21126), .ZN(n21129) );
  NOR4_X1 U24049 ( .A1(n21132), .A2(n21131), .A3(n21130), .A4(n21129), .ZN(
        n21183) );
  INV_X1 U24050 ( .A(DATAI_2_), .ZN(n21135) );
  INV_X1 U24051 ( .A(keyinput68), .ZN(n21134) );
  AOI22_X1 U24052 ( .A1(n21135), .A2(keyinput20), .B1(P1_D_C_N_REG_SCAN_IN), 
        .B2(n21134), .ZN(n21133) );
  OAI221_X1 U24053 ( .B1(n21135), .B2(keyinput20), .C1(n21134), .C2(
        P1_D_C_N_REG_SCAN_IN), .A(n21133), .ZN(n21148) );
  AOI22_X1 U24054 ( .A1(n21138), .A2(keyinput57), .B1(n21137), .B2(keyinput49), 
        .ZN(n21136) );
  OAI221_X1 U24055 ( .B1(n21138), .B2(keyinput57), .C1(n21137), .C2(keyinput49), .A(n21136), .ZN(n21147) );
  INV_X1 U24056 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n21140) );
  AOI22_X1 U24057 ( .A1(n21141), .A2(keyinput98), .B1(n21140), .B2(keyinput1), 
        .ZN(n21139) );
  OAI221_X1 U24058 ( .B1(n21141), .B2(keyinput98), .C1(n21140), .C2(keyinput1), 
        .A(n21139), .ZN(n21146) );
  AOI22_X1 U24059 ( .A1(n21144), .A2(keyinput58), .B1(keyinput102), .B2(n21143), .ZN(n21142) );
  OAI221_X1 U24060 ( .B1(n21144), .B2(keyinput58), .C1(n21143), .C2(
        keyinput102), .A(n21142), .ZN(n21145) );
  NOR4_X1 U24061 ( .A1(n21148), .A2(n21147), .A3(n21146), .A4(n21145), .ZN(
        n21182) );
  INV_X1 U24062 ( .A(keyinput69), .ZN(n21151) );
  INV_X1 U24063 ( .A(keyinput123), .ZN(n21150) );
  AOI22_X1 U24064 ( .A1(n21151), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(
        P3_DATAWIDTH_REG_11__SCAN_IN), .B2(n21150), .ZN(n21149) );
  OAI221_X1 U24065 ( .B1(n21151), .B2(P3_LWORD_REG_7__SCAN_IN), .C1(n21150), 
        .C2(P3_DATAWIDTH_REG_11__SCAN_IN), .A(n21149), .ZN(n21164) );
  AOI22_X1 U24066 ( .A1(n21154), .A2(keyinput21), .B1(n21153), .B2(keyinput92), 
        .ZN(n21152) );
  OAI221_X1 U24067 ( .B1(n21154), .B2(keyinput21), .C1(n21153), .C2(keyinput92), .A(n21152), .ZN(n21163) );
  INV_X1 U24068 ( .A(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n21156) );
  AOI22_X1 U24069 ( .A1(n21157), .A2(keyinput81), .B1(keyinput43), .B2(n21156), 
        .ZN(n21155) );
  OAI221_X1 U24070 ( .B1(n21157), .B2(keyinput81), .C1(n21156), .C2(keyinput43), .A(n21155), .ZN(n21162) );
  INV_X1 U24071 ( .A(keyinput112), .ZN(n21160) );
  INV_X1 U24072 ( .A(keyinput32), .ZN(n21159) );
  AOI22_X1 U24073 ( .A1(n21160), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n21159), .ZN(n21158) );
  OAI221_X1 U24074 ( .B1(n21160), .B2(P3_UWORD_REG_7__SCAN_IN), .C1(n21159), 
        .C2(P1_DATAO_REG_30__SCAN_IN), .A(n21158), .ZN(n21161) );
  NOR4_X1 U24075 ( .A1(n21164), .A2(n21163), .A3(n21162), .A4(n21161), .ZN(
        n21181) );
  AOI22_X1 U24076 ( .A1(n21167), .A2(keyinput116), .B1(n21166), .B2(
        keyinput121), .ZN(n21165) );
  OAI221_X1 U24077 ( .B1(n21167), .B2(keyinput116), .C1(n21166), .C2(
        keyinput121), .A(n21165), .ZN(n21179) );
  AOI22_X1 U24078 ( .A1(n21170), .A2(keyinput97), .B1(keyinput111), .B2(n21169), .ZN(n21168) );
  OAI221_X1 U24079 ( .B1(n21170), .B2(keyinput97), .C1(n21169), .C2(
        keyinput111), .A(n21168), .ZN(n21178) );
  INV_X1 U24080 ( .A(keyinput54), .ZN(n21172) );
  AOI22_X1 U24081 ( .A1(n11382), .A2(keyinput64), .B1(P2_DATAO_REG_27__SCAN_IN), .B2(n21172), .ZN(n21171) );
  OAI221_X1 U24082 ( .B1(n11382), .B2(keyinput64), .C1(n21172), .C2(
        P2_DATAO_REG_27__SCAN_IN), .A(n21171), .ZN(n21177) );
  INV_X1 U24083 ( .A(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n21175) );
  INV_X1 U24084 ( .A(keyinput122), .ZN(n21174) );
  AOI22_X1 U24085 ( .A1(n21175), .A2(keyinput10), .B1(P1_UWORD_REG_10__SCAN_IN), .B2(n21174), .ZN(n21173) );
  OAI221_X1 U24086 ( .B1(n21175), .B2(keyinput10), .C1(n21174), .C2(
        P1_UWORD_REG_10__SCAN_IN), .A(n21173), .ZN(n21176) );
  NOR4_X1 U24087 ( .A1(n21179), .A2(n21178), .A3(n21177), .A4(n21176), .ZN(
        n21180) );
  NAND4_X1 U24088 ( .A1(n21183), .A2(n21182), .A3(n21181), .A4(n21180), .ZN(
        n21184) );
  NOR4_X1 U24089 ( .A1(n21187), .A2(n21186), .A3(n21185), .A4(n21184), .ZN(
        n21188) );
  NAND4_X1 U24090 ( .A1(n21191), .A2(n21190), .A3(n21189), .A4(n21188), .ZN(
        n21192) );
  AOI211_X1 U24091 ( .C1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .C2(n21194), .A(
        n21193), .B(n21192), .ZN(n21207) );
  AOI22_X1 U24092 ( .A1(n21198), .A2(n21197), .B1(n21196), .B2(n21195), .ZN(
        n21203) );
  AOI22_X1 U24093 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n21201), .B1(
        n21200), .B2(n21199), .ZN(n21202) );
  OAI211_X1 U24094 ( .C1(n21205), .C2(n21204), .A(n21203), .B(n21202), .ZN(
        n21206) );
  XOR2_X1 U24095 ( .A(n21207), .B(n21206), .Z(P1_U3105) );
  INV_X1 U11206 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18793) );
  NAND2_X1 U11227 ( .A1(n11508), .A2(n11507), .ZN(n14077) );
  AND2_X2 U11277 ( .A1(n13880), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13647) );
  BUF_X2 U11192 ( .A(n15736), .Z(n9724) );
  CLKBUF_X2 U11249 ( .A(n11799), .Z(n9751) );
  INV_X1 U11250 ( .A(n15645), .ZN(n15694) );
  NAND2_X1 U11272 ( .A1(n20189), .A2(n12974), .ZN(n12623) );
  CLKBUF_X1 U11273 ( .A(n10473), .Z(n10480) );
  NAND3_X1 U11294 ( .A1(n9857), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14341), .ZN(n14323) );
  CLKBUF_X1 U11323 ( .A(n11139), .Z(n13000) );
  CLKBUF_X1 U11393 ( .A(n13170), .Z(n9741) );
  CLKBUF_X1 U11454 ( .A(n12426), .Z(n13405) );
  CLKBUF_X1 U11464 ( .A(n15847), .Z(n9725) );
  CLKBUF_X1 U11521 ( .A(n16484), .Z(n16487) );
  CLKBUF_X1 U11522 ( .A(n17476), .Z(n17480) );
endmodule

