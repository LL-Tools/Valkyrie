

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297;

  OR2_X1 U4906 ( .A1(n9285), .A2(n9265), .ZN(n9263) );
  NAND2_X1 U4907 ( .A1(n7404), .A2(n7307), .ZN(n9871) );
  NAND2_X1 U4908 ( .A1(n5990), .A2(n9492), .ZN(n6261) );
  INV_X1 U4910 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U4911 ( .A(n7842), .ZN(n5031) );
  INV_X1 U4912 ( .A(n5782), .ZN(n5638) );
  OR2_X1 U4913 ( .A1(n8472), .A2(n5930), .ZN(n8473) );
  OAI21_X1 U4914 ( .B1(n8041), .B2(n5577), .A(n5576), .ZN(n5589) );
  INV_X1 U4915 ( .A(n7941), .ZN(n7983) );
  AOI21_X1 U4916 ( .B1(n9141), .B2(n9147), .A(n6326), .ZN(n6337) );
  OR2_X1 U4917 ( .A1(n9166), .A2(n9183), .ZN(n9164) );
  NAND2_X1 U4918 ( .A1(n6498), .A2(n6428), .ZN(n8772) );
  INV_X1 U4919 ( .A(n8845), .ZN(n9763) );
  INV_X1 U4920 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6121) );
  XNOR2_X1 U4921 ( .A(n5667), .B(P2_IR_REG_22__SCAN_IN), .ZN(n5689) );
  OAI211_X2 U4922 ( .C1(n8772), .C2(n6436), .A(n6062), .B(n6061), .ZN(n9700)
         );
  XNOR2_X1 U4923 ( .A(n6347), .B(n6346), .ZN(n6356) );
  INV_X1 U4924 ( .A(n7451), .ZN(n5050) );
  INV_X1 U4925 ( .A(n7027), .ZN(n9779) );
  BUF_X1 U4926 ( .A(n6561), .Z(n9215) );
  NAND2_X2 U4927 ( .A1(n8302), .A2(n8308), .ZN(n8301) );
  NOR2_X4 U4928 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6077) );
  OAI21_X2 U4929 ( .B1(n8390), .B2(n4758), .A(n4755), .ZN(n8354) );
  NAND2_X2 U4930 ( .A1(n8408), .A2(n5731), .ZN(n8390) );
  NAND2_X2 U4931 ( .A1(n4965), .A2(n4966), .ZN(n8365) );
  OR2_X2 U4932 ( .A1(n6765), .A2(n6764), .ZN(n6981) );
  NAND2_X2 U4933 ( .A1(n6000), .A2(n6003), .ZN(n6372) );
  INV_X1 U4934 ( .A(n6261), .ZN(n4403) );
  INV_X2 U4935 ( .A(n6261), .ZN(n6097) );
  AND2_X4 U4936 ( .A1(n4555), .A2(n4554), .ZN(n5061) );
  OAI222_X1 U4937 ( .A1(n5030), .A2(n8130), .B1(n8025), .B2(n9490), .C1(n8651), 
        .C2(n5762), .ZN(P2_U3328) );
  INV_X1 U4938 ( .A(n5030), .ZN(n5029) );
  NAND2_X1 U4939 ( .A1(n6134), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6062) );
  OAI21_X2 U4940 ( .B1(n9305), .B2(n9317), .A(n9299), .ZN(n9277) );
  OAI21_X2 U4941 ( .B1(n5044), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5667) );
  OAI21_X2 U4942 ( .B1(n8752), .B2(n8755), .A(n8753), .ZN(n8689) );
  NAND2_X1 U4943 ( .A1(n8682), .A2(n8680), .ZN(n4635) );
  MUX2_X1 U4944 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n6420), .S(n9809), .Z(n6417)
         );
  MUX2_X1 U4945 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n6420), .S(n10189), .Z(n6421) );
  OAI21_X1 U4946 ( .B1(n9192), .B2(n4445), .A(n4924), .ZN(n4923) );
  NAND2_X1 U4947 ( .A1(n5723), .A2(n5936), .ZN(n7338) );
  NAND2_X1 U4948 ( .A1(n6143), .A2(n6142), .ZN(n9796) );
  NAND2_X1 U4949 ( .A1(n6667), .A2(n7408), .ZN(n6677) );
  NAND2_X2 U4950 ( .A1(n7409), .A2(n7981), .ZN(n6675) );
  INV_X2 U4951 ( .A(n7890), .ZN(n7981) );
  INV_X1 U4952 ( .A(n8949), .ZN(n8944) );
  OAI211_X1 U4953 ( .C1(n6739), .C2(n8192), .A(n5094), .B(n5093), .ZN(n8545)
         );
  INV_X1 U4954 ( .A(n9748), .ZN(n9734) );
  NAND4_X2 U4955 ( .A1(n6076), .A2(n6075), .A3(n6074), .A4(n6073), .ZN(n6589)
         );
  NAND2_X1 U4956 ( .A1(n6739), .A2(n5061), .ZN(n5106) );
  BUF_X2 U4957 ( .A(n6100), .Z(n6374) );
  NAND2_X2 U4958 ( .A1(n6372), .A2(n9047), .ZN(n6498) );
  MUX2_X1 U4959 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5054), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5056) );
  AND2_X1 U4960 ( .A1(n5052), .A2(n5021), .ZN(n5024) );
  AND4_X1 U4961 ( .A1(n4991), .A2(n5019), .A3(n5145), .A4(n4463), .ZN(n5052)
         );
  INV_X8 U4962 ( .A(n5061), .ZN(n6428) );
  INV_X2 U4963 ( .A(P2_STATE_REG_SCAN_IN), .ZN(n8130) );
  OAI21_X1 U4964 ( .B1(n5968), .B2(n5967), .A(n7540), .ZN(n5973) );
  AND2_X1 U4965 ( .A1(n5786), .A2(n5785), .ZN(n5968) );
  NAND2_X1 U4966 ( .A1(n4635), .A2(n4634), .ZN(n8745) );
  OR2_X1 U4967 ( .A1(n5692), .A2(n5691), .ZN(n5693) );
  AOI211_X1 U4968 ( .C1(n8565), .C2(n8520), .A(n8313), .B(n8312), .ZN(n8314)
         );
  OAI21_X1 U4969 ( .B1(n8285), .B2(n8284), .A(n9843), .ZN(n8291) );
  NAND2_X1 U4970 ( .A1(n4889), .A2(n4888), .ZN(n4887) );
  NAND2_X1 U4971 ( .A1(n8953), .A2(n9013), .ZN(n4888) );
  INV_X1 U4972 ( .A(n8952), .ZN(n4889) );
  NAND3_X1 U4973 ( .A1(n7943), .A2(n4871), .A3(n4872), .ZN(n8705) );
  NAND2_X1 U4974 ( .A1(n4599), .A2(n4598), .ZN(n8953) );
  AOI21_X1 U4975 ( .B1(n4770), .B2(n9843), .A(n4767), .ZN(n8567) );
  NAND2_X1 U4976 ( .A1(n4602), .A2(n4600), .ZN(n4599) );
  OR2_X1 U4977 ( .A1(n8945), .A2(n4603), .ZN(n4602) );
  INV_X1 U4978 ( .A(n4923), .ZN(n9141) );
  NAND2_X1 U4979 ( .A1(n8442), .A2(n4995), .ZN(n8420) );
  INV_X1 U4980 ( .A(n8708), .ZN(n4872) );
  AND2_X1 U4981 ( .A1(n8505), .A2(n8504), .ZN(n8507) );
  NOR2_X1 U4982 ( .A1(n8113), .A2(n4794), .ZN(n4793) );
  INV_X1 U4983 ( .A(n9340), .ZN(n4700) );
  OR2_X1 U4984 ( .A1(n7776), .A2(n8768), .ZN(n9340) );
  AOI21_X1 U4985 ( .B1(n7132), .B2(n4835), .A(n4834), .ZN(n4833) );
  INV_X2 U4986 ( .A(n8549), .ZN(n9860) );
  NAND2_X1 U4987 ( .A1(n5351), .A2(n5350), .ZN(n9525) );
  INV_X1 U4988 ( .A(n9769), .ZN(n6988) );
  CLKBUF_X1 U4989 ( .A(n8730), .Z(n8767) );
  NAND2_X1 U4990 ( .A1(n6137), .A2(n6136), .ZN(n7124) );
  NAND2_X1 U4991 ( .A1(n6125), .A2(n6124), .ZN(n9769) );
  XNOR2_X1 U4992 ( .A(n6579), .B(n6972), .ZN(n6629) );
  NAND2_X1 U4993 ( .A1(n5214), .A2(n5213), .ZN(n5227) );
  XNOR2_X1 U4994 ( .A(n5196), .B(n5195), .ZN(n6441) );
  NAND2_X1 U4995 ( .A1(n4533), .A2(n4879), .ZN(n5211) );
  INV_X1 U4996 ( .A(n7986), .ZN(n6972) );
  OAI211_X1 U4997 ( .C1(n6438), .C2(n8772), .A(n6053), .B(n4686), .ZN(n8845)
         );
  AND2_X2 U4998 ( .A1(n6558), .A2(n6557), .ZN(n5005) );
  AND3_X1 U4999 ( .A1(n6082), .A2(n4808), .A3(n4805), .ZN(n9732) );
  AND3_X1 U5000 ( .A1(n6118), .A2(n6117), .A3(n4532), .ZN(n7027) );
  NAND4_X1 U5001 ( .A1(n6105), .A2(n6104), .A3(n6103), .A4(n6102), .ZN(n9044)
         );
  INV_X2 U5002 ( .A(n5106), .ZN(n5764) );
  NAND2_X1 U5003 ( .A1(n5049), .A2(n5048), .ZN(n7451) );
  AND4_X1 U5004 ( .A1(n6049), .A2(n6048), .A3(n6050), .A4(n4619), .ZN(n6896)
         );
  XNOR2_X1 U5005 ( .A(n5039), .B(n5040), .ZN(n7310) );
  AND4_X1 U5006 ( .A1(n5126), .A2(n5125), .A3(n5124), .A4(n5123), .ZN(n7868)
         );
  OAI211_X1 U5007 ( .C1(n8772), .C2(n6430), .A(n6095), .B(n6094), .ZN(n6707)
         );
  AND2_X2 U5008 ( .A1(n6501), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  AND4_X1 U5009 ( .A1(n5101), .A2(n5100), .A3(n5099), .A4(n5098), .ZN(n6956)
         );
  NAND4_X2 U5010 ( .A1(n6092), .A2(n6091), .A3(n6090), .A4(n6089), .ZN(n9748)
         );
  INV_X2 U5011 ( .A(n8772), .ZN(n8780) );
  AND2_X2 U5012 ( .A1(n5029), .A2(n7842), .ZN(n4430) );
  INV_X2 U5013 ( .A(n6498), .ZN(n6243) );
  NAND2_X1 U5014 ( .A1(n6389), .A2(n6397), .ZN(n6558) );
  INV_X1 U5015 ( .A(n5689), .ZN(n7404) );
  XNOR2_X1 U5016 ( .A(n5045), .B(n4499), .ZN(n7307) );
  CLKBUF_X3 U5017 ( .A(n6098), .Z(n6313) );
  CLKBUF_X1 U5018 ( .A(n5705), .Z(n8646) );
  NAND2_X1 U5019 ( .A1(n5023), .A2(n5028), .ZN(n7842) );
  NAND2_X1 U5020 ( .A1(n6006), .A2(n6001), .ZN(n9047) );
  NOR2_X2 U5021 ( .A1(n6023), .A2(n6015), .ZN(n6344) );
  INV_X1 U5022 ( .A(n5226), .ZN(n4404) );
  NAND2_X1 U5023 ( .A1(n5027), .A2(n5026), .ZN(n5028) );
  MUX2_X1 U5024 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6005), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n6006) );
  MUX2_X1 U5025 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6002), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n6003) );
  AOI21_X1 U5026 ( .B1(n6000), .B2(n4439), .A(n4605), .ZN(n4604) );
  OR2_X1 U5027 ( .A1(n5989), .A2(n6121), .ZN(n5988) );
  AND2_X1 U5028 ( .A1(n5987), .A2(n4461), .ZN(n5989) );
  NAND2_X2 U5029 ( .A1(n6428), .A2(P1_U3084), .ZN(n9494) );
  NAND2_X2 U5030 ( .A1(n5061), .A2(n8130), .ZN(n8025) );
  NAND2_X1 U5031 ( .A1(n4804), .A2(n5037), .ZN(n4803) );
  NAND2_X1 U5032 ( .A1(n5020), .A2(n4763), .ZN(n4762) );
  NAND2_X1 U5033 ( .A1(n5025), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5026) );
  INV_X4 U5034 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U5035 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n4722) );
  NOR2_X1 U5036 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4723) );
  NOR2_X1 U5037 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4641) );
  NOR2_X1 U5038 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4501) );
  INV_X1 U5039 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5009) );
  NOR2_X1 U5040 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n4605) );
  INV_X1 U5041 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5666) );
  INV_X1 U5042 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5373) );
  NOR2_X2 U5043 ( .A1(n7158), .A2(n7233), .ZN(n7379) );
  NOR2_X2 U5044 ( .A1(n9545), .A2(n4937), .ZN(n9311) );
  NOR2_X2 U5045 ( .A1(n9332), .A2(n9331), .ZN(n9545) );
  AND2_X1 U5046 ( .A1(n9487), .A2(n9492), .ZN(n6098) );
  NAND2_X1 U5047 ( .A1(n6097), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6076) );
  OAI22_X2 U5048 ( .A1(n7817), .A2(n4857), .B1(n4859), .B2(n7905), .ZN(n8752)
         );
  OAI21_X2 U5049 ( .B1(n4667), .B2(n4666), .A(n4664), .ZN(n5170) );
  AOI21_X2 U5050 ( .B1(n7908), .B2(n7907), .A(n8688), .ZN(n8698) );
  NOR2_X2 U5051 ( .A1(n8689), .A2(n8690), .ZN(n8688) );
  AND2_X1 U5052 ( .A1(n5029), .A2(n7842), .ZN(n4405) );
  AND2_X1 U5053 ( .A1(n5029), .A2(n7842), .ZN(n4406) );
  AND2_X4 U5054 ( .A1(n5030), .A2(n7842), .ZN(n5120) );
  XNOR2_X2 U5055 ( .A(n5022), .B(n7846), .ZN(n5030) );
  AND2_X1 U5056 ( .A1(n5031), .A2(n5029), .ZN(n4407) );
  AND2_X2 U5057 ( .A1(n5031), .A2(n5029), .ZN(n4408) );
  AND2_X1 U5058 ( .A1(n5031), .A2(n5029), .ZN(n5121) );
  OAI21_X1 U5059 ( .B1(n5228), .B2(n4571), .A(n4569), .ZN(n4568) );
  NOR2_X1 U5060 ( .A1(n4680), .A2(n4570), .ZN(n4569) );
  INV_X1 U5061 ( .A(n5255), .ZN(n4570) );
  INV_X1 U5062 ( .A(n4681), .ZN(n4680) );
  OR2_X1 U5063 ( .A1(n8267), .A2(n8155), .ZN(n5858) );
  NAND2_X1 U5064 ( .A1(n7800), .A2(n5858), .ZN(n8529) );
  INV_X1 U5065 ( .A(n6739), .ZN(n6524) );
  INV_X1 U5066 ( .A(n4925), .ZN(n4924) );
  NAND2_X1 U5067 ( .A1(n4557), .A2(n4558), .ZN(n5366) );
  NAND2_X1 U5068 ( .A1(n8858), .A2(n8857), .ZN(n8863) );
  AOI21_X1 U5069 ( .B1(n4612), .B2(n4611), .A(n4610), .ZN(n4609) );
  AND2_X1 U5070 ( .A1(n8894), .A2(n8949), .ZN(n4611) );
  INV_X1 U5071 ( .A(n8991), .ZN(n4610) );
  OAI21_X1 U5072 ( .B1(n8893), .B2(n8892), .A(n4613), .ZN(n4612) );
  INV_X1 U5073 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5404) );
  INV_X1 U5074 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U5075 ( .A1(n5326), .A2(n5325), .ZN(n5329) );
  INV_X1 U5076 ( .A(SI_13_), .ZN(n5325) );
  NOR2_X1 U5077 ( .A1(n5295), .A2(n4682), .ZN(n4681) );
  INV_X1 U5078 ( .A(n5281), .ZN(n4682) );
  INV_X1 U5079 ( .A(n5294), .ZN(n5295) );
  OAI21_X1 U5080 ( .B1(n5228), .B2(n4571), .A(n5255), .ZN(n4565) );
  INV_X1 U5081 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5215) );
  INV_X1 U5082 ( .A(n5293), .ZN(n4787) );
  NOR2_X1 U5083 ( .A1(n8589), .A2(n8584), .ZN(n4656) );
  OR2_X1 U5084 ( .A1(n8594), .A2(n8429), .ZN(n5894) );
  NAND2_X1 U5085 ( .A1(n8407), .A2(n8429), .ZN(n4975) );
  OR2_X1 U5086 ( .A1(n8605), .A2(n8428), .ZN(n5876) );
  NOR2_X1 U5087 ( .A1(n4985), .A2(n8275), .ZN(n4984) );
  INV_X1 U5088 ( .A(n4988), .ZN(n4985) );
  NAND2_X1 U5089 ( .A1(n8485), .A2(n4987), .ZN(n4986) );
  INV_X1 U5090 ( .A(n4990), .ZN(n4987) );
  OR2_X1 U5091 ( .A1(n7704), .A2(n7703), .ZN(n5842) );
  INV_X1 U5092 ( .A(n9871), .ZN(n5687) );
  NOR2_X1 U5093 ( .A1(n5330), .A2(n4803), .ZN(n5043) );
  NAND2_X1 U5094 ( .A1(n10198), .A2(n5009), .ZN(n4488) );
  INV_X1 U5095 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5010) );
  AOI21_X1 U5096 ( .B1(n6760), .B2(n6759), .A(n6758), .ZN(n6765) );
  OR2_X1 U5097 ( .A1(n8665), .A2(n7922), .ZN(n7921) );
  NAND3_X1 U5098 ( .A1(n6981), .A2(n6766), .A3(n6769), .ZN(n6982) );
  AND2_X1 U5099 ( .A1(n4825), .A2(n4827), .ZN(n4824) );
  OR2_X1 U5100 ( .A1(n9258), .A2(n4529), .ZN(n4524) );
  INV_X1 U5101 ( .A(n4530), .ZN(n4529) );
  AND2_X1 U5102 ( .A1(n4527), .A2(n8918), .ZN(n4526) );
  NAND2_X1 U5103 ( .A1(n4530), .A2(n4528), .ZN(n4527) );
  INV_X1 U5104 ( .A(n8962), .ZN(n4528) );
  INV_X1 U5105 ( .A(n6409), .ZN(n6397) );
  NAND2_X1 U5106 ( .A1(n5748), .A2(n5747), .ZN(n5759) );
  NAND2_X1 U5107 ( .A1(n4896), .A2(n4900), .ZN(n5748) );
  AND2_X1 U5108 ( .A1(n5004), .A2(n4957), .ZN(n4956) );
  NOR2_X1 U5109 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n4957) );
  AND2_X1 U5110 ( .A1(n5517), .A2(n5501), .ZN(n5515) );
  NAND2_X1 U5111 ( .A1(n4582), .A2(n5452), .ZN(n5469) );
  NAND2_X1 U5112 ( .A1(n4562), .A2(n5365), .ZN(n5402) );
  OR2_X1 U5113 ( .A1(n5324), .A2(n4561), .ZN(n4557) );
  INV_X1 U5114 ( .A(n5347), .ZN(n4561) );
  OAI21_X1 U5115 ( .B1(n5227), .B2(n4563), .A(n4567), .ZN(n4677) );
  INV_X1 U5116 ( .A(n4568), .ZN(n4567) );
  XNOR2_X1 U5117 ( .A(n5297), .B(SI_11_), .ZN(n5294) );
  INV_X1 U5118 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6013) );
  NAND2_X1 U5119 ( .A1(n4669), .A2(n4670), .ZN(n5692) );
  AOI21_X1 U5120 ( .B1(n4672), .B2(n4797), .A(n4671), .ZN(n4670) );
  INV_X1 U5121 ( .A(n5629), .ZN(n4671) );
  NAND3_X1 U5122 ( .A1(n6673), .A2(n9871), .A3(n7307), .ZN(n5051) );
  INV_X1 U5123 ( .A(n5121), .ZN(n5645) );
  NOR2_X1 U5124 ( .A1(n8293), .A2(n8292), .ZN(n4648) );
  AOI21_X1 U5125 ( .B1(n4972), .B2(n4970), .A(n4969), .ZN(n4968) );
  INV_X1 U5126 ( .A(n4973), .ZN(n4970) );
  INV_X1 U5127 ( .A(n4972), .ZN(n4971) );
  AOI21_X1 U5128 ( .B1(n8277), .B2(n8457), .A(n8276), .ZN(n8441) );
  AND4_X1 U5129 ( .A1(n5168), .A2(n5167), .A3(n5166), .A4(n5165), .ZN(n7276)
         );
  NOR2_X1 U5130 ( .A1(n7276), .A2(n9882), .ZN(n4981) );
  NAND2_X1 U5131 ( .A1(n5038), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5046) );
  INV_X1 U5132 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4910) );
  INV_X1 U5133 ( .A(n7935), .ZN(n7988) );
  AND2_X1 U5134 ( .A1(n9487), .A2(n5991), .ZN(n6100) );
  AND2_X1 U5135 ( .A1(n9220), .A2(n9228), .ZN(n6295) );
  NAND2_X1 U5136 ( .A1(n7770), .A2(n4414), .ZN(n9330) );
  INV_X1 U5137 ( .A(n4949), .ZN(n4948) );
  AOI21_X1 U5138 ( .B1(n4949), .B2(n4947), .A(n4952), .ZN(n4946) );
  AND2_X1 U5139 ( .A1(n7618), .A2(n9041), .ZN(n4952) );
  AND2_X1 U5140 ( .A1(n6372), .A2(n6394), .ZN(n9791) );
  NOR2_X1 U5141 ( .A1(n4640), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4639) );
  INV_X1 U5142 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4628) );
  NAND2_X1 U5143 ( .A1(n5338), .A2(n5337), .ZN(n8267) );
  INV_X1 U5144 ( .A(n8861), .ZN(n4597) );
  NAND2_X1 U5145 ( .A1(n4592), .A2(n4591), .ZN(n8874) );
  NAND2_X1 U5146 ( .A1(n8866), .A2(n8944), .ZN(n4591) );
  NAND2_X1 U5147 ( .A1(n4593), .A2(n8949), .ZN(n4592) );
  NAND2_X1 U5148 ( .A1(n5847), .A2(n4536), .ZN(n5849) );
  AOI21_X1 U5149 ( .B1(n5846), .B2(n5922), .A(n4537), .ZN(n4536) );
  AND2_X1 U5150 ( .A1(n5845), .A2(n5911), .ZN(n4537) );
  NAND2_X1 U5151 ( .A1(n5868), .A2(n4551), .ZN(n4548) );
  OAI21_X1 U5152 ( .B1(n4607), .B2(n4606), .A(n4417), .ZN(n8919) );
  INV_X1 U5153 ( .A(n8918), .ZN(n4606) );
  AOI21_X1 U5154 ( .B1(n8916), .B2(n8962), .A(n4608), .ZN(n4607) );
  INV_X1 U5155 ( .A(n5739), .ZN(n4902) );
  NOR2_X1 U5156 ( .A1(n8031), .A2(n4668), .ZN(n5379) );
  INV_X1 U5157 ( .A(n8028), .ZN(n4668) );
  NAND2_X1 U5158 ( .A1(n4542), .A2(n5909), .ZN(n4541) );
  NAND2_X1 U5159 ( .A1(n4546), .A2(n4543), .ZN(n4542) );
  AND2_X1 U5160 ( .A1(n5905), .A2(n4544), .ZN(n4543) );
  OR2_X1 U5161 ( .A1(n8325), .A2(n4433), .ZN(n4539) );
  AND2_X1 U5162 ( .A1(n7351), .A2(n5829), .ZN(n4743) );
  AND2_X1 U5163 ( .A1(n8672), .A2(n4853), .ZN(n4852) );
  INV_X1 U5164 ( .A(n7899), .ZN(n4861) );
  NOR2_X1 U5165 ( .A1(n9220), .A2(n4695), .ZN(n4694) );
  AND2_X1 U5166 ( .A1(n4697), .A2(n9305), .ZN(n4699) );
  INV_X1 U5167 ( .A(n4701), .ZN(n4697) );
  NAND2_X1 U5168 ( .A1(n8845), .A2(n6896), .ZN(n8973) );
  INV_X1 U5169 ( .A(n4901), .ZN(n4900) );
  OAI21_X1 U5170 ( .B1(n5737), .B2(n4902), .A(n5743), .ZN(n4901) );
  INV_X1 U5171 ( .A(n5195), .ZN(n4881) );
  INV_X1 U5172 ( .A(n5173), .ZN(n4880) );
  OR2_X1 U5173 ( .A1(n7629), .A2(n4787), .ZN(n4786) );
  INV_X1 U5174 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5331) );
  OR2_X1 U5175 ( .A1(n8318), .A2(n8564), .ZN(n8293) );
  OR2_X1 U5176 ( .A1(n8564), .A2(n8286), .ZN(n5913) );
  OR2_X1 U5177 ( .A1(n8576), .A2(n8357), .ZN(n5905) );
  INV_X1 U5178 ( .A(n5732), .ZN(n4757) );
  AND2_X1 U5179 ( .A1(n4735), .A2(n4734), .ZN(n4733) );
  INV_X1 U5180 ( .A(n5863), .ZN(n4739) );
  OR2_X1 U5181 ( .A1(n8538), .A2(n8503), .ZN(n5863) );
  AND2_X1 U5182 ( .A1(n5854), .A2(n5853), .ZN(n7751) );
  NAND2_X1 U5183 ( .A1(n7704), .A2(n7703), .ZN(n5844) );
  NOR2_X1 U5184 ( .A1(n5163), .A2(n5162), .ZN(n5187) );
  NAND2_X1 U5185 ( .A1(n8176), .A2(n6949), .ZN(n5805) );
  INV_X1 U5186 ( .A(n7307), .ZN(n5804) );
  NAND2_X1 U5187 ( .A1(n8024), .A2(n7890), .ZN(n6667) );
  NAND2_X1 U5188 ( .A1(n8458), .A2(n5729), .ZN(n4724) );
  OR2_X1 U5189 ( .A1(n5675), .A2(n7702), .ZN(n5680) );
  AND2_X1 U5190 ( .A1(n7682), .A2(n5671), .ZN(n5675) );
  INV_X1 U5191 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5020) );
  INV_X1 U5192 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4763) );
  NAND2_X1 U5193 ( .A1(n5668), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U5194 ( .A1(n5082), .A2(n4641), .ZN(n5103) );
  NAND2_X1 U5196 ( .A1(n4852), .A2(n4849), .ZN(n4848) );
  NOR2_X1 U5197 ( .A1(n4850), .A2(n4842), .ZN(n4841) );
  INV_X1 U5198 ( .A(n7923), .ZN(n4842) );
  INV_X1 U5199 ( .A(n4852), .ZN(n4850) );
  INV_X1 U5200 ( .A(n4480), .ZN(n4851) );
  NOR2_X1 U5201 ( .A1(n4851), .A2(n4849), .ZN(n4845) );
  OR2_X1 U5202 ( .A1(n4851), .A2(n4852), .ZN(n4844) );
  AND2_X1 U5203 ( .A1(n7818), .A2(n4861), .ZN(n4860) );
  OR2_X1 U5204 ( .A1(n7818), .A2(n4861), .ZN(n4859) );
  NAND2_X1 U5205 ( .A1(n9363), .A2(n8942), .ZN(n4603) );
  OR2_X1 U5206 ( .A1(n6320), .A2(n9977), .ZN(n6330) );
  OR2_X1 U5207 ( .A1(n9249), .A2(n7932), .ZN(n9224) );
  AND2_X1 U5208 ( .A1(n8888), .A2(n4505), .ZN(n4504) );
  NAND2_X1 U5209 ( .A1(n8872), .A2(n8789), .ZN(n4505) );
  INV_X1 U5210 ( .A(n4818), .ZN(n4817) );
  INV_X1 U5211 ( .A(n6126), .ZN(n4945) );
  AND2_X1 U5212 ( .A1(n8857), .A2(n8977), .ZN(n4818) );
  OR2_X1 U5213 ( .A1(n9467), .A2(n9389), .ZN(n8961) );
  INV_X1 U5214 ( .A(n8772), .ZN(n4807) );
  INV_X1 U5215 ( .A(n6434), .ZN(n4806) );
  OAI21_X1 U5216 ( .B1(n5609), .B2(n5608), .A(n5607), .ZN(n5631) );
  AND2_X1 U5217 ( .A1(n5579), .A2(n5566), .ZN(n5578) );
  INV_X1 U5218 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6351) );
  NAND2_X1 U5219 ( .A1(n5538), .A2(n5537), .ZN(n5559) );
  NAND2_X1 U5220 ( .A1(n5518), .A2(n5517), .ZN(n5532) );
  NAND2_X1 U5221 ( .A1(n4575), .A2(n4573), .ZN(n5518) );
  AOI21_X1 U5222 ( .B1(n4576), .B2(n4579), .A(n4574), .ZN(n4573) );
  NAND2_X1 U5223 ( .A1(n5406), .A2(n5405), .ZN(n5431) );
  AOI21_X1 U5224 ( .B1(n5347), .B2(n4560), .A(n4559), .ZN(n4558) );
  INV_X1 U5225 ( .A(n5329), .ZN(n4559) );
  INV_X1 U5226 ( .A(n5321), .ZN(n4676) );
  NAND2_X1 U5227 ( .A1(n5258), .A2(n5257), .ZN(n5281) );
  INV_X1 U5228 ( .A(SI_10_), .ZN(n5257) );
  OAI21_X1 U5229 ( .B1(n5227), .B2(n4566), .A(n4564), .ZN(n5280) );
  NAND2_X1 U5230 ( .A1(n4404), .A2(n5002), .ZN(n4566) );
  INV_X1 U5231 ( .A(n4565), .ZN(n4564) );
  NAND2_X1 U5232 ( .A1(n5217), .A2(n5216), .ZN(n5228) );
  NAND2_X1 U5233 ( .A1(n6077), .A2(n4501), .ZN(n6106) );
  INV_X1 U5234 ( .A(n9885), .ZN(n7356) );
  NAND2_X1 U5235 ( .A1(n5547), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5569) );
  INV_X1 U5236 ( .A(n5641), .ZN(n8055) );
  NOR2_X1 U5237 ( .A1(n7109), .A2(n4781), .ZN(n4780) );
  INV_X1 U5238 ( .A(n5186), .ZN(n4781) );
  INV_X1 U5239 ( .A(n7290), .ZN(n4645) );
  INV_X1 U5240 ( .A(n4775), .ZN(n4774) );
  OAI21_X1 U5241 ( .B1(n4780), .B2(n4776), .A(n7169), .ZN(n4775) );
  INV_X1 U5242 ( .A(n4777), .ZN(n4776) );
  OAI21_X1 U5243 ( .B1(n7630), .B2(n4787), .A(n4426), .ZN(n7737) );
  INV_X1 U5244 ( .A(n5353), .ZN(n5339) );
  OR2_X1 U5245 ( .A1(n8083), .A2(n4796), .ZN(n4795) );
  INV_X1 U5246 ( .A(n8082), .ZN(n4796) );
  NAND2_X1 U5247 ( .A1(n4675), .A2(n5378), .ZN(n5387) );
  INV_X1 U5248 ( .A(n5396), .ZN(n4675) );
  NAND2_X1 U5249 ( .A1(n5050), .A2(n5689), .ZN(n6673) );
  NAND2_X1 U5250 ( .A1(n8178), .A2(n4717), .ZN(n8190) );
  OR2_X1 U5251 ( .A1(n6735), .A2(n7892), .ZN(n4717) );
  OR2_X1 U5252 ( .A1(n6800), .A2(n6799), .ZN(n4719) );
  INV_X1 U5253 ( .A(n4648), .ZN(n8294) );
  NAND2_X1 U5254 ( .A1(n5751), .A2(n5750), .ZN(n8292) );
  NAND2_X1 U5255 ( .A1(n5794), .A2(n5790), .ZN(n8282) );
  NAND2_X1 U5256 ( .A1(n8311), .A2(n8530), .ZN(n4768) );
  NAND2_X1 U5257 ( .A1(n5913), .A2(n5914), .ZN(n8308) );
  XNOR2_X1 U5258 ( .A(n8569), .B(n8062), .ZN(n8325) );
  AND2_X1 U5259 ( .A1(n8373), .A2(n5896), .ZN(n4759) );
  NAND2_X1 U5260 ( .A1(n8390), .A2(n5732), .ZN(n8393) );
  AND2_X1 U5261 ( .A1(n4975), .A2(n8278), .ZN(n4973) );
  NAND2_X1 U5262 ( .A1(n4452), .A2(n4975), .ZN(n4972) );
  OR2_X1 U5263 ( .A1(n8447), .A2(n8428), .ZN(n4995) );
  OR2_X1 U5264 ( .A1(n8452), .A2(n8605), .ZN(n8443) );
  NAND2_X1 U5265 ( .A1(n4983), .A2(n4982), .ZN(n8451) );
  NOR2_X1 U5266 ( .A1(n8490), .A2(n8615), .ZN(n8468) );
  NAND2_X1 U5267 ( .A1(n4989), .A2(n8501), .ZN(n4988) );
  NAND2_X1 U5268 ( .A1(n5438), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5481) );
  AOI21_X1 U5269 ( .B1(n4738), .B2(n8526), .A(n4736), .ZN(n4735) );
  INV_X1 U5270 ( .A(n5864), .ZN(n4736) );
  AND2_X1 U5271 ( .A1(n8626), .A2(n8532), .ZN(n4990) );
  OR2_X1 U5272 ( .A1(n8507), .A2(n4986), .ZN(n8482) );
  NOR2_X1 U5273 ( .A1(n8267), .A2(n8538), .ZN(n4651) );
  NAND2_X1 U5274 ( .A1(n7805), .A2(n4415), .ZN(n8514) );
  NAND2_X1 U5275 ( .A1(n4747), .A2(n4419), .ZN(n7800) );
  NOR2_X1 U5276 ( .A1(n9920), .A2(n4661), .ZN(n4659) );
  NOR2_X1 U5277 ( .A1(n7762), .A2(n9525), .ZN(n7805) );
  NOR2_X1 U5278 ( .A1(n5725), .A2(n4765), .ZN(n4764) );
  INV_X1 U5279 ( .A(n5835), .ZN(n4765) );
  AND2_X1 U5280 ( .A1(n5842), .A2(n5844), .ZN(n7562) );
  NAND2_X1 U5281 ( .A1(n7497), .A2(n7495), .ZN(n7559) );
  AND4_X1 U5282 ( .A1(n5208), .A2(n5207), .A3(n5206), .A4(n5205), .ZN(n7506)
         );
  AOI21_X1 U5283 ( .B1(n4449), .B2(n7276), .A(n4980), .ZN(n4979) );
  NOR2_X1 U5284 ( .A1(n7259), .A2(n7349), .ZN(n4980) );
  INV_X1 U5285 ( .A(n8502), .ZN(n8530) );
  AND2_X1 U5286 ( .A1(n6727), .A2(n8646), .ZN(n8533) );
  NAND2_X1 U5287 ( .A1(n7338), .A2(n7351), .ZN(n7337) );
  AND2_X1 U5288 ( .A1(n5825), .A2(n5820), .ZN(n7351) );
  NAND2_X1 U5289 ( .A1(n7325), .A2(n6952), .ZN(n4960) );
  NOR2_X1 U5290 ( .A1(n4964), .A2(n4963), .ZN(n4962) );
  AND4_X1 U5291 ( .A1(n5144), .A2(n5143), .A3(n5142), .A4(n5141), .ZN(n7258)
         );
  NAND2_X1 U5292 ( .A1(n7334), .A2(n7333), .ZN(n7332) );
  OR2_X1 U5293 ( .A1(n6526), .A2(n8646), .ZN(n8502) );
  NAND2_X1 U5294 ( .A1(n5805), .A2(n5807), .ZN(n6910) );
  OR2_X1 U5295 ( .A1(n9524), .A2(n5804), .ZN(n7264) );
  INV_X1 U5296 ( .A(n8563), .ZN(n4746) );
  AND2_X1 U5297 ( .A1(n5240), .A2(n5239), .ZN(n9899) );
  OR2_X1 U5298 ( .A1(n9871), .A2(n7451), .ZN(n5688) );
  NAND2_X1 U5299 ( .A1(n6425), .A2(n9868), .ZN(n9862) );
  INV_X1 U5300 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5025) );
  XNOR2_X1 U5301 ( .A(n5053), .B(n5021), .ZN(n5705) );
  NAND2_X1 U5302 ( .A1(n5055), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5053) );
  NAND2_X1 U5303 ( .A1(n5684), .A2(n5683), .ZN(n5686) );
  INV_X1 U5304 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5042) );
  NAND2_X1 U5305 ( .A1(n5046), .A2(n10255), .ZN(n5049) );
  NAND2_X1 U5306 ( .A1(n4801), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5455) );
  NOR2_X1 U5307 ( .A1(n4422), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n4802) );
  INV_X1 U5308 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5008) );
  INV_X1 U5309 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5411) );
  XNOR2_X1 U5310 ( .A(n6972), .B(n6564), .ZN(n6614) );
  AOI21_X1 U5311 ( .B1(n4634), .B2(n4632), .A(n4477), .ZN(n4631) );
  INV_X1 U5312 ( .A(n8680), .ZN(n4632) );
  INV_X1 U5313 ( .A(n4634), .ZN(n4633) );
  AOI21_X1 U5314 ( .B1(n4833), .B2(n4836), .A(n4830), .ZN(n4829) );
  XNOR2_X1 U5315 ( .A(n6617), .B(n6972), .ZN(n6751) );
  NOR2_X1 U5316 ( .A1(n4836), .A2(n4625), .ZN(n4624) );
  NOR2_X1 U5317 ( .A1(n7653), .A2(n4874), .ZN(n4873) );
  INV_X1 U5318 ( .A(n7641), .ZN(n4874) );
  XNOR2_X1 U5319 ( .A(n6588), .B(n6972), .ZN(n6592) );
  AOI22_X1 U5320 ( .A1(n6590), .A2(n6589), .B1(n7811), .B2(n7862), .ZN(n6591)
         );
  INV_X1 U5321 ( .A(n6627), .ZN(n6580) );
  INV_X1 U5322 ( .A(n6629), .ZN(n6582) );
  CLKBUF_X1 U5323 ( .A(n6982), .Z(n6767) );
  AND2_X1 U5324 ( .A1(n8746), .A2(n4469), .ZN(n4634) );
  NOR2_X1 U5325 ( .A1(n9024), .A2(n6348), .ZN(n4884) );
  NAND2_X1 U5326 ( .A1(n7061), .A2(n9679), .ZN(n7200) );
  INV_X1 U5327 ( .A(n4510), .ZN(n4509) );
  OAI21_X1 U5328 ( .B1(n6338), .B2(n4513), .A(n4511), .ZN(n4510) );
  NAND2_X1 U5329 ( .A1(n9135), .A2(n4512), .ZN(n4511) );
  NAND2_X1 U5330 ( .A1(n9134), .A2(n9132), .ZN(n4513) );
  NAND2_X1 U5331 ( .A1(n4821), .A2(n9010), .ZN(n4820) );
  INV_X1 U5332 ( .A(n4824), .ZN(n4821) );
  OR2_X1 U5333 ( .A1(n9178), .A2(n8825), .ZN(n4826) );
  INV_X1 U5334 ( .A(n4828), .ZN(n4827) );
  OAI21_X1 U5335 ( .B1(n8825), .B2(n8932), .A(n8837), .ZN(n4828) );
  NAND2_X1 U5336 ( .A1(n4423), .A2(n4409), .ZN(n4927) );
  OR2_X1 U5337 ( .A1(n4434), .A2(n8838), .ZN(n9156) );
  NAND2_X1 U5338 ( .A1(n4409), .A2(n6297), .ZN(n4928) );
  OR2_X1 U5339 ( .A1(n9185), .A2(n9197), .ZN(n9175) );
  AND2_X1 U5340 ( .A1(n8957), .A2(n8956), .ZN(n9194) );
  AOI21_X1 U5341 ( .B1(n8959), .B2(n4815), .A(n4814), .ZN(n4813) );
  INV_X1 U5342 ( .A(n8961), .ZN(n4815) );
  INV_X1 U5343 ( .A(n8958), .ZN(n4814) );
  NAND2_X1 U5344 ( .A1(n4524), .A2(n4441), .ZN(n4812) );
  NAND2_X1 U5345 ( .A1(n4932), .A2(n4931), .ZN(n9207) );
  AOI21_X1 U5346 ( .B1(n4933), .B2(n4935), .A(n4476), .ZN(n4931) );
  OR2_X1 U5347 ( .A1(n7932), .A2(n9471), .ZN(n4996) );
  NAND2_X1 U5348 ( .A1(n9240), .A2(n9239), .ZN(n9238) );
  NAND2_X1 U5349 ( .A1(n9273), .A2(n8914), .ZN(n9258) );
  NAND2_X1 U5350 ( .A1(n6228), .A2(n6227), .ZN(n9332) );
  OR2_X1 U5351 ( .A1(n9484), .A2(n9339), .ZN(n4994) );
  NAND2_X1 U5352 ( .A1(n4519), .A2(n4521), .ZN(n7770) );
  NAND2_X1 U5353 ( .A1(n4520), .A2(n8894), .ZN(n4519) );
  INV_X1 U5354 ( .A(n7686), .ZN(n4520) );
  AND2_X1 U5355 ( .A1(n8803), .A2(n8896), .ZN(n8991) );
  NAND2_X1 U5356 ( .A1(n7686), .A2(n6366), .ZN(n7688) );
  AND2_X1 U5357 ( .A1(n8804), .A2(n8890), .ZN(n8990) );
  NOR2_X1 U5358 ( .A1(n8965), .A2(n4950), .ZN(n4949) );
  NAND2_X1 U5359 ( .A1(n7476), .A2(n8986), .ZN(n7475) );
  AOI21_X1 U5360 ( .B1(n4940), .B2(n4942), .A(n4432), .ZN(n4939) );
  NAND2_X1 U5361 ( .A1(n8864), .A2(n8875), .ZN(n6150) );
  NAND2_X1 U5362 ( .A1(n6151), .A2(n6150), .ZN(n7088) );
  NAND2_X1 U5363 ( .A1(n6944), .A2(n4818), .ZN(n6894) );
  NAND2_X1 U5364 ( .A1(n6364), .A2(n4410), .ZN(n6944) );
  NAND2_X1 U5365 ( .A1(n4920), .A2(n6085), .ZN(n4919) );
  NAND2_X1 U5366 ( .A1(n8775), .A2(n8774), .ZN(n9110) );
  NAND2_X1 U5367 ( .A1(n6180), .A2(n6179), .ZN(n9553) );
  INV_X1 U5368 ( .A(n9791), .ZN(n9733) );
  INV_X1 U5369 ( .A(n9361), .ZN(n9794) );
  NAND2_X1 U5370 ( .A1(n6398), .A2(n6397), .ZN(n9718) );
  NOR2_X1 U5371 ( .A1(n4895), .A2(n5777), .ZN(n4893) );
  INV_X1 U5372 ( .A(n5777), .ZN(n4892) );
  XNOR2_X1 U5373 ( .A(n5778), .B(n5761), .ZN(n8776) );
  XNOR2_X1 U5374 ( .A(n5744), .B(n5743), .ZN(n7885) );
  NAND2_X1 U5375 ( .A1(n4899), .A2(n5739), .ZN(n5744) );
  NAND2_X1 U5376 ( .A1(n5738), .A2(n5737), .ZN(n4899) );
  NOR2_X1 U5377 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6385) );
  AND2_X1 U5378 ( .A1(n4639), .A2(n4637), .ZN(n4636) );
  INV_X1 U5379 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4637) );
  NAND2_X1 U5380 ( .A1(n6351), .A2(n6391), .ZN(n4640) );
  XNOR2_X1 U5381 ( .A(n4556), .B(n5578), .ZN(n7539) );
  OAI21_X1 U5382 ( .B1(n5559), .B2(n5558), .A(n5560), .ZN(n4556) );
  NAND2_X1 U5383 ( .A1(n6345), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6347) );
  NAND2_X1 U5384 ( .A1(n4572), .A2(n4576), .ZN(n5516) );
  OR2_X1 U5385 ( .A1(n5432), .A2(n4579), .ZN(n4572) );
  OAI21_X1 U5386 ( .B1(n6241), .B2(P1_IR_REG_18__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6242) );
  NAND2_X1 U5387 ( .A1(n4918), .A2(n5471), .ZN(n5496) );
  NAND2_X1 U5388 ( .A1(n5469), .A2(n5468), .ZN(n4918) );
  NAND2_X1 U5389 ( .A1(n4677), .A2(n4678), .ZN(n5322) );
  AND2_X1 U5390 ( .A1(n6009), .A2(n6051), .ZN(n6119) );
  AOI21_X1 U5391 ( .B1(n5150), .B2(n4665), .A(n4447), .ZN(n4664) );
  INV_X1 U5392 ( .A(n8169), .ZN(n9830) );
  NAND2_X1 U5393 ( .A1(n4792), .A2(n4791), .ZN(n4790) );
  INV_X1 U5394 ( .A(n5095), .ZN(n4791) );
  AND2_X1 U5395 ( .A1(n8068), .A2(n8138), .ZN(n8058) );
  NAND2_X1 U5396 ( .A1(n4779), .A2(n4778), .ZN(n4777) );
  INV_X1 U5397 ( .A(n5202), .ZN(n4779) );
  INV_X1 U5398 ( .A(n5201), .ZN(n4778) );
  NAND2_X1 U5399 ( .A1(n7100), .A2(n4780), .ZN(n4773) );
  INV_X1 U5400 ( .A(n8423), .ZN(n8601) );
  NAND2_X1 U5401 ( .A1(n5581), .A2(n5580), .ZN(n8584) );
  AND3_X1 U5402 ( .A1(n5573), .A2(n5572), .A3(n5571), .ZN(n8414) );
  AND4_X1 U5403 ( .A1(n5526), .A2(n5525), .A3(n5524), .A4(n5523), .ZN(n8413)
         );
  INV_X1 U5404 ( .A(n6920), .ZN(n5160) );
  AND3_X1 U5405 ( .A1(n5180), .A2(n5179), .A3(n5178), .ZN(n9882) );
  AND4_X1 U5406 ( .A1(n5193), .A2(n5192), .A3(n5191), .A4(n5190), .ZN(n7357)
         );
  INV_X1 U5407 ( .A(n8138), .ZN(n9826) );
  AND2_X1 U5408 ( .A1(n6796), .A2(n4720), .ZN(n6800) );
  NAND2_X1 U5409 ( .A1(n6797), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4720) );
  AND2_X1 U5410 ( .A1(n5336), .A2(n5372), .ZN(n8224) );
  OAI21_X1 U5411 ( .B1(n8255), .B2(n8254), .A(n4716), .ZN(n4715) );
  AOI21_X1 U5412 ( .B1(n8257), .B2(n8258), .A(n8256), .ZN(n4716) );
  OAI21_X1 U5413 ( .B1(n8262), .B2(n4911), .A(n8261), .ZN(n4714) );
  INV_X1 U5414 ( .A(n8254), .ZN(n8253) );
  INV_X1 U5415 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n7846) );
  INV_X1 U5416 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10015) );
  NOR2_X1 U5417 ( .A1(n4866), .A2(n7995), .ZN(n4864) );
  NOR2_X1 U5418 ( .A1(n4437), .A2(n4867), .ZN(n4866) );
  INV_X1 U5419 ( .A(n4869), .ZN(n4867) );
  NAND2_X1 U5420 ( .A1(n4869), .A2(n4870), .ZN(n4868) );
  INV_X1 U5421 ( .A(n7965), .ZN(n4870) );
  NAND2_X1 U5422 ( .A1(n6208), .A2(n6207), .ZN(n7824) );
  NAND2_X1 U5423 ( .A1(n8735), .A2(n5007), .ZN(n4620) );
  NOR2_X1 U5424 ( .A1(n4416), .A2(n4438), .ZN(n4532) );
  NOR2_X1 U5425 ( .A1(n6479), .A2(n6512), .ZN(n6482) );
  XOR2_X1 U5426 ( .A(n7202), .B(n7200), .Z(n7062) );
  AND2_X1 U5427 ( .A1(n6416), .A2(n6415), .ZN(n9486) );
  NAND2_X1 U5428 ( .A1(n6001), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6002) );
  INV_X1 U5429 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4912) );
  OAI21_X1 U5430 ( .B1(n8863), .B2(n8862), .A(n4595), .ZN(n4594) );
  NOR2_X1 U5431 ( .A1(n4597), .A2(n4596), .ZN(n4595) );
  NAND2_X1 U5432 ( .A1(n4553), .A2(n4552), .ZN(n5837) );
  NAND2_X1 U5433 ( .A1(n5836), .A2(n5911), .ZN(n4553) );
  NAND2_X1 U5434 ( .A1(n4587), .A2(n4947), .ZN(n8889) );
  NOR2_X1 U5435 ( .A1(n4614), .A2(n6365), .ZN(n4613) );
  INV_X1 U5436 ( .A(n8891), .ZN(n4614) );
  NAND2_X1 U5437 ( .A1(n5849), .A2(n5943), .ZN(n5850) );
  AND2_X1 U5438 ( .A1(n8528), .A2(n5859), .ZN(n4549) );
  INV_X1 U5439 ( .A(n5872), .ZN(n4551) );
  OAI21_X1 U5440 ( .B1(n8895), .B2(n8949), .A(n4609), .ZN(n8901) );
  INV_X1 U5441 ( .A(n8917), .ZN(n4608) );
  AND2_X1 U5442 ( .A1(n5885), .A2(n5881), .ZN(n4550) );
  NAND2_X1 U5443 ( .A1(n4545), .A2(n5911), .ZN(n4544) );
  INV_X1 U5444 ( .A(n5906), .ZN(n4545) );
  INV_X1 U5445 ( .A(n8788), .ZN(n4811) );
  NAND2_X1 U5446 ( .A1(n9327), .A2(n4698), .ZN(n4701) );
  NOR2_X1 U5447 ( .A1(n4898), .A2(n4902), .ZN(n4897) );
  INV_X1 U5448 ( .A(n5632), .ZN(n4898) );
  NAND2_X1 U5449 ( .A1(n5631), .A2(n5630), .ZN(n5633) );
  AND2_X1 U5450 ( .A1(n4908), .A2(n5578), .ZN(n4907) );
  NAND2_X1 U5451 ( .A1(n5558), .A2(n5560), .ZN(n4908) );
  INV_X1 U5452 ( .A(n5560), .ZN(n4905) );
  INV_X1 U5453 ( .A(n5515), .ZN(n4574) );
  INV_X1 U5454 ( .A(n5497), .ZN(n4914) );
  NOR2_X1 U5455 ( .A1(n5495), .A2(n4917), .ZN(n4916) );
  INV_X1 U5456 ( .A(n5471), .ZN(n4917) );
  NOR2_X1 U5457 ( .A1(n4915), .A2(n4581), .ZN(n4580) );
  INV_X1 U5458 ( .A(n5452), .ZN(n4581) );
  INV_X1 U5459 ( .A(n4916), .ZN(n4915) );
  NOR2_X1 U5460 ( .A1(n5453), .A2(n4584), .ZN(n4583) );
  INV_X1 U5461 ( .A(n5431), .ZN(n4584) );
  INV_X1 U5462 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5434) );
  INV_X1 U5463 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5433) );
  INV_X1 U5464 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n5367) );
  INV_X1 U5465 ( .A(SI_14_), .ZN(n10080) );
  INV_X1 U5466 ( .A(SI_9_), .ZN(n5229) );
  NOR2_X1 U5467 ( .A1(n4785), .A2(n4443), .ZN(n4784) );
  INV_X1 U5468 ( .A(n5395), .ZN(n4785) );
  AOI21_X1 U5469 ( .B1(n4541), .B2(n4540), .A(n4539), .ZN(n5917) );
  OR2_X1 U5470 ( .A1(n8581), .A2(n8140), .ZN(n5906) );
  OR2_X1 U5471 ( .A1(n5521), .A2(n8076), .ZN(n5549) );
  OR2_X1 U5472 ( .A1(n8601), .A2(n8413), .ZN(n5889) );
  NAND2_X1 U5473 ( .A1(n4662), .A2(n9916), .ZN(n4661) );
  NOR2_X1 U5474 ( .A1(n7704), .A2(n7517), .ZN(n4662) );
  NAND2_X1 U5475 ( .A1(n7517), .A2(n9830), .ZN(n5835) );
  NAND2_X1 U5476 ( .A1(n4741), .A2(n5829), .ZN(n4740) );
  NAND2_X1 U5477 ( .A1(n5825), .A2(n4978), .ZN(n4741) );
  INV_X1 U5478 ( .A(n6952), .ZN(n4964) );
  INV_X1 U5479 ( .A(n6950), .ZN(n4963) );
  NOR2_X1 U5480 ( .A1(n7513), .A2(n7517), .ZN(n7568) );
  OR2_X1 U5481 ( .A1(n7367), .A2(n7494), .ZN(n7513) );
  NOR2_X1 U5482 ( .A1(n7340), .A2(n7349), .ZN(n7341) );
  NAND2_X1 U5483 ( .A1(n4644), .A2(n7449), .ZN(n7340) );
  INV_X1 U5484 ( .A(n7013), .ZN(n4644) );
  NAND2_X1 U5485 ( .A1(n4646), .A2(n4645), .ZN(n7013) );
  INV_X1 U5486 ( .A(n7327), .ZN(n4646) );
  NAND2_X1 U5487 ( .A1(n7328), .A2(n4727), .ZN(n7327) );
  INV_X1 U5488 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5021) );
  INV_X1 U5489 ( .A(n4762), .ZN(n4761) );
  INV_X1 U5490 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5683) );
  INV_X1 U5491 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5037) );
  INV_X1 U5492 ( .A(n5036), .ZN(n4804) );
  NAND2_X1 U5493 ( .A1(n5303), .A2(n5015), .ZN(n5330) );
  INV_X1 U5494 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5334) );
  INV_X1 U5495 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4642) );
  INV_X1 U5496 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4643) );
  INV_X1 U5497 ( .A(n7133), .ZN(n4835) );
  INV_X1 U5498 ( .A(n7180), .ZN(n4834) );
  INV_X1 U5499 ( .A(n6983), .ZN(n4625) );
  NAND2_X1 U5500 ( .A1(n9110), .A2(n9113), .ZN(n8946) );
  NAND2_X1 U5501 ( .A1(n4411), .A2(n9363), .ZN(n4704) );
  INV_X1 U5502 ( .A(n9132), .ZN(n4512) );
  NAND2_X1 U5503 ( .A1(n9010), .A2(n4823), .ZN(n4822) );
  NAND2_X1 U5504 ( .A1(n8939), .A2(n9132), .ZN(n8998) );
  OAI21_X1 U5505 ( .B1(n4927), .B2(n4434), .A(n4926), .ZN(n4925) );
  INV_X1 U5506 ( .A(n8838), .ZN(n4926) );
  INV_X1 U5507 ( .A(n4996), .ZN(n4935) );
  INV_X1 U5508 ( .A(n4934), .ZN(n4933) );
  OAI21_X1 U5509 ( .B1(n9239), .B2(n4935), .A(n6285), .ZN(n4934) );
  NAND2_X1 U5510 ( .A1(n9467), .A2(n9247), .ZN(n6285) );
  NAND2_X1 U5511 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(n6278), .ZN(n6289) );
  INV_X1 U5512 ( .A(n6288), .ZN(n6278) );
  AND2_X1 U5513 ( .A1(n9244), .A2(n4531), .ZN(n4530) );
  INV_X1 U5514 ( .A(n4810), .ZN(n4809) );
  OAI21_X1 U5515 ( .B1(n4414), .B2(n4811), .A(n8907), .ZN(n4810) );
  NAND2_X1 U5516 ( .A1(n4518), .A2(n4523), .ZN(n4517) );
  NAND2_X1 U5517 ( .A1(n7379), .A2(n4418), .ZN(n4690) );
  NOR2_X1 U5518 ( .A1(n9553), .A2(n7392), .ZN(n4689) );
  INV_X1 U5519 ( .A(n4941), .ZN(n4940) );
  OAI21_X1 U5520 ( .B1(n6150), .B2(n4942), .A(n6164), .ZN(n4941) );
  INV_X1 U5521 ( .A(n6152), .ZN(n4942) );
  NAND2_X1 U5522 ( .A1(n6248), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n4619) );
  NAND2_X1 U5523 ( .A1(n9248), .A2(n4691), .ZN(n9183) );
  NOR2_X1 U5524 ( .A1(n9185), .A2(n4693), .ZN(n4691) );
  NAND2_X1 U5525 ( .A1(n9248), .A2(n4694), .ZN(n9213) );
  NAND2_X1 U5526 ( .A1(n4700), .A2(n4420), .ZN(n9285) );
  NAND2_X1 U5527 ( .A1(n4700), .A2(n4699), .ZN(n9304) );
  NOR2_X1 U5528 ( .A1(n9340), .A2(n4701), .ZN(n9318) );
  NOR2_X1 U5529 ( .A1(n9340), .A2(n9539), .ZN(n9342) );
  NOR2_X1 U5530 ( .A1(n4690), .A2(n7645), .ZN(n7692) );
  NAND2_X1 U5531 ( .A1(n8976), .A2(n8974), .ZN(n6893) );
  AND2_X1 U5532 ( .A1(n5739), .A2(n5637), .ZN(n5737) );
  OAI21_X1 U5533 ( .B1(n5597), .B2(n5596), .A(n5595), .ZN(n5609) );
  OAI21_X1 U5534 ( .B1(n5559), .B2(n4906), .A(n4903), .ZN(n5597) );
  AOI21_X1 U5535 ( .B1(n4907), .B2(n4905), .A(n4904), .ZN(n4903) );
  INV_X1 U5536 ( .A(n4907), .ZN(n4906) );
  INV_X1 U5537 ( .A(n5579), .ZN(n4904) );
  AOI21_X1 U5538 ( .B1(n4580), .B2(n4578), .A(n4577), .ZN(n4576) );
  INV_X1 U5539 ( .A(n4583), .ZN(n4578) );
  INV_X1 U5540 ( .A(n4913), .ZN(n4577) );
  AOI21_X1 U5541 ( .B1(n5467), .B2(n4916), .A(n4914), .ZN(n4913) );
  INV_X1 U5542 ( .A(n4580), .ZN(n4579) );
  INV_X1 U5543 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6341) );
  INV_X1 U5544 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6342) );
  OAI21_X1 U5545 ( .B1(n5402), .B2(n5401), .A(n5400), .ZN(n5430) );
  AND2_X1 U5546 ( .A1(n5431), .A2(n5408), .ZN(n5429) );
  NAND2_X1 U5547 ( .A1(n5300), .A2(n5299), .ZN(n5323) );
  AND2_X1 U5548 ( .A1(n5329), .A2(n5328), .ZN(n5347) );
  AOI21_X1 U5549 ( .B1(n4681), .B2(n4679), .A(n4446), .ZN(n4678) );
  INV_X1 U5550 ( .A(n5001), .ZN(n4679) );
  NAND2_X1 U5551 ( .A1(n5219), .A2(n5228), .ZN(n5226) );
  AOI21_X1 U5552 ( .B1(n5195), .B2(n4880), .A(n4448), .ZN(n4879) );
  INV_X1 U5553 ( .A(n5133), .ZN(n4665) );
  XNOR2_X1 U5554 ( .A(n8267), .B(n8055), .ZN(n5384) );
  AND2_X1 U5555 ( .A1(n8067), .A2(n5655), .ZN(n5691) );
  INV_X1 U5556 ( .A(n5494), .ZN(n4794) );
  CLKBUF_X1 U5557 ( .A(n8047), .Z(n4494) );
  INV_X1 U5558 ( .A(n4795), .ZN(n4673) );
  AND2_X1 U5559 ( .A1(n5650), .A2(n5649), .ZN(n8062) );
  NAND2_X1 U5560 ( .A1(n8180), .A2(n8179), .ZN(n8178) );
  NOR2_X1 U5561 ( .A1(n7141), .A2(n4708), .ZN(n7144) );
  AND2_X1 U5562 ( .A1(n7147), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4708) );
  NAND2_X1 U5563 ( .A1(n7144), .A2(n7143), .ZN(n7602) );
  NAND2_X1 U5564 ( .A1(n7602), .A2(n4707), .ZN(n8216) );
  OR2_X1 U5565 ( .A1(n7611), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4707) );
  NAND2_X1 U5566 ( .A1(n8216), .A2(n8217), .ZN(n8215) );
  NOR2_X1 U5567 ( .A1(n8283), .A2(n8282), .ZN(n8284) );
  AND2_X1 U5568 ( .A1(n8283), .A2(n8282), .ZN(n8285) );
  AND2_X1 U5569 ( .A1(n5752), .A2(n5698), .ZN(n8305) );
  AND2_X1 U5570 ( .A1(n8402), .A2(n4652), .ZN(n8341) );
  NOR2_X1 U5571 ( .A1(n8576), .A2(n4654), .ZN(n4652) );
  NAND2_X1 U5572 ( .A1(n8341), .A2(n8324), .ZN(n8318) );
  OR2_X1 U5573 ( .A1(n8581), .A2(n8375), .ZN(n8280) );
  OR2_X1 U5574 ( .A1(n5582), .A2(n10119), .ZN(n5617) );
  AOI21_X1 U5575 ( .B1(n4757), .B2(n4759), .A(n4756), .ZN(n4755) );
  INV_X1 U5576 ( .A(n4759), .ZN(n4758) );
  INV_X1 U5577 ( .A(n5901), .ZN(n4756) );
  INV_X1 U5578 ( .A(n8350), .ZN(n8353) );
  AND2_X1 U5579 ( .A1(n5623), .A2(n5622), .ZN(n8357) );
  NAND2_X1 U5580 ( .A1(n5906), .A2(n5907), .ZN(n8350) );
  NAND2_X1 U5581 ( .A1(n8351), .A2(n8350), .ZN(n8349) );
  NAND2_X1 U5582 ( .A1(n8402), .A2(n4656), .ZN(n8366) );
  NAND2_X1 U5583 ( .A1(n8402), .A2(n8389), .ZN(n8383) );
  AND2_X1 U5584 ( .A1(n8421), .A2(n8407), .ZN(n8402) );
  NOR2_X1 U5585 ( .A1(n8443), .A2(n8601), .ZN(n8421) );
  AND2_X1 U5586 ( .A1(n5885), .A2(n8436), .ZN(n8460) );
  AOI21_X1 U5587 ( .B1(n4731), .B2(n4735), .A(n4730), .ZN(n4729) );
  NOR2_X1 U5588 ( .A1(n4738), .A2(n8485), .ZN(n4731) );
  NAND2_X1 U5589 ( .A1(n7805), .A2(n4649), .ZN(n8490) );
  AND2_X1 U5590 ( .A1(n4415), .A2(n4989), .ZN(n4649) );
  INV_X1 U5591 ( .A(n5419), .ZN(n5417) );
  NAND2_X1 U5592 ( .A1(n8527), .A2(n5863), .ZN(n8499) );
  AND4_X1 U5593 ( .A1(n5394), .A2(n5393), .A3(n5392), .A4(n5391), .ZN(n8503)
         );
  NAND2_X1 U5594 ( .A1(n8529), .A2(n8528), .ZN(n8527) );
  AND2_X1 U5595 ( .A1(n7805), .A2(n9518), .ZN(n8536) );
  AOI21_X1 U5596 ( .B1(n4750), .B2(n4754), .A(n4749), .ZN(n4748) );
  INV_X1 U5597 ( .A(n5853), .ZN(n4749) );
  NAND2_X1 U5598 ( .A1(n9852), .A2(n4958), .ZN(n8271) );
  NOR2_X1 U5599 ( .A1(n7795), .A2(n4959), .ZN(n4958) );
  INV_X1 U5600 ( .A(n7707), .ZN(n4959) );
  INV_X1 U5601 ( .A(n7751), .ZN(n7755) );
  NAND2_X1 U5602 ( .A1(n4752), .A2(n5932), .ZN(n7756) );
  NAND2_X1 U5603 ( .A1(n4753), .A2(n5931), .ZN(n4752) );
  INV_X1 U5604 ( .A(n7710), .ZN(n4753) );
  AND4_X1 U5605 ( .A1(n5316), .A2(n5315), .A3(n5314), .A4(n5313), .ZN(n7757)
         );
  AND2_X1 U5606 ( .A1(n5932), .A2(n5931), .ZN(n7790) );
  NAND2_X1 U5607 ( .A1(n9852), .A2(n7707), .ZN(n7796) );
  NOR2_X1 U5608 ( .A1(n7513), .A2(n4660), .ZN(n9854) );
  INV_X1 U5609 ( .A(n4662), .ZN(n4660) );
  NAND2_X1 U5610 ( .A1(n7505), .A2(n5835), .ZN(n7563) );
  AND2_X1 U5611 ( .A1(n5242), .A2(n5241), .ZN(n5264) );
  AND2_X1 U5612 ( .A1(n5187), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5242) );
  AND2_X1 U5613 ( .A1(n5836), .A2(n5835), .ZN(n7498) );
  AND4_X1 U5614 ( .A1(n5272), .A2(n5271), .A3(n5270), .A4(n5269), .ZN(n7703)
         );
  NAND2_X1 U5615 ( .A1(n6951), .A2(n6950), .ZN(n7334) );
  NOR2_X1 U5616 ( .A1(n5680), .A2(P2_D_REG_0__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U5617 ( .A1(n5640), .A2(n5639), .ZN(n8569) );
  NAND2_X1 U5618 ( .A1(n5544), .A2(n5543), .ZN(n8594) );
  OR2_X1 U5619 ( .A1(n8507), .A2(n8506), .ZN(n8630) );
  OR2_X1 U5620 ( .A1(n5782), .A2(n6429), .ZN(n5114) );
  NOR2_X1 U5621 ( .A1(n7262), .A2(n6665), .ZN(n6703) );
  NOR2_X1 U5622 ( .A1(n5663), .A2(n4762), .ZN(n4493) );
  NOR2_X1 U5623 ( .A1(n5330), .A2(n5036), .ZN(n5409) );
  AND2_X1 U5624 ( .A1(n4991), .A2(n5145), .ZN(n5303) );
  CLKBUF_X1 U5625 ( .A(n5145), .Z(n5146) );
  CLKBUF_X1 U5626 ( .A(n5103), .Z(n5104) );
  CLKBUF_X1 U5627 ( .A(n5082), .Z(n5083) );
  NAND2_X1 U5628 ( .A1(n6974), .A2(n6975), .ZN(n7133) );
  XOR2_X1 U5629 ( .A(n7982), .B(n7994), .Z(n7965) );
  INV_X1 U5630 ( .A(n8716), .ZN(n4853) );
  NAND2_X1 U5631 ( .A1(n6222), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6233) );
  INV_X1 U5632 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6157) );
  OR2_X1 U5633 ( .A1(n6158), .A2(n6157), .ZN(n6169) );
  AND2_X1 U5634 ( .A1(n6257), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U5635 ( .A1(n7637), .A2(n7636), .ZN(n4875) );
  OR2_X1 U5636 ( .A1(n6196), .A2(n6195), .ZN(n6209) );
  NOR2_X1 U5637 ( .A1(n4851), .A2(n4847), .ZN(n4846) );
  NAND2_X1 U5638 ( .A1(n4848), .A2(n7937), .ZN(n4847) );
  AND2_X1 U5639 ( .A1(n4844), .A2(n7938), .ZN(n4622) );
  OR2_X1 U5640 ( .A1(n6169), .A2(n7252), .ZN(n6182) );
  NOR2_X1 U5641 ( .A1(n6182), .A2(n6181), .ZN(n6184) );
  AND3_X1 U5642 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6115) );
  CLKBUF_X1 U5643 ( .A(n7120), .Z(n6984) );
  NAND2_X1 U5644 ( .A1(n4858), .A2(n4862), .ZN(n4857) );
  INV_X1 U5645 ( .A(n4860), .ZN(n4858) );
  AND2_X1 U5646 ( .A1(n4859), .A2(n7905), .ZN(n4856) );
  NOR2_X1 U5647 ( .A1(n8951), .A2(n4601), .ZN(n4600) );
  OAI21_X1 U5648 ( .B1(n9363), .B2(n8949), .A(n8943), .ZN(n4601) );
  NAND2_X1 U5649 ( .A1(n8945), .A2(n4470), .ZN(n4598) );
  NOR2_X1 U5650 ( .A1(n9017), .A2(n8954), .ZN(n4885) );
  INV_X1 U5651 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5974) );
  NOR2_X1 U5652 ( .A1(n9577), .A2(n6478), .ZN(n9598) );
  OR2_X1 U5653 ( .A1(n9085), .A2(n9086), .ZN(n9098) );
  NOR3_X1 U5654 ( .A1(n9164), .A2(n4704), .A3(n9117), .ZN(n9116) );
  NOR2_X1 U5655 ( .A1(n9142), .A2(n8006), .ZN(n9124) );
  AND2_X1 U5656 ( .A1(n6330), .A2(n6321), .ZN(n9144) );
  OR2_X1 U5657 ( .A1(n9164), .A2(n9370), .ZN(n9142) );
  OR2_X1 U5658 ( .A1(n9176), .A2(n9155), .ZN(n9158) );
  AND2_X1 U5659 ( .A1(n9178), .A2(n8932), .ZN(n9176) );
  NAND2_X1 U5660 ( .A1(n4525), .A2(n4530), .ZN(n9242) );
  NAND2_X1 U5661 ( .A1(n9258), .A2(n8962), .ZN(n4525) );
  AND2_X1 U5662 ( .A1(n8963), .A2(n8962), .ZN(n9257) );
  NAND2_X1 U5663 ( .A1(n9274), .A2(n9276), .ZN(n9273) );
  AND2_X1 U5664 ( .A1(n8911), .A2(n8914), .ZN(n9276) );
  OR2_X1 U5665 ( .A1(n6233), .A2(n8699), .ZN(n6235) );
  NOR2_X1 U5666 ( .A1(n6235), .A2(n6019), .ZN(n6246) );
  AOI21_X1 U5667 ( .B1(n9311), .B2(n6240), .A(n4936), .ZN(n9298) );
  NOR2_X1 U5668 ( .A1(n9428), .A2(n9541), .ZN(n4936) );
  AND2_X1 U5669 ( .A1(n9292), .A2(n8905), .ZN(n9310) );
  AND2_X1 U5670 ( .A1(n9539), .A2(n9431), .ZN(n4937) );
  OR2_X1 U5671 ( .A1(n7824), .A2(n9432), .ZN(n6215) );
  NAND2_X1 U5672 ( .A1(n4503), .A2(n4502), .ZN(n7546) );
  AOI21_X1 U5673 ( .B1(n4504), .B2(n4506), .A(n8887), .ZN(n4502) );
  INV_X1 U5674 ( .A(n8872), .ZN(n4506) );
  NAND2_X1 U5675 ( .A1(n7376), .A2(n8869), .ZN(n7477) );
  NAND2_X1 U5676 ( .A1(n7379), .A2(n4689), .ZN(n7482) );
  NAND2_X1 U5677 ( .A1(n7379), .A2(n7385), .ZN(n7484) );
  AND2_X1 U5678 ( .A1(n8869), .A2(n8871), .ZN(n7377) );
  NAND2_X1 U5679 ( .A1(n4817), .A2(n8974), .ZN(n4816) );
  NAND2_X1 U5680 ( .A1(n4451), .A2(n6364), .ZN(n4515) );
  OR2_X1 U5681 ( .A1(n7085), .A2(n6150), .ZN(n7086) );
  NAND2_X1 U5682 ( .A1(n4685), .A2(n4684), .ZN(n7158) );
  INV_X1 U5683 ( .A(n9796), .ZN(n4684) );
  INV_X1 U5684 ( .A(n7094), .ZN(n4685) );
  INV_X1 U5685 ( .A(n6150), .ZN(n8982) );
  OAI21_X1 U5686 ( .B1(n9765), .B2(n4945), .A(n4943), .ZN(n6139) );
  OR2_X1 U5687 ( .A1(n7028), .A2(n7124), .ZN(n7094) );
  NAND2_X1 U5688 ( .A1(n9765), .A2(n4431), .ZN(n6892) );
  NAND2_X1 U5689 ( .A1(n6938), .A2(n6988), .ZN(n7028) );
  NOR2_X1 U5690 ( .A1(n6780), .A2(n6785), .ZN(n6940) );
  AND2_X1 U5691 ( .A1(n9763), .A2(n6940), .ZN(n6938) );
  AND2_X1 U5692 ( .A1(n6348), .A2(n6698), .ZN(n9695) );
  CLKBUF_X1 U5693 ( .A(n8966), .Z(n9705) );
  NAND2_X1 U5694 ( .A1(n6308), .A2(n6307), .ZN(n9166) );
  NAND2_X1 U5695 ( .A1(n6368), .A2(n8961), .ZN(n9210) );
  NAND2_X1 U5696 ( .A1(n4524), .A2(n4526), .ZN(n6368) );
  INV_X1 U5697 ( .A(n9789), .ZN(n9759) );
  OR2_X1 U5698 ( .A1(n8949), .A2(n9025), .ZN(n9801) );
  NAND2_X1 U5699 ( .A1(n6243), .A2(n9060), .ZN(n4808) );
  INV_X1 U5700 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4953) );
  XNOR2_X1 U5701 ( .A(n5759), .B(n5749), .ZN(n8781) );
  NAND2_X1 U5702 ( .A1(n5987), .A2(n4954), .ZN(n6001) );
  AND2_X1 U5703 ( .A1(n5004), .A2(n4955), .ZN(n4954) );
  INV_X1 U5704 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4955) );
  XNOR2_X1 U5705 ( .A(n5738), .B(n5737), .ZN(n7743) );
  XNOR2_X1 U5706 ( .A(n5631), .B(n5630), .ZN(n7700) );
  XNOR2_X1 U5707 ( .A(n5609), .B(n5608), .ZN(n7681) );
  NAND2_X1 U5708 ( .A1(n5987), .A2(n6351), .ZN(n6390) );
  AND2_X1 U5709 ( .A1(n6355), .A2(n6350), .ZN(n9021) );
  OR2_X1 U5710 ( .A1(n6204), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U5711 ( .A1(n4683), .A2(n5281), .ZN(n5296) );
  NAND2_X1 U5712 ( .A1(n5280), .A2(n5001), .ZN(n4683) );
  XNOR2_X1 U5713 ( .A(n4538), .B(n5002), .ZN(n6455) );
  OAI21_X1 U5714 ( .B1(n5227), .B2(n5226), .A(n5228), .ZN(n4538) );
  INV_X1 U5715 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6010) );
  NOR2_X2 U5716 ( .A1(n6106), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6009) );
  XNOR2_X1 U5717 ( .A(n5384), .B(n5383), .ZN(n8031) );
  NAND2_X1 U5718 ( .A1(n7539), .A2(n5764), .ZN(n5568) );
  AND2_X1 U5719 ( .A1(n5278), .A2(n7312), .ZN(n4799) );
  NAND2_X1 U5720 ( .A1(n4800), .A2(n7312), .ZN(n9828) );
  NAND2_X1 U5721 ( .A1(n5477), .A2(n5476), .ZN(n8611) );
  NAND2_X1 U5722 ( .A1(n5741), .A2(n5740), .ZN(n8564) );
  AOI21_X1 U5723 ( .B1(n6671), .B2(n9922), .A(n5076), .ZN(n7972) );
  NAND2_X1 U5724 ( .A1(n4788), .A2(n5077), .ZN(n7971) );
  INV_X1 U5725 ( .A(n4789), .ZN(n4788) );
  AND3_X1 U5726 ( .A1(n5553), .A2(n5552), .A3(n5551), .ZN(n8429) );
  AND4_X1 U5727 ( .A1(n5510), .A2(n5509), .A3(n5508), .A4(n5507), .ZN(n8428)
         );
  AND4_X1 U5728 ( .A1(n5360), .A2(n5359), .A3(n5358), .A4(n5357), .ZN(n8032)
         );
  NAND2_X1 U5729 ( .A1(n7628), .A2(n5293), .ZN(n7673) );
  NAND2_X1 U5730 ( .A1(n5591), .A2(n5590), .ZN(n8085) );
  NAND2_X1 U5731 ( .A1(n7034), .A2(n5139), .ZN(n6921) );
  AOI21_X1 U5732 ( .B1(n4774), .B2(n4776), .A(n4442), .ZN(n4772) );
  NAND2_X1 U5733 ( .A1(n4494), .A2(n5494), .ZN(n8114) );
  NAND2_X1 U5734 ( .A1(n5503), .A2(n5502), .ZN(n8605) );
  NAND2_X1 U5735 ( .A1(n7630), .A2(n7629), .ZN(n7628) );
  AND4_X2 U5736 ( .A1(n5034), .A2(n5033), .A3(n5032), .A4(n5035), .ZN(n8024)
         );
  NAND2_X1 U5737 ( .A1(n4408), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5032) );
  NAND2_X1 U5738 ( .A1(n5457), .A2(n5456), .ZN(n8615) );
  OR2_X1 U5739 ( .A1(n7978), .A2(n9921), .ZN(n9829) );
  NAND2_X1 U5740 ( .A1(n4674), .A2(n4672), .ZN(n8139) );
  AND2_X1 U5741 ( .A1(n5704), .A2(n5690), .ZN(n8138) );
  AND4_X1 U5742 ( .A1(n5346), .A2(n5345), .A3(n5344), .A4(n5343), .ZN(n8155)
         );
  AND4_X1 U5743 ( .A1(n5424), .A2(n5423), .A3(n5422), .A4(n5421), .ZN(n8154)
         );
  OR2_X1 U5744 ( .A1(n8142), .A2(n8500), .ZN(n9832) );
  OR2_X1 U5745 ( .A1(n8142), .A2(n8502), .ZN(n9831) );
  AND2_X1 U5746 ( .A1(n5388), .A2(n5387), .ZN(n8148) );
  INV_X1 U5747 ( .A(n9829), .ZN(n8158) );
  INV_X1 U5748 ( .A(P2_U3966), .ZN(n8177) );
  INV_X1 U5749 ( .A(n4719), .ZN(n6819) );
  NAND2_X1 U5750 ( .A1(n6820), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4718) );
  NOR2_X1 U5751 ( .A1(n6847), .A2(n4710), .ZN(n6859) );
  AND2_X1 U5752 ( .A1(n6851), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4710) );
  NOR2_X1 U5753 ( .A1(n6859), .A2(n6858), .ZN(n6857) );
  NOR2_X1 U5754 ( .A1(n6857), .A2(n4709), .ZN(n6823) );
  AND2_X1 U5755 ( .A1(n6862), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4709) );
  NOR2_X1 U5756 ( .A1(n6823), .A2(n6822), .ZN(n6835) );
  NOR2_X1 U5757 ( .A1(n6872), .A2(n4712), .ZN(n6887) );
  AND2_X1 U5758 ( .A1(n6873), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4712) );
  NOR2_X1 U5759 ( .A1(n6887), .A2(n6886), .ZN(n6885) );
  NOR2_X1 U5760 ( .A1(n6885), .A2(n4711), .ZN(n6876) );
  AND2_X1 U5761 ( .A1(n6890), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4711) );
  NOR2_X1 U5762 ( .A1(n6876), .A2(n6875), .ZN(n7075) );
  AND2_X1 U5763 ( .A1(n6731), .A2(n8646), .ZN(n8256) );
  XNOR2_X1 U5764 ( .A(n4647), .B(n8556), .ZN(n8558) );
  NAND2_X1 U5765 ( .A1(n4769), .A2(n4768), .ZN(n4767) );
  NAND2_X1 U5766 ( .A1(n8310), .A2(n8533), .ZN(n4769) );
  INV_X1 U5767 ( .A(n8569), .ZN(n8324) );
  NAND2_X1 U5768 ( .A1(n8393), .A2(n4759), .ZN(n8372) );
  OAI21_X1 U5769 ( .B1(n8420), .B2(n4971), .A(n4968), .ZN(n8381) );
  NAND2_X1 U5770 ( .A1(n4967), .A2(n4972), .ZN(n8382) );
  NAND2_X1 U5771 ( .A1(n8420), .A2(n4973), .ZN(n4967) );
  INV_X1 U5772 ( .A(n8594), .ZN(n8407) );
  AND2_X1 U5773 ( .A1(n4974), .A2(n4435), .ZN(n8401) );
  NAND2_X1 U5774 ( .A1(n8420), .A2(n8278), .ZN(n4974) );
  AND2_X1 U5775 ( .A1(n5520), .A2(n5519), .ZN(n8423) );
  NAND2_X1 U5776 ( .A1(n8482), .A2(n4988), .ZN(n8467) );
  NAND2_X1 U5777 ( .A1(n4728), .A2(n4735), .ZN(n8486) );
  OR2_X1 U5778 ( .A1(n8529), .A2(n4737), .ZN(n4728) );
  NOR2_X1 U5779 ( .A1(n8507), .A2(n4990), .ZN(n8483) );
  NAND2_X1 U5780 ( .A1(n7805), .A2(n4651), .ZN(n8512) );
  NAND2_X1 U5781 ( .A1(n7559), .A2(n7558), .ZN(n7560) );
  INV_X1 U5782 ( .A(n9899), .ZN(n7517) );
  NAND2_X1 U5783 ( .A1(n7337), .A2(n5825), .ZN(n7275) );
  OAI21_X1 U5784 ( .B1(n7260), .B2(n4981), .A(n4979), .ZN(n7355) );
  NAND2_X1 U5785 ( .A1(n7260), .A2(n7259), .ZN(n7350) );
  NAND2_X1 U5786 ( .A1(n7332), .A2(n6952), .ZN(n6953) );
  OR2_X1 U5787 ( .A1(n9855), .A2(n9922), .ZN(n8551) );
  OR2_X1 U5788 ( .A1(n5106), .A2(n6434), .ZN(n5093) );
  INV_X1 U5789 ( .A(n8496), .ZN(n9847) );
  INV_X1 U5790 ( .A(n8551), .ZN(n8520) );
  NAND2_X1 U5791 ( .A1(n8549), .A2(n7267), .ZN(n8543) );
  AND2_X2 U5792 ( .A1(n6703), .A2(n7270), .ZN(n9945) );
  AOI211_X1 U5793 ( .C1(n9853), .C2(n9511), .A(n9510), .B(n9509), .ZN(n9532)
         );
  INV_X1 U5794 ( .A(n8562), .ZN(n4585) );
  AND2_X2 U5795 ( .A1(n6703), .A2(n7263), .ZN(n9930) );
  AND2_X1 U5796 ( .A1(n5966), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9868) );
  INV_X1 U5797 ( .A(n9863), .ZN(n9865) );
  NAND2_X1 U5798 ( .A1(n5023), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5022) );
  NAND2_X1 U5799 ( .A1(n5686), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5670) );
  INV_X1 U5800 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n10195) );
  INV_X1 U5801 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7308) );
  INV_X1 U5802 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4499) );
  INV_X1 U5803 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7311) );
  NAND2_X1 U5804 ( .A1(n5049), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5039) );
  INV_X1 U5805 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7045) );
  INV_X1 U5806 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6539) );
  INV_X1 U5807 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6511) );
  INV_X1 U5808 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6456) );
  OR2_X1 U5809 ( .A1(n5238), .A2(n5237), .ZN(n6874) );
  INV_X1 U5810 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6442) );
  INV_X1 U5811 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6439) );
  INV_X1 U5812 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6444) );
  XNOR2_X1 U5813 ( .A(n5057), .B(n5058), .ZN(n6735) );
  NAND2_X1 U5814 ( .A1(n4832), .A2(n7132), .ZN(n7181) );
  NAND2_X1 U5815 ( .A1(n6984), .A2(n7133), .ZN(n4832) );
  NOR2_X1 U5816 ( .A1(n4496), .A2(n7818), .ZN(n7900) );
  AND2_X1 U5817 ( .A1(n4496), .A2(n7818), .ZN(n7906) );
  CLKBUF_X1 U5819 ( .A(n7521), .Z(n7240) );
  NAND2_X1 U5820 ( .A1(n4630), .A2(n4629), .ZN(n8010) );
  AOI21_X1 U5821 ( .B1(n4631), .B2(n4633), .A(n4475), .ZN(n4629) );
  AND2_X1 U5822 ( .A1(n4854), .A2(n4853), .ZN(n8674) );
  NAND2_X1 U5823 ( .A1(n4843), .A2(n8715), .ZN(n4854) );
  AND2_X1 U5824 ( .A1(n4877), .A2(n6766), .ZN(n6768) );
  NAND2_X1 U5825 ( .A1(n4871), .A2(n7943), .ZN(n8707) );
  INV_X1 U5826 ( .A(n9778), .ZN(n7300) );
  NAND2_X1 U5827 ( .A1(n6256), .A2(n6255), .ZN(n9265) );
  OAI21_X1 U5828 ( .B1(n6599), .B2(n6693), .A(n9301), .ZN(n8730) );
  NAND2_X1 U5829 ( .A1(n4498), .A2(n4497), .ZN(n5006) );
  INV_X1 U5830 ( .A(n6591), .ZN(n4497) );
  INV_X1 U5831 ( .A(n6592), .ZN(n4498) );
  INV_X1 U5832 ( .A(n6628), .ZN(n6583) );
  OR2_X1 U5833 ( .A1(n7914), .A2(n7913), .ZN(n4855) );
  INV_X1 U5834 ( .A(n9793), .ZN(n7188) );
  INV_X1 U5835 ( .A(n8759), .ZN(n8739) );
  NAND2_X1 U5836 ( .A1(n4884), .A2(n4618), .ZN(n4617) );
  NAND2_X1 U5837 ( .A1(n4885), .A2(n4886), .ZN(n4618) );
  INV_X1 U5838 ( .A(n8955), .ZN(n4886) );
  NAND2_X1 U5839 ( .A1(n9026), .A2(n6348), .ZN(n4883) );
  NAND2_X1 U5840 ( .A1(n6087), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6091) );
  NOR2_X1 U5841 ( .A1(n6651), .A2(n6650), .ZN(n9627) );
  NOR2_X1 U5842 ( .A1(n6655), .A2(n9654), .ZN(n7055) );
  AOI21_X1 U5843 ( .B1(n7203), .B2(n7202), .A(n7201), .ZN(n7206) );
  AOI21_X1 U5844 ( .B1(n9071), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9070), .ZN(
        n9073) );
  NAND2_X1 U5845 ( .A1(n4413), .A2(n4513), .ZN(n4508) );
  NAND2_X1 U5846 ( .A1(n6370), .A2(n4421), .ZN(n4507) );
  NAND2_X1 U5847 ( .A1(n4826), .A2(n4827), .ZN(n9146) );
  OAI21_X1 U5848 ( .B1(n9192), .B2(n4928), .A(n4927), .ZN(n9154) );
  NAND2_X1 U5849 ( .A1(n4929), .A2(n6297), .ZN(n9174) );
  NAND2_X1 U5850 ( .A1(n9192), .A2(n4429), .ZN(n4929) );
  NAND2_X1 U5851 ( .A1(n4812), .A2(n4813), .ZN(n9193) );
  NAND2_X1 U5852 ( .A1(n6287), .A2(n6286), .ZN(n9220) );
  NAND2_X1 U5853 ( .A1(n9238), .A2(n4996), .ZN(n9223) );
  NAND2_X1 U5854 ( .A1(n6268), .A2(n6267), .ZN(n9249) );
  NAND2_X1 U5855 ( .A1(n6018), .A2(n6017), .ZN(n9421) );
  NAND2_X1 U5856 ( .A1(n9330), .A2(n8788), .ZN(n9293) );
  NAND2_X1 U5857 ( .A1(n7688), .A2(n8894), .ZN(n7771) );
  NAND2_X1 U5858 ( .A1(n6219), .A2(n6218), .ZN(n8768) );
  INV_X1 U5859 ( .A(n4951), .ZN(n7548) );
  AND2_X1 U5860 ( .A1(n7475), .A2(n4949), .ZN(n7465) );
  NAND2_X1 U5861 ( .A1(n9716), .A2(n9699), .ZN(n9326) );
  NAND2_X1 U5862 ( .A1(n7088), .A2(n6152), .ZN(n7157) );
  NAND2_X1 U5863 ( .A1(n6894), .A2(n8974), .ZN(n7022) );
  NAND2_X1 U5864 ( .A1(n6364), .A2(n8849), .ZN(n6941) );
  NAND2_X1 U5865 ( .A1(n6243), .A2(n4687), .ZN(n4686) );
  INV_X1 U5866 ( .A(n9594), .ZN(n4687) );
  INV_X1 U5867 ( .A(n9215), .ZN(n9704) );
  NAND2_X1 U5868 ( .A1(n9719), .A2(n6554), .ZN(n9301) );
  INV_X1 U5869 ( .A(n9326), .ZN(n9347) );
  INV_X2 U5870 ( .A(n10187), .ZN(n10189) );
  INV_X1 U5871 ( .A(n9110), .ZN(n9443) );
  INV_X1 U5872 ( .A(n9220), .ZN(n9464) );
  INV_X1 U5873 ( .A(n9249), .ZN(n9471) );
  INV_X2 U5874 ( .A(n9807), .ZN(n9809) );
  INV_X1 U5875 ( .A(n9720), .ZN(n9721) );
  XNOR2_X1 U5876 ( .A(n5781), .B(n5780), .ZN(n8771) );
  NAND2_X1 U5877 ( .A1(n4412), .A2(n6384), .ZN(n6388) );
  NOR2_X1 U5878 ( .A1(n6386), .A2(n6385), .ZN(n6387) );
  NOR2_X1 U5879 ( .A1(n5985), .A2(n6121), .ZN(n6384) );
  NAND2_X1 U5880 ( .A1(n4838), .A2(n4412), .ZN(n7748) );
  MUX2_X1 U5881 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4839), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n4838) );
  INV_X1 U5882 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10172) );
  XNOR2_X1 U5883 ( .A(n4837), .B(n6383), .ZN(n7600) );
  INV_X1 U5884 ( .A(n4640), .ZN(n4638) );
  INV_X1 U5885 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7405) );
  INV_X1 U5886 ( .A(n9021), .ZN(n8954) );
  INV_X1 U5887 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7215) );
  CLKBUF_X1 U5888 ( .A(n6356), .Z(n6348) );
  INV_X1 U5889 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7139) );
  AND2_X1 U5890 ( .A1(n6192), .A2(n6204), .ZN(n9668) );
  INV_X1 U5891 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6532) );
  INV_X1 U5892 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10261) );
  INV_X1 U5893 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6457) );
  INV_X1 U5894 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6453) );
  INV_X1 U5895 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6440) );
  NAND2_X1 U5896 ( .A1(n4882), .A2(n5173), .ZN(n5196) );
  NAND2_X1 U5897 ( .A1(n5170), .A2(n5169), .ZN(n4882) );
  INV_X1 U5898 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6437) );
  XNOR2_X1 U5899 ( .A(n5170), .B(n5169), .ZN(n6438) );
  INV_X1 U5900 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10262) );
  NAND2_X1 U5901 ( .A1(n4667), .A2(n5133), .ZN(n5151) );
  NOR2_X1 U5902 ( .A1(n7441), .A2(n10288), .ZN(n9973) );
  AOI21_X1 U5903 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9971), .ZN(n9970) );
  NOR2_X1 U5904 ( .A1(n9970), .A2(n9969), .ZN(n9968) );
  NAND2_X1 U5905 ( .A1(n7100), .A2(n5186), .ZN(n7110) );
  NAND2_X1 U5906 ( .A1(n4773), .A2(n4777), .ZN(n7170) );
  NAND2_X1 U5907 ( .A1(n5119), .A2(n5118), .ZN(n7037) );
  OAI21_X1 U5908 ( .B1(n8259), .B2(n5050), .A(n4713), .ZN(P2_U3264) );
  AOI21_X1 U5909 ( .B1(n4715), .B2(n5050), .A(n4714), .ZN(n4713) );
  NAND2_X1 U5910 ( .A1(n7335), .A2(n4726), .ZN(P2_U3293) );
  AND2_X1 U5911 ( .A1(n7336), .A2(n4482), .ZN(n4726) );
  NAND2_X1 U5912 ( .A1(n4745), .A2(n4744), .ZN(P2_U3549) );
  OR2_X1 U5913 ( .A1(n9945), .A2(n10254), .ZN(n4744) );
  NAND2_X1 U5914 ( .A1(n8632), .A2(n9945), .ZN(n4745) );
  OAI222_X1 U5915 ( .A1(n8651), .A2(n7683), .B1(n8025), .B2(n7747), .C1(
        P2_U3152), .C2(n7682), .ZN(P2_U3333) );
  OAI222_X1 U5916 ( .A1(n8651), .A2(n10195), .B1(n8025), .B2(n7406), .C1(n7404), .C2(n8130), .ZN(P2_U3336) );
  OAI222_X1 U5917 ( .A1(n8651), .A2(n7308), .B1(P2_U3152), .B2(n7307), .C1(
        n8025), .C2(n7306), .ZN(P2_U3337) );
  OAI222_X1 U5918 ( .A1(n8651), .A2(n7311), .B1(n8130), .B2(n7310), .C1(n8025), 
        .C2(n7309), .ZN(P2_U3338) );
  OAI222_X1 U5919 ( .A1(n8651), .A2(n7045), .B1(n8025), .B2(n7140), .C1(n7451), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI222_X1 U5920 ( .A1(n8651), .A2(n6689), .B1(n8025), .B2(n6688), .C1(n8130), 
        .C2(n7726), .ZN(P2_U3343) );
  OAI222_X1 U5921 ( .A1(n8651), .A2(n6543), .B1(n8025), .B2(n6544), .C1(n7609), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  OAI222_X1 U5922 ( .A1(n8651), .A2(n6539), .B1(n8025), .B2(n6540), .C1(n7155), 
        .C2(n8130), .ZN(P2_U3345) );
  OAI222_X1 U5923 ( .A1(n8651), .A2(n10015), .B1(n8025), .B2(n6531), .C1(
        P2_U3152), .C2(n6530), .ZN(P2_U3346) );
  OAI222_X1 U5924 ( .A1(n8651), .A2(n6511), .B1(n8025), .B2(n6510), .C1(n7077), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  OAI222_X1 U5925 ( .A1(n8651), .A2(n6456), .B1(n8025), .B2(n6458), .C1(n6874), 
        .C2(n8130), .ZN(P2_U3349) );
  OAI222_X1 U5926 ( .A1(n8651), .A2(n6450), .B1(n8025), .B2(n6449), .C1(n8130), 
        .C2(n6448), .ZN(P2_U3351) );
  NAND2_X1 U5927 ( .A1(n4868), .A2(n8744), .ZN(n4865) );
  AND2_X1 U5928 ( .A1(n8750), .A2(n4478), .ZN(n4492) );
  AOI21_X1 U5929 ( .B1(n4635), .B2(n4469), .A(n8746), .ZN(n4489) );
  MUX2_X1 U5930 ( .A(n9106), .B(n9105), .S(n9215), .Z(n9107) );
  OR2_X1 U5931 ( .A1(n9185), .A2(n9161), .ZN(n4409) );
  AND2_X1 U5932 ( .A1(n6933), .A2(n8849), .ZN(n4410) );
  AND2_X1 U5933 ( .A1(n4706), .A2(n4705), .ZN(n4411) );
  AND2_X1 U5934 ( .A1(n6498), .A2(n5061), .ZN(n6134) );
  NAND2_X1 U5935 ( .A1(n5987), .A2(n4636), .ZN(n4412) );
  AND2_X1 U5936 ( .A1(n4509), .A2(n9706), .ZN(n4413) );
  AND2_X1 U5937 ( .A1(n9331), .A2(n8803), .ZN(n4414) );
  OR2_X1 U5938 ( .A1(n9370), .A2(n7875), .ZN(n9010) );
  INV_X1 U5939 ( .A(n7184), .ZN(n4830) );
  AND2_X1 U5940 ( .A1(n4651), .A2(n4650), .ZN(n4415) );
  INV_X1 U5941 ( .A(n8485), .ZN(n4734) );
  INV_X1 U5942 ( .A(n8391), .ZN(n4969) );
  AND2_X1 U5943 ( .A1(n6313), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4416) );
  AND3_X1 U5944 ( .A1(n4450), .A2(n8957), .A3(n8932), .ZN(n4417) );
  INV_X1 U5945 ( .A(n7354), .ZN(n4978) );
  NAND2_X1 U5946 ( .A1(n6232), .A2(n6231), .ZN(n9428) );
  AND2_X1 U5947 ( .A1(n4689), .A2(n4688), .ZN(n4418) );
  AND2_X1 U5948 ( .A1(n4748), .A2(n7801), .ZN(n4419) );
  NAND2_X1 U5949 ( .A1(n5614), .A2(n5613), .ZN(n8576) );
  INV_X1 U5950 ( .A(n9185), .ZN(n9456) );
  NAND2_X1 U5951 ( .A1(n6299), .A2(n6298), .ZN(n9185) );
  AND2_X1 U5952 ( .A1(n4699), .A2(n4702), .ZN(n4420) );
  AND2_X1 U5953 ( .A1(n4413), .A2(n4444), .ZN(n4421) );
  OR2_X1 U5954 ( .A1(n4803), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n4422) );
  NAND2_X1 U5955 ( .A1(n9173), .A2(n4462), .ZN(n4423) );
  NOR2_X1 U5956 ( .A1(n7755), .A2(n4751), .ZN(n4750) );
  NAND2_X1 U5957 ( .A1(n4885), .A2(n7407), .ZN(n4424) );
  INV_X1 U5958 ( .A(n8006), .ZN(n4706) );
  AND2_X1 U5959 ( .A1(n4891), .A2(n4486), .ZN(n4425) );
  INV_X1 U5960 ( .A(n6590), .ZN(n7941) );
  NAND2_X1 U5961 ( .A1(n5148), .A2(n10198), .ZN(n5175) );
  AND2_X1 U5962 ( .A1(n4786), .A2(n7672), .ZN(n4426) );
  NAND2_X1 U5963 ( .A1(n6077), .A2(n5974), .ZN(n6079) );
  NAND2_X1 U5964 ( .A1(n5083), .A2(n5008), .ZN(n5086) );
  AND2_X1 U5965 ( .A1(n4938), .A2(n4939), .ZN(n4427) );
  AND2_X1 U5966 ( .A1(n8946), .A2(n8779), .ZN(n4428) );
  OR2_X1 U5967 ( .A1(n9460), .A2(n8659), .ZN(n4429) );
  INV_X1 U5968 ( .A(n9492), .ZN(n5991) );
  NAND2_X1 U5969 ( .A1(n7843), .A2(n4604), .ZN(n9492) );
  INV_X1 U5970 ( .A(n5987), .ZN(n6350) );
  AND2_X1 U5971 ( .A1(n5146), .A2(n5009), .ZN(n5148) );
  INV_X1 U5972 ( .A(n7645), .ZN(n7671) );
  NAND2_X1 U5973 ( .A1(n6194), .A2(n6193), .ZN(n7645) );
  INV_X1 U5974 ( .A(n9117), .ZN(n9447) );
  NAND2_X1 U5975 ( .A1(n8778), .A2(n8777), .ZN(n9117) );
  INV_X1 U5976 ( .A(n8986), .ZN(n4947) );
  AND2_X1 U5977 ( .A1(n6893), .A2(n6114), .ZN(n4431) );
  AND2_X1 U5978 ( .A1(n7233), .A2(n9792), .ZN(n4432) );
  AND2_X1 U5979 ( .A1(n5910), .A2(n5922), .ZN(n4433) );
  INV_X1 U5980 ( .A(n8825), .ZN(n4823) );
  NAND2_X1 U5981 ( .A1(n6008), .A2(n6007), .ZN(n9199) );
  NOR2_X1 U5982 ( .A1(n9166), .A2(n9180), .ZN(n4434) );
  NAND2_X1 U5983 ( .A1(n5024), .A2(n5025), .ZN(n5023) );
  NAND2_X1 U5984 ( .A1(n8601), .A2(n8438), .ZN(n4435) );
  AND2_X1 U5985 ( .A1(n4719), .A2(n4718), .ZN(n4436) );
  NOR2_X1 U5986 ( .A1(n7965), .A2(n4477), .ZN(n4437) );
  AND2_X1 U5987 ( .A1(n6097), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n4438) );
  NAND2_X1 U5988 ( .A1(n6168), .A2(n6167), .ZN(n7392) );
  NAND2_X1 U5989 ( .A1(n5263), .A2(n5262), .ZN(n7704) );
  INV_X1 U5990 ( .A(n7905), .ZN(n4862) );
  INV_X1 U5991 ( .A(n8589), .ZN(n8389) );
  NAND2_X1 U5992 ( .A1(n5568), .A2(n5567), .ZN(n8589) );
  NAND2_X1 U5993 ( .A1(n8402), .A2(n4653), .ZN(n4657) );
  NAND2_X1 U5994 ( .A1(n9248), .A2(n4692), .ZN(n4696) );
  NAND2_X1 U5995 ( .A1(n5376), .A2(n5375), .ZN(n8538) );
  XNOR2_X1 U5996 ( .A(n5364), .B(n10080), .ZN(n5363) );
  INV_X1 U5997 ( .A(n4703), .ZN(n9125) );
  OR2_X1 U5998 ( .A1(n9164), .A2(n4704), .ZN(n4703) );
  INV_X1 U5999 ( .A(n4738), .ZN(n4737) );
  NOR2_X1 U6000 ( .A1(n5727), .A2(n4739), .ZN(n4738) );
  AND2_X1 U6001 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n4439) );
  NAND2_X1 U6002 ( .A1(n5798), .A2(n5815), .ZN(n7333) );
  AND2_X1 U6003 ( .A1(n5858), .A2(n5857), .ZN(n7801) );
  INV_X1 U6004 ( .A(n4522), .ZN(n4521) );
  OAI21_X1 U6005 ( .B1(n6366), .B2(n4523), .A(n8991), .ZN(n4522) );
  AND2_X1 U6006 ( .A1(n4826), .A2(n4824), .ZN(n4440) );
  INV_X1 U6007 ( .A(n5931), .ZN(n4754) );
  AND2_X1 U6008 ( .A1(n4526), .A2(n8959), .ZN(n4441) );
  INV_X1 U6009 ( .A(n9127), .ZN(n9363) );
  NAND2_X1 U6010 ( .A1(n8783), .A2(n8782), .ZN(n9127) );
  INV_X1 U6011 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6391) );
  AND2_X1 U6012 ( .A1(n5225), .A2(n5224), .ZN(n4442) );
  AND2_X1 U6013 ( .A1(n4426), .A2(n4787), .ZN(n4443) );
  NAND2_X1 U6014 ( .A1(n6338), .A2(n9135), .ZN(n4444) );
  INV_X1 U6015 ( .A(n4654), .ZN(n4653) );
  NAND2_X1 U6016 ( .A1(n4656), .A2(n4655), .ZN(n4654) );
  INV_X1 U6017 ( .A(n4693), .ZN(n4692) );
  NAND2_X1 U6018 ( .A1(n4694), .A2(n9460), .ZN(n4693) );
  INV_X1 U6019 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6383) );
  INV_X1 U6020 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5015) );
  OR2_X1 U6021 ( .A1(n4928), .A2(n4434), .ZN(n4445) );
  AND2_X1 U6022 ( .A1(n5298), .A2(SI_11_), .ZN(n4446) );
  AND2_X1 U6023 ( .A1(n5153), .A2(SI_4_), .ZN(n4447) );
  AND2_X1 U6024 ( .A1(n5198), .A2(SI_6_), .ZN(n4448) );
  NAND2_X1 U6025 ( .A1(n7259), .A2(n7349), .ZN(n4449) );
  AND2_X1 U6026 ( .A1(n8902), .A2(n9312), .ZN(n9331) );
  AND3_X1 U6027 ( .A1(n8958), .A2(n8944), .A3(n8961), .ZN(n4450) );
  AND2_X1 U6028 ( .A1(n4410), .A2(n8974), .ZN(n4451) );
  NAND2_X1 U6029 ( .A1(n8279), .A2(n4435), .ZN(n4452) );
  INV_X1 U6030 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n10198) );
  OR2_X1 U6031 ( .A1(n8622), .A2(n8501), .ZN(n5869) );
  INV_X1 U6032 ( .A(n5869), .ZN(n4730) );
  NAND2_X1 U6033 ( .A1(n9010), .A2(n8835), .ZN(n9147) );
  INV_X1 U6034 ( .A(n9147), .ZN(n4825) );
  AND2_X1 U6035 ( .A1(n4813), .A2(n8957), .ZN(n4453) );
  AND2_X1 U6036 ( .A1(n4678), .A2(n4676), .ZN(n4454) );
  INV_X1 U6037 ( .A(n5002), .ZN(n4571) );
  AND2_X1 U6038 ( .A1(n4558), .A2(n5363), .ZN(n4455) );
  AND2_X1 U6039 ( .A1(n5138), .A2(n5118), .ZN(n4456) );
  AND2_X1 U6040 ( .A1(n5725), .A2(n7558), .ZN(n4457) );
  AND2_X1 U6041 ( .A1(n7529), .A2(n7522), .ZN(n4458) );
  NOR2_X1 U6042 ( .A1(n4522), .A2(n4811), .ZN(n4518) );
  AND2_X1 U6043 ( .A1(n4746), .A2(n4585), .ZN(n4459) );
  AND2_X1 U6044 ( .A1(n8393), .A2(n5896), .ZN(n4460) );
  AND2_X1 U6045 ( .A1(n4956), .A2(n4953), .ZN(n4461) );
  NAND2_X1 U6046 ( .A1(n6710), .A2(n9732), .ZN(n6085) );
  OR2_X1 U6047 ( .A1(n4429), .A2(n4930), .ZN(n4462) );
  AND2_X1 U6048 ( .A1(n4761), .A2(n4760), .ZN(n4463) );
  AND2_X1 U6049 ( .A1(n4809), .A2(n4517), .ZN(n4464) );
  NOR2_X1 U6050 ( .A1(n8389), .A2(n8414), .ZN(n4465) );
  NOR2_X1 U6051 ( .A1(n8471), .A2(n8274), .ZN(n4466) );
  INV_X1 U6052 ( .A(n6086), .ZN(n6087) );
  NAND2_X1 U6053 ( .A1(n6245), .A2(n6244), .ZN(n9289) );
  INV_X1 U6054 ( .A(n9289), .ZN(n4702) );
  OR2_X1 U6055 ( .A1(n9215), .A2(n9034), .ZN(n8949) );
  AND2_X1 U6056 ( .A1(n9248), .A2(n9467), .ZN(n4467) );
  OR2_X1 U6057 ( .A1(n5663), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4468) );
  OR2_X1 U6058 ( .A1(n7824), .A2(n8758), .ZN(n8894) );
  INV_X1 U6059 ( .A(n5120), .ZN(n5203) );
  AND2_X1 U6060 ( .A1(n6277), .A2(n6276), .ZN(n9467) );
  INV_X1 U6061 ( .A(n9467), .ZN(n4695) );
  OAI22_X1 U6062 ( .A1(n8771), .A2(n5106), .B1(n5782), .B2(n7847), .ZN(n8556)
         );
  OR2_X1 U6063 ( .A1(n7954), .A2(n7953), .ZN(n4469) );
  NAND2_X1 U6064 ( .A1(n6319), .A2(n6318), .ZN(n9370) );
  INV_X1 U6065 ( .A(n9370), .ZN(n4705) );
  AND2_X1 U6066 ( .A1(n9038), .A2(n8944), .ZN(n4470) );
  NAND2_X1 U6067 ( .A1(n4875), .A2(n7641), .ZN(n7652) );
  OR2_X1 U6068 ( .A1(n7392), .A2(n7533), .ZN(n8869) );
  OR2_X1 U6069 ( .A1(n9920), .A2(n7757), .ZN(n5932) );
  INV_X1 U6070 ( .A(n5932), .ZN(n4751) );
  AND2_X1 U6071 ( .A1(n7770), .A2(n8803), .ZN(n4471) );
  NOR2_X1 U6072 ( .A1(n8030), .A2(n8031), .ZN(n4472) );
  NOR2_X1 U6073 ( .A1(n4798), .A2(n8082), .ZN(n4797) );
  NAND2_X1 U6074 ( .A1(n6328), .A2(n6327), .ZN(n8006) );
  NAND2_X1 U6075 ( .A1(n7793), .A2(n7797), .ZN(n4473) );
  AND2_X1 U6076 ( .A1(n4747), .A2(n4748), .ZN(n4474) );
  INV_X1 U6077 ( .A(n6297), .ZN(n4930) );
  OR2_X1 U6078 ( .A1(n9199), .A2(n9388), .ZN(n6297) );
  INV_X1 U6079 ( .A(n8894), .ZN(n4523) );
  NOR2_X1 U6080 ( .A1(n7994), .A2(n7993), .ZN(n4475) );
  NOR2_X1 U6081 ( .A1(n9467), .A2(n9247), .ZN(n4476) );
  AND2_X1 U6082 ( .A1(n7960), .A2(n7959), .ZN(n4477) );
  AOI21_X1 U6083 ( .B1(n8776), .B2(n5764), .A(n5763), .ZN(n9508) );
  OR2_X1 U6084 ( .A1(n9452), .A2(n8751), .ZN(n4478) );
  NOR2_X1 U6085 ( .A1(n8135), .A2(n4673), .ZN(n4672) );
  AND2_X1 U6086 ( .A1(n4782), .A2(n8149), .ZN(n4479) );
  INV_X1 U6087 ( .A(n5043), .ZN(n5413) );
  NAND2_X1 U6088 ( .A1(n7006), .A2(n7009), .ZN(n7260) );
  NAND2_X1 U6089 ( .A1(n6388), .A2(n6387), .ZN(n6409) );
  NAND2_X1 U6090 ( .A1(n6892), .A2(n6126), .ZN(n7023) );
  AND2_X1 U6091 ( .A1(n7501), .A2(n5796), .ZN(n7491) );
  NAND2_X1 U6092 ( .A1(n6030), .A2(n6029), .ZN(n9539) );
  INV_X1 U6093 ( .A(n9539), .ZN(n4698) );
  NAND2_X1 U6094 ( .A1(n5437), .A2(n5436), .ZN(n8622) );
  INV_X1 U6095 ( .A(n8622), .ZN(n4989) );
  OR2_X1 U6096 ( .A1(n7934), .A2(n7933), .ZN(n4480) );
  INV_X1 U6097 ( .A(n8715), .ZN(n4849) );
  NAND2_X1 U6098 ( .A1(n9769), .A2(n7027), .ZN(n8974) );
  INV_X1 U6099 ( .A(n8974), .ZN(n4596) );
  OR2_X1 U6100 ( .A1(n4661), .A2(n7513), .ZN(n4481) );
  INV_X1 U6101 ( .A(n7132), .ZN(n4836) );
  NAND2_X1 U6102 ( .A1(n5603), .A2(n5602), .ZN(n8581) );
  INV_X1 U6103 ( .A(n8581), .ZN(n4655) );
  OR2_X1 U6104 ( .A1(n8496), .A2(n4727), .ZN(n4482) );
  NAND2_X1 U6105 ( .A1(n4876), .A2(n7522), .ZN(n7527) );
  INV_X1 U6106 ( .A(n4895), .ZN(n4894) );
  NOR2_X1 U6107 ( .A1(n5757), .A2(n5760), .ZN(n4895) );
  NOR2_X1 U6108 ( .A1(n5758), .A2(SI_29_), .ZN(n4483) );
  AND2_X1 U6109 ( .A1(n6944), .A2(n8977), .ZN(n4484) );
  AND2_X1 U6110 ( .A1(n9765), .A2(n6114), .ZN(n4485) );
  NAND2_X1 U6111 ( .A1(n6041), .A2(n6040), .ZN(n7618) );
  INV_X1 U6112 ( .A(n7618), .ZN(n4688) );
  INV_X1 U6113 ( .A(n8024), .ZN(n7409) );
  NOR2_X1 U6114 ( .A1(n6599), .A2(n6598), .ZN(n8744) );
  NAND2_X1 U6115 ( .A1(n5307), .A2(n5306), .ZN(n9920) );
  INV_X1 U6116 ( .A(n9920), .ZN(n4663) );
  NAND2_X1 U6117 ( .A1(n5416), .A2(n5415), .ZN(n8626) );
  INV_X1 U6118 ( .A(n8626), .ZN(n4650) );
  AND2_X1 U6119 ( .A1(n8955), .A2(n6371), .ZN(n9784) );
  AND2_X1 U6120 ( .A1(n6623), .A2(n6620), .ZN(n6757) );
  OAI211_X1 U6121 ( .C1(n6569), .C2(n6694), .A(n6568), .B(n6567), .ZN(n6603)
         );
  OR2_X1 U6122 ( .A1(n5776), .A2(SI_30_), .ZN(n4486) );
  INV_X1 U6123 ( .A(n6072), .ZN(n4922) );
  OR2_X1 U6124 ( .A1(n9137), .A2(n9136), .ZN(n4487) );
  INV_X1 U6125 ( .A(n7407), .ZN(n9034) );
  INV_X1 U6126 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4911) );
  INV_X1 U6127 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4760) );
  OAI222_X1 U6128 ( .A1(n8651), .A2(n6439), .B1(n8025), .B2(n6438), .C1(
        P2_U3152), .C2(n6811), .ZN(P2_U3353) );
  OAI222_X1 U6129 ( .A1(n8651), .A2(n6442), .B1(n8025), .B2(n6441), .C1(n8130), 
        .C2(n6813), .ZN(P2_U3352) );
  OAI222_X1 U6130 ( .A1(n8651), .A2(n6444), .B1(n8025), .B2(n6443), .C1(
        P2_U3152), .C2(n6806), .ZN(P2_U3354) );
  NAND2_X2 U6131 ( .A1(n6428), .A2(n8130), .ZN(n8651) );
  NAND2_X1 U6132 ( .A1(n5908), .A2(n5922), .ZN(n4540) );
  OAI222_X1 U6133 ( .A1(n8651), .A2(n8650), .B1(n8649), .B2(n8130), .C1(n8025), 
        .C2(n8648), .ZN(P2_U3331) );
  AOI21_X1 U6134 ( .B1(n4984), .B2(n4986), .A(n4466), .ZN(n4982) );
  AOI21_X1 U6135 ( .B1(n4968), .B2(n4971), .A(n4465), .ZN(n4966) );
  NOR2_X2 U6136 ( .A1(n4488), .A2(n4721), .ZN(n4991) );
  NAND2_X1 U6137 ( .A1(n9850), .A2(n9849), .ZN(n9852) );
  AOI21_X1 U6138 ( .B1(n4979), .B2(n4981), .A(n4978), .ZN(n4977) );
  MUX2_X1 U6139 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8632), .S(n9930), .Z(
        P2_U3517) );
  NAND2_X1 U6140 ( .A1(n8559), .A2(n9927), .ZN(n4586) );
  NAND2_X1 U6141 ( .A1(n8270), .A2(n8271), .ZN(n8525) );
  NAND2_X1 U6142 ( .A1(n7559), .A2(n4457), .ZN(n7706) );
  NAND2_X1 U6143 ( .A1(n6951), .A2(n4962), .ZN(n4961) );
  NAND2_X2 U6144 ( .A1(n6739), .A2(n6428), .ZN(n5782) );
  NAND2_X1 U6145 ( .A1(n7101), .A2(n7102), .ZN(n7100) );
  NAND2_X1 U6146 ( .A1(n5250), .A2(n5249), .ZN(n4800) );
  NAND2_X1 U6147 ( .A1(n5070), .A2(n7972), .ZN(n4789) );
  NAND2_X1 U6148 ( .A1(n5493), .A2(n5492), .ZN(n8047) );
  OAI21_X1 U6149 ( .B1(n8012), .B2(n8013), .A(n4790), .ZN(n7867) );
  OAI22_X1 U6150 ( .A1(n8101), .A2(n8100), .B1(n5448), .B2(n5447), .ZN(n8129)
         );
  NOR2_X2 U6151 ( .A1(n6081), .A2(n6080), .ZN(n9060) );
  NAND2_X2 U6152 ( .A1(n8663), .A2(n7921), .ZN(n7924) );
  OAI21_X2 U6153 ( .B1(n8653), .B2(n7942), .A(n8654), .ZN(n7943) );
  NAND2_X1 U6154 ( .A1(n4491), .A2(n4622), .ZN(n8724) );
  OAI21_X1 U6155 ( .B1(n4490), .B2(n4489), .A(n4492), .ZN(P1_U3238) );
  NAND2_X1 U6156 ( .A1(n8745), .A2(n8744), .ZN(n4490) );
  NAND2_X1 U6157 ( .A1(n7521), .A2(n7520), .ZN(n4876) );
  OAI21_X1 U6158 ( .B1(n8735), .B2(n5007), .A(n8733), .ZN(n4621) );
  NAND2_X1 U6159 ( .A1(n8714), .A2(n4845), .ZN(n4491) );
  AND2_X2 U6160 ( .A1(n6119), .A2(n6010), .ZN(n6012) );
  NAND2_X1 U6161 ( .A1(n6012), .A2(n6011), .ZN(n6140) );
  NAND2_X1 U6162 ( .A1(n7924), .A2(n7923), .ZN(n8714) );
  NAND2_X1 U6163 ( .A1(n4840), .A2(n4846), .ZN(n8723) );
  INV_X1 U6164 ( .A(n6012), .ZN(n6122) );
  NAND2_X1 U6165 ( .A1(n5724), .A2(n7498), .ZN(n7505) );
  NAND2_X4 U6166 ( .A1(n8649), .A2(n5705), .ZN(n6739) );
  INV_X1 U6167 ( .A(n4493), .ZN(n5673) );
  NAND2_X1 U6168 ( .A1(n4724), .A2(n5876), .ZN(n8426) );
  NAND2_X1 U6169 ( .A1(n4586), .A2(n4459), .ZN(n8632) );
  NAND2_X1 U6170 ( .A1(n8291), .A2(n8290), .ZN(n8563) );
  NAND2_X1 U6171 ( .A1(n4766), .A2(n5842), .ZN(n9841) );
  NAND2_X1 U6172 ( .A1(n5736), .A2(n5735), .ZN(n8309) );
  NAND2_X1 U6173 ( .A1(n4732), .A2(n4729), .ZN(n8472) );
  NAND2_X2 U6174 ( .A1(n8705), .A2(n7947), .ZN(n8682) );
  NAND2_X1 U6175 ( .A1(n4876), .A2(n4458), .ZN(n7580) );
  NAND2_X1 U6176 ( .A1(n4875), .A2(n4873), .ZN(n7813) );
  NAND2_X1 U6177 ( .A1(n6594), .A2(n6593), .ZN(n7857) );
  AND2_X2 U6178 ( .A1(n7813), .A2(n7812), .ZN(n7817) );
  NAND2_X1 U6179 ( .A1(n6583), .A2(n6582), .ZN(n6584) );
  INV_X1 U6180 ( .A(n4944), .ZN(n4943) );
  OAI21_X2 U6181 ( .B1(n7476), .B2(n4948), .A(n4946), .ZN(n4951) );
  AOI22_X2 U6182 ( .A1(n9256), .A2(n6265), .B1(n9284), .B2(n9474), .ZN(n9240)
         );
  OAI21_X2 U6183 ( .B1(n8698), .B2(n8697), .A(n4855), .ZN(n8735) );
  NAND2_X1 U6184 ( .A1(n8120), .A2(n5557), .ZN(n8041) );
  NAND2_X1 U6185 ( .A1(n4495), .A2(n6096), .ZN(n6776) );
  NAND3_X1 U6186 ( .A1(n4921), .A2(n4919), .A3(n6709), .ZN(n4495) );
  NAND2_X2 U6187 ( .A1(n6112), .A2(n6113), .ZN(n9765) );
  NAND2_X1 U6188 ( .A1(n4807), .A2(n4806), .ZN(n4805) );
  INV_X1 U6189 ( .A(n4920), .ZN(n6084) );
  NAND2_X1 U6190 ( .A1(n6083), .A2(n6085), .ZN(n4920) );
  NAND2_X1 U6191 ( .A1(n6577), .A2(n6578), .ZN(n6579) );
  NAND2_X1 U6192 ( .A1(n6982), .A2(n6981), .ZN(n4626) );
  AND2_X1 U6193 ( .A1(n6009), .A2(n4628), .ZN(n4627) );
  OR2_X1 U6194 ( .A1(n6569), .A2(n9732), .ZN(n6586) );
  NAND2_X1 U6195 ( .A1(n5043), .A2(n5000), .ZN(n5044) );
  NAND2_X1 U6196 ( .A1(n4789), .A2(n5077), .ZN(n8012) );
  NAND2_X1 U6197 ( .A1(n4674), .A2(n4795), .ZN(n8136) );
  NAND2_X2 U6198 ( .A1(n9836), .A2(n5279), .ZN(n7630) );
  NAND2_X1 U6199 ( .A1(n7295), .A2(n7239), .ZN(n7521) );
  NAND3_X1 U6200 ( .A1(n7293), .A2(n7294), .A3(n7297), .ZN(n7295) );
  INV_X1 U6201 ( .A(n4833), .ZN(n4623) );
  NAND2_X1 U6202 ( .A1(n7857), .A2(n6595), .ZN(n6760) );
  NAND2_X1 U6203 ( .A1(n4831), .A2(n4829), .ZN(n7228) );
  AND2_X2 U6204 ( .A1(n4627), .A2(n5984), .ZN(n5987) );
  NAND2_X1 U6205 ( .A1(n7376), .A2(n4504), .ZN(n4503) );
  OAI211_X1 U6206 ( .C1(n6370), .C2(n4508), .A(n4487), .B(n4507), .ZN(n9366)
         );
  NAND2_X1 U6207 ( .A1(n6370), .A2(n6338), .ZN(n9133) );
  NAND2_X1 U6208 ( .A1(n4514), .A2(n8861), .ZN(n7085) );
  NAND3_X1 U6209 ( .A1(n4816), .A2(n8981), .A3(n4515), .ZN(n4514) );
  NAND2_X1 U6210 ( .A1(n7686), .A2(n4518), .ZN(n4516) );
  NAND2_X1 U6211 ( .A1(n4516), .A2(n4464), .ZN(n6367) );
  OAI21_X1 U6212 ( .B1(n9258), .B2(n8913), .A(n8962), .ZN(n9243) );
  NAND2_X1 U6213 ( .A1(n8913), .A2(n8962), .ZN(n4531) );
  NAND2_X1 U6214 ( .A1(n4534), .A2(n5170), .ZN(n4533) );
  NAND2_X1 U6215 ( .A1(n5129), .A2(n5130), .ZN(n4667) );
  NOR2_X1 U6216 ( .A1(n4881), .A2(n4535), .ZN(n4534) );
  INV_X1 U6217 ( .A(n5169), .ZN(n4535) );
  NAND3_X1 U6218 ( .A1(n5904), .A2(n5903), .A3(n8353), .ZN(n4546) );
  NAND2_X1 U6219 ( .A1(n4547), .A2(n4548), .ZN(n5883) );
  NAND4_X1 U6220 ( .A1(n5861), .A2(n4551), .A3(n5860), .A4(n4549), .ZN(n4547)
         );
  AOI21_X1 U6221 ( .B1(n5883), .B2(n4550), .A(n5875), .ZN(n5877) );
  NAND3_X1 U6222 ( .A1(n5835), .A2(n5922), .A3(n5844), .ZN(n4552) );
  MUX2_X1 U6223 ( .A(n6427), .B(n6429), .S(n5061), .Z(n5131) );
  NAND3_X1 U6224 ( .A1(n4909), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4554) );
  NAND3_X1 U6225 ( .A1(n4911), .A2(n4912), .A3(n4910), .ZN(n4555) );
  NAND2_X1 U6226 ( .A1(n4557), .A2(n4455), .ZN(n4562) );
  NAND2_X1 U6227 ( .A1(n5324), .A2(n5323), .ZN(n5348) );
  INV_X1 U6228 ( .A(n5323), .ZN(n4560) );
  NAND2_X1 U6229 ( .A1(n4404), .A2(n5002), .ZN(n4563) );
  NAND2_X1 U6230 ( .A1(n5432), .A2(n4576), .ZN(n4575) );
  NAND2_X1 U6231 ( .A1(n5432), .A2(n4583), .ZN(n4582) );
  NAND2_X1 U6232 ( .A1(n5432), .A2(n5431), .ZN(n5454) );
  MUX2_X1 U6233 ( .A(n10262), .B(n6444), .S(n5061), .Z(n5152) );
  NAND2_X1 U6234 ( .A1(n4588), .A2(n8949), .ZN(n4587) );
  NAND2_X1 U6235 ( .A1(n4589), .A2(n8871), .ZN(n4588) );
  NAND2_X1 U6236 ( .A1(n8870), .A2(n4590), .ZN(n4589) );
  AND2_X1 U6237 ( .A1(n8869), .A2(n8868), .ZN(n4590) );
  NAND3_X1 U6238 ( .A1(n4594), .A2(n8864), .A3(n8865), .ZN(n4593) );
  AND2_X1 U6239 ( .A1(n4884), .A2(n4424), .ZN(n4616) );
  OAI211_X1 U6240 ( .C1(n4887), .C2(n4617), .A(n4883), .B(n4615), .ZN(n9037)
         );
  NAND2_X1 U6241 ( .A1(n4887), .A2(n4616), .ZN(n4615) );
  INV_X2 U6242 ( .A(n6896), .ZN(n9768) );
  AND2_X2 U6243 ( .A1(n4621), .A2(n4620), .ZN(n8663) );
  AND2_X2 U6244 ( .A1(n8724), .A2(n7939), .ZN(n8653) );
  NAND2_X1 U6245 ( .A1(n4626), .A2(n6983), .ZN(n7120) );
  AOI21_X1 U6246 ( .B1(n4626), .B2(n4624), .A(n4623), .ZN(n7183) );
  NAND2_X1 U6247 ( .A1(n5984), .A2(n6009), .ZN(n6353) );
  NAND2_X1 U6248 ( .A1(n8682), .A2(n4631), .ZN(n4630) );
  AND2_X1 U6249 ( .A1(n5987), .A2(n4638), .ZN(n6382) );
  NAND2_X1 U6250 ( .A1(n5987), .A2(n4639), .ZN(n6381) );
  AND2_X2 U6251 ( .A1(n4643), .A2(n4642), .ZN(n5082) );
  NAND3_X1 U6252 ( .A1(n4991), .A2(n5019), .A3(n5145), .ZN(n5663) );
  OAI21_X1 U6253 ( .B1(n8558), .B2(n9922), .A(n8557), .ZN(n8631) );
  NAND2_X1 U6254 ( .A1(n4648), .A2(n9508), .ZN(n4647) );
  INV_X1 U6255 ( .A(n4657), .ZN(n8358) );
  INV_X1 U6256 ( .A(n7513), .ZN(n4658) );
  NAND2_X1 U6257 ( .A1(n4658), .A2(n4659), .ZN(n7762) );
  INV_X1 U6258 ( .A(n5150), .ZN(n4666) );
  NAND2_X1 U6259 ( .A1(n8085), .A2(n4672), .ZN(n4669) );
  OR2_X2 U6260 ( .A1(n8085), .A2(n4797), .ZN(n4674) );
  NAND3_X1 U6261 ( .A1(n5387), .A2(n5388), .A3(n8151), .ZN(n4782) );
  NAND2_X1 U6262 ( .A1(n4677), .A2(n4454), .ZN(n5324) );
  MUX2_X1 U6263 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n5061), .Z(n5088) );
  MUX2_X1 U6264 ( .A(n6433), .B(n6431), .S(n5061), .Z(n5109) );
  INV_X1 U6265 ( .A(n4690), .ZN(n7552) );
  INV_X1 U6266 ( .A(n4696), .ZN(n9198) );
  MUX2_X1 U6267 ( .A(n7892), .B(P2_REG2_REG_1__SCAN_IN), .S(n6735), .Z(n8180)
         );
  NAND3_X1 U6268 ( .A1(n4723), .A2(n4722), .A3(n5010), .ZN(n4721) );
  OR2_X2 U6269 ( .A1(n8426), .A2(n8425), .ZN(n8408) );
  INV_X1 U6270 ( .A(n5720), .ZN(n4727) );
  NAND2_X1 U6271 ( .A1(n4727), .A2(n8175), .ZN(n5815) );
  NAND2_X1 U6272 ( .A1(n4727), .A2(n6956), .ZN(n6952) );
  NAND3_X1 U6273 ( .A1(n9876), .A2(n9875), .A3(n4725), .ZN(n9877) );
  NAND2_X1 U6274 ( .A1(n9886), .A2(n5720), .ZN(n4725) );
  OAI211_X1 U6275 ( .C1(n7328), .C2(n4727), .A(n9853), .B(n7327), .ZN(n9875)
         );
  OAI22_X1 U6276 ( .A1(n9832), .A2(n7868), .B1(n9829), .B2(n4727), .ZN(n7869)
         );
  NAND2_X1 U6277 ( .A1(n8529), .A2(n4733), .ZN(n4732) );
  NAND2_X1 U6278 ( .A1(n4742), .A2(n4740), .ZN(n7360) );
  NAND2_X1 U6279 ( .A1(n4743), .A2(n7338), .ZN(n4742) );
  NAND2_X1 U6280 ( .A1(n7710), .A2(n4750), .ZN(n4747) );
  NAND2_X1 U6281 ( .A1(n7505), .A2(n4764), .ZN(n4766) );
  NOR2_X1 U6282 ( .A1(n8567), .A2(n9860), .ZN(n8312) );
  XNOR2_X1 U6283 ( .A(n8309), .B(n8308), .ZN(n4770) );
  NAND2_X1 U6284 ( .A1(n8459), .A2(n8460), .ZN(n8458) );
  NAND2_X1 U6285 ( .A1(n5733), .A2(n5906), .ZN(n8338) );
  NAND2_X1 U6286 ( .A1(n5734), .A2(n5905), .ZN(n8326) );
  NAND2_X1 U6287 ( .A1(n7360), .A2(n7491), .ZN(n7503) );
  OAI21_X2 U6288 ( .B1(n9841), .B2(n5726), .A(n5942), .ZN(n7710) );
  NAND2_X1 U6289 ( .A1(n7324), .A2(n7325), .ZN(n7323) );
  MUX2_X1 U6290 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9495), .S(n6498), .Z(n9694) );
  NAND2_X1 U6291 ( .A1(n7100), .A2(n4774), .ZN(n4771) );
  NAND2_X1 U6292 ( .A1(n4771), .A2(n4772), .ZN(n7316) );
  NAND2_X1 U6293 ( .A1(n8092), .A2(n5428), .ZN(n8101) );
  NAND3_X1 U6294 ( .A1(n4782), .A2(n8093), .A3(n8149), .ZN(n8092) );
  NAND2_X1 U6295 ( .A1(n4783), .A2(n4784), .ZN(n5399) );
  NAND2_X1 U6296 ( .A1(n7630), .A2(n4426), .ZN(n4783) );
  NAND2_X1 U6297 ( .A1(n5119), .A2(n4456), .ZN(n7034) );
  AND2_X1 U6298 ( .A1(n5077), .A2(n5070), .ZN(n7973) );
  INV_X1 U6299 ( .A(n5096), .ZN(n4792) );
  NAND2_X1 U6300 ( .A1(n8047), .A2(n4793), .ZN(n5514) );
  INV_X1 U6301 ( .A(n8083), .ZN(n4798) );
  NAND2_X1 U6302 ( .A1(n4800), .A2(n4799), .ZN(n9836) );
  NAND2_X1 U6303 ( .A1(n5303), .A2(n4802), .ZN(n4801) );
  INV_X1 U6304 ( .A(n9732), .ZN(n7862) );
  NAND2_X1 U6305 ( .A1(n4812), .A2(n4453), .ZN(n6369) );
  OR2_X1 U6306 ( .A1(n9178), .A2(n4822), .ZN(n4819) );
  NAND2_X1 U6307 ( .A1(n4819), .A2(n4820), .ZN(n6370) );
  NAND2_X1 U6308 ( .A1(n7120), .A2(n4833), .ZN(n4831) );
  NOR2_X1 U6309 ( .A1(n7748), .A2(n7600), .ZN(n6389) );
  OR2_X1 U6310 ( .A1(n6382), .A2(n6121), .ZN(n4837) );
  NAND2_X1 U6311 ( .A1(n6381), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4839) );
  NAND2_X1 U6312 ( .A1(n7924), .A2(n4841), .ZN(n4840) );
  CLKBUF_X1 U6313 ( .A(n8714), .Z(n4843) );
  OAI21_X2 U6314 ( .B1(n7817), .B2(n4860), .A(n4856), .ZN(n8753) );
  NAND2_X1 U6315 ( .A1(n8745), .A2(n4864), .ZN(n4863) );
  OAI211_X1 U6316 ( .C1(n8745), .C2(n4865), .A(n7970), .B(n4863), .ZN(P1_U3212) );
  NAND2_X1 U6317 ( .A1(n7965), .A2(n4477), .ZN(n4869) );
  NAND2_X1 U6318 ( .A1(n8653), .A2(n7942), .ZN(n4871) );
  CLKBUF_X1 U6319 ( .A(n6981), .Z(n4877) );
  NAND2_X1 U6320 ( .A1(n8779), .A2(n8833), .ZN(n4878) );
  NAND2_X1 U6321 ( .A1(n4878), .A2(n9110), .ZN(n9019) );
  NAND2_X1 U6322 ( .A1(n5759), .A2(n4893), .ZN(n4890) );
  OAI21_X1 U6323 ( .B1(n5759), .B2(n4483), .A(n4894), .ZN(n5778) );
  NAND2_X1 U6324 ( .A1(n4890), .A2(n4425), .ZN(n5781) );
  NAND3_X1 U6325 ( .A1(n4894), .A2(n4483), .A3(n4892), .ZN(n4891) );
  NAND2_X1 U6326 ( .A1(n5633), .A2(n5632), .ZN(n5738) );
  NAND2_X1 U6327 ( .A1(n5633), .A2(n4897), .ZN(n4896) );
  INV_X2 U6328 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4909) );
  INV_X1 U6329 ( .A(n5061), .ZN(n5060) );
  NAND2_X1 U6330 ( .A1(n6072), .A2(n6085), .ZN(n4921) );
  NAND2_X1 U6331 ( .A1(n6993), .A2(n6085), .ZN(n6708) );
  NAND2_X1 U6332 ( .A1(n4922), .A2(n6084), .ZN(n6993) );
  NAND2_X1 U6333 ( .A1(n9240), .A2(n4933), .ZN(n4932) );
  NAND2_X1 U6334 ( .A1(n6151), .A2(n4940), .ZN(n4938) );
  OAI21_X1 U6335 ( .B1(n4431), .B2(n4945), .A(n7024), .ZN(n4944) );
  NAND2_X1 U6336 ( .A1(n7475), .A2(n6189), .ZN(n7463) );
  INV_X1 U6337 ( .A(n6189), .ZN(n4950) );
  NAND2_X1 U6338 ( .A1(n5987), .A2(n4956), .ZN(n6000) );
  NAND2_X1 U6339 ( .A1(n5987), .A2(n5004), .ZN(n6004) );
  NAND2_X1 U6340 ( .A1(n6675), .A2(n6667), .ZN(n6669) );
  OAI211_X2 U6341 ( .C1(n6739), .C2(n6735), .A(n5065), .B(n5064), .ZN(n7890)
         );
  NAND3_X1 U6342 ( .A1(n4961), .A2(n6954), .A3(n4960), .ZN(n7005) );
  NAND2_X1 U6343 ( .A1(n8420), .A2(n4968), .ZN(n4965) );
  NAND2_X1 U6344 ( .A1(n7260), .A2(n4979), .ZN(n4976) );
  NAND2_X1 U6345 ( .A1(n4976), .A2(n4977), .ZN(n7359) );
  NAND2_X1 U6346 ( .A1(n8507), .A2(n4984), .ZN(n4983) );
  NOR2_X2 U6347 ( .A1(n9249), .A2(n9263), .ZN(n9248) );
  NAND2_X1 U6348 ( .A1(n5430), .A2(n5429), .ZN(n5432) );
  CLKBUF_X1 U6349 ( .A(n7637), .Z(n7586) );
  OR2_X1 U6350 ( .A1(n6261), .A2(n6054), .ZN(n6057) );
  CLKBUF_X1 U6351 ( .A(n6760), .Z(n6596) );
  INV_X1 U6352 ( .A(n6004), .ZN(n6386) );
  OR2_X1 U6353 ( .A1(n7796), .A2(n7790), .ZN(n7750) );
  NAND2_X1 U6354 ( .A1(n6575), .A2(n6604), .ZN(n6628) );
  AOI21_X1 U6355 ( .B1(n8611), .B2(n8477), .A(n8451), .ZN(n8276) );
  OAI22_X1 U6356 ( .A1(n8365), .A2(n8373), .B1(n8584), .B2(n8395), .ZN(n8351)
         );
  INV_X1 U6357 ( .A(n6101), .ZN(n6086) );
  NAND2_X2 U6358 ( .A1(n7265), .A2(n8344), .ZN(n8549) );
  AND2_X1 U6359 ( .A1(n5159), .A2(n5158), .ZN(n4992) );
  AND3_X1 U6360 ( .A1(n6343), .A2(n6342), .A3(n6341), .ZN(n4993) );
  INV_X1 U6361 ( .A(n8488), .ZN(n9843) );
  INV_X1 U6362 ( .A(n9039), .ZN(n9362) );
  OR2_X1 U6363 ( .A1(n4706), .A2(n9439), .ZN(n4997) );
  OR2_X1 U6364 ( .A1(n4706), .A2(n9483), .ZN(n4998) );
  AND3_X1 U6365 ( .A1(n8065), .A2(n8067), .A3(n8138), .ZN(n4999) );
  AND4_X1 U6366 ( .A1(n5042), .A2(n5041), .A3(n10255), .A4(n5040), .ZN(n5000)
         );
  AND2_X1 U6367 ( .A1(n5281), .A2(n5260), .ZN(n5001) );
  AND2_X1 U6368 ( .A1(n5255), .A2(n5232), .ZN(n5002) );
  OR2_X1 U6369 ( .A1(n8288), .A2(n8287), .ZN(n5003) );
  INV_X1 U6370 ( .A(n9161), .ZN(n9197) );
  AND4_X1 U6371 ( .A1(n5986), .A2(n5985), .A3(n6391), .A4(n6383), .ZN(n5004)
         );
  INV_X1 U6372 ( .A(n7377), .ZN(n6175) );
  NAND2_X2 U6373 ( .A1(n6779), .A2(n9301), .ZN(n9716) );
  XNOR2_X1 U6374 ( .A(n7986), .B(n7915), .ZN(n5007) );
  INV_X1 U6375 ( .A(n6134), .ZN(n6153) );
  INV_X1 U6376 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5985) );
  INV_X1 U6377 ( .A(n8425), .ZN(n5730) );
  INV_X1 U6378 ( .A(n5505), .ZN(n5504) );
  INV_X1 U6379 ( .A(n6954), .ZN(n5721) );
  INV_X1 U6380 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n10260) );
  INV_X1 U6381 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5256) );
  INV_X1 U6382 ( .A(n5549), .ZN(n5547) );
  INV_X1 U6383 ( .A(n7491), .ZN(n7492) );
  INV_X1 U6384 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5041) );
  INV_X1 U6385 ( .A(n5532), .ZN(n5534) );
  INV_X1 U6386 ( .A(n5467), .ZN(n5468) );
  INV_X1 U6387 ( .A(SI_12_), .ZN(n5299) );
  INV_X1 U6388 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6011) );
  OR2_X1 U6389 ( .A1(n5389), .A2(n8152), .ZN(n5419) );
  INV_X1 U6390 ( .A(n7036), .ZN(n5138) );
  OR2_X1 U6391 ( .A1(n5311), .A2(n5310), .ZN(n5353) );
  OR2_X1 U6392 ( .A1(n5697), .A2(n8060), .ZN(n5752) );
  OR2_X1 U6393 ( .A1(n5569), .A2(n8042), .ZN(n5582) );
  NAND2_X1 U6394 ( .A1(n7493), .A2(n7492), .ZN(n7497) );
  OAI21_X1 U6395 ( .B1(n5680), .B2(P2_D_REG_1__SCAN_IN), .A(n5679), .ZN(n7261)
         );
  INV_X1 U6396 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6127) );
  INV_X1 U6397 ( .A(n8744), .ZN(n7995) );
  INV_X1 U6398 ( .A(n7958), .ZN(n7959) );
  NAND2_X1 U6399 ( .A1(n8665), .A2(n7922), .ZN(n7923) );
  INV_X1 U6400 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6181) );
  AND2_X1 U6401 ( .A1(n6220), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6222) );
  OR2_X1 U6402 ( .A1(n6330), .A2(n6329), .ZN(n6373) );
  NAND2_X1 U6403 ( .A1(n6269), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6279) );
  NOR2_X1 U6404 ( .A1(n6209), .A2(n10232), .ZN(n6220) );
  INV_X1 U6405 ( .A(n9160), .ZN(n7875) );
  INV_X1 U6406 ( .A(n8841), .ZN(n8957) );
  INV_X1 U6407 ( .A(n9260), .ZN(n7932) );
  OR2_X1 U6408 ( .A1(n8768), .A2(n9540), .ZN(n6227) );
  AND2_X1 U6409 ( .A1(n7645), .A2(n9040), .ZN(n6202) );
  OR2_X1 U6410 ( .A1(n5355), .A2(n5340), .ZN(n5389) );
  INV_X1 U6411 ( .A(n9827), .ZN(n5278) );
  OR2_X1 U6412 ( .A1(n5481), .A2(n5480), .ZN(n5505) );
  AND2_X1 U6413 ( .A1(n5969), .A2(n6727), .ZN(n7977) );
  AOI21_X1 U6414 ( .B1(n5161), .B2(n5160), .A(n4992), .ZN(n7101) );
  AND2_X1 U6415 ( .A1(n9921), .A2(n6526), .ZN(n5690) );
  NAND2_X1 U6416 ( .A1(n9922), .A2(n6674), .ZN(n5785) );
  OR2_X1 U6417 ( .A1(n8321), .A2(n5645), .ZN(n5650) );
  INV_X1 U6418 ( .A(n6727), .ZN(n6526) );
  AND2_X1 U6419 ( .A1(n5689), .A2(n5804), .ZN(n6727) );
  OR2_X1 U6420 ( .A1(n9862), .A2(n7264), .ZN(n8344) );
  INV_X1 U6421 ( .A(n9921), .ZN(n9886) );
  AND2_X1 U6422 ( .A1(n6674), .A2(n6673), .ZN(n8488) );
  OR3_X1 U6423 ( .A1(n7598), .A2(n7682), .A3(n7702), .ZN(n6425) );
  NOR2_X1 U6424 ( .A1(n6128), .A2(n6127), .ZN(n6144) );
  NOR2_X1 U6425 ( .A1(n7996), .A2(n7995), .ZN(n7997) );
  NAND2_X1 U6426 ( .A1(n7183), .A2(n4830), .ZN(n7293) );
  INV_X1 U6427 ( .A(n8762), .ZN(n8737) );
  OR2_X1 U6428 ( .A1(n6552), .A2(n9485), .ZN(n6599) );
  AND3_X1 U6429 ( .A1(n6465), .A2(n6464), .A3(n6463), .ZN(n9113) );
  AND2_X1 U6430 ( .A1(n6246), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6257) );
  INV_X1 U6431 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7252) );
  AND2_X1 U6432 ( .A1(n7407), .A2(n8954), .ZN(n6698) );
  INV_X1 U6433 ( .A(n8998), .ZN(n6338) );
  INV_X1 U6434 ( .A(n9228), .ZN(n9196) );
  INV_X1 U6435 ( .A(n9431), .ZN(n9316) );
  INV_X1 U6436 ( .A(n9432), .ZN(n8758) );
  AND2_X1 U6437 ( .A1(n8879), .A2(n8873), .ZN(n8965) );
  INV_X1 U6438 ( .A(n9695), .ZN(n9319) );
  AND2_X1 U6439 ( .A1(n9695), .A2(n9704), .ZN(n6554) );
  INV_X1 U6440 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n10232) );
  NAND2_X1 U6441 ( .A1(n8773), .A2(n8780), .ZN(n8775) );
  NAND2_X1 U6442 ( .A1(n9028), .A2(n6698), .ZN(n9782) );
  AND2_X1 U6443 ( .A1(n9719), .A2(n6545), .ZN(n6690) );
  AND2_X1 U6444 ( .A1(n5632), .A2(n5612), .ZN(n5630) );
  OAI21_X1 U6445 ( .B1(n8324), .B2(n9829), .A(n5712), .ZN(n5713) );
  NAND2_X1 U6446 ( .A1(n5264), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5311) );
  INV_X1 U6447 ( .A(n8533), .ZN(n8500) );
  AND2_X1 U6448 ( .A1(n7268), .A2(n5688), .ZN(n9921) );
  AND3_X1 U6449 ( .A1(n5767), .A2(n5766), .A3(n5765), .ZN(n7854) );
  AND4_X1 U6450 ( .A1(n5444), .A2(n5443), .A3(n5442), .A4(n5441), .ZN(n8501)
         );
  AND4_X1 U6451 ( .A1(n5289), .A2(n5288), .A3(n5287), .A4(n5286), .ZN(n9833)
         );
  INV_X1 U6452 ( .A(n6813), .ZN(n6862) );
  AND2_X1 U6453 ( .A1(n6741), .A2(n6740), .ZN(n8258) );
  INV_X1 U6454 ( .A(n9882), .ZN(n7349) );
  INV_X1 U6455 ( .A(n8344), .ZN(n9845) );
  NOR2_X1 U6456 ( .A1(n9864), .A2(n5678), .ZN(n7270) );
  INV_X1 U6457 ( .A(n9927), .ZN(n8624) );
  NAND2_X1 U6458 ( .A1(n8508), .A2(n9524), .ZN(n9927) );
  INV_X1 U6459 ( .A(n5680), .ZN(n9861) );
  NAND2_X1 U6460 ( .A1(n5006), .A2(n6595), .ZN(n7860) );
  INV_X1 U6461 ( .A(n8765), .ZN(n8749) );
  AND4_X1 U6462 ( .A1(n6284), .A2(n6283), .A3(n6282), .A4(n6281), .ZN(n9247)
         );
  INV_X1 U6463 ( .A(n6374), .ZN(n6264) );
  AND2_X1 U6464 ( .A1(n6500), .A2(n7744), .ZN(n9100) );
  INV_X1 U6465 ( .A(n9600), .ZN(n9687) );
  INV_X1 U6466 ( .A(n9686), .ZN(n9651) );
  AND2_X1 U6467 ( .A1(n9561), .A2(n9047), .ZN(n9686) );
  XNOR2_X1 U6468 ( .A(n9123), .B(n9134), .ZN(n9360) );
  AND2_X1 U6469 ( .A1(n8868), .A2(n8867), .ZN(n8983) );
  INV_X1 U6470 ( .A(n9333), .ZN(n9300) );
  INV_X1 U6471 ( .A(n9486), .ZN(n6691) );
  INV_X1 U6472 ( .A(n9784), .ZN(n9706) );
  INV_X1 U6473 ( .A(n9782), .ZN(n9795) );
  NAND2_X1 U6474 ( .A1(n9712), .A2(n9801), .ZN(n9789) );
  INV_X1 U6475 ( .A(n9485), .ZN(n9719) );
  AND2_X1 U6476 ( .A1(n6206), .A2(n6216), .ZN(n9677) );
  AND2_X1 U6477 ( .A1(n6166), .A2(n6177), .ZN(n6646) );
  INV_X1 U6478 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6051) );
  XNOR2_X1 U6479 ( .A(n5090), .B(n5063), .ZN(n5089) );
  INV_X1 U6480 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10107) );
  INV_X1 U6481 ( .A(n8262), .ZN(n8235) );
  NAND2_X1 U6482 ( .A1(n5709), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9840) );
  NAND2_X1 U6483 ( .A1(n8066), .A2(n4999), .ZN(n8071) );
  INV_X1 U6484 ( .A(n8062), .ZN(n8311) );
  NAND2_X1 U6485 ( .A1(n6724), .A2(n9868), .ZN(n8164) );
  INV_X1 U6486 ( .A(n7357), .ZN(n8171) );
  NAND2_X1 U6487 ( .A1(n8549), .A2(n7269), .ZN(n8496) );
  INV_X1 U6488 ( .A(n9945), .ZN(n9943) );
  INV_X1 U6489 ( .A(n9930), .ZN(n9928) );
  NOR2_X1 U6490 ( .A1(n9862), .A2(n9861), .ZN(n9863) );
  AND2_X1 U6491 ( .A1(n7598), .A2(n7702), .ZN(n9864) );
  XNOR2_X1 U6492 ( .A(n5670), .B(n5669), .ZN(n7598) );
  INV_X1 U6493 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6689) );
  NAND2_X1 U6494 ( .A1(n8010), .A2(n7998), .ZN(n8008) );
  AND2_X1 U6495 ( .A1(n6551), .A2(n6607), .ZN(n8765) );
  INV_X1 U6496 ( .A(n9247), .ZN(n9389) );
  INV_X1 U6497 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9507) );
  OR2_X1 U6498 ( .A1(P1_U3083), .A2(n6501), .ZN(n9691) );
  NAND2_X1 U6499 ( .A1(n9122), .A2(n6340), .ZN(n7884) );
  NAND3_X1 U6500 ( .A1(n9716), .A2(n6774), .A3(n7986), .ZN(n9333) );
  NAND2_X1 U6501 ( .A1(n10189), .A2(n9795), .ZN(n9439) );
  OR2_X1 U6502 ( .A1(n6419), .A2(n6691), .ZN(n10187) );
  INV_X1 U6503 ( .A(n9166), .ZN(n9452) );
  INV_X1 U6504 ( .A(n9265), .ZN(n9474) );
  NAND2_X1 U6505 ( .A1(n9809), .A2(n9795), .ZN(n9483) );
  OR2_X1 U6506 ( .A1(n6419), .A2(n9486), .ZN(n9807) );
  AND2_X1 U6507 ( .A1(n9719), .A2(n9718), .ZN(n9720) );
  NAND2_X1 U6508 ( .A1(n6558), .A2(n6393), .ZN(n9485) );
  INV_X1 U6509 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10219) );
  INV_X1 U6510 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10193) );
  INV_X1 U6511 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6461) );
  NOR2_X1 U6512 ( .A1(n10290), .A2(n10289), .ZN(n10288) );
  NOR2_X1 U6513 ( .A1(n9973), .A2(n9972), .ZN(n9971) );
  INV_X1 U6514 ( .A(n8164), .ZN(P2_U3966) );
  NAND2_X1 U6515 ( .A1(n6422), .A2(n4997), .ZN(P1_U3551) );
  NAND2_X1 U6516 ( .A1(n6418), .A2(n4998), .ZN(P1_U3519) );
  NOR2_X2 U6517 ( .A1(n5103), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5145) );
  NOR2_X1 U6518 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5014) );
  NOR2_X1 U6519 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5013) );
  NOR2_X1 U6520 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5012) );
  NOR2_X1 U6521 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5011) );
  NAND4_X1 U6522 ( .A1(n5014), .A2(n5013), .A3(n5012), .A4(n5011), .ZN(n5018)
         );
  NOR2_X1 U6523 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5016) );
  INV_X2 U6524 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n10255) );
  NAND4_X1 U6525 ( .A1(n5016), .A2(n5015), .A3(n10255), .A4(n5666), .ZN(n5017)
         );
  NOR2_X2 U6526 ( .A1(n5018), .A2(n5017), .ZN(n5019) );
  OAI21_X1 U6527 ( .B1(n5024), .B2(n5411), .A(P2_IR_REG_29__SCAN_IN), .ZN(
        n5027) );
  AND2_X4 U6528 ( .A1(n5030), .A2(n5031), .ZN(n5584) );
  NAND2_X1 U6529 ( .A1(n5584), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5035) );
  NAND2_X1 U6530 ( .A1(n5120), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5034) );
  NAND2_X1 U6531 ( .A1(n4406), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5033) );
  NAND3_X1 U6532 ( .A1(n5331), .A2(n5334), .A3(n5373), .ZN(n5036) );
  NAND2_X1 U6533 ( .A1(n5455), .A2(n5041), .ZN(n5038) );
  INV_X1 U6534 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5040) );
  NAND2_X1 U6535 ( .A1(n5044), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5045) );
  NAND2_X1 U6536 ( .A1(n7310), .A2(n5687), .ZN(n5361) );
  NOR2_X1 U6537 ( .A1(n8024), .A2(n6683), .ZN(n5066) );
  INV_X1 U6538 ( .A(n5046), .ZN(n5047) );
  NAND2_X1 U6539 ( .A1(n5047), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n5048) );
  NAND2_X1 U6540 ( .A1(n7310), .A2(n5804), .ZN(n7266) );
  NAND2_X4 U6541 ( .A1(n5051), .A2(n7266), .ZN(n5641) );
  INV_X1 U6542 ( .A(n5052), .ZN(n5055) );
  NAND2_X1 U6543 ( .A1(n5673), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5054) );
  NAND2_X2 U6544 ( .A1(n5056), .A2(n5055), .ZN(n8649) );
  INV_X1 U6545 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5058) );
  NAND2_X1 U6546 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5057) );
  AND2_X1 U6547 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5059) );
  NAND2_X1 U6548 ( .A1(n5060), .A2(n5059), .ZN(n6069) );
  NAND3_X1 U6549 ( .A1(n5061), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n5062) );
  NAND2_X1 U6550 ( .A1(n6069), .A2(n5062), .ZN(n5090) );
  INV_X1 U6551 ( .A(SI_1_), .ZN(n5063) );
  XNOR2_X1 U6552 ( .A(n5089), .B(n5088), .ZN(n6436) );
  OR2_X1 U6553 ( .A1(n5106), .A2(n6436), .ZN(n5065) );
  INV_X1 U6554 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6432) );
  OR2_X1 U6555 ( .A1(n5782), .A2(n6432), .ZN(n5064) );
  XNOR2_X1 U6556 ( .A(n5641), .B(n7890), .ZN(n5067) );
  NAND2_X1 U6557 ( .A1(n5066), .A2(n5067), .ZN(n5070) );
  INV_X1 U6558 ( .A(n5066), .ZN(n5069) );
  INV_X1 U6559 ( .A(n5067), .ZN(n5068) );
  NAND2_X1 U6560 ( .A1(n5069), .A2(n5068), .ZN(n5077) );
  NAND2_X1 U6561 ( .A1(n5584), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5074) );
  NAND2_X1 U6562 ( .A1(n4405), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5073) );
  NAND2_X1 U6563 ( .A1(n5120), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5072) );
  NAND2_X1 U6564 ( .A1(n4407), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5071) );
  NAND4_X1 U6565 ( .A1(n5074), .A2(n5073), .A3(n5072), .A4(n5071), .ZN(n5716)
         );
  NAND2_X1 U6566 ( .A1(n5061), .A2(SI_0_), .ZN(n5075) );
  XNOR2_X1 U6567 ( .A(n5075), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8652) );
  MUX2_X1 U6568 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8652), .S(n6739), .Z(n8020) );
  NAND2_X1 U6569 ( .A1(n5716), .A2(n8020), .ZN(n6668) );
  INV_X1 U6570 ( .A(n6668), .ZN(n6671) );
  NOR2_X1 U6571 ( .A1(n5641), .A2(n8020), .ZN(n5076) );
  NAND2_X1 U6572 ( .A1(n4430), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5081) );
  NAND2_X1 U6573 ( .A1(n5120), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5080) );
  NAND2_X1 U6574 ( .A1(n4408), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5079) );
  NAND2_X1 U6575 ( .A1(n5584), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5078) );
  AND4_X2 U6576 ( .A1(n5081), .A2(n5080), .A3(n5079), .A4(n5078), .ZN(n5717)
         );
  INV_X1 U6577 ( .A(n5361), .ZN(n6683) );
  OR2_X1 U6578 ( .A1(n5717), .A2(n6683), .ZN(n5095) );
  NOR2_X1 U6579 ( .A1(n5083), .A2(n5411), .ZN(n5084) );
  MUX2_X1 U6580 ( .A(n5411), .B(n5084), .S(P2_IR_REG_2__SCAN_IN), .Z(n5085) );
  INV_X1 U6581 ( .A(n5085), .ZN(n5087) );
  NAND2_X1 U6582 ( .A1(n5087), .A2(n5086), .ZN(n8192) );
  INV_X1 U6583 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6431) );
  OR2_X1 U6584 ( .A1(n5782), .A2(n6431), .ZN(n5094) );
  NAND2_X1 U6585 ( .A1(n5089), .A2(n5088), .ZN(n5092) );
  NAND2_X1 U6586 ( .A1(n5090), .A2(SI_1_), .ZN(n5091) );
  NAND2_X1 U6587 ( .A1(n5092), .A2(n5091), .ZN(n5108) );
  INV_X1 U6588 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6433) );
  XNOR2_X1 U6589 ( .A(n5109), .B(SI_2_), .ZN(n5107) );
  XNOR2_X1 U6590 ( .A(n5108), .B(n5107), .ZN(n6434) );
  INV_X1 U6591 ( .A(n8545), .ZN(n6949) );
  XNOR2_X1 U6592 ( .A(n5641), .B(n6949), .ZN(n5096) );
  XNOR2_X1 U6593 ( .A(n5095), .B(n5096), .ZN(n8013) );
  NAND2_X1 U6594 ( .A1(n5120), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5101) );
  NAND2_X1 U6595 ( .A1(n4430), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5100) );
  INV_X1 U6596 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5097) );
  NAND2_X1 U6597 ( .A1(n4408), .A2(n5097), .ZN(n5099) );
  NAND2_X1 U6598 ( .A1(n5584), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5098) );
  OR2_X1 U6599 ( .A1(n6956), .A2(n6683), .ZN(n5115) );
  NAND2_X1 U6600 ( .A1(n5086), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5102) );
  MUX2_X1 U6601 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5102), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5105) );
  NAND2_X1 U6602 ( .A1(n5105), .A2(n5104), .ZN(n6790) );
  INV_X1 U6603 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6429) );
  NAND2_X1 U6604 ( .A1(n5108), .A2(n5107), .ZN(n5112) );
  INV_X1 U6605 ( .A(n5109), .ZN(n5110) );
  NAND2_X1 U6606 ( .A1(n5110), .A2(SI_2_), .ZN(n5111) );
  NAND2_X1 U6607 ( .A1(n5112), .A2(n5111), .ZN(n5130) );
  INV_X1 U6608 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6427) );
  XNOR2_X1 U6609 ( .A(n5131), .B(SI_3_), .ZN(n5129) );
  XNOR2_X1 U6610 ( .A(n5130), .B(n5129), .ZN(n6430) );
  OR2_X1 U6611 ( .A1(n5106), .A2(n6430), .ZN(n5113) );
  OAI211_X1 U6612 ( .C1(n6739), .C2(n6790), .A(n5114), .B(n5113), .ZN(n5720)
         );
  XNOR2_X1 U6613 ( .A(n5641), .B(n5720), .ZN(n5116) );
  XNOR2_X1 U6614 ( .A(n5115), .B(n5116), .ZN(n7866) );
  NAND2_X1 U6615 ( .A1(n7867), .A2(n7866), .ZN(n5119) );
  INV_X1 U6616 ( .A(n5115), .ZN(n5117) );
  NAND2_X1 U6617 ( .A1(n5117), .A2(n5116), .ZN(n5118) );
  NAND2_X1 U6618 ( .A1(n5120), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5126) );
  NAND2_X1 U6619 ( .A1(n4430), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5125) );
  AND2_X1 U6620 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5140) );
  NOR2_X1 U6621 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5122) );
  NOR2_X1 U6622 ( .A1(n5140), .A2(n5122), .ZN(n7038) );
  NAND2_X1 U6623 ( .A1(n4408), .A2(n7038), .ZN(n5124) );
  NAND2_X1 U6624 ( .A1(n5584), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5123) );
  OR2_X1 U6625 ( .A1(n7868), .A2(n6683), .ZN(n5137) );
  NAND2_X1 U6626 ( .A1(n5104), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5128) );
  INV_X1 U6627 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5127) );
  XNOR2_X1 U6628 ( .A(n5128), .B(n5127), .ZN(n6806) );
  INV_X1 U6629 ( .A(n5131), .ZN(n5132) );
  NAND2_X1 U6630 ( .A1(n5132), .A2(SI_3_), .ZN(n5133) );
  XNOR2_X1 U6631 ( .A(n5152), .B(SI_4_), .ZN(n5150) );
  XNOR2_X1 U6632 ( .A(n5151), .B(n5150), .ZN(n6443) );
  OR2_X1 U6633 ( .A1(n5106), .A2(n6443), .ZN(n5135) );
  OR2_X1 U6634 ( .A1(n5782), .A2(n6444), .ZN(n5134) );
  OAI211_X1 U6635 ( .C1(n6739), .C2(n6806), .A(n5135), .B(n5134), .ZN(n7290)
         );
  XNOR2_X1 U6636 ( .A(n5641), .B(n4645), .ZN(n5136) );
  NAND2_X1 U6637 ( .A1(n5137), .A2(n5136), .ZN(n5139) );
  OAI21_X1 U6638 ( .B1(n5137), .B2(n5136), .A(n5139), .ZN(n7036) );
  INV_X1 U6639 ( .A(n6921), .ZN(n5161) );
  NAND2_X1 U6640 ( .A1(n5120), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5144) );
  NAND2_X1 U6641 ( .A1(n4430), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5143) );
  NAND2_X1 U6642 ( .A1(n5140), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5163) );
  OAI21_X1 U6643 ( .B1(n5140), .B2(P2_REG3_REG_5__SCAN_IN), .A(n5163), .ZN(
        n6925) );
  INV_X1 U6644 ( .A(n6925), .ZN(n7450) );
  NAND2_X1 U6645 ( .A1(n4408), .A2(n7450), .ZN(n5142) );
  NAND2_X1 U6646 ( .A1(n5584), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5141) );
  OR2_X1 U6647 ( .A1(n7258), .A2(n6683), .ZN(n5156) );
  NOR2_X1 U6648 ( .A1(n5146), .A2(n5411), .ZN(n5147) );
  MUX2_X1 U6649 ( .A(n5411), .B(n5147), .S(P2_IR_REG_5__SCAN_IN), .Z(n5149) );
  OR2_X1 U6650 ( .A1(n5149), .A2(n5148), .ZN(n6811) );
  INV_X1 U6651 ( .A(n5152), .ZN(n5153) );
  MUX2_X1 U6652 ( .A(n6439), .B(n6437), .S(n6428), .Z(n5171) );
  XNOR2_X1 U6653 ( .A(n5171), .B(SI_5_), .ZN(n5169) );
  OR2_X1 U6654 ( .A1(n5106), .A2(n6438), .ZN(n5155) );
  OR2_X1 U6655 ( .A1(n5782), .A2(n6439), .ZN(n5154) );
  OAI211_X1 U6656 ( .C1(n6739), .C2(n6811), .A(n5155), .B(n5154), .ZN(n7015)
         );
  INV_X1 U6657 ( .A(n7015), .ZN(n7449) );
  XNOR2_X1 U6658 ( .A(n5641), .B(n7449), .ZN(n5157) );
  XNOR2_X1 U6659 ( .A(n5156), .B(n5157), .ZN(n6920) );
  INV_X1 U6660 ( .A(n5156), .ZN(n5159) );
  INV_X1 U6661 ( .A(n5157), .ZN(n5158) );
  NAND2_X1 U6662 ( .A1(n5120), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5168) );
  INV_X1 U6663 ( .A(n4430), .ZN(n5268) );
  NAND2_X1 U6664 ( .A1(n4430), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5167) );
  INV_X1 U6665 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5162) );
  AND2_X1 U6666 ( .A1(n5163), .A2(n5162), .ZN(n5164) );
  NOR2_X1 U6667 ( .A1(n5187), .A2(n5164), .ZN(n7344) );
  NAND2_X1 U6668 ( .A1(n4408), .A2(n7344), .ZN(n5166) );
  NAND2_X1 U6669 ( .A1(n5584), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5165) );
  NOR2_X1 U6670 ( .A1(n7276), .A2(n9853), .ZN(n5181) );
  INV_X1 U6671 ( .A(n5171), .ZN(n5172) );
  NAND2_X1 U6672 ( .A1(n5172), .A2(SI_5_), .ZN(n5173) );
  MUX2_X1 U6673 ( .A(n6442), .B(n6440), .S(n6428), .Z(n5197) );
  XNOR2_X1 U6674 ( .A(n5197), .B(SI_6_), .ZN(n5195) );
  OR2_X1 U6675 ( .A1(n5106), .A2(n6441), .ZN(n5180) );
  OR2_X1 U6676 ( .A1(n5782), .A2(n6442), .ZN(n5179) );
  NOR2_X1 U6677 ( .A1(n5148), .A2(n5411), .ZN(n5174) );
  MUX2_X1 U6678 ( .A(n5411), .B(n5174), .S(P2_IR_REG_6__SCAN_IN), .Z(n5177) );
  INV_X1 U6679 ( .A(n5175), .ZN(n5176) );
  OR2_X1 U6680 ( .A1(n5177), .A2(n5176), .ZN(n6813) );
  NAND2_X1 U6681 ( .A1(n6524), .A2(n6862), .ZN(n5178) );
  XNOR2_X1 U6682 ( .A(n7349), .B(n5641), .ZN(n5182) );
  NAND2_X1 U6683 ( .A1(n5181), .A2(n5182), .ZN(n5185) );
  INV_X1 U6684 ( .A(n5181), .ZN(n5184) );
  INV_X1 U6685 ( .A(n5182), .ZN(n5183) );
  NAND2_X1 U6686 ( .A1(n5184), .A2(n5183), .ZN(n5186) );
  AND2_X1 U6687 ( .A1(n5185), .A2(n5186), .ZN(n7102) );
  NAND2_X1 U6688 ( .A1(n4430), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5193) );
  NAND2_X1 U6689 ( .A1(n5584), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5192) );
  NOR2_X1 U6690 ( .A1(n5187), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5188) );
  OR2_X1 U6691 ( .A1(n5242), .A2(n5188), .ZN(n7273) );
  INV_X1 U6692 ( .A(n7273), .ZN(n5189) );
  NAND2_X1 U6693 ( .A1(n4408), .A2(n5189), .ZN(n5191) );
  NAND2_X1 U6694 ( .A1(n5120), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5190) );
  INV_X2 U6695 ( .A(n9922), .ZN(n9853) );
  OR2_X1 U6696 ( .A1(n7357), .A2(n9853), .ZN(n5201) );
  NAND2_X1 U6697 ( .A1(n5175), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5194) );
  XNOR2_X1 U6698 ( .A(n5194), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6836) );
  INV_X1 U6699 ( .A(n6836), .ZN(n6448) );
  INV_X1 U6700 ( .A(n5197), .ZN(n5198) );
  MUX2_X1 U6701 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6428), .Z(n5212) );
  XNOR2_X1 U6702 ( .A(n5212), .B(SI_7_), .ZN(n5209) );
  XNOR2_X1 U6703 ( .A(n5211), .B(n5209), .ZN(n6446) );
  NAND2_X1 U6704 ( .A1(n6446), .A2(n5764), .ZN(n5200) );
  NAND2_X1 U6705 ( .A1(n5638), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n5199) );
  OAI211_X1 U6706 ( .C1(n6739), .C2(n6448), .A(n5200), .B(n5199), .ZN(n9885)
         );
  XNOR2_X1 U6707 ( .A(n5641), .B(n7356), .ZN(n5202) );
  XNOR2_X1 U6708 ( .A(n5201), .B(n5202), .ZN(n7109) );
  NAND2_X1 U6709 ( .A1(n5120), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5208) );
  NAND2_X1 U6710 ( .A1(n4430), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5207) );
  INV_X1 U6711 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5204) );
  XNOR2_X1 U6712 ( .A(n5242), .B(n5204), .ZN(n7171) );
  NAND2_X1 U6713 ( .A1(n5121), .A2(n7171), .ZN(n5206) );
  NAND2_X1 U6714 ( .A1(n5584), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5205) );
  OR2_X1 U6715 ( .A1(n7506), .A2(n6683), .ZN(n5223) );
  INV_X1 U6716 ( .A(n5209), .ZN(n5210) );
  NAND2_X1 U6717 ( .A1(n5211), .A2(n5210), .ZN(n5214) );
  NAND2_X1 U6718 ( .A1(n5212), .A2(SI_7_), .ZN(n5213) );
  MUX2_X1 U6719 ( .A(n5215), .B(n6453), .S(n6428), .Z(n5217) );
  INV_X1 U6720 ( .A(SI_8_), .ZN(n5216) );
  INV_X1 U6721 ( .A(n5217), .ZN(n5218) );
  NAND2_X1 U6722 ( .A1(n5218), .A2(SI_8_), .ZN(n5219) );
  XNOR2_X1 U6723 ( .A(n5227), .B(n5226), .ZN(n6451) );
  NAND2_X1 U6724 ( .A1(n6451), .A2(n5764), .ZN(n5222) );
  OR2_X1 U6725 ( .A1(n5175), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5233) );
  NAND2_X1 U6726 ( .A1(n5233), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5220) );
  XNOR2_X1 U6727 ( .A(n5220), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6873) );
  AOI22_X1 U6728 ( .A1(n5638), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6524), .B2(
        n6873), .ZN(n5221) );
  NAND2_X1 U6729 ( .A1(n5222), .A2(n5221), .ZN(n7494) );
  XNOR2_X1 U6730 ( .A(n7494), .B(n5641), .ZN(n5224) );
  XNOR2_X1 U6731 ( .A(n5223), .B(n5224), .ZN(n7169) );
  INV_X1 U6732 ( .A(n5223), .ZN(n5225) );
  INV_X1 U6733 ( .A(n7316), .ZN(n5250) );
  MUX2_X1 U6734 ( .A(n6456), .B(n6457), .S(n6428), .Z(n5230) );
  NAND2_X1 U6735 ( .A1(n5230), .A2(n5229), .ZN(n5255) );
  INV_X1 U6736 ( .A(n5230), .ZN(n5231) );
  NAND2_X1 U6737 ( .A1(n5231), .A2(SI_9_), .ZN(n5232) );
  NAND2_X1 U6738 ( .A1(n6455), .A2(n5764), .ZN(n5240) );
  NOR2_X1 U6739 ( .A1(n5233), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5236) );
  NOR2_X1 U6740 ( .A1(n5236), .A2(n5411), .ZN(n5234) );
  MUX2_X1 U6741 ( .A(n5411), .B(n5234), .S(P2_IR_REG_9__SCAN_IN), .Z(n5238) );
  INV_X1 U6742 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5235) );
  NAND2_X1 U6743 ( .A1(n5236), .A2(n5235), .ZN(n5282) );
  INV_X1 U6744 ( .A(n5282), .ZN(n5237) );
  INV_X1 U6745 ( .A(n6874), .ZN(n6890) );
  AOI22_X1 U6746 ( .A1(n5638), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6524), .B2(
        n6890), .ZN(n5239) );
  XNOR2_X1 U6747 ( .A(n9899), .B(n8055), .ZN(n5251) );
  NAND2_X1 U6748 ( .A1(n5120), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5248) );
  AND2_X1 U6749 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n5241) );
  AOI21_X1 U6750 ( .B1(n5242), .B2(P2_REG3_REG_8__SCAN_IN), .A(
        P2_REG3_REG_9__SCAN_IN), .ZN(n5243) );
  OR2_X1 U6751 ( .A1(n5264), .A2(n5243), .ZN(n7511) );
  INV_X1 U6752 ( .A(n7511), .ZN(n5244) );
  NAND2_X1 U6753 ( .A1(n5121), .A2(n5244), .ZN(n5247) );
  NAND2_X1 U6754 ( .A1(n5584), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5246) );
  NAND2_X1 U6755 ( .A1(n4430), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5245) );
  NAND4_X1 U6756 ( .A1(n5248), .A2(n5247), .A3(n5246), .A4(n5245), .ZN(n8169)
         );
  AND2_X1 U6757 ( .A1(n8169), .A2(n9922), .ZN(n5252) );
  AND2_X1 U6758 ( .A1(n5251), .A2(n5252), .ZN(n7313) );
  INV_X1 U6759 ( .A(n7313), .ZN(n5249) );
  INV_X1 U6760 ( .A(n5251), .ZN(n5254) );
  INV_X1 U6761 ( .A(n5252), .ZN(n5253) );
  NAND2_X1 U6762 ( .A1(n5254), .A2(n5253), .ZN(n7312) );
  MUX2_X1 U6763 ( .A(n5256), .B(n6461), .S(n6428), .Z(n5258) );
  INV_X1 U6764 ( .A(n5258), .ZN(n5259) );
  NAND2_X1 U6765 ( .A1(n5259), .A2(SI_10_), .ZN(n5260) );
  XNOR2_X1 U6766 ( .A(n5280), .B(n5001), .ZN(n6459) );
  NAND2_X1 U6767 ( .A1(n6459), .A2(n5764), .ZN(n5263) );
  NAND2_X1 U6768 ( .A1(n5282), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5261) );
  XNOR2_X1 U6769 ( .A(n5261), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7076) );
  AOI22_X1 U6770 ( .A1(n5638), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6524), .B2(
        n7076), .ZN(n5262) );
  XNOR2_X1 U6771 ( .A(n7704), .B(n5641), .ZN(n5273) );
  NAND2_X1 U6772 ( .A1(n5120), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5272) );
  INV_X1 U6773 ( .A(n5264), .ZN(n5265) );
  INV_X1 U6774 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10205) );
  NAND2_X1 U6775 ( .A1(n5265), .A2(n10205), .ZN(n5266) );
  NAND2_X1 U6776 ( .A1(n5311), .A2(n5266), .ZN(n9839) );
  INV_X1 U6777 ( .A(n9839), .ZN(n5267) );
  NAND2_X1 U6778 ( .A1(n5121), .A2(n5267), .ZN(n5271) );
  NAND2_X1 U6779 ( .A1(n5584), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5270) );
  INV_X1 U6780 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7567) );
  OR2_X1 U6781 ( .A1(n5268), .A2(n7567), .ZN(n5269) );
  NOR2_X1 U6782 ( .A1(n7703), .A2(n9853), .ZN(n5274) );
  NAND2_X1 U6783 ( .A1(n5273), .A2(n5274), .ZN(n5279) );
  INV_X1 U6784 ( .A(n5273), .ZN(n5276) );
  INV_X1 U6785 ( .A(n5274), .ZN(n5275) );
  NAND2_X1 U6786 ( .A1(n5276), .A2(n5275), .ZN(n5277) );
  NAND2_X1 U6787 ( .A1(n5279), .A2(n5277), .ZN(n9827) );
  MUX2_X1 U6788 ( .A(n6511), .B(n10261), .S(n6428), .Z(n5297) );
  XNOR2_X1 U6789 ( .A(n5296), .B(n5294), .ZN(n6509) );
  NAND2_X1 U6790 ( .A1(n6509), .A2(n5764), .ZN(n5285) );
  OAI21_X1 U6791 ( .B1(n5282), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5283) );
  XNOR2_X1 U6792 ( .A(n5283), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8206) );
  AOI22_X1 U6793 ( .A1(n5638), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6524), .B2(
        n8206), .ZN(n5284) );
  NAND2_X1 U6794 ( .A1(n5285), .A2(n5284), .ZN(n9848) );
  XNOR2_X1 U6795 ( .A(n9848), .B(n8055), .ZN(n5290) );
  NAND2_X1 U6796 ( .A1(n5120), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U6797 ( .A1(n4430), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5288) );
  XNOR2_X1 U6798 ( .A(n5311), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n9846) );
  NAND2_X1 U6799 ( .A1(n5121), .A2(n9846), .ZN(n5287) );
  NAND2_X1 U6800 ( .A1(n5584), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5286) );
  NOR2_X1 U6801 ( .A1(n9833), .A2(n9853), .ZN(n5291) );
  XNOR2_X1 U6802 ( .A(n5290), .B(n5291), .ZN(n7629) );
  INV_X1 U6803 ( .A(n5290), .ZN(n5292) );
  NAND2_X1 U6804 ( .A1(n5292), .A2(n5291), .ZN(n5293) );
  INV_X1 U6805 ( .A(n5297), .ZN(n5298) );
  MUX2_X1 U6806 ( .A(n10015), .B(n6532), .S(n6428), .Z(n5300) );
  INV_X1 U6807 ( .A(n5300), .ZN(n5301) );
  NAND2_X1 U6808 ( .A1(n5301), .A2(SI_12_), .ZN(n5302) );
  NAND2_X1 U6809 ( .A1(n5323), .A2(n5302), .ZN(n5321) );
  XNOR2_X1 U6810 ( .A(n5322), .B(n5321), .ZN(n6529) );
  NAND2_X1 U6811 ( .A1(n6529), .A2(n5764), .ZN(n5307) );
  INV_X1 U6812 ( .A(n5303), .ZN(n5304) );
  NAND2_X1 U6813 ( .A1(n5304), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5305) );
  XNOR2_X1 U6814 ( .A(n5305), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7147) );
  AOI22_X1 U6815 ( .A1(n5638), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6524), .B2(
        n7147), .ZN(n5306) );
  XNOR2_X1 U6816 ( .A(n9920), .B(n8055), .ZN(n5317) );
  NAND2_X1 U6817 ( .A1(n4430), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U6818 ( .A1(n5120), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5315) );
  INV_X1 U6819 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5309) );
  INV_X1 U6820 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5308) );
  OAI21_X1 U6821 ( .B1(n5311), .B2(n5309), .A(n5308), .ZN(n5312) );
  NAND2_X1 U6822 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n5310) );
  AND2_X1 U6823 ( .A1(n5312), .A2(n5353), .ZN(n7712) );
  NAND2_X1 U6824 ( .A1(n5121), .A2(n7712), .ZN(n5314) );
  NAND2_X1 U6825 ( .A1(n5584), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5313) );
  OR2_X1 U6826 ( .A1(n7757), .A2(n9853), .ZN(n5318) );
  NAND2_X1 U6827 ( .A1(n5317), .A2(n5318), .ZN(n7672) );
  INV_X1 U6828 ( .A(n5317), .ZN(n5320) );
  INV_X1 U6829 ( .A(n5318), .ZN(n5319) );
  NAND2_X1 U6830 ( .A1(n5320), .A2(n5319), .ZN(n7736) );
  MUX2_X1 U6831 ( .A(n6539), .B(n10193), .S(n6428), .Z(n5326) );
  INV_X1 U6832 ( .A(n5326), .ZN(n5327) );
  NAND2_X1 U6833 ( .A1(n5327), .A2(SI_13_), .ZN(n5328) );
  MUX2_X1 U6834 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6428), .Z(n5364) );
  XNOR2_X1 U6835 ( .A(n5366), .B(n5363), .ZN(n6542) );
  NAND2_X1 U6836 ( .A1(n6542), .A2(n5764), .ZN(n5338) );
  NAND2_X1 U6837 ( .A1(n5330), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U6838 ( .A1(n5349), .A2(n5331), .ZN(n5332) );
  NAND2_X1 U6839 ( .A1(n5332), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5335) );
  INV_X1 U6840 ( .A(n5335), .ZN(n5333) );
  NAND2_X1 U6841 ( .A1(n5333), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U6842 ( .A1(n5335), .A2(n5334), .ZN(n5372) );
  AOI22_X1 U6843 ( .A1(n5638), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6524), .B2(
        n8224), .ZN(n5337) );
  NAND2_X1 U6844 ( .A1(n5120), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U6845 ( .A1(n5339), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5355) );
  INV_X1 U6846 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U6847 ( .A1(n5355), .A2(n5340), .ZN(n5341) );
  AND2_X1 U6848 ( .A1(n5389), .A2(n5341), .ZN(n8034) );
  NAND2_X1 U6849 ( .A1(n5121), .A2(n8034), .ZN(n5345) );
  NAND2_X1 U6850 ( .A1(n5584), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5344) );
  INV_X1 U6851 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5342) );
  OR2_X1 U6852 ( .A1(n5268), .A2(n5342), .ZN(n5343) );
  INV_X1 U6853 ( .A(n8155), .ZN(n8531) );
  NAND2_X1 U6854 ( .A1(n8531), .A2(n9922), .ZN(n5383) );
  XNOR2_X1 U6855 ( .A(n5348), .B(n5347), .ZN(n6538) );
  NAND2_X1 U6856 ( .A1(n6538), .A2(n5764), .ZN(n5351) );
  XNOR2_X1 U6857 ( .A(n5349), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7611) );
  AOI22_X1 U6858 ( .A1(n5638), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6524), .B2(
        n7611), .ZN(n5350) );
  XNOR2_X1 U6859 ( .A(n9525), .B(n5641), .ZN(n5381) );
  NAND2_X1 U6860 ( .A1(n5584), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5360) );
  INV_X1 U6861 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U6862 ( .A1(n5353), .A2(n5352), .ZN(n5354) );
  AND2_X1 U6863 ( .A1(n5355), .A2(n5354), .ZN(n7764) );
  NAND2_X1 U6864 ( .A1(n5121), .A2(n7764), .ZN(n5359) );
  NAND2_X1 U6865 ( .A1(n5120), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5358) );
  INV_X1 U6866 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5356) );
  OR2_X1 U6867 ( .A1(n5268), .A2(n5356), .ZN(n5357) );
  INV_X1 U6868 ( .A(n8032), .ZN(n8165) );
  CLKBUF_X3 U6869 ( .A(n5361), .Z(n9922) );
  NAND2_X1 U6870 ( .A1(n8165), .A2(n9922), .ZN(n5380) );
  INV_X1 U6871 ( .A(n5380), .ZN(n5362) );
  NAND2_X1 U6872 ( .A1(n5381), .A2(n5362), .ZN(n8028) );
  AND2_X1 U6873 ( .A1(n7736), .A2(n5379), .ZN(n5395) );
  NAND2_X1 U6874 ( .A1(n5364), .A2(SI_14_), .ZN(n5365) );
  MUX2_X1 U6875 ( .A(n6689), .B(n5367), .S(n6428), .Z(n5369) );
  INV_X1 U6876 ( .A(SI_15_), .ZN(n5368) );
  NAND2_X1 U6877 ( .A1(n5369), .A2(n5368), .ZN(n5400) );
  INV_X1 U6878 ( .A(n5369), .ZN(n5370) );
  NAND2_X1 U6879 ( .A1(n5370), .A2(SI_15_), .ZN(n5371) );
  NAND2_X1 U6880 ( .A1(n5400), .A2(n5371), .ZN(n5401) );
  XNOR2_X1 U6881 ( .A(n5402), .B(n5401), .ZN(n6634) );
  NAND2_X1 U6882 ( .A1(n6634), .A2(n5764), .ZN(n5376) );
  NAND2_X1 U6883 ( .A1(n5372), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5374) );
  XNOR2_X1 U6884 ( .A(n5374), .B(n5373), .ZN(n7726) );
  INV_X1 U6885 ( .A(n7726), .ZN(n7605) );
  AOI22_X1 U6886 ( .A1(n5638), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6524), .B2(
        n7605), .ZN(n5375) );
  XNOR2_X1 U6887 ( .A(n8538), .B(n8055), .ZN(n5378) );
  AND2_X1 U6888 ( .A1(n5395), .A2(n5378), .ZN(n5377) );
  NAND2_X1 U6889 ( .A1(n7737), .A2(n5377), .ZN(n5388) );
  INV_X1 U6890 ( .A(n5378), .ZN(n5397) );
  INV_X1 U6891 ( .A(n5379), .ZN(n5382) );
  XNOR2_X1 U6892 ( .A(n5381), .B(n5380), .ZN(n8026) );
  OR2_X1 U6893 ( .A1(n5382), .A2(n8026), .ZN(n5386) );
  NAND2_X1 U6894 ( .A1(n5384), .A2(n5383), .ZN(n5385) );
  AND2_X1 U6895 ( .A1(n5386), .A2(n5385), .ZN(n5396) );
  NAND2_X1 U6896 ( .A1(n4430), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5394) );
  NAND2_X1 U6897 ( .A1(n5120), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5393) );
  INV_X1 U6898 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8152) );
  NAND2_X1 U6899 ( .A1(n5389), .A2(n8152), .ZN(n5390) );
  AND2_X1 U6900 ( .A1(n5419), .A2(n5390), .ZN(n8537) );
  NAND2_X1 U6901 ( .A1(n5121), .A2(n8537), .ZN(n5392) );
  NAND2_X1 U6902 ( .A1(n5584), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5391) );
  NOR2_X1 U6903 ( .A1(n8503), .A2(n9853), .ZN(n8151) );
  AND2_X1 U6904 ( .A1(n5397), .A2(n5396), .ZN(n5398) );
  NAND2_X1 U6905 ( .A1(n5399), .A2(n5398), .ZN(n8149) );
  MUX2_X1 U6906 ( .A(n5404), .B(n5403), .S(n6428), .Z(n5406) );
  INV_X1 U6907 ( .A(SI_16_), .ZN(n5405) );
  INV_X1 U6908 ( .A(n5406), .ZN(n5407) );
  NAND2_X1 U6909 ( .A1(n5407), .A2(SI_16_), .ZN(n5408) );
  XNOR2_X1 U6910 ( .A(n5430), .B(n5429), .ZN(n6659) );
  NAND2_X1 U6911 ( .A1(n6659), .A2(n5764), .ZN(n5416) );
  NOR2_X1 U6912 ( .A1(n5409), .A2(n5411), .ZN(n5410) );
  MUX2_X1 U6913 ( .A(n5411), .B(n5410), .S(P2_IR_REG_16__SCAN_IN), .Z(n5412)
         );
  INV_X1 U6914 ( .A(n5412), .ZN(n5414) );
  AND2_X1 U6915 ( .A1(n5414), .A2(n5413), .ZN(n7835) );
  AOI22_X1 U6916 ( .A1(n5638), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6524), .B2(
        n7835), .ZN(n5415) );
  XNOR2_X1 U6917 ( .A(n8626), .B(n8055), .ZN(n5427) );
  NAND2_X1 U6918 ( .A1(n4430), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U6919 ( .A1(n5120), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5423) );
  NAND2_X1 U6920 ( .A1(n5417), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5439) );
  INV_X1 U6921 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5418) );
  NAND2_X1 U6922 ( .A1(n5419), .A2(n5418), .ZN(n5420) );
  AND2_X1 U6923 ( .A1(n5439), .A2(n5420), .ZN(n8515) );
  NAND2_X1 U6924 ( .A1(n5121), .A2(n8515), .ZN(n5422) );
  NAND2_X1 U6925 ( .A1(n5584), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5421) );
  NOR2_X1 U6926 ( .A1(n8154), .A2(n9853), .ZN(n5425) );
  XNOR2_X1 U6927 ( .A(n5427), .B(n5425), .ZN(n8093) );
  INV_X1 U6928 ( .A(n5425), .ZN(n5426) );
  NAND2_X1 U6929 ( .A1(n5427), .A2(n5426), .ZN(n5428) );
  MUX2_X1 U6930 ( .A(n5434), .B(n5433), .S(n6428), .Z(n5450) );
  XNOR2_X1 U6931 ( .A(n5450), .B(SI_17_), .ZN(n5449) );
  XNOR2_X1 U6932 ( .A(n5454), .B(n5449), .ZN(n6720) );
  NAND2_X1 U6933 ( .A1(n6720), .A2(n5764), .ZN(n5437) );
  NAND2_X1 U6934 ( .A1(n5413), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5435) );
  XNOR2_X1 U6935 ( .A(n5435), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8238) );
  AOI22_X1 U6936 ( .A1(n5638), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6524), .B2(
        n8238), .ZN(n5436) );
  XNOR2_X1 U6937 ( .A(n8622), .B(n5641), .ZN(n5445) );
  NAND2_X1 U6938 ( .A1(n4430), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U6939 ( .A1(n5584), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5443) );
  INV_X1 U6940 ( .A(n5439), .ZN(n5438) );
  INV_X1 U6941 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8102) );
  NAND2_X1 U6942 ( .A1(n5439), .A2(n8102), .ZN(n5440) );
  AND2_X1 U6943 ( .A1(n5481), .A2(n5440), .ZN(n8493) );
  NAND2_X1 U6944 ( .A1(n5121), .A2(n8493), .ZN(n5442) );
  NAND2_X1 U6945 ( .A1(n5120), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5441) );
  NOR2_X1 U6946 ( .A1(n8501), .A2(n9853), .ZN(n5446) );
  XNOR2_X1 U6947 ( .A(n5445), .B(n5446), .ZN(n8100) );
  INV_X1 U6948 ( .A(n5445), .ZN(n5448) );
  INV_X1 U6949 ( .A(n5446), .ZN(n5447) );
  INV_X1 U6950 ( .A(n5449), .ZN(n5453) );
  INV_X1 U6951 ( .A(n5450), .ZN(n5451) );
  NAND2_X1 U6952 ( .A1(n5451), .A2(SI_17_), .ZN(n5452) );
  MUX2_X1 U6953 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6428), .Z(n5470) );
  XNOR2_X1 U6954 ( .A(n5470), .B(SI_18_), .ZN(n5467) );
  XNOR2_X1 U6955 ( .A(n5469), .B(n5467), .ZN(n6964) );
  NAND2_X1 U6956 ( .A1(n6964), .A2(n5764), .ZN(n5457) );
  XNOR2_X1 U6957 ( .A(n5455), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8250) );
  AOI22_X1 U6958 ( .A1(n5638), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6524), .B2(
        n8250), .ZN(n5456) );
  XNOR2_X1 U6959 ( .A(n5641), .B(n8615), .ZN(n5464) );
  NAND2_X1 U6960 ( .A1(n4430), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U6961 ( .A1(n5584), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5460) );
  XNOR2_X1 U6962 ( .A(n5481), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n8469) );
  NAND2_X1 U6963 ( .A1(n5121), .A2(n8469), .ZN(n5459) );
  NAND2_X1 U6964 ( .A1(n5120), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5458) );
  NAND4_X1 U6965 ( .A1(n5461), .A2(n5460), .A3(n5459), .A4(n5458), .ZN(n8461)
         );
  NAND2_X1 U6966 ( .A1(n8461), .A2(n9922), .ZN(n5462) );
  XNOR2_X1 U6967 ( .A(n5464), .B(n5462), .ZN(n8128) );
  NAND2_X1 U6968 ( .A1(n8129), .A2(n8128), .ZN(n5466) );
  INV_X1 U6969 ( .A(n5462), .ZN(n5463) );
  NAND2_X1 U6970 ( .A1(n5464), .A2(n5463), .ZN(n5465) );
  NAND2_X1 U6971 ( .A1(n5466), .A2(n5465), .ZN(n8050) );
  INV_X1 U6972 ( .A(n8050), .ZN(n5493) );
  NAND2_X1 U6973 ( .A1(n5470), .A2(SI_18_), .ZN(n5471) );
  MUX2_X1 U6974 ( .A(n7045), .B(n7139), .S(n6428), .Z(n5473) );
  INV_X1 U6975 ( .A(SI_19_), .ZN(n5472) );
  NAND2_X1 U6976 ( .A1(n5473), .A2(n5472), .ZN(n5497) );
  INV_X1 U6977 ( .A(n5473), .ZN(n5474) );
  NAND2_X1 U6978 ( .A1(n5474), .A2(SI_19_), .ZN(n5475) );
  NAND2_X1 U6979 ( .A1(n5497), .A2(n5475), .ZN(n5495) );
  XNOR2_X1 U6980 ( .A(n5496), .B(n5495), .ZN(n7044) );
  NAND2_X1 U6981 ( .A1(n7044), .A2(n5764), .ZN(n5477) );
  AOI22_X1 U6982 ( .A1(n5638), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5050), .B2(
        n6524), .ZN(n5476) );
  XNOR2_X1 U6983 ( .A(n8611), .B(n8055), .ZN(n5487) );
  NAND2_X1 U6984 ( .A1(n4430), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5486) );
  INV_X1 U6985 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5479) );
  INV_X1 U6986 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5478) );
  OAI21_X1 U6987 ( .B1(n5481), .B2(n5479), .A(n5478), .ZN(n5482) );
  NAND2_X1 U6988 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n5480) );
  AND2_X1 U6989 ( .A1(n5482), .A2(n5505), .ZN(n8455) );
  NAND2_X1 U6990 ( .A1(n5121), .A2(n8455), .ZN(n5485) );
  NAND2_X1 U6991 ( .A1(n5584), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U6992 ( .A1(n5120), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5483) );
  NAND4_X1 U6993 ( .A1(n5486), .A2(n5485), .A3(n5484), .A4(n5483), .ZN(n8477)
         );
  NAND2_X1 U6994 ( .A1(n8477), .A2(n9922), .ZN(n5488) );
  NAND2_X1 U6995 ( .A1(n5487), .A2(n5488), .ZN(n5494) );
  INV_X1 U6996 ( .A(n5487), .ZN(n5490) );
  INV_X1 U6997 ( .A(n5488), .ZN(n5489) );
  NAND2_X1 U6998 ( .A1(n5490), .A2(n5489), .ZN(n5491) );
  NAND2_X1 U6999 ( .A1(n5494), .A2(n5491), .ZN(n8049) );
  INV_X1 U7000 ( .A(n8049), .ZN(n5492) );
  MUX2_X1 U7001 ( .A(n7311), .B(n7215), .S(n6428), .Z(n5499) );
  INV_X1 U7002 ( .A(SI_20_), .ZN(n5498) );
  NAND2_X1 U7003 ( .A1(n5499), .A2(n5498), .ZN(n5517) );
  INV_X1 U7004 ( .A(n5499), .ZN(n5500) );
  NAND2_X1 U7005 ( .A1(n5500), .A2(SI_20_), .ZN(n5501) );
  XNOR2_X1 U7006 ( .A(n5516), .B(n5515), .ZN(n7214) );
  NAND2_X1 U7007 ( .A1(n7214), .A2(n5764), .ZN(n5503) );
  NAND2_X1 U7008 ( .A1(n5638), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5502) );
  XNOR2_X1 U7009 ( .A(n8605), .B(n5641), .ZN(n5512) );
  NAND2_X1 U7010 ( .A1(n4430), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U7011 ( .A1(n5584), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5509) );
  NAND2_X1 U7012 ( .A1(n5504), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5521) );
  INV_X1 U7013 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10067) );
  NAND2_X1 U7014 ( .A1(n5505), .A2(n10067), .ZN(n5506) );
  AND2_X1 U7015 ( .A1(n5521), .A2(n5506), .ZN(n8445) );
  NAND2_X1 U7016 ( .A1(n5121), .A2(n8445), .ZN(n5508) );
  INV_X1 U7017 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n10010) );
  OR2_X1 U7018 ( .A1(n5203), .A2(n10010), .ZN(n5507) );
  NOR2_X1 U7019 ( .A1(n8428), .A2(n9853), .ZN(n5511) );
  XNOR2_X1 U7020 ( .A(n5512), .B(n5511), .ZN(n8113) );
  NAND2_X1 U7021 ( .A1(n5512), .A2(n5511), .ZN(n5513) );
  NAND2_X1 U7022 ( .A1(n5514), .A2(n5513), .ZN(n8075) );
  MUX2_X1 U7023 ( .A(n7308), .B(n10219), .S(n6428), .Z(n5535) );
  XNOR2_X1 U7024 ( .A(n5535), .B(SI_21_), .ZN(n5533) );
  XNOR2_X1 U7025 ( .A(n5532), .B(n5533), .ZN(n7213) );
  NAND2_X1 U7026 ( .A1(n7213), .A2(n5764), .ZN(n5520) );
  NAND2_X1 U7027 ( .A1(n5638), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5519) );
  XNOR2_X1 U7028 ( .A(n8423), .B(n5641), .ZN(n5527) );
  NAND2_X1 U7029 ( .A1(n4430), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U7030 ( .A1(n5120), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5525) );
  INV_X1 U7031 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8076) );
  NAND2_X1 U7032 ( .A1(n5521), .A2(n8076), .ZN(n5522) );
  AND2_X1 U7033 ( .A1(n5549), .A2(n5522), .ZN(n8430) );
  NAND2_X1 U7034 ( .A1(n5121), .A2(n8430), .ZN(n5524) );
  NAND2_X1 U7035 ( .A1(n5584), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5523) );
  NOR2_X1 U7036 ( .A1(n8413), .A2(n9853), .ZN(n5528) );
  XNOR2_X1 U7037 ( .A(n5527), .B(n5528), .ZN(n8074) );
  NAND2_X1 U7038 ( .A1(n8075), .A2(n8074), .ZN(n5531) );
  INV_X1 U7039 ( .A(n5527), .ZN(n5529) );
  NAND2_X1 U7040 ( .A1(n5529), .A2(n5528), .ZN(n5530) );
  NAND2_X1 U7041 ( .A1(n5531), .A2(n5530), .ZN(n5556) );
  NAND2_X1 U7042 ( .A1(n5534), .A2(n5533), .ZN(n5538) );
  INV_X1 U7043 ( .A(n5535), .ZN(n5536) );
  NAND2_X1 U7044 ( .A1(n5536), .A2(SI_21_), .ZN(n5537) );
  MUX2_X1 U7045 ( .A(n10195), .B(n7405), .S(n6428), .Z(n5540) );
  INV_X1 U7046 ( .A(SI_22_), .ZN(n5539) );
  NAND2_X1 U7047 ( .A1(n5540), .A2(n5539), .ZN(n5560) );
  INV_X1 U7048 ( .A(n5540), .ZN(n5541) );
  NAND2_X1 U7049 ( .A1(n5541), .A2(SI_22_), .ZN(n5542) );
  NAND2_X1 U7050 ( .A1(n5560), .A2(n5542), .ZN(n5558) );
  XNOR2_X1 U7051 ( .A(n5559), .B(n5558), .ZN(n7403) );
  NAND2_X1 U7052 ( .A1(n7403), .A2(n5764), .ZN(n5544) );
  OR2_X1 U7053 ( .A1(n5782), .A2(n10195), .ZN(n5543) );
  XNOR2_X1 U7054 ( .A(n8594), .B(n8055), .ZN(n5554) );
  XNOR2_X1 U7055 ( .A(n5556), .B(n5554), .ZN(n8122) );
  NAND2_X1 U7056 ( .A1(n5120), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U7057 ( .A1(n4430), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5545) );
  AND2_X1 U7058 ( .A1(n5546), .A2(n5545), .ZN(n5553) );
  INV_X1 U7059 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U7060 ( .A1(n5549), .A2(n5548), .ZN(n5550) );
  NAND2_X1 U7061 ( .A1(n5569), .A2(n5550), .ZN(n8404) );
  OR2_X1 U7062 ( .A1(n5645), .A2(n8404), .ZN(n5552) );
  NAND2_X1 U7063 ( .A1(n5584), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5551) );
  INV_X1 U7064 ( .A(n8429), .ZN(n8396) );
  NAND2_X1 U7065 ( .A1(n8396), .A2(n9922), .ZN(n8121) );
  NAND2_X1 U7066 ( .A1(n8122), .A2(n8121), .ZN(n8120) );
  INV_X1 U7067 ( .A(n5554), .ZN(n5555) );
  OR2_X1 U7068 ( .A1(n5556), .A2(n5555), .ZN(n5557) );
  INV_X1 U7069 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5562) );
  INV_X1 U7070 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5561) );
  MUX2_X1 U7071 ( .A(n5562), .B(n5561), .S(n6428), .Z(n5564) );
  INV_X1 U7072 ( .A(SI_23_), .ZN(n5563) );
  NAND2_X1 U7073 ( .A1(n5564), .A2(n5563), .ZN(n5579) );
  INV_X1 U7074 ( .A(n5564), .ZN(n5565) );
  NAND2_X1 U7075 ( .A1(n5565), .A2(SI_23_), .ZN(n5566) );
  NAND2_X1 U7076 ( .A1(n5638), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5567) );
  XNOR2_X1 U7077 ( .A(n8589), .B(n8055), .ZN(n8039) );
  INV_X1 U7078 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8042) );
  NAND2_X1 U7079 ( .A1(n5569), .A2(n8042), .ZN(n5570) );
  NAND2_X1 U7080 ( .A1(n5582), .A2(n5570), .ZN(n8386) );
  OR2_X1 U7081 ( .A1(n8386), .A2(n5645), .ZN(n5573) );
  AOI22_X1 U7082 ( .A1(n5120), .A2(P2_REG0_REG_23__SCAN_IN), .B1(n4430), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U7083 ( .A1(n5584), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5571) );
  INV_X1 U7084 ( .A(n8414), .ZN(n8374) );
  NAND2_X1 U7085 ( .A1(n8374), .A2(n9922), .ZN(n8038) );
  AND2_X1 U7086 ( .A1(n8039), .A2(n8038), .ZN(n5577) );
  INV_X1 U7087 ( .A(n8039), .ZN(n5575) );
  INV_X1 U7088 ( .A(n8038), .ZN(n5574) );
  NAND2_X1 U7089 ( .A1(n5575), .A2(n5574), .ZN(n5576) );
  INV_X1 U7090 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7597) );
  MUX2_X1 U7091 ( .A(n7597), .B(n10172), .S(n6428), .Z(n5593) );
  XNOR2_X1 U7092 ( .A(n5593), .B(SI_24_), .ZN(n5592) );
  XNOR2_X1 U7093 ( .A(n5597), .B(n5592), .ZN(n7596) );
  NAND2_X1 U7094 ( .A1(n7596), .A2(n5764), .ZN(n5581) );
  NAND2_X1 U7095 ( .A1(n5638), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5580) );
  XNOR2_X1 U7096 ( .A(n8584), .B(n8055), .ZN(n5587) );
  XNOR2_X1 U7097 ( .A(n5589), .B(n5587), .ZN(n8108) );
  INV_X1 U7098 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10119) );
  NAND2_X1 U7099 ( .A1(n5582), .A2(n10119), .ZN(n5583) );
  NAND2_X1 U7100 ( .A1(n5617), .A2(n5583), .ZN(n8368) );
  AOI22_X1 U7101 ( .A1(n5120), .A2(P2_REG0_REG_24__SCAN_IN), .B1(n4406), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n5586) );
  NAND2_X1 U7102 ( .A1(n5584), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5585) );
  OAI211_X1 U7103 ( .C1(n8368), .C2(n5645), .A(n5586), .B(n5585), .ZN(n8395)
         );
  AND2_X1 U7104 ( .A1(n8395), .A2(n9922), .ZN(n8107) );
  NAND2_X1 U7105 ( .A1(n8108), .A2(n8107), .ZN(n5591) );
  INV_X1 U7106 ( .A(n5587), .ZN(n5588) );
  NAND2_X1 U7107 ( .A1(n5589), .A2(n5588), .ZN(n5590) );
  INV_X1 U7108 ( .A(n5592), .ZN(n5596) );
  INV_X1 U7109 ( .A(n5593), .ZN(n5594) );
  NAND2_X1 U7110 ( .A1(n5594), .A2(SI_24_), .ZN(n5595) );
  INV_X1 U7111 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7683) );
  INV_X1 U7112 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7746) );
  MUX2_X1 U7113 ( .A(n7683), .B(n7746), .S(n6428), .Z(n5599) );
  INV_X1 U7114 ( .A(SI_25_), .ZN(n5598) );
  NAND2_X1 U7115 ( .A1(n5599), .A2(n5598), .ZN(n5607) );
  INV_X1 U7116 ( .A(n5599), .ZN(n5600) );
  NAND2_X1 U7117 ( .A1(n5600), .A2(SI_25_), .ZN(n5601) );
  NAND2_X1 U7118 ( .A1(n5607), .A2(n5601), .ZN(n5608) );
  NAND2_X1 U7119 ( .A1(n7681), .A2(n5764), .ZN(n5603) );
  NAND2_X1 U7120 ( .A1(n5638), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5602) );
  XNOR2_X1 U7121 ( .A(n8581), .B(n5641), .ZN(n8083) );
  XNOR2_X1 U7122 ( .A(n5617), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n8359) );
  INV_X1 U7123 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n10204) );
  NAND2_X1 U7124 ( .A1(n5584), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U7125 ( .A1(n4430), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5604) );
  OAI211_X1 U7126 ( .C1(n5203), .C2(n10204), .A(n5605), .B(n5604), .ZN(n5606)
         );
  AOI21_X1 U7127 ( .B1(n8359), .B2(n5121), .A(n5606), .ZN(n8140) );
  OR2_X1 U7128 ( .A1(n8140), .A2(n9853), .ZN(n8082) );
  INV_X1 U7129 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7701) );
  INV_X1 U7130 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7896) );
  MUX2_X1 U7131 ( .A(n7701), .B(n7896), .S(n6428), .Z(n5610) );
  NAND2_X1 U7132 ( .A1(n5610), .A2(n9981), .ZN(n5632) );
  INV_X1 U7133 ( .A(n5610), .ZN(n5611) );
  NAND2_X1 U7134 ( .A1(n5611), .A2(SI_26_), .ZN(n5612) );
  NAND2_X1 U7135 ( .A1(n7700), .A2(n5764), .ZN(n5614) );
  NAND2_X1 U7136 ( .A1(n5638), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5613) );
  XNOR2_X1 U7137 ( .A(n8576), .B(n5641), .ZN(n5624) );
  INV_X1 U7138 ( .A(n5617), .ZN(n5616) );
  AND2_X1 U7139 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_26__SCAN_IN), 
        .ZN(n5615) );
  NAND2_X1 U7140 ( .A1(n5616), .A2(n5615), .ZN(n5643) );
  INV_X1 U7141 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8086) );
  INV_X1 U7142 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8141) );
  OAI21_X1 U7143 ( .B1(n5617), .B2(n8086), .A(n8141), .ZN(n5618) );
  AND2_X1 U7144 ( .A1(n5643), .A2(n5618), .ZN(n8342) );
  NAND2_X1 U7145 ( .A1(n8342), .A2(n5121), .ZN(n5623) );
  INV_X1 U7146 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n10138) );
  INV_X1 U7147 ( .A(n5584), .ZN(n5755) );
  NAND2_X1 U7148 ( .A1(n5120), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5620) );
  NAND2_X1 U7149 ( .A1(n4430), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5619) );
  OAI211_X1 U7150 ( .C1(n10138), .C2(n5755), .A(n5620), .B(n5619), .ZN(n5621)
         );
  INV_X1 U7151 ( .A(n5621), .ZN(n5622) );
  NOR2_X1 U7152 ( .A1(n8357), .A2(n9853), .ZN(n5625) );
  NAND2_X1 U7153 ( .A1(n5624), .A2(n5625), .ZN(n5629) );
  INV_X1 U7154 ( .A(n5624), .ZN(n5627) );
  INV_X1 U7155 ( .A(n5625), .ZN(n5626) );
  NAND2_X1 U7156 ( .A1(n5627), .A2(n5626), .ZN(n5628) );
  NAND2_X1 U7157 ( .A1(n5629), .A2(n5628), .ZN(n8135) );
  INV_X1 U7158 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8650) );
  INV_X1 U7159 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9998) );
  MUX2_X1 U7160 ( .A(n8650), .B(n9998), .S(n6428), .Z(n5635) );
  INV_X1 U7161 ( .A(SI_27_), .ZN(n5634) );
  NAND2_X1 U7162 ( .A1(n5635), .A2(n5634), .ZN(n5739) );
  INV_X1 U7163 ( .A(n5635), .ZN(n5636) );
  NAND2_X1 U7164 ( .A1(n5636), .A2(SI_27_), .ZN(n5637) );
  NAND2_X1 U7165 ( .A1(n7743), .A2(n5764), .ZN(n5640) );
  NAND2_X1 U7166 ( .A1(n5638), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5639) );
  XNOR2_X1 U7167 ( .A(n8569), .B(n5641), .ZN(n5651) );
  INV_X1 U7168 ( .A(n5643), .ZN(n5642) );
  NAND2_X1 U7169 ( .A1(n5642), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5697) );
  INV_X1 U7170 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10069) );
  NAND2_X1 U7171 ( .A1(n5643), .A2(n10069), .ZN(n5644) );
  NAND2_X1 U7172 ( .A1(n5697), .A2(n5644), .ZN(n8321) );
  INV_X1 U7173 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n10252) );
  NAND2_X1 U7174 ( .A1(n4406), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5647) );
  NAND2_X1 U7175 ( .A1(n5120), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5646) );
  OAI211_X1 U7176 ( .C1(n10252), .C2(n5755), .A(n5647), .B(n5646), .ZN(n5648)
         );
  INV_X1 U7177 ( .A(n5648), .ZN(n5649) );
  NOR2_X1 U7178 ( .A1(n8062), .A2(n9853), .ZN(n5652) );
  NAND2_X1 U7179 ( .A1(n5651), .A2(n5652), .ZN(n8067) );
  INV_X1 U7180 ( .A(n5651), .ZN(n5654) );
  INV_X1 U7181 ( .A(n5652), .ZN(n5653) );
  NAND2_X1 U7182 ( .A1(n5654), .A2(n5653), .ZN(n5655) );
  NAND2_X1 U7183 ( .A1(n5692), .A2(n5691), .ZN(n8066) );
  NOR4_X1 U7184 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n5659) );
  NOR4_X1 U7185 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n5658) );
  NOR4_X1 U7186 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n5657) );
  NOR4_X1 U7187 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n5656) );
  NAND4_X1 U7188 ( .A1(n5659), .A2(n5658), .A3(n5657), .A4(n5656), .ZN(n5677)
         );
  NOR4_X1 U7189 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n10245) );
  NOR2_X1 U7190 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .ZN(
        n5662) );
  NOR4_X1 U7191 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n5661) );
  NOR4_X1 U7192 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5660) );
  NAND4_X1 U7193 ( .A1(n10245), .A2(n5662), .A3(n5661), .A4(n5660), .ZN(n5676)
         );
  NAND2_X1 U7194 ( .A1(n5663), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5664) );
  MUX2_X1 U7195 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5664), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5665) );
  NAND2_X1 U7196 ( .A1(n5665), .A2(n4468), .ZN(n7682) );
  NAND2_X1 U7197 ( .A1(n5667), .A2(n5666), .ZN(n5668) );
  INV_X1 U7198 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5669) );
  XNOR2_X1 U7199 ( .A(n7598), .B(P2_B_REG_SCAN_IN), .ZN(n5671) );
  NAND2_X1 U7200 ( .A1(n4468), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5672) );
  MUX2_X1 U7201 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5672), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5674) );
  NAND2_X1 U7202 ( .A1(n5674), .A2(n5673), .ZN(n7702) );
  OAI21_X1 U7203 ( .B1(n5677), .B2(n5676), .A(n9861), .ZN(n6664) );
  AND2_X1 U7204 ( .A1(n7702), .A2(n7682), .ZN(n9867) );
  INV_X1 U7205 ( .A(n9867), .ZN(n5679) );
  INV_X1 U7206 ( .A(n7261), .ZN(n5681) );
  AND2_X1 U7207 ( .A1(n7270), .A2(n5681), .ZN(n5682) );
  NAND2_X1 U7208 ( .A1(n6664), .A2(n5682), .ZN(n5695) );
  OR2_X1 U7209 ( .A1(n5684), .A2(n5683), .ZN(n5685) );
  NAND2_X1 U7210 ( .A1(n5686), .A2(n5685), .ZN(n5966) );
  NOR2_X1 U7211 ( .A1(n5695), .A2(n9862), .ZN(n5704) );
  INV_X1 U7212 ( .A(n7310), .ZN(n5959) );
  NAND2_X1 U7213 ( .A1(n5959), .A2(n5687), .ZN(n7268) );
  NAND3_X1 U7214 ( .A1(n8066), .A2(n8138), .A3(n5693), .ZN(n5715) );
  NOR2_X1 U7215 ( .A1(n5689), .A2(n7451), .ZN(n5694) );
  NAND2_X1 U7216 ( .A1(n7310), .A2(n5694), .ZN(n9524) );
  NAND2_X1 U7217 ( .A1(n5695), .A2(n7264), .ZN(n5708) );
  INV_X1 U7218 ( .A(n9862), .ZN(n5696) );
  NAND2_X1 U7219 ( .A1(n5708), .A2(n5696), .ZN(n7978) );
  INV_X1 U7220 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8060) );
  NAND2_X1 U7221 ( .A1(n5697), .A2(n8060), .ZN(n5698) );
  INV_X1 U7222 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n5701) );
  NAND2_X1 U7223 ( .A1(n5120), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U7224 ( .A1(n4406), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5699) );
  OAI211_X1 U7225 ( .C1(n5701), .C2(n5755), .A(n5700), .B(n5699), .ZN(n5702)
         );
  AOI21_X1 U7226 ( .B1(n8305), .B2(n5121), .A(n5702), .ZN(n8286) );
  NAND2_X1 U7227 ( .A1(n7310), .A2(n7451), .ZN(n5969) );
  INV_X1 U7228 ( .A(n5969), .ZN(n5703) );
  NAND2_X1 U7229 ( .A1(n5704), .A2(n5703), .ZN(n8142) );
  OAI22_X1 U7230 ( .A1(n8286), .A2(n9832), .B1(n9831), .B2(n8357), .ZN(n5711)
         );
  INV_X1 U7231 ( .A(n7977), .ZN(n5706) );
  AND3_X1 U7232 ( .A1(n5706), .A2(n6425), .A3(n5966), .ZN(n5707) );
  NAND2_X1 U7233 ( .A1(n5708), .A2(n5707), .ZN(n5709) );
  OAI22_X1 U7234 ( .A1(n9840), .A2(n8321), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10069), .ZN(n5710) );
  NOR2_X1 U7235 ( .A1(n5711), .A2(n5710), .ZN(n5712) );
  INV_X1 U7236 ( .A(n5713), .ZN(n5714) );
  NAND2_X1 U7237 ( .A1(n5715), .A2(n5714), .ZN(P2_U3216) );
  INV_X1 U7238 ( .A(n5716), .ZN(n6680) );
  NAND2_X1 U7239 ( .A1(n6680), .A2(n8020), .ZN(n7408) );
  NAND2_X1 U7240 ( .A1(n6677), .A2(n6675), .ZN(n6909) );
  INV_X1 U7241 ( .A(n6909), .ZN(n5719) );
  INV_X1 U7242 ( .A(n5717), .ZN(n8176) );
  NAND2_X1 U7243 ( .A1(n5717), .A2(n8545), .ZN(n5807) );
  INV_X1 U7244 ( .A(n6910), .ZN(n5718) );
  NAND2_X1 U7245 ( .A1(n5719), .A2(n5718), .ZN(n6907) );
  NAND2_X1 U7246 ( .A1(n6907), .A2(n5807), .ZN(n7324) );
  NAND2_X1 U7247 ( .A1(n6956), .A2(n5720), .ZN(n5798) );
  INV_X1 U7248 ( .A(n6956), .ZN(n8175) );
  INV_X1 U7249 ( .A(n7333), .ZN(n7325) );
  NAND2_X1 U7250 ( .A1(n7323), .A2(n5798), .ZN(n6955) );
  INV_X1 U7251 ( .A(n6955), .ZN(n5722) );
  NAND2_X1 U7252 ( .A1(n7868), .A2(n7290), .ZN(n5799) );
  INV_X1 U7253 ( .A(n7868), .ZN(n8174) );
  NAND2_X1 U7254 ( .A1(n8174), .A2(n4645), .ZN(n7008) );
  NAND2_X1 U7255 ( .A1(n5799), .A2(n7008), .ZN(n6954) );
  NAND2_X1 U7256 ( .A1(n5722), .A2(n5721), .ZN(n7007) );
  INV_X1 U7257 ( .A(n7258), .ZN(n8173) );
  NAND2_X1 U7258 ( .A1(n8173), .A2(n7449), .ZN(n5935) );
  AND2_X1 U7259 ( .A1(n5935), .A2(n7008), .ZN(n5816) );
  NAND2_X1 U7260 ( .A1(n7007), .A2(n5816), .ZN(n5723) );
  NAND2_X1 U7261 ( .A1(n7258), .A2(n7015), .ZN(n5936) );
  NAND2_X1 U7262 ( .A1(n7276), .A2(n7349), .ZN(n5825) );
  INV_X1 U7263 ( .A(n7276), .ZN(n8172) );
  NAND2_X1 U7264 ( .A1(n8172), .A2(n9882), .ZN(n5820) );
  NAND2_X1 U7265 ( .A1(n7357), .A2(n9885), .ZN(n5839) );
  NAND2_X1 U7266 ( .A1(n8171), .A2(n7356), .ZN(n5829) );
  NAND2_X1 U7267 ( .A1(n5839), .A2(n5829), .ZN(n7354) );
  NAND2_X1 U7268 ( .A1(n7506), .A2(n7494), .ZN(n7501) );
  INV_X1 U7269 ( .A(n7506), .ZN(n8170) );
  INV_X1 U7270 ( .A(n7494), .ZN(n9892) );
  NAND2_X1 U7271 ( .A1(n8170), .A2(n9892), .ZN(n5796) );
  NAND2_X1 U7272 ( .A1(n7503), .A2(n7501), .ZN(n5724) );
  NAND2_X1 U7273 ( .A1(n9899), .A2(n8169), .ZN(n5836) );
  INV_X1 U7274 ( .A(n7562), .ZN(n5725) );
  OR2_X1 U7275 ( .A1(n9848), .A2(n9833), .ZN(n5943) );
  INV_X1 U7276 ( .A(n5943), .ZN(n5726) );
  NAND2_X1 U7277 ( .A1(n9848), .A2(n9833), .ZN(n5942) );
  NAND2_X1 U7278 ( .A1(n9920), .A2(n7757), .ZN(n5931) );
  OR2_X1 U7279 ( .A1(n9525), .A2(n8032), .ZN(n5854) );
  NAND2_X1 U7280 ( .A1(n9525), .A2(n8032), .ZN(n5853) );
  NAND2_X1 U7281 ( .A1(n8267), .A2(n8155), .ZN(n5857) );
  INV_X1 U7282 ( .A(n7801), .ZN(n7799) );
  NAND2_X1 U7283 ( .A1(n8538), .A2(n8503), .ZN(n5862) );
  NAND2_X1 U7284 ( .A1(n5863), .A2(n5862), .ZN(n8526) );
  INV_X1 U7285 ( .A(n8526), .ZN(n8528) );
  OR2_X1 U7286 ( .A1(n8626), .A2(n8154), .ZN(n5865) );
  INV_X1 U7287 ( .A(n5865), .ZN(n5727) );
  NAND2_X1 U7288 ( .A1(n8626), .A2(n8154), .ZN(n5864) );
  NAND2_X1 U7289 ( .A1(n8622), .A2(n8501), .ZN(n5870) );
  NAND2_X1 U7290 ( .A1(n5869), .A2(n5870), .ZN(n8485) );
  INV_X1 U7291 ( .A(n8461), .ZN(n8274) );
  OR2_X1 U7292 ( .A1(n8615), .A2(n8274), .ZN(n5881) );
  NAND2_X1 U7293 ( .A1(n8615), .A2(n8274), .ZN(n5873) );
  NAND2_X1 U7294 ( .A1(n5881), .A2(n5873), .ZN(n5930) );
  NAND2_X1 U7295 ( .A1(n8473), .A2(n5873), .ZN(n8459) );
  INV_X1 U7296 ( .A(n8477), .ZN(n8277) );
  OR2_X1 U7297 ( .A1(n8611), .A2(n8277), .ZN(n5885) );
  NAND2_X1 U7298 ( .A1(n8611), .A2(n8277), .ZN(n8436) );
  NAND2_X1 U7299 ( .A1(n8605), .A2(n8428), .ZN(n5888) );
  NAND2_X1 U7300 ( .A1(n5876), .A2(n5888), .ZN(n8440) );
  INV_X1 U7301 ( .A(n8436), .ZN(n5728) );
  NOR2_X1 U7302 ( .A1(n8440), .A2(n5728), .ZN(n5729) );
  NAND2_X1 U7303 ( .A1(n8601), .A2(n8413), .ZN(n8410) );
  NAND2_X1 U7304 ( .A1(n5889), .A2(n8410), .ZN(n8425) );
  NAND2_X1 U7305 ( .A1(n8594), .A2(n8429), .ZN(n5879) );
  NAND2_X1 U7306 ( .A1(n5894), .A2(n5879), .ZN(n8279) );
  INV_X1 U7307 ( .A(n8410), .ZN(n5891) );
  NOR2_X1 U7308 ( .A1(n8279), .A2(n5891), .ZN(n5731) );
  OR2_X1 U7309 ( .A1(n8589), .A2(n8414), .ZN(n5897) );
  NAND2_X1 U7310 ( .A1(n8589), .A2(n8414), .ZN(n5896) );
  NAND2_X1 U7311 ( .A1(n5897), .A2(n5896), .ZN(n8391) );
  INV_X1 U7312 ( .A(n5894), .ZN(n8392) );
  NOR2_X1 U7313 ( .A1(n8391), .A2(n8392), .ZN(n5732) );
  XNOR2_X1 U7314 ( .A(n8584), .B(n8395), .ZN(n8373) );
  INV_X1 U7315 ( .A(n8395), .ZN(n8356) );
  OR2_X1 U7316 ( .A1(n8584), .A2(n8356), .ZN(n5901) );
  NAND2_X1 U7317 ( .A1(n8581), .A2(n8140), .ZN(n5907) );
  NAND2_X1 U7318 ( .A1(n8354), .A2(n8353), .ZN(n5733) );
  NAND2_X1 U7319 ( .A1(n8576), .A2(n8357), .ZN(n5909) );
  NAND2_X1 U7320 ( .A1(n5905), .A2(n5909), .ZN(n8334) );
  INV_X1 U7321 ( .A(n8334), .ZN(n8337) );
  NAND2_X1 U7322 ( .A1(n8338), .A2(n8337), .ZN(n5734) );
  INV_X1 U7323 ( .A(n8325), .ZN(n5952) );
  NAND2_X1 U7324 ( .A1(n8326), .A2(n5952), .ZN(n5736) );
  OR2_X1 U7325 ( .A1(n8569), .A2(n8062), .ZN(n5735) );
  INV_X1 U7326 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n10222) );
  INV_X1 U7327 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7886) );
  MUX2_X1 U7328 ( .A(n10222), .B(n7886), .S(n6428), .Z(n5746) );
  XNOR2_X1 U7329 ( .A(n5746), .B(SI_28_), .ZN(n5743) );
  NAND2_X1 U7330 ( .A1(n7885), .A2(n5764), .ZN(n5741) );
  OR2_X1 U7331 ( .A1(n5782), .A2(n10222), .ZN(n5740) );
  NAND2_X1 U7332 ( .A1(n8564), .A2(n8286), .ZN(n5914) );
  INV_X1 U7333 ( .A(n8308), .ZN(n5954) );
  NAND2_X1 U7334 ( .A1(n8309), .A2(n5954), .ZN(n5742) );
  NAND2_X1 U7335 ( .A1(n5742), .A2(n5913), .ZN(n8283) );
  INV_X1 U7336 ( .A(SI_28_), .ZN(n5745) );
  NAND2_X1 U7337 ( .A1(n5746), .A2(n5745), .ZN(n5747) );
  INV_X1 U7338 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n10016) );
  INV_X1 U7339 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10218) );
  MUX2_X1 U7340 ( .A(n10016), .B(n10218), .S(n6428), .Z(n5757) );
  XNOR2_X1 U7341 ( .A(n5757), .B(SI_29_), .ZN(n5749) );
  NAND2_X1 U7342 ( .A1(n8781), .A2(n5764), .ZN(n5751) );
  OR2_X1 U7343 ( .A1(n5782), .A2(n10016), .ZN(n5750) );
  INV_X1 U7344 ( .A(n5752), .ZN(n8295) );
  INV_X1 U7345 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n10254) );
  NAND2_X1 U7346 ( .A1(n5120), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U7347 ( .A1(n4430), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5753) );
  OAI211_X1 U7348 ( .C1(n10254), .C2(n5755), .A(n5754), .B(n5753), .ZN(n5756)
         );
  AOI21_X1 U7349 ( .B1(n8295), .B2(n5121), .A(n5756), .ZN(n8163) );
  OR2_X1 U7350 ( .A1(n8292), .A2(n8163), .ZN(n5794) );
  NAND2_X1 U7351 ( .A1(n8292), .A2(n8163), .ZN(n5790) );
  INV_X1 U7352 ( .A(SI_29_), .ZN(n5760) );
  INV_X1 U7353 ( .A(n5757), .ZN(n5758) );
  MUX2_X1 U7354 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n6428), .Z(n5776) );
  XNOR2_X1 U7355 ( .A(n5776), .B(SI_30_), .ZN(n5761) );
  INV_X1 U7356 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n5762) );
  NOR2_X1 U7357 ( .A1(n5782), .A2(n5762), .ZN(n5763) );
  NAND2_X1 U7358 ( .A1(n5120), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5767) );
  NAND2_X1 U7359 ( .A1(n4406), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5766) );
  NAND2_X1 U7360 ( .A1(n5584), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U7361 ( .A1(n7854), .A2(n5804), .ZN(n5768) );
  OAI21_X1 U7362 ( .B1(n9508), .B2(n5768), .A(n5790), .ZN(n5773) );
  INV_X1 U7363 ( .A(n5768), .ZN(n5772) );
  INV_X1 U7364 ( .A(n9508), .ZN(n7851) );
  NAND2_X1 U7365 ( .A1(n5120), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5771) );
  NAND2_X1 U7366 ( .A1(n4430), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5770) );
  NAND2_X1 U7367 ( .A1(n5584), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5769) );
  AND3_X1 U7368 ( .A1(n5771), .A2(n5770), .A3(n5769), .ZN(n8288) );
  OR2_X1 U7369 ( .A1(n7851), .A2(n8288), .ZN(n5920) );
  OAI22_X1 U7370 ( .A1(n8284), .A2(n5773), .B1(n5772), .B2(n5920), .ZN(n5783)
         );
  INV_X1 U7371 ( .A(n5776), .ZN(n5775) );
  INV_X1 U7372 ( .A(SI_30_), .ZN(n5774) );
  NOR2_X1 U7373 ( .A1(n5775), .A2(n5774), .ZN(n5777) );
  MUX2_X1 U7374 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n6428), .Z(n5779) );
  XNOR2_X1 U7375 ( .A(n5779), .B(SI_31_), .ZN(n5780) );
  INV_X1 U7376 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n7847) );
  NOR2_X1 U7377 ( .A1(n8556), .A2(n7854), .ZN(n5923) );
  INV_X1 U7378 ( .A(n8288), .ZN(n8162) );
  NOR2_X1 U7379 ( .A1(n9508), .A2(n8162), .ZN(n5795) );
  NOR2_X1 U7380 ( .A1(n5923), .A2(n5795), .ZN(n5928) );
  INV_X1 U7381 ( .A(n8556), .ZN(n7852) );
  INV_X1 U7382 ( .A(n7854), .ZN(n8161) );
  NOR2_X1 U7383 ( .A1(n7852), .A2(n8161), .ZN(n5924) );
  AOI21_X1 U7384 ( .B1(n5783), .B2(n5928), .A(n5924), .ZN(n5784) );
  XNOR2_X1 U7385 ( .A(n5784), .B(n7451), .ZN(n5786) );
  NAND2_X1 U7386 ( .A1(n5959), .A2(n5804), .ZN(n6674) );
  INV_X1 U7387 ( .A(n5920), .ZN(n5787) );
  NOR2_X1 U7388 ( .A1(n5924), .A2(n5787), .ZN(n5929) );
  NOR2_X1 U7389 ( .A1(n7451), .A2(n7307), .ZN(n5788) );
  NAND2_X1 U7390 ( .A1(n5788), .A2(n7404), .ZN(n5922) );
  MUX2_X1 U7391 ( .A(n5928), .B(n5929), .S(n5922), .Z(n5927) );
  INV_X1 U7392 ( .A(n5913), .ZN(n5789) );
  AOI21_X1 U7393 ( .B1(n5789), .B2(n5922), .A(n8282), .ZN(n5915) );
  OAI21_X1 U7394 ( .B1(n8324), .B2(n8311), .A(n5914), .ZN(n5792) );
  INV_X1 U7395 ( .A(n5790), .ZN(n5791) );
  AOI21_X1 U7396 ( .B1(n5915), .B2(n5792), .A(n5791), .ZN(n5793) );
  MUX2_X1 U7397 ( .A(n5794), .B(n5793), .S(n5922), .Z(n5921) );
  INV_X1 U7398 ( .A(n5795), .ZN(n5919) );
  INV_X1 U7399 ( .A(n5905), .ZN(n5910) );
  AND2_X1 U7400 ( .A1(n5836), .A2(n5796), .ZN(n5833) );
  INV_X1 U7401 ( .A(n5922), .ZN(n5911) );
  AND2_X1 U7402 ( .A1(n5936), .A2(n5799), .ZN(n5797) );
  MUX2_X1 U7403 ( .A(n5797), .B(n5816), .S(n5922), .Z(n5819) );
  NAND2_X1 U7404 ( .A1(n5799), .A2(n5798), .ZN(n5801) );
  NAND2_X1 U7405 ( .A1(n5936), .A2(n5825), .ZN(n5800) );
  AOI21_X1 U7406 ( .B1(n5819), .B2(n5801), .A(n5800), .ZN(n5813) );
  INV_X1 U7407 ( .A(n8020), .ZN(n9870) );
  NAND2_X1 U7408 ( .A1(n5716), .A2(n9870), .ZN(n8017) );
  NAND2_X1 U7409 ( .A1(n6675), .A2(n8017), .ZN(n5802) );
  NAND3_X1 U7410 ( .A1(n5807), .A2(n6667), .A3(n5802), .ZN(n5803) );
  NAND2_X1 U7411 ( .A1(n5803), .A2(n5805), .ZN(n5810) );
  AND2_X1 U7412 ( .A1(n8017), .A2(n5804), .ZN(n5806) );
  OAI211_X1 U7413 ( .C1(n6677), .C2(n5806), .A(n5805), .B(n6675), .ZN(n5808)
         );
  NAND2_X1 U7414 ( .A1(n5808), .A2(n5807), .ZN(n5809) );
  MUX2_X1 U7415 ( .A(n5810), .B(n5809), .S(n5922), .Z(n5811) );
  NAND3_X1 U7416 ( .A1(n5811), .A2(n7325), .A3(n5819), .ZN(n5812) );
  OAI21_X1 U7417 ( .B1(n5911), .B2(n5813), .A(n5812), .ZN(n5814) );
  NAND2_X1 U7418 ( .A1(n5814), .A2(n5820), .ZN(n5824) );
  INV_X1 U7419 ( .A(n5935), .ZN(n5818) );
  NAND2_X1 U7420 ( .A1(n5816), .A2(n5815), .ZN(n5817) );
  OAI21_X1 U7421 ( .B1(n5819), .B2(n5818), .A(n5817), .ZN(n5821) );
  NAND2_X1 U7422 ( .A1(n5821), .A2(n5820), .ZN(n5822) );
  NAND2_X1 U7423 ( .A1(n5822), .A2(n5911), .ZN(n5823) );
  NAND2_X1 U7424 ( .A1(n5824), .A2(n5823), .ZN(n5828) );
  NOR2_X1 U7425 ( .A1(n5825), .A2(n5922), .ZN(n5826) );
  NOR2_X1 U7426 ( .A1(n5826), .A2(n7354), .ZN(n5827) );
  NAND2_X1 U7427 ( .A1(n5828), .A2(n5827), .ZN(n5841) );
  AND2_X1 U7428 ( .A1(n7491), .A2(n5829), .ZN(n5831) );
  INV_X1 U7429 ( .A(n7501), .ZN(n5830) );
  AOI21_X1 U7430 ( .B1(n5841), .B2(n5831), .A(n5830), .ZN(n5832) );
  MUX2_X1 U7431 ( .A(n5833), .B(n5832), .S(n5911), .Z(n5834) );
  NAND2_X1 U7432 ( .A1(n5834), .A2(n5835), .ZN(n5838) );
  AND2_X1 U7433 ( .A1(n5837), .A2(n5842), .ZN(n5840) );
  NAND2_X1 U7434 ( .A1(n5838), .A2(n5840), .ZN(n5847) );
  NAND4_X1 U7435 ( .A1(n5841), .A2(n7491), .A3(n5840), .A4(n5839), .ZN(n5843)
         );
  NAND3_X1 U7436 ( .A1(n5843), .A2(n5943), .A3(n5842), .ZN(n5846) );
  NAND2_X1 U7437 ( .A1(n5942), .A2(n5844), .ZN(n5845) );
  NAND3_X1 U7438 ( .A1(n5849), .A2(n5931), .A3(n5942), .ZN(n5848) );
  NAND2_X1 U7439 ( .A1(n5848), .A2(n5932), .ZN(n5852) );
  AOI21_X1 U7440 ( .B1(n5850), .B2(n5931), .A(n4751), .ZN(n5851) );
  MUX2_X1 U7441 ( .A(n5852), .B(n5851), .S(n5911), .Z(n5856) );
  MUX2_X1 U7442 ( .A(n5854), .B(n5853), .S(n5922), .Z(n5855) );
  OAI211_X1 U7443 ( .C1(n5856), .C2(n7755), .A(n7801), .B(n5855), .ZN(n5861)
         );
  NAND2_X1 U7444 ( .A1(n5865), .A2(n5864), .ZN(n8504) );
  INV_X1 U7445 ( .A(n8504), .ZN(n5860) );
  MUX2_X1 U7446 ( .A(n5858), .B(n5857), .S(n5911), .Z(n5859) );
  MUX2_X1 U7447 ( .A(n5863), .B(n5862), .S(n5922), .Z(n5867) );
  MUX2_X1 U7448 ( .A(n5865), .B(n5864), .S(n5922), .Z(n5866) );
  OAI211_X1 U7449 ( .C1(n5867), .C2(n8504), .A(n4734), .B(n5866), .ZN(n5868)
         );
  NAND2_X1 U7450 ( .A1(n5873), .A2(n5870), .ZN(n5871) );
  MUX2_X1 U7451 ( .A(n4730), .B(n5871), .S(n5911), .Z(n5872) );
  INV_X1 U7452 ( .A(n5885), .ZN(n5874) );
  OAI211_X1 U7453 ( .C1(n5874), .C2(n5873), .A(n5888), .B(n8436), .ZN(n5875)
         );
  NAND2_X1 U7454 ( .A1(n5889), .A2(n5876), .ZN(n5884) );
  OAI211_X1 U7455 ( .C1(n5877), .C2(n5884), .A(n5879), .B(n8410), .ZN(n5878)
         );
  MUX2_X1 U7456 ( .A(n5879), .B(n5878), .S(n5922), .Z(n5880) );
  NAND2_X1 U7457 ( .A1(n5880), .A2(n4969), .ZN(n5900) );
  INV_X1 U7458 ( .A(n5881), .ZN(n5882) );
  OAI21_X1 U7459 ( .B1(n5883), .B2(n5882), .A(n8436), .ZN(n5887) );
  INV_X1 U7460 ( .A(n5884), .ZN(n5886) );
  NAND3_X1 U7461 ( .A1(n5887), .A2(n5886), .A3(n5885), .ZN(n5893) );
  INV_X1 U7462 ( .A(n5888), .ZN(n5890) );
  OAI21_X1 U7463 ( .B1(n5891), .B2(n5890), .A(n5889), .ZN(n5892) );
  AOI21_X1 U7464 ( .B1(n5893), .B2(n5892), .A(n5922), .ZN(n5895) );
  MUX2_X1 U7465 ( .A(n5922), .B(n5895), .S(n5894), .Z(n5899) );
  MUX2_X1 U7466 ( .A(n5897), .B(n5896), .S(n5922), .Z(n5898) );
  OAI211_X1 U7467 ( .C1(n5900), .C2(n5899), .A(n8373), .B(n5898), .ZN(n5904)
         );
  NAND2_X1 U7468 ( .A1(n8584), .A2(n8356), .ZN(n5902) );
  MUX2_X1 U7469 ( .A(n5902), .B(n5901), .S(n5922), .Z(n5903) );
  NAND2_X1 U7470 ( .A1(n5909), .A2(n5907), .ZN(n5908) );
  NAND3_X1 U7471 ( .A1(n8324), .A2(n5911), .A3(n8311), .ZN(n5912) );
  NAND2_X1 U7472 ( .A1(n5913), .A2(n5912), .ZN(n5916) );
  OAI211_X1 U7473 ( .C1(n5917), .C2(n5916), .A(n5915), .B(n5914), .ZN(n5918)
         );
  NAND4_X1 U7474 ( .A1(n5921), .A2(n5920), .A3(n5919), .A4(n5918), .ZN(n5926)
         );
  MUX2_X1 U7475 ( .A(n5924), .B(n5923), .S(n5922), .Z(n5925) );
  AOI21_X1 U7476 ( .B1(n5927), .B2(n5926), .A(n5925), .ZN(n5960) );
  INV_X1 U7477 ( .A(n5960), .ZN(n5965) );
  OAI21_X1 U7478 ( .B1(n5959), .B2(n6673), .A(n9922), .ZN(n5964) );
  INV_X1 U7479 ( .A(n5928), .ZN(n5957) );
  INV_X1 U7480 ( .A(n5929), .ZN(n5956) );
  INV_X1 U7481 ( .A(n8373), .ZN(n8364) );
  INV_X1 U7482 ( .A(n8279), .ZN(n8409) );
  INV_X1 U7483 ( .A(n5930), .ZN(n8474) );
  OR2_X1 U7484 ( .A1(n6954), .A2(n7333), .ZN(n5934) );
  NAND3_X1 U7485 ( .A1(n6675), .A2(n8017), .A3(n5959), .ZN(n5933) );
  NOR2_X1 U7486 ( .A1(n5934), .A2(n5933), .ZN(n5939) );
  NAND2_X1 U7487 ( .A1(n5936), .A2(n5935), .ZN(n7009) );
  INV_X1 U7488 ( .A(n7009), .ZN(n5938) );
  NOR2_X1 U7489 ( .A1(n6677), .A2(n6910), .ZN(n5937) );
  NAND4_X1 U7490 ( .A1(n5939), .A2(n5938), .A3(n7351), .A4(n5937), .ZN(n5940)
         );
  NOR2_X1 U7491 ( .A1(n5940), .A2(n7354), .ZN(n5941) );
  NAND4_X1 U7492 ( .A1(n5941), .A2(n7562), .A3(n7498), .A4(n7491), .ZN(n5944)
         );
  NAND2_X1 U7493 ( .A1(n5943), .A2(n5942), .ZN(n9849) );
  NOR2_X1 U7494 ( .A1(n5944), .A2(n9849), .ZN(n5945) );
  AND4_X1 U7495 ( .A1(n7801), .A2(n7751), .A3(n7790), .A4(n5945), .ZN(n5946)
         );
  NAND2_X1 U7496 ( .A1(n8528), .A2(n5946), .ZN(n5947) );
  NOR2_X1 U7497 ( .A1(n8504), .A2(n5947), .ZN(n5948) );
  NAND4_X1 U7498 ( .A1(n8460), .A2(n4734), .A3(n8474), .A4(n5948), .ZN(n5949)
         );
  NOR2_X1 U7499 ( .A1(n8440), .A2(n5949), .ZN(n5950) );
  NAND4_X1 U7500 ( .A1(n4969), .A2(n8409), .A3(n5730), .A4(n5950), .ZN(n5951)
         );
  NOR3_X1 U7501 ( .A1(n8350), .A2(n8364), .A3(n5951), .ZN(n5953) );
  NAND4_X1 U7502 ( .A1(n5954), .A2(n8337), .A3(n5953), .A4(n5952), .ZN(n5955)
         );
  NOR4_X1 U7503 ( .A1(n5957), .A2(n5956), .A3(n8282), .A4(n5955), .ZN(n5958)
         );
  XNOR2_X1 U7504 ( .A(n5958), .B(n7451), .ZN(n5962) );
  AOI21_X1 U7505 ( .B1(n5960), .B2(n6673), .A(n5959), .ZN(n5961) );
  AOI21_X1 U7506 ( .B1(n5962), .B2(n7307), .A(n5961), .ZN(n5963) );
  AOI21_X1 U7507 ( .B1(n5965), .B2(n5964), .A(n5963), .ZN(n5967) );
  NOR2_X1 U7508 ( .A1(n5966), .A2(P2_U3152), .ZN(n7540) );
  NOR4_X1 U7509 ( .A1(n9862), .A2(n8649), .A3(n5969), .A4(n8502), .ZN(n5971)
         );
  INV_X1 U7510 ( .A(n7540), .ZN(n6726) );
  OAI21_X1 U7511 ( .B1(n6726), .B2(n5689), .A(P2_B_REG_SCAN_IN), .ZN(n5970) );
  OR2_X1 U7512 ( .A1(n5971), .A2(n5970), .ZN(n5972) );
  NAND2_X1 U7513 ( .A1(n5973), .A2(n5972), .ZN(P2_U3244) );
  NOR2_X1 U7514 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5978) );
  NOR2_X1 U7515 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5977) );
  NOR2_X1 U7516 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5976) );
  NOR2_X1 U7517 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5975) );
  NAND4_X1 U7518 ( .A1(n5978), .A2(n5977), .A3(n5976), .A4(n5975), .ZN(n6015)
         );
  NOR2_X1 U7519 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5982) );
  NOR2_X1 U7520 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5981) );
  NOR2_X1 U7521 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5980) );
  NOR2_X1 U7522 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5979) );
  NAND4_X1 U7523 ( .A1(n5982), .A2(n5981), .A3(n5980), .A4(n5979), .ZN(n5983)
         );
  NOR2_X1 U7524 ( .A1(n6015), .A2(n5983), .ZN(n5984) );
  NOR2_X1 U7525 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5986) );
  XNOR2_X2 U7526 ( .A(n5988), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9487) );
  INV_X1 U7527 ( .A(n9487), .ZN(n5990) );
  INV_X1 U7528 ( .A(n5989), .ZN(n7843) );
  NAND2_X1 U7529 ( .A1(n4403), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5999) );
  NOR2_X2 U7530 ( .A1(n9487), .A2(n9492), .ZN(n6101) );
  INV_X2 U7531 ( .A(n6086), .ZN(n6248) );
  NAND2_X1 U7532 ( .A1(n6087), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U7533 ( .A1(n6115), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U7534 ( .A1(n6144), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U7535 ( .A1(n6184), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6196) );
  INV_X1 U7536 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6195) );
  INV_X1 U7537 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8699) );
  INV_X1 U7538 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6019) );
  INV_X1 U7539 ( .A(n6279), .ZN(n5992) );
  NAND2_X1 U7540 ( .A1(n5992), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6288) );
  INV_X1 U7541 ( .A(n6289), .ZN(n5993) );
  NAND2_X1 U7542 ( .A1(n5993), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6301) );
  INV_X1 U7543 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5994) );
  NAND2_X1 U7544 ( .A1(n6289), .A2(n5994), .ZN(n5995) );
  AND2_X1 U7545 ( .A1(n6301), .A2(n5995), .ZN(n9200) );
  NAND2_X1 U7546 ( .A1(n6374), .A2(n9200), .ZN(n5997) );
  NAND2_X1 U7547 ( .A1(n6313), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5996) );
  NAND4_X1 U7548 ( .A1(n5999), .A2(n5998), .A3(n5997), .A4(n5996), .ZN(n9388)
         );
  INV_X1 U7549 ( .A(n9388), .ZN(n8659) );
  NAND2_X1 U7550 ( .A1(n6004), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U7551 ( .A1(n7596), .A2(n8780), .ZN(n6008) );
  NAND2_X1 U7552 ( .A1(n6266), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6007) );
  INV_X1 U7553 ( .A(n9199), .ZN(n9460) );
  NAND2_X1 U7554 ( .A1(n6964), .A2(n8780), .ZN(n6018) );
  INV_X1 U7555 ( .A(n6153), .ZN(n6266) );
  INV_X1 U7556 ( .A(n6140), .ZN(n6014) );
  NAND2_X1 U7557 ( .A1(n6014), .A2(n6013), .ZN(n6023) );
  NAND2_X1 U7558 ( .A1(n6344), .A2(n6342), .ZN(n6241) );
  NAND2_X1 U7559 ( .A1(n6241), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6016) );
  XNOR2_X1 U7560 ( .A(n6016), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9093) );
  AOI22_X1 U7561 ( .A1(n6266), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9093), .B2(
        n6243), .ZN(n6017) );
  INV_X1 U7562 ( .A(n9421), .ZN(n9305) );
  AND2_X1 U7563 ( .A1(n6235), .A2(n6019), .ZN(n6020) );
  OR2_X1 U7564 ( .A1(n6020), .A2(n6246), .ZN(n9302) );
  AOI22_X1 U7565 ( .A1(n6097), .A2(P1_REG0_REG_18__SCAN_IN), .B1(n6313), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n6022) );
  NAND2_X1 U7566 ( .A1(n6248), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6021) );
  OAI211_X1 U7567 ( .C1(n9302), .C2(n6264), .A(n6022), .B(n6021), .ZN(n9411)
         );
  INV_X1 U7568 ( .A(n9411), .ZN(n9317) );
  NAND2_X1 U7569 ( .A1(n6659), .A2(n8780), .ZN(n6030) );
  INV_X1 U7570 ( .A(n6023), .ZN(n6026) );
  NOR2_X1 U7571 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n10247) );
  NOR2_X1 U7572 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n6024) );
  AND2_X1 U7573 ( .A1(n10247), .A2(n6024), .ZN(n6025) );
  NAND2_X1 U7574 ( .A1(n6026), .A2(n6025), .ZN(n6190) );
  INV_X1 U7575 ( .A(n6190), .ZN(n6027) );
  INV_X1 U7576 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10236) );
  NAND2_X1 U7577 ( .A1(n6027), .A2(n10236), .ZN(n6204) );
  OAI21_X1 U7578 ( .B1(n6216), .B2(P1_IR_REG_15__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6028) );
  XNOR2_X1 U7579 ( .A(n6028), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9071) );
  AOI22_X1 U7580 ( .A1(n9071), .A2(n6243), .B1(n6254), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n6029) );
  OR2_X1 U7581 ( .A1(n6222), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6031) );
  AND2_X1 U7582 ( .A1(n6233), .A2(n6031), .ZN(n9334) );
  NAND2_X1 U7583 ( .A1(n9334), .A2(n6374), .ZN(n6035) );
  NAND2_X1 U7584 ( .A1(n6097), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7585 ( .A1(n6313), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6033) );
  NAND2_X1 U7586 ( .A1(n6248), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6032) );
  NAND4_X1 U7587 ( .A1(n6035), .A2(n6034), .A3(n6033), .A4(n6032), .ZN(n9431)
         );
  NAND2_X1 U7588 ( .A1(n6529), .A2(n8780), .ZN(n6041) );
  INV_X1 U7589 ( .A(n6153), .ZN(n6254) );
  OAI21_X1 U7590 ( .B1(n6023), .B2(P1_IR_REG_9__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6165) );
  INV_X1 U7591 ( .A(n10247), .ZN(n6036) );
  NAND2_X1 U7592 ( .A1(n6036), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U7593 ( .A1(n6165), .A2(n6037), .ZN(n6039) );
  INV_X1 U7594 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6038) );
  XNOR2_X1 U7595 ( .A(n6039), .B(n6038), .ZN(n7048) );
  AOI22_X1 U7596 ( .A1(n6266), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7048), .B2(
        n6243), .ZN(n6040) );
  NAND2_X1 U7597 ( .A1(n4403), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6046) );
  NAND2_X1 U7598 ( .A1(n6248), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6045) );
  OR2_X1 U7599 ( .A1(n6184), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6042) );
  AND2_X1 U7600 ( .A1(n6042), .A2(n6196), .ZN(n7587) );
  NAND2_X1 U7601 ( .A1(n6374), .A2(n7587), .ZN(n6044) );
  NAND2_X1 U7602 ( .A1(n6313), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6043) );
  NAND4_X1 U7603 ( .A1(n6046), .A2(n6045), .A3(n6044), .A4(n6043), .ZN(n9041)
         );
  NAND2_X1 U7604 ( .A1(n4403), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6050) );
  AOI21_X1 U7605 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6047) );
  NOR2_X1 U7606 ( .A1(n6047), .A2(n6115), .ZN(n6750) );
  NAND2_X1 U7607 ( .A1(n6374), .A2(n6750), .ZN(n6049) );
  NAND2_X1 U7608 ( .A1(n6313), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6048) );
  OR2_X1 U7609 ( .A1(n6009), .A2(n6121), .ZN(n6052) );
  XNOR2_X1 U7610 ( .A(n6052), .B(n6051), .ZN(n9594) );
  NAND2_X1 U7611 ( .A1(n6134), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7612 ( .A1(n9768), .A2(n9763), .ZN(n8977) );
  AND2_X1 U7613 ( .A1(n8973), .A2(n8977), .ZN(n6933) );
  INV_X1 U7614 ( .A(n6933), .ZN(n6113) );
  NAND2_X1 U7615 ( .A1(n6100), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6058) );
  INV_X1 U7616 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6054) );
  NAND2_X1 U7617 ( .A1(n6098), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6056) );
  NAND2_X1 U7618 ( .A1(n6101), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6055) );
  NAND4_X2 U7619 ( .A1(n6058), .A2(n6057), .A3(n6056), .A4(n6055), .ZN(n6576)
         );
  INV_X1 U7620 ( .A(n6576), .ZN(n6996) );
  NAND2_X1 U7621 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6059) );
  XNOR2_X1 U7622 ( .A(n6059), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6490) );
  INV_X1 U7623 ( .A(n6490), .ZN(n6060) );
  OR2_X1 U7624 ( .A1(n6498), .A2(n6060), .ZN(n6061) );
  NAND2_X1 U7625 ( .A1(n6996), .A2(n9700), .ZN(n6360) );
  INV_X1 U7626 ( .A(n9700), .ZN(n9727) );
  NAND2_X1 U7627 ( .A1(n6576), .A2(n9727), .ZN(n8795) );
  NAND2_X1 U7628 ( .A1(n6360), .A2(n8795), .ZN(n8966) );
  INV_X1 U7629 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9725) );
  OR2_X1 U7630 ( .A1(n6261), .A2(n9725), .ZN(n6066) );
  NAND2_X1 U7631 ( .A1(n6098), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7632 ( .A1(n6100), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7633 ( .A1(n6101), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6063) );
  NAND4_X1 U7634 ( .A1(n6066), .A2(n6065), .A3(n6064), .A4(n6063), .ZN(n6572)
         );
  NAND2_X1 U7635 ( .A1(n6428), .A2(SI_0_), .ZN(n6068) );
  INV_X1 U7636 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U7637 ( .A1(n6068), .A2(n6067), .ZN(n6070) );
  AND2_X1 U7638 ( .A1(n6070), .A2(n6069), .ZN(n9495) );
  AND2_X1 U7639 ( .A1(n6572), .A2(n9694), .ZN(n9693) );
  NAND2_X1 U7640 ( .A1(n8966), .A2(n9693), .ZN(n9692) );
  NAND2_X1 U7641 ( .A1(n6576), .A2(n9700), .ZN(n6071) );
  NAND2_X1 U7642 ( .A1(n9692), .A2(n6071), .ZN(n6072) );
  NAND2_X1 U7643 ( .A1(n6100), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7644 ( .A1(n6098), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U7645 ( .A1(n6101), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6073) );
  INV_X1 U7646 ( .A(n6589), .ZN(n6710) );
  NAND2_X1 U7647 ( .A1(n6134), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6082) );
  NOR2_X1 U7648 ( .A1(n6077), .A2(n6121), .ZN(n6078) );
  MUX2_X1 U7649 ( .A(n6121), .B(n6078), .S(P1_IR_REG_2__SCAN_IN), .Z(n6081) );
  INV_X1 U7650 ( .A(n6079), .ZN(n6080) );
  NAND2_X1 U7651 ( .A1(n6589), .A2(n7862), .ZN(n6083) );
  NAND2_X1 U7652 ( .A1(n6097), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U7653 ( .A1(n6098), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6090) );
  INV_X1 U7654 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U7655 ( .A1(n6100), .A2(n6088), .ZN(n6089) );
  NAND2_X1 U7656 ( .A1(n6134), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U7657 ( .A1(n6079), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6093) );
  XNOR2_X1 U7658 ( .A(n6093), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9501) );
  NAND2_X1 U7659 ( .A1(n6243), .A2(n9501), .ZN(n6094) );
  NAND2_X1 U7660 ( .A1(n9734), .A2(n6707), .ZN(n8850) );
  INV_X1 U7661 ( .A(n6707), .ZN(n9742) );
  NAND2_X1 U7662 ( .A1(n9748), .A2(n9742), .ZN(n8799) );
  NAND2_X1 U7663 ( .A1(n8850), .A2(n8799), .ZN(n6709) );
  NAND2_X1 U7664 ( .A1(n9734), .A2(n9742), .ZN(n6096) );
  NAND2_X1 U7665 ( .A1(n4403), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7666 ( .A1(n6098), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6104) );
  INV_X1 U7667 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6099) );
  XNOR2_X1 U7668 ( .A(n6099), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n6610) );
  NAND2_X1 U7669 ( .A1(n6100), .A2(n6610), .ZN(n6103) );
  NAND2_X1 U7670 ( .A1(n6101), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6102) );
  INV_X1 U7671 ( .A(n9044), .ZN(n6942) );
  NAND2_X1 U7672 ( .A1(n6134), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7673 ( .A1(n6106), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6107) );
  XNOR2_X1 U7674 ( .A(n6107), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U7675 ( .A1(n6243), .A2(n6487), .ZN(n6108) );
  OAI211_X2 U7676 ( .C1(n8772), .C2(n6443), .A(n6109), .B(n6108), .ZN(n6785)
         );
  NAND2_X1 U7677 ( .A1(n6942), .A2(n6785), .ZN(n8849) );
  INV_X1 U7678 ( .A(n6785), .ZN(n9751) );
  NAND2_X1 U7679 ( .A1(n9044), .A2(n9751), .ZN(n8971) );
  NAND2_X1 U7680 ( .A1(n8849), .A2(n8971), .ZN(n6777) );
  NAND2_X1 U7681 ( .A1(n6776), .A2(n6777), .ZN(n6111) );
  NAND2_X1 U7682 ( .A1(n6942), .A2(n9751), .ZN(n6110) );
  NAND2_X1 U7683 ( .A1(n6111), .A2(n6110), .ZN(n6934) );
  INV_X1 U7684 ( .A(n6934), .ZN(n6112) );
  NAND2_X1 U7685 ( .A1(n9768), .A2(n8845), .ZN(n6114) );
  OAI21_X1 U7686 ( .B1(n6115), .B2(P1_REG3_REG_6__SCAN_IN), .A(n6128), .ZN(
        n6992) );
  INV_X1 U7687 ( .A(n6992), .ZN(n6116) );
  NAND2_X1 U7688 ( .A1(n6374), .A2(n6116), .ZN(n6118) );
  NAND2_X1 U7689 ( .A1(n6248), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6117) );
  OR2_X1 U7690 ( .A1(n6441), .A2(n8772), .ZN(n6125) );
  NOR2_X1 U7691 ( .A1(n6119), .A2(n6121), .ZN(n6120) );
  MUX2_X1 U7692 ( .A(n6121), .B(n6120), .S(P1_IR_REG_6__SCAN_IN), .Z(n6123) );
  OR2_X1 U7693 ( .A1(n6123), .A2(n6012), .ZN(n9611) );
  INV_X1 U7694 ( .A(n9611), .ZN(n6495) );
  AOI22_X1 U7695 ( .A1(n6254), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6243), .B2(
        n6495), .ZN(n6124) );
  NAND2_X1 U7696 ( .A1(n6988), .A2(n9779), .ZN(n8976) );
  NAND2_X1 U7697 ( .A1(n7027), .A2(n6988), .ZN(n6126) );
  NAND2_X1 U7698 ( .A1(n6097), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6133) );
  NAND2_X1 U7699 ( .A1(n6248), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6132) );
  AND2_X1 U7700 ( .A1(n6128), .A2(n6127), .ZN(n6129) );
  NOR2_X1 U7701 ( .A1(n6144), .A2(n6129), .ZN(n7137) );
  NAND2_X1 U7702 ( .A1(n6374), .A2(n7137), .ZN(n6131) );
  NAND2_X1 U7703 ( .A1(n6313), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6130) );
  NAND4_X1 U7704 ( .A1(n6133), .A2(n6132), .A3(n6131), .A4(n6130), .ZN(n9793)
         );
  NAND2_X1 U7705 ( .A1(n6446), .A2(n8780), .ZN(n6137) );
  NAND2_X1 U7706 ( .A1(n6122), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6135) );
  XNOR2_X1 U7707 ( .A(n6135), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6518) );
  AOI22_X1 U7708 ( .A1(n6254), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6243), .B2(
        n6518), .ZN(n6136) );
  OR2_X1 U7709 ( .A1(n7188), .A2(n7124), .ZN(n8865) );
  NAND2_X1 U7710 ( .A1(n7124), .A2(n7188), .ZN(n8861) );
  NAND2_X1 U7711 ( .A1(n8865), .A2(n8861), .ZN(n7024) );
  OR2_X1 U7712 ( .A1(n7124), .A2(n9793), .ZN(n6138) );
  NAND2_X1 U7713 ( .A1(n6139), .A2(n6138), .ZN(n7090) );
  INV_X1 U7714 ( .A(n7090), .ZN(n6151) );
  NAND2_X1 U7715 ( .A1(n6451), .A2(n8780), .ZN(n6143) );
  NAND2_X1 U7716 ( .A1(n6140), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6141) );
  XNOR2_X1 U7717 ( .A(n6141), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6649) );
  AOI22_X1 U7718 ( .A1(n6254), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6243), .B2(
        n6649), .ZN(n6142) );
  NAND2_X1 U7719 ( .A1(n4403), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7720 ( .A1(n6248), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6148) );
  OR2_X1 U7721 ( .A1(n6144), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6145) );
  AND2_X1 U7722 ( .A1(n6158), .A2(n6145), .ZN(n7190) );
  NAND2_X1 U7723 ( .A1(n6374), .A2(n7190), .ZN(n6147) );
  NAND2_X1 U7724 ( .A1(n6313), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6146) );
  NAND4_X1 U7725 ( .A1(n6149), .A2(n6148), .A3(n6147), .A4(n6146), .ZN(n9778)
         );
  OR2_X1 U7726 ( .A1(n9796), .A2(n7300), .ZN(n8864) );
  NAND2_X1 U7727 ( .A1(n9796), .A2(n7300), .ZN(n8875) );
  NAND2_X1 U7728 ( .A1(n9796), .A2(n9778), .ZN(n6152) );
  NAND2_X1 U7729 ( .A1(n6455), .A2(n8780), .ZN(n6156) );
  NAND2_X1 U7730 ( .A1(n6023), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6154) );
  XNOR2_X1 U7731 ( .A(n6154), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6652) );
  AOI22_X1 U7732 ( .A1(n6254), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6243), .B2(
        n6652), .ZN(n6155) );
  NAND2_X1 U7733 ( .A1(n6156), .A2(n6155), .ZN(n7233) );
  NAND2_X1 U7734 ( .A1(n6097), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U7735 ( .A1(n6248), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U7736 ( .A1(n6158), .A2(n6157), .ZN(n6159) );
  AND2_X1 U7737 ( .A1(n6169), .A2(n6159), .ZN(n7302) );
  NAND2_X1 U7738 ( .A1(n6374), .A2(n7302), .ZN(n6161) );
  NAND2_X1 U7739 ( .A1(n6313), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6160) );
  NAND4_X1 U7740 ( .A1(n6163), .A2(n6162), .A3(n6161), .A4(n6160), .ZN(n9792)
         );
  OR2_X1 U7741 ( .A1(n7233), .A2(n9792), .ZN(n6164) );
  NAND2_X1 U7742 ( .A1(n6459), .A2(n8780), .ZN(n6168) );
  INV_X1 U7743 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n10055) );
  OR2_X1 U7744 ( .A1(n6165), .A2(n10055), .ZN(n6166) );
  NAND2_X1 U7745 ( .A1(n6165), .A2(n10055), .ZN(n6177) );
  AOI22_X1 U7746 ( .A1(n6254), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6243), .B2(
        n6646), .ZN(n6167) );
  NAND2_X1 U7747 ( .A1(n6248), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U7748 ( .A1(n4403), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7749 ( .A1(n6169), .A2(n7252), .ZN(n6170) );
  AND2_X1 U7750 ( .A1(n6182), .A2(n6170), .ZN(n7251) );
  NAND2_X1 U7751 ( .A1(n6374), .A2(n7251), .ZN(n6172) );
  NAND2_X1 U7752 ( .A1(n6313), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6171) );
  NAND4_X1 U7753 ( .A1(n6174), .A2(n6173), .A3(n6172), .A4(n6171), .ZN(n9043)
         );
  INV_X1 U7754 ( .A(n9043), .ZN(n7533) );
  NAND2_X1 U7755 ( .A1(n7392), .A2(n7533), .ZN(n8871) );
  NAND2_X1 U7756 ( .A1(n4427), .A2(n6175), .ZN(n7375) );
  OR2_X1 U7757 ( .A1(n7392), .A2(n9043), .ZN(n6176) );
  NAND2_X1 U7758 ( .A1(n7375), .A2(n6176), .ZN(n7476) );
  NAND2_X1 U7759 ( .A1(n6509), .A2(n8780), .ZN(n6180) );
  NAND2_X1 U7760 ( .A1(n6177), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6178) );
  XNOR2_X1 U7761 ( .A(n6178), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9645) );
  AOI22_X1 U7762 ( .A1(n6266), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9645), .B2(
        n6243), .ZN(n6179) );
  NAND2_X1 U7763 ( .A1(n6248), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U7764 ( .A1(n6097), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6187) );
  AND2_X1 U7765 ( .A1(n6182), .A2(n6181), .ZN(n6183) );
  NOR2_X1 U7766 ( .A1(n6184), .A2(n6183), .ZN(n7535) );
  NAND2_X1 U7767 ( .A1(n6374), .A2(n7535), .ZN(n6186) );
  NAND2_X1 U7768 ( .A1(n6313), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6185) );
  NAND4_X1 U7769 ( .A1(n6188), .A2(n6187), .A3(n6186), .A4(n6185), .ZN(n9042)
         );
  INV_X1 U7770 ( .A(n9042), .ZN(n7470) );
  OR2_X1 U7771 ( .A1(n9553), .A2(n7470), .ZN(n7459) );
  NAND2_X1 U7772 ( .A1(n9553), .A2(n7470), .ZN(n8872) );
  NAND2_X1 U7773 ( .A1(n7459), .A2(n8872), .ZN(n8986) );
  OR2_X1 U7774 ( .A1(n9553), .A2(n9042), .ZN(n6189) );
  INV_X1 U7775 ( .A(n9041), .ZN(n7551) );
  OR2_X1 U7776 ( .A1(n7618), .A2(n7551), .ZN(n8879) );
  NAND2_X1 U7777 ( .A1(n7618), .A2(n7551), .ZN(n8873) );
  NAND2_X1 U7778 ( .A1(n6538), .A2(n8780), .ZN(n6194) );
  NAND2_X1 U7779 ( .A1(n6190), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6191) );
  MUX2_X1 U7780 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6191), .S(
        P1_IR_REG_13__SCAN_IN), .Z(n6192) );
  AOI22_X1 U7781 ( .A1(n6266), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n9668), .B2(
        n6243), .ZN(n6193) );
  NAND2_X1 U7782 ( .A1(n6248), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6201) );
  NAND2_X1 U7783 ( .A1(n6097), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U7784 ( .A1(n6196), .A2(n6195), .ZN(n6197) );
  AND2_X1 U7785 ( .A1(n6209), .A2(n6197), .ZN(n7659) );
  NAND2_X1 U7786 ( .A1(n6374), .A2(n7659), .ZN(n6199) );
  NAND2_X1 U7787 ( .A1(n6313), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6198) );
  NAND4_X1 U7788 ( .A1(n6201), .A2(n6200), .A3(n6199), .A4(n6198), .ZN(n9040)
         );
  INV_X1 U7789 ( .A(n9040), .ZN(n7592) );
  NAND2_X1 U7790 ( .A1(n7671), .A2(n7592), .ZN(n6203) );
  AOI21_X1 U7791 ( .B1(n4951), .B2(n6203), .A(n6202), .ZN(n7685) );
  NAND2_X1 U7792 ( .A1(n6542), .A2(n8780), .ZN(n6208) );
  NAND2_X1 U7793 ( .A1(n6204), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6205) );
  MUX2_X1 U7794 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6205), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n6206) );
  AOI22_X1 U7795 ( .A1(n6243), .A2(n9677), .B1(n6254), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U7796 ( .A1(n6097), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6214) );
  NAND2_X1 U7797 ( .A1(n6313), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6213) );
  AND2_X1 U7798 ( .A1(n6209), .A2(n10232), .ZN(n6210) );
  NOR2_X1 U7799 ( .A1(n6220), .A2(n6210), .ZN(n7820) );
  NAND2_X1 U7800 ( .A1(n6374), .A2(n7820), .ZN(n6212) );
  NAND2_X1 U7801 ( .A1(n6248), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6211) );
  NAND4_X1 U7802 ( .A1(n6214), .A2(n6213), .A3(n6212), .A4(n6211), .ZN(n9432)
         );
  NAND2_X1 U7803 ( .A1(n7824), .A2(n8758), .ZN(n8891) );
  NAND2_X1 U7804 ( .A1(n8894), .A2(n8891), .ZN(n8964) );
  NAND2_X1 U7805 ( .A1(n7685), .A2(n8964), .ZN(n7684) );
  NAND2_X1 U7806 ( .A1(n7684), .A2(n6215), .ZN(n7772) );
  NAND2_X1 U7807 ( .A1(n6634), .A2(n8780), .ZN(n6219) );
  NAND2_X1 U7808 ( .A1(n6216), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6217) );
  XNOR2_X1 U7809 ( .A(n6217), .B(P1_IR_REG_15__SCAN_IN), .ZN(n7202) );
  AOI22_X1 U7810 ( .A1(n7202), .A2(n6243), .B1(n6266), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n6218) );
  INV_X1 U7811 ( .A(n8768), .ZN(n9484) );
  NAND2_X1 U7812 ( .A1(n6248), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6226) );
  NAND2_X1 U7813 ( .A1(n4403), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6225) );
  NOR2_X1 U7814 ( .A1(n6220), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6221) );
  OR2_X1 U7815 ( .A1(n6222), .A2(n6221), .ZN(n8764) );
  INV_X1 U7816 ( .A(n8764), .ZN(n7773) );
  NAND2_X1 U7817 ( .A1(n6374), .A2(n7773), .ZN(n6224) );
  NAND2_X1 U7818 ( .A1(n6313), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6223) );
  NAND4_X1 U7819 ( .A1(n6226), .A2(n6225), .A3(n6224), .A4(n6223), .ZN(n9540)
         );
  INV_X1 U7820 ( .A(n9540), .ZN(n9339) );
  NAND2_X1 U7821 ( .A1(n7772), .A2(n4994), .ZN(n6228) );
  OR2_X1 U7822 ( .A1(n9539), .A2(n9316), .ZN(n8902) );
  NAND2_X1 U7823 ( .A1(n9539), .A2(n9316), .ZN(n9312) );
  NAND2_X1 U7824 ( .A1(n6720), .A2(n8780), .ZN(n6232) );
  INV_X1 U7825 ( .A(n6344), .ZN(n6229) );
  NAND2_X1 U7826 ( .A1(n6229), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6230) );
  XNOR2_X1 U7827 ( .A(n6230), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9082) );
  AOI22_X1 U7828 ( .A1(n6266), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6243), .B2(
        n9082), .ZN(n6231) );
  NAND2_X1 U7829 ( .A1(n6233), .A2(n8699), .ZN(n6234) );
  NAND2_X1 U7830 ( .A1(n6235), .A2(n6234), .ZN(n9322) );
  NAND2_X1 U7831 ( .A1(n4403), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U7832 ( .A1(n6248), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6236) );
  AND2_X1 U7833 ( .A1(n6237), .A2(n6236), .ZN(n6239) );
  NAND2_X1 U7834 ( .A1(n6313), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6238) );
  OAI211_X1 U7835 ( .C1(n9322), .C2(n6264), .A(n6239), .B(n6238), .ZN(n9541)
         );
  NAND2_X1 U7836 ( .A1(n9428), .A2(n9541), .ZN(n6240) );
  INV_X1 U7837 ( .A(n9428), .ZN(n9327) );
  INV_X1 U7838 ( .A(n9541), .ZN(n8693) );
  OR2_X1 U7839 ( .A1(n9421), .A2(n9317), .ZN(n8912) );
  NAND2_X1 U7840 ( .A1(n9421), .A2(n9317), .ZN(n8906) );
  NAND2_X1 U7841 ( .A1(n8912), .A2(n8906), .ZN(n9297) );
  NAND2_X1 U7842 ( .A1(n9298), .A2(n9297), .ZN(n9299) );
  NAND2_X1 U7843 ( .A1(n7044), .A2(n8780), .ZN(n6245) );
  XNOR2_X1 U7844 ( .A(n6242), .B(n6341), .ZN(n6561) );
  AOI22_X1 U7845 ( .A1(n9704), .A2(n6243), .B1(n6266), .B2(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n6244) );
  NOR2_X1 U7846 ( .A1(n6246), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6247) );
  OR2_X1 U7847 ( .A1(n6257), .A2(n6247), .ZN(n9278) );
  INV_X1 U7848 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9418) );
  NAND2_X1 U7849 ( .A1(n4403), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6250) );
  NAND2_X1 U7850 ( .A1(n6313), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6249) );
  OAI211_X1 U7851 ( .C1(n9418), .C2(n6086), .A(n6250), .B(n6249), .ZN(n6251)
         );
  INV_X1 U7852 ( .A(n6251), .ZN(n6252) );
  OAI21_X1 U7853 ( .B1(n9278), .B2(n6264), .A(n6252), .ZN(n9295) );
  INV_X1 U7854 ( .A(n9295), .ZN(n8736) );
  NAND2_X1 U7855 ( .A1(n4702), .A2(n8736), .ZN(n6253) );
  AOI22_X2 U7856 ( .A1(n9277), .A2(n6253), .B1(n9295), .B2(n9289), .ZN(n9256)
         );
  NAND2_X1 U7857 ( .A1(n7214), .A2(n8780), .ZN(n6256) );
  NAND2_X1 U7858 ( .A1(n6254), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6255) );
  NOR2_X1 U7859 ( .A1(n6257), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6258) );
  OR2_X1 U7860 ( .A1(n6269), .A2(n6258), .ZN(n9266) );
  INV_X1 U7861 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10136) );
  NAND2_X1 U7862 ( .A1(n6248), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6260) );
  NAND2_X1 U7863 ( .A1(n6313), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6259) );
  OAI211_X1 U7864 ( .C1(n6261), .C2(n10136), .A(n6260), .B(n6259), .ZN(n6262)
         );
  INV_X1 U7865 ( .A(n6262), .ZN(n6263) );
  OAI21_X1 U7866 ( .B1(n9266), .B2(n6264), .A(n6263), .ZN(n9412) );
  NAND2_X1 U7867 ( .A1(n9265), .A2(n9412), .ZN(n6265) );
  INV_X1 U7868 ( .A(n9412), .ZN(n9284) );
  NAND2_X1 U7869 ( .A1(n7213), .A2(n8780), .ZN(n6268) );
  NAND2_X1 U7870 ( .A1(n6266), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6267) );
  OR2_X1 U7871 ( .A1(n6269), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6270) );
  AND2_X1 U7872 ( .A1(n6270), .A2(n6279), .ZN(n9250) );
  NAND2_X1 U7873 ( .A1(n9250), .A2(n6374), .ZN(n6275) );
  INV_X1 U7874 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9404) );
  NAND2_X1 U7875 ( .A1(n6097), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6272) );
  NAND2_X1 U7876 ( .A1(n6313), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6271) );
  OAI211_X1 U7877 ( .C1(n6086), .C2(n9404), .A(n6272), .B(n6271), .ZN(n6273)
         );
  INV_X1 U7878 ( .A(n6273), .ZN(n6274) );
  NAND2_X1 U7879 ( .A1(n6275), .A2(n6274), .ZN(n9260) );
  NAND2_X1 U7880 ( .A1(n9249), .A2(n7932), .ZN(n8917) );
  NAND2_X1 U7881 ( .A1(n9224), .A2(n8917), .ZN(n9239) );
  NAND2_X1 U7882 ( .A1(n7403), .A2(n8780), .ZN(n6277) );
  NAND2_X1 U7883 ( .A1(n6266), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6276) );
  NAND2_X1 U7884 ( .A1(n6248), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6284) );
  NAND2_X1 U7885 ( .A1(n6097), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6283) );
  INV_X1 U7886 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6280) );
  AOI21_X1 U7887 ( .B1(n6280), .B2(n6279), .A(n6278), .ZN(n9232) );
  NAND2_X1 U7888 ( .A1(n6374), .A2(n9232), .ZN(n6282) );
  NAND2_X1 U7889 ( .A1(n6313), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6281) );
  NAND2_X1 U7890 ( .A1(n7539), .A2(n8780), .ZN(n6287) );
  NAND2_X1 U7891 ( .A1(n6266), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6286) );
  NAND2_X1 U7892 ( .A1(n4403), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6294) );
  NAND2_X1 U7893 ( .A1(n6313), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6293) );
  INV_X1 U7894 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n10223) );
  NAND2_X1 U7895 ( .A1(n10223), .A2(n6288), .ZN(n6290) );
  AND2_X1 U7896 ( .A1(n6290), .A2(n6289), .ZN(n9214) );
  NAND2_X1 U7897 ( .A1(n6374), .A2(n9214), .ZN(n6292) );
  NAND2_X1 U7898 ( .A1(n6248), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6291) );
  NAND4_X1 U7899 ( .A1(n6294), .A2(n6293), .A3(n6292), .A4(n6291), .ZN(n9228)
         );
  NAND2_X1 U7900 ( .A1(n9464), .A2(n9196), .ZN(n6296) );
  AOI21_X2 U7901 ( .B1(n9207), .B2(n6296), .A(n6295), .ZN(n9192) );
  NAND2_X1 U7902 ( .A1(n7681), .A2(n8780), .ZN(n6299) );
  NAND2_X1 U7903 ( .A1(n6266), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6298) );
  NAND2_X1 U7904 ( .A1(n6248), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U7905 ( .A1(n4403), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6305) );
  INV_X1 U7906 ( .A(n6301), .ZN(n6300) );
  NAND2_X1 U7907 ( .A1(n6300), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6311) );
  INV_X1 U7908 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n10196) );
  NAND2_X1 U7909 ( .A1(n6301), .A2(n10196), .ZN(n6302) );
  AND2_X1 U7910 ( .A1(n6311), .A2(n6302), .ZN(n9186) );
  NAND2_X1 U7911 ( .A1(n6374), .A2(n9186), .ZN(n6304) );
  NAND2_X1 U7912 ( .A1(n6313), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6303) );
  NAND4_X1 U7913 ( .A1(n6306), .A2(n6305), .A3(n6304), .A4(n6303), .ZN(n9161)
         );
  NAND2_X1 U7914 ( .A1(n9185), .A2(n9197), .ZN(n8932) );
  NAND2_X1 U7915 ( .A1(n9175), .A2(n8932), .ZN(n9173) );
  NAND2_X1 U7916 ( .A1(n7700), .A2(n8780), .ZN(n6308) );
  NAND2_X1 U7917 ( .A1(n6266), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6307) );
  NAND2_X1 U7918 ( .A1(n6087), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6317) );
  NAND2_X1 U7919 ( .A1(n6097), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6316) );
  INV_X1 U7920 ( .A(n6311), .ZN(n6309) );
  NAND2_X1 U7921 ( .A1(n6309), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6320) );
  INV_X1 U7922 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6310) );
  NAND2_X1 U7923 ( .A1(n6311), .A2(n6310), .ZN(n6312) );
  AND2_X1 U7924 ( .A1(n6320), .A2(n6312), .ZN(n9167) );
  NAND2_X1 U7925 ( .A1(n6374), .A2(n9167), .ZN(n6315) );
  NAND2_X1 U7926 ( .A1(n6313), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6314) );
  NAND4_X1 U7927 ( .A1(n6317), .A2(n6316), .A3(n6315), .A4(n6314), .ZN(n9180)
         );
  AND2_X1 U7928 ( .A1(n9166), .A2(n9180), .ZN(n8838) );
  NAND2_X1 U7929 ( .A1(n7743), .A2(n8780), .ZN(n6319) );
  NAND2_X1 U7930 ( .A1(n6266), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6318) );
  NAND2_X1 U7931 ( .A1(n4403), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6325) );
  NAND2_X1 U7932 ( .A1(n6313), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6324) );
  INV_X1 U7933 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9977) );
  NAND2_X1 U7934 ( .A1(n6320), .A2(n9977), .ZN(n6321) );
  NAND2_X1 U7935 ( .A1(n6374), .A2(n9144), .ZN(n6323) );
  NAND2_X1 U7936 ( .A1(n6087), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6322) );
  NAND4_X1 U7937 ( .A1(n6325), .A2(n6324), .A3(n6323), .A4(n6322), .ZN(n9160)
         );
  NAND2_X1 U7938 ( .A1(n9370), .A2(n7875), .ZN(n8835) );
  NOR2_X1 U7939 ( .A1(n9370), .A2(n9160), .ZN(n6326) );
  NAND2_X1 U7940 ( .A1(n7885), .A2(n8780), .ZN(n6328) );
  NAND2_X1 U7941 ( .A1(n6266), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6327) );
  NAND2_X1 U7942 ( .A1(n6248), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U7943 ( .A1(n6097), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6335) );
  INV_X1 U7944 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6329) );
  NAND2_X1 U7945 ( .A1(n6330), .A2(n6329), .ZN(n6331) );
  NAND2_X1 U7946 ( .A1(n6373), .A2(n6331), .ZN(n8001) );
  INV_X1 U7947 ( .A(n8001), .ZN(n6332) );
  NAND2_X1 U7948 ( .A1(n6374), .A2(n6332), .ZN(n6334) );
  NAND2_X1 U7949 ( .A1(n6313), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6333) );
  NAND4_X1 U7950 ( .A1(n6336), .A2(n6335), .A3(n6334), .A4(n6333), .ZN(n9039)
         );
  OR2_X1 U7951 ( .A1(n8006), .A2(n9362), .ZN(n8939) );
  NAND2_X1 U7952 ( .A1(n8006), .A2(n9362), .ZN(n9132) );
  NAND2_X1 U7953 ( .A1(n6337), .A2(n8998), .ZN(n9122) );
  INV_X1 U7954 ( .A(n6337), .ZN(n6339) );
  NAND2_X1 U7955 ( .A1(n6339), .A2(n6338), .ZN(n6340) );
  INV_X1 U7956 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6343) );
  NAND2_X1 U7957 ( .A1(n6344), .A2(n4993), .ZN(n6345) );
  INV_X1 U7958 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6346) );
  NAND2_X1 U7959 ( .A1(n9215), .A2(n6348), .ZN(n9028) );
  NAND2_X1 U7960 ( .A1(n6350), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6349) );
  MUX2_X1 U7961 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6349), .S(
        P1_IR_REG_22__SCAN_IN), .Z(n6352) );
  NAND2_X1 U7962 ( .A1(n6352), .A2(n6390), .ZN(n7407) );
  NAND2_X1 U7963 ( .A1(n6353), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6354) );
  MUX2_X1 U7964 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6354), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n6355) );
  NAND2_X1 U7965 ( .A1(n9034), .A2(n9021), .ZN(n6597) );
  OR2_X1 U7966 ( .A1(n9028), .A2(n6597), .ZN(n6774) );
  NAND2_X2 U7967 ( .A1(n6356), .A2(n9021), .ZN(n6562) );
  NAND2_X1 U7968 ( .A1(n6562), .A2(n7407), .ZN(n6357) );
  AND2_X1 U7969 ( .A1(n6357), .A2(n9215), .ZN(n6358) );
  NAND2_X1 U7970 ( .A1(n6774), .A2(n6358), .ZN(n9712) );
  INV_X1 U7971 ( .A(n6348), .ZN(n9025) );
  INV_X1 U7972 ( .A(n6572), .ZN(n6359) );
  NAND2_X1 U7973 ( .A1(n6359), .A2(n9694), .ZN(n9708) );
  NAND2_X1 U7974 ( .A1(n9708), .A2(n6360), .ZN(n6361) );
  NAND2_X1 U7975 ( .A1(n6361), .A2(n8795), .ZN(n6994) );
  OR2_X1 U7976 ( .A1(n6084), .A2(n6994), .ZN(n6363) );
  NAND2_X1 U7977 ( .A1(n6710), .A2(n7862), .ZN(n6362) );
  NAND2_X1 U7978 ( .A1(n6363), .A2(n6362), .ZN(n9006) );
  NAND2_X1 U7979 ( .A1(n9006), .A2(n8799), .ZN(n8852) );
  NAND2_X1 U7980 ( .A1(n8852), .A2(n8850), .ZN(n8843) );
  INV_X1 U7981 ( .A(n6777), .ZN(n6775) );
  NAND2_X1 U7982 ( .A1(n8843), .A2(n6775), .ZN(n6364) );
  INV_X1 U7983 ( .A(n6893), .ZN(n8857) );
  INV_X1 U7984 ( .A(n7024), .ZN(n8981) );
  NAND2_X1 U7985 ( .A1(n7086), .A2(n8864), .ZN(n7161) );
  INV_X1 U7986 ( .A(n9792), .ZN(n7393) );
  OR2_X1 U7987 ( .A1(n7233), .A2(n7393), .ZN(n8868) );
  NAND2_X1 U7988 ( .A1(n7233), .A2(n7393), .ZN(n8867) );
  NAND2_X1 U7989 ( .A1(n7161), .A2(n8983), .ZN(n7160) );
  NAND2_X1 U7990 ( .A1(n7160), .A2(n8868), .ZN(n7378) );
  NAND2_X1 U7991 ( .A1(n7378), .A2(n7377), .ZN(n7376) );
  AND2_X1 U7992 ( .A1(n8879), .A2(n7459), .ZN(n8888) );
  OR2_X1 U7993 ( .A1(n7645), .A2(n7592), .ZN(n8804) );
  NAND2_X1 U7994 ( .A1(n7645), .A2(n7592), .ZN(n8890) );
  NAND2_X1 U7995 ( .A1(n7546), .A2(n8990), .ZN(n7686) );
  INV_X1 U7996 ( .A(n8890), .ZN(n6365) );
  NOR2_X1 U7997 ( .A1(n8964), .A2(n6365), .ZN(n6366) );
  OR2_X1 U7998 ( .A1(n8768), .A2(n9339), .ZN(n8803) );
  NAND2_X1 U7999 ( .A1(n8768), .A2(n9339), .ZN(n8896) );
  INV_X1 U8000 ( .A(n9331), .ZN(n8993) );
  NAND2_X1 U8001 ( .A1(n9428), .A2(n8693), .ZN(n8905) );
  AND2_X1 U8002 ( .A1(n8905), .A2(n9312), .ZN(n8788) );
  OR2_X1 U8003 ( .A1(n9428), .A2(n8693), .ZN(n9292) );
  AND2_X1 U8004 ( .A1(n8912), .A2(n9292), .ZN(n8907) );
  NAND2_X1 U8005 ( .A1(n6367), .A2(n8906), .ZN(n9274) );
  OR2_X1 U8006 ( .A1(n9289), .A2(n8736), .ZN(n8911) );
  NAND2_X1 U8007 ( .A1(n9289), .A2(n8736), .ZN(n8914) );
  AND2_X1 U8008 ( .A1(n9265), .A2(n9284), .ZN(n8913) );
  OR2_X1 U8009 ( .A1(n9265), .A2(n9284), .ZN(n8962) );
  INV_X1 U8010 ( .A(n9239), .ZN(n9244) );
  NAND2_X1 U8011 ( .A1(n9467), .A2(n9389), .ZN(n8960) );
  AND2_X1 U8012 ( .A1(n8960), .A2(n9224), .ZN(n8918) );
  OR2_X1 U8013 ( .A1(n9220), .A2(n9196), .ZN(n8959) );
  NAND2_X1 U8014 ( .A1(n9220), .A2(n9196), .ZN(n8958) );
  AND2_X1 U8015 ( .A1(n9199), .A2(n8659), .ZN(n8841) );
  OR2_X1 U8016 ( .A1(n9199), .A2(n8659), .ZN(n8956) );
  NAND2_X1 U8017 ( .A1(n6369), .A2(n8956), .ZN(n9178) );
  INV_X1 U8018 ( .A(n9180), .ZN(n9148) );
  OR2_X1 U8019 ( .A1(n9166), .A2(n9148), .ZN(n8836) );
  NAND2_X1 U8020 ( .A1(n8836), .A2(n9175), .ZN(n8825) );
  NAND2_X1 U8021 ( .A1(n9166), .A2(n9148), .ZN(n8837) );
  INV_X1 U8022 ( .A(n9010), .ZN(n8827) );
  OAI21_X1 U8023 ( .B1(n6370), .B2(n6338), .A(n9133), .ZN(n7882) );
  OR2_X1 U8024 ( .A1(n9215), .A2(n7407), .ZN(n8955) );
  OR2_X1 U8025 ( .A1(n6348), .A2(n8954), .ZN(n6371) );
  NOR2_X1 U8026 ( .A1(n9700), .A2(n9694), .ZN(n9697) );
  NAND2_X1 U8027 ( .A1(n9697), .A2(n9732), .ZN(n6998) );
  OR2_X1 U8028 ( .A1(n6998), .A2(n6707), .ZN(n6780) );
  INV_X1 U8029 ( .A(n7392), .ZN(n7385) );
  INV_X1 U8030 ( .A(n7824), .ZN(n7789) );
  NAND2_X1 U8031 ( .A1(n7692), .A2(n7789), .ZN(n7776) );
  AOI211_X1 U8032 ( .C1(n8006), .C2(n9142), .A(n9319), .B(n9124), .ZN(n7873)
         );
  OR2_X1 U8033 ( .A1(n6372), .A2(n6597), .ZN(n9361) );
  NAND2_X1 U8034 ( .A1(n4403), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6378) );
  NAND2_X1 U8035 ( .A1(n6313), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6377) );
  INV_X1 U8036 ( .A(n6373), .ZN(n9128) );
  NAND2_X1 U8037 ( .A1(n6374), .A2(n9128), .ZN(n6376) );
  NAND2_X1 U8038 ( .A1(n6087), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6375) );
  NAND4_X1 U8039 ( .A1(n6378), .A2(n6377), .A3(n6376), .A4(n6375), .ZN(n9038)
         );
  INV_X1 U8040 ( .A(n9038), .ZN(n8942) );
  INV_X1 U8041 ( .A(n6597), .ZN(n6394) );
  OAI22_X1 U8042 ( .A1(n7875), .A2(n9361), .B1(n8942), .B2(n9733), .ZN(n6379)
         );
  AOI211_X1 U8043 ( .C1(n7882), .C2(n9706), .A(n7873), .B(n6379), .ZN(n6380)
         );
  OAI21_X1 U8044 ( .B1(n7884), .B2(n9759), .A(n6380), .ZN(n6420) );
  NAND2_X1 U8045 ( .A1(n6390), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6392) );
  XNOR2_X1 U8046 ( .A(n6392), .B(n6391), .ZN(n7543) );
  AND2_X1 U8047 ( .A1(n7543), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6393) );
  NAND2_X1 U8048 ( .A1(n9028), .A2(n6394), .ZN(n6545) );
  NAND2_X1 U8049 ( .A1(n7748), .A2(P1_B_REG_SCAN_IN), .ZN(n6396) );
  INV_X1 U8050 ( .A(n7600), .ZN(n6395) );
  MUX2_X1 U8051 ( .A(n6396), .B(P1_B_REG_SCAN_IN), .S(n6395), .Z(n6398) );
  NOR4_X1 U8052 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6402) );
  NOR4_X1 U8053 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6401) );
  NOR4_X1 U8054 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n6400) );
  NOR4_X1 U8055 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n6399) );
  NAND4_X1 U8056 ( .A1(n6402), .A2(n6401), .A3(n6400), .A4(n6399), .ZN(n6407)
         );
  NOR2_X1 U8057 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .ZN(
        n10246) );
  NOR4_X1 U8058 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n6405) );
  NOR4_X1 U8059 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6404) );
  NOR4_X1 U8060 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n6403) );
  NAND4_X1 U8061 ( .A1(n10246), .A2(n6405), .A3(n6404), .A4(n6403), .ZN(n6406)
         );
  NOR2_X1 U8062 ( .A1(n6407), .A2(n6406), .ZN(n6408) );
  NOR2_X1 U8063 ( .A1(n9718), .A2(n6408), .ZN(n6546) );
  INV_X1 U8064 ( .A(n6546), .ZN(n6412) );
  NAND2_X1 U8065 ( .A1(n6409), .A2(n7748), .ZN(n6410) );
  OAI21_X1 U8066 ( .B1(n9718), .B2(P1_D_REG_1__SCAN_IN), .A(n6410), .ZN(n6547)
         );
  INV_X1 U8067 ( .A(n6554), .ZN(n6411) );
  NAND4_X1 U8068 ( .A1(n6690), .A2(n6412), .A3(n6547), .A4(n6411), .ZN(n6419)
         );
  INV_X1 U8069 ( .A(n9718), .ZN(n6414) );
  INV_X1 U8070 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U8071 ( .A1(n6414), .A2(n6413), .ZN(n6416) );
  NAND2_X1 U8072 ( .A1(n6409), .A2(n7600), .ZN(n6415) );
  INV_X1 U8073 ( .A(n6417), .ZN(n6418) );
  INV_X1 U8074 ( .A(n6421), .ZN(n6422) );
  NAND2_X1 U8075 ( .A1(n6558), .A2(n6597), .ZN(n6423) );
  NAND2_X1 U8076 ( .A1(n6423), .A2(n7543), .ZN(n6500) );
  NAND2_X1 U8077 ( .A1(n6500), .A2(n6498), .ZN(n6424) );
  NAND2_X1 U8078 ( .A1(n6424), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8079 ( .A(n6425), .ZN(n6724) );
  INV_X1 U8080 ( .A(n7543), .ZN(n6426) );
  NOR2_X1 U8081 ( .A1(n6558), .A2(n6426), .ZN(n6501) );
  INV_X1 U8082 ( .A(n9501), .ZN(n6474) );
  NOR2_X1 U8083 ( .A1(n6428), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9488) );
  INV_X1 U8084 ( .A(n9488), .ZN(n9491) );
  OAI222_X1 U8085 ( .A1(n6474), .A2(P1_U3084), .B1(n9494), .B2(n6430), .C1(
        n6427), .C2(n9491), .ZN(P1_U3350) );
  INV_X1 U8086 ( .A(n6487), .ZN(n9575) );
  OAI222_X1 U8087 ( .A1(n9575), .A2(P1_U3084), .B1(n9494), .B2(n6443), .C1(
        n10262), .C2(n9491), .ZN(P1_U3349) );
  OAI222_X1 U8088 ( .A1(n8130), .A2(n6790), .B1(n8025), .B2(n6430), .C1(n6429), 
        .C2(n8651), .ZN(P2_U3355) );
  OAI222_X1 U8089 ( .A1(P2_U3152), .A2(n8192), .B1(n8025), .B2(n6434), .C1(
        n6431), .C2(n8651), .ZN(P2_U3356) );
  OAI222_X1 U8090 ( .A1(P2_U3152), .A2(n6735), .B1(n8025), .B2(n6436), .C1(
        n6432), .C2(n8651), .ZN(P2_U3357) );
  INV_X1 U8091 ( .A(n9060), .ZN(n6471) );
  OAI222_X1 U8092 ( .A1(n6471), .A2(P1_U3084), .B1(n9494), .B2(n6434), .C1(
        n6433), .C2(n9491), .ZN(P1_U3351) );
  INV_X1 U8093 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6435) );
  OAI222_X1 U8094 ( .A1(n6060), .A2(P1_U3084), .B1(n9494), .B2(n6436), .C1(
        n6435), .C2(n9491), .ZN(P1_U3352) );
  OAI222_X1 U8095 ( .A1(n9594), .A2(P1_U3084), .B1(n9494), .B2(n6438), .C1(
        n6437), .C2(n9491), .ZN(P1_U3348) );
  OAI222_X1 U8096 ( .A1(n9611), .A2(P1_U3084), .B1(n9494), .B2(n6441), .C1(
        n6440), .C2(n9491), .ZN(P1_U3347) );
  NAND2_X1 U8097 ( .A1(n9485), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6445) );
  OAI21_X1 U8098 ( .B1(n6547), .B2(n9485), .A(n6445), .ZN(P1_U3441) );
  INV_X1 U8099 ( .A(n6518), .ZN(n6467) );
  INV_X1 U8100 ( .A(n6446), .ZN(n6449) );
  INV_X1 U8101 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6447) );
  OAI222_X1 U8102 ( .A1(n6467), .A2(P1_U3084), .B1(n9494), .B2(n6449), .C1(
        n6447), .C2(n9491), .ZN(P1_U3346) );
  INV_X1 U8103 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6450) );
  INV_X1 U8104 ( .A(n6451), .ZN(n6454) );
  INV_X1 U8105 ( .A(n8651), .ZN(n7541) );
  AOI22_X1 U8106 ( .A1(n6873), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n7541), .ZN(n6452) );
  OAI21_X1 U8107 ( .B1(n6454), .B2(n8025), .A(n6452), .ZN(P2_U3350) );
  INV_X1 U8108 ( .A(n6649), .ZN(n6504) );
  OAI222_X1 U8109 ( .A1(n6504), .A2(P1_U3084), .B1(n9494), .B2(n6454), .C1(
        n6453), .C2(n9491), .ZN(P1_U3345) );
  INV_X1 U8110 ( .A(n6455), .ZN(n6458) );
  INV_X1 U8111 ( .A(n6652), .ZN(n9622) );
  OAI222_X1 U8112 ( .A1(P1_U3084), .A2(n9622), .B1(n9494), .B2(n6458), .C1(
        n6457), .C2(n9491), .ZN(P1_U3344) );
  INV_X1 U8113 ( .A(n6459), .ZN(n6462) );
  AOI22_X1 U8114 ( .A1(n7076), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n7541), .ZN(n6460) );
  OAI21_X1 U8115 ( .B1(n6462), .B2(n8025), .A(n6460), .ZN(P2_U3348) );
  INV_X1 U8116 ( .A(n6646), .ZN(n9633) );
  OAI222_X1 U8117 ( .A1(P1_U3084), .A2(n9633), .B1(n9494), .B2(n6462), .C1(
        n6461), .C2(n9491), .ZN(P1_U3343) );
  NAND2_X1 U8118 ( .A1(n6087), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6465) );
  NAND2_X1 U8119 ( .A1(n6313), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U8120 ( .A1(n6097), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6463) );
  INV_X1 U8121 ( .A(n9113), .ZN(n8833) );
  NAND2_X1 U8122 ( .A1(P1_U4006), .A2(n8833), .ZN(n6466) );
  OAI21_X1 U8123 ( .B1(P1_U4006), .B2(n7847), .A(n6466), .ZN(P1_U3586) );
  NOR2_X1 U8124 ( .A1(n6518), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6479) );
  INV_X1 U8125 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6468) );
  AOI22_X1 U8126 ( .A1(n6518), .A2(n6468), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n6467), .ZN(n6514) );
  INV_X1 U8127 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10013) );
  INV_X1 U8128 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9980) );
  NAND2_X1 U8129 ( .A1(n9501), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6476) );
  XNOR2_X1 U8130 ( .A(n9060), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n9053) );
  INV_X1 U8131 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6469) );
  MUX2_X1 U8132 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6469), .S(n6490), .Z(n9569)
         );
  AND2_X1 U8133 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9570) );
  NAND2_X1 U8134 ( .A1(n9569), .A2(n9570), .ZN(n9568) );
  NAND2_X1 U8135 ( .A1(n6490), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6470) );
  NAND2_X1 U8136 ( .A1(n9568), .A2(n6470), .ZN(n9052) );
  INV_X1 U8137 ( .A(n9052), .ZN(n6472) );
  INV_X1 U8138 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10250) );
  OAI22_X1 U8139 ( .A1(n9053), .A2(n6472), .B1(n6471), .B2(n10250), .ZN(n9503)
         );
  INV_X1 U8140 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6475) );
  INV_X1 U8141 ( .A(n6476), .ZN(n6473) );
  AOI21_X1 U8142 ( .B1(n6475), .B2(n6474), .A(n6473), .ZN(n9504) );
  NAND2_X1 U8143 ( .A1(n9503), .A2(n9504), .ZN(n9502) );
  NAND2_X1 U8144 ( .A1(n6476), .A2(n9502), .ZN(n9579) );
  INV_X1 U8145 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6477) );
  AOI22_X1 U8146 ( .A1(n6487), .A2(n6477), .B1(P1_REG2_REG_4__SCAN_IN), .B2(
        n9575), .ZN(n9578) );
  NOR2_X1 U8147 ( .A1(n9579), .A2(n9578), .ZN(n9577) );
  NOR2_X1 U8148 ( .A1(n6487), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6478) );
  MUX2_X1 U8149 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9980), .S(n9594), .Z(n9597)
         );
  NOR2_X1 U8150 ( .A1(n9598), .A2(n9597), .ZN(n9596) );
  AOI21_X1 U8151 ( .B1(n9594), .B2(n9980), .A(n9596), .ZN(n9615) );
  MUX2_X1 U8152 ( .A(n10013), .B(P1_REG2_REG_6__SCAN_IN), .S(n9611), .Z(n9614)
         );
  NAND2_X1 U8153 ( .A1(n9615), .A2(n9614), .ZN(n9613) );
  OAI21_X1 U8154 ( .B1(n9611), .B2(n10013), .A(n9613), .ZN(n6513) );
  NOR2_X1 U8155 ( .A1(n6514), .A2(n6513), .ZN(n6512) );
  INV_X1 U8156 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6480) );
  AOI22_X1 U8157 ( .A1(n6649), .A2(n6480), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n6504), .ZN(n6481) );
  NOR2_X1 U8158 ( .A1(n6482), .A2(n6481), .ZN(n6650) );
  AOI21_X1 U8159 ( .B1(n6482), .B2(n6481), .A(n6650), .ZN(n6508) );
  NOR2_X1 U8160 ( .A1(n9047), .A2(P1_U3084), .ZN(n7744) );
  INV_X1 U8161 ( .A(n6372), .ZN(n9049) );
  NAND2_X1 U8162 ( .A1(n9100), .A2(n9049), .ZN(n9600) );
  INV_X1 U8163 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9824) );
  AOI22_X1 U8164 ( .A1(n6649), .A2(P1_REG1_REG_8__SCAN_IN), .B1(n9824), .B2(
        n6504), .ZN(n6497) );
  NOR2_X1 U8165 ( .A1(n6518), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6483) );
  AOI21_X1 U8166 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n6518), .A(n6483), .ZN(
        n6517) );
  NOR2_X1 U8167 ( .A1(P1_REG1_REG_6__SCAN_IN), .A2(n6495), .ZN(n6484) );
  AOI21_X1 U8168 ( .B1(n6495), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6484), .ZN(
        n9606) );
  INV_X1 U8169 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6485) );
  OR2_X1 U8170 ( .A1(n9594), .A2(n6485), .ZN(n6494) );
  MUX2_X1 U8171 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6485), .S(n9594), .Z(n9589)
         );
  OR2_X1 U8172 ( .A1(n6487), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6492) );
  NOR2_X1 U8173 ( .A1(n6487), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6486) );
  AOI21_X1 U8174 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n6487), .A(n6486), .ZN(
        n9574) );
  INV_X1 U8175 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6488) );
  MUX2_X1 U8176 ( .A(n6488), .B(P1_REG1_REG_1__SCAN_IN), .S(n6490), .Z(n9564)
         );
  INV_X1 U8177 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9810) );
  INV_X1 U8178 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6489) );
  NOR3_X1 U8179 ( .A1(n9564), .A2(n9810), .A3(n6489), .ZN(n9563) );
  AOI21_X1 U8180 ( .B1(n6490), .B2(P1_REG1_REG_1__SCAN_IN), .A(n9563), .ZN(
        n9056) );
  XNOR2_X1 U8181 ( .A(n9060), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9055) );
  NOR2_X1 U8182 ( .A1(n9056), .A2(n9055), .ZN(n9054) );
  AOI21_X1 U8183 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(n9060), .A(n9054), .ZN(
        n9498) );
  XNOR2_X1 U8184 ( .A(n9501), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9497) );
  NOR2_X1 U8185 ( .A1(n9498), .A2(n9497), .ZN(n9496) );
  AOI21_X1 U8186 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n9501), .A(n9496), .ZN(
        n9573) );
  NAND2_X1 U8187 ( .A1(n9574), .A2(n9573), .ZN(n6491) );
  NAND2_X1 U8188 ( .A1(n6492), .A2(n6491), .ZN(n9588) );
  NOR2_X1 U8189 ( .A1(n9589), .A2(n9588), .ZN(n9587) );
  INV_X1 U8190 ( .A(n9587), .ZN(n6493) );
  AND2_X1 U8191 ( .A1(n6494), .A2(n6493), .ZN(n9605) );
  NAND2_X1 U8192 ( .A1(n9606), .A2(n9605), .ZN(n9604) );
  OAI21_X1 U8193 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n6495), .A(n9604), .ZN(
        n6516) );
  NAND2_X1 U8194 ( .A1(n6517), .A2(n6516), .ZN(n6515) );
  OAI21_X1 U8195 ( .B1(n6518), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6515), .ZN(
        n6496) );
  NAND2_X1 U8196 ( .A1(n6497), .A2(n6496), .ZN(n6638) );
  OAI21_X1 U8197 ( .B1(n6497), .B2(n6496), .A(n6638), .ZN(n6506) );
  AND2_X1 U8198 ( .A1(n6498), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6499) );
  AND2_X1 U8199 ( .A1(n6500), .A2(n6499), .ZN(n9561) );
  NAND2_X1 U8200 ( .A1(n9100), .A2(n6372), .ZN(n9634) );
  INV_X1 U8201 ( .A(n9691), .ZN(n9649) );
  NAND2_X1 U8202 ( .A1(n9649), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n6503) );
  INV_X1 U8203 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6502) );
  OR2_X1 U8204 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6502), .ZN(n7186) );
  OAI211_X1 U8205 ( .C1(n6504), .C2(n9634), .A(n6503), .B(n7186), .ZN(n6505)
         );
  AOI21_X1 U8206 ( .B1(n6506), .B2(n9686), .A(n6505), .ZN(n6507) );
  OAI21_X1 U8207 ( .B1(n6508), .B2(n9600), .A(n6507), .ZN(P1_U3249) );
  INV_X1 U8208 ( .A(n9645), .ZN(n9653) );
  INV_X1 U8209 ( .A(n6509), .ZN(n6510) );
  OAI222_X1 U8210 ( .A1(P1_U3084), .A2(n9653), .B1(n9494), .B2(n6510), .C1(
        n10261), .C2(n9491), .ZN(P1_U3342) );
  INV_X1 U8211 ( .A(n8206), .ZN(n7077) );
  AOI21_X1 U8212 ( .B1(n6514), .B2(n6513), .A(n6512), .ZN(n6523) );
  OAI21_X1 U8213 ( .B1(n6517), .B2(n6516), .A(n6515), .ZN(n6521) );
  INV_X1 U8214 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7433) );
  INV_X1 U8215 ( .A(n9634), .ZN(n9678) );
  NAND2_X1 U8216 ( .A1(n9678), .A2(n6518), .ZN(n6519) );
  NAND2_X1 U8217 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7116) );
  OAI211_X1 U8218 ( .C1(n7433), .C2(n9691), .A(n6519), .B(n7116), .ZN(n6520)
         );
  AOI21_X1 U8219 ( .B1(n9686), .B2(n6521), .A(n6520), .ZN(n6522) );
  OAI21_X1 U8220 ( .B1(n6523), .B2(n9600), .A(n6522), .ZN(P1_U3248) );
  NAND2_X1 U8221 ( .A1(n9862), .A2(n6726), .ZN(n6525) );
  NAND2_X1 U8222 ( .A1(n6525), .A2(n6524), .ZN(n6528) );
  OR2_X1 U8223 ( .A1(n9862), .A2(n6526), .ZN(n6527) );
  AND2_X1 U8224 ( .A1(n6528), .A2(n6527), .ZN(n8262) );
  NOR2_X1 U8225 ( .A1(n8235), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8226 ( .A(n6529), .ZN(n6531) );
  INV_X1 U8227 ( .A(n7147), .ZN(n6530) );
  INV_X1 U8228 ( .A(n7048), .ZN(n6645) );
  OAI222_X1 U8229 ( .A1(n9491), .A2(n6532), .B1(n9494), .B2(n6531), .C1(
        P1_U3084), .C2(n6645), .ZN(P1_U3341) );
  NAND2_X1 U8230 ( .A1(n6101), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6535) );
  NAND2_X1 U8231 ( .A1(n6313), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6534) );
  NAND2_X1 U8232 ( .A1(n6097), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6533) );
  AND3_X1 U8233 ( .A1(n6535), .A2(n6534), .A3(n6533), .ZN(n9137) );
  INV_X1 U8234 ( .A(n9137), .ZN(n8830) );
  NAND2_X1 U8235 ( .A1(P1_U4006), .A2(n8830), .ZN(n6536) );
  OAI21_X1 U8236 ( .B1(P1_U4006), .B2(n5762), .A(n6536), .ZN(P1_U3585) );
  INV_X1 U8237 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n10266) );
  NAND2_X1 U8238 ( .A1(P1_U4006), .A2(n6572), .ZN(n6537) );
  OAI21_X1 U8239 ( .B1(P1_U4006), .B2(n10266), .A(n6537), .ZN(P1_U3555) );
  INV_X1 U8240 ( .A(n6538), .ZN(n6540) );
  INV_X1 U8241 ( .A(n7611), .ZN(n7155) );
  INV_X1 U8242 ( .A(n9668), .ZN(n6541) );
  OAI222_X1 U8243 ( .A1(P1_U3084), .A2(n6541), .B1(n9494), .B2(n6540), .C1(
        n10193), .C2(n9491), .ZN(P1_U3340) );
  INV_X1 U8244 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6543) );
  INV_X1 U8245 ( .A(n6542), .ZN(n6544) );
  INV_X1 U8246 ( .A(n8224), .ZN(n7609) );
  INV_X1 U8247 ( .A(n9677), .ZN(n7059) );
  INV_X1 U8248 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10192) );
  OAI222_X1 U8249 ( .A1(P1_U3084), .A2(n7059), .B1(n9494), .B2(n6544), .C1(
        n10192), .C2(n9491), .ZN(P1_U3339) );
  AND3_X1 U8250 ( .A1(n6545), .A2(n6558), .A3(n7543), .ZN(n6548) );
  NOR2_X1 U8251 ( .A1(n6547), .A2(n6546), .ZN(n6692) );
  NAND2_X1 U8252 ( .A1(n6692), .A2(n9486), .ZN(n6552) );
  NAND2_X1 U8253 ( .A1(n6552), .A2(n9782), .ZN(n6606) );
  NAND2_X1 U8254 ( .A1(n6548), .A2(n6606), .ZN(n6549) );
  NAND2_X1 U8255 ( .A1(n6549), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6551) );
  NAND2_X1 U8256 ( .A1(n9025), .A2(n6698), .ZN(n6693) );
  NOR2_X1 U8257 ( .A1(n6693), .A2(n9485), .ZN(n6550) );
  NAND2_X1 U8258 ( .A1(n6552), .A2(n6550), .ZN(n6607) );
  INV_X1 U8259 ( .A(n6599), .ZN(n6553) );
  NOR2_X1 U8260 ( .A1(n6774), .A2(n6372), .ZN(n9031) );
  NAND2_X1 U8261 ( .A1(n6553), .A2(n9031), .ZN(n8759) );
  NOR2_X1 U8262 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6088), .ZN(n9500) );
  INV_X1 U8263 ( .A(n8730), .ZN(n8751) );
  OR2_X1 U8264 ( .A1(n6774), .A2(n9049), .ZN(n6555) );
  NOR2_X2 U8265 ( .A1(n6599), .A2(n6555), .ZN(n8762) );
  OAI22_X1 U8266 ( .A1(n9742), .A2(n8751), .B1(n8737), .B2(n6942), .ZN(n6556)
         );
  AOI211_X1 U8267 ( .C1(n8739), .C2(n6589), .A(n9500), .B(n6556), .ZN(n6602)
         );
  INV_X1 U8268 ( .A(n6562), .ZN(n6557) );
  NAND2_X1 U8269 ( .A1(n9748), .A2(n5005), .ZN(n6560) );
  NAND2_X2 U8270 ( .A1(n6558), .A2(n6562), .ZN(n6569) );
  INV_X4 U8271 ( .A(n6569), .ZN(n7989) );
  NAND2_X1 U8272 ( .A1(n7989), .A2(n6707), .ZN(n6559) );
  NAND2_X1 U8273 ( .A1(n6560), .A2(n6559), .ZN(n6564) );
  NAND2_X1 U8274 ( .A1(n6561), .A2(n9034), .ZN(n6563) );
  NAND2_X4 U8275 ( .A1(n6563), .A2(n6562), .ZN(n7986) );
  NOR2_X2 U8276 ( .A1(n6569), .A2(n6698), .ZN(n6590) );
  NAND2_X1 U8277 ( .A1(n6590), .A2(n9748), .ZN(n6566) );
  INV_X4 U8278 ( .A(n7935), .ZN(n7901) );
  NAND2_X1 U8279 ( .A1(n7901), .A2(n6707), .ZN(n6565) );
  NAND2_X1 U8280 ( .A1(n6566), .A2(n6565), .ZN(n6612) );
  XNOR2_X1 U8281 ( .A(n6614), .B(n6612), .ZN(n6754) );
  INV_X1 U8282 ( .A(n9694), .ZN(n6694) );
  NAND2_X1 U8283 ( .A1(n6572), .A2(n5005), .ZN(n6568) );
  INV_X1 U8284 ( .A(n6558), .ZN(n6571) );
  NAND2_X1 U8285 ( .A1(n6571), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6567) );
  INV_X1 U8286 ( .A(n6603), .ZN(n6570) );
  NAND2_X1 U8287 ( .A1(n6570), .A2(n7986), .ZN(n6575) );
  AOI22_X1 U8288 ( .A1(n5005), .A2(n9694), .B1(n6571), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n6574) );
  NAND2_X1 U8289 ( .A1(n6590), .A2(n6572), .ZN(n6573) );
  AND2_X1 U8290 ( .A1(n6574), .A2(n6573), .ZN(n6605) );
  NAND2_X1 U8291 ( .A1(n6605), .A2(n6603), .ZN(n6604) );
  NAND2_X1 U8292 ( .A1(n6576), .A2(n5005), .ZN(n6578) );
  NAND2_X1 U8293 ( .A1(n7989), .A2(n9700), .ZN(n6577) );
  NAND2_X1 U8294 ( .A1(n6628), .A2(n6629), .ZN(n6581) );
  INV_X2 U8295 ( .A(n5005), .ZN(n7935) );
  INV_X1 U8296 ( .A(n7935), .ZN(n7811) );
  AOI22_X1 U8297 ( .A1(n6590), .A2(n6576), .B1(n7811), .B2(n9700), .ZN(n6627)
         );
  NAND2_X1 U8298 ( .A1(n6581), .A2(n6580), .ZN(n6585) );
  NAND2_X1 U8299 ( .A1(n6585), .A2(n6584), .ZN(n7859) );
  INV_X1 U8300 ( .A(n7859), .ZN(n6594) );
  NAND2_X1 U8301 ( .A1(n6589), .A2(n5005), .ZN(n6587) );
  NAND2_X1 U8302 ( .A1(n6587), .A2(n6586), .ZN(n6588) );
  NAND2_X1 U8303 ( .A1(n6592), .A2(n6591), .ZN(n6595) );
  INV_X1 U8304 ( .A(n7860), .ZN(n6593) );
  NAND2_X1 U8305 ( .A1(n6596), .A2(n6754), .ZN(n6621) );
  OAI21_X1 U8306 ( .B1(n6754), .B2(n6596), .A(n6621), .ZN(n6600) );
  NAND2_X1 U8307 ( .A1(n9782), .A2(n6597), .ZN(n6598) );
  NAND2_X1 U8308 ( .A1(n6600), .A2(n8744), .ZN(n6601) );
  OAI211_X1 U8309 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n8765), .A(n6602), .B(
        n6601), .ZN(P1_U3216) );
  OAI21_X1 U8310 ( .B1(n6605), .B2(n6603), .A(n6604), .ZN(n9046) );
  AOI22_X1 U8311 ( .A1(n8744), .A2(n9046), .B1(n8762), .B2(n6576), .ZN(n6609)
         );
  NAND3_X1 U8312 ( .A1(n6607), .A2(n6606), .A3(n6690), .ZN(n7861) );
  AOI22_X1 U8313 ( .A1(n8767), .A2(n9694), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n7861), .ZN(n6608) );
  NAND2_X1 U8314 ( .A1(n6609), .A2(n6608), .ZN(P1_U3230) );
  INV_X1 U8315 ( .A(n6610), .ZN(n6783) );
  AND2_X1 U8316 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9582) );
  OAI22_X1 U8317 ( .A1(n9751), .A2(n8751), .B1(n8737), .B2(n6896), .ZN(n6611)
         );
  AOI211_X1 U8318 ( .C1(n8739), .C2(n9748), .A(n9582), .B(n6611), .ZN(n6626)
         );
  INV_X1 U8319 ( .A(n6612), .ZN(n6613) );
  NAND2_X1 U8320 ( .A1(n6614), .A2(n6613), .ZN(n6620) );
  AND2_X1 U8321 ( .A1(n6620), .A2(n6621), .ZN(n6624) );
  NAND2_X1 U8322 ( .A1(n9044), .A2(n5005), .ZN(n6616) );
  NAND2_X1 U8323 ( .A1(n7989), .A2(n6785), .ZN(n6615) );
  NAND2_X1 U8324 ( .A1(n6616), .A2(n6615), .ZN(n6617) );
  NAND2_X1 U8325 ( .A1(n6590), .A2(n9044), .ZN(n6619) );
  NAND2_X1 U8326 ( .A1(n5005), .A2(n6785), .ZN(n6618) );
  NAND2_X1 U8327 ( .A1(n6619), .A2(n6618), .ZN(n6752) );
  XNOR2_X1 U8328 ( .A(n6751), .B(n6752), .ZN(n6623) );
  NAND2_X1 U8329 ( .A1(n6621), .A2(n6757), .ZN(n6622) );
  OAI211_X1 U8330 ( .C1(n6624), .C2(n6623), .A(n6622), .B(n8744), .ZN(n6625)
         );
  OAI211_X1 U8331 ( .C1(n8765), .C2(n6783), .A(n6626), .B(n6625), .ZN(P1_U3228) );
  XNOR2_X1 U8332 ( .A(n6628), .B(n6627), .ZN(n6630) );
  XNOR2_X1 U8333 ( .A(n6629), .B(n6630), .ZN(n6633) );
  AOI22_X1 U8334 ( .A1(n8739), .A2(n6572), .B1(n8762), .B2(n6589), .ZN(n6632)
         );
  AOI22_X1 U8335 ( .A1(n8767), .A2(n9700), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n7861), .ZN(n6631) );
  OAI211_X1 U8336 ( .C1(n6633), .C2(n7995), .A(n6632), .B(n6631), .ZN(P1_U3220) );
  INV_X1 U8337 ( .A(n6634), .ZN(n6688) );
  AOI22_X1 U8338 ( .A1(n7202), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n9488), .ZN(n6635) );
  OAI21_X1 U8339 ( .B1(n6688), .B2(n9494), .A(n6635), .ZN(P1_U3338) );
  INV_X1 U8340 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6636) );
  MUX2_X1 U8341 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6636), .S(n7048), .Z(n6642)
         );
  INV_X1 U8342 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6637) );
  MUX2_X1 U8343 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n6637), .S(n9645), .Z(n9650)
         );
  OAI21_X1 U8344 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6649), .A(n6638), .ZN(
        n9619) );
  INV_X1 U8345 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6639) );
  MUX2_X1 U8346 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n6639), .S(n6652), .Z(n9620)
         );
  NAND2_X1 U8347 ( .A1(n9619), .A2(n9620), .ZN(n9618) );
  OAI21_X1 U8348 ( .B1(n6652), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9618), .ZN(
        n9631) );
  INV_X1 U8349 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6640) );
  MUX2_X1 U8350 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6640), .S(n6646), .Z(n9632)
         );
  NAND2_X1 U8351 ( .A1(n9631), .A2(n9632), .ZN(n9630) );
  OAI21_X1 U8352 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n6646), .A(n9630), .ZN(
        n9652) );
  NAND2_X1 U8353 ( .A1(n9650), .A2(n9652), .ZN(n9647) );
  OAI21_X1 U8354 ( .B1(n9645), .B2(P1_REG1_REG_11__SCAN_IN), .A(n9647), .ZN(
        n6641) );
  NAND2_X1 U8355 ( .A1(n6642), .A2(n6641), .ZN(n7047) );
  OAI21_X1 U8356 ( .B1(n6642), .B2(n6641), .A(n7047), .ZN(n6643) );
  NAND2_X1 U8357 ( .A1(n9686), .A2(n6643), .ZN(n6644) );
  NAND2_X1 U8358 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7588) );
  OAI211_X1 U8359 ( .C1(n6645), .C2(n9634), .A(n6644), .B(n7588), .ZN(n6657)
         );
  NAND2_X1 U8360 ( .A1(n6646), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6654) );
  INV_X1 U8361 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6647) );
  MUX2_X1 U8362 ( .A(n6647), .B(P1_REG2_REG_10__SCAN_IN), .S(n6646), .Z(n6648)
         );
  INV_X1 U8363 ( .A(n6648), .ZN(n9639) );
  INV_X1 U8364 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7217) );
  NOR2_X1 U8365 ( .A1(n6649), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6651) );
  MUX2_X1 U8366 ( .A(n7217), .B(P1_REG2_REG_9__SCAN_IN), .S(n6652), .Z(n6653)
         );
  INV_X1 U8367 ( .A(n6653), .ZN(n9626) );
  NAND2_X1 U8368 ( .A1(n9627), .A2(n9626), .ZN(n9625) );
  OAI21_X1 U8369 ( .B1(n7217), .B2(n9622), .A(n9625), .ZN(n9640) );
  NAND2_X1 U8370 ( .A1(n9639), .A2(n9640), .ZN(n9638) );
  NAND2_X1 U8371 ( .A1(n6654), .A2(n9638), .ZN(n9657) );
  INV_X1 U8372 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10029) );
  NOR2_X1 U8373 ( .A1(n9653), .A2(n10029), .ZN(n9656) );
  OAI22_X1 U8374 ( .A1(n9657), .A2(n9656), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n9645), .ZN(n9654) );
  NAND2_X1 U8375 ( .A1(n7048), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7057) );
  OAI21_X1 U8376 ( .B1(n7048), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7057), .ZN(
        n6655) );
  AOI211_X1 U8377 ( .C1(n9654), .C2(n6655), .A(n7055), .B(n9600), .ZN(n6656)
         );
  AOI211_X1 U8378 ( .C1(n9649), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n6657), .B(
        n6656), .ZN(n6658) );
  INV_X1 U8379 ( .A(n6658), .ZN(P1_U3253) );
  INV_X1 U8380 ( .A(n6659), .ZN(n6662) );
  AOI22_X1 U8381 ( .A1(n7835), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n7541), .ZN(n6660) );
  OAI21_X1 U8382 ( .B1(n6662), .B2(n8025), .A(n6660), .ZN(P2_U3342) );
  AOI22_X1 U8383 ( .A1(n9071), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9488), .ZN(n6661) );
  OAI21_X1 U8384 ( .B1(n6662), .B2(n9494), .A(n6661), .ZN(P1_U3337) );
  NOR2_X1 U8385 ( .A1(n9862), .A2(n7977), .ZN(n6663) );
  NAND2_X1 U8386 ( .A1(n6664), .A2(n6663), .ZN(n7262) );
  NAND2_X1 U8387 ( .A1(n7264), .A2(n7261), .ZN(n6665) );
  INV_X1 U8388 ( .A(n7270), .ZN(n7263) );
  INV_X1 U8389 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6687) );
  XNOR2_X1 U8390 ( .A(n5689), .B(n7266), .ZN(n6666) );
  NAND2_X1 U8391 ( .A1(n6666), .A2(n7451), .ZN(n8508) );
  INV_X1 U8392 ( .A(n6669), .ZN(n6672) );
  NAND2_X1 U8393 ( .A1(n6669), .A2(n6668), .ZN(n6903) );
  INV_X1 U8394 ( .A(n6903), .ZN(n6670) );
  AOI21_X1 U8395 ( .B1(n6672), .B2(n6671), .A(n6670), .ZN(n7895) );
  INV_X1 U8396 ( .A(n7408), .ZN(n6679) );
  INV_X1 U8397 ( .A(n6675), .ZN(n6676) );
  NOR2_X1 U8398 ( .A1(n6677), .A2(n6676), .ZN(n6678) );
  AOI211_X1 U8399 ( .C1(n6679), .C2(n6669), .A(n8488), .B(n6678), .ZN(n6681)
         );
  OAI22_X1 U8400 ( .A1(n6680), .A2(n8502), .B1(n5717), .B2(n8500), .ZN(n7975)
         );
  NOR2_X1 U8401 ( .A1(n6681), .A2(n7975), .ZN(n7891) );
  NAND2_X1 U8402 ( .A1(n7981), .A2(n9870), .ZN(n6905) );
  NAND2_X1 U8403 ( .A1(n7890), .A2(n8020), .ZN(n6682) );
  NAND3_X1 U8404 ( .A1(n6905), .A2(n6683), .A3(n6682), .ZN(n7888) );
  INV_X1 U8405 ( .A(n7888), .ZN(n6684) );
  AOI21_X1 U8406 ( .B1(n7890), .B2(n9886), .A(n6684), .ZN(n6685) );
  OAI211_X1 U8407 ( .C1(n8624), .C2(n7895), .A(n7891), .B(n6685), .ZN(n6704)
         );
  NAND2_X1 U8408 ( .A1(n6704), .A2(n9930), .ZN(n6686) );
  OAI21_X1 U8409 ( .B1(n9930), .B2(n6687), .A(n6686), .ZN(P2_U3454) );
  INV_X1 U8410 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9045) );
  NAND3_X1 U8411 ( .A1(n6692), .A2(n6691), .A3(n6690), .ZN(n6779) );
  INV_X1 U8412 ( .A(n6693), .ZN(n9699) );
  NAND2_X1 U8413 ( .A1(n9347), .A2(n9694), .ZN(n6702) );
  INV_X1 U8414 ( .A(n9708), .ZN(n8967) );
  NAND2_X1 U8415 ( .A1(n6572), .A2(n6694), .ZN(n8968) );
  INV_X1 U8416 ( .A(n8968), .ZN(n6696) );
  INV_X1 U8417 ( .A(n6698), .ZN(n6695) );
  OAI211_X1 U8418 ( .C1(n8967), .C2(n6696), .A(n6774), .B(n6695), .ZN(n6697)
         );
  OAI21_X1 U8419 ( .B1(n6996), .B2(n9733), .A(n6697), .ZN(n9724) );
  INV_X1 U8420 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6699) );
  NAND2_X1 U8421 ( .A1(n9694), .A2(n6698), .ZN(n9722) );
  OAI22_X1 U8422 ( .A1(n9301), .A2(n6699), .B1(n9704), .B2(n9722), .ZN(n6700)
         );
  OAI21_X1 U8423 ( .B1(n9724), .B2(n6700), .A(n9716), .ZN(n6701) );
  OAI211_X1 U8424 ( .C1(n9045), .C2(n9716), .A(n6702), .B(n6701), .ZN(P1_U3291) );
  INV_X1 U8425 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6734) );
  NAND2_X1 U8426 ( .A1(n6704), .A2(n9945), .ZN(n6705) );
  OAI21_X1 U8427 ( .B1(n9945), .B2(n6734), .A(n6705), .ZN(P2_U3521) );
  INV_X1 U8428 ( .A(n6780), .ZN(n6706) );
  AOI211_X1 U8429 ( .C1(n6707), .C2(n6998), .A(n9319), .B(n6706), .ZN(n9740)
         );
  XOR2_X1 U8430 ( .A(n6709), .B(n6708), .Z(n6714) );
  XOR2_X1 U8431 ( .A(n6709), .B(n9006), .Z(n6712) );
  OAI22_X1 U8432 ( .A1(n6942), .A2(n9733), .B1(n6710), .B2(n9361), .ZN(n6711)
         );
  AOI21_X1 U8433 ( .B1(n6712), .B2(n9706), .A(n6711), .ZN(n6713) );
  OAI21_X1 U8434 ( .B1(n6714), .B2(n9712), .A(n6713), .ZN(n9743) );
  AOI21_X1 U8435 ( .B1(n9740), .B2(n9215), .A(n9743), .ZN(n6719) );
  INV_X1 U8436 ( .A(n9716), .ZN(n9241) );
  NOR2_X1 U8437 ( .A1(n9215), .A2(n6562), .ZN(n9715) );
  NAND2_X1 U8438 ( .A1(n9716), .A2(n9715), .ZN(n7489) );
  INV_X1 U8439 ( .A(n7489), .ZN(n6717) );
  INV_X1 U8440 ( .A(n6714), .ZN(n9745) );
  INV_X1 U8441 ( .A(n9716), .ZN(n9208) );
  INV_X1 U8442 ( .A(n9301), .ZN(n9701) );
  AOI22_X1 U8443 ( .A1(n9208), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9701), .B2(
        n6088), .ZN(n6715) );
  OAI21_X1 U8444 ( .B1(n9742), .B2(n9326), .A(n6715), .ZN(n6716) );
  AOI21_X1 U8445 ( .B1(n6717), .B2(n9745), .A(n6716), .ZN(n6718) );
  OAI21_X1 U8446 ( .B1(n6719), .B2(n9241), .A(n6718), .ZN(P1_U3288) );
  INV_X1 U8447 ( .A(n6720), .ZN(n6723) );
  AOI22_X1 U8448 ( .A1(n9082), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9488), .ZN(n6721) );
  OAI21_X1 U8449 ( .B1(n6723), .B2(n9494), .A(n6721), .ZN(P1_U3336) );
  AOI22_X1 U8450 ( .A1(n8238), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n7541), .ZN(n6722) );
  OAI21_X1 U8451 ( .B1(n6723), .B2(n8025), .A(n6722), .ZN(P2_U3341) );
  NAND2_X1 U8452 ( .A1(n6724), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6725) );
  OAI211_X1 U8453 ( .C1(n9862), .C2(n6727), .A(n6726), .B(n6725), .ZN(n6741)
         );
  NAND2_X1 U8454 ( .A1(n6741), .A2(n6739), .ZN(n6728) );
  NAND2_X1 U8455 ( .A1(n6728), .A2(n8177), .ZN(n6731) );
  INV_X1 U8456 ( .A(n8256), .ZN(n7156) );
  INV_X1 U8457 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10028) );
  MUX2_X1 U8458 ( .A(n10028), .B(P2_REG2_REG_3__SCAN_IN), .S(n6790), .Z(n6733)
         );
  INV_X1 U8459 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n8548) );
  INV_X1 U8460 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7892) );
  XNOR2_X1 U8461 ( .A(n8192), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n8191) );
  NAND2_X1 U8462 ( .A1(n8190), .A2(n8191), .ZN(n8189) );
  OAI21_X1 U8463 ( .B1(n8548), .B2(n8192), .A(n8189), .ZN(n6732) );
  INV_X1 U8464 ( .A(n8649), .ZN(n6730) );
  INV_X1 U8465 ( .A(n8646), .ZN(n6729) );
  NAND3_X1 U8466 ( .A1(n6731), .A2(n6730), .A3(n6729), .ZN(n8254) );
  NAND2_X1 U8467 ( .A1(n6732), .A2(n6733), .ZN(n6796) );
  OAI211_X1 U8468 ( .C1(n6733), .C2(n6732), .A(n8253), .B(n6796), .ZN(n6749)
         );
  INV_X1 U8469 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6746) );
  XNOR2_X1 U8470 ( .A(n6790), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n6743) );
  XNOR2_X1 U8471 ( .A(n8192), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n8196) );
  MUX2_X1 U8472 ( .A(n6734), .B(P2_REG1_REG_1__SCAN_IN), .S(n6735), .Z(n8184)
         );
  AND2_X1 U8473 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n8183) );
  NAND2_X1 U8474 ( .A1(n8184), .A2(n8183), .ZN(n8182) );
  INV_X1 U8475 ( .A(n6735), .ZN(n8181) );
  NAND2_X1 U8476 ( .A1(n8181), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6736) );
  NAND2_X1 U8477 ( .A1(n8182), .A2(n6736), .ZN(n8195) );
  NAND2_X1 U8478 ( .A1(n8196), .A2(n8195), .ZN(n8194) );
  INV_X1 U8479 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6737) );
  OR2_X1 U8480 ( .A1(n8192), .A2(n6737), .ZN(n6738) );
  NAND2_X1 U8481 ( .A1(n8194), .A2(n6738), .ZN(n6742) );
  AND2_X1 U8482 ( .A1(n6739), .A2(n8649), .ZN(n6740) );
  NAND2_X1 U8483 ( .A1(n6742), .A2(n6743), .ZN(n6792) );
  OAI211_X1 U8484 ( .C1(n6743), .C2(n6742), .A(n8258), .B(n6792), .ZN(n6745)
         );
  NAND2_X1 U8485 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3152), .ZN(n6744) );
  OAI211_X1 U8486 ( .C1(n8262), .C2(n6746), .A(n6745), .B(n6744), .ZN(n6747)
         );
  INV_X1 U8487 ( .A(n6747), .ZN(n6748) );
  OAI211_X1 U8488 ( .C1(n7156), .C2(n6790), .A(n6749), .B(n6748), .ZN(P2_U3248) );
  INV_X1 U8489 ( .A(n6750), .ZN(n6932) );
  AOI22_X1 U8490 ( .A1(n7983), .A2(n9768), .B1(n7901), .B2(n8845), .ZN(n6769)
         );
  INV_X1 U8491 ( .A(n6751), .ZN(n6753) );
  NAND2_X1 U8492 ( .A1(n6753), .A2(n6752), .ZN(n6755) );
  AND2_X1 U8493 ( .A1(n6754), .A2(n6755), .ZN(n6759) );
  INV_X1 U8494 ( .A(n6755), .ZN(n6756) );
  NOR2_X1 U8495 ( .A1(n6757), .A2(n6756), .ZN(n6758) );
  NAND2_X1 U8496 ( .A1(n9768), .A2(n7901), .ZN(n6762) );
  NAND2_X1 U8497 ( .A1(n7989), .A2(n8845), .ZN(n6761) );
  NAND2_X1 U8498 ( .A1(n6762), .A2(n6761), .ZN(n6763) );
  XNOR2_X1 U8499 ( .A(n6763), .B(n7986), .ZN(n6764) );
  NAND2_X1 U8500 ( .A1(n6765), .A2(n6764), .ZN(n6766) );
  OAI21_X1 U8501 ( .B1(n6769), .B2(n6768), .A(n6767), .ZN(n6770) );
  NAND2_X1 U8502 ( .A1(n6770), .A2(n8744), .ZN(n6773) );
  AND2_X1 U8503 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9591) );
  OAI22_X1 U8504 ( .A1(n9763), .A2(n8751), .B1(n8737), .B2(n7027), .ZN(n6771)
         );
  AOI211_X1 U8505 ( .C1(n8739), .C2(n9044), .A(n9591), .B(n6771), .ZN(n6772)
         );
  OAI211_X1 U8506 ( .C1(n8765), .C2(n6932), .A(n6773), .B(n6772), .ZN(P1_U3225) );
  XNOR2_X1 U8507 ( .A(n6776), .B(n6775), .ZN(n9755) );
  XNOR2_X1 U8508 ( .A(n8843), .B(n6777), .ZN(n6778) );
  NOR2_X1 U8509 ( .A1(n6778), .A2(n9784), .ZN(n9753) );
  NAND2_X1 U8510 ( .A1(n9716), .A2(n9794), .ZN(n9338) );
  NOR2_X2 U8511 ( .A1(n6779), .A2(n9704), .ZN(n9321) );
  INV_X1 U8512 ( .A(n9321), .ZN(n9344) );
  NAND2_X1 U8513 ( .A1(n6780), .A2(n6785), .ZN(n6781) );
  NAND2_X1 U8514 ( .A1(n6781), .A2(n9695), .ZN(n6782) );
  OR2_X1 U8515 ( .A1(n6940), .A2(n6782), .ZN(n9750) );
  OAI22_X1 U8516 ( .A1(n9344), .A2(n9750), .B1(n6783), .B2(n9301), .ZN(n6784)
         );
  AOI21_X1 U8517 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n9241), .A(n6784), .ZN(
        n6787) );
  AND2_X1 U8518 ( .A1(n9716), .A2(n9791), .ZN(n9335) );
  AOI22_X1 U8519 ( .A1(n9347), .A2(n6785), .B1(n9335), .B2(n9768), .ZN(n6786)
         );
  OAI211_X1 U8520 ( .C1(n9734), .C2(n9338), .A(n6787), .B(n6786), .ZN(n6788)
         );
  AOI21_X1 U8521 ( .B1(n9753), .B2(n9716), .A(n6788), .ZN(n6789) );
  OAI21_X1 U8522 ( .B1(n9333), .B2(n9755), .A(n6789), .ZN(P1_U3287) );
  INV_X1 U8523 ( .A(n6806), .ZN(n6820) );
  XNOR2_X1 U8524 ( .A(n6806), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n6794) );
  INV_X1 U8525 ( .A(n6790), .ZN(n6797) );
  NAND2_X1 U8526 ( .A1(n6797), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6791) );
  NAND2_X1 U8527 ( .A1(n6792), .A2(n6791), .ZN(n6793) );
  NAND2_X1 U8528 ( .A1(n6793), .A2(n6794), .ZN(n6808) );
  OAI211_X1 U8529 ( .C1(n6794), .C2(n6793), .A(n8258), .B(n6808), .ZN(n6795)
         );
  NAND2_X1 U8530 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7039) );
  OAI211_X1 U8531 ( .C1(n8262), .C2(n10107), .A(n6795), .B(n7039), .ZN(n6802)
         );
  INV_X1 U8532 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6798) );
  MUX2_X1 U8533 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6798), .S(n6806), .Z(n6799)
         );
  AOI211_X1 U8534 ( .C1(n6800), .C2(n6799), .A(n6819), .B(n8254), .ZN(n6801)
         );
  AOI211_X1 U8535 ( .C1(n8256), .C2(n6820), .A(n6802), .B(n6801), .ZN(n6803)
         );
  INV_X1 U8536 ( .A(n6803), .ZN(P2_U3249) );
  INV_X1 U8537 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10009) );
  OR2_X1 U8538 ( .A1(n6836), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6804) );
  NAND2_X1 U8539 ( .A1(n6836), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6827) );
  AND2_X1 U8540 ( .A1(n6804), .A2(n6827), .ZN(n6816) );
  INV_X1 U8541 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6805) );
  OR2_X1 U8542 ( .A1(n6806), .A2(n6805), .ZN(n6807) );
  NAND2_X1 U8543 ( .A1(n6808), .A2(n6807), .ZN(n6844) );
  INV_X1 U8544 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6810) );
  INV_X1 U8545 ( .A(n6811), .ZN(n6851) );
  NAND2_X1 U8546 ( .A1(n6851), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6812) );
  INV_X1 U8547 ( .A(n6812), .ZN(n6809) );
  AOI21_X1 U8548 ( .B1(n6811), .B2(n6810), .A(n6809), .ZN(n6845) );
  NAND2_X1 U8549 ( .A1(n6844), .A2(n6845), .ZN(n6843) );
  NAND2_X1 U8550 ( .A1(n6843), .A2(n6812), .ZN(n6854) );
  XNOR2_X1 U8551 ( .A(n6813), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n6855) );
  NAND2_X1 U8552 ( .A1(n6854), .A2(n6855), .ZN(n6853) );
  NAND2_X1 U8553 ( .A1(n6862), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6814) );
  NAND2_X1 U8554 ( .A1(n6853), .A2(n6814), .ZN(n6815) );
  NAND2_X1 U8555 ( .A1(n6815), .A2(n6816), .ZN(n6828) );
  OAI211_X1 U8556 ( .C1(n6816), .C2(n6815), .A(n8258), .B(n6828), .ZN(n6818)
         );
  NAND2_X1 U8557 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3152), .ZN(n6817) );
  OAI211_X1 U8558 ( .C1(n8262), .C2(n10009), .A(n6818), .B(n6817), .ZN(n6825)
         );
  NAND2_X1 U8559 ( .A1(n6851), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6821) );
  OAI21_X1 U8560 ( .B1(n6851), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6821), .ZN(
        n6848) );
  NOR2_X1 U8561 ( .A1(n4436), .A2(n6848), .ZN(n6847) );
  XNOR2_X1 U8562 ( .A(n6862), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n6858) );
  INV_X1 U8563 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7279) );
  MUX2_X1 U8564 ( .A(n7279), .B(P2_REG2_REG_7__SCAN_IN), .S(n6836), .Z(n6822)
         );
  AOI211_X1 U8565 ( .C1(n6823), .C2(n6822), .A(n8254), .B(n6835), .ZN(n6824)
         );
  AOI211_X1 U8566 ( .C1(n8256), .C2(n6836), .A(n6825), .B(n6824), .ZN(n6826)
         );
  INV_X1 U8567 ( .A(n6826), .ZN(P2_U3252) );
  INV_X1 U8568 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n6834) );
  AND2_X1 U8569 ( .A1(n6828), .A2(n6827), .ZN(n6831) );
  INV_X1 U8570 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6829) );
  MUX2_X1 U8571 ( .A(n6829), .B(P2_REG1_REG_8__SCAN_IN), .S(n6873), .Z(n6830)
         );
  NOR2_X1 U8572 ( .A1(n6831), .A2(n6830), .ZN(n6865) );
  AOI21_X1 U8573 ( .B1(n6831), .B2(n6830), .A(n6865), .ZN(n6832) );
  NAND2_X1 U8574 ( .A1(n8258), .A2(n6832), .ZN(n6833) );
  NAND2_X1 U8575 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(n8130), .ZN(n7172) );
  OAI211_X1 U8576 ( .C1(n8262), .C2(n6834), .A(n6833), .B(n7172), .ZN(n6841)
         );
  AOI21_X1 U8577 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n6836), .A(n6835), .ZN(
        n6839) );
  NAND2_X1 U8578 ( .A1(n6873), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6837) );
  OAI21_X1 U8579 ( .B1(n6873), .B2(P2_REG2_REG_8__SCAN_IN), .A(n6837), .ZN(
        n6838) );
  NOR2_X1 U8580 ( .A1(n6839), .A2(n6838), .ZN(n6872) );
  AOI211_X1 U8581 ( .C1(n6839), .C2(n6838), .A(n6872), .B(n8254), .ZN(n6840)
         );
  AOI211_X1 U8582 ( .C1(n8256), .C2(n6873), .A(n6841), .B(n6840), .ZN(n6842)
         );
  INV_X1 U8583 ( .A(n6842), .ZN(P2_U3253) );
  INV_X1 U8584 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10234) );
  OAI211_X1 U8585 ( .C1(n6845), .C2(n6844), .A(n8258), .B(n6843), .ZN(n6846)
         );
  NAND2_X1 U8586 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6922) );
  OAI211_X1 U8587 ( .C1(n8262), .C2(n10234), .A(n6846), .B(n6922), .ZN(n6850)
         );
  AOI211_X1 U8588 ( .C1(n4436), .C2(n6848), .A(n6847), .B(n8254), .ZN(n6849)
         );
  AOI211_X1 U8589 ( .C1(n8256), .C2(n6851), .A(n6850), .B(n6849), .ZN(n6852)
         );
  INV_X1 U8590 ( .A(n6852), .ZN(P2_U3250) );
  INV_X1 U8591 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7428) );
  OAI211_X1 U8592 ( .C1(n6855), .C2(n6854), .A(n8258), .B(n6853), .ZN(n6856)
         );
  NAND2_X1 U8593 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(n8130), .ZN(n7104) );
  OAI211_X1 U8594 ( .C1(n8262), .C2(n7428), .A(n6856), .B(n7104), .ZN(n6861)
         );
  AOI211_X1 U8595 ( .C1(n6859), .C2(n6858), .A(n6857), .B(n8254), .ZN(n6860)
         );
  AOI211_X1 U8596 ( .C1(n8256), .C2(n6862), .A(n6861), .B(n6860), .ZN(n6863)
         );
  INV_X1 U8597 ( .A(n6863), .ZN(P2_U3251) );
  INV_X1 U8598 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10158) );
  INV_X1 U8599 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6864) );
  MUX2_X1 U8600 ( .A(n6864), .B(P2_REG1_REG_10__SCAN_IN), .S(n7076), .Z(n6868)
         );
  AOI21_X1 U8601 ( .B1(n6873), .B2(P2_REG1_REG_8__SCAN_IN), .A(n6865), .ZN(
        n6881) );
  INV_X1 U8602 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6866) );
  MUX2_X1 U8603 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6866), .S(n6874), .Z(n6882)
         );
  NOR2_X1 U8604 ( .A1(n6881), .A2(n6882), .ZN(n6880) );
  AOI21_X1 U8605 ( .B1(n6890), .B2(P2_REG1_REG_9__SCAN_IN), .A(n6880), .ZN(
        n6867) );
  NOR2_X1 U8606 ( .A1(n6867), .A2(n6868), .ZN(n7068) );
  AOI21_X1 U8607 ( .B1(n6868), .B2(n6867), .A(n7068), .ZN(n6869) );
  NAND2_X1 U8608 ( .A1(n8258), .A2(n6869), .ZN(n6871) );
  NAND2_X1 U8609 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(n8130), .ZN(n6870) );
  OAI211_X1 U8610 ( .C1(n8262), .C2(n10158), .A(n6871), .B(n6870), .ZN(n6878)
         );
  INV_X1 U8611 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7512) );
  MUX2_X1 U8612 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7512), .S(n6874), .Z(n6886)
         );
  MUX2_X1 U8613 ( .A(n7567), .B(P2_REG2_REG_10__SCAN_IN), .S(n7076), .Z(n6875)
         );
  AOI211_X1 U8614 ( .C1(n6876), .C2(n6875), .A(n7075), .B(n8254), .ZN(n6877)
         );
  AOI211_X1 U8615 ( .C1(n8256), .C2(n7076), .A(n6878), .B(n6877), .ZN(n6879)
         );
  INV_X1 U8616 ( .A(n6879), .ZN(P2_U3255) );
  INV_X1 U8617 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7440) );
  AOI21_X1 U8618 ( .B1(n6882), .B2(n6881), .A(n6880), .ZN(n6883) );
  NAND2_X1 U8619 ( .A1(n8258), .A2(n6883), .ZN(n6884) );
  NAND2_X1 U8620 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7317) );
  OAI211_X1 U8621 ( .C1(n8262), .C2(n7440), .A(n6884), .B(n7317), .ZN(n6889)
         );
  AOI211_X1 U8622 ( .C1(n6887), .C2(n6886), .A(n6885), .B(n8254), .ZN(n6888)
         );
  AOI211_X1 U8623 ( .C1(n8256), .C2(n6890), .A(n6889), .B(n6888), .ZN(n6891)
         );
  INV_X1 U8624 ( .A(n6891), .ZN(P2_U3254) );
  OAI21_X1 U8625 ( .B1(n4485), .B2(n6893), .A(n6892), .ZN(n9777) );
  INV_X1 U8626 ( .A(n9777), .ZN(n9774) );
  OAI21_X1 U8627 ( .B1(n8857), .B2(n4484), .A(n6894), .ZN(n6895) );
  NAND2_X1 U8628 ( .A1(n6895), .A2(n9706), .ZN(n9773) );
  MUX2_X1 U8629 ( .A(n9773), .B(n10013), .S(n9241), .Z(n6901) );
  OAI211_X1 U8630 ( .C1(n6938), .C2(n6988), .A(n9695), .B(n7028), .ZN(n9771)
         );
  INV_X1 U8631 ( .A(n9771), .ZN(n6899) );
  OAI22_X1 U8632 ( .A1(n9326), .A2(n6988), .B1(n9301), .B2(n6992), .ZN(n6898)
         );
  INV_X1 U8633 ( .A(n9335), .ZN(n9283) );
  OAI22_X1 U8634 ( .A1(n9283), .A2(n7188), .B1(n6896), .B2(n9338), .ZN(n6897)
         );
  AOI211_X1 U8635 ( .C1(n9321), .C2(n6899), .A(n6898), .B(n6897), .ZN(n6900)
         );
  OAI211_X1 U8636 ( .C1(n9774), .C2(n9333), .A(n6901), .B(n6900), .ZN(P1_U3285) );
  NAND2_X1 U8637 ( .A1(n8024), .A2(n7981), .ZN(n6902) );
  NAND2_X1 U8638 ( .A1(n6903), .A2(n6902), .ZN(n6904) );
  NAND2_X1 U8639 ( .A1(n6904), .A2(n6910), .ZN(n6951) );
  OAI21_X1 U8640 ( .B1(n6904), .B2(n6910), .A(n6951), .ZN(n8546) );
  AND2_X1 U8641 ( .A1(n6905), .A2(n8545), .ZN(n6906) );
  NOR2_X1 U8642 ( .A1(n6905), .A2(n8545), .ZN(n7328) );
  OR2_X1 U8643 ( .A1(n6906), .A2(n7328), .ZN(n8550) );
  OAI22_X1 U8644 ( .A1(n8550), .A2(n9922), .B1(n6949), .B2(n9921), .ZN(n6912)
         );
  INV_X1 U8645 ( .A(n6907), .ZN(n6908) );
  AOI21_X1 U8646 ( .B1(n6910), .B2(n6909), .A(n6908), .ZN(n6911) );
  OAI222_X1 U8647 ( .A1(n8500), .A2(n6956), .B1(n8502), .B2(n8024), .C1(n8488), 
        .C2(n6911), .ZN(n8547) );
  AOI211_X1 U8648 ( .C1(n9927), .C2(n8546), .A(n6912), .B(n8547), .ZN(n6929)
         );
  NAND2_X1 U8649 ( .A1(n9943), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6913) );
  OAI21_X1 U8650 ( .B1(n6929), .B2(n9943), .A(n6913), .ZN(P2_U3522) );
  INV_X1 U8651 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6914) );
  INV_X1 U8652 ( .A(n8258), .ZN(n7612) );
  OAI211_X1 U8653 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n7612), .A(n7156), .B(
        P2_IR_REG_0__SCAN_IN), .ZN(n6915) );
  AOI21_X1 U8654 ( .B1(n8253), .B2(n6914), .A(n6915), .ZN(n6919) );
  AOI21_X1 U8655 ( .B1(n8258), .B2(P2_REG1_REG_0__SCAN_IN), .A(
        P2_IR_REG_0__SCAN_IN), .ZN(n6918) );
  AOI22_X1 U8656 ( .A1(n8235), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n6917) );
  NAND3_X1 U8657 ( .A1(n6915), .A2(n8253), .A3(P2_REG2_REG_0__SCAN_IN), .ZN(
        n6916) );
  OAI211_X1 U8658 ( .C1(n6919), .C2(n6918), .A(n6917), .B(n6916), .ZN(P2_U3245) );
  XNOR2_X1 U8659 ( .A(n6921), .B(n6920), .ZN(n6928) );
  INV_X1 U8660 ( .A(n8142), .ZN(n7976) );
  OAI22_X1 U8661 ( .A1(n7868), .A2(n8502), .B1(n7276), .B2(n8500), .ZN(n7011)
         );
  INV_X1 U8662 ( .A(n6922), .ZN(n6923) );
  AOI21_X1 U8663 ( .B1(n7976), .B2(n7011), .A(n6923), .ZN(n6924) );
  OAI21_X1 U8664 ( .B1(n6925), .B2(n9840), .A(n6924), .ZN(n6926) );
  AOI21_X1 U8665 ( .B1(n8158), .B2(n7015), .A(n6926), .ZN(n6927) );
  OAI21_X1 U8666 ( .B1(n6928), .B2(n9826), .A(n6927), .ZN(P2_U3229) );
  INV_X1 U8667 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6931) );
  OR2_X1 U8668 ( .A1(n6929), .A2(n9928), .ZN(n6930) );
  OAI21_X1 U8669 ( .B1(n9930), .B2(n6931), .A(n6930), .ZN(P2_U3457) );
  OAI22_X1 U8670 ( .A1(n9716), .A2(n9980), .B1(n6932), .B2(n9301), .ZN(n6937)
         );
  INV_X1 U8671 ( .A(n9765), .ZN(n6935) );
  AND2_X1 U8672 ( .A1(n6934), .A2(n6933), .ZN(n9760) );
  NOR3_X1 U8673 ( .A1(n6935), .A2(n9760), .A3(n9333), .ZN(n6936) );
  AOI211_X1 U8674 ( .C1(n9347), .C2(n8845), .A(n6937), .B(n6936), .ZN(n6948)
         );
  INV_X1 U8675 ( .A(n6938), .ZN(n6939) );
  OAI211_X1 U8676 ( .C1(n9763), .C2(n6940), .A(n6939), .B(n9695), .ZN(n9761)
         );
  AOI21_X1 U8677 ( .B1(n6941), .B2(n6113), .A(n9784), .ZN(n6945) );
  OAI22_X1 U8678 ( .A1(n6942), .A2(n9361), .B1(n7027), .B2(n9733), .ZN(n6943)
         );
  AOI21_X1 U8679 ( .B1(n6945), .B2(n6944), .A(n6943), .ZN(n9762) );
  OAI21_X1 U8680 ( .B1(n9704), .B2(n9761), .A(n9762), .ZN(n6946) );
  NAND2_X1 U8681 ( .A1(n6946), .A2(n9716), .ZN(n6947) );
  NAND2_X1 U8682 ( .A1(n6948), .A2(n6947), .ZN(P1_U3286) );
  INV_X1 U8683 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6963) );
  NAND2_X1 U8684 ( .A1(n5717), .A2(n6949), .ZN(n6950) );
  OAI21_X1 U8685 ( .B1(n6953), .B2(n6954), .A(n7005), .ZN(n7287) );
  INV_X1 U8686 ( .A(n7287), .ZN(n6961) );
  XNOR2_X1 U8687 ( .A(n6955), .B(n5721), .ZN(n6958) );
  OAI22_X1 U8688 ( .A1(n6956), .A2(n8502), .B1(n7258), .B2(n8500), .ZN(n6957)
         );
  AOI21_X1 U8689 ( .B1(n6958), .B2(n9843), .A(n6957), .ZN(n7285) );
  NAND2_X1 U8690 ( .A1(n7327), .A2(n7290), .ZN(n6959) );
  AND2_X1 U8691 ( .A1(n7013), .A2(n6959), .ZN(n7283) );
  AOI22_X1 U8692 ( .A1(n7283), .A2(n9853), .B1(n7290), .B2(n9886), .ZN(n6960)
         );
  OAI211_X1 U8693 ( .C1(n6961), .C2(n8624), .A(n7285), .B(n6960), .ZN(n6968)
         );
  NAND2_X1 U8694 ( .A1(n6968), .A2(n9930), .ZN(n6962) );
  OAI21_X1 U8695 ( .B1(n9930), .B2(n6963), .A(n6962), .ZN(P2_U3463) );
  INV_X1 U8696 ( .A(n6964), .ZN(n6967) );
  AOI22_X1 U8697 ( .A1(n8250), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n7541), .ZN(n6965) );
  OAI21_X1 U8698 ( .B1(n6967), .B2(n8025), .A(n6965), .ZN(P2_U3340) );
  AOI22_X1 U8699 ( .A1(n9093), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9488), .ZN(n6966) );
  OAI21_X1 U8700 ( .B1(n6967), .B2(n9494), .A(n6966), .ZN(P1_U3335) );
  NAND2_X1 U8701 ( .A1(n6968), .A2(n9945), .ZN(n6969) );
  OAI21_X1 U8702 ( .B1(n9945), .B2(n6805), .A(n6969), .ZN(P2_U3524) );
  INV_X1 U8703 ( .A(n6767), .ZN(n6980) );
  INV_X1 U8704 ( .A(n4877), .ZN(n6979) );
  NAND2_X1 U8705 ( .A1(n9769), .A2(n7989), .ZN(n6971) );
  NAND2_X1 U8706 ( .A1(n9779), .A2(n7901), .ZN(n6970) );
  NAND2_X1 U8707 ( .A1(n6971), .A2(n6970), .ZN(n6973) );
  XNOR2_X1 U8708 ( .A(n6973), .B(n4500), .ZN(n6974) );
  AOI22_X1 U8709 ( .A1(n7983), .A2(n9779), .B1(n7901), .B2(n9769), .ZN(n6975)
         );
  INV_X1 U8710 ( .A(n6974), .ZN(n6977) );
  INV_X1 U8711 ( .A(n6975), .ZN(n6976) );
  NAND2_X1 U8712 ( .A1(n6977), .A2(n6976), .ZN(n6978) );
  AND2_X1 U8713 ( .A1(n7133), .A2(n6978), .ZN(n6983) );
  NOR3_X1 U8714 ( .A1(n6980), .A2(n6979), .A3(n6983), .ZN(n6986) );
  INV_X1 U8715 ( .A(n6984), .ZN(n6985) );
  OAI21_X1 U8716 ( .B1(n6986), .B2(n6985), .A(n8744), .ZN(n6991) );
  INV_X1 U8717 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6987) );
  NOR2_X1 U8718 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6987), .ZN(n9608) );
  OAI22_X1 U8719 ( .A1(n6988), .A2(n8751), .B1(n8737), .B2(n7188), .ZN(n6989)
         );
  AOI211_X1 U8720 ( .C1(n8739), .C2(n9768), .A(n9608), .B(n6989), .ZN(n6990)
         );
  OAI211_X1 U8721 ( .C1(n8765), .C2(n6992), .A(n6991), .B(n6990), .ZN(P1_U3237) );
  OAI21_X1 U8722 ( .B1(n4922), .B2(n6084), .A(n6993), .ZN(n9731) );
  XNOR2_X1 U8723 ( .A(n6084), .B(n6994), .ZN(n6995) );
  NAND2_X1 U8724 ( .A1(n6995), .A2(n9706), .ZN(n9737) );
  OAI22_X1 U8725 ( .A1(n9737), .A2(n9241), .B1(n9338), .B2(n6996), .ZN(n7002)
         );
  AOI22_X1 U8726 ( .A1(n9347), .A2(n7862), .B1(n9335), .B2(n9748), .ZN(n7000)
         );
  OR2_X1 U8727 ( .A1(n9697), .A2(n9732), .ZN(n6997) );
  AND3_X1 U8728 ( .A1(n6998), .A2(n9695), .A3(n6997), .ZN(n9735) );
  AOI22_X1 U8729 ( .A1(n9321), .A2(n9735), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n9701), .ZN(n6999) );
  OAI211_X1 U8730 ( .C1(n10250), .C2(n9716), .A(n7000), .B(n6999), .ZN(n7001)
         );
  AOI211_X1 U8731 ( .C1(n9300), .C2(n9731), .A(n7002), .B(n7001), .ZN(n7003)
         );
  INV_X1 U8732 ( .A(n7003), .ZN(P1_U3289) );
  INV_X1 U8733 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7019) );
  NAND2_X1 U8734 ( .A1(n7868), .A2(n4645), .ZN(n7004) );
  NAND2_X1 U8735 ( .A1(n7005), .A2(n7004), .ZN(n7006) );
  OAI21_X1 U8736 ( .B1(n7006), .B2(n7009), .A(n7260), .ZN(n7457) );
  INV_X1 U8737 ( .A(n7457), .ZN(n7017) );
  NAND2_X1 U8738 ( .A1(n7007), .A2(n7008), .ZN(n7010) );
  XNOR2_X1 U8739 ( .A(n7010), .B(n7009), .ZN(n7012) );
  AOI21_X1 U8740 ( .B1(n7012), .B2(n9843), .A(n7011), .ZN(n7454) );
  AOI21_X1 U8741 ( .B1(n7013), .B2(n7015), .A(n9922), .ZN(n7014) );
  AND2_X1 U8742 ( .A1(n7340), .A2(n7014), .ZN(n7452) );
  AOI21_X1 U8743 ( .B1(n7015), .B2(n9886), .A(n7452), .ZN(n7016) );
  OAI211_X1 U8744 ( .C1(n7017), .C2(n8624), .A(n7454), .B(n7016), .ZN(n7020)
         );
  NAND2_X1 U8745 ( .A1(n7020), .A2(n9930), .ZN(n7018) );
  OAI21_X1 U8746 ( .B1(n9930), .B2(n7019), .A(n7018), .ZN(P2_U3466) );
  NAND2_X1 U8747 ( .A1(n7020), .A2(n9945), .ZN(n7021) );
  OAI21_X1 U8748 ( .B1(n9945), .B2(n6810), .A(n7021), .ZN(P2_U3525) );
  XNOR2_X1 U8749 ( .A(n7022), .B(n7024), .ZN(n9785) );
  NOR2_X1 U8750 ( .A1(n9241), .A2(n9784), .ZN(n7881) );
  INV_X1 U8751 ( .A(n7881), .ZN(n9350) );
  XNOR2_X1 U8752 ( .A(n7023), .B(n7024), .ZN(n9788) );
  NAND2_X1 U8753 ( .A1(n9788), .A2(n9300), .ZN(n7033) );
  AOI22_X1 U8754 ( .A1(n9208), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7137), .B2(
        n9701), .ZN(n7026) );
  NAND2_X1 U8755 ( .A1(n9335), .A2(n9778), .ZN(n7025) );
  OAI211_X1 U8756 ( .C1(n7027), .C2(n9338), .A(n7026), .B(n7025), .ZN(n7031)
         );
  INV_X1 U8757 ( .A(n7028), .ZN(n7029) );
  INV_X1 U8758 ( .A(n7124), .ZN(n9783) );
  OAI211_X1 U8759 ( .C1(n7029), .C2(n9783), .A(n9695), .B(n7094), .ZN(n9781)
         );
  NOR2_X1 U8760 ( .A1(n9781), .A2(n9344), .ZN(n7030) );
  AOI211_X1 U8761 ( .C1(n9347), .C2(n7124), .A(n7031), .B(n7030), .ZN(n7032)
         );
  OAI211_X1 U8762 ( .C1(n9785), .C2(n9350), .A(n7033), .B(n7032), .ZN(P1_U3284) );
  INV_X1 U8763 ( .A(n7034), .ZN(n7035) );
  AOI21_X1 U8764 ( .B1(n7037), .B2(n7036), .A(n7035), .ZN(n7043) );
  INV_X1 U8765 ( .A(n9831), .ZN(n7320) );
  INV_X1 U8766 ( .A(n7038), .ZN(n7288) );
  OAI21_X1 U8767 ( .B1(n9840), .B2(n7288), .A(n7039), .ZN(n7041) );
  OAI22_X1 U8768 ( .A1(n9832), .A2(n7258), .B1(n4645), .B2(n9829), .ZN(n7040)
         );
  AOI211_X1 U8769 ( .C1(n7320), .C2(n8175), .A(n7041), .B(n7040), .ZN(n7042)
         );
  OAI21_X1 U8770 ( .B1(n7043), .B2(n9826), .A(n7042), .ZN(P2_U3232) );
  INV_X1 U8771 ( .A(n7044), .ZN(n7140) );
  INV_X1 U8772 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10203) );
  INV_X1 U8773 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7051) );
  MUX2_X1 U8774 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n7051), .S(n9677), .Z(n9684)
         );
  INV_X1 U8775 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7046) );
  MUX2_X1 U8776 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7046), .S(n9668), .Z(n7049)
         );
  OAI21_X1 U8777 ( .B1(n7048), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7047), .ZN(
        n9671) );
  NAND2_X1 U8778 ( .A1(n7049), .A2(n9671), .ZN(n9670) );
  OR2_X1 U8779 ( .A1(n9668), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7050) );
  NAND2_X1 U8780 ( .A1(n9670), .A2(n7050), .ZN(n9683) );
  NAND2_X1 U8781 ( .A1(n9684), .A2(n9683), .ZN(n9682) );
  NAND2_X1 U8782 ( .A1(n7059), .A2(n7051), .ZN(n7052) );
  NAND2_X1 U8783 ( .A1(n9682), .A2(n7052), .ZN(n7194) );
  XOR2_X1 U8784 ( .A(n7202), .B(n7194), .Z(n7053) );
  NOR2_X1 U8785 ( .A1(n7053), .A2(n10203), .ZN(n7195) );
  AOI211_X1 U8786 ( .C1(n10203), .C2(n7053), .A(n9651), .B(n7195), .ZN(n7067)
         );
  INV_X1 U8787 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10070) );
  INV_X1 U8788 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7054) );
  XNOR2_X1 U8789 ( .A(n9668), .B(n7054), .ZN(n9664) );
  INV_X1 U8790 ( .A(n7055), .ZN(n7056) );
  NAND2_X1 U8791 ( .A1(n7057), .A2(n7056), .ZN(n9663) );
  NAND2_X1 U8792 ( .A1(n9664), .A2(n9663), .ZN(n9662) );
  NAND2_X1 U8793 ( .A1(n9668), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7058) );
  NAND2_X1 U8794 ( .A1(n9662), .A2(n7058), .ZN(n7060) );
  OR2_X1 U8795 ( .A1(n7060), .A2(n9677), .ZN(n7061) );
  XNOR2_X1 U8796 ( .A(n7060), .B(n7059), .ZN(n9681) );
  INV_X1 U8797 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9680) );
  NAND2_X1 U8798 ( .A1(n9681), .A2(n9680), .ZN(n9679) );
  NOR2_X1 U8799 ( .A1(n7062), .A2(n10070), .ZN(n7201) );
  AOI211_X1 U8800 ( .C1(n10070), .C2(n7062), .A(n9600), .B(n7201), .ZN(n7066)
         );
  INV_X1 U8801 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7064) );
  NAND2_X1 U8802 ( .A1(n9678), .A2(n7202), .ZN(n7063) );
  NAND2_X1 U8803 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8757) );
  OAI211_X1 U8804 ( .C1(n7064), .C2(n9691), .A(n7063), .B(n8757), .ZN(n7065)
         );
  OR3_X1 U8805 ( .A1(n7067), .A2(n7066), .A3(n7065), .ZN(P1_U3256) );
  INV_X1 U8806 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n10083) );
  AOI21_X1 U8807 ( .B1(n7076), .B2(P2_REG1_REG_10__SCAN_IN), .A(n7068), .ZN(
        n8208) );
  INV_X1 U8808 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7069) );
  MUX2_X1 U8809 ( .A(n7069), .B(P2_REG1_REG_11__SCAN_IN), .S(n8206), .Z(n8209)
         );
  NOR2_X1 U8810 ( .A1(n8208), .A2(n8209), .ZN(n8207) );
  AOI21_X1 U8811 ( .B1(n8206), .B2(P2_REG1_REG_11__SCAN_IN), .A(n8207), .ZN(
        n7072) );
  INV_X1 U8812 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7070) );
  MUX2_X1 U8813 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7070), .S(n7147), .Z(n7071)
         );
  NAND2_X1 U8814 ( .A1(n7072), .A2(n7071), .ZN(n7146) );
  OAI21_X1 U8815 ( .B1(n7072), .B2(n7071), .A(n7146), .ZN(n7073) );
  NAND2_X1 U8816 ( .A1(n8258), .A2(n7073), .ZN(n7074) );
  NAND2_X1 U8817 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(n8130), .ZN(n7675) );
  OAI211_X1 U8818 ( .C1(n8262), .C2(n10083), .A(n7074), .B(n7675), .ZN(n7083)
         );
  AOI21_X1 U8819 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7076), .A(n7075), .ZN(
        n8203) );
  INV_X1 U8820 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7078) );
  AOI22_X1 U8821 ( .A1(n8206), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7078), .B2(
        n7077), .ZN(n8202) );
  NAND2_X1 U8822 ( .A1(n8203), .A2(n8202), .ZN(n8201) );
  OAI21_X1 U8823 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n8206), .A(n8201), .ZN(
        n7081) );
  INV_X1 U8824 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7079) );
  MUX2_X1 U8825 ( .A(n7079), .B(P2_REG2_REG_12__SCAN_IN), .S(n7147), .Z(n7080)
         );
  NOR2_X1 U8826 ( .A1(n7081), .A2(n7080), .ZN(n7141) );
  AOI211_X1 U8827 ( .C1(n7081), .C2(n7080), .A(n8254), .B(n7141), .ZN(n7082)
         );
  AOI211_X1 U8828 ( .C1(n8256), .C2(n7147), .A(n7083), .B(n7082), .ZN(n7084)
         );
  INV_X1 U8829 ( .A(n7084), .ZN(P2_U3257) );
  AOI21_X1 U8830 ( .B1(n7085), .B2(n6150), .A(n9784), .ZN(n7087) );
  NAND2_X1 U8831 ( .A1(n7087), .A2(n7086), .ZN(n9800) );
  INV_X1 U8832 ( .A(n7088), .ZN(n7089) );
  AOI21_X1 U8833 ( .B1(n8982), .B2(n7090), .A(n7089), .ZN(n9806) );
  NAND2_X1 U8834 ( .A1(n9806), .A2(n9300), .ZN(n7099) );
  INV_X1 U8835 ( .A(n7190), .ZN(n7091) );
  OAI22_X1 U8836 ( .A1(n9716), .A2(n6480), .B1(n7091), .B2(n9301), .ZN(n7092)
         );
  AOI21_X1 U8837 ( .B1(n9335), .B2(n9792), .A(n7092), .ZN(n7093) );
  OAI21_X1 U8838 ( .B1(n7188), .B2(n9338), .A(n7093), .ZN(n7097) );
  AOI21_X1 U8839 ( .B1(n7094), .B2(n9796), .A(n9319), .ZN(n7095) );
  NAND2_X1 U8840 ( .A1(n7095), .A2(n7158), .ZN(n9798) );
  NOR2_X1 U8841 ( .A1(n9798), .A2(n9344), .ZN(n7096) );
  AOI211_X1 U8842 ( .C1(n9347), .C2(n9796), .A(n7097), .B(n7096), .ZN(n7098)
         );
  OAI211_X1 U8843 ( .C1(n9208), .C2(n9800), .A(n7099), .B(n7098), .ZN(P1_U3283) );
  OAI21_X1 U8844 ( .B1(n7102), .B2(n7101), .A(n7100), .ZN(n7107) );
  OAI22_X1 U8845 ( .A1(n9832), .A2(n7357), .B1(n9882), .B2(n9829), .ZN(n7106)
         );
  INV_X1 U8846 ( .A(n9840), .ZN(n8144) );
  NAND2_X1 U8847 ( .A1(n8144), .A2(n7344), .ZN(n7103) );
  OAI211_X1 U8848 ( .C1(n9831), .C2(n7258), .A(n7104), .B(n7103), .ZN(n7105)
         );
  AOI211_X1 U8849 ( .C1(n7107), .C2(n8138), .A(n7106), .B(n7105), .ZN(n7108)
         );
  INV_X1 U8850 ( .A(n7108), .ZN(P2_U3241) );
  XNOR2_X1 U8851 ( .A(n7110), .B(n7109), .ZN(n7115) );
  INV_X1 U8852 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7111) );
  OAI22_X1 U8853 ( .A1(n9840), .A2(n7273), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7111), .ZN(n7113) );
  OAI22_X1 U8854 ( .A1(n9832), .A2(n7506), .B1(n7356), .B2(n9829), .ZN(n7112)
         );
  AOI211_X1 U8855 ( .C1(n7320), .C2(n8172), .A(n7113), .B(n7112), .ZN(n7114)
         );
  OAI21_X1 U8856 ( .B1(n7115), .B2(n9826), .A(n7114), .ZN(P2_U3215) );
  INV_X1 U8857 ( .A(n7116), .ZN(n7117) );
  AOI21_X1 U8858 ( .B1(n8739), .B2(n9779), .A(n7117), .ZN(n7119) );
  NAND2_X1 U8859 ( .A1(n8767), .A2(n7124), .ZN(n7118) );
  OAI211_X1 U8860 ( .C1(n7300), .C2(n8737), .A(n7119), .B(n7118), .ZN(n7136)
         );
  NAND2_X1 U8861 ( .A1(n7124), .A2(n7989), .ZN(n7122) );
  NAND2_X1 U8862 ( .A1(n9793), .A2(n7901), .ZN(n7121) );
  NAND2_X1 U8863 ( .A1(n7122), .A2(n7121), .ZN(n7123) );
  XNOR2_X1 U8864 ( .A(n7123), .B(n4500), .ZN(n7127) );
  NAND2_X1 U8865 ( .A1(n7124), .A2(n7901), .ZN(n7126) );
  NAND2_X1 U8866 ( .A1(n7983), .A2(n9793), .ZN(n7125) );
  AND2_X1 U8867 ( .A1(n7126), .A2(n7125), .ZN(n7128) );
  NAND2_X1 U8868 ( .A1(n7127), .A2(n7128), .ZN(n7180) );
  INV_X1 U8869 ( .A(n7127), .ZN(n7130) );
  INV_X1 U8870 ( .A(n7128), .ZN(n7129) );
  NAND2_X1 U8871 ( .A1(n7130), .A2(n7129), .ZN(n7131) );
  AND2_X1 U8872 ( .A1(n7180), .A2(n7131), .ZN(n7132) );
  NAND3_X1 U8873 ( .A1(n6984), .A2(n7133), .A3(n4836), .ZN(n7134) );
  AOI21_X1 U8874 ( .B1(n7181), .B2(n7134), .A(n7995), .ZN(n7135) );
  AOI211_X1 U8875 ( .C1(n7137), .C2(n8749), .A(n7136), .B(n7135), .ZN(n7138)
         );
  INV_X1 U8876 ( .A(n7138), .ZN(P1_U3211) );
  OAI222_X1 U8877 ( .A1(P1_U3084), .A2(n9215), .B1(n9494), .B2(n7140), .C1(
        n7139), .C2(n9491), .ZN(P1_U3334) );
  NOR2_X1 U8878 ( .A1(n7611), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7142) );
  AOI21_X1 U8879 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n7611), .A(n7142), .ZN(
        n7143) );
  OAI21_X1 U8880 ( .B1(n7144), .B2(n7143), .A(n7602), .ZN(n7145) );
  NAND2_X1 U8881 ( .A1(n7145), .A2(n8253), .ZN(n7154) );
  INV_X1 U8882 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10116) );
  AOI22_X1 U8883 ( .A1(n7611), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n10116), .B2(
        n7155), .ZN(n7149) );
  OAI21_X1 U8884 ( .B1(n7147), .B2(P2_REG1_REG_12__SCAN_IN), .A(n7146), .ZN(
        n7148) );
  NAND2_X1 U8885 ( .A1(n7149), .A2(n7148), .ZN(n7610) );
  OAI21_X1 U8886 ( .B1(n7149), .B2(n7148), .A(n7610), .ZN(n7152) );
  AND2_X1 U8887 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7739) );
  INV_X1 U8888 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7150) );
  NOR2_X1 U8889 ( .A1(n8262), .A2(n7150), .ZN(n7151) );
  AOI211_X1 U8890 ( .C1(n8258), .C2(n7152), .A(n7739), .B(n7151), .ZN(n7153)
         );
  OAI211_X1 U8891 ( .C1(n7156), .C2(n7155), .A(n7154), .B(n7153), .ZN(P2_U3258) );
  XOR2_X1 U8892 ( .A(n7157), .B(n8983), .Z(n7226) );
  AOI211_X1 U8893 ( .C1(n7233), .C2(n7158), .A(n9319), .B(n7379), .ZN(n7224)
         );
  OAI22_X1 U8894 ( .A1(n7300), .A2(n9361), .B1(n7533), .B2(n9733), .ZN(n7159)
         );
  NOR2_X1 U8895 ( .A1(n7224), .A2(n7159), .ZN(n7162) );
  OAI211_X1 U8896 ( .C1(n7161), .C2(n8983), .A(n7160), .B(n9706), .ZN(n7221)
         );
  OAI211_X1 U8897 ( .C1(n7226), .C2(n9759), .A(n7162), .B(n7221), .ZN(n7167)
         );
  INV_X1 U8898 ( .A(n7233), .ZN(n7305) );
  INV_X1 U8899 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7163) );
  OAI22_X1 U8900 ( .A1(n9483), .A2(n7305), .B1(n9809), .B2(n7163), .ZN(n7164)
         );
  AOI21_X1 U8901 ( .B1(n7167), .B2(n9809), .A(n7164), .ZN(n7165) );
  INV_X1 U8902 ( .A(n7165), .ZN(P1_U3481) );
  OAI22_X1 U8903 ( .A1(n9439), .A2(n7305), .B1(n10189), .B2(n6639), .ZN(n7166)
         );
  AOI21_X1 U8904 ( .B1(n7167), .B2(n10189), .A(n7166), .ZN(n7168) );
  INV_X1 U8905 ( .A(n7168), .ZN(P1_U3532) );
  XNOR2_X1 U8906 ( .A(n7170), .B(n7169), .ZN(n7176) );
  INV_X1 U8907 ( .A(n7171), .ZN(n7365) );
  OAI21_X1 U8908 ( .B1(n9840), .B2(n7365), .A(n7172), .ZN(n7174) );
  OAI22_X1 U8909 ( .A1(n9832), .A2(n9830), .B1(n9892), .B2(n9829), .ZN(n7173)
         );
  AOI211_X1 U8910 ( .C1(n7320), .C2(n8171), .A(n7174), .B(n7173), .ZN(n7175)
         );
  OAI21_X1 U8911 ( .B1(n7176), .B2(n9826), .A(n7175), .ZN(P2_U3223) );
  NAND2_X1 U8912 ( .A1(n9796), .A2(n7989), .ZN(n7178) );
  NAND2_X1 U8913 ( .A1(n9778), .A2(n7901), .ZN(n7177) );
  NAND2_X1 U8914 ( .A1(n7178), .A2(n7177), .ZN(n7179) );
  XNOR2_X1 U8915 ( .A(n7179), .B(n7986), .ZN(n7227) );
  AND2_X1 U8916 ( .A1(n7983), .A2(n9778), .ZN(n7182) );
  AOI21_X1 U8917 ( .B1(n9796), .B2(n7901), .A(n7182), .ZN(n7184) );
  NAND2_X1 U8918 ( .A1(n7293), .A2(n7228), .ZN(n7185) );
  XOR2_X1 U8919 ( .A(n7227), .B(n7185), .Z(n7193) );
  NAND2_X1 U8920 ( .A1(n8762), .A2(n9792), .ZN(n7187) );
  OAI211_X1 U8921 ( .C1(n7188), .C2(n8759), .A(n7187), .B(n7186), .ZN(n7189)
         );
  AOI21_X1 U8922 ( .B1(n8749), .B2(n7190), .A(n7189), .ZN(n7192) );
  NAND2_X1 U8923 ( .A1(n8730), .A2(n9796), .ZN(n7191) );
  OAI211_X1 U8924 ( .C1(n7193), .C2(n7995), .A(n7192), .B(n7191), .ZN(P1_U3219) );
  INV_X1 U8925 ( .A(n7194), .ZN(n7196) );
  AOI21_X1 U8926 ( .B1(n7196), .B2(n7202), .A(n7195), .ZN(n7199) );
  INV_X1 U8927 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7197) );
  MUX2_X1 U8928 ( .A(n7197), .B(P1_REG1_REG_16__SCAN_IN), .S(n9071), .Z(n7198)
         );
  NOR2_X1 U8929 ( .A1(n7199), .A2(n7198), .ZN(n9067) );
  AOI211_X1 U8930 ( .C1(n7199), .C2(n7198), .A(n9067), .B(n9651), .ZN(n7212)
         );
  INV_X1 U8931 ( .A(n7200), .ZN(n7203) );
  INV_X1 U8932 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7204) );
  MUX2_X1 U8933 ( .A(n7204), .B(P1_REG2_REG_16__SCAN_IN), .S(n9071), .Z(n7205)
         );
  NOR2_X1 U8934 ( .A1(n7206), .A2(n7205), .ZN(n9070) );
  AOI211_X1 U8935 ( .C1(n7206), .C2(n7205), .A(n9070), .B(n9600), .ZN(n7211)
         );
  INV_X1 U8936 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7209) );
  NAND2_X1 U8937 ( .A1(n9678), .A2(n9071), .ZN(n7208) );
  NAND2_X1 U8938 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n7207) );
  OAI211_X1 U8939 ( .C1(n7209), .C2(n9691), .A(n7208), .B(n7207), .ZN(n7210)
         );
  OR3_X1 U8940 ( .A1(n7212), .A2(n7211), .A3(n7210), .ZN(P1_U3257) );
  INV_X1 U8941 ( .A(n7213), .ZN(n7306) );
  OAI222_X1 U8942 ( .A1(n8954), .A2(P1_U3084), .B1(n9494), .B2(n7306), .C1(
        n10219), .C2(n9491), .ZN(P1_U3332) );
  INV_X1 U8943 ( .A(n7214), .ZN(n7309) );
  OAI222_X1 U8944 ( .A1(n6348), .A2(P1_U3084), .B1(n9494), .B2(n7309), .C1(
        n7215), .C2(n9491), .ZN(P1_U3333) );
  INV_X1 U8945 ( .A(n7302), .ZN(n7216) );
  OAI22_X1 U8946 ( .A1(n9716), .A2(n7217), .B1(n7216), .B2(n9301), .ZN(n7219)
         );
  NOR2_X1 U8947 ( .A1(n9338), .A2(n7300), .ZN(n7218) );
  AOI211_X1 U8948 ( .C1(n9335), .C2(n9043), .A(n7219), .B(n7218), .ZN(n7220)
         );
  OAI21_X1 U8949 ( .B1(n7305), .B2(n9326), .A(n7220), .ZN(n7223) );
  NOR2_X1 U8950 ( .A1(n7221), .A2(n9241), .ZN(n7222) );
  AOI211_X1 U8951 ( .C1(n7224), .C2(n9321), .A(n7223), .B(n7222), .ZN(n7225)
         );
  OAI21_X1 U8952 ( .B1(n9333), .B2(n7226), .A(n7225), .ZN(P1_U3282) );
  NAND2_X1 U8953 ( .A1(n7228), .A2(n7227), .ZN(n7294) );
  NAND2_X1 U8954 ( .A1(n7233), .A2(n7989), .ZN(n7230) );
  NAND2_X1 U8955 ( .A1(n9792), .A2(n7901), .ZN(n7229) );
  NAND2_X1 U8956 ( .A1(n7230), .A2(n7229), .ZN(n7231) );
  XNOR2_X1 U8957 ( .A(n7231), .B(n4500), .ZN(n7234) );
  AND2_X1 U8958 ( .A1(n7983), .A2(n9792), .ZN(n7232) );
  AOI21_X1 U8959 ( .B1(n7233), .B2(n7901), .A(n7232), .ZN(n7235) );
  NAND2_X1 U8960 ( .A1(n7234), .A2(n7235), .ZN(n7239) );
  INV_X1 U8961 ( .A(n7234), .ZN(n7237) );
  INV_X1 U8962 ( .A(n7235), .ZN(n7236) );
  NAND2_X1 U8963 ( .A1(n7237), .A2(n7236), .ZN(n7238) );
  AND2_X1 U8964 ( .A1(n7239), .A2(n7238), .ZN(n7297) );
  NAND2_X1 U8965 ( .A1(n7392), .A2(n7989), .ZN(n7242) );
  NAND2_X1 U8966 ( .A1(n9043), .A2(n7901), .ZN(n7241) );
  NAND2_X1 U8967 ( .A1(n7242), .A2(n7241), .ZN(n7243) );
  XNOR2_X1 U8968 ( .A(n7243), .B(n7986), .ZN(n7246) );
  NAND2_X1 U8969 ( .A1(n7392), .A2(n7901), .ZN(n7245) );
  NAND2_X1 U8970 ( .A1(n7983), .A2(n9043), .ZN(n7244) );
  NAND2_X1 U8971 ( .A1(n7245), .A2(n7244), .ZN(n7247) );
  NAND2_X1 U8972 ( .A1(n7246), .A2(n7247), .ZN(n7520) );
  INV_X1 U8973 ( .A(n7246), .ZN(n7249) );
  INV_X1 U8974 ( .A(n7247), .ZN(n7248) );
  NAND2_X1 U8975 ( .A1(n7249), .A2(n7248), .ZN(n7522) );
  NAND2_X1 U8976 ( .A1(n7520), .A2(n7522), .ZN(n7250) );
  XNOR2_X1 U8977 ( .A(n7240), .B(n7250), .ZN(n7257) );
  INV_X1 U8978 ( .A(n7251), .ZN(n7390) );
  NOR2_X1 U8979 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7252), .ZN(n9636) );
  AOI21_X1 U8980 ( .B1(n8739), .B2(n9792), .A(n9636), .ZN(n7254) );
  NAND2_X1 U8981 ( .A1(n8762), .A2(n9042), .ZN(n7253) );
  OAI211_X1 U8982 ( .C1(n8765), .C2(n7390), .A(n7254), .B(n7253), .ZN(n7255)
         );
  AOI21_X1 U8983 ( .B1(n7392), .B2(n8767), .A(n7255), .ZN(n7256) );
  OAI21_X1 U8984 ( .B1(n7257), .B2(n7995), .A(n7256), .ZN(P1_U3215) );
  NAND2_X1 U8985 ( .A1(n7258), .A2(n7449), .ZN(n7259) );
  XNOR2_X1 U8986 ( .A(n7355), .B(n7354), .ZN(n9891) );
  INV_X1 U8987 ( .A(n9891), .ZN(n7282) );
  NOR2_X1 U8988 ( .A1(n7262), .A2(n7261), .ZN(n7272) );
  NAND2_X1 U8989 ( .A1(n7272), .A2(n7263), .ZN(n7265) );
  OR2_X1 U8990 ( .A1(n7266), .A2(n7451), .ZN(n7371) );
  NAND2_X1 U8991 ( .A1(n8508), .A2(n7371), .ZN(n7267) );
  INV_X1 U8992 ( .A(n7268), .ZN(n7269) );
  NOR2_X1 U8993 ( .A1(n7270), .A2(n5050), .ZN(n7271) );
  NAND2_X1 U8994 ( .A1(n7272), .A2(n7271), .ZN(n9855) );
  NAND2_X1 U8995 ( .A1(n7341), .A2(n7356), .ZN(n7367) );
  OAI21_X1 U8996 ( .B1(n7341), .B2(n7356), .A(n7367), .ZN(n9889) );
  OAI22_X1 U8997 ( .A1(n8551), .A2(n9889), .B1(n7273), .B2(n8344), .ZN(n7274)
         );
  AOI21_X1 U8998 ( .B1(n9847), .B2(n9885), .A(n7274), .ZN(n7281) );
  XNOR2_X1 U8999 ( .A(n7275), .B(n4978), .ZN(n7278) );
  OAI22_X1 U9000 ( .A1(n7276), .A2(n8502), .B1(n7506), .B2(n8500), .ZN(n7277)
         );
  AOI21_X1 U9001 ( .B1(n7278), .B2(n9843), .A(n7277), .ZN(n9888) );
  MUX2_X1 U9002 ( .A(n7279), .B(n9888), .S(n8549), .Z(n7280) );
  OAI211_X1 U9003 ( .C1(n7282), .C2(n8543), .A(n7281), .B(n7280), .ZN(P2_U3289) );
  INV_X1 U9004 ( .A(n8543), .ZN(n9857) );
  INV_X1 U9005 ( .A(n7283), .ZN(n7284) );
  OAI22_X1 U9006 ( .A1(n9860), .A2(n7285), .B1(n8551), .B2(n7284), .ZN(n7286)
         );
  AOI21_X1 U9007 ( .B1(n9857), .B2(n7287), .A(n7286), .ZN(n7292) );
  OAI22_X1 U9008 ( .A1(n8549), .A2(n6798), .B1(n7288), .B2(n8344), .ZN(n7289)
         );
  AOI21_X1 U9009 ( .B1(n9847), .B2(n7290), .A(n7289), .ZN(n7291) );
  NAND2_X1 U9010 ( .A1(n7292), .A2(n7291), .ZN(P2_U3292) );
  AND2_X1 U9011 ( .A1(n7294), .A2(n7293), .ZN(n7296) );
  OAI21_X1 U9012 ( .B1(n7297), .B2(n7296), .A(n7295), .ZN(n7298) );
  NAND2_X1 U9013 ( .A1(n7298), .A2(n8744), .ZN(n7304) );
  NAND2_X1 U9014 ( .A1(n8762), .A2(n9043), .ZN(n7299) );
  NAND2_X1 U9015 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9621) );
  OAI211_X1 U9016 ( .C1(n7300), .C2(n8759), .A(n7299), .B(n9621), .ZN(n7301)
         );
  AOI21_X1 U9017 ( .B1(n8749), .B2(n7302), .A(n7301), .ZN(n7303) );
  OAI211_X1 U9018 ( .C1(n7305), .C2(n8751), .A(n7304), .B(n7303), .ZN(P1_U3229) );
  INV_X1 U9019 ( .A(n7312), .ZN(n7314) );
  NOR2_X1 U9020 ( .A1(n7314), .A2(n7313), .ZN(n7315) );
  XNOR2_X1 U9021 ( .A(n7316), .B(n7315), .ZN(n7322) );
  OAI21_X1 U9022 ( .B1(n9840), .B2(n7511), .A(n7317), .ZN(n7319) );
  OAI22_X1 U9023 ( .A1(n9832), .A2(n7703), .B1(n9899), .B2(n9829), .ZN(n7318)
         );
  AOI211_X1 U9024 ( .C1(n7320), .C2(n8170), .A(n7319), .B(n7318), .ZN(n7321)
         );
  OAI21_X1 U9025 ( .B1(n7322), .B2(n9826), .A(n7321), .ZN(P2_U3233) );
  OAI21_X1 U9026 ( .B1(n7325), .B2(n7324), .A(n7323), .ZN(n7326) );
  AOI222_X1 U9027 ( .A1(n9843), .A2(n7326), .B1(n8174), .B2(n8533), .C1(n8176), 
        .C2(n8530), .ZN(n9876) );
  INV_X1 U9028 ( .A(n9876), .ZN(n7331) );
  OAI22_X1 U9029 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(n8344), .B1(n8549), .B2(
        n10028), .ZN(n7330) );
  NOR2_X1 U9030 ( .A1(n9855), .A2(n9875), .ZN(n7329) );
  AOI211_X1 U9031 ( .C1(n7331), .C2(n8549), .A(n7330), .B(n7329), .ZN(n7336)
         );
  OAI21_X1 U9032 ( .B1(n7334), .B2(n7333), .A(n7332), .ZN(n9878) );
  NAND2_X1 U9033 ( .A1(n9857), .A2(n9878), .ZN(n7335) );
  OAI21_X1 U9034 ( .B1(n7351), .B2(n7338), .A(n7337), .ZN(n7339) );
  AOI222_X1 U9035 ( .A1(n9843), .A2(n7339), .B1(n8171), .B2(n8533), .C1(n8173), 
        .C2(n8530), .ZN(n9881) );
  INV_X1 U9036 ( .A(n7340), .ZN(n7343) );
  INV_X1 U9037 ( .A(n7341), .ZN(n7342) );
  OAI211_X1 U9038 ( .C1(n9882), .C2(n7343), .A(n7342), .B(n9853), .ZN(n9880)
         );
  INV_X1 U9039 ( .A(n7344), .ZN(n7345) );
  OAI22_X1 U9040 ( .A1(n9855), .A2(n9880), .B1(n7345), .B2(n8344), .ZN(n7348)
         );
  INV_X1 U9041 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7346) );
  NOR2_X1 U9042 ( .A1(n8549), .A2(n7346), .ZN(n7347) );
  AOI211_X1 U9043 ( .C1(n9847), .C2(n7349), .A(n7348), .B(n7347), .ZN(n7353)
         );
  XOR2_X1 U9044 ( .A(n7351), .B(n7350), .Z(n9884) );
  NAND2_X1 U9045 ( .A1(n9884), .A2(n9857), .ZN(n7352) );
  OAI211_X1 U9046 ( .C1(n9881), .C2(n9860), .A(n7353), .B(n7352), .ZN(P2_U3290) );
  NAND2_X1 U9047 ( .A1(n7357), .A2(n7356), .ZN(n7358) );
  NAND2_X1 U9048 ( .A1(n7359), .A2(n7358), .ZN(n7490) );
  XNOR2_X1 U9049 ( .A(n7490), .B(n7492), .ZN(n9895) );
  INV_X1 U9050 ( .A(n8508), .ZN(n7510) );
  OAI21_X1 U9051 ( .B1(n7491), .B2(n7360), .A(n7503), .ZN(n7361) );
  NAND2_X1 U9052 ( .A1(n7361), .A2(n9843), .ZN(n7363) );
  AOI22_X1 U9053 ( .A1(n8171), .A2(n8530), .B1(n8533), .B2(n8169), .ZN(n7362)
         );
  NAND2_X1 U9054 ( .A1(n7363), .A2(n7362), .ZN(n7364) );
  AOI21_X1 U9055 ( .B1(n9895), .B2(n7510), .A(n7364), .ZN(n9897) );
  INV_X1 U9056 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7366) );
  OAI22_X1 U9057 ( .A1(n8549), .A2(n7366), .B1(n7365), .B2(n8344), .ZN(n7370)
         );
  NAND2_X1 U9058 ( .A1(n7367), .A2(n7494), .ZN(n7368) );
  NAND2_X1 U9059 ( .A1(n7513), .A2(n7368), .ZN(n9893) );
  NOR2_X1 U9060 ( .A1(n8551), .A2(n9893), .ZN(n7369) );
  AOI211_X1 U9061 ( .C1(n9847), .C2(n7494), .A(n7370), .B(n7369), .ZN(n7374)
         );
  INV_X1 U9062 ( .A(n7371), .ZN(n7372) );
  AND2_X1 U9063 ( .A1(n8549), .A2(n7372), .ZN(n8521) );
  NAND2_X1 U9064 ( .A1(n9895), .A2(n8521), .ZN(n7373) );
  OAI211_X1 U9065 ( .C1(n9897), .C2(n9860), .A(n7374), .B(n7373), .ZN(P2_U3288) );
  OAI21_X1 U9066 ( .B1(n4427), .B2(n6175), .A(n7375), .ZN(n7401) );
  OAI211_X1 U9067 ( .C1(n7378), .C2(n7377), .A(n7376), .B(n9706), .ZN(n7398)
         );
  AOI22_X1 U9068 ( .A1(n9794), .A2(n9792), .B1(n9042), .B2(n9791), .ZN(n7380)
         );
  OAI211_X1 U9069 ( .C1(n7379), .C2(n7385), .A(n9695), .B(n7484), .ZN(n7389)
         );
  NAND3_X1 U9070 ( .A1(n7398), .A2(n7380), .A3(n7389), .ZN(n7381) );
  AOI21_X1 U9071 ( .B1(n7401), .B2(n9789), .A(n7381), .ZN(n7388) );
  INV_X1 U9072 ( .A(n9439), .ZN(n7382) );
  AOI22_X1 U9073 ( .A1(n7382), .A2(n7392), .B1(n10187), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7383) );
  OAI21_X1 U9074 ( .B1(n7388), .B2(n10187), .A(n7383), .ZN(P1_U3533) );
  INV_X1 U9075 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7384) );
  OAI22_X1 U9076 ( .A1(n7385), .A2(n9483), .B1(n9809), .B2(n7384), .ZN(n7386)
         );
  INV_X1 U9077 ( .A(n7386), .ZN(n7387) );
  OAI21_X1 U9078 ( .B1(n7388), .B2(n9807), .A(n7387), .ZN(P1_U3484) );
  OR2_X1 U9079 ( .A1(n7389), .A2(n9344), .ZN(n7397) );
  OAI22_X1 U9080 ( .A1(n9716), .A2(n6647), .B1(n7390), .B2(n9301), .ZN(n7391)
         );
  AOI21_X1 U9081 ( .B1(n9335), .B2(n9042), .A(n7391), .ZN(n7396) );
  NAND2_X1 U9082 ( .A1(n9347), .A2(n7392), .ZN(n7395) );
  OR2_X1 U9083 ( .A1(n9338), .A2(n7393), .ZN(n7394) );
  NAND4_X1 U9084 ( .A1(n7397), .A2(n7396), .A3(n7395), .A4(n7394), .ZN(n7400)
         );
  NOR2_X1 U9085 ( .A1(n7398), .A2(n9241), .ZN(n7399) );
  AOI211_X1 U9086 ( .C1(n9300), .C2(n7401), .A(n7400), .B(n7399), .ZN(n7402)
         );
  INV_X1 U9087 ( .A(n7402), .ZN(P1_U3281) );
  INV_X1 U9088 ( .A(n7403), .ZN(n7406) );
  OAI222_X1 U9089 ( .A1(P1_U3084), .A2(n7407), .B1(n9494), .B2(n7406), .C1(
        n7405), .C2(n9491), .ZN(P1_U3331) );
  NAND2_X1 U9090 ( .A1(n7408), .A2(n8017), .ZN(n9873) );
  INV_X1 U9091 ( .A(n9873), .ZN(n7414) );
  AOI22_X1 U9092 ( .A1(n9873), .A2(n9843), .B1(n8533), .B2(n7409), .ZN(n9869)
         );
  NAND2_X1 U9093 ( .A1(n9845), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7410) );
  AOI21_X1 U9094 ( .B1(n9869), .B2(n7410), .A(n9860), .ZN(n7411) );
  AOI21_X1 U9095 ( .B1(n9860), .B2(P2_REG2_REG_0__SCAN_IN), .A(n7411), .ZN(
        n7413) );
  OAI21_X1 U9096 ( .B1(n9847), .B2(n8520), .A(n8020), .ZN(n7412) );
  OAI211_X1 U9097 ( .C1(n7414), .C2(n8543), .A(n7413), .B(n7412), .ZN(P2_U3296) );
  INV_X1 U9098 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10286) );
  NOR2_X1 U9099 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7415) );
  AOI21_X1 U9100 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7415), .ZN(n9952) );
  NOR2_X1 U9101 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7416) );
  AOI21_X1 U9102 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7416), .ZN(n9955) );
  NOR2_X1 U9103 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7417) );
  AOI21_X1 U9104 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7417), .ZN(n9958) );
  NOR2_X1 U9105 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(P2_ADDR_REG_14__SCAN_IN), 
        .ZN(n7418) );
  AOI21_X1 U9106 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n7418), .ZN(n9961) );
  NOR2_X1 U9107 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .ZN(n7419) );
  AOI21_X1 U9108 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n7419), .ZN(n9964) );
  NOR2_X1 U9109 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(P1_ADDR_REG_4__SCAN_IN), 
        .ZN(n7425) );
  INV_X1 U9110 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9586) );
  AOI22_X1 U9111 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n9586), .B1(
        P1_ADDR_REG_4__SCAN_IN), .B2(n10107), .ZN(n10297) );
  NAND2_X1 U9112 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7423) );
  XNOR2_X1 U9113 ( .A(n9507), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(n10295) );
  NAND2_X1 U9114 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7421) );
  XOR2_X1 U9115 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10293) );
  AOI21_X1 U9116 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9946) );
  INV_X1 U9117 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10233) );
  NAND3_X1 U9118 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9948) );
  OAI21_X1 U9119 ( .B1(n9946), .B2(n10233), .A(n9948), .ZN(n10292) );
  NAND2_X1 U9120 ( .A1(n10293), .A2(n10292), .ZN(n7420) );
  NAND2_X1 U9121 ( .A1(n7421), .A2(n7420), .ZN(n10294) );
  NAND2_X1 U9122 ( .A1(n10295), .A2(n10294), .ZN(n7422) );
  NAND2_X1 U9123 ( .A1(n7423), .A2(n7422), .ZN(n10296) );
  NOR2_X1 U9124 ( .A1(n10297), .A2(n10296), .ZN(n7424) );
  NOR2_X1 U9125 ( .A1(n7425), .A2(n7424), .ZN(n7426) );
  NOR2_X1 U9126 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7426), .ZN(n10280) );
  AND2_X1 U9127 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7426), .ZN(n10281) );
  NOR2_X1 U9128 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10281), .ZN(n7427) );
  NOR2_X1 U9129 ( .A1(n10280), .A2(n7427), .ZN(n7429) );
  NAND2_X1 U9130 ( .A1(n7429), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7431) );
  XNOR2_X1 U9131 ( .A(n7429), .B(n7428), .ZN(n10279) );
  NAND2_X1 U9132 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n10279), .ZN(n7430) );
  NAND2_X1 U9133 ( .A1(n7431), .A2(n7430), .ZN(n7432) );
  NAND2_X1 U9134 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7432), .ZN(n7435) );
  XNOR2_X1 U9135 ( .A(n7433), .B(n7432), .ZN(n10283) );
  NAND2_X1 U9136 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10283), .ZN(n7434) );
  NAND2_X1 U9137 ( .A1(n7435), .A2(n7434), .ZN(n7436) );
  NAND2_X1 U9138 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7436), .ZN(n7438) );
  XOR2_X1 U9139 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7436), .Z(n10291) );
  NAND2_X1 U9140 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10291), .ZN(n7437) );
  NAND2_X1 U9141 ( .A1(n7438), .A2(n7437), .ZN(n7439) );
  AND2_X1 U9142 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7439), .ZN(n7441) );
  INV_X1 U9143 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10290) );
  XOR2_X1 U9144 ( .A(n7440), .B(n7439), .Z(n10289) );
  NAND2_X1 U9145 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7442) );
  OAI21_X1 U9146 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n7442), .ZN(n9972) );
  NAND2_X1 U9147 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7443) );
  OAI21_X1 U9148 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7443), .ZN(n9969) );
  AOI21_X1 U9149 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9968), .ZN(n9967) );
  NOR2_X1 U9150 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7444) );
  AOI21_X1 U9151 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7444), .ZN(n9966) );
  NAND2_X1 U9152 ( .A1(n9967), .A2(n9966), .ZN(n9965) );
  OAI21_X1 U9153 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9965), .ZN(n9963) );
  NAND2_X1 U9154 ( .A1(n9964), .A2(n9963), .ZN(n9962) );
  OAI21_X1 U9155 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9962), .ZN(n9960) );
  NAND2_X1 U9156 ( .A1(n9961), .A2(n9960), .ZN(n9959) );
  OAI21_X1 U9157 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9959), .ZN(n9957) );
  NAND2_X1 U9158 ( .A1(n9958), .A2(n9957), .ZN(n9956) );
  OAI21_X1 U9159 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9956), .ZN(n9954) );
  NAND2_X1 U9160 ( .A1(n9955), .A2(n9954), .ZN(n9953) );
  OAI21_X1 U9161 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9953), .ZN(n9951) );
  NAND2_X1 U9162 ( .A1(n9952), .A2(n9951), .ZN(n9950) );
  OAI21_X1 U9163 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9950), .ZN(n10285) );
  NOR2_X1 U9164 ( .A1(n10286), .A2(n10285), .ZN(n7445) );
  NAND2_X1 U9165 ( .A1(n10286), .A2(n10285), .ZN(n10284) );
  OAI21_X1 U9166 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7445), .A(n10284), .ZN(
        n7447) );
  XNOR2_X1 U9167 ( .A(n4912), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7446) );
  XNOR2_X1 U9168 ( .A(n7447), .B(n7446), .ZN(ADD_1071_U4) );
  INV_X1 U9169 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7448) );
  OAI22_X1 U9170 ( .A1(n8496), .A2(n7449), .B1(n7448), .B2(n8549), .ZN(n7456)
         );
  AOI22_X1 U9171 ( .A1(n7452), .A2(n7451), .B1(n9845), .B2(n7450), .ZN(n7453)
         );
  AOI21_X1 U9172 ( .B1(n7454), .B2(n7453), .A(n9860), .ZN(n7455) );
  AOI211_X1 U9173 ( .C1(n9857), .C2(n7457), .A(n7456), .B(n7455), .ZN(n7458)
         );
  INV_X1 U9174 ( .A(n7458), .ZN(P2_U3291) );
  INV_X1 U9175 ( .A(n7459), .ZN(n7460) );
  OAI21_X1 U9176 ( .B1(n7477), .B2(n7460), .A(n8872), .ZN(n7461) );
  XNOR2_X1 U9177 ( .A(n7461), .B(n8965), .ZN(n7462) );
  NAND2_X1 U9178 ( .A1(n7462), .A2(n9706), .ZN(n7621) );
  AND2_X1 U9179 ( .A1(n7463), .A2(n8965), .ZN(n7464) );
  NOR2_X1 U9180 ( .A1(n7465), .A2(n7464), .ZN(n7623) );
  NAND2_X1 U9181 ( .A1(n7482), .A2(n7618), .ZN(n7466) );
  NAND2_X1 U9182 ( .A1(n7466), .A2(n9695), .ZN(n7467) );
  OR2_X1 U9183 ( .A1(n7467), .A2(n7552), .ZN(n7619) );
  AOI22_X1 U9184 ( .A1(n9208), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7587), .B2(
        n9701), .ZN(n7469) );
  NAND2_X1 U9185 ( .A1(n9335), .A2(n9040), .ZN(n7468) );
  OAI211_X1 U9186 ( .C1(n7470), .C2(n9338), .A(n7469), .B(n7468), .ZN(n7471)
         );
  AOI21_X1 U9187 ( .B1(n7618), .B2(n9347), .A(n7471), .ZN(n7472) );
  OAI21_X1 U9188 ( .B1(n7619), .B2(n9344), .A(n7472), .ZN(n7473) );
  AOI21_X1 U9189 ( .B1(n7623), .B2(n9300), .A(n7473), .ZN(n7474) );
  OAI21_X1 U9190 ( .B1(n9241), .B2(n7621), .A(n7474), .ZN(P1_U3279) );
  OAI21_X1 U9191 ( .B1(n7476), .B2(n8986), .A(n7475), .ZN(n7478) );
  INV_X1 U9192 ( .A(n7478), .ZN(n9556) );
  XNOR2_X1 U9193 ( .A(n7477), .B(n4947), .ZN(n7481) );
  INV_X1 U9194 ( .A(n9712), .ZN(n9805) );
  NAND2_X1 U9195 ( .A1(n7478), .A2(n9805), .ZN(n7480) );
  AOI22_X1 U9196 ( .A1(n9794), .A2(n9043), .B1(n9041), .B2(n9791), .ZN(n7479)
         );
  OAI211_X1 U9197 ( .C1(n9784), .C2(n7481), .A(n7480), .B(n7479), .ZN(n9551)
         );
  NAND2_X1 U9198 ( .A1(n9551), .A2(n9716), .ZN(n7488) );
  INV_X1 U9199 ( .A(n7482), .ZN(n7483) );
  AOI211_X1 U9200 ( .C1(n9553), .C2(n7484), .A(n9319), .B(n7483), .ZN(n9552)
         );
  INV_X1 U9201 ( .A(n9553), .ZN(n7538) );
  AOI22_X1 U9202 ( .A1(n9208), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7535), .B2(
        n9701), .ZN(n7485) );
  OAI21_X1 U9203 ( .B1(n7538), .B2(n9326), .A(n7485), .ZN(n7486) );
  AOI21_X1 U9204 ( .B1(n9552), .B2(n9321), .A(n7486), .ZN(n7487) );
  OAI211_X1 U9205 ( .C1(n9556), .C2(n7489), .A(n7488), .B(n7487), .ZN(P1_U3280) );
  INV_X1 U9206 ( .A(n7490), .ZN(n7493) );
  NAND2_X1 U9207 ( .A1(n8170), .A2(n7494), .ZN(n7496) );
  INV_X1 U9208 ( .A(n7498), .ZN(n7502) );
  AND2_X1 U9209 ( .A1(n7496), .A2(n7502), .ZN(n7495) );
  NAND2_X1 U9210 ( .A1(n7497), .A2(n7496), .ZN(n7499) );
  NAND2_X1 U9211 ( .A1(n7499), .A2(n7498), .ZN(n7500) );
  NAND2_X1 U9212 ( .A1(n7559), .A2(n7500), .ZN(n9902) );
  NAND3_X1 U9213 ( .A1(n7503), .A2(n7502), .A3(n7501), .ZN(n7504) );
  AOI21_X1 U9214 ( .B1(n7505), .B2(n7504), .A(n8488), .ZN(n7508) );
  OAI22_X1 U9215 ( .A1(n7506), .A2(n8502), .B1(n7703), .B2(n8500), .ZN(n7507)
         );
  OR2_X1 U9216 ( .A1(n7508), .A2(n7507), .ZN(n7509) );
  AOI21_X1 U9217 ( .B1(n9902), .B2(n7510), .A(n7509), .ZN(n9904) );
  OAI22_X1 U9218 ( .A1(n8549), .A2(n7512), .B1(n7511), .B2(n8344), .ZN(n7516)
         );
  AND2_X1 U9219 ( .A1(n7513), .A2(n7517), .ZN(n7514) );
  OR2_X1 U9220 ( .A1(n7514), .A2(n7568), .ZN(n9900) );
  NOR2_X1 U9221 ( .A1(n9900), .A2(n8551), .ZN(n7515) );
  AOI211_X1 U9222 ( .C1(n9847), .C2(n7517), .A(n7516), .B(n7515), .ZN(n7519)
         );
  NAND2_X1 U9223 ( .A1(n9902), .A2(n8521), .ZN(n7518) );
  OAI211_X1 U9224 ( .C1(n9904), .C2(n9860), .A(n7519), .B(n7518), .ZN(P2_U3287) );
  NAND2_X1 U9225 ( .A1(n9553), .A2(n7989), .ZN(n7524) );
  NAND2_X1 U9226 ( .A1(n9042), .A2(n5005), .ZN(n7523) );
  NAND2_X1 U9227 ( .A1(n7524), .A2(n7523), .ZN(n7525) );
  XNOR2_X1 U9228 ( .A(n7525), .B(n4500), .ZN(n7575) );
  AND2_X1 U9229 ( .A1(n7983), .A2(n9042), .ZN(n7526) );
  AOI21_X1 U9230 ( .B1(n9553), .B2(n7901), .A(n7526), .ZN(n7576) );
  XNOR2_X1 U9231 ( .A(n7575), .B(n7576), .ZN(n7528) );
  AOI21_X1 U9232 ( .B1(n7527), .B2(n7528), .A(n7995), .ZN(n7530) );
  INV_X1 U9233 ( .A(n7528), .ZN(n7529) );
  NAND2_X1 U9234 ( .A1(n7530), .A2(n7580), .ZN(n7537) );
  NAND2_X1 U9235 ( .A1(n8762), .A2(n9041), .ZN(n7532) );
  AND2_X1 U9236 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9644) );
  INV_X1 U9237 ( .A(n9644), .ZN(n7531) );
  OAI211_X1 U9238 ( .C1(n7533), .C2(n8759), .A(n7532), .B(n7531), .ZN(n7534)
         );
  AOI21_X1 U9239 ( .B1(n8749), .B2(n7535), .A(n7534), .ZN(n7536) );
  OAI211_X1 U9240 ( .C1(n7538), .C2(n8751), .A(n7537), .B(n7536), .ZN(P1_U3234) );
  INV_X1 U9241 ( .A(n7539), .ZN(n7545) );
  AOI21_X1 U9242 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n7541), .A(n7540), .ZN(
        n7542) );
  OAI21_X1 U9243 ( .B1(n7545), .B2(n8025), .A(n7542), .ZN(P2_U3335) );
  NOR2_X1 U9244 ( .A1(n7543), .A2(P1_U3084), .ZN(n9030) );
  AOI21_X1 U9245 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9488), .A(n9030), .ZN(
        n7544) );
  OAI21_X1 U9246 ( .B1(n7545), .B2(n9494), .A(n7544), .ZN(P1_U3330) );
  OAI21_X1 U9247 ( .B1(n8990), .B2(n7546), .A(n7686), .ZN(n7547) );
  NAND2_X1 U9248 ( .A1(n7547), .A2(n9706), .ZN(n7664) );
  INV_X1 U9249 ( .A(n8990), .ZN(n8883) );
  XNOR2_X1 U9250 ( .A(n7548), .B(n8883), .ZN(n7666) );
  NAND2_X1 U9251 ( .A1(n7666), .A2(n9300), .ZN(n7557) );
  AOI22_X1 U9252 ( .A1(n9241), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7659), .B2(
        n9701), .ZN(n7550) );
  NAND2_X1 U9253 ( .A1(n9335), .A2(n9432), .ZN(n7549) );
  OAI211_X1 U9254 ( .C1(n7551), .C2(n9338), .A(n7550), .B(n7549), .ZN(n7555)
         );
  OAI21_X1 U9255 ( .B1(n7552), .B2(n7671), .A(n9695), .ZN(n7553) );
  OR2_X1 U9256 ( .A1(n7553), .A2(n7692), .ZN(n7662) );
  NOR2_X1 U9257 ( .A1(n7662), .A2(n9344), .ZN(n7554) );
  AOI211_X1 U9258 ( .C1(n9347), .C2(n7645), .A(n7555), .B(n7554), .ZN(n7556)
         );
  OAI211_X1 U9259 ( .C1(n9241), .C2(n7664), .A(n7557), .B(n7556), .ZN(P1_U3278) );
  NAND2_X1 U9260 ( .A1(n9899), .A2(n9830), .ZN(n7558) );
  NAND2_X1 U9261 ( .A1(n7560), .A2(n7562), .ZN(n7561) );
  NAND2_X1 U9262 ( .A1(n7706), .A2(n7561), .ZN(n9906) );
  INV_X1 U9263 ( .A(n8521), .ZN(n7574) );
  XNOR2_X1 U9264 ( .A(n7563), .B(n7562), .ZN(n7565) );
  OAI22_X1 U9265 ( .A1(n9830), .A2(n8502), .B1(n9833), .B2(n8500), .ZN(n7564)
         );
  AOI21_X1 U9266 ( .B1(n7565), .B2(n9843), .A(n7564), .ZN(n7566) );
  OAI21_X1 U9267 ( .B1(n9906), .B2(n8508), .A(n7566), .ZN(n9909) );
  NAND2_X1 U9268 ( .A1(n9909), .A2(n8549), .ZN(n7573) );
  OAI22_X1 U9269 ( .A1(n8549), .A2(n7567), .B1(n9839), .B2(n8344), .ZN(n7571)
         );
  INV_X1 U9270 ( .A(n7704), .ZN(n9907) );
  NOR2_X1 U9271 ( .A1(n7568), .A2(n9907), .ZN(n7569) );
  OR2_X1 U9272 ( .A1(n9854), .A2(n7569), .ZN(n9908) );
  NOR2_X1 U9273 ( .A1(n9908), .A2(n8551), .ZN(n7570) );
  AOI211_X1 U9274 ( .C1(n9847), .C2(n7704), .A(n7571), .B(n7570), .ZN(n7572)
         );
  OAI211_X1 U9275 ( .C1(n9906), .C2(n7574), .A(n7573), .B(n7572), .ZN(P2_U3286) );
  INV_X1 U9276 ( .A(n7575), .ZN(n7578) );
  INV_X1 U9277 ( .A(n7576), .ZN(n7577) );
  NAND2_X1 U9278 ( .A1(n7578), .A2(n7577), .ZN(n7579) );
  NAND2_X1 U9279 ( .A1(n7580), .A2(n7579), .ZN(n7637) );
  NAND2_X1 U9280 ( .A1(n7618), .A2(n7989), .ZN(n7582) );
  NAND2_X1 U9281 ( .A1(n9041), .A2(n5005), .ZN(n7581) );
  NAND2_X1 U9282 ( .A1(n7582), .A2(n7581), .ZN(n7583) );
  XNOR2_X1 U9283 ( .A(n7583), .B(n4500), .ZN(n7638) );
  AND2_X1 U9284 ( .A1(n7983), .A2(n9041), .ZN(n7584) );
  AOI21_X1 U9285 ( .B1(n7618), .B2(n7901), .A(n7584), .ZN(n7635) );
  INV_X1 U9286 ( .A(n7635), .ZN(n7639) );
  XNOR2_X1 U9287 ( .A(n7638), .B(n7639), .ZN(n7585) );
  XNOR2_X1 U9288 ( .A(n7586), .B(n7585), .ZN(n7595) );
  NAND2_X1 U9289 ( .A1(n8749), .A2(n7587), .ZN(n7591) );
  INV_X1 U9290 ( .A(n7588), .ZN(n7589) );
  AOI21_X1 U9291 ( .B1(n8739), .B2(n9042), .A(n7589), .ZN(n7590) );
  OAI211_X1 U9292 ( .C1(n7592), .C2(n8737), .A(n7591), .B(n7590), .ZN(n7593)
         );
  AOI21_X1 U9293 ( .B1(n7618), .B2(n8767), .A(n7593), .ZN(n7594) );
  OAI21_X1 U9294 ( .B1(n7595), .B2(n7995), .A(n7594), .ZN(P1_U3222) );
  INV_X1 U9295 ( .A(n7596), .ZN(n7599) );
  OAI222_X1 U9296 ( .A1(n8130), .A2(n7598), .B1(n8025), .B2(n7599), .C1(n7597), 
        .C2(n8651), .ZN(P2_U3334) );
  OAI222_X1 U9297 ( .A1(n7600), .A2(P1_U3084), .B1(n9494), .B2(n7599), .C1(
        n10172), .C2(n9491), .ZN(P1_U3329) );
  NOR2_X1 U9298 ( .A1(n8224), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7601) );
  AOI21_X1 U9299 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8224), .A(n7601), .ZN(
        n8217) );
  OAI21_X1 U9300 ( .B1(n8224), .B2(P2_REG2_REG_14__SCAN_IN), .A(n8215), .ZN(
        n7725) );
  XNOR2_X1 U9301 ( .A(n7725), .B(n7605), .ZN(n7604) );
  INV_X1 U9302 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7603) );
  NAND2_X1 U9303 ( .A1(n7604), .A2(n7603), .ZN(n7727) );
  OAI21_X1 U9304 ( .B1(n7604), .B2(n7603), .A(n7727), .ZN(n7616) );
  INV_X1 U9305 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7608) );
  NAND2_X1 U9306 ( .A1(n8256), .A2(n7605), .ZN(n7607) );
  NAND2_X1 U9307 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n7606) );
  OAI211_X1 U9308 ( .C1(n8262), .C2(n7608), .A(n7607), .B(n7606), .ZN(n7615)
         );
  INV_X1 U9309 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9523) );
  AOI22_X1 U9310 ( .A1(n8224), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n9523), .B2(
        n7609), .ZN(n8222) );
  OAI21_X1 U9311 ( .B1(n7611), .B2(P2_REG1_REG_13__SCAN_IN), .A(n7610), .ZN(
        n8221) );
  NAND2_X1 U9312 ( .A1(n8222), .A2(n8221), .ZN(n8220) );
  OAI21_X1 U9313 ( .B1(n8224), .B2(P2_REG1_REG_14__SCAN_IN), .A(n8220), .ZN(
        n7718) );
  XNOR2_X1 U9314 ( .A(n7718), .B(n7726), .ZN(n7613) );
  INV_X1 U9315 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10209) );
  NOR2_X1 U9316 ( .A1(n10209), .A2(n7613), .ZN(n7719) );
  AOI211_X1 U9317 ( .C1(n7613), .C2(n10209), .A(n7719), .B(n7612), .ZN(n7614)
         );
  AOI211_X1 U9318 ( .C1(n8253), .C2(n7616), .A(n7615), .B(n7614), .ZN(n7617)
         );
  INV_X1 U9319 ( .A(n7617), .ZN(P2_U3260) );
  INV_X1 U9320 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7624) );
  AOI22_X1 U9321 ( .A1(n9794), .A2(n9042), .B1(n9040), .B2(n9791), .ZN(n7620)
         );
  NAND3_X1 U9322 ( .A1(n7621), .A2(n7620), .A3(n7619), .ZN(n7622) );
  AOI21_X1 U9323 ( .B1(n7623), .B2(n9789), .A(n7622), .ZN(n7626) );
  MUX2_X1 U9324 ( .A(n7624), .B(n7626), .S(n9809), .Z(n7625) );
  OAI21_X1 U9325 ( .B1(n4688), .B2(n9483), .A(n7625), .ZN(P1_U3490) );
  MUX2_X1 U9326 ( .A(n6636), .B(n7626), .S(n10189), .Z(n7627) );
  OAI21_X1 U9327 ( .B1(n4688), .B2(n9439), .A(n7627), .ZN(P1_U3535) );
  INV_X1 U9328 ( .A(n9848), .ZN(n9916) );
  OAI211_X1 U9329 ( .C1(n7630), .C2(n7629), .A(n7628), .B(n8138), .ZN(n7634)
         );
  OAI22_X1 U9330 ( .A1(n7757), .A2(n8500), .B1(n7703), .B2(n8502), .ZN(n9842)
         );
  NOR2_X1 U9331 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5309), .ZN(n8205) );
  INV_X1 U9332 ( .A(n9846), .ZN(n7631) );
  NOR2_X1 U9333 ( .A1(n9840), .A2(n7631), .ZN(n7632) );
  AOI211_X1 U9334 ( .C1(n7976), .C2(n9842), .A(n8205), .B(n7632), .ZN(n7633)
         );
  OAI211_X1 U9335 ( .C1(n9916), .C2(n9829), .A(n7634), .B(n7633), .ZN(P2_U3238) );
  NAND2_X1 U9336 ( .A1(n7638), .A2(n7635), .ZN(n7636) );
  INV_X1 U9337 ( .A(n7638), .ZN(n7640) );
  NAND2_X1 U9338 ( .A1(n7640), .A2(n7639), .ZN(n7641) );
  NAND2_X1 U9339 ( .A1(n7645), .A2(n7989), .ZN(n7643) );
  NAND2_X1 U9340 ( .A1(n9040), .A2(n7901), .ZN(n7642) );
  NAND2_X1 U9341 ( .A1(n7643), .A2(n7642), .ZN(n7644) );
  XNOR2_X1 U9342 ( .A(n7644), .B(n7986), .ZN(n7648) );
  NAND2_X1 U9343 ( .A1(n7645), .A2(n7901), .ZN(n7647) );
  NAND2_X1 U9344 ( .A1(n7983), .A2(n9040), .ZN(n7646) );
  NAND2_X1 U9345 ( .A1(n7647), .A2(n7646), .ZN(n7649) );
  AND2_X1 U9346 ( .A1(n7648), .A2(n7649), .ZN(n7653) );
  INV_X1 U9347 ( .A(n7648), .ZN(n7651) );
  INV_X1 U9348 ( .A(n7649), .ZN(n7650) );
  NAND2_X1 U9349 ( .A1(n7651), .A2(n7650), .ZN(n7812) );
  INV_X1 U9350 ( .A(n7812), .ZN(n7655) );
  OAI21_X1 U9351 ( .B1(n7655), .B2(n7653), .A(n7652), .ZN(n7654) );
  OAI21_X1 U9352 ( .B1(n7813), .B2(n7655), .A(n7654), .ZN(n7656) );
  NAND2_X1 U9353 ( .A1(n7656), .A2(n8744), .ZN(n7661) );
  AND2_X1 U9354 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9667) );
  AOI21_X1 U9355 ( .B1(n8739), .B2(n9041), .A(n9667), .ZN(n7657) );
  OAI21_X1 U9356 ( .B1(n8758), .B2(n8737), .A(n7657), .ZN(n7658) );
  AOI21_X1 U9357 ( .B1(n7659), .B2(n8749), .A(n7658), .ZN(n7660) );
  OAI211_X1 U9358 ( .C1(n7671), .C2(n8751), .A(n7661), .B(n7660), .ZN(P1_U3232) );
  INV_X1 U9359 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7667) );
  AOI22_X1 U9360 ( .A1(n9794), .A2(n9041), .B1(n9432), .B2(n9791), .ZN(n7663)
         );
  NAND3_X1 U9361 ( .A1(n7664), .A2(n7663), .A3(n7662), .ZN(n7665) );
  AOI21_X1 U9362 ( .B1(n7666), .B2(n9789), .A(n7665), .ZN(n7669) );
  MUX2_X1 U9363 ( .A(n7667), .B(n7669), .S(n9809), .Z(n7668) );
  OAI21_X1 U9364 ( .B1(n7671), .B2(n9483), .A(n7668), .ZN(P1_U3493) );
  MUX2_X1 U9365 ( .A(n7046), .B(n7669), .S(n10189), .Z(n7670) );
  OAI21_X1 U9366 ( .B1(n7671), .B2(n9439), .A(n7670), .ZN(P1_U3536) );
  NAND2_X1 U9367 ( .A1(n7672), .A2(n7736), .ZN(n7674) );
  XOR2_X1 U9368 ( .A(n7674), .B(n7673), .Z(n7680) );
  INV_X1 U9369 ( .A(n7712), .ZN(n7676) );
  OAI21_X1 U9370 ( .B1(n9840), .B2(n7676), .A(n7675), .ZN(n7678) );
  OAI22_X1 U9371 ( .A1(n9833), .A2(n9831), .B1(n9832), .B2(n8032), .ZN(n7677)
         );
  AOI211_X1 U9372 ( .C1(n8158), .C2(n9920), .A(n7678), .B(n7677), .ZN(n7679)
         );
  OAI21_X1 U9373 ( .B1(n7680), .B2(n9826), .A(n7679), .ZN(P2_U3226) );
  INV_X1 U9374 ( .A(n7681), .ZN(n7747) );
  OAI21_X1 U9375 ( .B1(n7685), .B2(n8964), .A(n7684), .ZN(n7784) );
  INV_X1 U9376 ( .A(n7784), .ZN(n7699) );
  NAND2_X1 U9377 ( .A1(n7686), .A2(n8890), .ZN(n7687) );
  NAND2_X1 U9378 ( .A1(n7687), .A2(n8964), .ZN(n7689) );
  NAND3_X1 U9379 ( .A1(n7689), .A2(n9706), .A3(n7688), .ZN(n7691) );
  AOI22_X1 U9380 ( .A1(n9794), .A2(n9040), .B1(n9540), .B2(n9791), .ZN(n7690)
         );
  NAND2_X1 U9381 ( .A1(n7691), .A2(n7690), .ZN(n7782) );
  INV_X1 U9382 ( .A(n7692), .ZN(n7694) );
  INV_X1 U9383 ( .A(n7776), .ZN(n7693) );
  AOI211_X1 U9384 ( .C1(n7824), .C2(n7694), .A(n9319), .B(n7693), .ZN(n7783)
         );
  NAND2_X1 U9385 ( .A1(n7783), .A2(n9321), .ZN(n7696) );
  AOI22_X1 U9386 ( .A1(n9241), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7820), .B2(
        n9701), .ZN(n7695) );
  OAI211_X1 U9387 ( .C1(n7789), .C2(n9326), .A(n7696), .B(n7695), .ZN(n7697)
         );
  AOI21_X1 U9388 ( .B1(n7782), .B2(n9716), .A(n7697), .ZN(n7698) );
  OAI21_X1 U9389 ( .B1(n7699), .B2(n9333), .A(n7698), .ZN(P1_U3277) );
  INV_X1 U9390 ( .A(n7700), .ZN(n7897) );
  OAI222_X1 U9391 ( .A1(P2_U3152), .A2(n7702), .B1(n8025), .B2(n7897), .C1(
        n7701), .C2(n8651), .ZN(P2_U3332) );
  INV_X1 U9392 ( .A(n7703), .ZN(n8168) );
  NAND2_X1 U9393 ( .A1(n7704), .A2(n8168), .ZN(n7705) );
  NAND2_X1 U9394 ( .A1(n7706), .A2(n7705), .ZN(n9850) );
  INV_X1 U9395 ( .A(n9833), .ZN(n8167) );
  NAND2_X1 U9396 ( .A1(n9848), .A2(n8167), .ZN(n7707) );
  INV_X1 U9397 ( .A(n7796), .ZN(n7709) );
  INV_X1 U9398 ( .A(n7790), .ZN(n7708) );
  OAI21_X1 U9399 ( .B1(n7709), .B2(n7708), .A(n7750), .ZN(n9926) );
  INV_X1 U9400 ( .A(n9926), .ZN(n7717) );
  XOR2_X1 U9401 ( .A(n7790), .B(n7710), .Z(n7711) );
  OAI222_X1 U9402 ( .A1(n8500), .A2(n8032), .B1(n8502), .B2(n9833), .C1(n7711), 
        .C2(n8488), .ZN(n9924) );
  XNOR2_X1 U9403 ( .A(n4481), .B(n9920), .ZN(n9923) );
  AOI22_X1 U9404 ( .A1(n9860), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7712), .B2(
        n9845), .ZN(n7714) );
  NAND2_X1 U9405 ( .A1(n9847), .A2(n9920), .ZN(n7713) );
  OAI211_X1 U9406 ( .C1(n9923), .C2(n8551), .A(n7714), .B(n7713), .ZN(n7715)
         );
  AOI21_X1 U9407 ( .B1(n9924), .B2(n8549), .A(n7715), .ZN(n7716) );
  OAI21_X1 U9408 ( .B1(n7717), .B2(n8543), .A(n7716), .ZN(P2_U3284) );
  NOR2_X1 U9409 ( .A1(n7726), .A2(n7718), .ZN(n7720) );
  NOR2_X1 U9410 ( .A1(n7720), .A2(n7719), .ZN(n7722) );
  XOR2_X1 U9411 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n7835), .Z(n7721) );
  NAND2_X1 U9412 ( .A1(n7721), .A2(n7722), .ZN(n7827) );
  OAI21_X1 U9413 ( .B1(n7722), .B2(n7721), .A(n7827), .ZN(n7734) );
  INV_X1 U9414 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7724) );
  NAND2_X1 U9415 ( .A1(n8256), .A2(n7835), .ZN(n7723) );
  NAND2_X1 U9416 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8095) );
  OAI211_X1 U9417 ( .C1(n8262), .C2(n7724), .A(n7723), .B(n8095), .ZN(n7733)
         );
  NAND2_X1 U9418 ( .A1(n7726), .A2(n7725), .ZN(n7728) );
  NAND2_X1 U9419 ( .A1(n7728), .A2(n7727), .ZN(n7731) );
  NAND2_X1 U9420 ( .A1(n7835), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7729) );
  OAI21_X1 U9421 ( .B1(n7835), .B2(P2_REG2_REG_16__SCAN_IN), .A(n7729), .ZN(
        n7730) );
  NOR2_X1 U9422 ( .A1(n7730), .A2(n7731), .ZN(n7834) );
  AOI211_X1 U9423 ( .C1(n7731), .C2(n7730), .A(n7834), .B(n8254), .ZN(n7732)
         );
  AOI211_X1 U9424 ( .C1(n7734), .C2(n8258), .A(n7733), .B(n7732), .ZN(n7735)
         );
  INV_X1 U9425 ( .A(n7735), .ZN(P2_U3261) );
  NAND2_X1 U9426 ( .A1(n7737), .A2(n7736), .ZN(n8027) );
  XNOR2_X1 U9427 ( .A(n8027), .B(n8026), .ZN(n7742) );
  OAI22_X1 U9428 ( .A1(n7757), .A2(n9831), .B1(n9832), .B2(n8155), .ZN(n7738)
         );
  AOI211_X1 U9429 ( .C1(n8144), .C2(n7764), .A(n7739), .B(n7738), .ZN(n7741)
         );
  NAND2_X1 U9430 ( .A1(n8158), .A2(n9525), .ZN(n7740) );
  OAI211_X1 U9431 ( .C1(n7742), .C2(n9826), .A(n7741), .B(n7740), .ZN(P2_U3236) );
  INV_X1 U9432 ( .A(n7743), .ZN(n8648) );
  AOI21_X1 U9433 ( .B1(n9488), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7744), .ZN(
        n7745) );
  OAI21_X1 U9434 ( .B1(n8648), .B2(n9494), .A(n7745), .ZN(P1_U3326) );
  OAI222_X1 U9435 ( .A1(P1_U3084), .A2(n7748), .B1(n9494), .B2(n7747), .C1(
        n7746), .C2(n9491), .ZN(P1_U3328) );
  INV_X1 U9436 ( .A(n7757), .ZN(n8166) );
  OR2_X1 U9437 ( .A1(n9920), .A2(n8166), .ZN(n7749) );
  AND2_X1 U9438 ( .A1(n7755), .A2(n7749), .ZN(n7791) );
  NAND2_X1 U9439 ( .A1(n7750), .A2(n7791), .ZN(n7754) );
  NAND2_X1 U9440 ( .A1(n7750), .A2(n7749), .ZN(n7752) );
  NAND2_X1 U9441 ( .A1(n7752), .A2(n7751), .ZN(n7753) );
  NAND2_X1 U9442 ( .A1(n7754), .A2(n7753), .ZN(n7761) );
  XNOR2_X1 U9443 ( .A(n7756), .B(n7755), .ZN(n7759) );
  OAI22_X1 U9444 ( .A1(n7757), .A2(n8502), .B1(n8155), .B2(n8500), .ZN(n7758)
         );
  AOI21_X1 U9445 ( .B1(n7759), .B2(n9843), .A(n7758), .ZN(n7760) );
  OAI21_X1 U9446 ( .B1(n7761), .B2(n8508), .A(n7760), .ZN(n9528) );
  INV_X1 U9447 ( .A(n9528), .ZN(n7769) );
  INV_X1 U9448 ( .A(n7761), .ZN(n9530) );
  AND2_X1 U9449 ( .A1(n7762), .A2(n9525), .ZN(n7763) );
  OR2_X1 U9450 ( .A1(n7763), .A2(n7805), .ZN(n9527) );
  AOI22_X1 U9451 ( .A1(n9860), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7764), .B2(
        n9845), .ZN(n7766) );
  NAND2_X1 U9452 ( .A1(n9847), .A2(n9525), .ZN(n7765) );
  OAI211_X1 U9453 ( .C1(n9527), .C2(n8551), .A(n7766), .B(n7765), .ZN(n7767)
         );
  AOI21_X1 U9454 ( .B1(n9530), .B2(n8521), .A(n7767), .ZN(n7768) );
  OAI21_X1 U9455 ( .B1(n7769), .B2(n9860), .A(n7768), .ZN(P2_U3283) );
  OAI211_X1 U9456 ( .C1(n7771), .C2(n8991), .A(n7770), .B(n9706), .ZN(n9435)
         );
  XOR2_X1 U9457 ( .A(n7772), .B(n8991), .Z(n9437) );
  NAND2_X1 U9458 ( .A1(n9437), .A2(n9300), .ZN(n7781) );
  AOI22_X1 U9459 ( .A1(n9241), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n7773), .B2(
        n9701), .ZN(n7775) );
  NAND2_X1 U9460 ( .A1(n9335), .A2(n9431), .ZN(n7774) );
  OAI211_X1 U9461 ( .C1(n8758), .C2(n9338), .A(n7775), .B(n7774), .ZN(n7779)
         );
  AOI21_X1 U9462 ( .B1(n7776), .B2(n8768), .A(n9319), .ZN(n7777) );
  NAND2_X1 U9463 ( .A1(n7777), .A2(n9340), .ZN(n9433) );
  NOR2_X1 U9464 ( .A1(n9433), .A2(n9344), .ZN(n7778) );
  AOI211_X1 U9465 ( .C1(n9347), .C2(n8768), .A(n7779), .B(n7778), .ZN(n7780)
         );
  OAI211_X1 U9466 ( .C1(n9208), .C2(n9435), .A(n7781), .B(n7780), .ZN(P1_U3276) );
  INV_X1 U9467 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n7785) );
  AOI211_X1 U9468 ( .C1(n7784), .C2(n9789), .A(n7783), .B(n7782), .ZN(n7787)
         );
  MUX2_X1 U9469 ( .A(n7785), .B(n7787), .S(n9809), .Z(n7786) );
  OAI21_X1 U9470 ( .B1(n7789), .B2(n9483), .A(n7786), .ZN(P1_U3496) );
  MUX2_X1 U9471 ( .A(n7051), .B(n7787), .S(n10189), .Z(n7788) );
  OAI21_X1 U9472 ( .B1(n7789), .B2(n9439), .A(n7788), .ZN(P1_U3537) );
  AND2_X1 U9473 ( .A1(n9525), .A2(n8165), .ZN(n7792) );
  OR2_X1 U9474 ( .A1(n7790), .A2(n7792), .ZN(n7794) );
  OR2_X1 U9475 ( .A1(n7796), .A2(n7794), .ZN(n7793) );
  OR2_X1 U9476 ( .A1(n7792), .A2(n7791), .ZN(n7797) );
  OR2_X1 U9477 ( .A1(n7794), .A2(n7801), .ZN(n7795) );
  OR2_X1 U9478 ( .A1(n7801), .A2(n7797), .ZN(n8268) );
  AND2_X1 U9479 ( .A1(n8271), .A2(n8268), .ZN(n7798) );
  OAI21_X1 U9480 ( .B1(n4473), .B2(n7799), .A(n7798), .ZN(n9522) );
  INV_X1 U9481 ( .A(n9522), .ZN(n7810) );
  OAI211_X1 U9482 ( .C1(n4474), .C2(n7801), .A(n7800), .B(n9843), .ZN(n7803)
         );
  INV_X1 U9483 ( .A(n8503), .ZN(n8272) );
  AOI22_X1 U9484 ( .A1(n8533), .A2(n8272), .B1(n8165), .B2(n8530), .ZN(n7802)
         );
  NAND2_X1 U9485 ( .A1(n7803), .A2(n7802), .ZN(n9520) );
  INV_X1 U9486 ( .A(n8267), .ZN(n9518) );
  INV_X1 U9487 ( .A(n8536), .ZN(n7804) );
  OAI21_X1 U9488 ( .B1(n9518), .B2(n7805), .A(n7804), .ZN(n9519) );
  AOI22_X1 U9489 ( .A1(n9860), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8034), .B2(
        n9845), .ZN(n7807) );
  NAND2_X1 U9490 ( .A1(n9847), .A2(n8267), .ZN(n7806) );
  OAI211_X1 U9491 ( .C1(n9519), .C2(n8551), .A(n7807), .B(n7806), .ZN(n7808)
         );
  AOI21_X1 U9492 ( .B1(n9520), .B2(n8549), .A(n7808), .ZN(n7809) );
  OAI21_X1 U9493 ( .B1(n7810), .B2(n8543), .A(n7809), .ZN(P2_U3282) );
  AOI22_X1 U9494 ( .A1(n7824), .A2(n7811), .B1(n7983), .B2(n9432), .ZN(n7899)
         );
  NAND2_X1 U9495 ( .A1(n7824), .A2(n7989), .ZN(n7815) );
  NAND2_X1 U9496 ( .A1(n9432), .A2(n7988), .ZN(n7814) );
  NAND2_X1 U9497 ( .A1(n7815), .A2(n7814), .ZN(n7816) );
  XNOR2_X1 U9498 ( .A(n7816), .B(n7986), .ZN(n7818) );
  NOR2_X1 U9499 ( .A1(n7900), .A2(n7906), .ZN(n7819) );
  XOR2_X1 U9500 ( .A(n7899), .B(n7819), .Z(n7826) );
  NAND2_X1 U9501 ( .A1(n8749), .A2(n7820), .ZN(n7822) );
  NOR2_X1 U9502 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10232), .ZN(n9676) );
  AOI21_X1 U9503 ( .B1(n8739), .B2(n9040), .A(n9676), .ZN(n7821) );
  OAI211_X1 U9504 ( .C1(n9339), .C2(n8737), .A(n7822), .B(n7821), .ZN(n7823)
         );
  AOI21_X1 U9505 ( .B1(n7824), .B2(n8767), .A(n7823), .ZN(n7825) );
  OAI21_X1 U9506 ( .B1(n7826), .B2(n7995), .A(n7825), .ZN(P1_U3213) );
  INV_X1 U9507 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7833) );
  OAI21_X1 U9508 ( .B1(n7835), .B2(P2_REG1_REG_16__SCAN_IN), .A(n7827), .ZN(
        n7829) );
  XNOR2_X1 U9509 ( .A(n8238), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n7828) );
  NOR2_X1 U9510 ( .A1(n7828), .A2(n7829), .ZN(n8237) );
  AOI21_X1 U9511 ( .B1(n7829), .B2(n7828), .A(n8237), .ZN(n7830) );
  NAND2_X1 U9512 ( .A1(n8258), .A2(n7830), .ZN(n7832) );
  NAND2_X1 U9513 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(n8130), .ZN(n7831) );
  OAI211_X1 U9514 ( .C1(n8262), .C2(n7833), .A(n7832), .B(n7831), .ZN(n7840)
         );
  AOI21_X1 U9515 ( .B1(n7835), .B2(P2_REG2_REG_16__SCAN_IN), .A(n7834), .ZN(
        n7838) );
  NAND2_X1 U9516 ( .A1(n8238), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7836) );
  OAI21_X1 U9517 ( .B1(n8238), .B2(P2_REG2_REG_17__SCAN_IN), .A(n7836), .ZN(
        n7837) );
  NOR2_X1 U9518 ( .A1(n7838), .A2(n7837), .ZN(n8229) );
  AOI211_X1 U9519 ( .C1(n7838), .C2(n7837), .A(n8229), .B(n8254), .ZN(n7839)
         );
  AOI211_X1 U9520 ( .C1(n8256), .C2(n8238), .A(n7840), .B(n7839), .ZN(n7841)
         );
  INV_X1 U9521 ( .A(n7841), .ZN(P2_U3262) );
  INV_X1 U9522 ( .A(n8781), .ZN(n9493) );
  OAI222_X1 U9523 ( .A1(n8025), .A2(n9493), .B1(P2_U3152), .B2(n7842), .C1(
        n10016), .C2(n8651), .ZN(P2_U3329) );
  NOR4_X1 U9524 ( .A1(n7843), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n6121), .ZN(n7844) );
  AOI21_X1 U9525 ( .B1(n9488), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n7844), .ZN(
        n7845) );
  OAI21_X1 U9526 ( .B1(n8771), .B2(n9494), .A(n7845), .ZN(P1_U3322) );
  NAND3_X1 U9527 ( .A1(n7846), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n7848) );
  OAI22_X1 U9528 ( .A1(n5023), .A2(n7848), .B1(n7847), .B2(n8651), .ZN(n7849)
         );
  INV_X1 U9529 ( .A(n7849), .ZN(n7850) );
  OAI21_X1 U9530 ( .B1(n8771), .B2(n8025), .A(n7850), .ZN(P2_U3327) );
  INV_X1 U9531 ( .A(n8538), .ZN(n9513) );
  INV_X1 U9532 ( .A(n8611), .ZN(n8457) );
  NAND2_X1 U9533 ( .A1(n8468), .A2(n8457), .ZN(n8452) );
  INV_X1 U9534 ( .A(n8576), .ZN(n8147) );
  INV_X1 U9535 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n10214) );
  INV_X1 U9536 ( .A(P2_B_REG_SCAN_IN), .ZN(n7853) );
  OAI21_X1 U9537 ( .B1(n8649), .B2(n7853), .A(n8533), .ZN(n8287) );
  NOR2_X1 U9538 ( .A1(n7854), .A2(n8287), .ZN(n9510) );
  NAND2_X1 U9539 ( .A1(n8549), .A2(n9510), .ZN(n8263) );
  OAI21_X1 U9540 ( .B1(n10214), .B2(n8549), .A(n8263), .ZN(n7855) );
  AOI21_X1 U9541 ( .B1(n8556), .B2(n9847), .A(n7855), .ZN(n7856) );
  OAI21_X1 U9542 ( .B1(n8558), .B2(n8551), .A(n7856), .ZN(P2_U3265) );
  INV_X1 U9543 ( .A(n7857), .ZN(n7858) );
  AOI21_X1 U9544 ( .B1(n7860), .B2(n7859), .A(n7858), .ZN(n7865) );
  AOI22_X1 U9545 ( .A1(n8739), .A2(n6576), .B1(n8762), .B2(n9748), .ZN(n7864)
         );
  AOI22_X1 U9546 ( .A1(n8767), .A2(n7862), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n7861), .ZN(n7863) );
  OAI211_X1 U9547 ( .C1(n7865), .C2(n7995), .A(n7864), .B(n7863), .ZN(P1_U3235) );
  XOR2_X1 U9548 ( .A(n7867), .B(n7866), .Z(n7870) );
  AOI21_X1 U9549 ( .B1(n8138), .B2(n7870), .A(n7869), .ZN(n7872) );
  AOI22_X1 U9550 ( .A1(n8144), .A2(n5097), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8130), .ZN(n7871) );
  OAI211_X1 U9551 ( .C1(n5717), .C2(n9831), .A(n7872), .B(n7871), .ZN(P2_U3220) );
  NAND2_X1 U9552 ( .A1(n7873), .A2(n9321), .ZN(n7879) );
  INV_X1 U9553 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n7874) );
  OAI22_X1 U9554 ( .A1(n9716), .A2(n7874), .B1(n8001), .B2(n9301), .ZN(n7877)
         );
  NOR2_X1 U9555 ( .A1(n9338), .A2(n7875), .ZN(n7876) );
  AOI211_X1 U9556 ( .C1(n9335), .C2(n9038), .A(n7877), .B(n7876), .ZN(n7878)
         );
  OAI211_X1 U9557 ( .C1(n4706), .C2(n9326), .A(n7879), .B(n7878), .ZN(n7880)
         );
  AOI21_X1 U9558 ( .B1(n7882), .B2(n7881), .A(n7880), .ZN(n7883) );
  OAI21_X1 U9559 ( .B1(n7884), .B2(n9333), .A(n7883), .ZN(P1_U3263) );
  INV_X1 U9560 ( .A(n7885), .ZN(n8647) );
  OAI222_X1 U9561 ( .A1(n6372), .A2(P1_U3084), .B1(n9494), .B2(n8647), .C1(
        n7886), .C2(n9491), .ZN(P1_U3325) );
  INV_X1 U9562 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7887) );
  OAI22_X1 U9563 ( .A1(n9855), .A2(n7888), .B1(n7887), .B2(n8344), .ZN(n7889)
         );
  AOI21_X1 U9564 ( .B1(n9847), .B2(n7890), .A(n7889), .ZN(n7894) );
  MUX2_X1 U9565 ( .A(n7892), .B(n7891), .S(n8549), .Z(n7893) );
  OAI211_X1 U9566 ( .C1(n7895), .C2(n8543), .A(n7894), .B(n7893), .ZN(P2_U3295) );
  OAI222_X1 U9567 ( .A1(n6409), .A2(P1_U3084), .B1(n9494), .B2(n7897), .C1(
        n7896), .C2(n9491), .ZN(P1_U3327) );
  AOI22_X1 U9568 ( .A1(n9539), .A2(n7988), .B1(n7983), .B2(n9431), .ZN(n7908)
         );
  AOI22_X1 U9569 ( .A1(n9539), .A2(n7989), .B1(n7901), .B2(n9431), .ZN(n7898)
         );
  XNOR2_X1 U9570 ( .A(n7898), .B(n7986), .ZN(n7907) );
  NAND2_X1 U9571 ( .A1(n8768), .A2(n7989), .ZN(n7903) );
  NAND2_X1 U9572 ( .A1(n9540), .A2(n7901), .ZN(n7902) );
  NAND2_X1 U9573 ( .A1(n7903), .A2(n7902), .ZN(n7904) );
  XNOR2_X1 U9574 ( .A(n7904), .B(n7986), .ZN(n7905) );
  AOI22_X1 U9575 ( .A1(n8768), .A2(n7988), .B1(n7983), .B2(n9540), .ZN(n8755)
         );
  XNOR2_X1 U9576 ( .A(n7907), .B(n7908), .ZN(n8690) );
  AOI22_X1 U9577 ( .A1(n9428), .A2(n7988), .B1(n7983), .B2(n9541), .ZN(n7912)
         );
  NAND2_X1 U9578 ( .A1(n9428), .A2(n7989), .ZN(n7910) );
  NAND2_X1 U9579 ( .A1(n9541), .A2(n7988), .ZN(n7909) );
  NAND2_X1 U9580 ( .A1(n7910), .A2(n7909), .ZN(n7911) );
  XNOR2_X1 U9581 ( .A(n7911), .B(n7986), .ZN(n7914) );
  XOR2_X1 U9582 ( .A(n7912), .B(n7914), .Z(n8697) );
  INV_X1 U9583 ( .A(n7912), .ZN(n7913) );
  AOI22_X1 U9584 ( .A1(n9421), .A2(n7989), .B1(n7988), .B2(n9411), .ZN(n7915)
         );
  AOI22_X1 U9585 ( .A1(n9421), .A2(n7988), .B1(n7983), .B2(n9411), .ZN(n8733)
         );
  NAND2_X1 U9586 ( .A1(n9289), .A2(n7989), .ZN(n7917) );
  NAND2_X1 U9587 ( .A1(n9295), .A2(n7988), .ZN(n7916) );
  NAND2_X1 U9588 ( .A1(n7917), .A2(n7916), .ZN(n7918) );
  XNOR2_X1 U9589 ( .A(n7918), .B(n7986), .ZN(n8665) );
  NAND2_X1 U9590 ( .A1(n9289), .A2(n7988), .ZN(n7920) );
  NAND2_X1 U9591 ( .A1(n9295), .A2(n7983), .ZN(n7919) );
  NAND2_X1 U9592 ( .A1(n7920), .A2(n7919), .ZN(n7922) );
  INV_X1 U9593 ( .A(n7922), .ZN(n8664) );
  NAND2_X1 U9594 ( .A1(n9265), .A2(n7989), .ZN(n7926) );
  NAND2_X1 U9595 ( .A1(n9412), .A2(n7988), .ZN(n7925) );
  NAND2_X1 U9596 ( .A1(n7926), .A2(n7925), .ZN(n7927) );
  XNOR2_X1 U9597 ( .A(n7927), .B(n4500), .ZN(n7930) );
  AND2_X1 U9598 ( .A1(n9412), .A2(n7983), .ZN(n7928) );
  AOI21_X1 U9599 ( .B1(n9265), .B2(n7988), .A(n7928), .ZN(n7929) );
  NAND2_X1 U9600 ( .A1(n7930), .A2(n7929), .ZN(n8715) );
  NOR2_X1 U9601 ( .A1(n7930), .A2(n7929), .ZN(n8716) );
  AOI22_X1 U9602 ( .A1(n9249), .A2(n7989), .B1(n7988), .B2(n9260), .ZN(n7931)
         );
  XOR2_X1 U9603 ( .A(n7986), .B(n7931), .Z(n7934) );
  OAI22_X1 U9604 ( .A1(n9471), .A2(n7935), .B1(n7932), .B2(n7941), .ZN(n7933)
         );
  NAND2_X1 U9605 ( .A1(n7934), .A2(n7933), .ZN(n8672) );
  OAI22_X1 U9606 ( .A1(n9467), .A2(n7935), .B1(n9247), .B2(n7941), .ZN(n7937)
         );
  AOI22_X1 U9607 ( .A1(n4695), .A2(n7989), .B1(n7988), .B2(n9389), .ZN(n7936)
         );
  XNOR2_X1 U9608 ( .A(n7936), .B(n7986), .ZN(n8725) );
  NAND2_X1 U9609 ( .A1(n8723), .A2(n8725), .ZN(n7939) );
  INV_X1 U9610 ( .A(n7937), .ZN(n7938) );
  AOI22_X1 U9611 ( .A1(n9220), .A2(n7989), .B1(n7988), .B2(n9228), .ZN(n7940)
         );
  XOR2_X1 U9612 ( .A(n7986), .B(n7940), .Z(n7942) );
  INV_X1 U9613 ( .A(n7942), .ZN(n8655) );
  OAI22_X1 U9614 ( .A1(n9464), .A2(n7935), .B1(n9196), .B2(n7941), .ZN(n8654)
         );
  AOI22_X1 U9615 ( .A1(n9199), .A2(n7989), .B1(n7988), .B2(n9388), .ZN(n7944)
         );
  XNOR2_X1 U9616 ( .A(n7944), .B(n7986), .ZN(n7946) );
  AOI22_X1 U9617 ( .A1(n9199), .A2(n7988), .B1(n7983), .B2(n9388), .ZN(n7945)
         );
  NAND2_X1 U9618 ( .A1(n7946), .A2(n7945), .ZN(n7947) );
  OAI21_X1 U9619 ( .B1(n7946), .B2(n7945), .A(n7947), .ZN(n8708) );
  NAND2_X1 U9620 ( .A1(n9185), .A2(n7989), .ZN(n7949) );
  NAND2_X1 U9621 ( .A1(n9161), .A2(n7988), .ZN(n7948) );
  NAND2_X1 U9622 ( .A1(n7949), .A2(n7948), .ZN(n7950) );
  XNOR2_X1 U9623 ( .A(n7950), .B(n7986), .ZN(n7954) );
  NAND2_X1 U9624 ( .A1(n9185), .A2(n7988), .ZN(n7952) );
  NAND2_X1 U9625 ( .A1(n7983), .A2(n9161), .ZN(n7951) );
  NAND2_X1 U9626 ( .A1(n7952), .A2(n7951), .ZN(n7953) );
  NAND2_X1 U9627 ( .A1(n7954), .A2(n7953), .ZN(n8680) );
  AND2_X1 U9628 ( .A1(n7983), .A2(n9180), .ZN(n7955) );
  AOI21_X1 U9629 ( .B1(n9166), .B2(n7988), .A(n7955), .ZN(n7958) );
  AOI22_X1 U9630 ( .A1(n9166), .A2(n7989), .B1(n7988), .B2(n9180), .ZN(n7956)
         );
  XNOR2_X1 U9631 ( .A(n7956), .B(n7986), .ZN(n7957) );
  XOR2_X1 U9632 ( .A(n7958), .B(n7957), .Z(n8746) );
  INV_X1 U9633 ( .A(n7957), .ZN(n7960) );
  AND2_X1 U9634 ( .A1(n7983), .A2(n9160), .ZN(n7961) );
  AOI21_X1 U9635 ( .B1(n9370), .B2(n7988), .A(n7961), .ZN(n7982) );
  NAND2_X1 U9636 ( .A1(n9370), .A2(n7989), .ZN(n7963) );
  NAND2_X1 U9637 ( .A1(n9160), .A2(n7988), .ZN(n7962) );
  NAND2_X1 U9638 ( .A1(n7963), .A2(n7962), .ZN(n7964) );
  XNOR2_X1 U9639 ( .A(n7964), .B(n7986), .ZN(n7994) );
  INV_X1 U9640 ( .A(n9144), .ZN(n7968) );
  OAI22_X1 U9641 ( .A1(n8759), .A2(n9148), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9977), .ZN(n7966) );
  AOI21_X1 U9642 ( .B1(n8762), .B2(n9039), .A(n7966), .ZN(n7967) );
  OAI21_X1 U9643 ( .B1(n8765), .B2(n7968), .A(n7967), .ZN(n7969) );
  AOI21_X1 U9644 ( .B1(n9370), .B2(n8767), .A(n7969), .ZN(n7970) );
  OAI21_X1 U9645 ( .B1(n7973), .B2(n7972), .A(n7971), .ZN(n7974) );
  AOI22_X1 U9646 ( .A1(n7976), .A2(n7975), .B1(n8138), .B2(n7974), .ZN(n7980)
         );
  OR2_X1 U9647 ( .A1(n7978), .A2(n7977), .ZN(n8019) );
  NAND2_X1 U9648 ( .A1(n8019), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n7979) );
  OAI211_X1 U9649 ( .C1(n7981), .C2(n9829), .A(n7980), .B(n7979), .ZN(P2_U3224) );
  INV_X1 U9650 ( .A(n7982), .ZN(n7993) );
  NAND2_X1 U9651 ( .A1(n8006), .A2(n7988), .ZN(n7985) );
  NAND2_X1 U9652 ( .A1(n7983), .A2(n9039), .ZN(n7984) );
  NAND2_X1 U9653 ( .A1(n7985), .A2(n7984), .ZN(n7987) );
  XNOR2_X1 U9654 ( .A(n7987), .B(n7986), .ZN(n7991) );
  AOI22_X1 U9655 ( .A1(n8006), .A2(n7989), .B1(n7988), .B2(n9039), .ZN(n7990)
         );
  XNOR2_X1 U9656 ( .A(n7991), .B(n7990), .ZN(n8003) );
  INV_X1 U9657 ( .A(n8003), .ZN(n7992) );
  NAND2_X1 U9658 ( .A1(n7992), .A2(n8744), .ZN(n8009) );
  NAND2_X1 U9659 ( .A1(n7994), .A2(n7993), .ZN(n8002) );
  INV_X1 U9660 ( .A(n8002), .ZN(n7996) );
  AND2_X1 U9661 ( .A1(n8003), .A2(n7997), .ZN(n7998) );
  AOI22_X1 U9662 ( .A1(n8739), .A2(n9160), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8000) );
  NAND2_X1 U9663 ( .A1(n8762), .A2(n9038), .ZN(n7999) );
  OAI211_X1 U9664 ( .C1(n8765), .C2(n8001), .A(n8000), .B(n7999), .ZN(n8005)
         );
  NOR3_X1 U9665 ( .A1(n8003), .A2(n7995), .A3(n8002), .ZN(n8004) );
  AOI211_X1 U9666 ( .C1(n8006), .C2(n8767), .A(n8005), .B(n8004), .ZN(n8007)
         );
  OAI211_X1 U9667 ( .C1(n8010), .C2(n8009), .A(n8008), .B(n8007), .ZN(P1_U3218) );
  INV_X1 U9668 ( .A(n9832), .ZN(n8011) );
  AOI22_X1 U9669 ( .A1(n8011), .A2(n8175), .B1(n8158), .B2(n8545), .ZN(n8016)
         );
  XOR2_X1 U9670 ( .A(n8012), .B(n8013), .Z(n8014) );
  AOI22_X1 U9671 ( .A1(n8138), .A2(n8014), .B1(n8019), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n8015) );
  OAI211_X1 U9672 ( .C1(n8024), .C2(n9831), .A(n8016), .B(n8015), .ZN(P2_U3239) );
  NOR3_X1 U9673 ( .A1(n9826), .A2(n9853), .A3(n8017), .ZN(n8018) );
  AOI21_X1 U9674 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n8019), .A(n8018), .ZN(
        n8023) );
  AOI21_X1 U9675 ( .B1(n9922), .B2(n5716), .A(n9826), .ZN(n8021) );
  OAI21_X1 U9676 ( .B1(n8021), .B2(n8158), .A(n8020), .ZN(n8022) );
  OAI211_X1 U9677 ( .C1(n8024), .C2(n9832), .A(n8023), .B(n8022), .ZN(P2_U3234) );
  INV_X1 U9678 ( .A(n8776), .ZN(n9490) );
  NAND2_X1 U9679 ( .A1(n8027), .A2(n8026), .ZN(n8029) );
  NAND2_X1 U9680 ( .A1(n8029), .A2(n8028), .ZN(n8030) );
  AOI21_X1 U9681 ( .B1(n8031), .B2(n8030), .A(n4472), .ZN(n8037) );
  AND2_X1 U9682 ( .A1(n8130), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8219) );
  OAI22_X1 U9683 ( .A1(n8503), .A2(n9832), .B1(n9831), .B2(n8032), .ZN(n8033)
         );
  AOI211_X1 U9684 ( .C1(n8144), .C2(n8034), .A(n8219), .B(n8033), .ZN(n8036)
         );
  NAND2_X1 U9685 ( .A1(n8158), .A2(n8267), .ZN(n8035) );
  OAI211_X1 U9686 ( .C1(n8037), .C2(n9826), .A(n8036), .B(n8035), .ZN(P2_U3217) );
  XNOR2_X1 U9687 ( .A(n8039), .B(n8038), .ZN(n8040) );
  XNOR2_X1 U9688 ( .A(n8041), .B(n8040), .ZN(n8046) );
  OAI22_X1 U9689 ( .A1(n9840), .A2(n8386), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8042), .ZN(n8044) );
  OAI22_X1 U9690 ( .A1(n8356), .A2(n9832), .B1(n9831), .B2(n8429), .ZN(n8043)
         );
  AOI211_X1 U9691 ( .C1(n8589), .C2(n8158), .A(n8044), .B(n8043), .ZN(n8045)
         );
  OAI21_X1 U9692 ( .B1(n8046), .B2(n9826), .A(n8045), .ZN(P2_U3218) );
  INV_X1 U9693 ( .A(n4494), .ZN(n8048) );
  AOI21_X1 U9694 ( .B1(n8050), .B2(n8049), .A(n8048), .ZN(n8054) );
  AND2_X1 U9695 ( .A1(n8130), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8260) );
  OAI22_X1 U9696 ( .A1(n8274), .A2(n9831), .B1(n9832), .B2(n8428), .ZN(n8051)
         );
  AOI211_X1 U9697 ( .C1(n8144), .C2(n8455), .A(n8260), .B(n8051), .ZN(n8053)
         );
  NAND2_X1 U9698 ( .A1(n8611), .A2(n8158), .ZN(n8052) );
  OAI211_X1 U9699 ( .C1(n8054), .C2(n9826), .A(n8053), .B(n8052), .ZN(P2_U3221) );
  INV_X1 U9700 ( .A(n8066), .ZN(n8059) );
  OR2_X1 U9701 ( .A1(n8286), .A2(n9853), .ZN(n8056) );
  XNOR2_X1 U9702 ( .A(n8056), .B(n8055), .ZN(n8057) );
  XNOR2_X1 U9703 ( .A(n8564), .B(n8057), .ZN(n8068) );
  NAND2_X1 U9704 ( .A1(n8059), .A2(n8058), .ZN(n8073) );
  INV_X1 U9705 ( .A(n8305), .ZN(n8061) );
  OAI22_X1 U9706 ( .A1(n9840), .A2(n8061), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8060), .ZN(n8064) );
  OAI22_X1 U9707 ( .A1(n8163), .A2(n9832), .B1(n9831), .B2(n8062), .ZN(n8063)
         );
  AOI211_X1 U9708 ( .C1(n8564), .C2(n8158), .A(n8064), .B(n8063), .ZN(n8072)
         );
  INV_X1 U9709 ( .A(n8068), .ZN(n8065) );
  INV_X1 U9710 ( .A(n8067), .ZN(n8069) );
  NAND3_X1 U9711 ( .A1(n8069), .A2(n8138), .A3(n8068), .ZN(n8070) );
  NAND4_X1 U9712 ( .A1(n8073), .A2(n8072), .A3(n8071), .A4(n8070), .ZN(
        P2_U3222) );
  XNOR2_X1 U9713 ( .A(n8075), .B(n8074), .ZN(n8081) );
  INV_X1 U9714 ( .A(n8430), .ZN(n8077) );
  OAI22_X1 U9715 ( .A1(n9840), .A2(n8077), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8076), .ZN(n8079) );
  OAI22_X1 U9716 ( .A1(n8428), .A2(n9831), .B1(n9832), .B2(n8429), .ZN(n8078)
         );
  AOI211_X1 U9717 ( .C1(n8601), .C2(n8158), .A(n8079), .B(n8078), .ZN(n8080)
         );
  OAI21_X1 U9718 ( .B1(n8081), .B2(n9826), .A(n8080), .ZN(P2_U3225) );
  XNOR2_X1 U9719 ( .A(n8083), .B(n8082), .ZN(n8084) );
  XNOR2_X1 U9720 ( .A(n8085), .B(n8084), .ZN(n8091) );
  INV_X1 U9721 ( .A(n8359), .ZN(n8087) );
  OAI22_X1 U9722 ( .A1(n9840), .A2(n8087), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8086), .ZN(n8089) );
  OAI22_X1 U9723 ( .A1(n8356), .A2(n9831), .B1(n9832), .B2(n8357), .ZN(n8088)
         );
  AOI211_X1 U9724 ( .C1(n8581), .C2(n8158), .A(n8089), .B(n8088), .ZN(n8090)
         );
  OAI21_X1 U9725 ( .B1(n8091), .B2(n9826), .A(n8090), .ZN(P2_U3227) );
  OAI21_X1 U9726 ( .B1(n4479), .B2(n8093), .A(n8092), .ZN(n8094) );
  NAND2_X1 U9727 ( .A1(n8094), .A2(n8138), .ZN(n8099) );
  INV_X1 U9728 ( .A(n8095), .ZN(n8097) );
  OAI22_X1 U9729 ( .A1(n8503), .A2(n9831), .B1(n9832), .B2(n8501), .ZN(n8096)
         );
  AOI211_X1 U9730 ( .C1(n8515), .C2(n8144), .A(n8097), .B(n8096), .ZN(n8098)
         );
  OAI211_X1 U9731 ( .C1(n4650), .C2(n9829), .A(n8099), .B(n8098), .ZN(P2_U3228) );
  XNOR2_X1 U9732 ( .A(n8101), .B(n8100), .ZN(n8106) );
  INV_X1 U9733 ( .A(n8154), .ZN(n8532) );
  AOI22_X1 U9734 ( .A1(n8532), .A2(n8530), .B1(n8533), .B2(n8461), .ZN(n8487)
         );
  OAI22_X1 U9735 ( .A1(n8142), .A2(n8487), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8102), .ZN(n8103) );
  AOI21_X1 U9736 ( .B1(n8493), .B2(n8144), .A(n8103), .ZN(n8105) );
  NAND2_X1 U9737 ( .A1(n8622), .A2(n8158), .ZN(n8104) );
  OAI211_X1 U9738 ( .C1(n8106), .C2(n9826), .A(n8105), .B(n8104), .ZN(P2_U3230) );
  XNOR2_X1 U9739 ( .A(n8108), .B(n8107), .ZN(n8112) );
  OAI22_X1 U9740 ( .A1(n9840), .A2(n8368), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10119), .ZN(n8110) );
  OAI22_X1 U9741 ( .A1(n8414), .A2(n9831), .B1(n9832), .B2(n8140), .ZN(n8109)
         );
  AOI211_X1 U9742 ( .C1(n8584), .C2(n8158), .A(n8110), .B(n8109), .ZN(n8111)
         );
  OAI21_X1 U9743 ( .B1(n8112), .B2(n9826), .A(n8111), .ZN(P2_U3231) );
  XNOR2_X1 U9744 ( .A(n8114), .B(n8113), .ZN(n8119) );
  INV_X1 U9745 ( .A(n8445), .ZN(n8115) );
  OAI22_X1 U9746 ( .A1(n9840), .A2(n8115), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10067), .ZN(n8117) );
  OAI22_X1 U9747 ( .A1(n8277), .A2(n9831), .B1(n9832), .B2(n8413), .ZN(n8116)
         );
  AOI211_X1 U9748 ( .C1(n8605), .C2(n8158), .A(n8117), .B(n8116), .ZN(n8118)
         );
  OAI21_X1 U9749 ( .B1(n8119), .B2(n9826), .A(n8118), .ZN(P2_U3235) );
  OAI21_X1 U9750 ( .B1(n8122), .B2(n8121), .A(n8120), .ZN(n8123) );
  NAND2_X1 U9751 ( .A1(n8123), .A2(n8138), .ZN(n8127) );
  NOR2_X1 U9752 ( .A1(n9840), .A2(n8404), .ZN(n8125) );
  OAI22_X1 U9753 ( .A1(n8413), .A2(n9831), .B1(n9832), .B2(n8414), .ZN(n8124)
         );
  AOI211_X1 U9754 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(n8130), .A(n8125), .B(
        n8124), .ZN(n8126) );
  OAI211_X1 U9755 ( .C1(n8407), .C2(n9829), .A(n8127), .B(n8126), .ZN(P2_U3237) );
  XNOR2_X1 U9756 ( .A(n8129), .B(n8128), .ZN(n8134) );
  AND2_X1 U9757 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8234) );
  OAI22_X1 U9758 ( .A1(n8501), .A2(n9831), .B1(n9832), .B2(n8277), .ZN(n8131)
         );
  AOI211_X1 U9759 ( .C1(n8144), .C2(n8469), .A(n8234), .B(n8131), .ZN(n8133)
         );
  NAND2_X1 U9760 ( .A1(n8615), .A2(n8158), .ZN(n8132) );
  OAI211_X1 U9761 ( .C1(n8134), .C2(n9826), .A(n8133), .B(n8132), .ZN(P2_U3240) );
  NAND2_X1 U9762 ( .A1(n8136), .A2(n8135), .ZN(n8137) );
  NAND3_X1 U9763 ( .A1(n8139), .A2(n8138), .A3(n8137), .ZN(n8146) );
  INV_X1 U9764 ( .A(n8140), .ZN(n8375) );
  AOI22_X1 U9765 ( .A1(n8311), .A2(n8533), .B1(n8530), .B2(n8375), .ZN(n8339)
         );
  OAI22_X1 U9766 ( .A1(n8142), .A2(n8339), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8141), .ZN(n8143) );
  AOI21_X1 U9767 ( .B1(n8342), .B2(n8144), .A(n8143), .ZN(n8145) );
  OAI211_X1 U9768 ( .C1(n8147), .C2(n9829), .A(n8146), .B(n8145), .ZN(P2_U3242) );
  NAND2_X1 U9769 ( .A1(n8149), .A2(n8148), .ZN(n8150) );
  XOR2_X1 U9770 ( .A(n8151), .B(n8150), .Z(n8160) );
  INV_X1 U9771 ( .A(n8537), .ZN(n8153) );
  OAI22_X1 U9772 ( .A1(n9840), .A2(n8153), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8152), .ZN(n8157) );
  OAI22_X1 U9773 ( .A1(n8155), .A2(n9831), .B1(n9832), .B2(n8154), .ZN(n8156)
         );
  AOI211_X1 U9774 ( .C1(n8158), .C2(n8538), .A(n8157), .B(n8156), .ZN(n8159)
         );
  OAI21_X1 U9775 ( .B1(n8160), .B2(n9826), .A(n8159), .ZN(P2_U3243) );
  MUX2_X1 U9776 ( .A(n8161), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8177), .Z(
        P2_U3583) );
  MUX2_X1 U9777 ( .A(n8162), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8177), .Z(
        P2_U3582) );
  INV_X1 U9778 ( .A(n8163), .ZN(n8310) );
  MUX2_X1 U9779 ( .A(n8310), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8177), .Z(
        P2_U3581) );
  INV_X1 U9780 ( .A(n8286), .ZN(n8327) );
  MUX2_X1 U9781 ( .A(n8327), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8177), .Z(
        P2_U3580) );
  MUX2_X1 U9782 ( .A(n8311), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8164), .Z(
        P2_U3579) );
  INV_X1 U9783 ( .A(n8357), .ZN(n8328) );
  MUX2_X1 U9784 ( .A(n8328), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8164), .Z(
        P2_U3578) );
  MUX2_X1 U9785 ( .A(n8375), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8164), .Z(
        P2_U3577) );
  MUX2_X1 U9786 ( .A(n8395), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8164), .Z(
        P2_U3576) );
  MUX2_X1 U9787 ( .A(n8374), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8164), .Z(
        P2_U3575) );
  MUX2_X1 U9788 ( .A(n8396), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8164), .Z(
        P2_U3574) );
  INV_X1 U9789 ( .A(n8413), .ZN(n8438) );
  MUX2_X1 U9790 ( .A(n8438), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8164), .Z(
        P2_U3573) );
  INV_X1 U9791 ( .A(n8428), .ZN(n8462) );
  MUX2_X1 U9792 ( .A(n8462), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8164), .Z(
        P2_U3572) );
  MUX2_X1 U9793 ( .A(n8477), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8164), .Z(
        P2_U3571) );
  MUX2_X1 U9794 ( .A(n8461), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8164), .Z(
        P2_U3570) );
  INV_X1 U9795 ( .A(n8501), .ZN(n8476) );
  MUX2_X1 U9796 ( .A(n8476), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8164), .Z(
        P2_U3569) );
  MUX2_X1 U9797 ( .A(n8532), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8164), .Z(
        P2_U3568) );
  MUX2_X1 U9798 ( .A(n8272), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8177), .Z(
        P2_U3567) );
  MUX2_X1 U9799 ( .A(n8531), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8177), .Z(
        P2_U3566) );
  MUX2_X1 U9800 ( .A(n8165), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8177), .Z(
        P2_U3565) );
  MUX2_X1 U9801 ( .A(n8166), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8177), .Z(
        P2_U3564) );
  MUX2_X1 U9802 ( .A(n8167), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8177), .Z(
        P2_U3563) );
  MUX2_X1 U9803 ( .A(n8168), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8177), .Z(
        P2_U3562) );
  MUX2_X1 U9804 ( .A(n8169), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8177), .Z(
        P2_U3561) );
  MUX2_X1 U9805 ( .A(n8170), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8177), .Z(
        P2_U3560) );
  MUX2_X1 U9806 ( .A(n8171), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8177), .Z(
        P2_U3559) );
  MUX2_X1 U9807 ( .A(n8172), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8177), .Z(
        P2_U3558) );
  MUX2_X1 U9808 ( .A(n8173), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8177), .Z(
        P2_U3557) );
  MUX2_X1 U9809 ( .A(n8174), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8177), .Z(
        P2_U3556) );
  MUX2_X1 U9810 ( .A(n8175), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8177), .Z(
        P2_U3555) );
  MUX2_X1 U9811 ( .A(n8176), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8177), .Z(
        P2_U3554) );
  MUX2_X1 U9812 ( .A(n7409), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8177), .Z(
        P2_U3553) );
  MUX2_X1 U9813 ( .A(n5716), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8177), .Z(
        P2_U3552) );
  AND2_X1 U9814 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n8179) );
  OAI211_X1 U9815 ( .C1(n8180), .C2(n8179), .A(n8253), .B(n8178), .ZN(n8188)
         );
  AOI22_X1 U9816 ( .A1(n8235), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(n8130), .ZN(n8187) );
  NAND2_X1 U9817 ( .A1(n8256), .A2(n8181), .ZN(n8186) );
  OAI211_X1 U9818 ( .C1(n8184), .C2(n8183), .A(n8258), .B(n8182), .ZN(n8185)
         );
  NAND4_X1 U9819 ( .A1(n8188), .A2(n8187), .A3(n8186), .A4(n8185), .ZN(
        P2_U3246) );
  OAI211_X1 U9820 ( .C1(n8191), .C2(n8190), .A(n8253), .B(n8189), .ZN(n8200)
         );
  AOI22_X1 U9821 ( .A1(n8235), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n8199) );
  INV_X1 U9822 ( .A(n8192), .ZN(n8193) );
  NAND2_X1 U9823 ( .A1(n8256), .A2(n8193), .ZN(n8198) );
  OAI211_X1 U9824 ( .C1(n8196), .C2(n8195), .A(n8258), .B(n8194), .ZN(n8197)
         );
  NAND4_X1 U9825 ( .A1(n8200), .A2(n8199), .A3(n8198), .A4(n8197), .ZN(
        P2_U3247) );
  OAI21_X1 U9826 ( .B1(n8203), .B2(n8202), .A(n8201), .ZN(n8204) );
  NAND2_X1 U9827 ( .A1(n8204), .A2(n8253), .ZN(n8214) );
  AOI21_X1 U9828 ( .B1(n8235), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8205), .ZN(
        n8213) );
  NAND2_X1 U9829 ( .A1(n8256), .A2(n8206), .ZN(n8212) );
  AOI21_X1 U9830 ( .B1(n8209), .B2(n8208), .A(n8207), .ZN(n8210) );
  NAND2_X1 U9831 ( .A1(n8258), .A2(n8210), .ZN(n8211) );
  NAND4_X1 U9832 ( .A1(n8214), .A2(n8213), .A3(n8212), .A4(n8211), .ZN(
        P2_U3256) );
  OAI21_X1 U9833 ( .B1(n8217), .B2(n8216), .A(n8215), .ZN(n8218) );
  NAND2_X1 U9834 ( .A1(n8218), .A2(n8253), .ZN(n8228) );
  AOI21_X1 U9835 ( .B1(n8235), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n8219), .ZN(
        n8227) );
  OAI21_X1 U9836 ( .B1(n8222), .B2(n8221), .A(n8220), .ZN(n8223) );
  NAND2_X1 U9837 ( .A1(n8223), .A2(n8258), .ZN(n8226) );
  NAND2_X1 U9838 ( .A1(n8256), .A2(n8224), .ZN(n8225) );
  NAND4_X1 U9839 ( .A1(n8228), .A2(n8227), .A3(n8226), .A4(n8225), .ZN(
        P2_U3259) );
  AOI21_X1 U9840 ( .B1(n8238), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8229), .ZN(
        n8231) );
  INV_X1 U9841 ( .A(n8250), .ZN(n8230) );
  NOR2_X1 U9842 ( .A1(n8231), .A2(n8230), .ZN(n8247) );
  AOI21_X1 U9843 ( .B1(n8231), .B2(n8230), .A(n8247), .ZN(n8233) );
  AND2_X1 U9844 ( .A1(n8233), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8246) );
  INV_X1 U9845 ( .A(n8246), .ZN(n8232) );
  OAI211_X1 U9846 ( .C1(P2_REG2_REG_18__SCAN_IN), .C2(n8233), .A(n8253), .B(
        n8232), .ZN(n8245) );
  AOI21_X1 U9847 ( .B1(n8235), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8234), .ZN(
        n8244) );
  NAND2_X1 U9848 ( .A1(n8256), .A2(n8250), .ZN(n8243) );
  INV_X1 U9849 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8236) );
  XNOR2_X1 U9850 ( .A(n8250), .B(n8236), .ZN(n8240) );
  AOI21_X1 U9851 ( .B1(n8238), .B2(P2_REG1_REG_17__SCAN_IN), .A(n8237), .ZN(
        n8239) );
  NAND2_X1 U9852 ( .A1(n8240), .A2(n8239), .ZN(n8249) );
  OAI21_X1 U9853 ( .B1(n8240), .B2(n8239), .A(n8249), .ZN(n8241) );
  NAND2_X1 U9854 ( .A1(n8258), .A2(n8241), .ZN(n8242) );
  NAND4_X1 U9855 ( .A1(n8245), .A2(n8244), .A3(n8243), .A4(n8242), .ZN(
        P2_U3263) );
  NOR2_X1 U9856 ( .A1(n8247), .A2(n8246), .ZN(n8248) );
  XNOR2_X1 U9857 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8248), .ZN(n8255) );
  OAI21_X1 U9858 ( .B1(n8250), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8249), .ZN(
        n8251) );
  XOR2_X1 U9859 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8251), .Z(n8257) );
  INV_X1 U9860 ( .A(n8257), .ZN(n8252) );
  AOI22_X1 U9861 ( .A1(n8255), .A2(n8253), .B1(n8252), .B2(n8258), .ZN(n8259)
         );
  INV_X1 U9862 ( .A(n8260), .ZN(n8261) );
  XNOR2_X1 U9863 ( .A(n9508), .B(n8294), .ZN(n9511) );
  NAND2_X1 U9864 ( .A1(n9511), .A2(n8520), .ZN(n8266) );
  INV_X1 U9865 ( .A(n8263), .ZN(n8264) );
  AOI21_X1 U9866 ( .B1(n9860), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8264), .ZN(
        n8265) );
  OAI211_X1 U9867 ( .C1(n9508), .C2(n8496), .A(n8266), .B(n8265), .ZN(P2_U3266) );
  OR2_X1 U9868 ( .A1(n8267), .A2(n8531), .ZN(n8269) );
  AND2_X1 U9869 ( .A1(n8269), .A2(n8268), .ZN(n8270) );
  NOR2_X1 U9870 ( .A1(n8538), .A2(n8272), .ZN(n8273) );
  AOI21_X1 U9871 ( .B1(n8525), .B2(n8526), .A(n8273), .ZN(n8505) );
  NOR2_X1 U9872 ( .A1(n8615), .A2(n8461), .ZN(n8275) );
  INV_X1 U9873 ( .A(n8615), .ZN(n8471) );
  NAND2_X1 U9874 ( .A1(n8441), .A2(n8440), .ZN(n8442) );
  INV_X1 U9875 ( .A(n8605), .ZN(n8447) );
  NAND2_X1 U9876 ( .A1(n8423), .A2(n8413), .ZN(n8278) );
  NAND2_X1 U9877 ( .A1(n8349), .A2(n8280), .ZN(n8335) );
  NAND2_X1 U9878 ( .A1(n8335), .A2(n8334), .ZN(n8333) );
  OAI21_X1 U9879 ( .B1(n8328), .B2(n8576), .A(n8333), .ZN(n8316) );
  NAND2_X1 U9880 ( .A1(n8316), .A2(n8325), .ZN(n8315) );
  OAI21_X1 U9881 ( .B1(n8311), .B2(n8569), .A(n8315), .ZN(n8302) );
  OAI21_X1 U9882 ( .B1(n8327), .B2(n8564), .A(n8301), .ZN(n8281) );
  XNOR2_X1 U9883 ( .A(n8281), .B(n8282), .ZN(n8559) );
  INV_X1 U9884 ( .A(n8559), .ZN(n8300) );
  OR2_X1 U9885 ( .A1(n8286), .A2(n8502), .ZN(n8289) );
  AND2_X1 U9886 ( .A1(n8289), .A2(n5003), .ZN(n8290) );
  INV_X1 U9887 ( .A(n8292), .ZN(n8560) );
  INV_X1 U9888 ( .A(n8293), .ZN(n8304) );
  OAI21_X1 U9889 ( .B1(n8560), .B2(n8304), .A(n8294), .ZN(n8561) );
  NOR2_X1 U9890 ( .A1(n8561), .A2(n8551), .ZN(n8298) );
  AOI22_X1 U9891 ( .A1(n9860), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8295), .B2(
        n9845), .ZN(n8296) );
  OAI21_X1 U9892 ( .B1(n8560), .B2(n8496), .A(n8296), .ZN(n8297) );
  AOI211_X1 U9893 ( .C1(n8563), .C2(n8549), .A(n8298), .B(n8297), .ZN(n8299)
         );
  OAI21_X1 U9894 ( .B1(n8300), .B2(n8543), .A(n8299), .ZN(P2_U3267) );
  OAI21_X1 U9895 ( .B1(n8302), .B2(n8308), .A(n8301), .ZN(n8303) );
  INV_X1 U9896 ( .A(n8303), .ZN(n8568) );
  AOI21_X1 U9897 ( .B1(n8564), .B2(n8318), .A(n8304), .ZN(n8565) );
  INV_X1 U9898 ( .A(n8564), .ZN(n8307) );
  AOI22_X1 U9899 ( .A1(n9860), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8305), .B2(
        n9845), .ZN(n8306) );
  OAI21_X1 U9900 ( .B1(n8307), .B2(n8496), .A(n8306), .ZN(n8313) );
  OAI21_X1 U9901 ( .B1(n8568), .B2(n8543), .A(n8314), .ZN(P2_U3268) );
  OAI21_X1 U9902 ( .B1(n8316), .B2(n8325), .A(n8315), .ZN(n8317) );
  INV_X1 U9903 ( .A(n8317), .ZN(n8573) );
  INV_X1 U9904 ( .A(n8341), .ZN(n8320) );
  INV_X1 U9905 ( .A(n8318), .ZN(n8319) );
  AOI21_X1 U9906 ( .B1(n8569), .B2(n8320), .A(n8319), .ZN(n8570) );
  INV_X1 U9907 ( .A(n8321), .ZN(n8322) );
  AOI22_X1 U9908 ( .A1(n9860), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8322), .B2(
        n9845), .ZN(n8323) );
  OAI21_X1 U9909 ( .B1(n8324), .B2(n8496), .A(n8323), .ZN(n8331) );
  XNOR2_X1 U9910 ( .A(n8326), .B(n8325), .ZN(n8329) );
  AOI222_X1 U9911 ( .A1(n9843), .A2(n8329), .B1(n8328), .B2(n8530), .C1(n8327), 
        .C2(n8533), .ZN(n8572) );
  NOR2_X1 U9912 ( .A1(n8572), .A2(n9860), .ZN(n8330) );
  AOI211_X1 U9913 ( .C1(n8570), .C2(n8520), .A(n8331), .B(n8330), .ZN(n8332)
         );
  OAI21_X1 U9914 ( .B1(n8573), .B2(n8543), .A(n8332), .ZN(P2_U3269) );
  OAI21_X1 U9915 ( .B1(n8335), .B2(n8334), .A(n8333), .ZN(n8336) );
  INV_X1 U9916 ( .A(n8336), .ZN(n8578) );
  AOI22_X1 U9917 ( .A1(n8576), .A2(n9847), .B1(n9860), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8348) );
  XNOR2_X1 U9918 ( .A(n8338), .B(n8337), .ZN(n8340) );
  OAI21_X1 U9919 ( .B1(n8340), .B2(n8488), .A(n8339), .ZN(n8574) );
  AOI211_X1 U9920 ( .C1(n8576), .C2(n4657), .A(n9922), .B(n8341), .ZN(n8575)
         );
  INV_X1 U9921 ( .A(n8575), .ZN(n8345) );
  INV_X1 U9922 ( .A(n8342), .ZN(n8343) );
  OAI22_X1 U9923 ( .A1(n8345), .A2(n5050), .B1(n8344), .B2(n8343), .ZN(n8346)
         );
  OAI21_X1 U9924 ( .B1(n8574), .B2(n8346), .A(n8549), .ZN(n8347) );
  OAI211_X1 U9925 ( .C1(n8578), .C2(n8543), .A(n8348), .B(n8347), .ZN(P2_U3270) );
  OAI21_X1 U9926 ( .B1(n8351), .B2(n8350), .A(n8349), .ZN(n8352) );
  INV_X1 U9927 ( .A(n8352), .ZN(n8583) );
  XNOR2_X1 U9928 ( .A(n8354), .B(n8353), .ZN(n8355) );
  OAI222_X1 U9929 ( .A1(n8500), .A2(n8357), .B1(n8502), .B2(n8356), .C1(n8488), 
        .C2(n8355), .ZN(n8579) );
  AOI211_X1 U9930 ( .C1(n8581), .C2(n8366), .A(n9922), .B(n8358), .ZN(n8580)
         );
  NOR2_X1 U9931 ( .A1(n9860), .A2(n5050), .ZN(n8492) );
  NAND2_X1 U9932 ( .A1(n8580), .A2(n8492), .ZN(n8361) );
  AOI22_X1 U9933 ( .A1(n9860), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8359), .B2(
        n9845), .ZN(n8360) );
  OAI211_X1 U9934 ( .C1(n4655), .C2(n8496), .A(n8361), .B(n8360), .ZN(n8362)
         );
  AOI21_X1 U9935 ( .B1(n8579), .B2(n8549), .A(n8362), .ZN(n8363) );
  OAI21_X1 U9936 ( .B1(n8583), .B2(n8543), .A(n8363), .ZN(P2_U3271) );
  XNOR2_X1 U9937 ( .A(n8365), .B(n8364), .ZN(n8588) );
  INV_X1 U9938 ( .A(n8366), .ZN(n8367) );
  AOI21_X1 U9939 ( .B1(n8584), .B2(n8383), .A(n8367), .ZN(n8585) );
  INV_X1 U9940 ( .A(n8584), .ZN(n8371) );
  INV_X1 U9941 ( .A(n8368), .ZN(n8369) );
  AOI22_X1 U9942 ( .A1(n9860), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8369), .B2(
        n9845), .ZN(n8370) );
  OAI21_X1 U9943 ( .B1(n8371), .B2(n8496), .A(n8370), .ZN(n8379) );
  OAI211_X1 U9944 ( .C1(n4460), .C2(n8373), .A(n8372), .B(n9843), .ZN(n8377)
         );
  AOI22_X1 U9945 ( .A1(n8375), .A2(n8533), .B1(n8530), .B2(n8374), .ZN(n8376)
         );
  AND2_X1 U9946 ( .A1(n8377), .A2(n8376), .ZN(n8587) );
  NOR2_X1 U9947 ( .A1(n8587), .A2(n9860), .ZN(n8378) );
  AOI211_X1 U9948 ( .C1(n8585), .C2(n8520), .A(n8379), .B(n8378), .ZN(n8380)
         );
  OAI21_X1 U9949 ( .B1(n8588), .B2(n8543), .A(n8380), .ZN(P2_U3272) );
  OAI21_X1 U9950 ( .B1(n8382), .B2(n8391), .A(n8381), .ZN(n8593) );
  INV_X1 U9951 ( .A(n8402), .ZN(n8385) );
  INV_X1 U9952 ( .A(n8383), .ZN(n8384) );
  AOI21_X1 U9953 ( .B1(n8589), .B2(n8385), .A(n8384), .ZN(n8590) );
  INV_X1 U9954 ( .A(n8386), .ZN(n8387) );
  AOI22_X1 U9955 ( .A1(n9860), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8387), .B2(
        n9845), .ZN(n8388) );
  OAI21_X1 U9956 ( .B1(n8389), .B2(n8496), .A(n8388), .ZN(n8399) );
  INV_X1 U9957 ( .A(n8390), .ZN(n8412) );
  OAI21_X1 U9958 ( .B1(n8412), .B2(n8392), .A(n8391), .ZN(n8394) );
  NAND2_X1 U9959 ( .A1(n8394), .A2(n8393), .ZN(n8397) );
  AOI222_X1 U9960 ( .A1(n9843), .A2(n8397), .B1(n8396), .B2(n8530), .C1(n8395), 
        .C2(n8533), .ZN(n8592) );
  NOR2_X1 U9961 ( .A1(n8592), .A2(n9860), .ZN(n8398) );
  AOI211_X1 U9962 ( .C1(n8590), .C2(n8520), .A(n8399), .B(n8398), .ZN(n8400)
         );
  OAI21_X1 U9963 ( .B1(n8593), .B2(n8543), .A(n8400), .ZN(P2_U3273) );
  XNOR2_X1 U9964 ( .A(n8401), .B(n8409), .ZN(n8598) );
  INV_X1 U9965 ( .A(n8421), .ZN(n8403) );
  AOI21_X1 U9966 ( .B1(n8594), .B2(n8403), .A(n8402), .ZN(n8595) );
  INV_X1 U9967 ( .A(n8404), .ZN(n8405) );
  AOI22_X1 U9968 ( .A1(n9860), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8405), .B2(
        n9845), .ZN(n8406) );
  OAI21_X1 U9969 ( .B1(n8407), .B2(n8496), .A(n8406), .ZN(n8418) );
  AOI21_X1 U9970 ( .B1(n8408), .B2(n8410), .A(n8409), .ZN(n8411) );
  NOR3_X1 U9971 ( .A1(n8412), .A2(n8411), .A3(n8488), .ZN(n8416) );
  OAI22_X1 U9972 ( .A1(n8414), .A2(n8500), .B1(n8413), .B2(n8502), .ZN(n8415)
         );
  NOR2_X1 U9973 ( .A1(n8416), .A2(n8415), .ZN(n8597) );
  NOR2_X1 U9974 ( .A1(n8597), .A2(n9860), .ZN(n8417) );
  AOI211_X1 U9975 ( .C1(n8595), .C2(n8520), .A(n8418), .B(n8417), .ZN(n8419)
         );
  OAI21_X1 U9976 ( .B1(n8598), .B2(n8543), .A(n8419), .ZN(P2_U3274) );
  XNOR2_X1 U9977 ( .A(n8420), .B(n8425), .ZN(n8603) );
  AOI211_X1 U9978 ( .C1(n8601), .C2(n8443), .A(n9922), .B(n8421), .ZN(n8600)
         );
  INV_X1 U9979 ( .A(n9855), .ZN(n8434) );
  INV_X1 U9980 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8422) );
  OAI22_X1 U9981 ( .A1(n8423), .A2(n8496), .B1(n8549), .B2(n8422), .ZN(n8433)
         );
  INV_X1 U9982 ( .A(n8408), .ZN(n8424) );
  AOI21_X1 U9983 ( .B1(n8426), .B2(n8425), .A(n8424), .ZN(n8427) );
  OAI222_X1 U9984 ( .A1(n8500), .A2(n8429), .B1(n8502), .B2(n8428), .C1(n8488), 
        .C2(n8427), .ZN(n8599) );
  AOI21_X1 U9985 ( .B1(n8430), .B2(n9845), .A(n8599), .ZN(n8431) );
  NOR2_X1 U9986 ( .A1(n8431), .A2(n9860), .ZN(n8432) );
  AOI211_X1 U9987 ( .C1(n8600), .C2(n8434), .A(n8433), .B(n8432), .ZN(n8435)
         );
  OAI21_X1 U9988 ( .B1(n8543), .B2(n8603), .A(n8435), .ZN(P2_U3275) );
  NAND2_X1 U9989 ( .A1(n8458), .A2(n8436), .ZN(n8437) );
  XOR2_X1 U9990 ( .A(n8440), .B(n8437), .Z(n8439) );
  AOI222_X1 U9991 ( .A1(n9843), .A2(n8439), .B1(n8438), .B2(n8533), .C1(n8477), 
        .C2(n8530), .ZN(n8608) );
  OR2_X1 U9992 ( .A1(n8441), .A2(n8440), .ZN(n8604) );
  NAND3_X1 U9993 ( .A1(n8604), .A2(n8442), .A3(n9857), .ZN(n8450) );
  INV_X1 U9994 ( .A(n8443), .ZN(n8444) );
  AOI21_X1 U9995 ( .B1(n8605), .B2(n8452), .A(n8444), .ZN(n8606) );
  AOI22_X1 U9996 ( .A1(n9860), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8445), .B2(
        n9845), .ZN(n8446) );
  OAI21_X1 U9997 ( .B1(n8447), .B2(n8496), .A(n8446), .ZN(n8448) );
  AOI21_X1 U9998 ( .B1(n8606), .B2(n8520), .A(n8448), .ZN(n8449) );
  OAI211_X1 U9999 ( .C1(n9860), .C2(n8608), .A(n8450), .B(n8449), .ZN(P2_U3276) );
  XOR2_X1 U10000 ( .A(n8460), .B(n8451), .Z(n8614) );
  INV_X1 U10001 ( .A(n8468), .ZN(n8454) );
  INV_X1 U10002 ( .A(n8452), .ZN(n8453) );
  AOI211_X1 U10003 ( .C1(n8611), .C2(n8454), .A(n9922), .B(n8453), .ZN(n8610)
         );
  AOI22_X1 U10004 ( .A1(n9860), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8455), .B2(
        n9845), .ZN(n8456) );
  OAI21_X1 U10005 ( .B1(n8457), .B2(n8496), .A(n8456), .ZN(n8465) );
  OAI21_X1 U10006 ( .B1(n8460), .B2(n8459), .A(n8458), .ZN(n8463) );
  AOI222_X1 U10007 ( .A1(n9843), .A2(n8463), .B1(n8462), .B2(n8533), .C1(n8461), .C2(n8530), .ZN(n8613) );
  NOR2_X1 U10008 ( .A1(n8613), .A2(n9860), .ZN(n8464) );
  AOI211_X1 U10009 ( .C1(n8610), .C2(n8492), .A(n8465), .B(n8464), .ZN(n8466)
         );
  OAI21_X1 U10010 ( .B1(n8543), .B2(n8614), .A(n8466), .ZN(P2_U3277) );
  XNOR2_X1 U10011 ( .A(n8467), .B(n8474), .ZN(n8619) );
  AOI21_X1 U10012 ( .B1(n8615), .B2(n8490), .A(n8468), .ZN(n8616) );
  AOI22_X1 U10013 ( .A1(n9860), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8469), .B2(
        n9845), .ZN(n8470) );
  OAI21_X1 U10014 ( .B1(n8471), .B2(n8496), .A(n8470), .ZN(n8480) );
  INV_X1 U10015 ( .A(n8472), .ZN(n8475) );
  OAI21_X1 U10016 ( .B1(n8475), .B2(n8474), .A(n8473), .ZN(n8478) );
  AOI222_X1 U10017 ( .A1(n9843), .A2(n8478), .B1(n8477), .B2(n8533), .C1(n8476), .C2(n8530), .ZN(n8618) );
  NOR2_X1 U10018 ( .A1(n8618), .A2(n9860), .ZN(n8479) );
  AOI211_X1 U10019 ( .C1(n8616), .C2(n8520), .A(n8480), .B(n8479), .ZN(n8481)
         );
  OAI21_X1 U10020 ( .B1(n8619), .B2(n8543), .A(n8481), .ZN(P2_U3278) );
  OAI21_X1 U10021 ( .B1(n8483), .B2(n8485), .A(n8482), .ZN(n8484) );
  INV_X1 U10022 ( .A(n8484), .ZN(n8625) );
  XNOR2_X1 U10023 ( .A(n8486), .B(n8485), .ZN(n8489) );
  OAI21_X1 U10024 ( .B1(n8489), .B2(n8488), .A(n8487), .ZN(n8620) );
  INV_X1 U10025 ( .A(n8490), .ZN(n8491) );
  AOI211_X1 U10026 ( .C1(n8622), .C2(n8514), .A(n9922), .B(n8491), .ZN(n8621)
         );
  NAND2_X1 U10027 ( .A1(n8621), .A2(n8492), .ZN(n8495) );
  AOI22_X1 U10028 ( .A1(n9860), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8493), .B2(
        n9845), .ZN(n8494) );
  OAI211_X1 U10029 ( .C1(n4989), .C2(n8496), .A(n8495), .B(n8494), .ZN(n8497)
         );
  AOI21_X1 U10030 ( .B1(n8620), .B2(n8549), .A(n8497), .ZN(n8498) );
  OAI21_X1 U10031 ( .B1(n8625), .B2(n8543), .A(n8498), .ZN(P2_U3279) );
  XNOR2_X1 U10032 ( .A(n8499), .B(n8504), .ZN(n8511) );
  OAI22_X1 U10033 ( .A1(n8503), .A2(n8502), .B1(n8501), .B2(n8500), .ZN(n8510)
         );
  NOR2_X1 U10034 ( .A1(n8505), .A2(n8504), .ZN(n8506) );
  NOR2_X1 U10035 ( .A1(n8630), .A2(n8508), .ZN(n8509) );
  AOI211_X1 U10036 ( .C1(n9843), .C2(n8511), .A(n8510), .B(n8509), .ZN(n8629)
         );
  NAND2_X1 U10037 ( .A1(n8512), .A2(n8626), .ZN(n8513) );
  AND2_X1 U10038 ( .A1(n8514), .A2(n8513), .ZN(n8627) );
  INV_X1 U10039 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8518) );
  NAND2_X1 U10040 ( .A1(n8626), .A2(n9847), .ZN(n8517) );
  NAND2_X1 U10041 ( .A1(n9845), .A2(n8515), .ZN(n8516) );
  OAI211_X1 U10042 ( .C1(n8549), .C2(n8518), .A(n8517), .B(n8516), .ZN(n8519)
         );
  AOI21_X1 U10043 ( .B1(n8627), .B2(n8520), .A(n8519), .ZN(n8524) );
  INV_X1 U10044 ( .A(n8630), .ZN(n8522) );
  NAND2_X1 U10045 ( .A1(n8522), .A2(n8521), .ZN(n8523) );
  OAI211_X1 U10046 ( .C1(n8629), .C2(n9860), .A(n8524), .B(n8523), .ZN(
        P2_U3280) );
  XNOR2_X1 U10047 ( .A(n8525), .B(n8526), .ZN(n9517) );
  INV_X1 U10048 ( .A(n9517), .ZN(n8544) );
  OAI211_X1 U10049 ( .C1(n8529), .C2(n8528), .A(n8527), .B(n9843), .ZN(n8535)
         );
  AOI22_X1 U10050 ( .A1(n8533), .A2(n8532), .B1(n8531), .B2(n8530), .ZN(n8534)
         );
  NAND2_X1 U10051 ( .A1(n8535), .A2(n8534), .ZN(n9515) );
  XNOR2_X1 U10052 ( .A(n8536), .B(n9513), .ZN(n9514) );
  AOI22_X1 U10053 ( .A1(n9860), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8537), .B2(
        n9845), .ZN(n8540) );
  NAND2_X1 U10054 ( .A1(n9847), .A2(n8538), .ZN(n8539) );
  OAI211_X1 U10055 ( .C1(n9514), .C2(n8551), .A(n8540), .B(n8539), .ZN(n8541)
         );
  AOI21_X1 U10056 ( .B1(n9515), .B2(n8549), .A(n8541), .ZN(n8542) );
  OAI21_X1 U10057 ( .B1(n8544), .B2(n8543), .A(n8542), .ZN(P2_U3281) );
  AOI22_X1 U10058 ( .A1(n9857), .A2(n8546), .B1(n9847), .B2(n8545), .ZN(n8555)
         );
  AOI22_X1 U10059 ( .A1(n8547), .A2(n8549), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n9845), .ZN(n8554) );
  OAI22_X1 U10060 ( .A1(n8551), .A2(n8550), .B1(n8549), .B2(n8548), .ZN(n8552)
         );
  INV_X1 U10061 ( .A(n8552), .ZN(n8553) );
  NAND3_X1 U10062 ( .A1(n8555), .A2(n8554), .A3(n8553), .ZN(P2_U3294) );
  AOI21_X1 U10063 ( .B1(n8556), .B2(n9886), .A(n9510), .ZN(n8557) );
  MUX2_X1 U10064 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8631), .S(n9945), .Z(
        P2_U3551) );
  OAI22_X1 U10065 ( .A1(n8561), .A2(n9922), .B1(n9921), .B2(n8560), .ZN(n8562)
         );
  AOI22_X1 U10066 ( .A1(n8565), .A2(n9853), .B1(n9886), .B2(n8564), .ZN(n8566)
         );
  OAI211_X1 U10067 ( .C1(n8568), .C2(n8624), .A(n8567), .B(n8566), .ZN(n8633)
         );
  MUX2_X1 U10068 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8633), .S(n9945), .Z(
        P2_U3548) );
  AOI22_X1 U10069 ( .A1(n8570), .A2(n9853), .B1(n8569), .B2(n9886), .ZN(n8571)
         );
  OAI211_X1 U10070 ( .C1(n8573), .C2(n8624), .A(n8572), .B(n8571), .ZN(n8634)
         );
  MUX2_X1 U10071 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8634), .S(n9945), .Z(
        P2_U3547) );
  AOI211_X1 U10072 ( .C1(n8576), .C2(n9886), .A(n8575), .B(n8574), .ZN(n8577)
         );
  OAI21_X1 U10073 ( .B1(n8578), .B2(n8624), .A(n8577), .ZN(n8635) );
  MUX2_X1 U10074 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8635), .S(n9945), .Z(
        P2_U3546) );
  AOI211_X1 U10075 ( .C1(n8581), .C2(n9886), .A(n8580), .B(n8579), .ZN(n8582)
         );
  OAI21_X1 U10076 ( .B1(n8583), .B2(n8624), .A(n8582), .ZN(n8636) );
  MUX2_X1 U10077 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8636), .S(n9945), .Z(
        P2_U3545) );
  AOI22_X1 U10078 ( .A1(n8585), .A2(n9853), .B1(n8584), .B2(n9886), .ZN(n8586)
         );
  OAI211_X1 U10079 ( .C1(n8588), .C2(n8624), .A(n8587), .B(n8586), .ZN(n8637)
         );
  MUX2_X1 U10080 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8637), .S(n9945), .Z(
        P2_U3544) );
  AOI22_X1 U10081 ( .A1(n8590), .A2(n9853), .B1(n8589), .B2(n9886), .ZN(n8591)
         );
  OAI211_X1 U10082 ( .C1(n8593), .C2(n8624), .A(n8592), .B(n8591), .ZN(n8638)
         );
  MUX2_X1 U10083 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8638), .S(n9945), .Z(
        P2_U3543) );
  AOI22_X1 U10084 ( .A1(n8595), .A2(n9853), .B1(n8594), .B2(n9886), .ZN(n8596)
         );
  OAI211_X1 U10085 ( .C1(n8598), .C2(n8624), .A(n8597), .B(n8596), .ZN(n8639)
         );
  MUX2_X1 U10086 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8639), .S(n9945), .Z(
        P2_U3542) );
  AOI211_X1 U10087 ( .C1(n8601), .C2(n9886), .A(n8600), .B(n8599), .ZN(n8602)
         );
  OAI21_X1 U10088 ( .B1(n8603), .B2(n8624), .A(n8602), .ZN(n8640) );
  MUX2_X1 U10089 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8640), .S(n9945), .Z(
        P2_U3541) );
  NAND3_X1 U10090 ( .A1(n8604), .A2(n8442), .A3(n9927), .ZN(n8609) );
  AOI22_X1 U10091 ( .A1(n8606), .A2(n9853), .B1(n8605), .B2(n9886), .ZN(n8607)
         );
  NAND3_X1 U10092 ( .A1(n8609), .A2(n8608), .A3(n8607), .ZN(n8641) );
  MUX2_X1 U10093 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8641), .S(n9945), .Z(
        P2_U3540) );
  AOI21_X1 U10094 ( .B1(n8611), .B2(n9886), .A(n8610), .ZN(n8612) );
  OAI211_X1 U10095 ( .C1(n8614), .C2(n8624), .A(n8613), .B(n8612), .ZN(n8642)
         );
  MUX2_X1 U10096 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8642), .S(n9945), .Z(
        P2_U3539) );
  AOI22_X1 U10097 ( .A1(n8616), .A2(n9853), .B1(n8615), .B2(n9886), .ZN(n8617)
         );
  OAI211_X1 U10098 ( .C1(n8619), .C2(n8624), .A(n8618), .B(n8617), .ZN(n8643)
         );
  MUX2_X1 U10099 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8643), .S(n9945), .Z(
        P2_U3538) );
  AOI211_X1 U10100 ( .C1(n8622), .C2(n9886), .A(n8621), .B(n8620), .ZN(n8623)
         );
  OAI21_X1 U10101 ( .B1(n8625), .B2(n8624), .A(n8623), .ZN(n8644) );
  MUX2_X1 U10102 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8644), .S(n9945), .Z(
        P2_U3537) );
  AOI22_X1 U10103 ( .A1(n8627), .A2(n9853), .B1(n8626), .B2(n9886), .ZN(n8628)
         );
  OAI211_X1 U10104 ( .C1(n9524), .C2(n8630), .A(n8629), .B(n8628), .ZN(n8645)
         );
  MUX2_X1 U10105 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8645), .S(n9945), .Z(
        P2_U3536) );
  MUX2_X1 U10106 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8631), .S(n9930), .Z(
        P2_U3519) );
  MUX2_X1 U10107 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8633), .S(n9930), .Z(
        P2_U3516) );
  MUX2_X1 U10108 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8634), .S(n9930), .Z(
        P2_U3515) );
  MUX2_X1 U10109 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8635), .S(n9930), .Z(
        P2_U3514) );
  MUX2_X1 U10110 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8636), .S(n9930), .Z(
        P2_U3513) );
  MUX2_X1 U10111 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8637), .S(n9930), .Z(
        P2_U3512) );
  MUX2_X1 U10112 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8638), .S(n9930), .Z(
        P2_U3511) );
  MUX2_X1 U10113 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8639), .S(n9930), .Z(
        P2_U3510) );
  MUX2_X1 U10114 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8640), .S(n9930), .Z(
        P2_U3509) );
  MUX2_X1 U10115 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8641), .S(n9930), .Z(
        P2_U3508) );
  MUX2_X1 U10116 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8642), .S(n9930), .Z(
        P2_U3507) );
  MUX2_X1 U10117 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8643), .S(n9930), .Z(
        P2_U3505) );
  MUX2_X1 U10118 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8644), .S(n9930), .Z(
        P2_U3502) );
  MUX2_X1 U10119 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8645), .S(n9930), .Z(
        P2_U3499) );
  OAI222_X1 U10120 ( .A1(n8025), .A2(n8647), .B1(n8130), .B2(n8646), .C1(
        n10222), .C2(n8651), .ZN(P2_U3330) );
  MUX2_X1 U10121 ( .A(n8652), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10122 ( .A(n8655), .B(n8654), .ZN(n8656) );
  XNOR2_X1 U10123 ( .A(n8653), .B(n8656), .ZN(n8662) );
  NAND2_X1 U10124 ( .A1(n8749), .A2(n9214), .ZN(n8658) );
  AOI22_X1 U10125 ( .A1(n8739), .A2(n9389), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8657) );
  OAI211_X1 U10126 ( .C1(n8659), .C2(n8737), .A(n8658), .B(n8657), .ZN(n8660)
         );
  AOI21_X1 U10127 ( .B1(n9220), .B2(n8730), .A(n8660), .ZN(n8661) );
  OAI21_X1 U10128 ( .B1(n8662), .B2(n7995), .A(n8661), .ZN(P1_U3214) );
  XNOR2_X1 U10129 ( .A(n8665), .B(n8664), .ZN(n8666) );
  XNOR2_X1 U10130 ( .A(n8663), .B(n8666), .ZN(n8671) );
  NAND2_X1 U10131 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9108) );
  OAI21_X1 U10132 ( .B1(n8759), .B2(n9317), .A(n9108), .ZN(n8667) );
  AOI21_X1 U10133 ( .B1(n8762), .B2(n9412), .A(n8667), .ZN(n8668) );
  OAI21_X1 U10134 ( .B1(n8765), .B2(n9278), .A(n8668), .ZN(n8669) );
  AOI21_X1 U10135 ( .B1(n9289), .B2(n8730), .A(n8669), .ZN(n8670) );
  OAI21_X1 U10136 ( .B1(n8671), .B2(n7995), .A(n8670), .ZN(P1_U3217) );
  NAND2_X1 U10137 ( .A1(n4480), .A2(n8672), .ZN(n8673) );
  XNOR2_X1 U10138 ( .A(n8674), .B(n8673), .ZN(n8679) );
  NAND2_X1 U10139 ( .A1(n8749), .A2(n9250), .ZN(n8676) );
  AOI22_X1 U10140 ( .A1(n8739), .A2(n9412), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8675) );
  OAI211_X1 U10141 ( .C1(n9247), .C2(n8737), .A(n8676), .B(n8675), .ZN(n8677)
         );
  AOI21_X1 U10142 ( .B1(n9249), .B2(n8767), .A(n8677), .ZN(n8678) );
  OAI21_X1 U10143 ( .B1(n8679), .B2(n7995), .A(n8678), .ZN(P1_U3221) );
  NAND2_X1 U10144 ( .A1(n4469), .A2(n8680), .ZN(n8681) );
  XNOR2_X1 U10145 ( .A(n8682), .B(n8681), .ZN(n8687) );
  NAND2_X1 U10146 ( .A1(n8749), .A2(n9186), .ZN(n8684) );
  AOI22_X1 U10147 ( .A1(n8739), .A2(n9388), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8683) );
  OAI211_X1 U10148 ( .C1(n9148), .C2(n8737), .A(n8684), .B(n8683), .ZN(n8685)
         );
  AOI21_X1 U10149 ( .B1(n9185), .B2(n8767), .A(n8685), .ZN(n8686) );
  OAI21_X1 U10150 ( .B1(n8687), .B2(n7995), .A(n8686), .ZN(P1_U3223) );
  AOI21_X1 U10151 ( .B1(n8690), .B2(n8689), .A(n8688), .ZN(n8696) );
  NAND2_X1 U10152 ( .A1(n8749), .A2(n9334), .ZN(n8692) );
  AOI22_X1 U10153 ( .A1(n8739), .A2(n9540), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3084), .ZN(n8691) );
  OAI211_X1 U10154 ( .C1(n8693), .C2(n8737), .A(n8692), .B(n8691), .ZN(n8694)
         );
  AOI21_X1 U10155 ( .B1(n9539), .B2(n8767), .A(n8694), .ZN(n8695) );
  OAI21_X1 U10156 ( .B1(n8696), .B2(n7995), .A(n8695), .ZN(P1_U3224) );
  XOR2_X1 U10157 ( .A(n8698), .B(n8697), .Z(n8704) );
  OAI22_X1 U10158 ( .A1(n8759), .A2(n9316), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8699), .ZN(n8700) );
  AOI21_X1 U10159 ( .B1(n8762), .B2(n9411), .A(n8700), .ZN(n8701) );
  OAI21_X1 U10160 ( .B1(n8765), .B2(n9322), .A(n8701), .ZN(n8702) );
  AOI21_X1 U10161 ( .B1(n9428), .B2(n8767), .A(n8702), .ZN(n8703) );
  OAI21_X1 U10162 ( .B1(n8704), .B2(n7995), .A(n8703), .ZN(P1_U3226) );
  INV_X1 U10163 ( .A(n8705), .ZN(n8706) );
  AOI21_X1 U10164 ( .B1(n8708), .B2(n8707), .A(n8706), .ZN(n8713) );
  NAND2_X1 U10165 ( .A1(n8749), .A2(n9200), .ZN(n8710) );
  AOI22_X1 U10166 ( .A1(n8739), .A2(n9228), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8709) );
  OAI211_X1 U10167 ( .C1(n9197), .C2(n8737), .A(n8710), .B(n8709), .ZN(n8711)
         );
  AOI21_X1 U10168 ( .B1(n9199), .B2(n8730), .A(n8711), .ZN(n8712) );
  OAI21_X1 U10169 ( .B1(n8713), .B2(n7995), .A(n8712), .ZN(P1_U3227) );
  NOR2_X1 U10170 ( .A1(n8716), .A2(n4849), .ZN(n8717) );
  XNOR2_X1 U10171 ( .A(n4843), .B(n8717), .ZN(n8722) );
  AOI22_X1 U10172 ( .A1(n8739), .A2(n9295), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8719) );
  NAND2_X1 U10173 ( .A1(n8762), .A2(n9260), .ZN(n8718) );
  OAI211_X1 U10174 ( .C1(n8765), .C2(n9266), .A(n8719), .B(n8718), .ZN(n8720)
         );
  AOI21_X1 U10175 ( .B1(n9265), .B2(n8730), .A(n8720), .ZN(n8721) );
  OAI21_X1 U10176 ( .B1(n8722), .B2(n7995), .A(n8721), .ZN(P1_U3231) );
  NAND2_X1 U10177 ( .A1(n8724), .A2(n8723), .ZN(n8726) );
  XNOR2_X1 U10178 ( .A(n8726), .B(n8725), .ZN(n8732) );
  NAND2_X1 U10179 ( .A1(n8749), .A2(n9232), .ZN(n8728) );
  AOI22_X1 U10180 ( .A1(n8739), .A2(n9260), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8727) );
  OAI211_X1 U10181 ( .C1(n9196), .C2(n8737), .A(n8728), .B(n8727), .ZN(n8729)
         );
  AOI21_X1 U10182 ( .B1(n4695), .B2(n8730), .A(n8729), .ZN(n8731) );
  OAI21_X1 U10183 ( .B1(n8732), .B2(n7995), .A(n8731), .ZN(P1_U3233) );
  XNOR2_X1 U10184 ( .A(n5007), .B(n8733), .ZN(n8734) );
  XNOR2_X1 U10185 ( .A(n8735), .B(n8734), .ZN(n8743) );
  NAND2_X1 U10186 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9091) );
  OAI21_X1 U10187 ( .B1(n8737), .B2(n8736), .A(n9091), .ZN(n8738) );
  AOI21_X1 U10188 ( .B1(n8739), .B2(n9541), .A(n8738), .ZN(n8740) );
  OAI21_X1 U10189 ( .B1(n8765), .B2(n9302), .A(n8740), .ZN(n8741) );
  AOI21_X1 U10190 ( .B1(n9421), .B2(n8767), .A(n8741), .ZN(n8742) );
  OAI21_X1 U10191 ( .B1(n8743), .B2(n7995), .A(n8742), .ZN(P1_U3236) );
  AOI22_X1 U10192 ( .A1(n8762), .A2(n9160), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8747) );
  OAI21_X1 U10193 ( .B1(n9197), .B2(n8759), .A(n8747), .ZN(n8748) );
  AOI21_X1 U10194 ( .B1(n9167), .B2(n8749), .A(n8748), .ZN(n8750) );
  INV_X1 U10195 ( .A(n8752), .ZN(n8754) );
  NAND2_X1 U10196 ( .A1(n8754), .A2(n8753), .ZN(n8756) );
  XNOR2_X1 U10197 ( .A(n8756), .B(n8755), .ZN(n8770) );
  INV_X1 U10198 ( .A(n8757), .ZN(n8761) );
  NOR2_X1 U10199 ( .A1(n8759), .A2(n8758), .ZN(n8760) );
  AOI211_X1 U10200 ( .C1(n8762), .C2(n9431), .A(n8761), .B(n8760), .ZN(n8763)
         );
  OAI21_X1 U10201 ( .B1(n8765), .B2(n8764), .A(n8763), .ZN(n8766) );
  AOI21_X1 U10202 ( .B1(n8768), .B2(n8767), .A(n8766), .ZN(n8769) );
  OAI21_X1 U10203 ( .B1(n8770), .B2(n7995), .A(n8769), .ZN(P1_U3239) );
  INV_X1 U10204 ( .A(n8771), .ZN(n8773) );
  NAND2_X1 U10205 ( .A1(n6254), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8774) );
  NAND2_X1 U10206 ( .A1(n8776), .A2(n8780), .ZN(n8778) );
  NAND2_X1 U10207 ( .A1(n6266), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8777) );
  OR2_X1 U10208 ( .A1(n9137), .A2(n9117), .ZN(n8779) );
  NAND2_X1 U10209 ( .A1(n8781), .A2(n8780), .ZN(n8783) );
  NAND2_X1 U10210 ( .A1(n6266), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8782) );
  OR2_X1 U10211 ( .A1(n9127), .A2(n8942), .ZN(n8784) );
  AND2_X1 U10212 ( .A1(n8784), .A2(n8939), .ZN(n8829) );
  INV_X1 U10213 ( .A(n8829), .ZN(n9016) );
  NAND2_X1 U10214 ( .A1(n9224), .A2(n8913), .ZN(n8785) );
  AND2_X1 U10215 ( .A1(n8785), .A2(n8917), .ZN(n8786) );
  NAND2_X1 U10216 ( .A1(n8961), .A2(n8786), .ZN(n8927) );
  INV_X1 U10217 ( .A(n8927), .ZN(n8787) );
  AND3_X1 U10218 ( .A1(n8787), .A2(n8958), .A3(n8914), .ZN(n8820) );
  INV_X1 U10219 ( .A(n8820), .ZN(n8794) );
  NAND2_X1 U10220 ( .A1(n8906), .A2(n8788), .ZN(n8814) );
  NAND2_X1 U10221 ( .A1(n8896), .A2(n8891), .ZN(n8811) );
  INV_X1 U10222 ( .A(n8869), .ZN(n8789) );
  OAI211_X1 U10223 ( .C1(n8789), .C2(n8867), .A(n8872), .B(n8871), .ZN(n8790)
         );
  INV_X1 U10224 ( .A(n8790), .ZN(n8791) );
  AND2_X1 U10225 ( .A1(n8791), .A2(n8873), .ZN(n8876) );
  NAND4_X1 U10226 ( .A1(n8890), .A2(n8876), .A3(n8875), .A4(n8861), .ZN(n8792)
         );
  OR3_X1 U10227 ( .A1(n8814), .A2(n8811), .A3(n8792), .ZN(n8793) );
  OR2_X1 U10228 ( .A1(n8794), .A2(n8793), .ZN(n8823) );
  INV_X1 U10229 ( .A(n8823), .ZN(n9009) );
  NAND2_X1 U10230 ( .A1(n8795), .A2(n8968), .ZN(n8796) );
  AOI211_X1 U10231 ( .C1(n9732), .C2(n6589), .A(n8954), .B(n8796), .ZN(n8798)
         );
  INV_X1 U10232 ( .A(n8850), .ZN(n8797) );
  NOR3_X1 U10233 ( .A1(n8798), .A2(n9006), .A3(n8797), .ZN(n8801) );
  AND2_X1 U10234 ( .A1(n8971), .A2(n8799), .ZN(n8978) );
  INV_X1 U10235 ( .A(n8978), .ZN(n8800) );
  OAI211_X1 U10236 ( .C1(n8801), .C2(n8800), .A(n8849), .B(n8973), .ZN(n8802)
         );
  AOI21_X1 U10237 ( .B1(n8802), .B2(n8977), .A(n4596), .ZN(n8824) );
  AND2_X1 U10238 ( .A1(n8976), .A2(n8865), .ZN(n8859) );
  NAND2_X1 U10239 ( .A1(n8902), .A2(n8803), .ZN(n8897) );
  AND2_X1 U10240 ( .A1(n8894), .A2(n8804), .ZN(n8885) );
  INV_X1 U10241 ( .A(n8885), .ZN(n8809) );
  INV_X1 U10242 ( .A(n8873), .ZN(n8887) );
  INV_X1 U10243 ( .A(n8876), .ZN(n8806) );
  AND3_X1 U10244 ( .A1(n8869), .A2(n8864), .A3(n8868), .ZN(n8805) );
  OR2_X1 U10245 ( .A1(n8806), .A2(n8805), .ZN(n8878) );
  OAI21_X1 U10246 ( .B1(n8888), .B2(n8887), .A(n8878), .ZN(n8807) );
  AND2_X1 U10247 ( .A1(n8807), .A2(n8890), .ZN(n8808) );
  NOR2_X1 U10248 ( .A1(n8809), .A2(n8808), .ZN(n8810) );
  NOR2_X1 U10249 ( .A1(n8811), .A2(n8810), .ZN(n8812) );
  NOR2_X1 U10250 ( .A1(n8897), .A2(n8812), .ZN(n8813) );
  NOR2_X1 U10251 ( .A1(n8814), .A2(n8813), .ZN(n8819) );
  AND2_X1 U10252 ( .A1(n8914), .A2(n8906), .ZN(n8924) );
  INV_X1 U10253 ( .A(n8924), .ZN(n8815) );
  AND2_X1 U10254 ( .A1(n8962), .A2(n8911), .ZN(n8922) );
  OAI211_X1 U10255 ( .C1(n8907), .C2(n8815), .A(n9224), .B(n8922), .ZN(n8816)
         );
  INV_X1 U10256 ( .A(n8816), .ZN(n8817) );
  OAI21_X1 U10257 ( .B1(n8927), .B2(n8817), .A(n8960), .ZN(n8818) );
  AOI22_X1 U10258 ( .A1(n8820), .A2(n8819), .B1(n8958), .B2(n8818), .ZN(n8822)
         );
  NAND2_X1 U10259 ( .A1(n8956), .A2(n8959), .ZN(n8842) );
  INV_X1 U10260 ( .A(n8842), .ZN(n8821) );
  OAI211_X1 U10261 ( .C1(n8859), .C2(n8823), .A(n8822), .B(n8821), .ZN(n9007)
         );
  AOI21_X1 U10262 ( .B1(n9009), .B2(n8824), .A(n9007), .ZN(n8826) );
  NAND2_X1 U10263 ( .A1(n8932), .A2(n8957), .ZN(n9011) );
  OAI211_X1 U10264 ( .C1(n8826), .C2(n9011), .A(n4825), .B(n4823), .ZN(n8832)
         );
  OAI211_X1 U10265 ( .C1(n8827), .C2(n8837), .A(n9132), .B(n8835), .ZN(n8828)
         );
  AOI22_X1 U10266 ( .A1(n8829), .A2(n8828), .B1(n8942), .B2(n9127), .ZN(n9014)
         );
  NOR2_X1 U10267 ( .A1(n9447), .A2(n8830), .ZN(n8999) );
  INV_X1 U10268 ( .A(n8999), .ZN(n8831) );
  OAI211_X1 U10269 ( .C1(n9016), .C2(n8832), .A(n9014), .B(n8831), .ZN(n8834)
         );
  AND2_X1 U10270 ( .A1(n9443), .A2(n8833), .ZN(n9017) );
  AOI21_X1 U10271 ( .B1(n4428), .B2(n8834), .A(n9017), .ZN(n9027) );
  NOR2_X1 U10272 ( .A1(n9027), .A2(n9215), .ZN(n9026) );
  OAI21_X1 U10273 ( .B1(n9137), .B2(n9113), .A(n9117), .ZN(n9013) );
  INV_X1 U10274 ( .A(n9019), .ZN(n8951) );
  MUX2_X1 U10275 ( .A(n8835), .B(n9010), .S(n8944), .Z(n8938) );
  MUX2_X1 U10276 ( .A(n8837), .B(n8836), .S(n8949), .Z(n8936) );
  NAND2_X1 U10277 ( .A1(n8957), .A2(n8842), .ZN(n8839) );
  NAND2_X1 U10278 ( .A1(n8839), .A2(n9175), .ZN(n8929) );
  NOR2_X1 U10279 ( .A1(n9228), .A2(n8944), .ZN(n8840) );
  AOI22_X1 U10280 ( .A1(n8841), .A2(n8949), .B1(n8840), .B2(n9220), .ZN(n8921)
         );
  NAND4_X1 U10281 ( .A1(n8932), .A2(n8944), .A3(n8842), .A4(n8957), .ZN(n8920)
         );
  NAND3_X1 U10282 ( .A1(n8843), .A2(n8971), .A3(n8949), .ZN(n8856) );
  OAI21_X1 U10283 ( .B1(n9768), .B2(n8944), .A(n8845), .ZN(n8844) );
  OAI21_X1 U10284 ( .B1(n9768), .B2(n8845), .A(n8844), .ZN(n8846) );
  OAI21_X1 U10285 ( .B1(n8849), .B2(n8944), .A(n8846), .ZN(n8847) );
  INV_X1 U10286 ( .A(n8847), .ZN(n8855) );
  AND2_X1 U10287 ( .A1(n8973), .A2(n8944), .ZN(n8851) );
  INV_X1 U10288 ( .A(n8851), .ZN(n8848) );
  OR2_X1 U10289 ( .A1(n8848), .A2(n8971), .ZN(n8854) );
  AND2_X1 U10290 ( .A1(n8850), .A2(n8849), .ZN(n8970) );
  NAND3_X1 U10291 ( .A1(n8852), .A2(n8851), .A3(n8970), .ZN(n8853) );
  NAND4_X1 U10292 ( .A1(n8856), .A2(n8855), .A3(n8854), .A4(n8853), .ZN(n8858)
         );
  NAND2_X1 U10293 ( .A1(n8863), .A2(n8859), .ZN(n8860) );
  NAND2_X1 U10294 ( .A1(n8860), .A2(n8861), .ZN(n8866) );
  INV_X1 U10295 ( .A(n8977), .ZN(n8862) );
  NAND3_X1 U10296 ( .A1(n8874), .A2(n8867), .A3(n8875), .ZN(n8870) );
  AND2_X1 U10297 ( .A1(n8873), .A2(n8872), .ZN(n8882) );
  INV_X1 U10298 ( .A(n8874), .ZN(n8877) );
  NAND3_X1 U10299 ( .A1(n8877), .A2(n8876), .A3(n8875), .ZN(n8880) );
  NAND4_X1 U10300 ( .A1(n8880), .A2(n8944), .A3(n8879), .A4(n8878), .ZN(n8881)
         );
  AOI21_X1 U10301 ( .B1(n8889), .B2(n8882), .A(n8881), .ZN(n8884) );
  OR2_X1 U10302 ( .A1(n8884), .A2(n8883), .ZN(n8893) );
  NAND2_X1 U10303 ( .A1(n8893), .A2(n8885), .ZN(n8886) );
  NAND2_X1 U10304 ( .A1(n8886), .A2(n8891), .ZN(n8895) );
  AOI21_X1 U10305 ( .B1(n8889), .B2(n8888), .A(n8887), .ZN(n8892) );
  NAND2_X1 U10306 ( .A1(n9312), .A2(n8896), .ZN(n8898) );
  MUX2_X1 U10307 ( .A(n8898), .B(n8897), .S(n8949), .Z(n8899) );
  INV_X1 U10308 ( .A(n8899), .ZN(n8900) );
  NAND2_X1 U10309 ( .A1(n8901), .A2(n8900), .ZN(n8904) );
  MUX2_X1 U10310 ( .A(n8902), .B(n9312), .S(n8949), .Z(n8903) );
  NAND3_X1 U10311 ( .A1(n8904), .A2(n9310), .A3(n8903), .ZN(n8910) );
  AND2_X1 U10312 ( .A1(n8906), .A2(n8905), .ZN(n8908) );
  MUX2_X1 U10313 ( .A(n8908), .B(n8907), .S(n8949), .Z(n8909) );
  NAND2_X1 U10314 ( .A1(n8910), .A2(n8909), .ZN(n8925) );
  NAND3_X1 U10315 ( .A1(n8925), .A2(n8912), .A3(n8911), .ZN(n8915) );
  INV_X1 U10316 ( .A(n8913), .ZN(n8963) );
  NAND3_X1 U10317 ( .A1(n8915), .A2(n8914), .A3(n8963), .ZN(n8916) );
  OAI211_X1 U10318 ( .C1(n8929), .C2(n8921), .A(n8920), .B(n8919), .ZN(n8931)
         );
  NAND2_X1 U10319 ( .A1(n9224), .A2(n8922), .ZN(n8923) );
  AOI21_X1 U10320 ( .B1(n8925), .B2(n8924), .A(n8923), .ZN(n8926) );
  OAI211_X1 U10321 ( .C1(n8927), .C2(n8926), .A(n8949), .B(n8960), .ZN(n8928)
         );
  NOR2_X1 U10322 ( .A1(n8929), .A2(n8928), .ZN(n8930) );
  NOR2_X1 U10323 ( .A1(n8931), .A2(n8930), .ZN(n8934) );
  MUX2_X1 U10324 ( .A(n9175), .B(n8932), .S(n8949), .Z(n8933) );
  NAND3_X1 U10325 ( .A1(n9156), .A2(n8934), .A3(n8933), .ZN(n8935) );
  NAND3_X1 U10326 ( .A1(n4825), .A2(n8936), .A3(n8935), .ZN(n8937) );
  NAND3_X1 U10327 ( .A1(n6338), .A2(n8938), .A3(n8937), .ZN(n8941) );
  MUX2_X1 U10328 ( .A(n9132), .B(n8939), .S(n8949), .Z(n8940) );
  AND2_X1 U10329 ( .A1(n8941), .A2(n8940), .ZN(n8945) );
  NAND2_X1 U10330 ( .A1(n9038), .A2(n8949), .ZN(n8943) );
  NAND3_X1 U10331 ( .A1(n9019), .A2(n8945), .A3(n9127), .ZN(n8948) );
  INV_X1 U10332 ( .A(n8946), .ZN(n8947) );
  AOI21_X1 U10333 ( .B1(n8948), .B2(n9013), .A(n8947), .ZN(n8950) );
  MUX2_X1 U10334 ( .A(n8951), .B(n8950), .S(n8949), .Z(n8952) );
  INV_X1 U10335 ( .A(n9017), .ZN(n9001) );
  INV_X1 U10336 ( .A(n9173), .ZN(n9179) );
  NAND2_X1 U10337 ( .A1(n8959), .A2(n8958), .ZN(n9211) );
  NAND2_X1 U10338 ( .A1(n8961), .A2(n8960), .ZN(n9225) );
  INV_X1 U10339 ( .A(n9310), .ZN(n9313) );
  INV_X1 U10340 ( .A(n8964), .ZN(n8989) );
  INV_X1 U10341 ( .A(n8965), .ZN(n8987) );
  OR2_X1 U10342 ( .A1(n9705), .A2(n8967), .ZN(n9707) );
  INV_X1 U10343 ( .A(n9707), .ZN(n8969) );
  NAND3_X1 U10344 ( .A1(n8969), .A2(n4920), .A3(n8968), .ZN(n8980) );
  INV_X1 U10345 ( .A(n8970), .ZN(n8972) );
  NAND3_X1 U10346 ( .A1(n8972), .A2(n8977), .A3(n8971), .ZN(n8975) );
  NAND3_X1 U10347 ( .A1(n8975), .A2(n8974), .A3(n8973), .ZN(n9004) );
  INV_X1 U10348 ( .A(n8976), .ZN(n8979) );
  NAND2_X1 U10349 ( .A1(n8978), .A2(n8977), .ZN(n9003) );
  NOR4_X1 U10350 ( .A1(n8980), .A2(n9004), .A3(n8979), .A4(n9003), .ZN(n8984)
         );
  NAND4_X1 U10351 ( .A1(n8984), .A2(n8983), .A3(n8982), .A4(n8981), .ZN(n8985)
         );
  NOR4_X1 U10352 ( .A1(n8987), .A2(n8986), .A3(n6175), .A4(n8985), .ZN(n8988)
         );
  NAND4_X1 U10353 ( .A1(n8991), .A2(n8990), .A3(n8989), .A4(n8988), .ZN(n8992)
         );
  NOR4_X1 U10354 ( .A1(n9297), .A2(n9313), .A3(n8993), .A4(n8992), .ZN(n8994)
         );
  NAND4_X1 U10355 ( .A1(n9244), .A2(n9257), .A3(n9276), .A4(n8994), .ZN(n8995)
         );
  NOR3_X1 U10356 ( .A1(n9211), .A2(n9225), .A3(n8995), .ZN(n8996) );
  NAND4_X1 U10357 ( .A1(n9156), .A2(n9179), .A3(n9194), .A4(n8996), .ZN(n8997)
         );
  NOR4_X1 U10358 ( .A1(n8999), .A2(n9147), .A3(n8998), .A4(n8997), .ZN(n9000)
         );
  XNOR2_X1 U10359 ( .A(n9127), .B(n9038), .ZN(n9134) );
  NAND4_X1 U10360 ( .A1(n9001), .A2(n4428), .A3(n9000), .A4(n9134), .ZN(n9002)
         );
  XNOR2_X1 U10361 ( .A(n9002), .B(n9704), .ZN(n9023) );
  INV_X1 U10362 ( .A(n9003), .ZN(n9005) );
  AOI21_X1 U10363 ( .B1(n9006), .B2(n9005), .A(n9004), .ZN(n9008) );
  AOI21_X1 U10364 ( .B1(n9009), .B2(n9008), .A(n9007), .ZN(n9012) );
  OAI211_X1 U10365 ( .C1(n9012), .C2(n9011), .A(n9010), .B(n4823), .ZN(n9015)
         );
  OAI211_X1 U10366 ( .C1(n9016), .C2(n9015), .A(n9014), .B(n9013), .ZN(n9018)
         );
  AOI21_X1 U10367 ( .B1(n9019), .B2(n9018), .A(n9017), .ZN(n9020) );
  NOR2_X1 U10368 ( .A1(n9020), .A2(n9704), .ZN(n9022) );
  MUX2_X1 U10369 ( .A(n9023), .B(n9022), .S(n9021), .Z(n9024) );
  INV_X1 U10370 ( .A(n9027), .ZN(n9029) );
  OAI21_X1 U10371 ( .B1(n9029), .B2(n9028), .A(n9030), .ZN(n9036) );
  INV_X1 U10372 ( .A(n9030), .ZN(n9033) );
  INV_X1 U10373 ( .A(n9047), .ZN(n9558) );
  NAND3_X1 U10374 ( .A1(n9031), .A2(n9719), .A3(n9558), .ZN(n9032) );
  OAI211_X1 U10375 ( .C1(n9034), .C2(n9033), .A(n9032), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9035) );
  OAI21_X1 U10376 ( .B1(n9037), .B2(n9036), .A(n9035), .ZN(P1_U3240) );
  MUX2_X1 U10377 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9038), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10378 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9039), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10379 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9160), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10380 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9180), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10381 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9161), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10382 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9388), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10383 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9228), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10384 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9389), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10385 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9260), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10386 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9412), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10387 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9295), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10388 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9411), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10389 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9541), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10390 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9431), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10391 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9540), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10392 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9432), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10393 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9040), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10394 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9041), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10395 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9042), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10396 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9043), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10397 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9792), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10398 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9778), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10399 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9793), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10400 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9779), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10401 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9768), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10402 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9044), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10403 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9748), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10404 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n6589), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10405 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6576), .S(P1_U4006), .Z(
        P1_U3556) );
  AOI21_X1 U10406 ( .B1(n9558), .B2(n9045), .A(n6372), .ZN(n9557) );
  INV_X1 U10407 ( .A(n9046), .ZN(n9048) );
  MUX2_X1 U10408 ( .A(n9570), .B(n9048), .S(n9047), .Z(n9050) );
  NAND2_X1 U10409 ( .A1(n9050), .A2(n9049), .ZN(n9051) );
  OAI211_X1 U10410 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9557), .A(n9051), .B(
        P1_U4006), .ZN(n9584) );
  XNOR2_X1 U10411 ( .A(n9053), .B(n9052), .ZN(n9058) );
  AOI21_X1 U10412 ( .B1(n9056), .B2(n9055), .A(n9054), .ZN(n9057) );
  AOI22_X1 U10413 ( .A1(n9687), .A2(n9058), .B1(n9686), .B2(n9057), .ZN(n9063)
         );
  AOI22_X1 U10414 ( .A1(n9678), .A2(n9060), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        P1_U3084), .ZN(n9062) );
  NAND2_X1 U10415 ( .A1(n9649), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n9061) );
  NAND4_X1 U10416 ( .A1(n9584), .A2(n9063), .A3(n9062), .A4(n9061), .ZN(
        P1_U3243) );
  INV_X1 U10417 ( .A(n9082), .ZN(n9066) );
  NAND2_X1 U10418 ( .A1(n9649), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9065) );
  NAND2_X1 U10419 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n9064) );
  OAI211_X1 U10420 ( .C1(n9634), .C2(n9066), .A(n9065), .B(n9064), .ZN(n9076)
         );
  AOI21_X1 U10421 ( .B1(n9071), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9067), .ZN(
        n9069) );
  XNOR2_X1 U10422 ( .A(n9082), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9068) );
  NOR2_X1 U10423 ( .A1(n9069), .A2(n9068), .ZN(n9078) );
  AOI211_X1 U10424 ( .C1(n9069), .C2(n9068), .A(n9078), .B(n9651), .ZN(n9075)
         );
  XNOR2_X1 U10425 ( .A(n9082), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n9072) );
  NOR2_X1 U10426 ( .A1(n9073), .A2(n9072), .ZN(n9081) );
  AOI211_X1 U10427 ( .C1(n9073), .C2(n9072), .A(n9081), .B(n9600), .ZN(n9074)
         );
  OR3_X1 U10428 ( .A1(n9076), .A2(n9075), .A3(n9074), .ZN(P1_U3258) );
  INV_X1 U10429 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9077) );
  XNOR2_X1 U10430 ( .A(n9093), .B(n9077), .ZN(n9080) );
  AOI21_X1 U10431 ( .B1(n9082), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9078), .ZN(
        n9079) );
  NAND2_X1 U10432 ( .A1(n9080), .A2(n9079), .ZN(n9095) );
  OAI21_X1 U10433 ( .B1(n9080), .B2(n9079), .A(n9095), .ZN(n9088) );
  AOI21_X1 U10434 ( .B1(n9082), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9081), .ZN(
        n9086) );
  NAND2_X1 U10435 ( .A1(n9093), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9097) );
  OR2_X1 U10436 ( .A1(n9093), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9083) );
  NAND2_X1 U10437 ( .A1(n9097), .A2(n9083), .ZN(n9085) );
  INV_X1 U10438 ( .A(n9098), .ZN(n9084) );
  AOI211_X1 U10439 ( .C1(n9086), .C2(n9085), .A(n9084), .B(n9600), .ZN(n9087)
         );
  AOI21_X1 U10440 ( .B1(n9686), .B2(n9088), .A(n9087), .ZN(n9092) );
  NAND2_X1 U10441 ( .A1(n9649), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n9090) );
  NAND2_X1 U10442 ( .A1(n9678), .A2(n9093), .ZN(n9089) );
  NAND4_X1 U10443 ( .A1(n9092), .A2(n9091), .A3(n9090), .A4(n9089), .ZN(
        P1_U3259) );
  OR2_X1 U10444 ( .A1(n9093), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U10445 ( .A1(n9095), .A2(n9094), .ZN(n9096) );
  XNOR2_X1 U10446 ( .A(n9096), .B(n9418), .ZN(n9104) );
  NAND2_X1 U10447 ( .A1(n9686), .A2(n9104), .ZN(n9102) );
  NAND2_X1 U10448 ( .A1(n9098), .A2(n9097), .ZN(n9099) );
  XNOR2_X1 U10449 ( .A(n9099), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9103) );
  NAND2_X1 U10450 ( .A1(n9103), .A2(n9100), .ZN(n9101) );
  NAND3_X1 U10451 ( .A1(n9102), .A2(n9634), .A3(n9101), .ZN(n9106) );
  OAI22_X1 U10452 ( .A1(n9651), .A2(n9104), .B1(n9103), .B2(n9600), .ZN(n9105)
         );
  INV_X1 U10453 ( .A(n9107), .ZN(n9109) );
  OAI211_X1 U10454 ( .C1(n4912), .C2(n9691), .A(n9109), .B(n9108), .ZN(
        P1_U3260) );
  XNOR2_X1 U10455 ( .A(n9116), .B(n9110), .ZN(n9111) );
  NAND2_X1 U10456 ( .A1(n9111), .A2(n9695), .ZN(n9352) );
  NAND2_X1 U10457 ( .A1(n9558), .A2(P1_B_REG_SCAN_IN), .ZN(n9112) );
  NAND2_X1 U10458 ( .A1(n9791), .A2(n9112), .ZN(n9136) );
  OR2_X1 U10459 ( .A1(n9113), .A2(n9136), .ZN(n9355) );
  NOR2_X1 U10460 ( .A1(n9241), .A2(n9355), .ZN(n9118) );
  NOR2_X1 U10461 ( .A1(n9443), .A2(n9326), .ZN(n9114) );
  AOI211_X1 U10462 ( .C1(n9208), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9118), .B(
        n9114), .ZN(n9115) );
  OAI21_X1 U10463 ( .B1(n9352), .B2(n9344), .A(n9115), .ZN(P1_U3261) );
  AOI211_X1 U10464 ( .C1(n9117), .C2(n4703), .A(n9319), .B(n9116), .ZN(n9357)
         );
  NAND2_X1 U10465 ( .A1(n9357), .A2(n9321), .ZN(n9120) );
  AOI21_X1 U10466 ( .B1(n9208), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9118), .ZN(
        n9119) );
  OAI211_X1 U10467 ( .C1(n9447), .C2(n9326), .A(n9120), .B(n9119), .ZN(
        P1_U3262) );
  NAND2_X1 U10468 ( .A1(n8006), .A2(n9039), .ZN(n9121) );
  NAND2_X1 U10469 ( .A1(n9122), .A2(n9121), .ZN(n9123) );
  INV_X1 U10470 ( .A(n9360), .ZN(n9140) );
  INV_X1 U10471 ( .A(n9124), .ZN(n9126) );
  AOI211_X1 U10472 ( .C1(n9127), .C2(n9126), .A(n9319), .B(n9125), .ZN(n9365)
         );
  NOR2_X1 U10473 ( .A1(n9363), .A2(n9326), .ZN(n9131) );
  AOI22_X1 U10474 ( .A1(n9208), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9128), .B2(
        n9701), .ZN(n9129) );
  OAI21_X1 U10475 ( .B1(n9362), .B2(n9338), .A(n9129), .ZN(n9130) );
  AOI211_X1 U10476 ( .C1(n9365), .C2(n9321), .A(n9131), .B(n9130), .ZN(n9139)
         );
  INV_X1 U10477 ( .A(n9134), .ZN(n9135) );
  NAND2_X1 U10478 ( .A1(n9366), .A2(n9716), .ZN(n9138) );
  OAI211_X1 U10479 ( .C1(n9140), .C2(n9333), .A(n9139), .B(n9138), .ZN(
        P1_U3355) );
  XOR2_X1 U10480 ( .A(n9147), .B(n9141), .Z(n9373) );
  INV_X1 U10481 ( .A(n9142), .ZN(n9143) );
  AOI211_X1 U10482 ( .C1(n9370), .C2(n9164), .A(n9319), .B(n9143), .ZN(n9369)
         );
  AOI22_X1 U10483 ( .A1(n9208), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9144), .B2(
        n9701), .ZN(n9145) );
  OAI21_X1 U10484 ( .B1(n4705), .B2(n9326), .A(n9145), .ZN(n9152) );
  AOI211_X1 U10485 ( .C1(n9147), .C2(n9146), .A(n9784), .B(n4440), .ZN(n9150)
         );
  OAI22_X1 U10486 ( .A1(n9148), .A2(n9361), .B1(n9362), .B2(n9733), .ZN(n9149)
         );
  NOR2_X1 U10487 ( .A1(n9150), .A2(n9149), .ZN(n9372) );
  NOR2_X1 U10488 ( .A1(n9372), .A2(n9241), .ZN(n9151) );
  AOI211_X1 U10489 ( .C1(n9321), .C2(n9369), .A(n9152), .B(n9151), .ZN(n9153)
         );
  OAI21_X1 U10490 ( .B1(n9373), .B2(n9333), .A(n9153), .ZN(P1_U3264) );
  XNOR2_X1 U10491 ( .A(n9154), .B(n9156), .ZN(n9376) );
  INV_X1 U10492 ( .A(n9376), .ZN(n9172) );
  INV_X1 U10493 ( .A(n9175), .ZN(n9155) );
  INV_X1 U10494 ( .A(n9156), .ZN(n9157) );
  XNOR2_X1 U10495 ( .A(n9158), .B(n9157), .ZN(n9159) );
  NAND2_X1 U10496 ( .A1(n9159), .A2(n9706), .ZN(n9163) );
  AOI22_X1 U10497 ( .A1(n9794), .A2(n9161), .B1(n9160), .B2(n9791), .ZN(n9162)
         );
  NAND2_X1 U10498 ( .A1(n9163), .A2(n9162), .ZN(n9374) );
  INV_X1 U10499 ( .A(n9164), .ZN(n9165) );
  AOI211_X1 U10500 ( .C1(n9166), .C2(n9183), .A(n9319), .B(n9165), .ZN(n9375)
         );
  NAND2_X1 U10501 ( .A1(n9375), .A2(n9321), .ZN(n9169) );
  AOI22_X1 U10502 ( .A1(n9208), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9167), .B2(
        n9701), .ZN(n9168) );
  OAI211_X1 U10503 ( .C1(n9452), .C2(n9326), .A(n9169), .B(n9168), .ZN(n9170)
         );
  AOI21_X1 U10504 ( .B1(n9374), .B2(n9716), .A(n9170), .ZN(n9171) );
  OAI21_X1 U10505 ( .B1(n9172), .B2(n9333), .A(n9171), .ZN(P1_U3265) );
  XNOR2_X1 U10506 ( .A(n9174), .B(n9173), .ZN(n9380) );
  INV_X1 U10507 ( .A(n9380), .ZN(n9191) );
  NAND2_X1 U10508 ( .A1(n9176), .A2(n9175), .ZN(n9177) );
  OAI211_X1 U10509 ( .C1(n9179), .C2(n9178), .A(n9177), .B(n9706), .ZN(n9182)
         );
  AOI22_X1 U10510 ( .A1(n9794), .A2(n9388), .B1(n9180), .B2(n9791), .ZN(n9181)
         );
  NAND2_X1 U10511 ( .A1(n9182), .A2(n9181), .ZN(n9378) );
  INV_X1 U10512 ( .A(n9183), .ZN(n9184) );
  AOI211_X1 U10513 ( .C1(n9185), .C2(n4696), .A(n9319), .B(n9184), .ZN(n9379)
         );
  NAND2_X1 U10514 ( .A1(n9379), .A2(n9321), .ZN(n9188) );
  AOI22_X1 U10515 ( .A1(n9241), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9186), .B2(
        n9701), .ZN(n9187) );
  OAI211_X1 U10516 ( .C1(n9456), .C2(n9326), .A(n9188), .B(n9187), .ZN(n9189)
         );
  AOI21_X1 U10517 ( .B1(n9378), .B2(n9716), .A(n9189), .ZN(n9190) );
  OAI21_X1 U10518 ( .B1(n9191), .B2(n9333), .A(n9190), .ZN(P1_U3266) );
  XOR2_X1 U10519 ( .A(n9194), .B(n9192), .Z(n9385) );
  INV_X1 U10520 ( .A(n9385), .ZN(n9206) );
  AOI22_X1 U10521 ( .A1(n9199), .A2(n9347), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9241), .ZN(n9205) );
  XOR2_X1 U10522 ( .A(n9194), .B(n9193), .Z(n9195) );
  OAI222_X1 U10523 ( .A1(n9733), .A2(n9197), .B1(n9361), .B2(n9196), .C1(n9195), .C2(n9784), .ZN(n9383) );
  AOI211_X1 U10524 ( .C1(n9199), .C2(n9213), .A(n9319), .B(n9198), .ZN(n9384)
         );
  INV_X1 U10525 ( .A(n9384), .ZN(n9202) );
  INV_X1 U10526 ( .A(n9200), .ZN(n9201) );
  OAI22_X1 U10527 ( .A1(n9202), .A2(n9704), .B1(n9301), .B2(n9201), .ZN(n9203)
         );
  OAI21_X1 U10528 ( .B1(n9383), .B2(n9203), .A(n9716), .ZN(n9204) );
  OAI211_X1 U10529 ( .C1(n9206), .C2(n9333), .A(n9205), .B(n9204), .ZN(
        P1_U3267) );
  XOR2_X1 U10530 ( .A(n9207), .B(n9211), .Z(n9394) );
  INV_X1 U10531 ( .A(n9394), .ZN(n9222) );
  AOI22_X1 U10532 ( .A1(n9335), .A2(n9388), .B1(n9208), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n9209) );
  OAI21_X1 U10533 ( .B1(n9247), .B2(n9338), .A(n9209), .ZN(n9219) );
  XOR2_X1 U10534 ( .A(n9211), .B(n9210), .Z(n9212) );
  NAND2_X1 U10535 ( .A1(n9212), .A2(n9706), .ZN(n9392) );
  OAI211_X1 U10536 ( .C1(n9464), .C2(n4467), .A(n9695), .B(n9213), .ZN(n9390)
         );
  INV_X1 U10537 ( .A(n9390), .ZN(n9216) );
  AOI22_X1 U10538 ( .A1(n9216), .A2(n9215), .B1(n9701), .B2(n9214), .ZN(n9217)
         );
  AOI21_X1 U10539 ( .B1(n9392), .B2(n9217), .A(n9241), .ZN(n9218) );
  AOI211_X1 U10540 ( .C1(n9347), .C2(n9220), .A(n9219), .B(n9218), .ZN(n9221)
         );
  OAI21_X1 U10541 ( .B1(n9222), .B2(n9333), .A(n9221), .ZN(P1_U3268) );
  XOR2_X1 U10542 ( .A(n9223), .B(n9225), .Z(n9398) );
  INV_X1 U10543 ( .A(n9398), .ZN(n9237) );
  NAND2_X1 U10544 ( .A1(n9242), .A2(n9224), .ZN(n9226) );
  XNOR2_X1 U10545 ( .A(n9226), .B(n9225), .ZN(n9227) );
  NAND2_X1 U10546 ( .A1(n9227), .A2(n9706), .ZN(n9230) );
  AOI22_X1 U10547 ( .A1(n9260), .A2(n9794), .B1(n9791), .B2(n9228), .ZN(n9229)
         );
  NAND2_X1 U10548 ( .A1(n9230), .A2(n9229), .ZN(n9396) );
  INV_X1 U10549 ( .A(n9248), .ZN(n9231) );
  AOI211_X1 U10550 ( .C1(n4695), .C2(n9231), .A(n9319), .B(n4467), .ZN(n9397)
         );
  NAND2_X1 U10551 ( .A1(n9397), .A2(n9321), .ZN(n9234) );
  AOI22_X1 U10552 ( .A1(n9241), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9232), .B2(
        n9701), .ZN(n9233) );
  OAI211_X1 U10553 ( .C1(n9467), .C2(n9326), .A(n9234), .B(n9233), .ZN(n9235)
         );
  AOI21_X1 U10554 ( .B1(n9396), .B2(n9716), .A(n9235), .ZN(n9236) );
  OAI21_X1 U10555 ( .B1(n9237), .B2(n9333), .A(n9236), .ZN(P1_U3269) );
  OAI21_X1 U10556 ( .B1(n9240), .B2(n9239), .A(n9238), .ZN(n9400) );
  AOI22_X1 U10557 ( .A1(n9249), .A2(n9347), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9241), .ZN(n9255) );
  OAI211_X1 U10558 ( .C1(n9244), .C2(n9243), .A(n9242), .B(n9706), .ZN(n9246)
         );
  NAND2_X1 U10559 ( .A1(n9412), .A2(n9794), .ZN(n9245) );
  OAI211_X1 U10560 ( .C1(n9247), .C2(n9733), .A(n9246), .B(n9245), .ZN(n9401)
         );
  AOI211_X1 U10561 ( .C1(n9249), .C2(n9263), .A(n9319), .B(n9248), .ZN(n9402)
         );
  INV_X1 U10562 ( .A(n9402), .ZN(n9252) );
  INV_X1 U10563 ( .A(n9250), .ZN(n9251) );
  OAI22_X1 U10564 ( .A1(n9252), .A2(n9704), .B1(n9301), .B2(n9251), .ZN(n9253)
         );
  OAI21_X1 U10565 ( .B1(n9401), .B2(n9253), .A(n9716), .ZN(n9254) );
  OAI211_X1 U10566 ( .C1(n9400), .C2(n9333), .A(n9255), .B(n9254), .ZN(
        P1_U3270) );
  XOR2_X1 U10567 ( .A(n9256), .B(n9257), .Z(n9408) );
  INV_X1 U10568 ( .A(n9408), .ZN(n9272) );
  XNOR2_X1 U10569 ( .A(n9258), .B(n9257), .ZN(n9259) );
  NAND2_X1 U10570 ( .A1(n9259), .A2(n9706), .ZN(n9262) );
  AOI22_X1 U10571 ( .A1(n9260), .A2(n9791), .B1(n9794), .B2(n9295), .ZN(n9261)
         );
  NAND2_X1 U10572 ( .A1(n9262), .A2(n9261), .ZN(n9406) );
  INV_X1 U10573 ( .A(n9263), .ZN(n9264) );
  AOI211_X1 U10574 ( .C1(n9265), .C2(n9285), .A(n9319), .B(n9264), .ZN(n9407)
         );
  NAND2_X1 U10575 ( .A1(n9407), .A2(n9321), .ZN(n9269) );
  INV_X1 U10576 ( .A(n9266), .ZN(n9267) );
  AOI22_X1 U10577 ( .A1(n9241), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9267), .B2(
        n9701), .ZN(n9268) );
  OAI211_X1 U10578 ( .C1(n9474), .C2(n9326), .A(n9269), .B(n9268), .ZN(n9270)
         );
  AOI21_X1 U10579 ( .B1(n9406), .B2(n9716), .A(n9270), .ZN(n9271) );
  OAI21_X1 U10580 ( .B1(n9272), .B2(n9333), .A(n9271), .ZN(P1_U3271) );
  OAI21_X1 U10581 ( .B1(n9274), .B2(n9276), .A(n9273), .ZN(n9275) );
  INV_X1 U10582 ( .A(n9275), .ZN(n9415) );
  XNOR2_X1 U10583 ( .A(n9277), .B(n9276), .ZN(n9417) );
  NAND2_X1 U10584 ( .A1(n9417), .A2(n9300), .ZN(n9291) );
  INV_X1 U10585 ( .A(n9338), .ZN(n9281) );
  INV_X1 U10586 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9279) );
  OAI22_X1 U10587 ( .A1(n9716), .A2(n9279), .B1(n9278), .B2(n9301), .ZN(n9280)
         );
  AOI21_X1 U10588 ( .B1(n9281), .B2(n9411), .A(n9280), .ZN(n9282) );
  OAI21_X1 U10589 ( .B1(n9284), .B2(n9283), .A(n9282), .ZN(n9288) );
  INV_X1 U10590 ( .A(n9304), .ZN(n9286) );
  OAI211_X1 U10591 ( .C1(n9286), .C2(n4702), .A(n9695), .B(n9285), .ZN(n9413)
         );
  NOR2_X1 U10592 ( .A1(n9413), .A2(n9344), .ZN(n9287) );
  AOI211_X1 U10593 ( .C1(n9347), .C2(n9289), .A(n9288), .B(n9287), .ZN(n9290)
         );
  OAI211_X1 U10594 ( .C1(n9415), .C2(n9350), .A(n9291), .B(n9290), .ZN(
        P1_U3272) );
  NAND2_X1 U10595 ( .A1(n9293), .A2(n9292), .ZN(n9294) );
  XNOR2_X1 U10596 ( .A(n9294), .B(n9297), .ZN(n9296) );
  AOI222_X1 U10597 ( .A1(n9706), .A2(n9296), .B1(n9295), .B2(n9791), .C1(n9541), .C2(n9794), .ZN(n9424) );
  OR2_X1 U10598 ( .A1(n9298), .A2(n9297), .ZN(n9420) );
  NAND3_X1 U10599 ( .A1(n9420), .A2(n9299), .A3(n9300), .ZN(n9309) );
  INV_X1 U10600 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9303) );
  OAI22_X1 U10601 ( .A1(n9716), .A2(n9303), .B1(n9302), .B2(n9301), .ZN(n9307)
         );
  OAI211_X1 U10602 ( .C1(n9318), .C2(n9305), .A(n9695), .B(n9304), .ZN(n9423)
         );
  NOR2_X1 U10603 ( .A1(n9423), .A2(n9344), .ZN(n9306) );
  AOI211_X1 U10604 ( .C1(n9347), .C2(n9421), .A(n9307), .B(n9306), .ZN(n9308)
         );
  OAI211_X1 U10605 ( .C1(n9241), .C2(n9424), .A(n9309), .B(n9308), .ZN(
        P1_U3273) );
  XNOR2_X1 U10606 ( .A(n9311), .B(n9310), .ZN(n9430) );
  NAND2_X1 U10607 ( .A1(n9330), .A2(n9312), .ZN(n9314) );
  XNOR2_X1 U10608 ( .A(n9314), .B(n9313), .ZN(n9315) );
  OAI222_X1 U10609 ( .A1(n9733), .A2(n9317), .B1(n9361), .B2(n9316), .C1(n9315), .C2(n9784), .ZN(n9426) );
  INV_X1 U10610 ( .A(n9342), .ZN(n9320) );
  AOI211_X1 U10611 ( .C1(n9428), .C2(n9320), .A(n9319), .B(n9318), .ZN(n9427)
         );
  NAND2_X1 U10612 ( .A1(n9427), .A2(n9321), .ZN(n9325) );
  INV_X1 U10613 ( .A(n9322), .ZN(n9323) );
  AOI22_X1 U10614 ( .A1(n9241), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9323), .B2(
        n9701), .ZN(n9324) );
  OAI211_X1 U10615 ( .C1(n9327), .C2(n9326), .A(n9325), .B(n9324), .ZN(n9328)
         );
  AOI21_X1 U10616 ( .B1(n9426), .B2(n9716), .A(n9328), .ZN(n9329) );
  OAI21_X1 U10617 ( .B1(n9430), .B2(n9333), .A(n9329), .ZN(P1_U3274) );
  OAI21_X1 U10618 ( .B1(n4471), .B2(n9331), .A(n9330), .ZN(n9548) );
  INV_X1 U10619 ( .A(n9548), .ZN(n9351) );
  AND2_X1 U10620 ( .A1(n9332), .A2(n9331), .ZN(n9544) );
  OR3_X1 U10621 ( .A1(n9545), .A2(n9544), .A3(n9333), .ZN(n9349) );
  AOI22_X1 U10622 ( .A1(n9241), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9334), .B2(
        n9701), .ZN(n9337) );
  NAND2_X1 U10623 ( .A1(n9335), .A2(n9541), .ZN(n9336) );
  OAI211_X1 U10624 ( .C1(n9339), .C2(n9338), .A(n9337), .B(n9336), .ZN(n9346)
         );
  NAND2_X1 U10625 ( .A1(n9340), .A2(n9539), .ZN(n9341) );
  NAND2_X1 U10626 ( .A1(n9341), .A2(n9695), .ZN(n9343) );
  OR2_X1 U10627 ( .A1(n9343), .A2(n9342), .ZN(n9543) );
  NOR2_X1 U10628 ( .A1(n9543), .A2(n9344), .ZN(n9345) );
  AOI211_X1 U10629 ( .C1(n9347), .C2(n9539), .A(n9346), .B(n9345), .ZN(n9348)
         );
  OAI211_X1 U10630 ( .C1(n9351), .C2(n9350), .A(n9349), .B(n9348), .ZN(
        P1_U3275) );
  INV_X1 U10631 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9353) );
  AND2_X1 U10632 ( .A1(n9352), .A2(n9355), .ZN(n9440) );
  MUX2_X1 U10633 ( .A(n9353), .B(n9440), .S(n10189), .Z(n9354) );
  OAI21_X1 U10634 ( .B1(n9443), .B2(n9439), .A(n9354), .ZN(P1_U3554) );
  INV_X1 U10635 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9358) );
  INV_X1 U10636 ( .A(n9355), .ZN(n9356) );
  NOR2_X1 U10637 ( .A1(n9357), .A2(n9356), .ZN(n9444) );
  MUX2_X1 U10638 ( .A(n9358), .B(n9444), .S(n10189), .Z(n9359) );
  OAI21_X1 U10639 ( .B1(n9447), .B2(n9439), .A(n9359), .ZN(P1_U3553) );
  NAND2_X1 U10640 ( .A1(n9360), .A2(n9789), .ZN(n9368) );
  OAI22_X1 U10641 ( .A1(n9363), .A2(n9782), .B1(n9362), .B2(n9361), .ZN(n9364)
         );
  NOR3_X1 U10642 ( .A1(n9366), .A2(n9365), .A3(n9364), .ZN(n9367) );
  NAND2_X1 U10643 ( .A1(n9368), .A2(n9367), .ZN(n9448) );
  MUX2_X1 U10644 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9448), .S(n10189), .Z(
        P1_U3552) );
  AOI21_X1 U10645 ( .B1(n9795), .B2(n9370), .A(n9369), .ZN(n9371) );
  OAI211_X1 U10646 ( .C1(n9373), .C2(n9759), .A(n9372), .B(n9371), .ZN(n9449)
         );
  MUX2_X1 U10647 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9449), .S(n10189), .Z(
        P1_U3550) );
  INV_X1 U10648 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10208) );
  AOI211_X1 U10649 ( .C1(n9376), .C2(n9789), .A(n9375), .B(n9374), .ZN(n9450)
         );
  MUX2_X1 U10650 ( .A(n10208), .B(n9450), .S(n10189), .Z(n9377) );
  OAI21_X1 U10651 ( .B1(n9452), .B2(n9439), .A(n9377), .ZN(P1_U3549) );
  INV_X1 U10652 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9381) );
  AOI211_X1 U10653 ( .C1(n9380), .C2(n9789), .A(n9379), .B(n9378), .ZN(n9453)
         );
  MUX2_X1 U10654 ( .A(n9381), .B(n9453), .S(n10189), .Z(n9382) );
  OAI21_X1 U10655 ( .B1(n9456), .B2(n9439), .A(n9382), .ZN(P1_U3548) );
  INV_X1 U10656 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9386) );
  AOI211_X1 U10657 ( .C1(n9385), .C2(n9789), .A(n9384), .B(n9383), .ZN(n9457)
         );
  MUX2_X1 U10658 ( .A(n9386), .B(n9457), .S(n10189), .Z(n9387) );
  OAI21_X1 U10659 ( .B1(n9460), .B2(n9439), .A(n9387), .ZN(P1_U3547) );
  INV_X1 U10660 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10197) );
  AOI22_X1 U10661 ( .A1(n9389), .A2(n9794), .B1(n9791), .B2(n9388), .ZN(n9391)
         );
  NAND3_X1 U10662 ( .A1(n9392), .A2(n9391), .A3(n9390), .ZN(n9393) );
  AOI21_X1 U10663 ( .B1(n9394), .B2(n9789), .A(n9393), .ZN(n9461) );
  MUX2_X1 U10664 ( .A(n10197), .B(n9461), .S(n10189), .Z(n9395) );
  OAI21_X1 U10665 ( .B1(n9464), .B2(n9439), .A(n9395), .ZN(P1_U3546) );
  INV_X1 U10666 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n10206) );
  AOI211_X1 U10667 ( .C1(n9398), .C2(n9789), .A(n9397), .B(n9396), .ZN(n9465)
         );
  MUX2_X1 U10668 ( .A(n10206), .B(n9465), .S(n10189), .Z(n9399) );
  OAI21_X1 U10669 ( .B1(n9467), .B2(n9439), .A(n9399), .ZN(P1_U3545) );
  INV_X1 U10670 ( .A(n9400), .ZN(n9403) );
  AOI211_X1 U10671 ( .C1(n9403), .C2(n9789), .A(n9402), .B(n9401), .ZN(n9468)
         );
  MUX2_X1 U10672 ( .A(n9404), .B(n9468), .S(n10189), .Z(n9405) );
  OAI21_X1 U10673 ( .B1(n9471), .B2(n9439), .A(n9405), .ZN(P1_U3544) );
  INV_X1 U10674 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9409) );
  AOI211_X1 U10675 ( .C1(n9408), .C2(n9789), .A(n9407), .B(n9406), .ZN(n9472)
         );
  MUX2_X1 U10676 ( .A(n9409), .B(n9472), .S(n10189), .Z(n9410) );
  OAI21_X1 U10677 ( .B1(n9474), .B2(n9439), .A(n9410), .ZN(P1_U3543) );
  AOI22_X1 U10678 ( .A1(n9412), .A2(n9791), .B1(n9794), .B2(n9411), .ZN(n9414)
         );
  OAI211_X1 U10679 ( .C1(n9415), .C2(n9784), .A(n9414), .B(n9413), .ZN(n9416)
         );
  AOI21_X1 U10680 ( .B1(n9417), .B2(n9789), .A(n9416), .ZN(n9475) );
  MUX2_X1 U10681 ( .A(n9418), .B(n9475), .S(n10189), .Z(n9419) );
  OAI21_X1 U10682 ( .B1(n4702), .B2(n9439), .A(n9419), .ZN(P1_U3542) );
  NAND3_X1 U10683 ( .A1(n9420), .A2(n9299), .A3(n9789), .ZN(n9425) );
  NAND2_X1 U10684 ( .A1(n9421), .A2(n9795), .ZN(n9422) );
  NAND4_X1 U10685 ( .A1(n9425), .A2(n9424), .A3(n9423), .A4(n9422), .ZN(n9478)
         );
  MUX2_X1 U10686 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9478), .S(n10189), .Z(
        P1_U3541) );
  AOI211_X1 U10687 ( .C1(n9795), .C2(n9428), .A(n9427), .B(n9426), .ZN(n9429)
         );
  OAI21_X1 U10688 ( .B1(n9430), .B2(n9759), .A(n9429), .ZN(n9479) );
  MUX2_X1 U10689 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9479), .S(n10189), .Z(
        P1_U3540) );
  AOI22_X1 U10690 ( .A1(n9794), .A2(n9432), .B1(n9431), .B2(n9791), .ZN(n9434)
         );
  NAND3_X1 U10691 ( .A1(n9435), .A2(n9434), .A3(n9433), .ZN(n9436) );
  AOI21_X1 U10692 ( .B1(n9437), .B2(n9789), .A(n9436), .ZN(n9480) );
  MUX2_X1 U10693 ( .A(n10203), .B(n9480), .S(n10189), .Z(n9438) );
  OAI21_X1 U10694 ( .B1(n9484), .B2(n9439), .A(n9438), .ZN(P1_U3538) );
  INV_X1 U10695 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9441) );
  MUX2_X1 U10696 ( .A(n9441), .B(n9440), .S(n9809), .Z(n9442) );
  OAI21_X1 U10697 ( .B1(n9443), .B2(n9483), .A(n9442), .ZN(P1_U3522) );
  INV_X1 U10698 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9445) );
  MUX2_X1 U10699 ( .A(n9445), .B(n9444), .S(n9809), .Z(n9446) );
  OAI21_X1 U10700 ( .B1(n9447), .B2(n9483), .A(n9446), .ZN(P1_U3521) );
  MUX2_X1 U10701 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9448), .S(n9809), .Z(
        P1_U3520) );
  MUX2_X1 U10702 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9449), .S(n9809), .Z(
        P1_U3518) );
  INV_X1 U10703 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10221) );
  MUX2_X1 U10704 ( .A(n10221), .B(n9450), .S(n9809), .Z(n9451) );
  OAI21_X1 U10705 ( .B1(n9452), .B2(n9483), .A(n9451), .ZN(P1_U3517) );
  INV_X1 U10706 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9454) );
  MUX2_X1 U10707 ( .A(n9454), .B(n9453), .S(n9809), .Z(n9455) );
  OAI21_X1 U10708 ( .B1(n9456), .B2(n9483), .A(n9455), .ZN(P1_U3516) );
  INV_X1 U10709 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9458) );
  MUX2_X1 U10710 ( .A(n9458), .B(n9457), .S(n9809), .Z(n9459) );
  OAI21_X1 U10711 ( .B1(n9460), .B2(n9483), .A(n9459), .ZN(P1_U3515) );
  INV_X1 U10712 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9462) );
  MUX2_X1 U10713 ( .A(n9462), .B(n9461), .S(n9809), .Z(n9463) );
  OAI21_X1 U10714 ( .B1(n9464), .B2(n9483), .A(n9463), .ZN(P1_U3514) );
  INV_X1 U10715 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10207) );
  MUX2_X1 U10716 ( .A(n10207), .B(n9465), .S(n9809), .Z(n9466) );
  OAI21_X1 U10717 ( .B1(n9467), .B2(n9483), .A(n9466), .ZN(P1_U3513) );
  INV_X1 U10718 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9469) );
  MUX2_X1 U10719 ( .A(n9469), .B(n9468), .S(n9809), .Z(n9470) );
  OAI21_X1 U10720 ( .B1(n9471), .B2(n9483), .A(n9470), .ZN(P1_U3512) );
  MUX2_X1 U10721 ( .A(n10136), .B(n9472), .S(n9809), .Z(n9473) );
  OAI21_X1 U10722 ( .B1(n9474), .B2(n9483), .A(n9473), .ZN(P1_U3511) );
  INV_X1 U10723 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9476) );
  MUX2_X1 U10724 ( .A(n9476), .B(n9475), .S(n9809), .Z(n9477) );
  OAI21_X1 U10725 ( .B1(n4702), .B2(n9483), .A(n9477), .ZN(P1_U3510) );
  MUX2_X1 U10726 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9478), .S(n9809), .Z(
        P1_U3508) );
  MUX2_X1 U10727 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9479), .S(n9809), .Z(
        P1_U3505) );
  INV_X1 U10728 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9481) );
  MUX2_X1 U10729 ( .A(n9481), .B(n9480), .S(n9809), .Z(n9482) );
  OAI21_X1 U10730 ( .B1(n9484), .B2(n9483), .A(n9482), .ZN(P1_U3499) );
  MUX2_X1 U10731 ( .A(n9486), .B(P1_D_REG_0__SCAN_IN), .S(n9485), .Z(P1_U3440)
         );
  AOI22_X1 U10732 ( .A1(n9487), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9488), .ZN(n9489) );
  OAI21_X1 U10733 ( .B1(n9490), .B2(n9494), .A(n9489), .ZN(P1_U3323) );
  OAI222_X1 U10734 ( .A1(n9494), .A2(n9493), .B1(n9492), .B2(P1_U3084), .C1(
        n10218), .C2(n9491), .ZN(P1_U3324) );
  MUX2_X1 U10735 ( .A(n9495), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI211_X1 U10736 ( .C1(n9498), .C2(n9497), .A(n9496), .B(n9651), .ZN(n9499)
         );
  AOI211_X1 U10737 ( .C1(n9678), .C2(n9501), .A(n9500), .B(n9499), .ZN(n9506)
         );
  OAI211_X1 U10738 ( .C1(n9504), .C2(n9503), .A(n9687), .B(n9502), .ZN(n9505)
         );
  OAI211_X1 U10739 ( .C1(n9507), .C2(n9691), .A(n9506), .B(n9505), .ZN(
        P1_U3244) );
  NOR2_X1 U10740 ( .A1(n9508), .A2(n9921), .ZN(n9509) );
  INV_X1 U10741 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9512) );
  AOI22_X1 U10742 ( .A1(n9945), .A2(n9532), .B1(n9512), .B2(n9943), .ZN(
        P2_U3550) );
  OAI22_X1 U10743 ( .A1(n9514), .A2(n9922), .B1(n9513), .B2(n9921), .ZN(n9516)
         );
  AOI211_X1 U10744 ( .C1(n9517), .C2(n9927), .A(n9516), .B(n9515), .ZN(n9534)
         );
  AOI22_X1 U10745 ( .A1(n9945), .A2(n9534), .B1(n10209), .B2(n9943), .ZN(
        P2_U3535) );
  OAI22_X1 U10746 ( .A1(n9519), .A2(n9922), .B1(n9518), .B2(n9921), .ZN(n9521)
         );
  AOI211_X1 U10747 ( .C1(n9522), .C2(n9927), .A(n9521), .B(n9520), .ZN(n9536)
         );
  AOI22_X1 U10748 ( .A1(n9945), .A2(n9536), .B1(n9523), .B2(n9943), .ZN(
        P2_U3534) );
  INV_X1 U10749 ( .A(n9524), .ZN(n9912) );
  INV_X1 U10750 ( .A(n9525), .ZN(n9526) );
  OAI22_X1 U10751 ( .A1(n9527), .A2(n9922), .B1(n9526), .B2(n9921), .ZN(n9529)
         );
  AOI211_X1 U10752 ( .C1(n9912), .C2(n9530), .A(n9529), .B(n9528), .ZN(n9538)
         );
  AOI22_X1 U10753 ( .A1(n9945), .A2(n9538), .B1(n10116), .B2(n9943), .ZN(
        P2_U3533) );
  INV_X1 U10754 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9531) );
  AOI22_X1 U10755 ( .A1(n9930), .A2(n9532), .B1(n9531), .B2(n9928), .ZN(
        P2_U3518) );
  INV_X1 U10756 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9533) );
  AOI22_X1 U10757 ( .A1(n9930), .A2(n9534), .B1(n9533), .B2(n9928), .ZN(
        P2_U3496) );
  INV_X1 U10758 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9535) );
  AOI22_X1 U10759 ( .A1(n9930), .A2(n9536), .B1(n9535), .B2(n9928), .ZN(
        P2_U3493) );
  INV_X1 U10760 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9537) );
  AOI22_X1 U10761 ( .A1(n9930), .A2(n9538), .B1(n9537), .B2(n9928), .ZN(
        P2_U3490) );
  AOI22_X1 U10762 ( .A1(n9541), .A2(n9791), .B1(n9540), .B2(n9794), .ZN(n9542)
         );
  OAI211_X1 U10763 ( .C1(n4698), .C2(n9782), .A(n9543), .B(n9542), .ZN(n9547)
         );
  NOR3_X1 U10764 ( .A1(n9545), .A2(n9544), .A3(n9759), .ZN(n9546) );
  AOI211_X1 U10765 ( .C1(n9706), .C2(n9548), .A(n9547), .B(n9546), .ZN(n9550)
         );
  AOI22_X1 U10766 ( .A1(n10189), .A2(n9550), .B1(n7197), .B2(n10187), .ZN(
        P1_U3539) );
  INV_X1 U10767 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9549) );
  AOI22_X1 U10768 ( .A1(n9809), .A2(n9550), .B1(n9549), .B2(n9807), .ZN(
        P1_U3502) );
  INV_X1 U10769 ( .A(n9551), .ZN(n9555) );
  AOI21_X1 U10770 ( .B1(n9795), .B2(n9553), .A(n9552), .ZN(n9554) );
  OAI211_X1 U10771 ( .C1(n9556), .C2(n9801), .A(n9555), .B(n9554), .ZN(n10188)
         );
  MUX2_X1 U10772 ( .A(n10188), .B(P1_REG0_REG_11__SCAN_IN), .S(n9807), .Z(
        P1_U3487) );
  XNOR2_X1 U10773 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XOR2_X1 U10774 ( .A(n4909), .B(P1_RD_REG_SCAN_IN), .Z(U126) );
  OAI21_X1 U10775 ( .B1(n9558), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9557), .ZN(
        n9559) );
  XNOR2_X1 U10776 ( .A(n9559), .B(P1_IR_REG_0__SCAN_IN), .ZN(n9560) );
  AOI22_X1 U10777 ( .A1(n9561), .A2(n9560), .B1(n9649), .B2(
        P1_ADDR_REG_0__SCAN_IN), .ZN(n9562) );
  OAI21_X1 U10778 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6699), .A(n9562), .ZN(
        P1_U3241) );
  INV_X1 U10779 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10096) );
  OAI22_X1 U10780 ( .A1(n9634), .A2(n6060), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10096), .ZN(n9567) );
  NAND2_X1 U10781 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9565) );
  AOI211_X1 U10782 ( .C1(n9565), .C2(n9564), .A(n9563), .B(n9651), .ZN(n9566)
         );
  AOI211_X1 U10783 ( .C1(P1_ADDR_REG_1__SCAN_IN), .C2(n9649), .A(n9567), .B(
        n9566), .ZN(n9572) );
  OAI211_X1 U10784 ( .C1(n9570), .C2(n9569), .A(n9687), .B(n9568), .ZN(n9571)
         );
  NAND2_X1 U10785 ( .A1(n9572), .A2(n9571), .ZN(P1_U3242) );
  XOR2_X1 U10786 ( .A(n9574), .B(n9573), .Z(n9576) );
  OAI22_X1 U10787 ( .A1(n9576), .A2(n9651), .B1(n9575), .B2(n9634), .ZN(n9583)
         );
  AOI21_X1 U10788 ( .B1(n9579), .B2(n9578), .A(n9577), .ZN(n9580) );
  NOR2_X1 U10789 ( .A1(n9600), .A2(n9580), .ZN(n9581) );
  NOR3_X1 U10790 ( .A1(n9583), .A2(n9582), .A3(n9581), .ZN(n9585) );
  OAI211_X1 U10791 ( .C1(n9586), .C2(n9691), .A(n9585), .B(n9584), .ZN(
        P1_U3245) );
  INV_X1 U10792 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9603) );
  AOI21_X1 U10793 ( .B1(n9589), .B2(n9588), .A(n9587), .ZN(n9590) );
  NAND2_X1 U10794 ( .A1(n9686), .A2(n9590), .ZN(n9593) );
  INV_X1 U10795 ( .A(n9591), .ZN(n9592) );
  OAI211_X1 U10796 ( .C1(n9594), .C2(n9634), .A(n9593), .B(n9592), .ZN(n9595)
         );
  INV_X1 U10797 ( .A(n9595), .ZN(n9602) );
  AOI21_X1 U10798 ( .B1(n9598), .B2(n9597), .A(n9596), .ZN(n9599) );
  OR2_X1 U10799 ( .A1(n9600), .A2(n9599), .ZN(n9601) );
  OAI211_X1 U10800 ( .C1(n9603), .C2(n9691), .A(n9602), .B(n9601), .ZN(
        P1_U3246) );
  INV_X1 U10801 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10150) );
  OAI21_X1 U10802 ( .B1(n9606), .B2(n9605), .A(n9604), .ZN(n9607) );
  NAND2_X1 U10803 ( .A1(n9686), .A2(n9607), .ZN(n9610) );
  INV_X1 U10804 ( .A(n9608), .ZN(n9609) );
  OAI211_X1 U10805 ( .C1(n9611), .C2(n9634), .A(n9610), .B(n9609), .ZN(n9612)
         );
  INV_X1 U10806 ( .A(n9612), .ZN(n9617) );
  OAI211_X1 U10807 ( .C1(n9615), .C2(n9614), .A(n9687), .B(n9613), .ZN(n9616)
         );
  OAI211_X1 U10808 ( .C1(n9691), .C2(n10150), .A(n9617), .B(n9616), .ZN(
        P1_U3247) );
  OAI21_X1 U10809 ( .B1(n9620), .B2(n9619), .A(n9618), .ZN(n9624) );
  OAI21_X1 U10810 ( .B1(n9634), .B2(n9622), .A(n9621), .ZN(n9623) );
  AOI21_X1 U10811 ( .B1(n9624), .B2(n9686), .A(n9623), .ZN(n9629) );
  OAI211_X1 U10812 ( .C1(n9627), .C2(n9626), .A(n9625), .B(n9687), .ZN(n9628)
         );
  OAI211_X1 U10813 ( .C1(n9691), .C2(n10290), .A(n9629), .B(n9628), .ZN(
        P1_U3250) );
  INV_X1 U10814 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9643) );
  OAI21_X1 U10815 ( .B1(n9632), .B2(n9631), .A(n9630), .ZN(n9637) );
  NOR2_X1 U10816 ( .A1(n9634), .A2(n9633), .ZN(n9635) );
  AOI211_X1 U10817 ( .C1(n9637), .C2(n9686), .A(n9636), .B(n9635), .ZN(n9642)
         );
  OAI211_X1 U10818 ( .C1(n9640), .C2(n9639), .A(n9687), .B(n9638), .ZN(n9641)
         );
  OAI211_X1 U10819 ( .C1(n9643), .C2(n9691), .A(n9642), .B(n9641), .ZN(
        P1_U3251) );
  AOI21_X1 U10820 ( .B1(n9678), .B2(n9645), .A(n9644), .ZN(n9646) );
  OAI21_X1 U10821 ( .B1(n9647), .B2(n9651), .A(n9646), .ZN(n9648) );
  AOI21_X1 U10822 ( .B1(n9649), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n9648), .ZN(
        n9661) );
  OR3_X1 U10823 ( .A1(n9652), .A2(n9651), .A3(n9650), .ZN(n9660) );
  NAND2_X1 U10824 ( .A1(n9653), .A2(n10029), .ZN(n9655) );
  OAI211_X1 U10825 ( .C1(n9657), .C2(n9655), .A(n9654), .B(n9687), .ZN(n9659)
         );
  NAND3_X1 U10826 ( .A1(n9657), .A2(n9656), .A3(n9687), .ZN(n9658) );
  NAND4_X1 U10827 ( .A1(n9661), .A2(n9660), .A3(n9659), .A4(n9658), .ZN(
        P1_U3252) );
  INV_X1 U10828 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10238) );
  OAI211_X1 U10829 ( .C1(n9664), .C2(n9663), .A(n9687), .B(n9662), .ZN(n9665)
         );
  INV_X1 U10830 ( .A(n9665), .ZN(n9666) );
  AOI211_X1 U10831 ( .C1(n9668), .C2(n9678), .A(n9667), .B(n9666), .ZN(n9675)
         );
  MUX2_X1 U10832 ( .A(n7046), .B(P1_REG1_REG_13__SCAN_IN), .S(n9668), .Z(n9669) );
  INV_X1 U10833 ( .A(n9669), .ZN(n9672) );
  OAI21_X1 U10834 ( .B1(n9672), .B2(n9671), .A(n9670), .ZN(n9673) );
  NAND2_X1 U10835 ( .A1(n9686), .A2(n9673), .ZN(n9674) );
  OAI211_X1 U10836 ( .C1(n9691), .C2(n10238), .A(n9675), .B(n9674), .ZN(
        P1_U3254) );
  INV_X1 U10837 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10159) );
  AOI21_X1 U10838 ( .B1(n9678), .B2(n9677), .A(n9676), .ZN(n9690) );
  OAI21_X1 U10839 ( .B1(n9681), .B2(n9680), .A(n9679), .ZN(n9688) );
  OAI21_X1 U10840 ( .B1(n9684), .B2(n9683), .A(n9682), .ZN(n9685) );
  AOI22_X1 U10841 ( .A1(n9688), .A2(n9687), .B1(n9686), .B2(n9685), .ZN(n9689)
         );
  OAI211_X1 U10842 ( .C1(n10159), .C2(n9691), .A(n9690), .B(n9689), .ZN(
        P1_U3255) );
  OAI21_X1 U10843 ( .B1(n9705), .B2(n9693), .A(n9692), .ZN(n9713) );
  INV_X1 U10844 ( .A(n9713), .ZN(n9730) );
  NAND2_X1 U10845 ( .A1(n9700), .A2(n9694), .ZN(n9696) );
  NAND2_X1 U10846 ( .A1(n9696), .A2(n9695), .ZN(n9698) );
  OR2_X1 U10847 ( .A1(n9698), .A2(n9697), .ZN(n9726) );
  NAND2_X1 U10848 ( .A1(n9700), .A2(n9699), .ZN(n9703) );
  NAND2_X1 U10849 ( .A1(n9701), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n9702) );
  OAI211_X1 U10850 ( .C1(n9726), .C2(n9704), .A(n9703), .B(n9702), .ZN(n9714)
         );
  AOI22_X1 U10851 ( .A1(n9794), .A2(n6572), .B1(n6589), .B2(n9791), .ZN(n9711)
         );
  INV_X1 U10852 ( .A(n9705), .ZN(n9709) );
  OAI211_X1 U10853 ( .C1(n9709), .C2(n9708), .A(n9707), .B(n9706), .ZN(n9710)
         );
  OAI211_X1 U10854 ( .C1(n9713), .C2(n9712), .A(n9711), .B(n9710), .ZN(n9728)
         );
  AOI211_X1 U10855 ( .C1(n9715), .C2(n9730), .A(n9714), .B(n9728), .ZN(n9717)
         );
  AOI22_X1 U10856 ( .A1(n9241), .A2(n6469), .B1(n9717), .B2(n9716), .ZN(
        P1_U3290) );
  AND2_X1 U10857 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9721), .ZN(P1_U3292) );
  AND2_X1 U10858 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9721), .ZN(P1_U3293) );
  AND2_X1 U10859 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9721), .ZN(P1_U3294) );
  AND2_X1 U10860 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9721), .ZN(P1_U3295) );
  AND2_X1 U10861 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9721), .ZN(P1_U3296) );
  AND2_X1 U10862 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9721), .ZN(P1_U3297) );
  INV_X1 U10863 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10132) );
  NOR2_X1 U10864 ( .A1(n9720), .A2(n10132), .ZN(P1_U3298) );
  AND2_X1 U10865 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9721), .ZN(P1_U3299) );
  AND2_X1 U10866 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9721), .ZN(P1_U3300) );
  AND2_X1 U10867 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9721), .ZN(P1_U3301) );
  AND2_X1 U10868 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9721), .ZN(P1_U3302) );
  AND2_X1 U10869 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9721), .ZN(P1_U3303) );
  AND2_X1 U10870 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9721), .ZN(P1_U3304) );
  AND2_X1 U10871 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9721), .ZN(P1_U3305) );
  AND2_X1 U10872 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9721), .ZN(P1_U3306) );
  INV_X1 U10873 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10240) );
  NOR2_X1 U10874 ( .A1(n9720), .A2(n10240), .ZN(P1_U3307) );
  INV_X1 U10875 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10040) );
  NOR2_X1 U10876 ( .A1(n9720), .A2(n10040), .ZN(P1_U3308) );
  AND2_X1 U10877 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9721), .ZN(P1_U3309) );
  AND2_X1 U10878 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9721), .ZN(P1_U3310) );
  AND2_X1 U10879 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9721), .ZN(P1_U3311) );
  AND2_X1 U10880 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9721), .ZN(P1_U3312) );
  AND2_X1 U10881 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9721), .ZN(P1_U3313) );
  AND2_X1 U10882 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9721), .ZN(P1_U3314) );
  AND2_X1 U10883 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9721), .ZN(P1_U3315) );
  AND2_X1 U10884 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9721), .ZN(P1_U3316) );
  AND2_X1 U10885 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9721), .ZN(P1_U3317) );
  INV_X1 U10886 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10012) );
  NOR2_X1 U10887 ( .A1(n9720), .A2(n10012), .ZN(P1_U3318) );
  AND2_X1 U10888 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9721), .ZN(P1_U3319) );
  INV_X1 U10889 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10053) );
  NOR2_X1 U10890 ( .A1(n9720), .A2(n10053), .ZN(P1_U3320) );
  AND2_X1 U10891 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9721), .ZN(P1_U3321) );
  INV_X1 U10892 ( .A(n9722), .ZN(n9723) );
  NOR2_X1 U10893 ( .A1(n9724), .A2(n9723), .ZN(n9811) );
  AOI22_X1 U10894 ( .A1(n9809), .A2(n9811), .B1(n9725), .B2(n9807), .ZN(
        P1_U3454) );
  INV_X1 U10895 ( .A(n9801), .ZN(n9746) );
  OAI21_X1 U10896 ( .B1(n9727), .B2(n9782), .A(n9726), .ZN(n9729) );
  AOI211_X1 U10897 ( .C1(n9746), .C2(n9730), .A(n9729), .B(n9728), .ZN(n9812)
         );
  AOI22_X1 U10898 ( .A1(n9809), .A2(n9812), .B1(n6054), .B2(n9807), .ZN(
        P1_U3457) );
  OAI21_X1 U10899 ( .B1(n9746), .B2(n9805), .A(n9731), .ZN(n9739) );
  OAI22_X1 U10900 ( .A1(n9734), .A2(n9733), .B1(n9732), .B2(n9782), .ZN(n9736)
         );
  AOI211_X1 U10901 ( .C1(n9794), .C2(n6576), .A(n9736), .B(n9735), .ZN(n9738)
         );
  AND3_X1 U10902 ( .A1(n9739), .A2(n9738), .A3(n9737), .ZN(n9814) );
  INV_X1 U10903 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10251) );
  AOI22_X1 U10904 ( .A1(n9809), .A2(n9814), .B1(n10251), .B2(n9807), .ZN(
        P1_U3460) );
  INV_X1 U10905 ( .A(n9740), .ZN(n9741) );
  OAI21_X1 U10906 ( .B1(n9742), .B2(n9782), .A(n9741), .ZN(n9744) );
  AOI211_X1 U10907 ( .C1(n9746), .C2(n9745), .A(n9744), .B(n9743), .ZN(n9816)
         );
  INV_X1 U10908 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9747) );
  AOI22_X1 U10909 ( .A1(n9809), .A2(n9816), .B1(n9747), .B2(n9807), .ZN(
        P1_U3463) );
  INV_X1 U10910 ( .A(n9755), .ZN(n9757) );
  AOI22_X1 U10911 ( .A1(n9794), .A2(n9748), .B1(n9768), .B2(n9791), .ZN(n9749)
         );
  OAI211_X1 U10912 ( .C1(n9751), .C2(n9782), .A(n9750), .B(n9749), .ZN(n9752)
         );
  NOR2_X1 U10913 ( .A1(n9753), .A2(n9752), .ZN(n9754) );
  OAI21_X1 U10914 ( .B1(n9755), .B2(n9801), .A(n9754), .ZN(n9756) );
  AOI21_X1 U10915 ( .B1(n9805), .B2(n9757), .A(n9756), .ZN(n9818) );
  INV_X1 U10916 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9758) );
  AOI22_X1 U10917 ( .A1(n9809), .A2(n9818), .B1(n9758), .B2(n9807), .ZN(
        P1_U3466) );
  NOR2_X1 U10918 ( .A1(n9760), .A2(n9759), .ZN(n9766) );
  OAI211_X1 U10919 ( .C1(n9763), .C2(n9782), .A(n9762), .B(n9761), .ZN(n9764)
         );
  AOI21_X1 U10920 ( .B1(n9766), .B2(n9765), .A(n9764), .ZN(n9819) );
  INV_X1 U10921 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9767) );
  AOI22_X1 U10922 ( .A1(n9809), .A2(n9819), .B1(n9767), .B2(n9807), .ZN(
        P1_U3469) );
  AOI22_X1 U10923 ( .A1(n9794), .A2(n9768), .B1(n9793), .B2(n9791), .ZN(n9772)
         );
  NAND2_X1 U10924 ( .A1(n9795), .A2(n9769), .ZN(n9770) );
  NAND4_X1 U10925 ( .A1(n9773), .A2(n9772), .A3(n9771), .A4(n9770), .ZN(n9776)
         );
  NOR2_X1 U10926 ( .A1(n9774), .A2(n9801), .ZN(n9775) );
  AOI211_X1 U10927 ( .C1(n9805), .C2(n9777), .A(n9776), .B(n9775), .ZN(n9821)
         );
  INV_X1 U10928 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10095) );
  AOI22_X1 U10929 ( .A1(n9809), .A2(n9821), .B1(n10095), .B2(n9807), .ZN(
        P1_U3472) );
  AOI22_X1 U10930 ( .A1(n9794), .A2(n9779), .B1(n9778), .B2(n9791), .ZN(n9780)
         );
  OAI211_X1 U10931 ( .C1(n9783), .C2(n9782), .A(n9781), .B(n9780), .ZN(n9787)
         );
  NOR2_X1 U10932 ( .A1(n9785), .A2(n9784), .ZN(n9786) );
  AOI211_X1 U10933 ( .C1(n9789), .C2(n9788), .A(n9787), .B(n9786), .ZN(n9823)
         );
  INV_X1 U10934 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9790) );
  AOI22_X1 U10935 ( .A1(n9809), .A2(n9823), .B1(n9790), .B2(n9807), .ZN(
        P1_U3475) );
  AOI22_X1 U10936 ( .A1(n9794), .A2(n9793), .B1(n9792), .B2(n9791), .ZN(n9799)
         );
  NAND2_X1 U10937 ( .A1(n9796), .A2(n9795), .ZN(n9797) );
  NAND4_X1 U10938 ( .A1(n9800), .A2(n9799), .A3(n9798), .A4(n9797), .ZN(n9804)
         );
  INV_X1 U10939 ( .A(n9806), .ZN(n9802) );
  NOR2_X1 U10940 ( .A1(n9802), .A2(n9801), .ZN(n9803) );
  AOI211_X1 U10941 ( .C1(n9806), .C2(n9805), .A(n9804), .B(n9803), .ZN(n9825)
         );
  INV_X1 U10942 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9808) );
  AOI22_X1 U10943 ( .A1(n9809), .A2(n9825), .B1(n9808), .B2(n9807), .ZN(
        P1_U3478) );
  AOI22_X1 U10944 ( .A1(n10189), .A2(n9811), .B1(n9810), .B2(n10187), .ZN(
        P1_U3523) );
  AOI22_X1 U10945 ( .A1(n10189), .A2(n9812), .B1(n6488), .B2(n10187), .ZN(
        P1_U3524) );
  INV_X1 U10946 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9813) );
  AOI22_X1 U10947 ( .A1(n10189), .A2(n9814), .B1(n9813), .B2(n10187), .ZN(
        P1_U3525) );
  INV_X1 U10948 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9815) );
  AOI22_X1 U10949 ( .A1(n10189), .A2(n9816), .B1(n9815), .B2(n10187), .ZN(
        P1_U3526) );
  INV_X1 U10950 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9817) );
  AOI22_X1 U10951 ( .A1(n10189), .A2(n9818), .B1(n9817), .B2(n10187), .ZN(
        P1_U3527) );
  AOI22_X1 U10952 ( .A1(n10189), .A2(n9819), .B1(n6485), .B2(n10187), .ZN(
        P1_U3528) );
  INV_X1 U10953 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9820) );
  AOI22_X1 U10954 ( .A1(n10189), .A2(n9821), .B1(n9820), .B2(n10187), .ZN(
        P1_U3529) );
  INV_X1 U10955 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9822) );
  AOI22_X1 U10956 ( .A1(n10189), .A2(n9823), .B1(n9822), .B2(n10187), .ZN(
        P1_U3530) );
  AOI22_X1 U10957 ( .A1(n10189), .A2(n9825), .B1(n9824), .B2(n10187), .ZN(
        P1_U3531) );
  AOI21_X1 U10958 ( .B1(n9828), .B2(n9827), .A(n9826), .ZN(n9837) );
  OAI22_X1 U10959 ( .A1(n9829), .A2(n9907), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10205), .ZN(n9835) );
  OAI22_X1 U10960 ( .A1(n9833), .A2(n9832), .B1(n9831), .B2(n9830), .ZN(n9834)
         );
  AOI211_X1 U10961 ( .C1(n9837), .C2(n9836), .A(n9835), .B(n9834), .ZN(n9838)
         );
  OAI21_X1 U10962 ( .B1(n9840), .B2(n9839), .A(n9838), .ZN(P2_U3219) );
  XNOR2_X1 U10963 ( .A(n9841), .B(n9849), .ZN(n9844) );
  AOI21_X1 U10964 ( .B1(n9844), .B2(n9843), .A(n9842), .ZN(n9915) );
  AOI222_X1 U10965 ( .A1(n9848), .A2(n9847), .B1(n9846), .B2(n9845), .C1(
        P2_REG2_REG_11__SCAN_IN), .C2(n9860), .ZN(n9859) );
  OR2_X1 U10966 ( .A1(n9850), .A2(n9849), .ZN(n9851) );
  AND2_X1 U10967 ( .A1(n9852), .A2(n9851), .ZN(n9918) );
  OAI211_X1 U10968 ( .C1(n9854), .C2(n9916), .A(n9853), .B(n4481), .ZN(n9914)
         );
  NOR2_X1 U10969 ( .A1(n9914), .A2(n9855), .ZN(n9856) );
  AOI21_X1 U10970 ( .B1(n9918), .B2(n9857), .A(n9856), .ZN(n9858) );
  OAI211_X1 U10971 ( .C1(n9860), .C2(n9915), .A(n9859), .B(n9858), .ZN(
        P2_U3285) );
  AND2_X1 U10972 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9865), .ZN(P2_U3297) );
  AND2_X1 U10973 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9865), .ZN(P2_U3298) );
  AND2_X1 U10974 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9865), .ZN(P2_U3299) );
  INV_X1 U10975 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n9975) );
  NOR2_X1 U10976 ( .A1(n9863), .A2(n9975), .ZN(P2_U3300) );
  AND2_X1 U10977 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9865), .ZN(P2_U3301) );
  AND2_X1 U10978 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9865), .ZN(P2_U3302) );
  INV_X1 U10979 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n10052) );
  NOR2_X1 U10980 ( .A1(n9863), .A2(n10052), .ZN(P2_U3303) );
  AND2_X1 U10981 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9865), .ZN(P2_U3304) );
  AND2_X1 U10982 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9865), .ZN(P2_U3305) );
  AND2_X1 U10983 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9865), .ZN(P2_U3306) );
  INV_X1 U10984 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n9988) );
  NOR2_X1 U10985 ( .A1(n9863), .A2(n9988), .ZN(P2_U3307) );
  AND2_X1 U10986 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9865), .ZN(P2_U3308) );
  AND2_X1 U10987 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9865), .ZN(P2_U3309) );
  AND2_X1 U10988 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9865), .ZN(P2_U3310) );
  AND2_X1 U10989 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9865), .ZN(P2_U3311) );
  AND2_X1 U10990 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9865), .ZN(P2_U3312) );
  INV_X1 U10991 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10064) );
  NOR2_X1 U10992 ( .A1(n9863), .A2(n10064), .ZN(P2_U3313) );
  AND2_X1 U10993 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9865), .ZN(P2_U3314) );
  AND2_X1 U10994 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9865), .ZN(P2_U3315) );
  INV_X1 U10995 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10133) );
  NOR2_X1 U10996 ( .A1(n9863), .A2(n10133), .ZN(P2_U3316) );
  AND2_X1 U10997 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9865), .ZN(P2_U3317) );
  AND2_X1 U10998 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9865), .ZN(P2_U3318) );
  INV_X1 U10999 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10106) );
  NOR2_X1 U11000 ( .A1(n9863), .A2(n10106), .ZN(P2_U3319) );
  AND2_X1 U11001 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9865), .ZN(P2_U3320) );
  AND2_X1 U11002 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9865), .ZN(P2_U3321) );
  AND2_X1 U11003 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9865), .ZN(P2_U3322) );
  INV_X1 U11004 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10145) );
  NOR2_X1 U11005 ( .A1(n9863), .A2(n10145), .ZN(P2_U3323) );
  AND2_X1 U11006 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9865), .ZN(P2_U3324) );
  AND2_X1 U11007 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9865), .ZN(P2_U3325) );
  AND2_X1 U11008 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9865), .ZN(P2_U3326) );
  INV_X1 U11009 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10161) );
  AOI22_X1 U11010 ( .A1(n9868), .A2(n9864), .B1(n10161), .B2(n9865), .ZN(
        P2_U3437) );
  INV_X1 U11011 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9866) );
  AOI22_X1 U11012 ( .A1(n9868), .A2(n9867), .B1(n9866), .B2(n9865), .ZN(
        P2_U3438) );
  OAI21_X1 U11013 ( .B1(n9871), .B2(n9870), .A(n9869), .ZN(n9872) );
  AOI21_X1 U11014 ( .B1(n9927), .B2(n9873), .A(n9872), .ZN(n9932) );
  INV_X1 U11015 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9874) );
  AOI22_X1 U11016 ( .A1(n9930), .A2(n9932), .B1(n9874), .B2(n9928), .ZN(
        P2_U3451) );
  AOI21_X1 U11017 ( .B1(n9927), .B2(n9878), .A(n9877), .ZN(n9934) );
  INV_X1 U11018 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9879) );
  AOI22_X1 U11019 ( .A1(n9930), .A2(n9934), .B1(n9879), .B2(n9928), .ZN(
        P2_U3460) );
  OAI211_X1 U11020 ( .C1(n9882), .C2(n9921), .A(n9881), .B(n9880), .ZN(n9883)
         );
  AOI21_X1 U11021 ( .B1(n9927), .B2(n9884), .A(n9883), .ZN(n9936) );
  INV_X1 U11022 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10043) );
  AOI22_X1 U11023 ( .A1(n9930), .A2(n9936), .B1(n10043), .B2(n9928), .ZN(
        P2_U3469) );
  NAND2_X1 U11024 ( .A1(n9886), .A2(n9885), .ZN(n9887) );
  OAI211_X1 U11025 ( .C1(n9922), .C2(n9889), .A(n9888), .B(n9887), .ZN(n9890)
         );
  AOI21_X1 U11026 ( .B1(n9927), .B2(n9891), .A(n9890), .ZN(n9938) );
  INV_X1 U11027 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10109) );
  AOI22_X1 U11028 ( .A1(n9930), .A2(n9938), .B1(n10109), .B2(n9928), .ZN(
        P2_U3472) );
  OAI22_X1 U11029 ( .A1(n9893), .A2(n9922), .B1(n9892), .B2(n9921), .ZN(n9894)
         );
  AOI21_X1 U11030 ( .B1(n9895), .B2(n9912), .A(n9894), .ZN(n9896) );
  AND2_X1 U11031 ( .A1(n9897), .A2(n9896), .ZN(n9939) );
  INV_X1 U11032 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9898) );
  AOI22_X1 U11033 ( .A1(n9930), .A2(n9939), .B1(n9898), .B2(n9928), .ZN(
        P2_U3475) );
  OAI22_X1 U11034 ( .A1(n9900), .A2(n9922), .B1(n9899), .B2(n9921), .ZN(n9901)
         );
  AOI21_X1 U11035 ( .B1(n9902), .B2(n9912), .A(n9901), .ZN(n9903) );
  AND2_X1 U11036 ( .A1(n9904), .A2(n9903), .ZN(n9940) );
  INV_X1 U11037 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9905) );
  AOI22_X1 U11038 ( .A1(n9930), .A2(n9940), .B1(n9905), .B2(n9928), .ZN(
        P2_U3478) );
  INV_X1 U11039 ( .A(n9906), .ZN(n9911) );
  OAI22_X1 U11040 ( .A1(n9908), .A2(n9922), .B1(n9907), .B2(n9921), .ZN(n9910)
         );
  AOI211_X1 U11041 ( .C1(n9912), .C2(n9911), .A(n9910), .B(n9909), .ZN(n9941)
         );
  INV_X1 U11042 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9913) );
  AOI22_X1 U11043 ( .A1(n9930), .A2(n9941), .B1(n9913), .B2(n9928), .ZN(
        P2_U3481) );
  OAI211_X1 U11044 ( .C1(n9916), .C2(n9921), .A(n9915), .B(n9914), .ZN(n9917)
         );
  AOI21_X1 U11045 ( .B1(n9918), .B2(n9927), .A(n9917), .ZN(n9942) );
  INV_X1 U11046 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9919) );
  AOI22_X1 U11047 ( .A1(n9930), .A2(n9942), .B1(n9919), .B2(n9928), .ZN(
        P2_U3484) );
  OAI22_X1 U11048 ( .A1(n9923), .A2(n9922), .B1(n4663), .B2(n9921), .ZN(n9925)
         );
  AOI211_X1 U11049 ( .C1(n9927), .C2(n9926), .A(n9925), .B(n9924), .ZN(n9944)
         );
  INV_X1 U11050 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9929) );
  AOI22_X1 U11051 ( .A1(n9930), .A2(n9944), .B1(n9929), .B2(n9928), .ZN(
        P2_U3487) );
  INV_X1 U11052 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9931) );
  AOI22_X1 U11053 ( .A1(n9945), .A2(n9932), .B1(n9931), .B2(n9943), .ZN(
        P2_U3520) );
  INV_X1 U11054 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9933) );
  AOI22_X1 U11055 ( .A1(n9945), .A2(n9934), .B1(n9933), .B2(n9943), .ZN(
        P2_U3523) );
  INV_X1 U11056 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9935) );
  AOI22_X1 U11057 ( .A1(n9945), .A2(n9936), .B1(n9935), .B2(n9943), .ZN(
        P2_U3526) );
  INV_X1 U11058 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9937) );
  AOI22_X1 U11059 ( .A1(n9945), .A2(n9938), .B1(n9937), .B2(n9943), .ZN(
        P2_U3527) );
  AOI22_X1 U11060 ( .A1(n9945), .A2(n9939), .B1(n6829), .B2(n9943), .ZN(
        P2_U3528) );
  AOI22_X1 U11061 ( .A1(n9945), .A2(n9940), .B1(n6866), .B2(n9943), .ZN(
        P2_U3529) );
  AOI22_X1 U11062 ( .A1(n9945), .A2(n9941), .B1(n6864), .B2(n9943), .ZN(
        P2_U3530) );
  AOI22_X1 U11063 ( .A1(n9945), .A2(n9942), .B1(n7069), .B2(n9943), .ZN(
        P2_U3531) );
  AOI22_X1 U11064 ( .A1(n9945), .A2(n9944), .B1(n7070), .B2(n9943), .ZN(
        P2_U3532) );
  INV_X1 U11065 ( .A(n9946), .ZN(n9947) );
  NAND2_X1 U11066 ( .A1(n9948), .A2(n9947), .ZN(n9949) );
  XOR2_X1 U11067 ( .A(n10233), .B(n9949), .Z(ADD_1071_U5) );
  XOR2_X1 U11068 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11069 ( .B1(n9952), .B2(n9951), .A(n9950), .ZN(ADD_1071_U56) );
  OAI21_X1 U11070 ( .B1(n9955), .B2(n9954), .A(n9953), .ZN(ADD_1071_U57) );
  OAI21_X1 U11071 ( .B1(n9958), .B2(n9957), .A(n9956), .ZN(ADD_1071_U58) );
  OAI21_X1 U11072 ( .B1(n9961), .B2(n9960), .A(n9959), .ZN(ADD_1071_U59) );
  OAI21_X1 U11073 ( .B1(n9964), .B2(n9963), .A(n9962), .ZN(ADD_1071_U60) );
  OAI21_X1 U11074 ( .B1(n9967), .B2(n9966), .A(n9965), .ZN(ADD_1071_U61) );
  AOI21_X1 U11075 ( .B1(n9970), .B2(n9969), .A(n9968), .ZN(ADD_1071_U62) );
  AOI21_X1 U11076 ( .B1(n9973), .B2(n9972), .A(n9971), .ZN(ADD_1071_U63) );
  AOI22_X1 U11077 ( .A1(n9975), .A2(keyinput108), .B1(keyinput97), .B2(n7567), 
        .ZN(n9974) );
  OAI221_X1 U11078 ( .B1(n9975), .B2(keyinput108), .C1(n7567), .C2(keyinput97), 
        .A(n9974), .ZN(n9985) );
  AOI22_X1 U11079 ( .A1(n10251), .A2(keyinput76), .B1(n9977), .B2(keyinput58), 
        .ZN(n9976) );
  OAI221_X1 U11080 ( .B1(n10251), .B2(keyinput76), .C1(n9977), .C2(keyinput58), 
        .A(n9976), .ZN(n9984) );
  AOI22_X1 U11081 ( .A1(n10266), .A2(keyinput90), .B1(n10261), .B2(keyinput1), 
        .ZN(n9978) );
  OAI221_X1 U11082 ( .B1(n10266), .B2(keyinput90), .C1(n10261), .C2(keyinput1), 
        .A(n9978), .ZN(n9983) );
  INV_X1 U11083 ( .A(SI_26_), .ZN(n9981) );
  AOI22_X1 U11084 ( .A1(n9981), .A2(keyinput54), .B1(keyinput56), .B2(n9980), 
        .ZN(n9979) );
  OAI221_X1 U11085 ( .B1(n9981), .B2(keyinput54), .C1(n9980), .C2(keyinput56), 
        .A(n9979), .ZN(n9982) );
  NOR4_X1 U11086 ( .A1(n9985), .A2(n9984), .A3(n9983), .A4(n9982), .ZN(n10026)
         );
  INV_X1 U11087 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9987) );
  AOI22_X1 U11088 ( .A1(n9988), .A2(keyinput7), .B1(keyinput68), .B2(n9987), 
        .ZN(n9986) );
  OAI221_X1 U11089 ( .B1(n9988), .B2(keyinput7), .C1(n9987), .C2(keyinput68), 
        .A(n9986), .ZN(n9996) );
  INV_X1 U11090 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n10253) );
  AOI22_X1 U11091 ( .A1(n10254), .A2(keyinput53), .B1(keyinput104), .B2(n10253), .ZN(n9989) );
  OAI221_X1 U11092 ( .B1(n10254), .B2(keyinput53), .C1(n10253), .C2(
        keyinput104), .A(n9989), .ZN(n9995) );
  INV_X1 U11093 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10249) );
  AOI22_X1 U11094 ( .A1(n10249), .A2(keyinput123), .B1(n10255), .B2(
        keyinput115), .ZN(n9990) );
  OAI221_X1 U11095 ( .B1(n10249), .B2(keyinput123), .C1(n10255), .C2(
        keyinput115), .A(n9990), .ZN(n9994) );
  XNOR2_X1 U11096 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput85), .ZN(n9992) );
  XNOR2_X1 U11097 ( .A(keyinput6), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n9991) );
  NAND2_X1 U11098 ( .A1(n9992), .A2(n9991), .ZN(n9993) );
  NOR4_X1 U11099 ( .A1(n9996), .A2(n9995), .A3(n9994), .A4(n9993), .ZN(n10025)
         );
  AOI22_X1 U11100 ( .A1(n9998), .A2(keyinput8), .B1(keyinput96), .B2(n10238), 
        .ZN(n9997) );
  OAI221_X1 U11101 ( .B1(n9998), .B2(keyinput8), .C1(n10238), .C2(keyinput96), 
        .A(n9997), .ZN(n10007) );
  INV_X1 U11102 ( .A(SI_24_), .ZN(n10000) );
  INV_X1 U11103 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10239) );
  AOI22_X1 U11104 ( .A1(n10000), .A2(keyinput86), .B1(keyinput59), .B2(n10239), 
        .ZN(n9999) );
  OAI221_X1 U11105 ( .B1(n10000), .B2(keyinput86), .C1(n10239), .C2(keyinput59), .A(n9999), .ZN(n10006) );
  AOI22_X1 U11106 ( .A1(n7070), .A2(keyinput47), .B1(n10204), .B2(keyinput105), 
        .ZN(n10001) );
  OAI221_X1 U11107 ( .B1(n7070), .B2(keyinput47), .C1(n10204), .C2(keyinput105), .A(n10001), .ZN(n10005) );
  XNOR2_X1 U11108 ( .A(P2_REG1_REG_27__SCAN_IN), .B(keyinput60), .ZN(n10003)
         );
  XNOR2_X1 U11109 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput110), .ZN(n10002) );
  NAND2_X1 U11110 ( .A1(n10003), .A2(n10002), .ZN(n10004) );
  NOR4_X1 U11111 ( .A1(n10007), .A2(n10006), .A3(n10005), .A4(n10004), .ZN(
        n10024) );
  AOI22_X1 U11112 ( .A1(n10010), .A2(keyinput24), .B1(keyinput57), .B2(n10009), 
        .ZN(n10008) );
  OAI221_X1 U11113 ( .B1(n10010), .B2(keyinput24), .C1(n10009), .C2(keyinput57), .A(n10008), .ZN(n10022) );
  AOI22_X1 U11114 ( .A1(n10013), .A2(keyinput42), .B1(n10012), .B2(keyinput70), 
        .ZN(n10011) );
  OAI221_X1 U11115 ( .B1(n10013), .B2(keyinput42), .C1(n10012), .C2(keyinput70), .A(n10011), .ZN(n10021) );
  AOI22_X1 U11116 ( .A1(n10016), .A2(keyinput94), .B1(n10015), .B2(keyinput52), 
        .ZN(n10014) );
  OAI221_X1 U11117 ( .B1(n10016), .B2(keyinput94), .C1(n10015), .C2(keyinput52), .A(n10014), .ZN(n10020) );
  XNOR2_X1 U11118 ( .A(P2_IR_REG_29__SCAN_IN), .B(keyinput40), .ZN(n10018) );
  XNOR2_X1 U11119 ( .A(P1_REG1_REG_15__SCAN_IN), .B(keyinput29), .ZN(n10017)
         );
  NAND2_X1 U11120 ( .A1(n10018), .A2(n10017), .ZN(n10019) );
  NOR4_X1 U11121 ( .A1(n10022), .A2(n10021), .A3(n10020), .A4(n10019), .ZN(
        n10023) );
  NAND4_X1 U11122 ( .A1(n10026), .A2(n10025), .A3(n10024), .A4(n10023), .ZN(
        n10186) );
  AOI22_X1 U11123 ( .A1(n10029), .A2(keyinput49), .B1(keyinput81), .B2(n10028), 
        .ZN(n10027) );
  OAI221_X1 U11124 ( .B1(n10029), .B2(keyinput49), .C1(n10028), .C2(keyinput81), .A(n10027), .ZN(n10038) );
  AOI22_X1 U11125 ( .A1(n10207), .A2(keyinput121), .B1(keyinput50), .B2(n10206), .ZN(n10030) );
  OAI221_X1 U11126 ( .B1(n10207), .B2(keyinput121), .C1(n10206), .C2(
        keyinput50), .A(n10030), .ZN(n10037) );
  XOR2_X1 U11127 ( .A(n10209), .B(keyinput14), .Z(n10035) );
  INV_X1 U11128 ( .A(SI_11_), .ZN(n10031) );
  XOR2_X1 U11129 ( .A(n10031), .B(keyinput72), .Z(n10034) );
  XNOR2_X1 U11130 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput0), .ZN(n10033) );
  XNOR2_X1 U11131 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput62), .ZN(n10032)
         );
  NAND4_X1 U11132 ( .A1(n10035), .A2(n10034), .A3(n10033), .A4(n10032), .ZN(
        n10036) );
  NOR3_X1 U11133 ( .A1(n10038), .A2(n10037), .A3(n10036), .ZN(n10078) );
  AOI22_X1 U11134 ( .A1(n10205), .A2(keyinput55), .B1(n10040), .B2(keyinput28), 
        .ZN(n10039) );
  OAI221_X1 U11135 ( .B1(n10205), .B2(keyinput55), .C1(n10040), .C2(keyinput28), .A(n10039), .ZN(n10050) );
  INV_X1 U11136 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n10042) );
  AOI22_X1 U11137 ( .A1(n10043), .A2(keyinput38), .B1(n10042), .B2(keyinput51), 
        .ZN(n10041) );
  OAI221_X1 U11138 ( .B1(n10043), .B2(keyinput38), .C1(n10042), .C2(keyinput51), .A(n10041), .ZN(n10049) );
  XNOR2_X1 U11139 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput100), .ZN(n10047) );
  XNOR2_X1 U11140 ( .A(P1_REG1_REG_26__SCAN_IN), .B(keyinput113), .ZN(n10046)
         );
  XNOR2_X1 U11141 ( .A(P2_IR_REG_27__SCAN_IN), .B(keyinput36), .ZN(n10045) );
  XNOR2_X1 U11142 ( .A(P1_REG0_REG_23__SCAN_IN), .B(keyinput125), .ZN(n10044)
         );
  NAND4_X1 U11143 ( .A1(n10047), .A2(n10046), .A3(n10045), .A4(n10044), .ZN(
        n10048) );
  NOR3_X1 U11144 ( .A1(n10050), .A2(n10049), .A3(n10048), .ZN(n10077) );
  AOI22_X1 U11145 ( .A1(n10053), .A2(keyinput33), .B1(keyinput117), .B2(n10052), .ZN(n10051) );
  OAI221_X1 U11146 ( .B1(n10053), .B2(keyinput33), .C1(n10052), .C2(
        keyinput117), .A(n10051), .ZN(n10062) );
  AOI22_X1 U11147 ( .A1(n10286), .A2(keyinput13), .B1(n10055), .B2(keyinput73), 
        .ZN(n10054) );
  OAI221_X1 U11148 ( .B1(n10286), .B2(keyinput13), .C1(n10055), .C2(keyinput73), .A(n10054), .ZN(n10061) );
  AOI22_X1 U11149 ( .A1(n4909), .A2(keyinput63), .B1(keyinput127), .B2(n10195), 
        .ZN(n10056) );
  OAI221_X1 U11150 ( .B1(n4909), .B2(keyinput63), .C1(n10195), .C2(keyinput127), .A(n10056), .ZN(n10060) );
  XNOR2_X1 U11151 ( .A(P1_REG3_REG_6__SCAN_IN), .B(keyinput82), .ZN(n10058) );
  XNOR2_X1 U11152 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput32), .ZN(n10057) );
  NAND2_X1 U11153 ( .A1(n10058), .A2(n10057), .ZN(n10059) );
  NOR4_X1 U11154 ( .A1(n10062), .A2(n10061), .A3(n10060), .A4(n10059), .ZN(
        n10076) );
  AOI22_X1 U11155 ( .A1(n10064), .A2(keyinput122), .B1(keyinput12), .B2(n6829), 
        .ZN(n10063) );
  OAI221_X1 U11156 ( .B1(n10064), .B2(keyinput122), .C1(n6829), .C2(keyinput12), .A(n10063), .ZN(n10074) );
  INV_X1 U11157 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n10194) );
  AOI22_X1 U11158 ( .A1(n10194), .A2(keyinput3), .B1(n8699), .B2(keyinput87), 
        .ZN(n10065) );
  OAI221_X1 U11159 ( .B1(n10194), .B2(keyinput3), .C1(n8699), .C2(keyinput87), 
        .A(n10065), .ZN(n10073) );
  AOI22_X1 U11160 ( .A1(n10067), .A2(keyinput89), .B1(n7197), .B2(keyinput27), 
        .ZN(n10066) );
  OAI221_X1 U11161 ( .B1(n10067), .B2(keyinput89), .C1(n7197), .C2(keyinput27), 
        .A(n10066), .ZN(n10072) );
  AOI22_X1 U11162 ( .A1(n10070), .A2(keyinput11), .B1(keyinput109), .B2(n10069), .ZN(n10068) );
  OAI221_X1 U11163 ( .B1(n10070), .B2(keyinput11), .C1(n10069), .C2(
        keyinput109), .A(n10068), .ZN(n10071) );
  NOR4_X1 U11164 ( .A1(n10074), .A2(n10073), .A3(n10072), .A4(n10071), .ZN(
        n10075) );
  NAND4_X1 U11165 ( .A1(n10078), .A2(n10077), .A3(n10076), .A4(n10075), .ZN(
        n10185) );
  AOI22_X1 U11166 ( .A1(n10196), .A2(keyinput21), .B1(n10080), .B2(keyinput126), .ZN(n10079) );
  OAI221_X1 U11167 ( .B1(n10196), .B2(keyinput21), .C1(n10080), .C2(
        keyinput126), .A(n10079), .ZN(n10081) );
  INV_X1 U11168 ( .A(n10081), .ZN(n10092) );
  INV_X1 U11169 ( .A(keyinput37), .ZN(n10082) );
  XNOR2_X1 U11170 ( .A(n10083), .B(n10082), .ZN(n10091) );
  INV_X1 U11171 ( .A(keyinput9), .ZN(n10084) );
  XNOR2_X1 U11172 ( .A(n10234), .B(n10084), .ZN(n10090) );
  XNOR2_X1 U11173 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput80), .ZN(n10088) );
  XNOR2_X1 U11174 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput67), .ZN(n10087) );
  XNOR2_X1 U11175 ( .A(P2_IR_REG_6__SCAN_IN), .B(keyinput98), .ZN(n10086) );
  XNOR2_X1 U11176 ( .A(P1_REG1_REG_23__SCAN_IN), .B(keyinput84), .ZN(n10085)
         );
  AND4_X1 U11177 ( .A1(n10088), .A2(n10087), .A3(n10086), .A4(n10085), .ZN(
        n10089) );
  AND4_X1 U11178 ( .A1(n10092), .A2(n10091), .A3(n10090), .A4(n10089), .ZN(
        n10130) );
  AOI22_X1 U11179 ( .A1(n10192), .A2(keyinput16), .B1(keyinput48), .B2(n6329), 
        .ZN(n10093) );
  OAI221_X1 U11180 ( .B1(n10192), .B2(keyinput16), .C1(n6329), .C2(keyinput48), 
        .A(n10093), .ZN(n10103) );
  AOI22_X1 U11181 ( .A1(n10095), .A2(keyinput92), .B1(n10193), .B2(keyinput95), 
        .ZN(n10094) );
  OAI221_X1 U11182 ( .B1(n10095), .B2(keyinput92), .C1(n10193), .C2(keyinput95), .A(n10094), .ZN(n10102) );
  XOR2_X1 U11183 ( .A(n10096), .B(keyinput17), .Z(n10100) );
  XNOR2_X1 U11184 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput18), .ZN(n10099)
         );
  XNOR2_X1 U11185 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(keyinput39), .ZN(n10098)
         );
  XNOR2_X1 U11186 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput30), .ZN(n10097) );
  NAND4_X1 U11187 ( .A1(n10100), .A2(n10099), .A3(n10098), .A4(n10097), .ZN(
        n10101) );
  NOR3_X1 U11188 ( .A1(n10103), .A2(n10102), .A3(n10101), .ZN(n10129) );
  INV_X1 U11189 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10216) );
  AOI22_X1 U11190 ( .A1(n7512), .A2(keyinput93), .B1(n10216), .B2(keyinput116), 
        .ZN(n10104) );
  OAI221_X1 U11191 ( .B1(n7512), .B2(keyinput93), .C1(n10216), .C2(keyinput116), .A(n10104), .ZN(n10114) );
  AOI22_X1 U11192 ( .A1(n10107), .A2(keyinput74), .B1(n10106), .B2(keyinput120), .ZN(n10105) );
  OAI221_X1 U11193 ( .B1(n10107), .B2(keyinput74), .C1(n10106), .C2(
        keyinput120), .A(n10105), .ZN(n10113) );
  AOI22_X1 U11194 ( .A1(n6485), .A2(keyinput111), .B1(keyinput118), .B2(n10109), .ZN(n10108) );
  OAI221_X1 U11195 ( .B1(n6485), .B2(keyinput111), .C1(n10109), .C2(
        keyinput118), .A(n10108), .ZN(n10112) );
  AOI22_X1 U11196 ( .A1(n10290), .A2(keyinput66), .B1(n7046), .B2(keyinput61), 
        .ZN(n10110) );
  OAI221_X1 U11197 ( .B1(n10290), .B2(keyinput66), .C1(n7046), .C2(keyinput61), 
        .A(n10110), .ZN(n10111) );
  NOR4_X1 U11198 ( .A1(n10114), .A2(n10113), .A3(n10112), .A4(n10111), .ZN(
        n10128) );
  AOI22_X1 U11199 ( .A1(n10116), .A2(keyinput19), .B1(n5309), .B2(keyinput101), 
        .ZN(n10115) );
  OAI221_X1 U11200 ( .B1(n10116), .B2(keyinput19), .C1(n5309), .C2(keyinput101), .A(n10115), .ZN(n10126) );
  INV_X1 U11201 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n10118) );
  AOI22_X1 U11202 ( .A1(n10119), .A2(keyinput102), .B1(n10118), .B2(keyinput69), .ZN(n10117) );
  OAI221_X1 U11203 ( .B1(n10119), .B2(keyinput102), .C1(n10118), .C2(
        keyinput69), .A(n10117), .ZN(n10125) );
  XNOR2_X1 U11204 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput77), .ZN(n10123) );
  XNOR2_X1 U11205 ( .A(P1_STATE_REG_SCAN_IN), .B(keyinput31), .ZN(n10122) );
  XNOR2_X1 U11206 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput5), .ZN(n10121) );
  XNOR2_X1 U11207 ( .A(keyinput78), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n10120) );
  NAND4_X1 U11208 ( .A1(n10123), .A2(n10122), .A3(n10121), .A4(n10120), .ZN(
        n10124) );
  NOR3_X1 U11209 ( .A1(n10126), .A2(n10125), .A3(n10124), .ZN(n10127) );
  NAND4_X1 U11210 ( .A1(n10130), .A2(n10129), .A3(n10128), .A4(n10127), .ZN(
        n10184) );
  AOI22_X1 U11211 ( .A1(n10133), .A2(keyinput45), .B1(n10132), .B2(keyinput88), 
        .ZN(n10131) );
  OAI221_X1 U11212 ( .B1(n10133), .B2(keyinput45), .C1(n10132), .C2(keyinput88), .A(n10131), .ZN(n10142) );
  AOI22_X1 U11213 ( .A1(n10219), .A2(keyinput25), .B1(keyinput83), .B2(n8060), 
        .ZN(n10134) );
  OAI221_X1 U11214 ( .B1(n10219), .B2(keyinput25), .C1(n8060), .C2(keyinput83), 
        .A(n10134), .ZN(n10141) );
  AOI22_X1 U11215 ( .A1(n7079), .A2(keyinput79), .B1(n10136), .B2(keyinput103), 
        .ZN(n10135) );
  OAI221_X1 U11216 ( .B1(n7079), .B2(keyinput79), .C1(n10136), .C2(keyinput103), .A(n10135), .ZN(n10140) );
  AOI22_X1 U11217 ( .A1(n10138), .A2(keyinput4), .B1(keyinput112), .B2(n7847), 
        .ZN(n10137) );
  OAI221_X1 U11218 ( .B1(n10138), .B2(keyinput4), .C1(n7847), .C2(keyinput112), 
        .A(n10137), .ZN(n10139) );
  NOR4_X1 U11219 ( .A1(n10142), .A2(n10141), .A3(n10140), .A4(n10139), .ZN(
        n10182) );
  AOI22_X1 U11220 ( .A1(n10232), .A2(keyinput91), .B1(keyinput106), .B2(n7204), 
        .ZN(n10143) );
  OAI221_X1 U11221 ( .B1(n10232), .B2(keyinput91), .C1(n7204), .C2(keyinput106), .A(n10143), .ZN(n10155) );
  AOI22_X1 U11222 ( .A1(n10214), .A2(keyinput15), .B1(n10145), .B2(keyinput75), 
        .ZN(n10144) );
  OAI221_X1 U11223 ( .B1(n10214), .B2(keyinput15), .C1(n10145), .C2(keyinput75), .A(n10144), .ZN(n10154) );
  INV_X1 U11224 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n10148) );
  INV_X1 U11225 ( .A(SI_31_), .ZN(n10147) );
  AOI22_X1 U11226 ( .A1(n10148), .A2(keyinput10), .B1(keyinput107), .B2(n10147), .ZN(n10146) );
  OAI221_X1 U11227 ( .B1(n10148), .B2(keyinput10), .C1(n10147), .C2(
        keyinput107), .A(n10146), .ZN(n10153) );
  INV_X1 U11228 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n10151) );
  AOI22_X1 U11229 ( .A1(n10151), .A2(keyinput65), .B1(keyinput23), .B2(n10150), 
        .ZN(n10149) );
  OAI221_X1 U11230 ( .B1(n10151), .B2(keyinput65), .C1(n10150), .C2(keyinput23), .A(n10149), .ZN(n10152) );
  NOR4_X1 U11231 ( .A1(n10155), .A2(n10154), .A3(n10153), .A4(n10152), .ZN(
        n10181) );
  AOI22_X1 U11232 ( .A1(n10223), .A2(keyinput35), .B1(keyinput64), .B2(n6798), 
        .ZN(n10156) );
  OAI221_X1 U11233 ( .B1(n10223), .B2(keyinput35), .C1(n6798), .C2(keyinput64), 
        .A(n10156), .ZN(n10167) );
  AOI22_X1 U11234 ( .A1(n10159), .A2(keyinput34), .B1(keyinput20), .B2(n10158), 
        .ZN(n10157) );
  OAI221_X1 U11235 ( .B1(n10159), .B2(keyinput34), .C1(n10158), .C2(keyinput20), .A(n10157), .ZN(n10166) );
  AOI22_X1 U11236 ( .A1(n10250), .A2(keyinput71), .B1(keyinput2), .B2(n10161), 
        .ZN(n10160) );
  OAI221_X1 U11237 ( .B1(n10250), .B2(keyinput71), .C1(n10161), .C2(keyinput2), 
        .A(n10160), .ZN(n10165) );
  XNOR2_X1 U11238 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput99), .ZN(n10163) );
  XNOR2_X1 U11239 ( .A(SI_1_), .B(keyinput44), .ZN(n10162) );
  NAND2_X1 U11240 ( .A1(n10163), .A2(n10162), .ZN(n10164) );
  NOR4_X1 U11241 ( .A1(n10167), .A2(n10166), .A3(n10165), .A4(n10164), .ZN(
        n10180) );
  INV_X1 U11242 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n10169) );
  AOI22_X1 U11243 ( .A1(n10240), .A2(keyinput41), .B1(keyinput124), .B2(n10169), .ZN(n10168) );
  OAI221_X1 U11244 ( .B1(n10240), .B2(keyinput41), .C1(n10169), .C2(
        keyinput124), .A(n10168), .ZN(n10178) );
  AOI22_X1 U11245 ( .A1(n10233), .A2(keyinput22), .B1(n10221), .B2(keyinput119), .ZN(n10170) );
  OAI221_X1 U11246 ( .B1(n10233), .B2(keyinput22), .C1(n10221), .C2(
        keyinput119), .A(n10170), .ZN(n10177) );
  AOI22_X1 U11247 ( .A1(n10172), .A2(keyinput46), .B1(keyinput26), .B2(n10222), 
        .ZN(n10171) );
  OAI221_X1 U11248 ( .B1(n10172), .B2(keyinput46), .C1(n10222), .C2(keyinput26), .A(n10171), .ZN(n10176) );
  XNOR2_X1 U11249 ( .A(P2_REG0_REG_24__SCAN_IN), .B(keyinput43), .ZN(n10174)
         );
  XNOR2_X1 U11250 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput114), .ZN(n10173) );
  NAND2_X1 U11251 ( .A1(n10174), .A2(n10173), .ZN(n10175) );
  NOR4_X1 U11252 ( .A1(n10178), .A2(n10177), .A3(n10176), .A4(n10175), .ZN(
        n10179) );
  NAND4_X1 U11253 ( .A1(n10182), .A2(n10181), .A3(n10180), .A4(n10179), .ZN(
        n10183) );
  NOR4_X1 U11254 ( .A1(n10186), .A2(n10185), .A3(n10184), .A4(n10183), .ZN(
        n10191) );
  AOI22_X1 U11255 ( .A1(n10189), .A2(n10188), .B1(P1_REG1_REG_11__SCAN_IN), 
        .B2(n10187), .ZN(n10190) );
  XNOR2_X1 U11256 ( .A(n10191), .B(n10190), .ZN(n10278) );
  NAND4_X1 U11257 ( .A1(P1_REG1_REG_16__SCAN_IN), .A2(P1_REG2_REG_15__SCAN_IN), 
        .A3(P2_REG3_REG_20__SCAN_IN), .A4(n8699), .ZN(n10202) );
  NAND4_X1 U11258 ( .A1(SI_14_), .A2(n10193), .A3(n10192), .A4(n6329), .ZN(
        n10201) );
  NAND4_X1 U11259 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_REG1_REG_8__SCAN_IN), 
        .A3(n10195), .A4(n10194), .ZN(n10200) );
  NAND4_X1 U11260 ( .A1(n10198), .A2(n10197), .A3(n10196), .A4(
        P2_REG3_REG_27__SCAN_IN), .ZN(n10199) );
  NOR4_X1 U11261 ( .A1(n10202), .A2(n10201), .A3(n10200), .A4(n10199), .ZN(
        n10276) );
  NAND4_X1 U11262 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(
        P1_DATAO_REG_29__SCAN_IN), .A3(n10204), .A4(n10203), .ZN(n10212) );
  NAND4_X1 U11263 ( .A1(n10208), .A2(n10207), .A3(n10206), .A4(n10205), .ZN(
        n10211) );
  NAND4_X1 U11264 ( .A1(P2_REG0_REG_20__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), 
        .A3(P2_REG2_REG_3__SCAN_IN), .A4(n10209), .ZN(n10210) );
  NOR4_X1 U11265 ( .A1(P2_REG0_REG_6__SCAN_IN), .A2(n10212), .A3(n10211), .A4(
        n10210), .ZN(n10213) );
  AND4_X1 U11266 ( .A1(n4760), .A2(P1_REG0_REG_23__SCAN_IN), .A3(
        P1_REG2_REG_24__SCAN_IN), .A4(n10213), .ZN(n10275) );
  NOR4_X1 U11267 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(P2_REG0_REG_19__SCAN_IN), 
        .A3(SI_31_), .A4(n10214), .ZN(n10215) );
  NAND3_X1 U11268 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_REG2_REG_18__SCAN_IN), 
        .A3(n10215), .ZN(n10231) );
  NAND4_X1 U11269 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_REG0_REG_7__SCAN_IN), 
        .A3(n10216), .A4(n7512), .ZN(n10217) );
  NOR3_X1 U11270 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(n10218), .A3(n10217), .ZN(
        n10229) );
  NAND4_X1 U11271 ( .A1(P1_REG0_REG_20__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .A3(P2_REG1_REG_26__SCAN_IN), .A4(P2_REG2_REG_12__SCAN_IN), .ZN(n10227) );
  NAND4_X1 U11272 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_REG3_REG_24__SCAN_IN), 
        .A3(n10219), .A4(n5309), .ZN(n10226) );
  INV_X1 U11273 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n10220) );
  NAND4_X1 U11274 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(n10222), .A3(n10221), 
        .A4(n10220), .ZN(n10225) );
  NAND4_X1 U11275 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(P2_D_REG_0__SCAN_IN), 
        .A3(P2_REG2_REG_4__SCAN_IN), .A4(n10223), .ZN(n10224) );
  NOR4_X1 U11276 ( .A1(n10227), .A2(n10226), .A3(n10225), .A4(n10224), .ZN(
        n10228) );
  NAND4_X1 U11277 ( .A1(P1_REG1_REG_13__SCAN_IN), .A2(P2_REG1_REG_13__SCAN_IN), 
        .A3(n10229), .A4(n10228), .ZN(n10230) );
  NOR4_X1 U11278 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(n10232), .A3(n10231), 
        .A4(n10230), .ZN(n10274) );
  NAND4_X1 U11279 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P2_ADDR_REG_7__SCAN_IN), 
        .A3(P1_ADDR_REG_14__SCAN_IN), .A4(n10290), .ZN(n10272) );
  NAND4_X1 U11280 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .A3(n10234), .A4(n10233), .ZN(n10271) );
  NAND4_X1 U11281 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), 
        .A3(P1_IR_REG_3__SCAN_IN), .A4(P1_U3084), .ZN(n10235) );
  NOR3_X1 U11282 ( .A1(n10236), .A2(P1_IR_REG_26__SCAN_IN), .A3(n10235), .ZN(
        n10237) );
  NAND3_X1 U11283 ( .A1(n10237), .A2(P1_IR_REG_14__SCAN_IN), .A3(
        P1_IR_REG_18__SCAN_IN), .ZN(n10243) );
  NAND4_X1 U11284 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .A3(n10239), .A4(n10238), .ZN(n10242) );
  NAND4_X1 U11285 ( .A1(P1_D_REG_0__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(n10240), .ZN(n10241) );
  NOR3_X1 U11286 ( .A1(n10243), .A2(n10242), .A3(n10241), .ZN(n10244) );
  NAND4_X1 U11287 ( .A1(n10247), .A2(n10246), .A3(n10245), .A4(n10244), .ZN(
        n10270) );
  NAND4_X1 U11288 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(P1_REG2_REG_6__SCAN_IN), 
        .A3(P1_REG1_REG_5__SCAN_IN), .A4(P1_REG2_REG_4__SCAN_IN), .ZN(n10248)
         );
  NOR3_X1 U11289 ( .A1(P1_REG0_REG_6__SCAN_IN), .A2(P1_REG2_REG_5__SCAN_IN), 
        .A3(n10248), .ZN(n10268) );
  NOR4_X1 U11290 ( .A1(SI_26_), .A2(P1_REG3_REG_27__SCAN_IN), .A3(
        P2_REG2_REG_7__SCAN_IN), .A4(n10249), .ZN(n10259) );
  NOR4_X1 U11291 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(n10251), .A3(n10250), .A4(
        n7567), .ZN(n10258) );
  NOR4_X1 U11292 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(SI_24_), .A3(
        P2_REG1_REG_12__SCAN_IN), .A4(n10252), .ZN(n10257) );
  NOR4_X1 U11293 ( .A1(P2_REG0_REG_22__SCAN_IN), .A2(n10255), .A3(n10254), 
        .A4(n10253), .ZN(n10256) );
  NAND4_X1 U11294 ( .A1(n10259), .A2(n10258), .A3(n10257), .A4(n10256), .ZN(
        n10265) );
  NAND4_X1 U11295 ( .A1(n4909), .A2(n10261), .A3(n10260), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n10264) );
  NAND4_X1 U11296 ( .A1(n10029), .A2(n10262), .A3(SI_11_), .A4(
        P1_REG3_REG_6__SCAN_IN), .ZN(n10263) );
  NOR3_X1 U11297 ( .A1(n10265), .A2(n10264), .A3(n10263), .ZN(n10267) );
  NAND4_X1 U11298 ( .A1(SI_1_), .A2(n10268), .A3(n10267), .A4(n10266), .ZN(
        n10269) );
  NOR4_X1 U11299 ( .A1(n10272), .A2(n10271), .A3(n10270), .A4(n10269), .ZN(
        n10273) );
  NAND4_X1 U11300 ( .A1(n10276), .A2(n10275), .A3(n10274), .A4(n10273), .ZN(
        n10277) );
  XNOR2_X1 U11301 ( .A(n10278), .B(n10277), .ZN(P1_U3534) );
  XOR2_X1 U11302 ( .A(n10279), .B(P1_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11303 ( .A1(n10281), .A2(n10280), .ZN(n10282) );
  XOR2_X1 U11304 ( .A(n10282), .B(P1_ADDR_REG_5__SCAN_IN), .Z(ADD_1071_U51) );
  XOR2_X1 U11305 ( .A(n10283), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  OAI21_X1 U11306 ( .B1(n10286), .B2(n10285), .A(n10284), .ZN(n10287) );
  XNOR2_X1 U11307 ( .A(n10287), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11308 ( .B1(n10290), .B2(n10289), .A(n10288), .ZN(ADD_1071_U47) );
  XOR2_X1 U11309 ( .A(n10291), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  XOR2_X1 U11310 ( .A(n10293), .B(n10292), .Z(ADD_1071_U54) );
  XOR2_X1 U11311 ( .A(n10295), .B(n10294), .Z(ADD_1071_U53) );
  XNOR2_X1 U11312 ( .A(n10297), .B(n10296), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4909 ( .A(n7817), .Z(n4496) );
  CLKBUF_X1 U5195 ( .A(n6972), .Z(n4500) );
endmodule

