

module b15_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD, 
        READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN, 
        M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN, 
        STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN, 
        W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N,
         BS16_N, READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN,
         CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN,
         REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN,
         FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3431, n3432, n3434, n3435, n3436, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116;

  OAI21_X1 U34650 ( .B1(n5306), .B2(n5305), .A(n5304), .ZN(n5721) );
  OR2_X1 U3466 ( .A1(n3455), .A2(n4492), .ZN(n4493) );
  INV_X1 U3467 ( .A(n6397), .ZN(n6410) );
  CLKBUF_X2 U34690 ( .A(n4229), .Z(n3435) );
  BUF_X2 U34700 ( .A(n3902), .Z(n5076) );
  BUF_X2 U34710 ( .A(n3896), .Z(n5051) );
  CLKBUF_X2 U34720 ( .A(n3952), .Z(n5068) );
  CLKBUF_X2 U34730 ( .A(n3590), .Z(n5088) );
  CLKBUF_X2 U34740 ( .A(n3628), .Z(n5063) );
  CLKBUF_X2 U3475 ( .A(n4273), .Z(n5080) );
  CLKBUF_X1 U3476 ( .A(n5037), .Z(n5078) );
  CLKBUF_X2 U3478 ( .A(n3668), .Z(n4586) );
  BUF_X1 U3479 ( .A(n3642), .Z(n6872) );
  AND4_X1 U3480 ( .A1(n3583), .A2(n3582), .A3(n3581), .A4(n3580), .ZN(n3589)
         );
  AND2_X2 U3481 ( .A1(n4592), .A2(n4687), .ZN(n3628) );
  NAND2_X1 U3483 ( .A1(n6914), .A2(n3651), .ZN(n4551) );
  AND2_X1 U3484 ( .A1(n3822), .A2(n3821), .ZN(n3835) );
  AND2_X1 U3485 ( .A1(n3553), .A2(n4136), .ZN(n4072) );
  NOR2_X1 U3486 ( .A1(n4037), .A2(n4036), .ZN(n4038) );
  AND4_X1 U3487 ( .A1(n3598), .A2(n3597), .A3(n3596), .A4(n3595), .ZN(n3441)
         );
  AND3_X1 U3488 ( .A1(n3586), .A2(n3585), .A3(n3584), .ZN(n3588) );
  OR2_X1 U3489 ( .A1(n4180), .A2(n4304), .ZN(n4187) );
  AND2_X1 U3490 ( .A1(n3640), .A2(n3639), .ZN(n3815) );
  AND2_X2 U3491 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4592) );
  NAND2_X1 U3492 ( .A1(n3990), .A2(n3989), .ZN(n4702) );
  OR2_X1 U3493 ( .A1(n4905), .A2(n4288), .ZN(n4289) );
  NAND2_X1 U3494 ( .A1(n3642), .A2(n3621), .ZN(n4131) );
  INV_X2 U3495 ( .A(n5782), .ZN(n5692) );
  OAI21_X1 U3496 ( .B1(n4180), .B2(n4046), .A(n4045), .ZN(n4047) );
  AND2_X1 U3497 ( .A1(n3579), .A2(n3578), .ZN(n5239) );
  INV_X1 U3498 ( .A(n3643), .ZN(n7000) );
  OAI21_X1 U3499 ( .B1(n5735), .B2(n7005), .A(n5734), .ZN(n5736) );
  INV_X1 U3500 ( .A(n6419), .ZN(n6391) );
  AOI211_X1 U3501 ( .C1(n5826), .C2(n6398), .A(n5762), .B(n5761), .ZN(n5763)
         );
  NAND2_X1 U3502 ( .A1(n4153), .A2(n6482), .ZN(n3918) );
  XNOR2_X2 U3503 ( .A(n3698), .B(n4548), .ZN(n4827) );
  AOI21_X2 U3504 ( .B1(n6541), .B2(n4085), .A(n3968), .ZN(n6087) );
  NAND2_X2 U3505 ( .A1(n3894), .A2(n3893), .ZN(n5924) );
  AND2_X1 U3506 ( .A1(n4591), .A2(n4690), .ZN(n3431) );
  AND2_X2 U3507 ( .A1(n4591), .A2(n4690), .ZN(n5036) );
  AND2_X2 U3508 ( .A1(n3479), .A2(n4687), .ZN(n3895) );
  AND2_X1 U3509 ( .A1(n3485), .A2(n4592), .ZN(n3432) );
  NOR2_X2 U3510 ( .A1(n5709), .A2(n4522), .ZN(n4525) );
  NAND2_X2 U3511 ( .A1(n5719), .A2(n5717), .ZN(n5709) );
  INV_X1 U3512 ( .A(n5166), .ZN(n5168) );
  CLKBUF_X1 U3513 ( .A(n5728), .Z(n5729) );
  AND2_X1 U3514 ( .A1(n5750), .A2(n4119), .ZN(n3447) );
  AND2_X1 U3515 ( .A1(n5791), .A2(n4114), .ZN(n5781) );
  INV_X1 U3516 ( .A(n4095), .ZN(n5782) );
  NAND2_X1 U3517 ( .A1(n4187), .A2(n4186), .ZN(n4654) );
  NAND2_X1 U3518 ( .A1(n4063), .A2(n4062), .ZN(n4088) );
  OAI21_X1 U3519 ( .B1(n5924), .B2(INSTADDRPOINTER_REG_1__SCAN_IN), .A(n5925), 
        .ZN(n3930) );
  AND2_X2 U3520 ( .A1(n4620), .A2(n4735), .ZN(n4721) );
  AND2_X1 U3521 ( .A1(n4638), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5925)
         );
  NOR2_X1 U3522 ( .A1(n4909), .A2(n4908), .ZN(n3742) );
  NAND2_X1 U3523 ( .A1(n4693), .A2(n3946), .ZN(n4676) );
  NAND2_X1 U3524 ( .A1(n3866), .A2(n3865), .ZN(n3932) );
  NAND2_X1 U3525 ( .A1(n3918), .A2(n3876), .ZN(n3931) );
  AND2_X1 U3526 ( .A1(n5193), .A2(n5192), .ZN(n5195) );
  OR2_X1 U3527 ( .A1(n4650), .A2(n4649), .ZN(n3715) );
  AND3_X1 U3528 ( .A1(n3803), .A2(n5240), .A3(n4595), .ZN(n4137) );
  AND2_X1 U3529 ( .A1(n4551), .A2(n3642), .ZN(n3817) );
  NOR2_X2 U3530 ( .A1(n3644), .A2(n7000), .ZN(n4668) );
  OR2_X1 U3531 ( .A1(n4131), .A2(n3820), .ZN(n3821) );
  NAND4_X2 U3532 ( .A1(n3495), .A2(n3494), .A3(n3493), .A4(n3492), .ZN(n3668)
         );
  AND4_X1 U3533 ( .A1(n3478), .A2(n3477), .A3(n3476), .A4(n3475), .ZN(n3494)
         );
  AND4_X1 U3534 ( .A1(n3483), .A2(n3482), .A3(n3481), .A4(n3480), .ZN(n3493)
         );
  BUF_X2 U3535 ( .A(n3853), .Z(n5087) );
  BUF_X2 U3536 ( .A(n3858), .Z(n5079) );
  BUF_X2 U3537 ( .A(n3895), .Z(n5077) );
  BUF_X2 U3538 ( .A(n3951), .Z(n3853) );
  INV_X2 U3539 ( .A(n3623), .ZN(n3434) );
  AND2_X2 U3541 ( .A1(n6137), .A2(n6482), .ZN(n6277) );
  OR2_X2 U3542 ( .A1(n6512), .A2(n5955), .ZN(n5952) );
  INV_X1 U3543 ( .A(n6541), .ZN(n3436) );
  OAI21_X1 U3545 ( .B1(n5169), .B2(n5168), .A(n5303), .ZN(n5735) );
  AND2_X1 U3546 ( .A1(n5414), .A2(n5416), .ZN(n3438) );
  AND2_X2 U3547 ( .A1(n5414), .A2(n5416), .ZN(n3439) );
  BUF_X4 U3548 ( .A(n4146), .Z(n6663) );
  AND2_X1 U3549 ( .A1(n5414), .A2(n5416), .ZN(n5407) );
  BUF_X2 U3550 ( .A(n5036), .Z(n5075) );
  AND2_X1 U3551 ( .A1(n3932), .A2(n3931), .ZN(n3962) );
  OAI21_X1 U3552 ( .B1(n5416), .B2(n5414), .A(n5415), .ZN(n6399) );
  NAND2_X1 U3553 ( .A1(n3730), .A2(n3729), .ZN(n4860) );
  AND2_X2 U3554 ( .A1(n6068), .A2(n5423), .ZN(n5422) );
  NAND2_X2 U3555 ( .A1(n3440), .A2(n3441), .ZN(n3637) );
  AND4_X1 U3556 ( .A1(n3594), .A2(n3593), .A3(n3592), .A4(n3591), .ZN(n3440)
         );
  AND2_X2 U3557 ( .A1(n4840), .A2(n4839), .ZN(n4842) );
  NAND2_X2 U3558 ( .A1(n3991), .A2(n4702), .ZN(n4037) );
  NAND2_X1 U3559 ( .A1(n5791), .A2(n3442), .ZN(n5750) );
  AND2_X1 U3560 ( .A1(n4114), .A2(n4117), .ZN(n3442) );
  AND2_X2 U3561 ( .A1(n5176), .A2(n5175), .ZN(n5174) );
  OAI211_X2 U3562 ( .C1(n5663), .C2(n5678), .A(n5662), .B(n5661), .ZN(n5664)
         );
  OAI21_X2 U3563 ( .B1(n4701), .B2(n4304), .A(n4286), .ZN(n4160) );
  XNOR2_X2 U3564 ( .A(n5225), .B(n5224), .ZN(n5683) );
  XNOR2_X2 U3565 ( .A(n4905), .B(n4288), .ZN(n4976) );
  NAND2_X1 U3566 ( .A1(n5782), .A2(n3443), .ZN(n3444) );
  NAND2_X1 U3567 ( .A1(n5004), .A2(n5003), .ZN(n3445) );
  NAND2_X1 U3568 ( .A1(n3444), .A2(n3445), .ZN(n5006) );
  INV_X1 U3569 ( .A(n5003), .ZN(n3443) );
  NAND2_X1 U3570 ( .A1(n5750), .A2(n4119), .ZN(n3446) );
  NAND2_X1 U3571 ( .A1(n5750), .A2(n4119), .ZN(n6124) );
  AOI21_X1 U3572 ( .B1(n3939), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3943), 
        .ZN(n3944) );
  XNOR2_X1 U3573 ( .A(n4047), .B(n4778), .ZN(n4776) );
  XNOR2_X1 U3574 ( .A(n4021), .B(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4846)
         );
  NAND4_X1 U3575 ( .A1(n3495), .A2(n3494), .A3(n3493), .A4(n3492), .ZN(n3448)
         );
  NOR2_X2 U3576 ( .A1(n4525), .A2(n5686), .ZN(n5003) );
  AND2_X1 U3577 ( .A1(n3485), .A2(n3484), .ZN(n3449) );
  AND2_X1 U3578 ( .A1(n3485), .A2(n3484), .ZN(n3450) );
  AND2_X1 U3579 ( .A1(n3485), .A2(n3484), .ZN(n3852) );
  OAI21_X2 U3581 ( .B1(n4845), .B2(n4846), .A(n4022), .ZN(n4775) );
  NAND2_X1 U3582 ( .A1(n6831), .A2(n4564), .ZN(n3452) );
  NAND2_X1 U3583 ( .A1(n6831), .A2(n4564), .ZN(n3453) );
  AOI21_X2 U3584 ( .B1(n5800), .B2(n4113), .A(n3463), .ZN(n5791) );
  AOI21_X2 U3585 ( .B1(n5728), .B2(n5730), .A(n4124), .ZN(n5719) );
  INV_X1 U3586 ( .A(n3965), .ZN(n3874) );
  INV_X1 U3587 ( .A(n4035), .ZN(n4036) );
  NAND2_X1 U3588 ( .A1(n4038), .A2(n4039), .ZN(n4065) );
  NAND2_X1 U3589 ( .A1(n4564), .A2(n6790), .ZN(n3660) );
  INV_X1 U3590 ( .A(n4304), .ZN(n4314) );
  OR2_X2 U3591 ( .A1(n3634), .A2(n3633), .ZN(n3925) );
  OR2_X1 U3592 ( .A1(n3913), .A2(n3874), .ZN(n3865) );
  NAND2_X1 U3593 ( .A1(n6545), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3873) );
  NAND2_X1 U3594 ( .A1(n6872), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3913) );
  OR2_X1 U3595 ( .A1(n3503), .A2(n6459), .ZN(n3513) );
  AOI22_X1 U3596 ( .A1(n3952), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3896), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3539) );
  AND2_X2 U3598 ( .A1(n6955), .A2(n3621), .ZN(n3644) );
  AND2_X1 U3599 ( .A1(n5279), .A2(n5281), .ZN(n5266) );
  AND2_X1 U3600 ( .A1(n5145), .A2(n5406), .ZN(n5289) );
  INV_X1 U3601 ( .A(n5149), .ZN(n5134) );
  BUF_X1 U3602 ( .A(n3621), .Z(n3889) );
  NAND2_X1 U3603 ( .A1(n6955), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4304) );
  INV_X1 U3604 ( .A(n4064), .ZN(n4062) );
  INV_X1 U3605 ( .A(n4065), .ZN(n4063) );
  OR2_X1 U3606 ( .A1(n3988), .A2(n3987), .ZN(n4016) );
  AND2_X1 U3607 ( .A1(n3889), .A2(n4586), .ZN(n4085) );
  INV_X1 U3608 ( .A(n3992), .ZN(n3991) );
  NAND2_X1 U3609 ( .A1(n3913), .A2(n3873), .ZN(n4071) );
  OAI21_X1 U3610 ( .B1(n6150), .B2(n6472), .A(n6478), .ZN(n6544) );
  OR2_X1 U3611 ( .A1(n5239), .A2(n6487), .ZN(n4619) );
  CLKBUF_X1 U3612 ( .A(n3840), .Z(n5236) );
  AND2_X1 U3613 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n4423), .ZN(n4424)
         );
  INV_X1 U3614 ( .A(n4422), .ZN(n4423) );
  NAND2_X1 U3615 ( .A1(n3837), .A2(n3836), .ZN(n3868) );
  INV_X1 U3616 ( .A(n5228), .ZN(n4550) );
  NAND2_X1 U3617 ( .A1(n4585), .A2(n4584), .ZN(n4665) );
  INV_X1 U3618 ( .A(n4562), .ZN(n6465) );
  INV_X1 U3619 ( .A(n4286), .ZN(n5220) );
  NAND2_X1 U3620 ( .A1(n3455), .A2(n5167), .ZN(n5303) );
  NAND2_X1 U3621 ( .A1(n4424), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4470)
         );
  INV_X1 U3622 ( .A(n4657), .ZN(n4191) );
  OR2_X1 U3623 ( .A1(n5692), .A2(n4118), .ZN(n4119) );
  NOR2_X2 U3624 ( .A1(n4860), .A2(n4859), .ZN(n4879) );
  NAND2_X1 U3625 ( .A1(n3678), .A2(n3677), .ZN(n6199) );
  NAND2_X1 U3626 ( .A1(n4141), .A2(n4550), .ZN(n6217) );
  NAND2_X1 U3627 ( .A1(n3924), .A2(n3923), .ZN(n4761) );
  NAND2_X1 U3628 ( .A1(n6482), .A2(n6544), .ZN(n6546) );
  INV_X1 U3629 ( .A(n6546), .ZN(n6999) );
  INV_X1 U3630 ( .A(n6578), .ZN(n6732) );
  INV_X1 U3631 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6709) );
  INV_X2 U3632 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6720) );
  AND2_X1 U3633 ( .A1(n6371), .A2(n4503), .ZN(n6419) );
  BUF_X1 U3635 ( .A(n4761), .Z(n6723) );
  INV_X1 U3636 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6736) );
  INV_X1 U3637 ( .A(n7085), .ZN(n7084) );
  AND2_X1 U3638 ( .A1(n6626), .A2(n6723), .ZN(n6971) );
  NAND2_X1 U3639 ( .A1(n5508), .A2(n5507), .ZN(n5509) );
  CLKBUF_X1 U3640 ( .A(n5085), .Z(n5042) );
  NOR2_X1 U3641 ( .A1(n3549), .A2(n3558), .ZN(n3564) );
  OR2_X1 U3642 ( .A1(n3542), .A2(n5240), .ZN(n3563) );
  INV_X1 U3643 ( .A(n3548), .ZN(n3508) );
  NAND2_X1 U3644 ( .A1(n3614), .A2(n6955), .ZN(n3617) );
  NAND2_X1 U3645 ( .A1(n4034), .A2(n4033), .ZN(n4039) );
  OR2_X1 U3646 ( .A1(n3864), .A2(n3863), .ZN(n3965) );
  AND2_X2 U3647 ( .A1(n3487), .A2(n4690), .ZN(n3590) );
  AND2_X2 U3648 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4687) );
  NOR2_X1 U3649 ( .A1(n3838), .A2(n6545), .ZN(n4494) );
  NAND2_X1 U3650 ( .A1(n3514), .A2(n4694), .ZN(n3569) );
  INV_X1 U3651 ( .A(n3513), .ZN(n3514) );
  OR2_X1 U3652 ( .A1(n5236), .A2(n3646), .ZN(n3670) );
  NAND2_X1 U3653 ( .A1(n3849), .A2(n3466), .ZN(n3850) );
  INV_X1 U3654 ( .A(n3617), .ZN(n3830) );
  AND2_X1 U3655 ( .A1(n5146), .A2(n5289), .ZN(n5279) );
  NOR2_X1 U3656 ( .A1(n4322), .A2(n6350), .ZN(n4350) );
  NOR2_X1 U3657 ( .A1(n4228), .A2(n4867), .ZN(n4244) );
  OAI21_X1 U3658 ( .B1(n4039), .B2(n4038), .A(n4065), .ZN(n4180) );
  NOR2_X1 U3659 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3486) );
  INV_X1 U3660 ( .A(n3962), .ZN(n3961) );
  AND2_X1 U3661 ( .A1(n4072), .A2(n4085), .ZN(n3577) );
  NAND2_X1 U3662 ( .A1(n3505), .A2(n3504), .ZN(n3576) );
  CLKBUF_X1 U3663 ( .A(n3838), .Z(n4597) );
  CLKBUF_X1 U3664 ( .A(n4494), .Z(n4495) );
  NOR2_X1 U3665 ( .A1(n4871), .A2(n6340), .ZN(n4946) );
  INV_X1 U3666 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5388) );
  XNOR2_X1 U3667 ( .A(n4693), .B(n4691), .ZN(n4593) );
  NAND2_X1 U3668 ( .A1(n6138), .A2(n4497), .ZN(n6371) );
  AND3_X1 U3669 ( .A1(n6269), .A2(n6485), .A3(n6473), .ZN(n4497) );
  AND2_X1 U3670 ( .A1(n5174), .A2(n5307), .ZN(n5309) );
  NOR2_X1 U3671 ( .A1(n4619), .A2(n4563), .ZN(n5956) );
  AND2_X1 U3672 ( .A1(n5257), .A2(n5154), .ZN(n5100) );
  AND2_X1 U3673 ( .A1(n4500), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5112)
         );
  INV_X1 U3674 ( .A(n5140), .ZN(n4500) );
  NAND2_X1 U3675 ( .A1(n5112), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5153)
         );
  AND2_X1 U3676 ( .A1(n4474), .A2(n4473), .ZN(n5406) );
  OR2_X1 U3677 ( .A1(n6411), .A2(n5141), .ZN(n4473) );
  AOI21_X1 U3678 ( .B1(n4445), .B2(n4444), .A(n4443), .ZN(n5416) );
  AND2_X1 U3679 ( .A1(n6398), .A2(n5154), .ZN(n4443) );
  AND2_X1 U3680 ( .A1(n4426), .A2(n4425), .ZN(n5764) );
  CLKBUF_X1 U3681 ( .A(n5425), .Z(n5426) );
  NOR2_X1 U3682 ( .A1(n4373), .A2(n4372), .ZN(n4374) );
  INV_X1 U3683 ( .A(n6065), .ZN(n4391) );
  CLKBUF_X1 U3684 ( .A(n5319), .Z(n5320) );
  AND2_X1 U3685 ( .A1(n4350), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4351)
         );
  NAND2_X1 U3686 ( .A1(n4351), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4373)
         );
  CLKBUF_X1 U3687 ( .A(n5318), .Z(n5335) );
  CLKBUF_X1 U3688 ( .A(n5333), .Z(n5334) );
  NAND2_X1 U3689 ( .A1(n4305), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4322)
         );
  CLKBUF_X1 U3690 ( .A(n5349), .Z(n5350) );
  CLKBUF_X1 U3691 ( .A(n5361), .Z(n5438) );
  NOR2_X1 U3692 ( .A1(n4300), .A2(n5823), .ZN(n4305) );
  NAND2_X1 U3693 ( .A1(n4285), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4300)
         );
  AND2_X1 U3694 ( .A1(n4244), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4259)
         );
  AND3_X1 U3696 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .A3(n4193), .ZN(n4214) );
  AOI21_X1 U3697 ( .B1(n4190), .B2(n4314), .A(n4189), .ZN(n4657) );
  NOR2_X1 U3698 ( .A1(n4181), .A2(n6100), .ZN(n4193) );
  NAND2_X1 U3699 ( .A1(n4174), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4181)
         );
  NOR2_X1 U3700 ( .A1(n4162), .A2(n5388), .ZN(n4174) );
  INV_X1 U3701 ( .A(n4612), .ZN(n4169) );
  NAND2_X1 U3702 ( .A1(n4150), .A2(n4149), .ZN(n4560) );
  INV_X1 U3703 ( .A(n4619), .ZN(n4893) );
  BUF_X1 U3704 ( .A(n3799), .Z(n5293) );
  INV_X1 U3705 ( .A(n5709), .ZN(n4125) );
  NOR2_X2 U3706 ( .A1(n5411), .A2(n4504), .ZN(n5176) );
  CLKBUF_X1 U3707 ( .A(n5417), .Z(n5884) );
  NOR2_X2 U3708 ( .A1(n6069), .A2(n6070), .ZN(n6068) );
  AND2_X1 U3709 ( .A1(n4086), .A2(n4085), .ZN(n4087) );
  INV_X1 U3710 ( .A(n5811), .ZN(n4110) );
  AND2_X1 U3711 ( .A1(n3750), .A2(n3749), .ZN(n5366) );
  NOR2_X2 U3712 ( .A1(n5367), .A2(n5366), .ZN(n5441) );
  AND2_X1 U3713 ( .A1(n5692), .A2(n6179), .ZN(n5811) );
  OR2_X1 U3714 ( .A1(n5692), .A2(n6179), .ZN(n5810) );
  OR2_X1 U3715 ( .A1(n5692), .A2(n6250), .ZN(n4953) );
  INV_X1 U3716 ( .A(n4824), .ZN(n3729) );
  INV_X1 U3717 ( .A(n4811), .ZN(n3730) );
  INV_X1 U3718 ( .A(n6217), .ZN(n5901) );
  AND2_X1 U3719 ( .A1(n3713), .A2(n3712), .ZN(n4650) );
  OR2_X2 U3720 ( .A1(n3945), .A2(n3944), .ZN(n4693) );
  AND2_X1 U3721 ( .A1(n6641), .A2(n6640), .ZN(n6653) );
  BUF_X1 U3722 ( .A(n4702), .Z(n6566) );
  INV_X1 U3723 ( .A(n6723), .ZN(n6696) );
  NAND2_X1 U3724 ( .A1(n6544), .A2(n6543), .ZN(n7001) );
  AOI21_X1 U3725 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6709), .A(n6546), .ZN(
        n6685) );
  AND2_X1 U3726 ( .A1(n6475), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3942) );
  AND2_X1 U3727 ( .A1(n6467), .A2(n6466), .ZN(n6468) );
  INV_X1 U3728 ( .A(n6152), .ZN(n6138) );
  OR2_X1 U3729 ( .A1(n4618), .A2(n4546), .ZN(n6152) );
  INV_X1 U3730 ( .A(n6395), .ZN(n6412) );
  CLKBUF_X1 U3731 ( .A(n4799), .Z(n4800) );
  INV_X1 U3732 ( .A(n3868), .ZN(n3869) );
  INV_X1 U3733 ( .A(n6390), .ZN(n6418) );
  NAND2_X1 U3734 ( .A1(n4534), .A2(n4533), .ZN(n4536) );
  AND2_X1 U3735 ( .A1(n6075), .A2(n5170), .ZN(n6072) );
  INV_X1 U3736 ( .A(n6060), .ZN(n6071) );
  INV_X1 U3737 ( .A(n6075), .ZN(n5445) );
  NAND2_X1 U3738 ( .A1(n6075), .A2(n7000), .ZN(n6060) );
  OAI21_X1 U3739 ( .B1(n5290), .B2(n5281), .A(n5280), .ZN(n5454) );
  NAND2_X1 U3740 ( .A1(n6514), .A2(n5171), .ZN(n6516) );
  AND2_X1 U3741 ( .A1(n6514), .A2(n4667), .ZN(n6534) );
  INV_X1 U3742 ( .A(n6514), .ZN(n6536) );
  NOR2_X2 U3743 ( .A1(n6536), .A2(n3662), .ZN(n6533) );
  NAND2_X1 U3744 ( .A1(n4760), .A2(n4666), .ZN(n6514) );
  OAI21_X1 U3745 ( .B1(n4665), .B2(n4664), .A(n6461), .ZN(n4666) );
  INV_X1 U3746 ( .A(n6534), .ZN(n5678) );
  NAND2_X1 U3747 ( .A1(n6514), .A2(n4668), .ZN(n5677) );
  OR2_X1 U3748 ( .A1(n4620), .A2(n6750), .ZN(n4760) );
  NOR2_X1 U3749 ( .A1(n5105), .A2(n4501), .ZN(n4502) );
  AOI21_X1 U3750 ( .B1(n5268), .B2(n5280), .A(n5267), .ZN(n5698) );
  INV_X1 U3751 ( .A(n6123), .ZN(n6101) );
  OR2_X1 U3752 ( .A1(n5877), .A2(n3685), .ZN(n5857) );
  OR2_X1 U3753 ( .A1(n6164), .A2(n4121), .ZN(n5848) );
  AND2_X1 U3754 ( .A1(n3682), .A2(n3681), .ZN(n6158) );
  NAND2_X1 U3755 ( .A1(n6199), .A2(n5930), .ZN(n5905) );
  AOI21_X1 U3756 ( .B1(n4958), .B2(n5901), .A(n4961), .ZN(n6249) );
  INV_X1 U3757 ( .A(n6223), .ZN(n6281) );
  OR2_X1 U3758 ( .A1(n4636), .A2(n4637), .ZN(n6165) );
  INV_X1 U3759 ( .A(n6663), .ZN(n6640) );
  INV_X1 U3760 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6649) );
  CLKBUF_X1 U3761 ( .A(n4676), .Z(n4677) );
  AND2_X1 U3762 ( .A1(n4700), .A2(n6546), .ZN(n5953) );
  NOR2_X1 U3763 ( .A1(n5239), .A2(n6744), .ZN(n5205) );
  AND2_X2 U3764 ( .A1(n3468), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4591)
         );
  INV_X1 U3765 ( .A(n5948), .ZN(n6430) );
  OR2_X1 U3766 ( .A1(n6713), .A2(n6712), .ZN(n7100) );
  OAI211_X1 U3767 ( .C1(n6704), .C2(n7092), .A(n6703), .B(n6702), .ZN(n7095)
         );
  OAI211_X1 U3768 ( .C1(n7078), .C2(n6744), .A(n6678), .B(n6742), .ZN(n7081)
         );
  AND2_X1 U3769 ( .A1(n6653), .A2(n6696), .ZN(n7080) );
  OAI211_X1 U3770 ( .C1(n7050), .C2(n6744), .A(n6623), .B(n6622), .ZN(n7053)
         );
  OAI21_X1 U3771 ( .B1(n7038), .B2(n6744), .A(n6604), .ZN(n7040) );
  AND2_X1 U3772 ( .A1(n5804), .A2(DATAI_26_), .ZN(n6821) );
  AND2_X1 U3773 ( .A1(n5804), .A2(DATAI_30_), .ZN(n6989) );
  INV_X1 U3774 ( .A(n6662), .ZN(n6735) );
  INV_X1 U3775 ( .A(n6775), .ZN(n6785) );
  INV_X1 U3776 ( .A(n6814), .ZN(n6826) );
  INV_X1 U3777 ( .A(n6855), .ZN(n6867) );
  INV_X1 U3778 ( .A(n6896), .ZN(n6908) );
  OR2_X1 U3779 ( .A1(n6552), .A2(n6696), .ZN(n7115) );
  INV_X1 U3780 ( .A(n7010), .ZN(n7013) );
  INV_X1 U3781 ( .A(n6940), .ZN(n6950) );
  INV_X1 U3782 ( .A(n6981), .ZN(n6994) );
  INV_X1 U3783 ( .A(n7076), .ZN(n7109) );
  INV_X1 U3784 ( .A(n5205), .ZN(n6478) );
  INV_X1 U3785 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6475) );
  NAND2_X1 U3786 ( .A1(n3942), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6487) );
  NOR2_X1 U3787 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6469) );
  INV_X1 U3788 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6482) );
  INV_X1 U3789 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6744) );
  AND2_X1 U3790 ( .A1(STATE_REG_1__SCAN_IN), .A2(n6501), .ZN(n6512) );
  NOR2_X1 U3791 ( .A1(n4096), .A2(n4921), .ZN(n3454) );
  AND2_X2 U3792 ( .A1(n3479), .A2(n4591), .ZN(n3902) );
  NAND2_X2 U3793 ( .A1(n6831), .A2(n4564), .ZN(n3693) );
  AND2_X2 U3794 ( .A1(n3479), .A2(n3487), .ZN(n3951) );
  INV_X1 U3795 ( .A(n5141), .ZN(n5154) );
  NOR2_X2 U3796 ( .A1(n7005), .A2(n6540), .ZN(n6725) );
  INV_X1 U3797 ( .A(n5320), .ZN(n6066) );
  AND2_X2 U3798 ( .A1(n5407), .A2(n5406), .ZN(n3455) );
  OR2_X1 U3799 ( .A1(n6383), .A2(n5189), .ZN(n3456) );
  NAND2_X1 U3800 ( .A1(n5166), .A2(n4493), .ZN(n5188) );
  AND4_X1 U3801 ( .A1(n3529), .A2(n3528), .A3(n3527), .A4(n3526), .ZN(n3457)
         );
  AND4_X1 U3802 ( .A1(n3537), .A2(n3536), .A3(n3535), .A4(n3534), .ZN(n3458)
         );
  NAND2_X1 U3803 ( .A1(n5692), .A2(n4126), .ZN(n3459) );
  AND2_X1 U3804 ( .A1(n3616), .A2(n3816), .ZN(n3460) );
  INV_X1 U3805 ( .A(n4388), .ZN(n5221) );
  AND2_X2 U3806 ( .A1(n6424), .A2(n4897), .ZN(n6123) );
  AND2_X1 U3807 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3461) );
  INV_X1 U3808 ( .A(READY_N), .ZN(n6500) );
  OR2_X1 U3809 ( .A1(n5768), .A2(n5767), .ZN(n5766) );
  INV_X1 U3810 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3500) );
  AND4_X1 U3811 ( .A1(n3541), .A2(n3540), .A3(n3539), .A4(n3538), .ZN(n3462)
         );
  AND2_X1 U3812 ( .A1(n5692), .A2(n6261), .ZN(n3463) );
  INV_X1 U3813 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4694) );
  AND4_X1 U3814 ( .A1(n3533), .A2(n3532), .A3(n3531), .A4(n3530), .ZN(n3464)
         );
  OR2_X1 U3815 ( .A1(n5707), .A2(n6223), .ZN(n3465) );
  OR2_X1 U3816 ( .A1(n3848), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3466)
         );
  NAND2_X2 U3817 ( .A1(n4088), .A2(n4087), .ZN(n4095) );
  INV_X1 U3818 ( .A(n3852), .ZN(n3623) );
  AND2_X2 U3819 ( .A1(n3484), .A2(n4591), .ZN(n3952) );
  INV_X1 U3820 ( .A(keyinput_4), .ZN(n5464) );
  NAND2_X1 U3821 ( .A1(n5465), .A2(n5464), .ZN(n5466) );
  NOR3_X1 U3822 ( .A1(n5479), .A2(n5478), .A3(n5477), .ZN(n5480) );
  AOI211_X1 U3823 ( .C1(DATAI_17_), .C2(keyinput_14), .A(n5484), .B(n5483), 
        .ZN(n5485) );
  AOI21_X1 U3824 ( .B1(keyinput_23), .B2(DATAI_8_), .A(n5493), .ZN(n5494) );
  OAI22_X1 U3825 ( .A1(n5614), .A2(keyinput_31), .B1(n5505), .B2(DATAI_0_), 
        .ZN(n5506) );
  INV_X1 U3826 ( .A(n5506), .ZN(n5507) );
  OAI22_X1 U3827 ( .A1(n6503), .A2(keyinput_33), .B1(n5511), .B2(NA_N), .ZN(
        n5512) );
  INV_X1 U3828 ( .A(n5512), .ZN(n5513) );
  NAND2_X1 U3829 ( .A1(n5514), .A2(n5513), .ZN(n5515) );
  AOI22_X1 U3830 ( .A1(n5519), .A2(n5518), .B1(READREQUEST_REG_SCAN_IN), .B2(
        keyinput_37), .ZN(n5520) );
  AOI211_X1 U3831 ( .C1(n5529), .C2(n5528), .A(n5527), .B(n5526), .ZN(n5530)
         );
  AOI21_X1 U3832 ( .B1(keyinput_48), .B2(n6056), .A(n5536), .ZN(n5537) );
  AND2_X1 U3833 ( .A1(n3815), .A2(n3814), .ZN(n3828) );
  INV_X1 U3834 ( .A(n3964), .ZN(n3914) );
  AOI21_X1 U3835 ( .B1(keyinput_56), .B2(n6027), .A(n5546), .ZN(n5547) );
  OR2_X1 U3837 ( .A1(n3909), .A2(n3908), .ZN(n4089) );
  OR2_X1 U3838 ( .A1(n4013), .A2(n4012), .ZN(n4040) );
  OR2_X1 U3839 ( .A1(n3958), .A2(n3957), .ZN(n3995) );
  AND2_X1 U3840 ( .A1(n4564), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3553) );
  INV_X1 U3841 ( .A(n3644), .ZN(n3813) );
  NAND2_X1 U3842 ( .A1(n3499), .A2(n3498), .ZN(n3507) );
  OR2_X1 U3843 ( .A1(n4059), .A2(n4058), .ZN(n4077) );
  NAND2_X1 U3844 ( .A1(n4200), .A2(n4085), .ZN(n4081) );
  OR2_X1 U3845 ( .A1(n3887), .A2(n3886), .ZN(n3964) );
  NAND2_X1 U3846 ( .A1(n3616), .A2(n6914), .ZN(n3802) );
  AND4_X1 U3847 ( .A1(n3835), .A2(n3834), .A3(n3833), .A4(n3832), .ZN(n3836)
         );
  AOI22_X1 U3848 ( .A1(n3952), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4229), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U3849 ( .A1(n3895), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3858), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3593) );
  AND2_X1 U3850 ( .A1(n4499), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5136)
         );
  OR2_X1 U3851 ( .A1(n5153), .A2(n5151), .ZN(n5103) );
  NOR2_X1 U3852 ( .A1(n4470), .A2(n5760), .ZN(n4471) );
  INV_X1 U3853 ( .A(n5337), .ZN(n4354) );
  AND2_X1 U3854 ( .A1(n3777), .A2(n3776), .ZN(n5882) );
  AND2_X1 U3855 ( .A1(n3735), .A2(n3734), .ZN(n4859) );
  OR2_X1 U3856 ( .A1(n4032), .A2(n4031), .ZN(n4043) );
  NAND2_X1 U3857 ( .A1(n3970), .A2(n3700), .ZN(n6089) );
  AND2_X1 U3858 ( .A1(n3919), .A2(n3920), .ZN(n3917) );
  OR2_X1 U3859 ( .A1(n4131), .A2(n4564), .ZN(n3636) );
  NAND2_X1 U3860 ( .A1(n5269), .A2(n5012), .ZN(n4533) );
  OR2_X1 U3861 ( .A1(n5269), .A2(n4531), .ZN(n4534) );
  NAND2_X1 U3862 ( .A1(n5136), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5140)
         );
  AND2_X1 U3863 ( .A1(n4061), .A2(n4060), .ZN(n4064) );
  OAI21_X1 U3864 ( .B1(n4167), .B2(n3467), .A(n4147), .ZN(n4148) );
  INV_X1 U3865 ( .A(n6143), .ZN(n5242) );
  OR2_X1 U3866 ( .A1(n5103), .A2(n5272), .ZN(n5105) );
  NAND2_X1 U3867 ( .A1(n4471), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4498)
         );
  NOR2_X1 U3868 ( .A1(n5204), .A2(n6482), .ZN(n5149) );
  INV_X1 U3869 ( .A(n4154), .ZN(n4388) );
  AOI21_X1 U3870 ( .B1(n4200), .B2(n4314), .A(n4199), .ZN(n4815) );
  NAND2_X1 U3871 ( .A1(n3978), .A2(n3977), .ZN(n4691) );
  NAND2_X1 U3872 ( .A1(n3577), .A2(n3576), .ZN(n3578) );
  INV_X1 U3873 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6717) );
  AND2_X1 U3874 ( .A1(n3844), .A2(n6681), .ZN(n6677) );
  NAND2_X1 U3875 ( .A1(n3918), .A2(n3917), .ZN(n3924) );
  INV_X1 U3876 ( .A(n4495), .ZN(n5229) );
  INV_X1 U3877 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6350) );
  AND2_X1 U3878 ( .A1(n4259), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4285)
         );
  NAND2_X1 U3879 ( .A1(n6296), .A2(n4865), .ZN(n6340) );
  OR2_X1 U3880 ( .A1(n4835), .A2(n4511), .ZN(n5249) );
  AOI211_X1 U3881 ( .C1(n6374), .C2(keyinput_62), .A(n5554), .B(n5553), .ZN(
        n5555) );
  OAI21_X1 U3882 ( .B1(n6124), .B2(n4123), .A(n4122), .ZN(n5728) );
  INV_X1 U3883 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5823) );
  NAND2_X1 U3884 ( .A1(n4214), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4228)
         );
  NAND2_X1 U3885 ( .A1(n5443), .A2(n3760), .ZN(n5342) );
  INV_X1 U3886 ( .A(n6165), .ZN(n5917) );
  OR2_X1 U3887 ( .A1(n4614), .A2(n3715), .ZN(n4660) );
  CLKBUF_X1 U3888 ( .A(n4614), .Z(n4651) );
  INV_X1 U3889 ( .A(n3687), .ZN(n5241) );
  OR2_X1 U3890 ( .A1(n6666), .A2(n6665), .ZN(n6682) );
  AND2_X1 U3891 ( .A1(n3436), .A2(n6640), .ZN(n6694) );
  INV_X1 U3892 ( .A(n6692), .ZN(n6697) );
  INV_X1 U3893 ( .A(n4564), .ZN(n6545) );
  INV_X2 U3894 ( .A(n3637), .ZN(n6955) );
  OR2_X1 U3895 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n5141) );
  NOR2_X1 U3896 ( .A1(n4619), .A2(n5229), .ZN(n4618) );
  NAND2_X1 U3897 ( .A1(n6371), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4835) );
  INV_X1 U3898 ( .A(n6348), .ZN(n6360) );
  INV_X1 U3899 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4867) );
  AND2_X1 U3900 ( .A1(n6371), .A2(n4513), .ZN(n6397) );
  INV_X1 U3901 ( .A(n5249), .ZN(n6296) );
  XNOR2_X1 U3902 ( .A(n4536), .B(n4535), .ZN(n5243) );
  INV_X1 U3903 ( .A(n6487), .ZN(n6461) );
  INV_X1 U3904 ( .A(n5303), .ZN(n5306) );
  INV_X1 U3905 ( .A(n6516), .ZN(n6537) );
  INV_X1 U3906 ( .A(n4760), .ZN(n4728) );
  AOI21_X1 U3907 ( .B1(n5408), .B2(n5415), .A(n3455), .ZN(n6535) );
  NAND2_X1 U3908 ( .A1(n4374), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4422)
         );
  CLKBUF_X1 U3909 ( .A(n4918), .Z(n4999) );
  NAND2_X1 U3910 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4162) );
  INV_X1 U3911 ( .A(n5848), .ZN(n6276) );
  AND2_X1 U3912 ( .A1(n5766), .A2(n5739), .ZN(n5759) );
  AND2_X1 U3913 ( .A1(n3656), .A2(n6461), .ZN(n4141) );
  AND2_X1 U3914 ( .A1(n4141), .A2(n3805), .ZN(n6280) );
  INV_X1 U3915 ( .A(n7105), .ZN(n7111) );
  INV_X1 U3916 ( .A(n7098), .ZN(n7101) );
  NOR2_X1 U3917 ( .A1(n6682), .A2(n6723), .ZN(n7094) );
  NOR2_X1 U3918 ( .A1(n6682), .A2(n6696), .ZN(n7085) );
  AND2_X1 U3919 ( .A1(n6653), .A2(n6723), .ZN(n7072) );
  AND2_X1 U3920 ( .A1(n6626), .A2(n6696), .ZN(n7065) );
  NAND2_X1 U3921 ( .A1(n6666), .A2(n6694), .ZN(n6615) );
  INV_X1 U3922 ( .A(n6974), .ZN(n7052) );
  NOR2_X2 U3923 ( .A1(n6615), .A2(n6696), .ZN(n7044) );
  INV_X1 U3924 ( .A(n7031), .ZN(n7033) );
  AND2_X1 U3925 ( .A1(n6568), .A2(n6640), .ZN(n7027) );
  INV_X1 U3926 ( .A(n7017), .ZN(n7018) );
  INV_X1 U3927 ( .A(n7115), .ZN(n7006) );
  INV_X1 U3928 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6459) );
  AND2_X1 U3929 ( .A1(n5236), .A2(n4496), .ZN(n4546) );
  OR2_X1 U3930 ( .A1(n4835), .A2(n4506), .ZN(n6390) );
  INV_X1 U3931 ( .A(n6415), .ZN(n6383) );
  AND2_X1 U3932 ( .A1(n6391), .A2(n4826), .ZN(n6318) );
  AND2_X1 U3933 ( .A1(n4555), .A2(n6461), .ZN(n6075) );
  INV_X2 U3934 ( .A(n6072), .ZN(n6061) );
  INV_X1 U3935 ( .A(n5956), .ZN(n5987) );
  NAND2_X1 U3936 ( .A1(n4893), .A2(n6465), .ZN(n4735) );
  INV_X1 U3937 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6100) );
  NAND2_X2 U3938 ( .A1(n4893), .A2(n6448), .ZN(n6424) );
  AND2_X1 U3939 ( .A1(n3673), .A2(n3672), .ZN(n6164) );
  INV_X1 U3940 ( .A(n6277), .ZN(n6269) );
  NAND2_X1 U3941 ( .A1(n4141), .A2(n4140), .ZN(n6223) );
  INV_X1 U3942 ( .A(n6280), .ZN(n6227) );
  INV_X1 U3943 ( .A(n4800), .ZN(n6607) );
  INV_X1 U3944 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5218) );
  OR2_X1 U3945 ( .A1(n6724), .A2(n6723), .ZN(n7105) );
  OR2_X1 U3946 ( .A1(n6724), .A2(n6696), .ZN(n7098) );
  INV_X1 U3947 ( .A(n7094), .ZN(n7091) );
  INV_X1 U3948 ( .A(n7080), .ZN(n6984) );
  INV_X1 U3949 ( .A(n7072), .ZN(n7069) );
  INV_X1 U3950 ( .A(n7065), .ZN(n6936) );
  OR2_X1 U3951 ( .A1(n6615), .A2(n6723), .ZN(n6974) );
  INV_X1 U3952 ( .A(n6971), .ZN(n7061) );
  INV_X1 U3953 ( .A(n6609), .ZN(n7049) );
  AOI22_X1 U3954 ( .A1(n6603), .A2(n6600), .B1(n6598), .B2(n6597), .ZN(n7043)
         );
  OR2_X1 U3955 ( .A1(n6592), .A2(n6696), .ZN(n7031) );
  INV_X1 U3956 ( .A(n7027), .ZN(n7024) );
  NAND2_X1 U3957 ( .A1(n6560), .A2(n6640), .ZN(n7017) );
  INV_X1 U3958 ( .A(n6772), .ZN(n6789) );
  OR2_X1 U3959 ( .A1(n6552), .A2(n6723), .ZN(n7010) );
  INV_X1 U3960 ( .A(n6468), .ZN(n6477) );
  INV_X1 U3961 ( .A(n6036), .ZN(n6030) );
  OR2_X1 U3962 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6509), .ZN(n6038) );
  OR2_X1 U3963 ( .A1(n4521), .A2(n4520), .ZN(U2803) );
  INV_X1 U3964 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4143) );
  INV_X1 U3965 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3467) );
  NOR2_X2 U3966 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n3474), .ZN(n3479)
         );
  NAND2_X1 U3968 ( .A1(n3951), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3473) );
  INV_X1 U3969 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3468) );
  NAND2_X1 U3970 ( .A1(n3902), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3472)
         );
  INV_X1 U3971 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3469) );
  NOR2_X2 U3972 ( .A1(n3469), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3485)
         );
  NOR2_X4 U3973 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4690) );
  AND2_X2 U3974 ( .A1(n3485), .A2(n4690), .ZN(n3622) );
  NAND2_X1 U3975 ( .A1(n5037), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3471) );
  NAND2_X1 U3976 ( .A1(n3628), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3470)
         );
  NAND2_X1 U3978 ( .A1(n5036), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3478) );
  INV_X1 U3979 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3474) );
  AND2_X2 U3980 ( .A1(n3474), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3484)
         );
  AND2_X2 U3981 ( .A1(n3484), .A2(n3487), .ZN(n3903) );
  NAND2_X1 U3982 ( .A1(n3903), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3477) );
  AND2_X2 U3983 ( .A1(n4591), .A2(n4592), .ZN(n3858) );
  NAND2_X1 U3984 ( .A1(n3858), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3476)
         );
  AND2_X2 U3985 ( .A1(n4690), .A2(n4687), .ZN(n4273) );
  NAND2_X1 U3986 ( .A1(n4273), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3475)
         );
  NAND2_X1 U3987 ( .A1(n3895), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3483)
         );
  AND2_X2 U3988 ( .A1(n3484), .A2(n4687), .ZN(n3896) );
  NAND2_X1 U3989 ( .A1(n3896), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3482)
         );
  NAND2_X1 U3990 ( .A1(n3432), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3481) );
  NAND2_X1 U3991 ( .A1(n3590), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3480) );
  NAND2_X1 U3992 ( .A1(n3952), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3491) );
  NAND2_X1 U3993 ( .A1(n3450), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3490) );
  AND2_X2 U3994 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4602) );
  AND2_X2 U3995 ( .A1(n4602), .A2(n3486), .ZN(n3600) );
  NAND2_X1 U3996 ( .A1(n4427), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3489) );
  NAND2_X1 U3998 ( .A1(n4229), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3488) );
  AND4_X2 U3999 ( .A1(n3491), .A2(n3490), .A3(n3489), .A4(n3488), .ZN(n3492)
         );
  XNOR2_X1 U4000 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .ZN(
        n6499) );
  OR2_X1 U4001 ( .A1(n6499), .A2(STATE_REG_0__SCAN_IN), .ZN(n6143) );
  XNOR2_X1 U4002 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3509) );
  NAND2_X1 U4003 ( .A1(n6709), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3548) );
  NAND2_X1 U4004 ( .A1(n3509), .A2(n3508), .ZN(n3497) );
  NAND2_X1 U4005 ( .A1(n6717), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3496) );
  NAND2_X1 U4006 ( .A1(n3497), .A2(n3496), .ZN(n3511) );
  XNOR2_X1 U4007 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3510) );
  NAND2_X1 U4008 ( .A1(n3511), .A2(n3510), .ZN(n3499) );
  NAND2_X1 U4009 ( .A1(n6649), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3498) );
  MUX2_X1 U4010 ( .A(n3500), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n3506) );
  NAND2_X1 U4011 ( .A1(n3507), .A2(n3506), .ZN(n3502) );
  NAND2_X1 U4012 ( .A1(n3500), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3501) );
  NAND2_X1 U4013 ( .A1(n3502), .A2(n3501), .ZN(n3503) );
  NAND2_X1 U4014 ( .A1(n3513), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3505) );
  NAND2_X1 U4015 ( .A1(n3503), .A2(n6459), .ZN(n3504) );
  XNOR2_X1 U4016 ( .A(n3507), .B(n3506), .ZN(n3568) );
  XNOR2_X1 U4017 ( .A(n3509), .B(n3508), .ZN(n3543) );
  XNOR2_X1 U4018 ( .A(n3511), .B(n3510), .ZN(n3558) );
  NOR3_X1 U4019 ( .A1(n3568), .A2(n3543), .A3(n3558), .ZN(n3512) );
  OR2_X1 U4020 ( .A1(n3576), .A2(n3512), .ZN(n3515) );
  NAND2_X1 U4021 ( .A1(n3515), .A2(n3569), .ZN(n5235) );
  NAND2_X1 U4022 ( .A1(n6500), .A2(n5235), .ZN(n4583) );
  AOI21_X1 U4023 ( .B1(n4586), .B2(n6143), .A(n4583), .ZN(n3612) );
  AOI22_X1 U4024 ( .A1(n3895), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3858), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3519) );
  AOI22_X1 U4025 ( .A1(n3896), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3432), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3518) );
  AOI22_X1 U4026 ( .A1(n3902), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3590), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3517) );
  AOI22_X1 U4027 ( .A1(n3853), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3628), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3516) );
  NAND4_X1 U4028 ( .A1(n3519), .A2(n3518), .A3(n3517), .A4(n3516), .ZN(n3525)
         );
  AOI22_X1 U4029 ( .A1(n3431), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5037), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3523) );
  AOI22_X1 U4030 ( .A1(n3952), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4229), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3522) );
  AOI22_X1 U4031 ( .A1(n3903), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3521) );
  BUF_X4 U4032 ( .A(n3600), .Z(n4427) );
  AOI22_X1 U4033 ( .A1(n3449), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4427), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3520) );
  NAND4_X1 U4034 ( .A1(n3523), .A2(n3522), .A3(n3521), .A4(n3520), .ZN(n3524)
         );
  OR2_X4 U4035 ( .A1(n3525), .A2(n3524), .ZN(n4564) );
  AOI22_X1 U4036 ( .A1(n3903), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3858), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3529) );
  AOI22_X1 U4037 ( .A1(n3952), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3622), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3528) );
  AOI22_X1 U4038 ( .A1(n3852), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4229), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3527) );
  AOI22_X1 U4039 ( .A1(n5036), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3526) );
  AOI22_X1 U4040 ( .A1(n3896), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3533) );
  AOI22_X1 U4041 ( .A1(n3902), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3590), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3532) );
  AOI22_X1 U4042 ( .A1(n3895), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3600), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3531) );
  AOI22_X1 U4043 ( .A1(n3951), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3628), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3530) );
  NAND2_X2 U4044 ( .A1(n3457), .A2(n3464), .ZN(n4136) );
  AOI22_X1 U4045 ( .A1(n3895), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3902), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4046 ( .A1(n3951), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3858), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3536) );
  AOI22_X1 U4047 ( .A1(n5036), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3600), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3535) );
  AOI22_X1 U4048 ( .A1(n3903), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4229), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3534) );
  AOI22_X1 U4049 ( .A1(n3852), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4050 ( .A1(n3622), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3590), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4051 ( .A1(n3432), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3628), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3538) );
  NAND2_X2 U4052 ( .A1(n3458), .A2(n3462), .ZN(n3621) );
  INV_X1 U4053 ( .A(n4072), .ZN(n3566) );
  INV_X1 U4054 ( .A(n4136), .ZN(n3642) );
  INV_X1 U4055 ( .A(n4071), .ZN(n3549) );
  INV_X2 U4056 ( .A(n3668), .ZN(n6750) );
  AND2_X1 U4057 ( .A1(n6750), .A2(n3889), .ZN(n3542) );
  NOR2_X2 U4058 ( .A1(n4564), .A2(n4586), .ZN(n5240) );
  OR2_X1 U4059 ( .A1(n3543), .A2(n6482), .ZN(n3550) );
  INV_X1 U4060 ( .A(n3550), .ZN(n3547) );
  NAND2_X1 U4061 ( .A1(n4071), .A2(n4586), .ZN(n3545) );
  NAND2_X1 U4062 ( .A1(n4072), .A2(n3543), .ZN(n3544) );
  AND3_X1 U4063 ( .A1(n3545), .A2(n3544), .A3(n3889), .ZN(n3551) );
  INV_X1 U4064 ( .A(n3551), .ZN(n3546) );
  OAI21_X1 U4065 ( .B1(n3577), .B2(n3547), .A(n3546), .ZN(n3561) );
  OAI21_X1 U4066 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6709), .A(n3548), 
        .ZN(n3552) );
  AOI211_X1 U4067 ( .C1(n3551), .C2(n3550), .A(n3552), .B(n3549), .ZN(n3557)
         );
  INV_X1 U4068 ( .A(n3552), .ZN(n3555) );
  INV_X1 U4069 ( .A(n3553), .ZN(n3554) );
  AOI21_X1 U4070 ( .B1(n3555), .B2(n4131), .A(n3554), .ZN(n3556) );
  OAI22_X1 U4071 ( .A1(n3557), .A2(n3577), .B1(n3556), .B2(n3563), .ZN(n3560)
         );
  AOI211_X1 U4072 ( .C1(n4072), .C2(n3558), .A(n3563), .B(n3564), .ZN(n3559)
         );
  AOI21_X1 U4073 ( .B1(n3561), .B2(n3560), .A(n3559), .ZN(n3562) );
  AOI21_X1 U4074 ( .B1(n3564), .B2(n3563), .A(n3562), .ZN(n3565) );
  AOI21_X1 U4075 ( .B1(n3566), .B2(n3568), .A(n3565), .ZN(n3567) );
  AOI21_X1 U4076 ( .B1(n3568), .B2(n3577), .A(n3567), .ZN(n3572) );
  NOR2_X1 U4077 ( .A1(n4072), .A2(n3569), .ZN(n3571) );
  INV_X1 U4078 ( .A(n3577), .ZN(n3570) );
  OAI22_X1 U4079 ( .A1(n3572), .A2(n3571), .B1(n3570), .B2(n3569), .ZN(n3573)
         );
  AOI21_X1 U4080 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6482), .A(n3573), 
        .ZN(n3575) );
  NAND2_X1 U4081 ( .A1(n4071), .A2(n3576), .ZN(n3574) );
  NAND2_X1 U4082 ( .A1(n3575), .A2(n3574), .ZN(n3579) );
  AOI22_X1 U4083 ( .A1(n3858), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3622), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3583) );
  AOI22_X1 U4084 ( .A1(n3897), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3582) );
  AOI22_X1 U4085 ( .A1(n3952), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3600), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U4086 ( .A1(n3903), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3628), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4087 ( .A1(n3450), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3896), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4088 ( .A1(n3895), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4229), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3585) );
  AOI22_X1 U4089 ( .A1(n3951), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3902), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3584) );
  AOI22_X1 U4090 ( .A1(n5036), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3590), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3587) );
  NAND3_X2 U4091 ( .A1(n3589), .A2(n3588), .A3(n3587), .ZN(n3643) );
  AOI22_X1 U4092 ( .A1(n3896), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3432), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3594) );
  AOI22_X1 U4093 ( .A1(n3902), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3590), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3592) );
  AOI22_X1 U4094 ( .A1(n3951), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3628), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4095 ( .A1(n3903), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4096 ( .A1(n3431), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3622), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4097 ( .A1(n3449), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3600), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3595) );
  AND2_X2 U4098 ( .A1(n3643), .A2(n3637), .ZN(n3616) );
  INV_X1 U4099 ( .A(n3616), .ZN(n3662) );
  NOR2_X1 U4100 ( .A1(n3616), .A2(n6545), .ZN(n3599) );
  NOR2_X1 U4101 ( .A1(n5239), .A2(n3599), .ZN(n3611) );
  AOI22_X1 U4102 ( .A1(n5036), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3622), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3604) );
  AOI22_X1 U4103 ( .A1(n3952), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4229), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3603) );
  AOI22_X1 U4104 ( .A1(n3903), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3602) );
  BUF_X2 U4105 ( .A(n3600), .Z(n5056) );
  AOI22_X1 U4106 ( .A1(n3852), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n5056), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3601) );
  NAND4_X1 U4107 ( .A1(n3604), .A2(n3603), .A3(n3602), .A4(n3601), .ZN(n3610)
         );
  AOI22_X1 U4108 ( .A1(n3895), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3858), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3608) );
  AOI22_X1 U4109 ( .A1(n3896), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3607) );
  AOI22_X1 U4110 ( .A1(n3902), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3590), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3606) );
  AOI22_X1 U4111 ( .A1(n3951), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3628), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3605) );
  NAND4_X1 U4112 ( .A1(n3608), .A2(n3607), .A3(n3606), .A4(n3605), .ZN(n3609)
         );
  OR2_X2 U4113 ( .A1(n3610), .A2(n3609), .ZN(n3816) );
  MUX2_X1 U4114 ( .A(n3612), .B(n3611), .S(n6790), .Z(n3613) );
  INV_X1 U4115 ( .A(n3613), .ZN(n3655) );
  AND2_X1 U4116 ( .A1(n4136), .A2(n3643), .ZN(n3614) );
  NAND2_X1 U4117 ( .A1(n3830), .A2(n3889), .ZN(n5204) );
  NOR2_X1 U4118 ( .A1(n5204), .A2(n6750), .ZN(n3648) );
  INV_X1 U4119 ( .A(n4131), .ZN(n3615) );
  NAND2_X1 U4120 ( .A1(n3615), .A2(n3460), .ZN(n3620) );
  INV_X2 U4121 ( .A(n3621), .ZN(n6914) );
  NAND2_X1 U4122 ( .A1(n3617), .A2(n3802), .ZN(n3618) );
  INV_X2 U4123 ( .A(n3816), .ZN(n6790) );
  NAND2_X1 U4124 ( .A1(n3618), .A2(n6790), .ZN(n3619) );
  NAND2_X1 U4125 ( .A1(n3620), .A2(n3619), .ZN(n3635) );
  AOI22_X1 U4126 ( .A1(n5036), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3622), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3627) );
  AOI22_X1 U4127 ( .A1(n3952), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4229), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4128 ( .A1(n3903), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4129 ( .A1(n3450), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5056), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3624) );
  NAND4_X1 U4130 ( .A1(n3627), .A2(n3626), .A3(n3625), .A4(n3624), .ZN(n3634)
         );
  AOI22_X1 U4131 ( .A1(n3895), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3858), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3632) );
  AOI22_X1 U4132 ( .A1(n3896), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3631) );
  AOI22_X1 U4133 ( .A1(n3902), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3590), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4134 ( .A1(n3951), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3628), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3629) );
  NAND4_X1 U4135 ( .A1(n3632), .A2(n3631), .A3(n3630), .A4(n3629), .ZN(n3633)
         );
  NAND2_X1 U4136 ( .A1(n3813), .A2(n3925), .ZN(n3831) );
  NAND2_X1 U4137 ( .A1(n3635), .A2(n3831), .ZN(n3812) );
  NOR2_X2 U4138 ( .A1(n3812), .A2(n3636), .ZN(n3840) );
  NAND2_X1 U4139 ( .A1(n3644), .A2(n6872), .ZN(n3640) );
  CLKBUF_X3 U4140 ( .A(n3643), .Z(n5170) );
  AND2_X1 U4141 ( .A1(n5170), .A2(n3925), .ZN(n3638) );
  AND2_X1 U4142 ( .A1(n3638), .A2(n4551), .ZN(n3639) );
  NAND2_X1 U4143 ( .A1(n5204), .A2(n6545), .ZN(n3641) );
  NAND3_X1 U4144 ( .A1(n3815), .A2(n3641), .A3(n6790), .ZN(n4132) );
  INV_X1 U4145 ( .A(n4132), .ZN(n4133) );
  NAND2_X1 U4146 ( .A1(n3817), .A2(n4668), .ZN(n3650) );
  AOI21_X1 U4147 ( .B1(n3644), .B2(n4586), .A(n6545), .ZN(n3645) );
  NAND2_X1 U4148 ( .A1(n3650), .A2(n3645), .ZN(n3665) );
  AND2_X1 U4149 ( .A1(n4133), .A2(n3665), .ZN(n3646) );
  INV_X1 U4150 ( .A(n3670), .ZN(n3647) );
  AOI21_X1 U4151 ( .B1(n5239), .B2(n3648), .A(n3647), .ZN(n4588) );
  OAI21_X1 U4152 ( .B1(n4586), .B2(n5242), .A(n6500), .ZN(n3649) );
  NOR2_X1 U4153 ( .A1(n5239), .A2(n3649), .ZN(n4582) );
  INV_X1 U4154 ( .A(n3650), .ZN(n3653) );
  NAND2_X1 U4155 ( .A1(n6790), .A2(n3925), .ZN(n3888) );
  NOR2_X1 U4156 ( .A1(n3888), .A2(n3651), .ZN(n3652) );
  NAND2_X1 U4157 ( .A1(n3653), .A2(n3652), .ZN(n3838) );
  INV_X1 U4158 ( .A(n4597), .ZN(n4579) );
  NAND2_X1 U4159 ( .A1(n4582), .A2(n4579), .ZN(n3654) );
  NAND3_X1 U4160 ( .A1(n3655), .A2(n4588), .A3(n3654), .ZN(n3656) );
  AND2_X1 U4161 ( .A1(n5236), .A2(n4586), .ZN(n5207) );
  NAND2_X1 U4162 ( .A1(n4141), .A2(n5207), .ZN(n3678) );
  INV_X1 U4163 ( .A(n3812), .ZN(n3658) );
  NAND2_X1 U4164 ( .A1(n4131), .A2(n4586), .ZN(n3657) );
  NAND2_X1 U4165 ( .A1(n3658), .A2(n3657), .ZN(n3659) );
  NAND2_X1 U4166 ( .A1(n3660), .A2(n3659), .ZN(n3837) );
  INV_X1 U4167 ( .A(n3815), .ZN(n3661) );
  INV_X4 U4168 ( .A(n3820), .ZN(n4531) );
  NAND2_X1 U4169 ( .A1(n3661), .A2(n4531), .ZN(n3664) );
  INV_X1 U4170 ( .A(n3925), .ZN(n6831) );
  NAND2_X1 U4171 ( .A1(n3662), .A2(n3888), .ZN(n3663) );
  AND4_X1 U4172 ( .A1(n3665), .A2(n3664), .A3(n3693), .A4(n3663), .ZN(n3666)
         );
  NAND2_X1 U4173 ( .A1(n3837), .A2(n3666), .ZN(n4594) );
  NAND2_X1 U4174 ( .A1(n4141), .A2(n4594), .ZN(n3677) );
  INV_X1 U4175 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U4176 ( .A1(n5940), .A2(n3678), .ZN(n5930) );
  INV_X1 U4177 ( .A(n5905), .ZN(n6181) );
  AND2_X1 U4178 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4115) );
  INV_X1 U4179 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3716) );
  INV_X1 U4180 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4852) );
  NOR2_X1 U4181 ( .A1(n4852), .A2(n4001), .ZN(n4851) );
  NAND2_X1 U4182 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4851), .ZN(n4792)
         );
  NOR2_X1 U4183 ( .A1(n3716), .A2(n4792), .ZN(n3671) );
  NAND3_X1 U4184 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n3671), .ZN(n6198) );
  NAND2_X1 U4185 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6232) );
  NOR2_X1 U4186 ( .A1(n6198), .A2(n6232), .ZN(n6219) );
  NAND3_X1 U4187 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n6219), .ZN(n4960) );
  INV_X1 U4188 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6179) );
  NAND3_X1 U4189 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n6174) );
  NOR2_X1 U4190 ( .A1(n6179), .A2(n6174), .ZN(n5916) );
  NAND3_X1 U4191 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n5916), .ZN(n5907) );
  NOR2_X1 U4192 ( .A1(n4960), .A2(n5907), .ZN(n5904) );
  NAND2_X1 U4193 ( .A1(n4115), .A2(n5904), .ZN(n3676) );
  INV_X1 U4194 ( .A(n3676), .ZN(n3667) );
  NAND2_X1 U4195 ( .A1(n6181), .A2(n3667), .ZN(n3673) );
  NAND2_X2 U4196 ( .A1(n4564), .A2(n3668), .ZN(n3687) );
  NOR2_X1 U4197 ( .A1(n5204), .A2(n3687), .ZN(n3669) );
  NAND2_X1 U4198 ( .A1(n3670), .A2(n3669), .ZN(n5228) );
  INV_X1 U4199 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5929) );
  OAI21_X1 U4200 ( .B1(n5929), .B2(n5940), .A(n3700), .ZN(n6183) );
  NAND2_X1 U4201 ( .A1(n3671), .A2(n6183), .ZN(n6195) );
  NOR2_X1 U4202 ( .A1(n6232), .A2(n6195), .ZN(n6218) );
  NAND3_X1 U4203 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n6218), .ZN(n4957) );
  NOR2_X1 U4204 ( .A1(n5907), .A2(n4957), .ZN(n5900) );
  NAND2_X1 U4205 ( .A1(n4115), .A2(n5900), .ZN(n3679) );
  OR2_X1 U4206 ( .A1(n6217), .A2(n3679), .ZN(n3672) );
  AND2_X1 U4207 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5893) );
  INV_X1 U4208 ( .A(n5893), .ZN(n3674) );
  NOR2_X1 U4209 ( .A1(n6164), .A2(n3674), .ZN(n5887) );
  AND2_X1 U4210 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5866) );
  INV_X1 U4211 ( .A(n5866), .ZN(n3675) );
  NAND2_X1 U4212 ( .A1(n5887), .A2(n3675), .ZN(n5872) );
  NOR2_X2 U4213 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6659) );
  AND2_X1 U4214 ( .A1(n6659), .A2(n6475), .ZN(n6137) );
  OAI22_X1 U4215 ( .A1(n3677), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .B1(n6277), 
        .B2(n4141), .ZN(n6222) );
  AOI21_X1 U4216 ( .B1(n6199), .B2(n3676), .A(n6222), .ZN(n3681) );
  NAND2_X1 U4217 ( .A1(n6217), .A2(n3677), .ZN(n4636) );
  INV_X1 U4218 ( .A(n3678), .ZN(n4637) );
  NAND2_X1 U4219 ( .A1(n3681), .A2(n5917), .ZN(n3684) );
  INV_X1 U4220 ( .A(n3679), .ZN(n3680) );
  OR2_X1 U4221 ( .A1(n6217), .A2(n3680), .ZN(n3682) );
  NAND2_X1 U4222 ( .A1(n6158), .A2(n5893), .ZN(n3683) );
  NAND2_X1 U4223 ( .A1(n3684), .A2(n3683), .ZN(n5891) );
  NAND2_X1 U4224 ( .A1(n5872), .A2(n5891), .ZN(n5877) );
  AND2_X1 U4225 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3806) );
  AOI21_X1 U4226 ( .B1(n6217), .B2(n5905), .A(n3806), .ZN(n3685) );
  NAND2_X1 U4227 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5852) );
  AND2_X1 U4228 ( .A1(n6165), .A2(n5852), .ZN(n3686) );
  NOR2_X1 U4229 ( .A1(n5857), .A2(n3686), .ZN(n5839) );
  INV_X1 U4230 ( .A(n3687), .ZN(n3706) );
  INV_X1 U4231 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3690) );
  NAND2_X1 U4232 ( .A1(n3706), .A2(n3690), .ZN(n3689) );
  NAND2_X1 U4233 ( .A1(n3452), .A2(n5929), .ZN(n3688) );
  NAND3_X1 U4234 ( .A1(n3689), .A2(n3820), .A3(n3688), .ZN(n3692) );
  NAND2_X1 U4235 ( .A1(n4531), .A2(n3690), .ZN(n3691) );
  NAND2_X1 U4236 ( .A1(n3692), .A2(n3691), .ZN(n3698) );
  NAND2_X1 U4237 ( .A1(n3453), .A2(EBX_REG_0__SCAN_IN), .ZN(n3696) );
  INV_X1 U4238 ( .A(EBX_REG_0__SCAN_IN), .ZN(n3694) );
  NAND2_X1 U4239 ( .A1(n3820), .A2(n3694), .ZN(n3695) );
  NAND2_X1 U4240 ( .A1(n3696), .A2(n3695), .ZN(n4548) );
  INV_X1 U4241 ( .A(n4548), .ZN(n3697) );
  NOR2_X1 U4242 ( .A1(n3698), .A2(n3697), .ZN(n3699) );
  AOI21_X2 U4243 ( .B1(n4827), .B2(n5241), .A(n3699), .ZN(n5193) );
  INV_X1 U4244 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3700) );
  NAND2_X1 U4245 ( .A1(n3693), .A2(n3700), .ZN(n3702) );
  INV_X1 U4246 ( .A(EBX_REG_2__SCAN_IN), .ZN(n3703) );
  NAND2_X1 U4247 ( .A1(n5241), .A2(n3703), .ZN(n3701) );
  NAND3_X1 U4248 ( .A1(n3702), .A2(n3451), .A3(n3701), .ZN(n3705) );
  NAND2_X1 U4249 ( .A1(n4531), .A2(n3703), .ZN(n3704) );
  NAND2_X1 U4250 ( .A1(n3705), .A2(n3704), .ZN(n5192) );
  NAND2_X2 U4251 ( .A1(n3693), .A2(n3451), .ZN(n4547) );
  NAND2_X2 U4252 ( .A1(n3706), .A2(n3451), .ZN(n3793) );
  MUX2_X1 U4253 ( .A(n3793), .B(n3451), .S(EBX_REG_3__SCAN_IN), .Z(n3707) );
  OAI21_X1 U4254 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n4547), .A(n3707), 
        .ZN(n3708) );
  INV_X1 U4255 ( .A(n3708), .ZN(n4615) );
  NAND2_X1 U4256 ( .A1(n5195), .A2(n4615), .ZN(n4614) );
  NAND2_X1 U4257 ( .A1(n3693), .A2(n4852), .ZN(n3710) );
  INV_X1 U4258 ( .A(EBX_REG_4__SCAN_IN), .ZN(n3711) );
  NAND2_X1 U4259 ( .A1(n5241), .A2(n3711), .ZN(n3709) );
  NAND3_X1 U4260 ( .A1(n3710), .A2(n3451), .A3(n3709), .ZN(n3713) );
  NAND2_X1 U4261 ( .A1(n4531), .A2(n3711), .ZN(n3712) );
  MUX2_X1 U4262 ( .A(n3793), .B(n3451), .S(EBX_REG_5__SCAN_IN), .Z(n3714) );
  OAI21_X1 U4263 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4547), .A(n3714), 
        .ZN(n4649) );
  NAND2_X1 U4264 ( .A1(n3693), .A2(n3716), .ZN(n3718) );
  INV_X1 U4265 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6324) );
  NAND2_X1 U4266 ( .A1(n5241), .A2(n6324), .ZN(n3717) );
  NAND3_X1 U4267 ( .A1(n3718), .A2(n3451), .A3(n3717), .ZN(n3720) );
  NAND2_X1 U4268 ( .A1(n4531), .A2(n6324), .ZN(n3719) );
  AND2_X1 U4269 ( .A1(n3720), .A2(n3719), .ZN(n4659) );
  NOR2_X2 U4270 ( .A1(n4660), .A2(n4659), .ZN(n4840) );
  MUX2_X1 U4271 ( .A(n3793), .B(n3451), .S(EBX_REG_7__SCAN_IN), .Z(n3721) );
  OAI21_X1 U4272 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n4547), .A(n3721), 
        .ZN(n3722) );
  INV_X1 U4273 ( .A(n3722), .ZN(n4839) );
  INV_X1 U4274 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U4275 ( .A1(n3693), .A2(n6209), .ZN(n3724) );
  INV_X1 U4276 ( .A(EBX_REG_8__SCAN_IN), .ZN(n3725) );
  NAND2_X1 U4277 ( .A1(n5241), .A2(n3725), .ZN(n3723) );
  NAND3_X1 U4278 ( .A1(n3724), .A2(n3451), .A3(n3723), .ZN(n3727) );
  NAND2_X1 U4279 ( .A1(n4531), .A2(n3725), .ZN(n3726) );
  NAND2_X1 U4280 ( .A1(n3727), .A2(n3726), .ZN(n4812) );
  NAND2_X1 U4281 ( .A1(n4842), .A2(n4812), .ZN(n4811) );
  MUX2_X1 U4282 ( .A(n3793), .B(n3451), .S(EBX_REG_9__SCAN_IN), .Z(n3728) );
  OAI21_X1 U4283 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n4547), .A(n3728), 
        .ZN(n4824) );
  NAND2_X1 U4284 ( .A1(n3693), .A2(n4100), .ZN(n3732) );
  INV_X1 U4285 ( .A(EBX_REG_10__SCAN_IN), .ZN(n3733) );
  NAND2_X1 U4286 ( .A1(n5241), .A2(n3733), .ZN(n3731) );
  NAND3_X1 U4287 ( .A1(n3732), .A2(n3451), .A3(n3731), .ZN(n3735) );
  NAND2_X1 U4288 ( .A1(n4531), .A2(n3733), .ZN(n3734) );
  MUX2_X1 U4289 ( .A(n3793), .B(n3451), .S(EBX_REG_11__SCAN_IN), .Z(n3736) );
  OAI21_X1 U4290 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n4547), .A(n3736), 
        .ZN(n4882) );
  INV_X1 U4291 ( .A(n4882), .ZN(n3737) );
  NAND2_X1 U4292 ( .A1(n4879), .A2(n3737), .ZN(n4909) );
  NAND2_X1 U4293 ( .A1(n3451), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3738) );
  NAND2_X1 U4294 ( .A1(n3693), .A2(n3738), .ZN(n3741) );
  INV_X1 U4295 ( .A(EBX_REG_12__SCAN_IN), .ZN(n3739) );
  NAND2_X1 U4296 ( .A1(n5241), .A2(n3739), .ZN(n3740) );
  AOI22_X1 U4297 ( .A1(n3741), .A2(n3740), .B1(n4531), .B2(n3739), .ZN(n4908)
         );
  INV_X1 U4298 ( .A(n3742), .ZN(n4979) );
  MUX2_X1 U4299 ( .A(n3793), .B(n3451), .S(EBX_REG_13__SCAN_IN), .Z(n3745) );
  INV_X1 U4300 ( .A(n4547), .ZN(n3743) );
  INV_X1 U4301 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U4302 ( .A1(n3743), .A2(n6173), .ZN(n3744) );
  NAND2_X1 U4303 ( .A1(n3745), .A2(n3744), .ZN(n4980) );
  OR2_X2 U4304 ( .A1(n4979), .A2(n4980), .ZN(n5367) );
  NAND2_X1 U4305 ( .A1(n3693), .A2(n6179), .ZN(n3747) );
  INV_X1 U4306 ( .A(EBX_REG_14__SCAN_IN), .ZN(n3748) );
  NAND2_X1 U4307 ( .A1(n5241), .A2(n3748), .ZN(n3746) );
  NAND3_X1 U4308 ( .A1(n3747), .A2(n3820), .A3(n3746), .ZN(n3750) );
  NAND2_X1 U4309 ( .A1(n4531), .A2(n3748), .ZN(n3749) );
  MUX2_X1 U4310 ( .A(n3793), .B(n3451), .S(EBX_REG_15__SCAN_IN), .Z(n3751) );
  OAI21_X1 U4311 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n4547), .A(n3751), 
        .ZN(n3752) );
  INV_X1 U4312 ( .A(n3752), .ZN(n5440) );
  AND2_X2 U4313 ( .A1(n5441), .A2(n5440), .ZN(n5443) );
  MUX2_X1 U4314 ( .A(n3793), .B(n3451), .S(EBX_REG_17__SCAN_IN), .Z(n3754) );
  OR2_X1 U4315 ( .A1(n4547), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3753)
         );
  NAND2_X1 U4316 ( .A1(n3754), .A2(n3753), .ZN(n5340) );
  INV_X1 U4317 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6262) );
  NAND2_X1 U4318 ( .A1(n3693), .A2(n6262), .ZN(n3756) );
  INV_X1 U4319 ( .A(EBX_REG_16__SCAN_IN), .ZN(n3757) );
  NAND2_X1 U4320 ( .A1(n5241), .A2(n3757), .ZN(n3755) );
  NAND3_X1 U4321 ( .A1(n3756), .A2(n3451), .A3(n3755), .ZN(n3759) );
  NAND2_X1 U4322 ( .A1(n4531), .A2(n3757), .ZN(n3758) );
  AND2_X1 U4323 ( .A1(n3759), .A2(n3758), .ZN(n5339) );
  NOR2_X1 U4324 ( .A1(n5340), .A2(n5339), .ZN(n3760) );
  INV_X1 U4325 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U4326 ( .A1(n3693), .A2(n5908), .ZN(n3762) );
  INV_X1 U4327 ( .A(EBX_REG_18__SCAN_IN), .ZN(n3763) );
  NAND2_X1 U4328 ( .A1(n5241), .A2(n3763), .ZN(n3761) );
  NAND3_X1 U4329 ( .A1(n3762), .A2(n3451), .A3(n3761), .ZN(n3765) );
  NAND2_X1 U4330 ( .A1(n4531), .A2(n3763), .ZN(n3764) );
  AND2_X1 U4331 ( .A1(n3765), .A2(n3764), .ZN(n5322) );
  OR2_X2 U4332 ( .A1(n5342), .A2(n5322), .ZN(n6069) );
  NAND2_X1 U4333 ( .A1(n3451), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3766) );
  OAI211_X1 U4334 ( .C1(n3687), .C2(EBX_REG_19__SCAN_IN), .A(n3693), .B(n3766), 
        .ZN(n3767) );
  OAI21_X1 U4335 ( .B1(n3793), .B2(EBX_REG_19__SCAN_IN), .A(n3767), .ZN(n6070)
         );
  NAND2_X1 U4336 ( .A1(n3451), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3768) );
  NAND2_X1 U4337 ( .A1(n3693), .A2(n3768), .ZN(n3770) );
  INV_X1 U4338 ( .A(EBX_REG_20__SCAN_IN), .ZN(n3771) );
  NAND2_X1 U4339 ( .A1(n5241), .A2(n3771), .ZN(n3769) );
  NAND2_X1 U4340 ( .A1(n3770), .A2(n3769), .ZN(n3773) );
  NAND2_X1 U4341 ( .A1(n4531), .A2(n3771), .ZN(n3772) );
  NAND2_X1 U4342 ( .A1(n3773), .A2(n3772), .ZN(n5423) );
  INV_X1 U4343 ( .A(n3793), .ZN(n3774) );
  INV_X1 U4344 ( .A(EBX_REG_21__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U4345 ( .A1(n3774), .A2(n6064), .ZN(n3777) );
  NAND2_X1 U4346 ( .A1(n3451), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3775) );
  OAI211_X1 U4347 ( .C1(n3687), .C2(EBX_REG_21__SCAN_IN), .A(n3693), .B(n3775), 
        .ZN(n3776) );
  NAND2_X1 U4348 ( .A1(n5422), .A2(n5882), .ZN(n5417) );
  INV_X1 U4349 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5757) );
  NAND2_X1 U4350 ( .A1(n3693), .A2(n5757), .ZN(n3779) );
  INV_X1 U4351 ( .A(EBX_REG_22__SCAN_IN), .ZN(n3780) );
  NAND2_X1 U4352 ( .A1(n5241), .A2(n3780), .ZN(n3778) );
  NAND3_X1 U4353 ( .A1(n3779), .A2(n3451), .A3(n3778), .ZN(n3782) );
  NAND2_X1 U4354 ( .A1(n4531), .A2(n3780), .ZN(n3781) );
  AND2_X1 U4355 ( .A1(n3782), .A2(n3781), .ZN(n5418) );
  OR2_X2 U4356 ( .A1(n5417), .A2(n5418), .ZN(n5420) );
  MUX2_X1 U4357 ( .A(n3793), .B(n3451), .S(EBX_REG_23__SCAN_IN), .Z(n3783) );
  OAI21_X1 U4358 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n4547), .A(n3783), 
        .ZN(n5409) );
  OR2_X2 U4359 ( .A1(n5420), .A2(n5409), .ZN(n5411) );
  INV_X1 U4360 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U4361 ( .A1(n3693), .A2(n5859), .ZN(n3785) );
  INV_X1 U4362 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5189) );
  NAND2_X1 U4363 ( .A1(n5241), .A2(n5189), .ZN(n3784) );
  NAND3_X1 U4364 ( .A1(n3785), .A2(n3451), .A3(n3784), .ZN(n3787) );
  NAND2_X1 U4365 ( .A1(n4531), .A2(n5189), .ZN(n3786) );
  AND2_X1 U4366 ( .A1(n3787), .A2(n3786), .ZN(n4504) );
  MUX2_X1 U4367 ( .A(n3793), .B(n3820), .S(EBX_REG_25__SCAN_IN), .Z(n3788) );
  OAI21_X1 U4368 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n4547), .A(n3788), 
        .ZN(n3789) );
  INV_X1 U4369 ( .A(n3789), .ZN(n5175) );
  INV_X1 U4370 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U4371 ( .A1(n3693), .A2(n5708), .ZN(n3790) );
  OAI211_X1 U4372 ( .C1(EBX_REG_26__SCAN_IN), .C2(n3687), .A(n3790), .B(n3451), 
        .ZN(n3792) );
  INV_X1 U4373 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U4374 ( .A1(n4531), .A2(n5405), .ZN(n3791) );
  NAND2_X1 U4375 ( .A1(n3792), .A2(n3791), .ZN(n5307) );
  MUX2_X1 U4376 ( .A(n3793), .B(n3451), .S(EBX_REG_27__SCAN_IN), .Z(n3794) );
  OAI21_X1 U4377 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n4547), .A(n3794), 
        .ZN(n3795) );
  INV_X1 U4378 ( .A(n3795), .ZN(n5292) );
  NAND2_X1 U4379 ( .A1(n5309), .A2(n5292), .ZN(n3799) );
  NAND2_X1 U4380 ( .A1(n3451), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3796) );
  NAND2_X1 U4381 ( .A1(n3693), .A2(n3796), .ZN(n3798) );
  INV_X1 U4382 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5402) );
  NAND2_X1 U4383 ( .A1(n5241), .A2(n5402), .ZN(n3797) );
  AOI22_X1 U4384 ( .A1(n3798), .A2(n3797), .B1(n4531), .B2(n5402), .ZN(n3800)
         );
  OR2_X2 U4385 ( .A1(n3799), .A2(n3800), .ZN(n5271) );
  NAND2_X1 U4386 ( .A1(n5293), .A2(n3800), .ZN(n3801) );
  NAND2_X1 U4387 ( .A1(n5271), .A2(n3801), .ZN(n5401) );
  AND2_X4 U4388 ( .A1(n6750), .A2(n4564), .ZN(n3818) );
  NAND2_X1 U4389 ( .A1(n4579), .A2(n3818), .ZN(n4562) );
  INV_X1 U4390 ( .A(n3802), .ZN(n3803) );
  NOR2_X1 U4391 ( .A1(n3925), .A2(n3816), .ZN(n4595) );
  NAND2_X1 U4392 ( .A1(n4137), .A2(n6872), .ZN(n3804) );
  NAND2_X1 U4393 ( .A1(n4562), .A2(n3804), .ZN(n3805) );
  NAND3_X1 U4394 ( .A1(n5866), .A2(n5893), .A3(n3806), .ZN(n4121) );
  INV_X1 U4395 ( .A(n5852), .ZN(n3807) );
  NAND2_X1 U4396 ( .A1(n6276), .A2(n3807), .ZN(n5843) );
  INV_X1 U4397 ( .A(n5843), .ZN(n3809) );
  XNOR2_X1 U4398 ( .A(n4143), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3808)
         );
  AND2_X1 U4399 ( .A1(n6277), .A2(REIP_REG_28__SCAN_IN), .ZN(n5701) );
  AOI21_X1 U4400 ( .B1(n3809), .B2(n3808), .A(n5701), .ZN(n3810) );
  OAI21_X1 U4401 ( .B1(n5401), .B2(n6227), .A(n3810), .ZN(n3811) );
  INV_X1 U4402 ( .A(n3811), .ZN(n4142) );
  OAI21_X1 U4403 ( .B1(n3812), .B2(n4586), .A(n6545), .ZN(n3824) );
  NAND2_X1 U4404 ( .A1(n3813), .A2(n4136), .ZN(n3814) );
  NAND2_X1 U4405 ( .A1(n6750), .A2(n6499), .ZN(n3839) );
  AOI21_X1 U4406 ( .B1(n3839), .B2(n6914), .A(n3816), .ZN(n3823) );
  NAND2_X1 U4407 ( .A1(n3817), .A2(n5170), .ZN(n3819) );
  NAND2_X1 U4408 ( .A1(n3819), .A2(n3818), .ZN(n3822) );
  NAND4_X1 U4409 ( .A1(n3824), .A2(n3828), .A3(n3823), .A4(n3835), .ZN(n3825)
         );
  NAND2_X1 U4410 ( .A1(n3825), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3845) );
  INV_X1 U4411 ( .A(n3845), .ZN(n3938) );
  NAND2_X1 U4412 ( .A1(n3938), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3827) );
  NAND2_X1 U4413 ( .A1(n6469), .A2(n6482), .ZN(n4896) );
  MUX2_X1 U4414 ( .A(n3942), .B(n4896), .S(n6709), .Z(n3826) );
  NAND2_X1 U4415 ( .A1(n3827), .A2(n3826), .ZN(n3867) );
  INV_X1 U4416 ( .A(n3828), .ZN(n3829) );
  NAND2_X1 U4417 ( .A1(n3829), .A2(n4586), .ZN(n3834) );
  NAND2_X1 U4418 ( .A1(n6469), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6134) );
  AOI21_X1 U4419 ( .B1(n3830), .B2(n4595), .A(n6134), .ZN(n3833) );
  NAND2_X1 U4420 ( .A1(n3831), .A2(n3818), .ZN(n3832) );
  NAND2_X2 U4421 ( .A1(n3867), .A2(n3868), .ZN(n3934) );
  INV_X1 U4422 ( .A(n3934), .ZN(n3851) );
  NAND2_X1 U4423 ( .A1(n4494), .A2(n3839), .ZN(n3842) );
  NAND2_X2 U4424 ( .A1(n3840), .A2(n6750), .ZN(n4135) );
  INV_X1 U4425 ( .A(n4137), .ZN(n3841) );
  NAND3_X1 U4426 ( .A1(n3842), .A2(n4135), .A3(n3841), .ZN(n3843) );
  NAND2_X1 U4427 ( .A1(n3843), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3846) );
  INV_X1 U4428 ( .A(n4896), .ZN(n3976) );
  NAND2_X1 U4429 ( .A1(n6717), .A2(n6709), .ZN(n3844) );
  NAND2_X1 U4430 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6681) );
  INV_X1 U4431 ( .A(n3942), .ZN(n3975) );
  AOI22_X1 U4432 ( .A1(n3976), .A2(n6677), .B1(n3975), .B2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3847) );
  OAI211_X1 U4433 ( .C1(n3845), .C2(n3467), .A(n3846), .B(n3847), .ZN(n3936)
         );
  INV_X1 U4434 ( .A(n3846), .ZN(n3849) );
  INV_X1 U4435 ( .A(n3847), .ZN(n3848) );
  NAND2_X1 U4436 ( .A1(n3936), .A2(n3850), .ZN(n3933) );
  XNOR2_X1 U4437 ( .A(n3851), .B(n3933), .ZN(n4799) );
  NAND2_X1 U4438 ( .A1(n4799), .A2(n6482), .ZN(n3866) );
  BUF_X1 U4439 ( .A(n3903), .Z(n5085) );
  AOI22_X1 U4440 ( .A1(n3434), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n5085), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4441 ( .A1(n5087), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4442 ( .A1(n5068), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4443 ( .A1(n5037), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3854) );
  NAND4_X1 U4444 ( .A1(n3857), .A2(n3856), .A3(n3855), .A4(n3854), .ZN(n3864)
         );
  AOI22_X1 U4445 ( .A1(n5077), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5036), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4446 ( .A1(n5079), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4447 ( .A1(n5080), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5056), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4448 ( .A1(n5086), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3859) );
  NAND4_X1 U4449 ( .A1(n3862), .A2(n3861), .A3(n3860), .A4(n3859), .ZN(n3863)
         );
  INV_X1 U4450 ( .A(n3867), .ZN(n3870) );
  NAND2_X1 U4451 ( .A1(n3870), .A2(n3869), .ZN(n3871) );
  AND2_X2 U4452 ( .A1(n3871), .A2(n3934), .ZN(n4153) );
  NAND2_X1 U4453 ( .A1(n4072), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3872) );
  OAI211_X1 U4454 ( .C1(n3874), .C2(n3873), .A(n3872), .B(n3913), .ZN(n3875)
         );
  INV_X1 U4455 ( .A(n3875), .ZN(n3876) );
  INV_X1 U4456 ( .A(n3931), .ZN(n3877) );
  XNOR2_X2 U4457 ( .A(n3932), .B(n3877), .ZN(n4146) );
  NAND2_X1 U4458 ( .A1(n4146), .A2(n4085), .ZN(n3894) );
  AOI22_X1 U4459 ( .A1(n5077), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n5078), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4460 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n5076), .B1(n5086), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4461 ( .A1(n5085), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4462 ( .A1(n3434), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4427), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3878) );
  NAND4_X1 U4463 ( .A1(n3881), .A2(n3880), .A3(n3879), .A4(n3878), .ZN(n3887)
         );
  AOI22_X1 U4464 ( .A1(n5068), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3858), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4465 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5036), .B1(n5088), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4466 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n5051), .B1(n5080), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4467 ( .A1(n5087), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3882) );
  NAND4_X1 U4468 ( .A1(n3885), .A2(n3884), .A3(n3883), .A4(n3882), .ZN(n3886)
         );
  XNOR2_X1 U4469 ( .A(n3965), .B(n3964), .ZN(n3891) );
  INV_X1 U4470 ( .A(n3818), .ZN(n4516) );
  INV_X1 U4471 ( .A(n3888), .ZN(n3890) );
  OAI211_X1 U4472 ( .C1(n3891), .C2(n4516), .A(n3890), .B(n3889), .ZN(n3892)
         );
  INV_X1 U4473 ( .A(n3892), .ZN(n3893) );
  NAND2_X1 U4474 ( .A1(n4072), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4475 ( .A1(n3434), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5078), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4476 ( .A1(n5077), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4477 ( .A1(n3858), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3897), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4478 ( .A1(n5088), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3898) );
  NAND4_X1 U4479 ( .A1(n3901), .A2(n3900), .A3(n3899), .A4(n3898), .ZN(n3909)
         );
  AOI22_X1 U4480 ( .A1(n5076), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5085), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4481 ( .A1(n3431), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4482 ( .A1(n5087), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4483 ( .A1(n5068), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4427), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3904) );
  NAND4_X1 U4484 ( .A1(n3907), .A2(n3906), .A3(n3905), .A4(n3904), .ZN(n3908)
         );
  NAND2_X1 U4485 ( .A1(n6872), .A2(n4089), .ZN(n4084) );
  OAI211_X1 U4486 ( .C1(n3914), .C2(n4564), .A(n4084), .B(
        STATE2_REG_0__SCAN_IN), .ZN(n3910) );
  INV_X1 U4487 ( .A(n3910), .ZN(n3911) );
  NAND2_X1 U4488 ( .A1(n3912), .A2(n3911), .ZN(n3919) );
  INV_X1 U4489 ( .A(n3913), .ZN(n3916) );
  XNOR2_X1 U4490 ( .A(n3914), .B(n4089), .ZN(n3915) );
  NAND2_X1 U4491 ( .A1(n3916), .A2(n3915), .ZN(n3920) );
  INV_X1 U4492 ( .A(n3919), .ZN(n3922) );
  INV_X1 U4493 ( .A(n3920), .ZN(n3921) );
  NAND2_X1 U4494 ( .A1(n3922), .A2(n3921), .ZN(n3923) );
  NAND2_X1 U4495 ( .A1(n4761), .A2(n4085), .ZN(n3928) );
  NAND2_X1 U4496 ( .A1(n6545), .A2(n3925), .ZN(n3966) );
  OAI21_X1 U4497 ( .B1(n4516), .B2(n3964), .A(n3966), .ZN(n3926) );
  INV_X1 U4498 ( .A(n3926), .ZN(n3927) );
  NAND2_X1 U4499 ( .A1(n3928), .A2(n3927), .ZN(n4638) );
  NAND2_X1 U4500 ( .A1(n5924), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3929)
         );
  NAND2_X1 U4501 ( .A1(n3930), .A2(n3929), .ZN(n3969) );
  NAND2_X1 U4502 ( .A1(n3969), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6088)
         );
  INV_X1 U4503 ( .A(n3933), .ZN(n3935) );
  NAND2_X1 U4504 ( .A1(n3935), .A2(n3934), .ZN(n3937) );
  NAND2_X1 U4505 ( .A1(n3937), .A2(n3936), .ZN(n3945) );
  INV_X1 U4507 ( .A(n6681), .ZN(n3940) );
  NAND2_X1 U4508 ( .A1(n3940), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6542) );
  NAND2_X1 U4509 ( .A1(n6681), .A2(n6649), .ZN(n3941) );
  NAND2_X1 U4510 ( .A1(n6542), .A2(n3941), .ZN(n6557) );
  OAI22_X1 U4511 ( .A1(n6557), .A2(n4896), .B1(n3942), .B2(n6649), .ZN(n3943)
         );
  NAND2_X1 U4512 ( .A1(n3945), .A2(n3944), .ZN(n3946) );
  AOI22_X1 U4513 ( .A1(n5077), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3950) );
  AOI22_X1 U4514 ( .A1(n5051), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5078), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4515 ( .A1(n5042), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4516 ( .A1(n5086), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3947) );
  NAND4_X1 U4517 ( .A1(n3950), .A2(n3949), .A3(n3948), .A4(n3947), .ZN(n3958)
         );
  AOI22_X1 U4518 ( .A1(n3434), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4519 ( .A1(n5087), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4520 ( .A1(n5068), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5056), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4521 ( .A1(n5079), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3953) );
  NAND4_X1 U4522 ( .A1(n3956), .A2(n3955), .A3(n3954), .A4(n3953), .ZN(n3957)
         );
  AOI22_X1 U4523 ( .A1(n4071), .A2(n3995), .B1(n4072), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3959) );
  OAI21_X2 U4524 ( .B1(n4676), .B2(STATE2_REG_0__SCAN_IN), .A(n3959), .ZN(
        n3963) );
  INV_X1 U4525 ( .A(n3963), .ZN(n3960) );
  NAND2_X1 U4526 ( .A1(n3961), .A2(n3960), .ZN(n6579) );
  NAND2_X1 U4527 ( .A1(n3963), .A2(n3962), .ZN(n3992) );
  NAND2_X1 U4528 ( .A1(n6579), .A2(n3992), .ZN(n4701) );
  INV_X1 U4529 ( .A(n4701), .ZN(n6541) );
  NAND2_X1 U4530 ( .A1(n3965), .A2(n3964), .ZN(n3997) );
  XNOR2_X1 U4531 ( .A(n3997), .B(n3995), .ZN(n3967) );
  OAI21_X1 U4532 ( .B1(n3967), .B2(n4516), .A(n3966), .ZN(n3968) );
  NAND2_X1 U4533 ( .A1(n6088), .A2(n6087), .ZN(n3971) );
  INV_X1 U4534 ( .A(n3969), .ZN(n3970) );
  NAND2_X1 U4535 ( .A1(n3971), .A2(n6089), .ZN(n4002) );
  INV_X1 U4536 ( .A(n4002), .ZN(n3972) );
  INV_X1 U4537 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4001) );
  NAND2_X1 U4538 ( .A1(n3972), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4768)
         );
  NAND2_X1 U4539 ( .A1(n3939), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3978) );
  NAND2_X1 U4540 ( .A1(n6542), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3974) );
  NAND3_X1 U4541 ( .A1(n3500), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6639) );
  INV_X1 U4542 ( .A(n6639), .ZN(n3973) );
  NAND2_X1 U4543 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3973), .ZN(n6627) );
  NAND2_X1 U4544 ( .A1(n3974), .A2(n6627), .ZN(n6676) );
  AOI22_X1 U4545 ( .A1(n6676), .A2(n3976), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3975), .ZN(n3977) );
  NAND2_X1 U4546 ( .A1(n4593), .A2(n6482), .ZN(n3990) );
  AOI22_X1 U4547 ( .A1(n5077), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5079), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4548 ( .A1(n5051), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4549 ( .A1(n5076), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4550 ( .A1(n3853), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3979) );
  NAND4_X1 U4551 ( .A1(n3982), .A2(n3981), .A3(n3980), .A4(n3979), .ZN(n3988)
         );
  AOI22_X1 U4552 ( .A1(n5075), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5078), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3986) );
  AOI22_X1 U4553 ( .A1(n5068), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U4554 ( .A1(n5042), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4555 ( .A1(n3434), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4427), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3983) );
  NAND4_X1 U4556 ( .A1(n3986), .A2(n3985), .A3(n3984), .A4(n3983), .ZN(n3987)
         );
  AOI22_X1 U4557 ( .A1(n4071), .A2(n4016), .B1(n4072), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3989) );
  INV_X1 U4558 ( .A(n4702), .ZN(n3993) );
  NAND2_X1 U4559 ( .A1(n3993), .A2(n3992), .ZN(n3994) );
  AND2_X2 U4560 ( .A1(n4037), .A2(n3994), .ZN(n6666) );
  INV_X1 U4561 ( .A(n3995), .ZN(n3996) );
  NAND2_X1 U4562 ( .A1(n3997), .A2(n3996), .ZN(n4017) );
  INV_X1 U4563 ( .A(n4016), .ZN(n3998) );
  XNOR2_X1 U4564 ( .A(n4017), .B(n3998), .ZN(n3999) );
  AND2_X1 U4565 ( .A1(n3999), .A2(n3818), .ZN(n4000) );
  AOI21_X1 U4566 ( .B1(n6666), .B2(n4085), .A(n4000), .ZN(n4769) );
  NAND2_X1 U4567 ( .A1(n4768), .A2(n4769), .ZN(n4003) );
  NAND2_X1 U4568 ( .A1(n4002), .A2(n4001), .ZN(n4767) );
  NAND2_X1 U4569 ( .A1(n4003), .A2(n4767), .ZN(n4845) );
  AOI22_X1 U4570 ( .A1(n5077), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n5079), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U4571 ( .A1(n5051), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U4572 ( .A1(n5076), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4005) );
  AOI22_X1 U4573 ( .A1(n3853), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4004) );
  NAND4_X1 U4574 ( .A1(n4007), .A2(n4006), .A3(n4005), .A4(n4004), .ZN(n4013)
         );
  AOI22_X1 U4575 ( .A1(n5075), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5078), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4576 ( .A1(n5068), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U4577 ( .A1(n5042), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U4578 ( .A1(n3434), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4427), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4008) );
  NAND4_X1 U4579 ( .A1(n4011), .A2(n4010), .A3(n4009), .A4(n4008), .ZN(n4012)
         );
  NAND2_X1 U4580 ( .A1(n4071), .A2(n4040), .ZN(n4015) );
  NAND2_X1 U4581 ( .A1(n4072), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4014) );
  NAND2_X1 U4582 ( .A1(n4015), .A2(n4014), .ZN(n4035) );
  XNOR2_X1 U4583 ( .A(n4037), .B(n4035), .ZN(n4179) );
  NAND2_X1 U4584 ( .A1(n4179), .A2(n4085), .ZN(n4020) );
  NAND2_X1 U4585 ( .A1(n4017), .A2(n4016), .ZN(n4042) );
  XNOR2_X1 U4586 ( .A(n4042), .B(n4040), .ZN(n4018) );
  NAND2_X1 U4587 ( .A1(n4018), .A2(n3818), .ZN(n4019) );
  NAND2_X1 U4588 ( .A1(n4020), .A2(n4019), .ZN(n4021) );
  NAND2_X1 U4589 ( .A1(n4021), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4022)
         );
  AOI22_X1 U4590 ( .A1(n5077), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U4591 ( .A1(n5042), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U4592 ( .A1(n5068), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U4593 ( .A1(n5088), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4023) );
  NAND4_X1 U4594 ( .A1(n4026), .A2(n4025), .A3(n4024), .A4(n4023), .ZN(n4032)
         );
  AOI22_X1 U4595 ( .A1(n5087), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n5078), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U4596 ( .A1(n5086), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U4597 ( .A1(n5079), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U4598 ( .A1(n3434), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4427), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4027) );
  NAND4_X1 U4599 ( .A1(n4030), .A2(n4029), .A3(n4028), .A4(n4027), .ZN(n4031)
         );
  NAND2_X1 U4600 ( .A1(n4071), .A2(n4043), .ZN(n4034) );
  NAND2_X1 U4601 ( .A1(n4072), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4033) );
  INV_X1 U4602 ( .A(n4085), .ZN(n4046) );
  INV_X1 U4603 ( .A(n4040), .ZN(n4041) );
  NOR2_X1 U4604 ( .A1(n4042), .A2(n4041), .ZN(n4044) );
  NAND2_X1 U4605 ( .A1(n4044), .A2(n4043), .ZN(n4076) );
  OAI211_X1 U4606 ( .C1(n4044), .C2(n4043), .A(n4076), .B(n3818), .ZN(n4045)
         );
  INV_X1 U4607 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4778) );
  NAND2_X1 U4608 ( .A1(n4775), .A2(n4776), .ZN(n4049) );
  NAND2_X1 U4609 ( .A1(n4047), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4048)
         );
  NAND2_X1 U4610 ( .A1(n4049), .A2(n4048), .ZN(n4788) );
  AOI22_X1 U4611 ( .A1(n5077), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n5079), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4053) );
  AOI22_X1 U4612 ( .A1(n5051), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4052) );
  AOI22_X1 U4613 ( .A1(n5076), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4051) );
  AOI22_X1 U4614 ( .A1(n3853), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4050) );
  NAND4_X1 U4615 ( .A1(n4053), .A2(n4052), .A3(n4051), .A4(n4050), .ZN(n4059)
         );
  AOI22_X1 U4616 ( .A1(n5075), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5078), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U4617 ( .A1(n5068), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U4618 ( .A1(n5042), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4055) );
  AOI22_X1 U4619 ( .A1(n3434), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4427), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4054) );
  NAND4_X1 U4620 ( .A1(n4057), .A2(n4056), .A3(n4055), .A4(n4054), .ZN(n4058)
         );
  NAND2_X1 U4621 ( .A1(n4071), .A2(n4077), .ZN(n4061) );
  NAND2_X1 U4622 ( .A1(n4072), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4060) );
  NAND2_X1 U4623 ( .A1(n4065), .A2(n4064), .ZN(n4190) );
  NAND3_X1 U4624 ( .A1(n4088), .A2(n4190), .A3(n4085), .ZN(n4068) );
  XNOR2_X1 U4625 ( .A(n4076), .B(n4077), .ZN(n4066) );
  NAND2_X1 U4626 ( .A1(n4066), .A2(n3818), .ZN(n4067) );
  NAND2_X1 U4627 ( .A1(n4068), .A2(n4067), .ZN(n4069) );
  OR2_X1 U4628 ( .A1(n4069), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4790)
         );
  NAND2_X1 U4629 ( .A1(n4788), .A2(n4790), .ZN(n4070) );
  NAND2_X1 U4630 ( .A1(n4069), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4789)
         );
  NAND2_X1 U4631 ( .A1(n4070), .A2(n4789), .ZN(n6107) );
  NAND2_X1 U4632 ( .A1(n4071), .A2(n4089), .ZN(n4074) );
  NAND2_X1 U4633 ( .A1(n4072), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4073) );
  NAND2_X1 U4634 ( .A1(n4074), .A2(n4073), .ZN(n4075) );
  XNOR2_X2 U4635 ( .A(n4088), .B(n4075), .ZN(n4200) );
  INV_X1 U4636 ( .A(n4076), .ZN(n4078) );
  NAND2_X1 U4637 ( .A1(n4078), .A2(n4077), .ZN(n4091) );
  XNOR2_X1 U4638 ( .A(n4091), .B(n4089), .ZN(n4079) );
  NAND2_X1 U4639 ( .A1(n4079), .A2(n3818), .ZN(n4080) );
  NAND2_X1 U4640 ( .A1(n4081), .A2(n4080), .ZN(n4082) );
  INV_X1 U4641 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6215) );
  XNOR2_X1 U4642 ( .A(n4082), .B(n6215), .ZN(n6106) );
  NAND2_X1 U4643 ( .A1(n6107), .A2(n6106), .ZN(n6109) );
  NAND2_X1 U4644 ( .A1(n4082), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4083)
         );
  NAND2_X1 U4645 ( .A1(n6109), .A2(n4083), .ZN(n4997) );
  INV_X1 U4646 ( .A(n4084), .ZN(n4086) );
  NAND2_X1 U4647 ( .A1(n3818), .A2(n4089), .ZN(n4090) );
  OR2_X1 U4648 ( .A1(n4091), .A2(n4090), .ZN(n4092) );
  NAND2_X1 U4649 ( .A1(n4095), .A2(n4092), .ZN(n4093) );
  XNOR2_X1 U4650 ( .A(n4093), .B(n6209), .ZN(n4996) );
  NAND2_X1 U4651 ( .A1(n4997), .A2(n4996), .ZN(n4918) );
  NAND2_X1 U4652 ( .A1(n4093), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4919)
         );
  INV_X1 U4653 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6244) );
  OR2_X1 U4654 ( .A1(n4095), .A2(n6244), .ZN(n4094) );
  AND2_X1 U4655 ( .A1(n4919), .A2(n4094), .ZN(n4097) );
  INV_X1 U4656 ( .A(n4094), .ZN(n4096) );
  XNOR2_X1 U4657 ( .A(n4095), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4921)
         );
  AOI21_X2 U4658 ( .B1(n4918), .B2(n4097), .A(n3454), .ZN(n4928) );
  NAND2_X1 U4659 ( .A1(n4928), .A2(n3461), .ZN(n4098) );
  NAND2_X1 U4660 ( .A1(n4098), .A2(n5692), .ZN(n4104) );
  INV_X1 U4661 ( .A(n4928), .ZN(n4102) );
  INV_X1 U4662 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4100) );
  INV_X1 U4663 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4099) );
  AND2_X1 U4664 ( .A1(n4100), .A2(n4099), .ZN(n4101) );
  NAND2_X1 U4665 ( .A1(n4102), .A2(n4101), .ZN(n4103) );
  NAND2_X1 U4666 ( .A1(n4104), .A2(n4103), .ZN(n4105) );
  INV_X1 U4667 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6250) );
  NAND2_X1 U4668 ( .A1(n4105), .A2(n4953), .ZN(n4107) );
  NAND2_X1 U4669 ( .A1(n5692), .A2(n4099), .ZN(n4106) );
  NAND2_X1 U4670 ( .A1(n4107), .A2(n4106), .ZN(n5821) );
  XNOR2_X1 U4671 ( .A(n4095), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5822)
         );
  NAND2_X1 U4672 ( .A1(n5821), .A2(n5822), .ZN(n4109) );
  NAND2_X1 U4673 ( .A1(n5692), .A2(n6173), .ZN(n4108) );
  NAND2_X1 U4674 ( .A1(n4109), .A2(n4108), .ZN(n5809) );
  INV_X1 U4675 ( .A(n5809), .ZN(n4111) );
  NAND2_X1 U4676 ( .A1(n4111), .A2(n4110), .ZN(n5800) );
  INV_X1 U4677 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6261) );
  NOR2_X1 U4678 ( .A1(n5692), .A2(n6261), .ZN(n5801) );
  INV_X1 U4679 ( .A(n5801), .ZN(n4112) );
  AND2_X1 U4680 ( .A1(n4112), .A2(n5810), .ZN(n4113) );
  NAND2_X1 U4681 ( .A1(n5692), .A2(n6262), .ZN(n4114) );
  INV_X1 U4682 ( .A(n4115), .ZN(n4116) );
  NAND2_X1 U4683 ( .A1(n5692), .A2(n4116), .ZN(n4117) );
  INV_X1 U4684 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6272) );
  AND3_X1 U4685 ( .A1(n6272), .A2(n6262), .A3(n5908), .ZN(n4118) );
  NOR2_X1 U4686 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5894) );
  NOR2_X1 U4687 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5740) );
  INV_X1 U4688 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5865) );
  AND4_X1 U4689 ( .A1(n5894), .A2(n5740), .A3(n5865), .A4(n5859), .ZN(n4120)
         );
  NOR2_X1 U4690 ( .A1(n5692), .A2(n4120), .ZN(n4123) );
  NAND2_X1 U4691 ( .A1(n5692), .A2(n4121), .ZN(n4122) );
  XNOR2_X1 U4692 ( .A(n5692), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5730)
         );
  INV_X1 U4693 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6285) );
  AND2_X1 U4694 ( .A1(n5692), .A2(n6285), .ZN(n4124) );
  NAND2_X1 U4695 ( .A1(n5692), .A2(n5708), .ZN(n5717) );
  INV_X1 U4696 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4126) );
  NAND2_X1 U4697 ( .A1(n4125), .A2(n3459), .ZN(n5688) );
  NAND2_X1 U4698 ( .A1(n5708), .A2(n4126), .ZN(n4523) );
  INV_X1 U4699 ( .A(n4523), .ZN(n4127) );
  OR2_X1 U4700 ( .A1(n5692), .A2(n4127), .ZN(n4128) );
  NAND2_X1 U4701 ( .A1(n5688), .A2(n4128), .ZN(n4130) );
  XNOR2_X1 U4702 ( .A(n5692), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4129)
         );
  XNOR2_X1 U4703 ( .A(n4130), .B(n4129), .ZN(n5707) );
  NOR2_X1 U4704 ( .A1(n4132), .A2(n4131), .ZN(n6448) );
  INV_X1 U4705 ( .A(n6448), .ZN(n4134) );
  NAND2_X1 U4706 ( .A1(n4133), .A2(n5240), .ZN(n4600) );
  AND2_X1 U4707 ( .A1(n4134), .A2(n4600), .ZN(n5230) );
  NAND2_X1 U4708 ( .A1(n4137), .A2(n4136), .ZN(n4139) );
  NAND2_X1 U4709 ( .A1(n4579), .A2(n5241), .ZN(n4138) );
  NAND4_X1 U4710 ( .A1(n5230), .A2(n4135), .A3(n4139), .A4(n4138), .ZN(n4140)
         );
  OAI211_X1 U4711 ( .C1(n4143), .C2(n5839), .A(n4142), .B(n3465), .ZN(U2990)
         );
  NAND2_X1 U4712 ( .A1(n6720), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4286) );
  NAND2_X1 U4713 ( .A1(n3616), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4167) );
  OAI21_X1 U4714 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n4162), .ZN(n6095) );
  AOI22_X1 U4715 ( .A1(n5220), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n5154), 
        .B2(n6095), .ZN(n4145) );
  NOR2_X2 U4716 ( .A1(n5170), .A2(n6720), .ZN(n4154) );
  NAND2_X1 U4717 ( .A1(n5221), .A2(EAX_REG_2__SCAN_IN), .ZN(n4144) );
  OAI211_X1 U4718 ( .C1(n4167), .C2(n5218), .A(n4145), .B(n4144), .ZN(n4159)
         );
  NAND2_X1 U4719 ( .A1(n4160), .A2(n4159), .ZN(n4158) );
  NAND2_X1 U4720 ( .A1(n6663), .A2(n4314), .ZN(n4150) );
  AOI22_X1 U4721 ( .A1(n5221), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6720), .ZN(n4147) );
  INV_X1 U4722 ( .A(n4148), .ZN(n4149) );
  NAND2_X1 U4723 ( .A1(n6955), .A2(n5170), .ZN(n4151) );
  OR2_X1 U4724 ( .A1(n4761), .A2(n4151), .ZN(n4152) );
  NAND2_X1 U4725 ( .A1(n4152), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4557) );
  INV_X1 U4726 ( .A(n4153), .ZN(n6629) );
  AOI22_X1 U4727 ( .A1(n4154), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6720), .ZN(n4156) );
  INV_X1 U4728 ( .A(n4167), .ZN(n4171) );
  NAND2_X1 U4729 ( .A1(n4171), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4155) );
  OAI211_X1 U4730 ( .C1(n6629), .C2(n4304), .A(n4156), .B(n4155), .ZN(n4556)
         );
  MUX2_X1 U4731 ( .A(n5141), .B(n4557), .S(n4556), .Z(n4157) );
  INV_X1 U4732 ( .A(n4157), .ZN(n4559) );
  NAND2_X1 U4733 ( .A1(n4560), .A2(n4559), .ZN(n4558) );
  NAND2_X1 U4734 ( .A1(n4158), .A2(n4558), .ZN(n4161) );
  OR2_X1 U4735 ( .A1(n4160), .A2(n4159), .ZN(n4670) );
  NAND2_X1 U4736 ( .A1(n4161), .A2(n4670), .ZN(n4611) );
  INV_X1 U4737 ( .A(n4611), .ZN(n4170) );
  INV_X1 U4738 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4601) );
  INV_X1 U4739 ( .A(n4162), .ZN(n4164) );
  INV_X1 U4740 ( .A(n4174), .ZN(n4163) );
  OAI21_X1 U4741 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n4164), .A(n4163), 
        .ZN(n5387) );
  AOI22_X1 U4742 ( .A1(n5154), .A2(n5387), .B1(n5220), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4166) );
  NAND2_X1 U4743 ( .A1(n5221), .A2(EAX_REG_3__SCAN_IN), .ZN(n4165) );
  OAI211_X1 U4744 ( .C1(n4167), .C2(n4601), .A(n4166), .B(n4165), .ZN(n4168)
         );
  AOI21_X1 U4745 ( .B1(n6666), .B2(n4314), .A(n4168), .ZN(n4612) );
  NAND2_X1 U4746 ( .A1(n4170), .A2(n4169), .ZN(n4610) );
  NAND2_X1 U4747 ( .A1(n4171), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4177) );
  INV_X1 U4748 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4172) );
  AOI21_X1 U4749 ( .B1(n4172), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4173) );
  AOI21_X1 U4750 ( .B1(n5221), .B2(EAX_REG_4__SCAN_IN), .A(n4173), .ZN(n4176)
         );
  OAI21_X1 U4751 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n4174), .A(n4181), 
        .ZN(n6299) );
  NOR2_X1 U4752 ( .A1(n6299), .A2(n5141), .ZN(n4175) );
  AOI21_X1 U4753 ( .B1(n4177), .B2(n4176), .A(n4175), .ZN(n4178) );
  AOI21_X1 U4754 ( .B1(n4179), .B2(n4314), .A(n4178), .ZN(n4644) );
  NOR2_X2 U4755 ( .A1(n4610), .A2(n4644), .ZN(n4645) );
  INV_X1 U4756 ( .A(n4181), .ZN(n4183) );
  INV_X1 U4757 ( .A(n4193), .ZN(n4182) );
  OAI21_X1 U4758 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n4183), .A(n4182), 
        .ZN(n6321) );
  NAND2_X1 U4759 ( .A1(n6321), .A2(n5154), .ZN(n4184) );
  OAI21_X1 U4760 ( .B1(n6100), .B2(n4286), .A(n4184), .ZN(n4185) );
  AOI21_X1 U4761 ( .B1(n5221), .B2(EAX_REG_5__SCAN_IN), .A(n4185), .ZN(n4186)
         );
  NAND2_X1 U4762 ( .A1(n4645), .A2(n4654), .ZN(n4653) );
  INV_X1 U4763 ( .A(n4653), .ZN(n4192) );
  INV_X1 U4764 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4727) );
  XNOR2_X1 U4765 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .B(n4193), .ZN(n6332) );
  AOI22_X1 U4766 ( .A1(n5154), .A2(n6332), .B1(n5220), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4188) );
  OAI21_X1 U4767 ( .B1(n4388), .B2(n4727), .A(n4188), .ZN(n4189) );
  NAND2_X1 U4768 ( .A1(n4192), .A2(n4191), .ZN(n4816) );
  INV_X1 U4769 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4730) );
  INV_X1 U4770 ( .A(n4214), .ZN(n4197) );
  INV_X1 U4771 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4195) );
  NAND2_X1 U4772 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n4193), .ZN(n4194)
         );
  NAND2_X1 U4773 ( .A1(n4195), .A2(n4194), .ZN(n4196) );
  NAND2_X1 U4774 ( .A1(n4197), .A2(n4196), .ZN(n6346) );
  AOI22_X1 U4775 ( .A1(n6346), .A2(n5154), .B1(n5220), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4198) );
  OAI21_X1 U4776 ( .B1(n4388), .B2(n4730), .A(n4198), .ZN(n4199) );
  NOR2_X2 U4777 ( .A1(n4816), .A2(n4815), .ZN(n4806) );
  AOI22_X1 U4778 ( .A1(n5068), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4204) );
  AOI22_X1 U4779 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n5076), .B1(n5086), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4203) );
  AOI22_X1 U4780 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n5042), .B1(n3435), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4202) );
  AOI22_X1 U4781 ( .A1(n5079), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4201) );
  NAND4_X1 U4782 ( .A1(n4204), .A2(n4203), .A3(n4202), .A4(n4201), .ZN(n4210)
         );
  AOI22_X1 U4783 ( .A1(n3434), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4208) );
  AOI22_X1 U4784 ( .A1(n5077), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4207) );
  AOI22_X1 U4785 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(n3853), .B1(n5080), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4206) );
  AOI22_X1 U4786 ( .A1(n5037), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n5056), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4205) );
  NAND4_X1 U4787 ( .A1(n4208), .A2(n4207), .A3(n4206), .A4(n4205), .ZN(n4209)
         );
  NOR2_X1 U4788 ( .A1(n4210), .A2(n4209), .ZN(n4213) );
  XNOR2_X1 U4789 ( .A(n4214), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5376) );
  AOI22_X1 U4790 ( .A1(n5376), .A2(n5154), .B1(n5220), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4212) );
  NAND2_X1 U4791 ( .A1(n5221), .A2(EAX_REG_8__SCAN_IN), .ZN(n4211) );
  OAI211_X1 U4792 ( .C1(n4304), .C2(n4213), .A(n4212), .B(n4211), .ZN(n4805)
         );
  AND2_X2 U4793 ( .A1(n4806), .A2(n4805), .ZN(n4808) );
  XNOR2_X1 U4794 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n4228), .ZN(n4926) );
  AOI22_X1 U4795 ( .A1(n5087), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4218) );
  AOI22_X1 U4796 ( .A1(n5076), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5042), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4217) );
  AOI22_X1 U4797 ( .A1(n3434), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4216) );
  AOI22_X1 U4798 ( .A1(n5079), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4215) );
  NAND4_X1 U4799 ( .A1(n4218), .A2(n4217), .A3(n4216), .A4(n4215), .ZN(n4224)
         );
  AOI22_X1 U4800 ( .A1(n5037), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4222) );
  AOI22_X1 U4801 ( .A1(n5051), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4221) );
  AOI22_X1 U4802 ( .A1(n5068), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4427), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4220) );
  AOI22_X1 U4803 ( .A1(n5077), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4219) );
  NAND4_X1 U4804 ( .A1(n4222), .A2(n4221), .A3(n4220), .A4(n4219), .ZN(n4223)
         );
  OR2_X1 U4805 ( .A1(n4224), .A2(n4223), .ZN(n4225) );
  AOI22_X1 U4806 ( .A1(n4314), .A2(n4225), .B1(n5220), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4227) );
  NAND2_X1 U4807 ( .A1(n4154), .A2(EAX_REG_9__SCAN_IN), .ZN(n4226) );
  OAI211_X1 U4808 ( .C1(n4926), .C2(n5141), .A(n4227), .B(n4226), .ZN(n4821)
         );
  NAND2_X1 U4809 ( .A1(n4808), .A2(n4821), .ZN(n4820) );
  XNOR2_X1 U4810 ( .A(n4244), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4939)
         );
  AOI22_X1 U4811 ( .A1(n5076), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5042), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4233) );
  AOI22_X1 U4812 ( .A1(n5075), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4229), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4232) );
  AOI22_X1 U4813 ( .A1(n5088), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4231) );
  AOI22_X1 U4814 ( .A1(n5068), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4427), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4230) );
  NAND4_X1 U4815 ( .A1(n4233), .A2(n4232), .A3(n4231), .A4(n4230), .ZN(n4239)
         );
  AOI22_X1 U4816 ( .A1(n3434), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5078), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4237) );
  AOI22_X1 U4817 ( .A1(n5077), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n5087), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4236) );
  AOI22_X1 U4818 ( .A1(n5079), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4235) );
  AOI22_X1 U4819 ( .A1(n5051), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4234) );
  NAND4_X1 U4820 ( .A1(n4237), .A2(n4236), .A3(n4235), .A4(n4234), .ZN(n4238)
         );
  OAI21_X1 U4821 ( .B1(n4239), .B2(n4238), .A(n4314), .ZN(n4242) );
  NAND2_X1 U4822 ( .A1(n4154), .A2(EAX_REG_10__SCAN_IN), .ZN(n4241) );
  NAND2_X1 U4823 ( .A1(n5220), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4240)
         );
  NAND3_X1 U4824 ( .A1(n4242), .A2(n4241), .A3(n4240), .ZN(n4243) );
  AOI21_X1 U4825 ( .B1(n4939), .B2(n5154), .A(n4243), .ZN(n4856) );
  OR2_X2 U4826 ( .A1(n4820), .A2(n4856), .ZN(n4877) );
  XNOR2_X1 U4827 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n4259), .ZN(n4933)
         );
  AOI22_X1 U4828 ( .A1(n5079), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4248) );
  AOI22_X1 U4829 ( .A1(n5085), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4247) );
  AOI22_X1 U4830 ( .A1(n5077), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4246) );
  AOI22_X1 U4831 ( .A1(n5068), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5056), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4245) );
  NAND4_X1 U4832 ( .A1(n4248), .A2(n4247), .A3(n4246), .A4(n4245), .ZN(n4254)
         );
  AOI22_X1 U4833 ( .A1(n5051), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5078), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4252) );
  AOI22_X1 U4834 ( .A1(n5087), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4251) );
  AOI22_X1 U4835 ( .A1(n3434), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4250) );
  AOI22_X1 U4836 ( .A1(n5075), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4249) );
  NAND4_X1 U4837 ( .A1(n4252), .A2(n4251), .A3(n4250), .A4(n4249), .ZN(n4253)
         );
  OAI21_X1 U4838 ( .B1(n4254), .B2(n4253), .A(n4314), .ZN(n4257) );
  NAND2_X1 U4839 ( .A1(n4154), .A2(EAX_REG_11__SCAN_IN), .ZN(n4256) );
  NAND2_X1 U4840 ( .A1(n5220), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4255)
         );
  NAND3_X1 U4841 ( .A1(n4257), .A2(n4256), .A3(n4255), .ZN(n4258) );
  AOI21_X1 U4842 ( .B1(n4933), .B2(n5154), .A(n4258), .ZN(n4876) );
  NOR2_X4 U4843 ( .A1(n4877), .A2(n4876), .ZN(n4907) );
  AOI22_X1 U4844 ( .A1(n4154), .A2(EAX_REG_12__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6720), .ZN(n4272) );
  XNOR2_X1 U4845 ( .A(n4285), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4971)
         );
  NAND2_X1 U4846 ( .A1(n4971), .A2(n5154), .ZN(n4271) );
  AOI22_X1 U4847 ( .A1(n5076), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5079), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4263) );
  AOI22_X1 U4848 ( .A1(n5087), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n5078), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4262) );
  AOI22_X1 U4849 ( .A1(n3435), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4261) );
  AOI22_X1 U4850 ( .A1(n3434), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n5056), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4260) );
  NAND4_X1 U4851 ( .A1(n4263), .A2(n4262), .A3(n4261), .A4(n4260), .ZN(n4269)
         );
  AOI22_X1 U4852 ( .A1(n5085), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4267) );
  AOI22_X1 U4853 ( .A1(n5068), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4266) );
  AOI22_X1 U4854 ( .A1(n5077), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4265) );
  AOI22_X1 U4855 ( .A1(n5075), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4264) );
  NAND4_X1 U4856 ( .A1(n4267), .A2(n4266), .A3(n4265), .A4(n4264), .ZN(n4268)
         );
  OAI21_X1 U4857 ( .B1(n4269), .B2(n4268), .A(n4314), .ZN(n4270) );
  OAI211_X1 U4858 ( .C1(n5154), .C2(n4272), .A(n4271), .B(n4270), .ZN(n4906)
         );
  NAND2_X2 U4859 ( .A1(n4907), .A2(n4906), .ZN(n4905) );
  AOI22_X1 U4860 ( .A1(n5077), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n5068), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4277) );
  AOI22_X1 U4861 ( .A1(n5079), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4276) );
  AOI22_X1 U4862 ( .A1(n3434), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4427), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4275) );
  AOI22_X1 U4863 ( .A1(n3435), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4274) );
  NAND4_X1 U4864 ( .A1(n4277), .A2(n4276), .A3(n4275), .A4(n4274), .ZN(n4283)
         );
  AOI22_X1 U4865 ( .A1(n5075), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5078), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4281) );
  AOI22_X1 U4866 ( .A1(n5085), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4280) );
  AOI22_X1 U4867 ( .A1(n5087), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4279) );
  AOI22_X1 U4868 ( .A1(n5076), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4278) );
  NAND4_X1 U4869 ( .A1(n4281), .A2(n4280), .A3(n4279), .A4(n4278), .ZN(n4282)
         );
  OR2_X1 U4870 ( .A1(n4283), .A2(n4282), .ZN(n4284) );
  NAND2_X1 U4871 ( .A1(n4314), .A2(n4284), .ZN(n4288) );
  XNOR2_X1 U4872 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(n4300), .ZN(n5825)
         );
  OAI22_X1 U4873 ( .A1(n5141), .A2(n5825), .B1(n4286), .B2(n5823), .ZN(n4287)
         );
  AOI21_X1 U4874 ( .B1(n4154), .B2(EAX_REG_13__SCAN_IN), .A(n4287), .ZN(n4977)
         );
  OAI21_X2 U4875 ( .B1(n4976), .B2(n4977), .A(n4289), .ZN(n5363) );
  AOI22_X1 U4876 ( .A1(n5042), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n5079), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4293) );
  AOI22_X1 U4877 ( .A1(n5077), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4292) );
  AOI22_X1 U4878 ( .A1(n5037), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4291) );
  AOI22_X1 U4879 ( .A1(n5088), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4290) );
  NAND4_X1 U4880 ( .A1(n4293), .A2(n4292), .A3(n4291), .A4(n4290), .ZN(n4299)
         );
  AOI22_X1 U4881 ( .A1(n5087), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n5068), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4297) );
  AOI22_X1 U4882 ( .A1(n5076), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4296) );
  AOI22_X1 U4883 ( .A1(n5075), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4295) );
  AOI22_X1 U4884 ( .A1(n3434), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4427), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4294) );
  NAND4_X1 U4885 ( .A1(n4297), .A2(n4296), .A3(n4295), .A4(n4294), .ZN(n4298)
         );
  NOR2_X1 U4886 ( .A1(n4299), .A2(n4298), .ZN(n4303) );
  XNOR2_X1 U4887 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4305), .ZN(n5816)
         );
  AOI22_X1 U4888 ( .A1(n5154), .A2(n5816), .B1(n5220), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4302) );
  NAND2_X1 U4889 ( .A1(n4154), .A2(EAX_REG_14__SCAN_IN), .ZN(n4301) );
  OAI211_X1 U4890 ( .C1(n4304), .C2(n4303), .A(n4302), .B(n4301), .ZN(n5362)
         );
  NAND2_X1 U4891 ( .A1(n5363), .A2(n5362), .ZN(n5361) );
  XNOR2_X1 U4892 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n4322), .ZN(n6353)
         );
  INV_X1 U4893 ( .A(n6353), .ZN(n4321) );
  AOI22_X1 U4894 ( .A1(n3853), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4309) );
  AOI22_X1 U4895 ( .A1(n5079), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5078), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4308) );
  AOI22_X1 U4896 ( .A1(n5080), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4427), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4307) );
  AOI22_X1 U4897 ( .A1(n5075), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4306) );
  NAND4_X1 U4898 ( .A1(n4309), .A2(n4308), .A3(n4307), .A4(n4306), .ZN(n4316)
         );
  AOI22_X1 U4899 ( .A1(n5068), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5085), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4313) );
  AOI22_X1 U4900 ( .A1(n5077), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4312) );
  AOI22_X1 U4901 ( .A1(n5051), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4311) );
  AOI22_X1 U4902 ( .A1(n3434), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4310) );
  NAND4_X1 U4903 ( .A1(n4313), .A2(n4312), .A3(n4311), .A4(n4310), .ZN(n4315)
         );
  OAI21_X1 U4904 ( .B1(n4316), .B2(n4315), .A(n4314), .ZN(n4319) );
  NAND2_X1 U4905 ( .A1(n4154), .A2(EAX_REG_15__SCAN_IN), .ZN(n4318) );
  NAND2_X1 U4906 ( .A1(n5220), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4317)
         );
  NAND3_X1 U4907 ( .A1(n4319), .A2(n4318), .A3(n4317), .ZN(n4320) );
  AOI21_X1 U4908 ( .B1(n4321), .B2(n5154), .A(n4320), .ZN(n5439) );
  NOR2_X2 U4909 ( .A1(n5361), .A2(n5439), .ZN(n5349) );
  INV_X1 U4910 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4323) );
  XNOR2_X1 U4911 ( .A(n4350), .B(n4323), .ZN(n5794) );
  AOI22_X1 U4912 ( .A1(n4154), .A2(EAX_REG_16__SCAN_IN), .B1(n5220), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4335) );
  AOI22_X1 U4913 ( .A1(n5075), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4327) );
  AOI22_X1 U4914 ( .A1(n5079), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4326) );
  AOI22_X1 U4915 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(n5085), .B1(n5080), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4325) );
  AOI22_X1 U4916 ( .A1(n5037), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4427), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4324) );
  NAND4_X1 U4917 ( .A1(n4327), .A2(n4326), .A3(n4325), .A4(n4324), .ZN(n4333)
         );
  AOI22_X1 U4918 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n5077), .B1(n3434), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4331) );
  AOI22_X1 U4919 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n5087), .B1(n5076), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4330) );
  AOI22_X1 U4920 ( .A1(n5068), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4329) );
  AOI22_X1 U4921 ( .A1(n5086), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4328) );
  NAND4_X1 U4922 ( .A1(n4331), .A2(n4330), .A3(n4329), .A4(n4328), .ZN(n4332)
         );
  OAI21_X1 U4923 ( .B1(n4333), .B2(n4332), .A(n5149), .ZN(n4334) );
  OAI211_X1 U4924 ( .C1(n5794), .C2(n5141), .A(n4335), .B(n4334), .ZN(n5351)
         );
  NAND2_X1 U4925 ( .A1(n5349), .A2(n5351), .ZN(n5333) );
  INV_X1 U4926 ( .A(n5333), .ZN(n4355) );
  AOI22_X1 U4927 ( .A1(n5068), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5085), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4339) );
  AOI22_X1 U4928 ( .A1(n5079), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4338) );
  AOI22_X1 U4929 ( .A1(n3434), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4427), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4337) );
  AOI22_X1 U4930 ( .A1(n5075), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4336) );
  NAND4_X1 U4931 ( .A1(n4339), .A2(n4338), .A3(n4337), .A4(n4336), .ZN(n4345)
         );
  AOI22_X1 U4932 ( .A1(n5087), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n5078), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4343) );
  AOI22_X1 U4933 ( .A1(n5076), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4342) );
  AOI22_X1 U4934 ( .A1(n5086), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4341) );
  AOI22_X1 U4935 ( .A1(n5077), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4340) );
  NAND4_X1 U4936 ( .A1(n4343), .A2(n4342), .A3(n4341), .A4(n4340), .ZN(n4344)
         );
  NOR2_X1 U4937 ( .A1(n4345), .A2(n4344), .ZN(n4349) );
  OAI21_X1 U4938 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6736), .A(n6720), 
        .ZN(n4346) );
  INV_X1 U4939 ( .A(n4346), .ZN(n4347) );
  AOI21_X1 U4940 ( .B1(n4154), .B2(EAX_REG_17__SCAN_IN), .A(n4347), .ZN(n4348)
         );
  OAI21_X1 U4941 ( .B1(n5134), .B2(n4349), .A(n4348), .ZN(n4353) );
  OAI21_X1 U4942 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n4351), .A(n4373), 
        .ZN(n6121) );
  OR2_X1 U4943 ( .A1(n5141), .A2(n6121), .ZN(n4352) );
  NAND2_X1 U4944 ( .A1(n4353), .A2(n4352), .ZN(n5337) );
  NAND2_X1 U4945 ( .A1(n4355), .A2(n4354), .ZN(n5318) );
  AOI22_X1 U4946 ( .A1(n5075), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5085), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4359) );
  AOI22_X1 U4947 ( .A1(n5077), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n5087), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4358) );
  AOI22_X1 U4948 ( .A1(n5076), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4357) );
  AOI22_X1 U4949 ( .A1(n3434), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4356) );
  NAND4_X1 U4950 ( .A1(n4359), .A2(n4358), .A3(n4357), .A4(n4356), .ZN(n4367)
         );
  AOI22_X1 U4951 ( .A1(n5068), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5079), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4365) );
  AOI22_X1 U4952 ( .A1(n5086), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4364) );
  AOI22_X1 U4953 ( .A1(n5037), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4363) );
  NAND2_X1 U4954 ( .A1(n5063), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4361) );
  NAND2_X1 U4955 ( .A1(n4427), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4360) );
  AND3_X1 U4956 ( .A1(n4361), .A2(n4360), .A3(n5141), .ZN(n4362) );
  NAND4_X1 U4957 ( .A1(n4365), .A2(n4364), .A3(n4363), .A4(n4362), .ZN(n4366)
         );
  NAND2_X1 U4958 ( .A1(n5134), .A2(n5141), .ZN(n4441) );
  OAI21_X1 U4959 ( .B1(n4367), .B2(n4366), .A(n4441), .ZN(n4369) );
  AOI22_X1 U4960 ( .A1(n5221), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6720), .ZN(n4368) );
  NAND2_X1 U4961 ( .A1(n4369), .A2(n4368), .ZN(n4371) );
  XNOR2_X1 U4962 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n4373), .ZN(n5786)
         );
  NAND2_X1 U4963 ( .A1(n5786), .A2(n5154), .ZN(n4370) );
  NAND2_X1 U4964 ( .A1(n4371), .A2(n4370), .ZN(n5321) );
  NOR2_X2 U4965 ( .A1(n5318), .A2(n5321), .ZN(n5319) );
  INV_X1 U4966 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4372) );
  OR2_X1 U4967 ( .A1(n4374), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4375)
         );
  NAND2_X1 U4968 ( .A1(n4375), .A2(n4422), .ZN(n6357) );
  AOI22_X1 U4969 ( .A1(n5042), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n5078), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4379) );
  AOI22_X1 U4970 ( .A1(n5087), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5079), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4378) );
  AOI22_X1 U4971 ( .A1(n5076), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4377) );
  AOI22_X1 U4972 ( .A1(n5075), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4376) );
  NAND4_X1 U4973 ( .A1(n4379), .A2(n4378), .A3(n4377), .A4(n4376), .ZN(n4385)
         );
  AOI22_X1 U4974 ( .A1(n5068), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4383) );
  AOI22_X1 U4975 ( .A1(n3435), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4382) );
  AOI22_X1 U4976 ( .A1(n3434), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4427), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4381) );
  AOI22_X1 U4977 ( .A1(n5077), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4380) );
  NAND4_X1 U4978 ( .A1(n4383), .A2(n4382), .A3(n4381), .A4(n4380), .ZN(n4384)
         );
  NOR2_X1 U4979 ( .A1(n4385), .A2(n4384), .ZN(n4386) );
  NOR2_X1 U4980 ( .A1(n5134), .A2(n4386), .ZN(n4390) );
  INV_X1 U4981 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4724) );
  NAND2_X1 U4982 ( .A1(n6720), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4387)
         );
  OAI211_X1 U4983 ( .C1(n4388), .C2(n4724), .A(n5141), .B(n4387), .ZN(n4389)
         );
  OAI22_X1 U4984 ( .A1(n6357), .A2(n5141), .B1(n4390), .B2(n4389), .ZN(n6065)
         );
  NAND2_X1 U4985 ( .A1(n5319), .A2(n4391), .ZN(n5427) );
  AOI22_X1 U4986 ( .A1(n5075), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n5078), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4395) );
  AOI22_X1 U4987 ( .A1(n5087), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4394) );
  AOI22_X1 U4988 ( .A1(n5051), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4393) );
  AOI22_X1 U4989 ( .A1(n3434), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4392) );
  NAND4_X1 U4990 ( .A1(n4395), .A2(n4394), .A3(n4393), .A4(n4392), .ZN(n4403)
         );
  AOI22_X1 U4991 ( .A1(n5068), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5085), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4401) );
  AOI22_X1 U4992 ( .A1(n5077), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n5079), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4400) );
  AOI22_X1 U4993 ( .A1(n3435), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4399) );
  NAND2_X1 U4994 ( .A1(n5076), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4397)
         );
  AOI21_X1 U4995 ( .B1(n4427), .B2(INSTQUEUE_REG_9__4__SCAN_IN), .A(n5154), 
        .ZN(n4396) );
  AND2_X1 U4996 ( .A1(n4397), .A2(n4396), .ZN(n4398) );
  NAND4_X1 U4997 ( .A1(n4401), .A2(n4400), .A3(n4399), .A4(n4398), .ZN(n4402)
         );
  OAI21_X1 U4998 ( .B1(n4403), .B2(n4402), .A(n4441), .ZN(n4405) );
  AOI22_X1 U4999 ( .A1(n5221), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6720), .ZN(n4404) );
  NAND2_X1 U5000 ( .A1(n4405), .A2(n4404), .ZN(n4407) );
  XNOR2_X1 U5001 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n4422), .ZN(n6369)
         );
  NAND2_X1 U5002 ( .A1(n6369), .A2(n5154), .ZN(n4406) );
  NAND2_X1 U5003 ( .A1(n4407), .A2(n4406), .ZN(n5428) );
  NOR2_X2 U5004 ( .A1(n5427), .A2(n5428), .ZN(n5425) );
  AOI22_X1 U5005 ( .A1(n5075), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5079), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4411) );
  AOI22_X1 U5006 ( .A1(n5077), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n5085), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4410) );
  AOI22_X1 U5007 ( .A1(n5076), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4409) );
  AOI22_X1 U5008 ( .A1(n3434), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4408) );
  NAND4_X1 U5009 ( .A1(n4411), .A2(n4410), .A3(n4409), .A4(n4408), .ZN(n4417)
         );
  AOI22_X1 U5010 ( .A1(n5037), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4415) );
  AOI22_X1 U5011 ( .A1(n5051), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4414) );
  AOI22_X1 U5012 ( .A1(n5068), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4427), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4413) );
  AOI22_X1 U5013 ( .A1(n3853), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4412) );
  NAND4_X1 U5014 ( .A1(n4415), .A2(n4414), .A3(n4413), .A4(n4412), .ZN(n4416)
         );
  NOR2_X1 U5015 ( .A1(n4417), .A2(n4416), .ZN(n4421) );
  NAND2_X1 U5016 ( .A1(n6720), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4418)
         );
  NAND2_X1 U5017 ( .A1(n5141), .A2(n4418), .ZN(n4419) );
  AOI21_X1 U5018 ( .B1(n4154), .B2(EAX_REG_21__SCAN_IN), .A(n4419), .ZN(n4420)
         );
  OAI21_X1 U5019 ( .B1(n5134), .B2(n4421), .A(n4420), .ZN(n4426) );
  OAI21_X1 U5020 ( .B1(n4424), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n4470), 
        .ZN(n6387) );
  OR2_X1 U5021 ( .A1(n6387), .A2(n5141), .ZN(n4425) );
  AND2_X2 U5022 ( .A1(n5425), .A2(n5764), .ZN(n5414) );
  AOI22_X1 U5023 ( .A1(n5079), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4433) );
  AOI22_X1 U5024 ( .A1(n5051), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4432) );
  NAND2_X1 U5025 ( .A1(n5076), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4429)
         );
  AOI21_X1 U5026 ( .B1(n4427), .B2(INSTQUEUE_REG_9__6__SCAN_IN), .A(n5154), 
        .ZN(n4428) );
  AND2_X1 U5027 ( .A1(n4429), .A2(n4428), .ZN(n4431) );
  AOI22_X1 U5028 ( .A1(n5077), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4430) );
  NAND4_X1 U5029 ( .A1(n4433), .A2(n4432), .A3(n4431), .A4(n4430), .ZN(n4439)
         );
  AOI22_X1 U5030 ( .A1(n5068), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5078), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4437) );
  AOI22_X1 U5031 ( .A1(n5075), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5042), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4436) );
  AOI22_X1 U5032 ( .A1(n5087), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4435) );
  AOI22_X1 U5033 ( .A1(n3434), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4434) );
  NAND4_X1 U5034 ( .A1(n4437), .A2(n4436), .A3(n4435), .A4(n4434), .ZN(n4438)
         );
  OR2_X1 U5035 ( .A1(n4439), .A2(n4438), .ZN(n4440) );
  NAND2_X1 U5036 ( .A1(n4441), .A2(n4440), .ZN(n4445) );
  INV_X1 U5037 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5760) );
  NOR2_X1 U5038 ( .A1(n5760), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4442) );
  AOI21_X1 U5039 ( .B1(n4154), .B2(EAX_REG_22__SCAN_IN), .A(n4442), .ZN(n4444)
         );
  XNOR2_X1 U5040 ( .A(n4470), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6398)
         );
  AOI22_X1 U5041 ( .A1(n5079), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n5078), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4449) );
  AOI22_X1 U5042 ( .A1(n5075), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4448) );
  AOI22_X1 U5043 ( .A1(n5080), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n5056), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4447) );
  AOI22_X1 U5044 ( .A1(n5086), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4446) );
  NAND4_X1 U5045 ( .A1(n4449), .A2(n4448), .A3(n4447), .A4(n4446), .ZN(n4455)
         );
  AOI22_X1 U5046 ( .A1(n5068), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5042), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4453) );
  AOI22_X1 U5047 ( .A1(n5077), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3853), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4452) );
  AOI22_X1 U5048 ( .A1(n5076), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4451) );
  AOI22_X1 U5049 ( .A1(n3434), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4450) );
  NAND4_X1 U5050 ( .A1(n4453), .A2(n4452), .A3(n4451), .A4(n4450), .ZN(n4454)
         );
  NOR2_X1 U5051 ( .A1(n4455), .A2(n4454), .ZN(n4475) );
  AOI22_X1 U5052 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n5042), .B1(n5088), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4459) );
  AOI22_X1 U5053 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n5086), .B1(n3435), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4458) );
  AOI22_X1 U5054 ( .A1(n5075), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5056), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4457) );
  AOI22_X1 U5055 ( .A1(n5051), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4456) );
  NAND4_X1 U5056 ( .A1(n4459), .A2(n4458), .A3(n4457), .A4(n4456), .ZN(n4465)
         );
  AOI22_X1 U5057 ( .A1(n5077), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n5079), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4463) );
  AOI22_X1 U5058 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n3853), .B1(n5076), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4462) );
  AOI22_X1 U5059 ( .A1(n3434), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5078), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4461) );
  AOI22_X1 U5060 ( .A1(n5068), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4460) );
  NAND4_X1 U5061 ( .A1(n4463), .A2(n4462), .A3(n4461), .A4(n4460), .ZN(n4464)
         );
  NOR2_X1 U5062 ( .A1(n4465), .A2(n4464), .ZN(n4476) );
  XNOR2_X1 U5063 ( .A(n4475), .B(n4476), .ZN(n4469) );
  NAND2_X1 U5064 ( .A1(n6720), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4466)
         );
  NAND2_X1 U5065 ( .A1(n5141), .A2(n4466), .ZN(n4467) );
  AOI21_X1 U5066 ( .B1(n4154), .B2(EAX_REG_23__SCAN_IN), .A(n4467), .ZN(n4468)
         );
  OAI21_X1 U5067 ( .B1(n5134), .B2(n4469), .A(n4468), .ZN(n4474) );
  OR2_X1 U5068 ( .A1(n4471), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4472)
         );
  NAND2_X1 U5069 ( .A1(n4498), .A2(n4472), .ZN(n6411) );
  OR2_X1 U5070 ( .A1(n4476), .A2(n4475), .ZN(n5050) );
  AOI22_X1 U5071 ( .A1(n3434), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4480) );
  AOI22_X1 U5072 ( .A1(n5077), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n5068), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4479) );
  AOI22_X1 U5073 ( .A1(n5079), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5078), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4478) );
  AOI22_X1 U5074 ( .A1(n5087), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n5056), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4477) );
  NAND4_X1 U5075 ( .A1(n4480), .A2(n4479), .A3(n4478), .A4(n4477), .ZN(n4486)
         );
  AOI22_X1 U5076 ( .A1(n5051), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4484) );
  AOI22_X1 U5077 ( .A1(n5076), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4483) );
  AOI22_X1 U5078 ( .A1(n5075), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4482) );
  AOI22_X1 U5079 ( .A1(n5042), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4481) );
  NAND4_X1 U5080 ( .A1(n4484), .A2(n4483), .A3(n4482), .A4(n4481), .ZN(n4485)
         );
  NOR2_X1 U5081 ( .A1(n4486), .A2(n4485), .ZN(n5049) );
  INV_X1 U5082 ( .A(n5049), .ZN(n4487) );
  XNOR2_X1 U5083 ( .A(n5050), .B(n4487), .ZN(n4491) );
  XNOR2_X1 U5084 ( .A(n4498), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5744)
         );
  NAND2_X1 U5085 ( .A1(n4154), .A2(EAX_REG_24__SCAN_IN), .ZN(n4489) );
  NAND2_X1 U5086 ( .A1(n5220), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4488)
         );
  OAI211_X1 U5087 ( .C1(n5744), .C2(n5141), .A(n4489), .B(n4488), .ZN(n4490)
         );
  AOI21_X1 U5088 ( .B1(n5149), .B2(n4491), .A(n4490), .ZN(n5144) );
  INV_X1 U5089 ( .A(n5144), .ZN(n4492) );
  NAND2_X1 U5090 ( .A1(n3455), .A2(n4492), .ZN(n5166) );
  AND2_X1 U5091 ( .A1(n5235), .A2(n6461), .ZN(n4496) );
  NOR2_X1 U5092 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6150) );
  NAND3_X1 U5093 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), 
        .A3(n6150), .ZN(n6485) );
  NOR2_X1 U5094 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6475), .ZN(n4894) );
  NAND2_X1 U5095 ( .A1(n5154), .A2(n4894), .ZN(n6473) );
  INV_X1 U5096 ( .A(n4498), .ZN(n4499) );
  INV_X1 U5097 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5151) );
  INV_X1 U5098 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5272) );
  INV_X1 U5099 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4501) );
  XNOR2_X1 U5100 ( .A(n4502), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5681)
         );
  NOR2_X1 U5101 ( .A1(n5681), .A2(n6475), .ZN(n4503) );
  AND2_X1 U5102 ( .A1(n5411), .A2(n4504), .ZN(n4505) );
  NOR2_X1 U5103 ( .A1(n5176), .A2(n4505), .ZN(n5862) );
  INV_X1 U5104 ( .A(n5862), .ZN(n4507) );
  NAND2_X1 U5105 ( .A1(n6736), .A2(n6500), .ZN(n4514) );
  NAND3_X1 U5106 ( .A1(n5241), .A2(n4514), .A3(EBX_REG_31__SCAN_IN), .ZN(n4506) );
  OAI22_X1 U5107 ( .A1(n5188), .A2(n6391), .B1(n4507), .B2(n6390), .ZN(n4521)
         );
  AND2_X2 U5108 ( .A1(n6371), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6395) );
  INV_X1 U5109 ( .A(n6371), .ZN(n5386) );
  NAND2_X1 U5110 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .ZN(
        n5352) );
  INV_X1 U5111 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6268) );
  NOR2_X1 U5112 ( .A1(n5352), .A2(n6268), .ZN(n5330) );
  NAND2_X1 U5113 ( .A1(n5330), .A2(REIP_REG_18__SCAN_IN), .ZN(n6359) );
  INV_X1 U5114 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6157) );
  NOR2_X1 U5115 ( .A1(n6359), .A2(n6157), .ZN(n6373) );
  NAND2_X1 U5116 ( .A1(REIP_REG_12__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .ZN(
        n5371) );
  INV_X1 U5117 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6011) );
  NOR2_X1 U5118 ( .A1(n5371), .A2(n6011), .ZN(n5329) );
  NAND3_X1 U5119 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6373), .A3(n5329), .ZN(
        n6385) );
  NAND2_X1 U5120 ( .A1(REIP_REG_6__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .ZN(
        n6338) );
  INV_X1 U5121 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6001) );
  NOR2_X1 U5122 ( .A1(n6338), .A2(n6001), .ZN(n4864) );
  INV_X1 U5123 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6309) );
  INV_X1 U5124 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6308) );
  NOR2_X1 U5125 ( .A1(n6309), .A2(n6308), .ZN(n4868) );
  INV_X1 U5126 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6003) );
  INV_X1 U5127 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6255) );
  INV_X1 U5128 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6225) );
  NOR3_X1 U5129 ( .A1(n6003), .A2(n6255), .A3(n6225), .ZN(n4947) );
  NAND2_X1 U5130 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .ZN(
        n5385) );
  INV_X1 U5131 ( .A(REIP_REG_3__SCAN_IN), .ZN(n5993) );
  NOR2_X1 U5132 ( .A1(n5385), .A2(n5993), .ZN(n6295) );
  NAND4_X1 U5133 ( .A1(n4864), .A2(n4868), .A3(n4947), .A4(n6295), .ZN(n5324)
         );
  NOR2_X1 U5134 ( .A1(n6385), .A2(n5324), .ZN(n6372) );
  NAND4_X1 U5135 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_23__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n6372), .ZN(n5181) );
  NAND2_X1 U5136 ( .A1(n4564), .A2(n5242), .ZN(n4508) );
  NAND2_X1 U5137 ( .A1(n3687), .A2(n4508), .ZN(n4510) );
  INV_X1 U5138 ( .A(n4514), .ZN(n4509) );
  NAND2_X1 U5139 ( .A1(n4510), .A2(n4509), .ZN(n4511) );
  NAND2_X1 U5140 ( .A1(n5249), .A2(n6371), .ZN(n6304) );
  OAI21_X1 U5141 ( .B1(n5386), .B2(n5181), .A(n6304), .ZN(n6423) );
  INV_X1 U5142 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U5143 ( .A1(n6296), .A2(n6023), .ZN(n5179) );
  OAI22_X1 U5144 ( .A1(n6423), .A2(n6023), .B1(n5181), .B2(n5179), .ZN(n4512)
         );
  AOI21_X1 U5145 ( .B1(PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n6395), .A(n4512), 
        .ZN(n4519) );
  AND2_X1 U5146 ( .A1(n5681), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4513) );
  NAND2_X1 U5147 ( .A1(n6397), .A2(n5744), .ZN(n4518) );
  NOR2_X1 U5148 ( .A1(n6143), .A2(n4514), .ZN(n6464) );
  NOR2_X1 U5149 ( .A1(n4835), .A2(n6464), .ZN(n5250) );
  INV_X1 U5150 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5398) );
  NAND3_X1 U5151 ( .A1(n4564), .A2(n4514), .A3(n5398), .ZN(n4515) );
  NAND2_X1 U5152 ( .A1(n4516), .A2(n4515), .ZN(n4517) );
  AND2_X2 U5153 ( .A1(n5250), .A2(n4517), .ZN(n6415) );
  NAND3_X1 U5154 ( .A1(n4519), .A2(n4518), .A3(n3456), .ZN(n4520) );
  NAND4_X1 U5155 ( .A1(n5692), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_28__SCAN_IN), .A4(INSTADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n4527) );
  AND2_X1 U5156 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U5157 ( .A1(n5834), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5007) );
  AND2_X1 U5158 ( .A1(n5692), .A2(n5007), .ZN(n4522) );
  NOR2_X1 U5159 ( .A1(n4523), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4524)
         );
  NOR2_X1 U5160 ( .A1(n5692), .A2(n4524), .ZN(n5686) );
  INV_X1 U5161 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5005) );
  INV_X1 U5162 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5691) );
  NAND4_X1 U5163 ( .A1(n5003), .A2(n5782), .A3(n5005), .A4(n5691), .ZN(n4526)
         );
  OAI21_X1 U5164 ( .B1(n4527), .B2(n5688), .A(n4526), .ZN(n4528) );
  XNOR2_X1 U5165 ( .A(n4528), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5685)
         );
  OR2_X1 U5166 ( .A1(n4547), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4530)
         );
  INV_X1 U5167 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4529) );
  NAND2_X1 U5168 ( .A1(n5241), .A2(n4529), .ZN(n4532) );
  NAND2_X1 U5169 ( .A1(n4530), .A2(n4532), .ZN(n5010) );
  MUX2_X1 U5170 ( .A(n5010), .B(n4532), .S(n4531), .Z(n5270) );
  NOR2_X4 U5171 ( .A1(n5271), .A2(n5270), .ZN(n5269) );
  AOI22_X1 U5172 ( .A1(n4547), .A2(EBX_REG_30__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n3687), .ZN(n5012) );
  OAI22_X1 U5173 ( .A1(n4547), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n3687), .ZN(n4535) );
  INV_X1 U5174 ( .A(n5243), .ZN(n4537) );
  NAND2_X1 U5175 ( .A1(n4537), .A2(n6280), .ZN(n4543) );
  INV_X1 U5176 ( .A(n5007), .ZN(n4538) );
  OAI21_X1 U5177 ( .B1(n4538), .B2(n5917), .A(n5839), .ZN(n5009) );
  INV_X1 U5178 ( .A(n5009), .ZN(n4539) );
  OAI21_X1 U5179 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5917), .A(n4539), 
        .ZN(n4541) );
  AND2_X1 U5180 ( .A1(n6277), .A2(REIP_REG_31__SCAN_IN), .ZN(n5679) );
  NOR4_X1 U5181 ( .A1(n5843), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5005), 
        .A4(n5007), .ZN(n4540) );
  AOI211_X1 U5182 ( .C1(n4541), .C2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n5679), .B(n4540), .ZN(n4542) );
  OAI211_X1 U5183 ( .C1(n5685), .C2(n6223), .A(n4543), .B(n4542), .ZN(U2987)
         );
  INV_X1 U5184 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6511) );
  INV_X1 U5185 ( .A(n4618), .ZN(n4545) );
  INV_X1 U5186 ( .A(n6137), .ZN(n4544) );
  OAI211_X1 U5187 ( .C1(n4546), .C2(n6511), .A(n4545), .B(n4544), .ZN(U2788)
         );
  OR2_X1 U5188 ( .A1(n4547), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4549)
         );
  NAND2_X1 U5189 ( .A1(n4549), .A2(n4548), .ZN(n6287) );
  NAND2_X1 U5190 ( .A1(n5239), .A2(n4550), .ZN(n4554) );
  INV_X1 U5191 ( .A(n4551), .ZN(n4552) );
  NAND4_X1 U5192 ( .A1(n4552), .A2(n6872), .A3(n7000), .A4(n4595), .ZN(n4663)
         );
  OR2_X1 U5193 ( .A1(n4663), .A2(n3687), .ZN(n4553) );
  NAND2_X1 U5194 ( .A1(n4554), .A2(n4553), .ZN(n4555) );
  XNOR2_X1 U5195 ( .A(n4557), .B(n4556), .ZN(n6077) );
  INV_X1 U5196 ( .A(n6077), .ZN(n6292) );
  OAI222_X1 U5197 ( .A1(n6287), .A2(n6060), .B1(n6061), .B2(n6292), .C1(n3694), 
        .C2(n6075), .ZN(U2859) );
  OAI21_X1 U5198 ( .B1(n4560), .B2(n4559), .A(n4558), .ZN(n6082) );
  XNOR2_X1 U5199 ( .A(n4827), .B(n5241), .ZN(n5928) );
  AOI22_X1 U5200 ( .A1(n6071), .A2(n5928), .B1(EBX_REG_1__SCAN_IN), .B2(n5445), 
        .ZN(n4561) );
  OAI21_X1 U5201 ( .B1(n6061), .B2(n6082), .A(n4561), .ZN(U2858) );
  INV_X1 U5202 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4566) );
  OAI21_X1 U5203 ( .B1(n5207), .B2(n6465), .A(n5242), .ZN(n4563) );
  NAND2_X1 U5204 ( .A1(n5956), .A2(n4564), .ZN(n4720) );
  AND2_X2 U5205 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4894), .ZN(n6154) );
  NOR2_X4 U5206 ( .A1(n6154), .A2(n5956), .ZN(n5969) );
  AOI22_X1 U5207 ( .A1(n6154), .A2(UWORD_REG_7__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4565) );
  OAI21_X1 U5208 ( .B1(n4566), .B2(n4720), .A(n4565), .ZN(U2900) );
  INV_X1 U5209 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4568) );
  AOI22_X1 U5210 ( .A1(n6154), .A2(UWORD_REG_5__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4567) );
  OAI21_X1 U5211 ( .B1(n4568), .B2(n4720), .A(n4567), .ZN(U2902) );
  INV_X1 U5212 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4570) );
  AOI22_X1 U5213 ( .A1(n6154), .A2(UWORD_REG_10__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4569) );
  OAI21_X1 U5214 ( .B1(n4570), .B2(n4720), .A(n4569), .ZN(U2897) );
  INV_X1 U5215 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4572) );
  AOI22_X1 U5216 ( .A1(n6154), .A2(UWORD_REG_9__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4571) );
  OAI21_X1 U5217 ( .B1(n4572), .B2(n4720), .A(n4571), .ZN(U2898) );
  INV_X1 U5218 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4574) );
  AOI22_X1 U5219 ( .A1(n6154), .A2(UWORD_REG_4__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4573) );
  OAI21_X1 U5220 ( .B1(n4574), .B2(n4720), .A(n4573), .ZN(U2903) );
  INV_X1 U5221 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4576) );
  AOI22_X1 U5222 ( .A1(n6154), .A2(UWORD_REG_8__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4575) );
  OAI21_X1 U5223 ( .B1(n4576), .B2(n4720), .A(n4575), .ZN(U2899) );
  INV_X1 U5224 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4578) );
  AOI22_X1 U5225 ( .A1(n6154), .A2(UWORD_REG_6__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4577) );
  OAI21_X1 U5226 ( .B1(n4578), .B2(n4720), .A(n4577), .ZN(U2901) );
  NOR2_X1 U5227 ( .A1(n6744), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6543) );
  OAI22_X1 U5228 ( .A1(n5207), .A2(n4579), .B1(n4495), .B2(n5242), .ZN(n4580)
         );
  INV_X1 U5229 ( .A(n4580), .ZN(n4581) );
  NAND2_X1 U5230 ( .A1(n4582), .A2(n4581), .ZN(n4590) );
  OR2_X1 U5231 ( .A1(n5239), .A2(n4600), .ZN(n4585) );
  OR2_X1 U5232 ( .A1(n4135), .A2(n4583), .ZN(n4584) );
  INV_X1 U5233 ( .A(n4665), .ZN(n4589) );
  AND2_X1 U5234 ( .A1(n6545), .A2(n4586), .ZN(n4833) );
  NAND2_X1 U5235 ( .A1(n4833), .A2(n6790), .ZN(n4587) );
  NAND4_X1 U5236 ( .A1(n4590), .A2(n4589), .A3(n4588), .A4(n4587), .ZN(n4685)
         );
  INV_X1 U5237 ( .A(n4685), .ZN(n6436) );
  INV_X1 U5238 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6451) );
  NOR2_X1 U5239 ( .A1(n6720), .A2(n6475), .ZN(n6472) );
  NAND2_X1 U5240 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6472), .ZN(n6476) );
  OAI22_X1 U5241 ( .A1(n6436), .A2(n6487), .B1(n6451), .B2(n6476), .ZN(n6428)
         );
  NOR2_X1 U5242 ( .A1(n6543), .A2(n6428), .ZN(n5948) );
  AOI21_X1 U5243 ( .B1(n6430), .B2(n5086), .A(n4591), .ZN(n4609) );
  INV_X1 U5244 ( .A(n4592), .ZN(n5934) );
  NAND2_X1 U5245 ( .A1(n5934), .A2(n5205), .ZN(n5941) );
  NAND2_X1 U5246 ( .A1(n6430), .A2(n5941), .ZN(n5212) );
  NAND2_X1 U5247 ( .A1(n5212), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4608) );
  INV_X1 U5248 ( .A(n4594), .ZN(n4599) );
  INV_X1 U5249 ( .A(n4595), .ZN(n4596) );
  AND3_X1 U5250 ( .A1(n4597), .A2(n4596), .A3(n4135), .ZN(n4598) );
  NAND2_X1 U5251 ( .A1(n4599), .A2(n4598), .ZN(n5939) );
  NAND2_X1 U5252 ( .A1(n6630), .A2(n5939), .ZN(n4606) );
  NAND2_X1 U5253 ( .A1(n5228), .A2(n4600), .ZN(n4681) );
  NAND2_X1 U5254 ( .A1(n5934), .A2(n5218), .ZN(n4678) );
  XNOR2_X1 U5255 ( .A(n4601), .B(n4678), .ZN(n4604) );
  XNOR2_X1 U5256 ( .A(n4602), .B(n4601), .ZN(n4603) );
  AOI22_X1 U5257 ( .A1(n4681), .A2(n4604), .B1(n5207), .B2(n4603), .ZN(n4605)
         );
  NAND2_X1 U5258 ( .A1(n4606), .A2(n4605), .ZN(n4675) );
  NAND3_X1 U5259 ( .A1(n6430), .A2(n6469), .A3(n4675), .ZN(n4607) );
  OAI211_X1 U5260 ( .C1(n4609), .C2(n6478), .A(n4608), .B(n4607), .ZN(U3456)
         );
  CLKBUF_X1 U5261 ( .A(n4611), .Z(n4672) );
  NAND2_X1 U5262 ( .A1(n4672), .A2(n4612), .ZN(n4613) );
  AND2_X1 U5263 ( .A1(n4610), .A2(n4613), .ZN(n5392) );
  INV_X1 U5264 ( .A(n5392), .ZN(n4669) );
  OR2_X1 U5265 ( .A1(n5195), .A2(n4615), .ZN(n4616) );
  AND2_X1 U5266 ( .A1(n4651), .A2(n4616), .ZN(n5394) );
  AOI22_X1 U5267 ( .A1(n6071), .A2(n5394), .B1(EBX_REG_3__SCAN_IN), .B2(n5445), 
        .ZN(n4617) );
  OAI21_X1 U5268 ( .B1(n4669), .B2(n6061), .A(n4617), .ZN(U2856) );
  NAND2_X1 U5269 ( .A1(n4618), .A2(n6500), .ZN(n4620) );
  NAND2_X1 U5270 ( .A1(n4728), .A2(DATAI_4_), .ZN(n4623) );
  INV_X2 U5271 ( .A(n4735), .ZN(n4758) );
  AOI22_X1 U5272 ( .A1(n4758), .A2(EAX_REG_20__SCAN_IN), .B1(n4721), .B2(
        UWORD_REG_4__SCAN_IN), .ZN(n4621) );
  NAND2_X1 U5273 ( .A1(n4623), .A2(n4621), .ZN(U2928) );
  AOI22_X1 U5274 ( .A1(n4758), .A2(EAX_REG_4__SCAN_IN), .B1(n4721), .B2(
        LWORD_REG_4__SCAN_IN), .ZN(n4622) );
  NAND2_X1 U5275 ( .A1(n4623), .A2(n4622), .ZN(U2943) );
  NAND2_X1 U5276 ( .A1(n4728), .A2(DATAI_2_), .ZN(n4749) );
  AOI22_X1 U5277 ( .A1(n4758), .A2(EAX_REG_2__SCAN_IN), .B1(n4721), .B2(
        LWORD_REG_2__SCAN_IN), .ZN(n4624) );
  NAND2_X1 U5278 ( .A1(n4749), .A2(n4624), .ZN(U2941) );
  NAND2_X1 U5279 ( .A1(n4728), .A2(DATAI_1_), .ZN(n4732) );
  AOI22_X1 U5280 ( .A1(n4758), .A2(EAX_REG_1__SCAN_IN), .B1(n4721), .B2(
        LWORD_REG_1__SCAN_IN), .ZN(n4625) );
  NAND2_X1 U5281 ( .A1(n4732), .A2(n4625), .ZN(U2940) );
  NAND2_X1 U5282 ( .A1(n4728), .A2(DATAI_0_), .ZN(n4751) );
  AOI22_X1 U5283 ( .A1(n4758), .A2(EAX_REG_0__SCAN_IN), .B1(n4721), .B2(
        LWORD_REG_0__SCAN_IN), .ZN(n4626) );
  NAND2_X1 U5284 ( .A1(n4751), .A2(n4626), .ZN(U2939) );
  INV_X1 U5285 ( .A(DATAI_14_), .ZN(n5676) );
  OR2_X1 U5286 ( .A1(n4760), .A2(n5676), .ZN(n4745) );
  AOI22_X1 U5287 ( .A1(n4758), .A2(EAX_REG_30__SCAN_IN), .B1(n4721), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n4627) );
  NAND2_X1 U5288 ( .A1(n4745), .A2(n4627), .ZN(U2938) );
  NAND2_X1 U5289 ( .A1(n4728), .A2(DATAI_3_), .ZN(n4723) );
  AOI22_X1 U5290 ( .A1(n4758), .A2(EAX_REG_3__SCAN_IN), .B1(n4721), .B2(
        LWORD_REG_3__SCAN_IN), .ZN(n4628) );
  NAND2_X1 U5291 ( .A1(n4723), .A2(n4628), .ZN(U2942) );
  NAND2_X1 U5292 ( .A1(n4728), .A2(DATAI_12_), .ZN(n4747) );
  AOI22_X1 U5293 ( .A1(n4758), .A2(EAX_REG_28__SCAN_IN), .B1(n4721), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n4629) );
  NAND2_X1 U5294 ( .A1(n4747), .A2(n4629), .ZN(U2936) );
  NAND2_X1 U5295 ( .A1(n4728), .A2(DATAI_11_), .ZN(n4757) );
  AOI22_X1 U5296 ( .A1(n4758), .A2(EAX_REG_27__SCAN_IN), .B1(n4721), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n4630) );
  NAND2_X1 U5297 ( .A1(n4757), .A2(n4630), .ZN(U2935) );
  NAND2_X1 U5298 ( .A1(n4728), .A2(DATAI_10_), .ZN(n4739) );
  AOI22_X1 U5299 ( .A1(n4758), .A2(EAX_REG_26__SCAN_IN), .B1(n4721), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n4631) );
  NAND2_X1 U5300 ( .A1(n4739), .A2(n4631), .ZN(U2934) );
  NAND2_X1 U5301 ( .A1(n4728), .A2(DATAI_9_), .ZN(n4755) );
  AOI22_X1 U5302 ( .A1(n4758), .A2(EAX_REG_25__SCAN_IN), .B1(n4721), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n4632) );
  NAND2_X1 U5303 ( .A1(n4755), .A2(n4632), .ZN(U2933) );
  NAND2_X1 U5304 ( .A1(n4728), .A2(DATAI_13_), .ZN(n4734) );
  AOI22_X1 U5305 ( .A1(n4758), .A2(EAX_REG_29__SCAN_IN), .B1(n4721), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n4633) );
  NAND2_X1 U5306 ( .A1(n4734), .A2(n4633), .ZN(U2937) );
  INV_X1 U5307 ( .A(DATAI_6_), .ZN(n4674) );
  OR2_X1 U5308 ( .A1(n4760), .A2(n4674), .ZN(n4726) );
  AOI22_X1 U5309 ( .A1(n4758), .A2(EAX_REG_22__SCAN_IN), .B1(n4721), .B2(
        UWORD_REG_6__SCAN_IN), .ZN(n4634) );
  NAND2_X1 U5310 ( .A1(n4726), .A2(n4634), .ZN(U2930) );
  INV_X1 U5311 ( .A(DATAI_8_), .ZN(n4818) );
  OR2_X1 U5312 ( .A1(n4760), .A2(n4818), .ZN(n4753) );
  AOI22_X1 U5313 ( .A1(n4758), .A2(EAX_REG_24__SCAN_IN), .B1(n4721), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n4635) );
  NAND2_X1 U5314 ( .A1(n4753), .A2(n4635), .ZN(U2932) );
  INV_X1 U5315 ( .A(n6222), .ZN(n6196) );
  OAI21_X1 U5316 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n6217), .A(n6196), 
        .ZN(n5923) );
  OAI22_X1 U5317 ( .A1(n5923), .A2(n4637), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n4636), .ZN(n4643) );
  NOR2_X1 U5318 ( .A1(n4638), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4639)
         );
  OR2_X1 U5319 ( .A1(n5925), .A2(n4639), .ZN(n6081) );
  INV_X1 U5320 ( .A(REIP_REG_0__SCAN_IN), .ZN(n4640) );
  OAI22_X1 U5321 ( .A1(n6223), .A2(n6081), .B1(n6269), .B2(n4640), .ZN(n4641)
         );
  INV_X1 U5322 ( .A(n4641), .ZN(n4642) );
  OAI211_X1 U5323 ( .C1(n6227), .C2(n6287), .A(n4643), .B(n4642), .ZN(U3018)
         );
  AND2_X1 U5324 ( .A1(n4610), .A2(n4644), .ZN(n4647) );
  CLKBUF_X1 U5325 ( .A(n4645), .Z(n4646) );
  OR2_X1 U5326 ( .A1(n4647), .A2(n4646), .ZN(n6300) );
  XNOR2_X1 U5327 ( .A(n4651), .B(n4650), .ZN(n4849) );
  INV_X1 U5328 ( .A(n4849), .ZN(n6293) );
  AOI22_X1 U5329 ( .A1(n6071), .A2(n6293), .B1(EBX_REG_4__SCAN_IN), .B2(n5445), 
        .ZN(n4648) );
  OAI21_X1 U5330 ( .B1(n6300), .B2(n6061), .A(n4648), .ZN(U2855) );
  OAI21_X1 U5331 ( .B1(n4651), .B2(n4650), .A(n4649), .ZN(n4652) );
  AND2_X1 U5332 ( .A1(n4652), .A2(n4660), .ZN(n4782) );
  INV_X1 U5333 ( .A(n4782), .ZN(n6313) );
  INV_X1 U5334 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4656) );
  CLKBUF_X1 U5335 ( .A(n4653), .Z(n4658) );
  OR2_X1 U5336 ( .A1(n4646), .A2(n4654), .ZN(n4655) );
  NAND2_X1 U5337 ( .A1(n4658), .A2(n4655), .ZN(n6317) );
  OAI222_X1 U5338 ( .A1(n6313), .A2(n6060), .B1(n4656), .B2(n6075), .C1(n6317), 
        .C2(n6061), .ZN(U2854) );
  XNOR2_X1 U5339 ( .A(n4658), .B(n4657), .ZN(n6326) );
  AND2_X1 U5340 ( .A1(n4660), .A2(n4659), .ZN(n4661) );
  NOR2_X1 U5341 ( .A1(n4840), .A2(n4661), .ZN(n6322) );
  AOI22_X1 U5342 ( .A1(n6071), .A2(n6322), .B1(EBX_REG_6__SCAN_IN), .B2(n5445), 
        .ZN(n4662) );
  OAI21_X1 U5343 ( .B1(n6326), .B2(n6061), .A(n4662), .ZN(U2853) );
  INV_X1 U5344 ( .A(n5240), .ZN(n5238) );
  NOR2_X1 U5345 ( .A1(n4663), .A2(n5238), .ZN(n4664) );
  INV_X1 U5346 ( .A(n4668), .ZN(n4667) );
  INV_X1 U5347 ( .A(DATAI_4_), .ZN(n5497) );
  INV_X1 U5348 ( .A(EAX_REG_4__SCAN_IN), .ZN(n5966) );
  OAI222_X1 U5349 ( .A1(n6300), .A2(n5678), .B1(n5677), .B2(n5497), .C1(n6514), 
        .C2(n5966), .ZN(U2887) );
  INV_X1 U5350 ( .A(DATAI_0_), .ZN(n5614) );
  INV_X1 U5351 ( .A(EAX_REG_0__SCAN_IN), .ZN(n5958) );
  OAI222_X1 U5352 ( .A1(n5678), .A2(n6292), .B1(n5677), .B2(n5614), .C1(n6514), 
        .C2(n5958), .ZN(U2891) );
  INV_X1 U5353 ( .A(DATAI_5_), .ZN(n4736) );
  INV_X1 U5354 ( .A(EAX_REG_5__SCAN_IN), .ZN(n5968) );
  OAI222_X1 U5355 ( .A1(n6317), .A2(n5678), .B1(n5677), .B2(n4736), .C1(n6514), 
        .C2(n5968), .ZN(U2886) );
  INV_X1 U5356 ( .A(DATAI_3_), .ZN(n5604) );
  INV_X1 U5357 ( .A(EAX_REG_3__SCAN_IN), .ZN(n5964) );
  OAI222_X1 U5358 ( .A1(n4669), .A2(n5678), .B1(n5677), .B2(n5604), .C1(n6514), 
        .C2(n5964), .ZN(U2888) );
  INV_X1 U5359 ( .A(DATAI_1_), .ZN(n5612) );
  INV_X1 U5360 ( .A(EAX_REG_1__SCAN_IN), .ZN(n5960) );
  OAI222_X1 U5361 ( .A1(n6082), .A2(n5678), .B1(n5677), .B2(n5612), .C1(n6514), 
        .C2(n5960), .ZN(U2890) );
  INV_X1 U5362 ( .A(n4670), .ZN(n4671) );
  NAND2_X1 U5363 ( .A1(n4671), .A2(n4558), .ZN(n4673) );
  NAND2_X1 U5364 ( .A1(n4673), .A2(n4672), .ZN(n6091) );
  INV_X1 U5365 ( .A(DATAI_2_), .ZN(n5603) );
  INV_X1 U5366 ( .A(EAX_REG_2__SCAN_IN), .ZN(n5962) );
  OAI222_X1 U5367 ( .A1(n6091), .A2(n5678), .B1(n5677), .B2(n5603), .C1(n6514), 
        .C2(n5962), .ZN(U2889) );
  OAI222_X1 U5368 ( .A1(n5678), .A2(n6326), .B1(n5677), .B2(n4674), .C1(n6514), 
        .C2(n4727), .ZN(U2885) );
  INV_X1 U5369 ( .A(n6630), .ZN(n6698) );
  MUX2_X1 U5370 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n4675), .S(n4685), 
        .Z(n6444) );
  INV_X1 U5371 ( .A(n5939), .ZN(n4683) );
  OAI21_X1 U5372 ( .B1(n5934), .B2(n5218), .A(n4678), .ZN(n4680) );
  XNOR2_X1 U5373 ( .A(n3467), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4679)
         );
  AOI22_X1 U5374 ( .A1(n4681), .A2(n4680), .B1(n5207), .B2(n4679), .ZN(n4682)
         );
  OAI21_X1 U5375 ( .B1(n4677), .B2(n4683), .A(n4682), .ZN(n5216) );
  NAND2_X1 U5376 ( .A1(n4685), .A2(n5216), .ZN(n4684) );
  OAI21_X1 U5377 ( .B1(n4685), .B2(n5218), .A(n4684), .ZN(n6439) );
  NAND3_X1 U5378 ( .A1(n6444), .A2(n6475), .A3(n6439), .ZN(n4689) );
  NOR2_X1 U5379 ( .A1(FLUSH_REG_SCAN_IN), .A2(n6475), .ZN(n4686) );
  NAND2_X1 U5380 ( .A1(n4687), .A2(n4686), .ZN(n4688) );
  NAND2_X1 U5381 ( .A1(n4689), .A2(n4688), .ZN(n6447) );
  INV_X1 U5382 ( .A(n4690), .ZN(n5942) );
  NAND2_X1 U5383 ( .A1(n6447), .A2(n5942), .ZN(n4699) );
  MUX2_X1 U5384 ( .A(n6436), .B(n6451), .S(STATE2_REG_1__SCAN_IN), .Z(n4698)
         );
  INV_X1 U5385 ( .A(n4691), .ZN(n4692) );
  NOR2_X1 U5386 ( .A1(n4693), .A2(n4692), .ZN(n4695) );
  XNOR2_X1 U5387 ( .A(n4695), .B(n4694), .ZN(n6426) );
  NOR2_X1 U5388 ( .A1(n4135), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4696) );
  AND2_X1 U5389 ( .A1(n6426), .A2(n4696), .ZN(n4697) );
  AOI21_X1 U5390 ( .B1(n4698), .B2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(n4697), 
        .ZN(n6456) );
  NAND2_X1 U5391 ( .A1(n4699), .A2(n6456), .ZN(n4763) );
  INV_X1 U5392 ( .A(n6476), .ZN(n6148) );
  OAI21_X1 U5393 ( .B1(n4763), .B2(FLUSH_REG_SCAN_IN), .A(n6148), .ZN(n4700)
         );
  INV_X1 U5394 ( .A(n5953), .ZN(n4787) );
  OAI21_X1 U5395 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6475), .A(n4787), .ZN(
        n4804) );
  INV_X1 U5396 ( .A(n6659), .ZN(n6710) );
  NOR2_X1 U5397 ( .A1(n5953), .A2(n6710), .ZN(n4784) );
  INV_X1 U5398 ( .A(n6666), .ZN(n6695) );
  NOR2_X1 U5399 ( .A1(n3436), .A2(n6736), .ZN(n4703) );
  NAND3_X1 U5400 ( .A1(n4703), .A2(n6566), .A3(n6640), .ZN(n6572) );
  NOR2_X1 U5401 ( .A1(n3436), .A2(n6566), .ZN(n6641) );
  NAND2_X1 U5402 ( .A1(n6663), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4785) );
  INV_X1 U5403 ( .A(n4785), .ZN(n6585) );
  NAND2_X1 U5404 ( .A1(n6641), .A2(n6585), .ZN(n6628) );
  OAI211_X1 U5405 ( .C1(n6695), .C2(n4703), .A(n6572), .B(n6628), .ZN(n4704)
         );
  AOI22_X1 U5406 ( .A1(n4784), .A2(n4704), .B1(n5953), .B2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4705) );
  OAI21_X1 U5407 ( .B1(n6698), .B2(n4804), .A(n4705), .ZN(U3462) );
  INV_X1 U5408 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4707) );
  AOI22_X1 U5409 ( .A1(n6154), .A2(UWORD_REG_14__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4706) );
  OAI21_X1 U5410 ( .B1(n4707), .B2(n4720), .A(n4706), .ZN(U2893) );
  INV_X1 U5411 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4709) );
  AOI22_X1 U5412 ( .A1(n6154), .A2(UWORD_REG_0__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4708) );
  OAI21_X1 U5413 ( .B1(n4709), .B2(n4720), .A(n4708), .ZN(U2907) );
  INV_X1 U5414 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4711) );
  AOI22_X1 U5415 ( .A1(n6154), .A2(UWORD_REG_2__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4710) );
  OAI21_X1 U5416 ( .B1(n4711), .B2(n4720), .A(n4710), .ZN(U2905) );
  INV_X1 U5417 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4713) );
  AOI22_X1 U5418 ( .A1(n6154), .A2(UWORD_REG_13__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4712) );
  OAI21_X1 U5419 ( .B1(n4713), .B2(n4720), .A(n4712), .ZN(U2894) );
  INV_X1 U5420 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4715) );
  AOI22_X1 U5421 ( .A1(n6154), .A2(UWORD_REG_12__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4714) );
  OAI21_X1 U5422 ( .B1(n4715), .B2(n4720), .A(n4714), .ZN(U2895) );
  INV_X1 U5423 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4717) );
  AOI22_X1 U5424 ( .A1(n6154), .A2(UWORD_REG_11__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4716) );
  OAI21_X1 U5425 ( .B1(n4717), .B2(n4720), .A(n4716), .ZN(U2896) );
  AOI22_X1 U5426 ( .A1(n6154), .A2(UWORD_REG_3__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4718) );
  OAI21_X1 U5427 ( .B1(n4724), .B2(n4720), .A(n4718), .ZN(U2904) );
  INV_X1 U5428 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6515) );
  AOI22_X1 U5429 ( .A1(n6154), .A2(UWORD_REG_1__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4719) );
  OAI21_X1 U5430 ( .B1(n6515), .B2(n4720), .A(n4719), .ZN(U2906) );
  NAND2_X1 U5431 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n4721), .ZN(n4722) );
  OAI211_X1 U5432 ( .C1(n4735), .C2(n4724), .A(n4723), .B(n4722), .ZN(U2927)
         );
  NAND2_X1 U5433 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n4721), .ZN(n4725) );
  OAI211_X1 U5434 ( .C1(n4735), .C2(n4727), .A(n4726), .B(n4725), .ZN(U2945)
         );
  NAND2_X1 U5435 ( .A1(n4728), .A2(DATAI_7_), .ZN(n4743) );
  NAND2_X1 U5436 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n4721), .ZN(n4729) );
  OAI211_X1 U5437 ( .C1(n4735), .C2(n4730), .A(n4743), .B(n4729), .ZN(U2946)
         );
  NAND2_X1 U5438 ( .A1(UWORD_REG_1__SCAN_IN), .A2(n4721), .ZN(n4731) );
  OAI211_X1 U5439 ( .C1(n4735), .C2(n6515), .A(n4732), .B(n4731), .ZN(U2925)
         );
  INV_X1 U5440 ( .A(EAX_REG_13__SCAN_IN), .ZN(n5983) );
  NAND2_X1 U5441 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n4721), .ZN(n4733) );
  OAI211_X1 U5442 ( .C1(n4735), .C2(n5983), .A(n4734), .B(n4733), .ZN(U2952)
         );
  OR2_X1 U5443 ( .A1(n4760), .A2(n4736), .ZN(n4741) );
  AOI22_X1 U5444 ( .A1(n4758), .A2(EAX_REG_5__SCAN_IN), .B1(n4721), .B2(
        LWORD_REG_5__SCAN_IN), .ZN(n4737) );
  NAND2_X1 U5445 ( .A1(n4741), .A2(n4737), .ZN(U2944) );
  AOI22_X1 U5446 ( .A1(n4758), .A2(EAX_REG_10__SCAN_IN), .B1(n4721), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n4738) );
  NAND2_X1 U5447 ( .A1(n4739), .A2(n4738), .ZN(U2949) );
  AOI22_X1 U5448 ( .A1(n4758), .A2(EAX_REG_21__SCAN_IN), .B1(n4721), .B2(
        UWORD_REG_5__SCAN_IN), .ZN(n4740) );
  NAND2_X1 U5449 ( .A1(n4741), .A2(n4740), .ZN(U2929) );
  AOI22_X1 U5450 ( .A1(n4758), .A2(EAX_REG_23__SCAN_IN), .B1(n4721), .B2(
        UWORD_REG_7__SCAN_IN), .ZN(n4742) );
  NAND2_X1 U5451 ( .A1(n4743), .A2(n4742), .ZN(U2931) );
  AOI22_X1 U5452 ( .A1(n4758), .A2(EAX_REG_14__SCAN_IN), .B1(n4721), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n4744) );
  NAND2_X1 U5453 ( .A1(n4745), .A2(n4744), .ZN(U2953) );
  AOI22_X1 U5454 ( .A1(n4758), .A2(EAX_REG_12__SCAN_IN), .B1(n4721), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n4746) );
  NAND2_X1 U5455 ( .A1(n4747), .A2(n4746), .ZN(U2951) );
  AOI22_X1 U5456 ( .A1(n4758), .A2(EAX_REG_18__SCAN_IN), .B1(n4721), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n4748) );
  NAND2_X1 U5457 ( .A1(n4749), .A2(n4748), .ZN(U2926) );
  AOI22_X1 U5458 ( .A1(n4758), .A2(EAX_REG_16__SCAN_IN), .B1(n4721), .B2(
        UWORD_REG_0__SCAN_IN), .ZN(n4750) );
  NAND2_X1 U5459 ( .A1(n4751), .A2(n4750), .ZN(U2924) );
  AOI22_X1 U5460 ( .A1(n4758), .A2(EAX_REG_8__SCAN_IN), .B1(n4721), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n4752) );
  NAND2_X1 U5461 ( .A1(n4753), .A2(n4752), .ZN(U2947) );
  AOI22_X1 U5462 ( .A1(n4758), .A2(EAX_REG_9__SCAN_IN), .B1(n4721), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n4754) );
  NAND2_X1 U5463 ( .A1(n4755), .A2(n4754), .ZN(U2948) );
  AOI22_X1 U5464 ( .A1(n4758), .A2(EAX_REG_11__SCAN_IN), .B1(n4721), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n4756) );
  NAND2_X1 U5465 ( .A1(n4757), .A2(n4756), .ZN(U2950) );
  INV_X1 U5466 ( .A(DATAI_15_), .ZN(n5674) );
  AOI22_X1 U5467 ( .A1(n4758), .A2(EAX_REG_15__SCAN_IN), .B1(n4721), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n4759) );
  OAI21_X1 U5468 ( .B1(n4760), .B2(n5674), .A(n4759), .ZN(U2954) );
  INV_X1 U5469 ( .A(n6472), .ZN(n4762) );
  OR2_X1 U5470 ( .A1(n4763), .A2(n4762), .ZN(n6483) );
  NAND2_X1 U5471 ( .A1(n5953), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4764) );
  OAI21_X1 U5472 ( .B1(n5953), .B2(n6483), .A(n4764), .ZN(n4765) );
  AOI21_X1 U5473 ( .B1(n4784), .B2(n6723), .A(n4765), .ZN(n4766) );
  OAI21_X1 U5474 ( .B1(n6629), .B2(n4804), .A(n4766), .ZN(U3465) );
  NAND2_X1 U5475 ( .A1(n4768), .A2(n4767), .ZN(n4770) );
  XNOR2_X1 U5476 ( .A(n4770), .B(n4769), .ZN(n4904) );
  NAND2_X1 U5477 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4771) );
  AOI21_X1 U5478 ( .B1(n6199), .B2(n4771), .A(n6222), .ZN(n6193) );
  OAI21_X1 U5479 ( .B1(n6217), .B2(n6183), .A(n6193), .ZN(n4847) );
  NOR3_X1 U5480 ( .A1(n3700), .A2(n5929), .A3(n5905), .ZN(n4777) );
  OR2_X1 U5481 ( .A1(n5901), .A2(n4777), .ZN(n6200) );
  NAND2_X1 U5482 ( .A1(n6183), .A2(n6200), .ZN(n4850) );
  INV_X1 U5483 ( .A(n4850), .ZN(n4772) );
  AOI22_X1 U5484 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4847), .B1(n4772), 
        .B2(n4001), .ZN(n4774) );
  NOR2_X1 U5485 ( .A1(n6269), .A2(n5993), .ZN(n4900) );
  AOI21_X1 U5486 ( .B1(n6280), .B2(n5394), .A(n4900), .ZN(n4773) );
  OAI211_X1 U5487 ( .C1(n4904), .C2(n6223), .A(n4774), .B(n4773), .ZN(U3015)
         );
  XNOR2_X1 U5488 ( .A(n4775), .B(n4776), .ZN(n6096) );
  NAND2_X1 U5489 ( .A1(n6277), .A2(REIP_REG_5__SCAN_IN), .ZN(n6098) );
  INV_X1 U5490 ( .A(n6098), .ZN(n4781) );
  OAI211_X1 U5491 ( .C1(n4777), .C2(n5901), .A(n6183), .B(n4851), .ZN(n4779)
         );
  AOI21_X1 U5492 ( .B1(n6165), .B2(n4792), .A(n4847), .ZN(n4793) );
  AOI21_X1 U5493 ( .B1(n4779), .B2(n4778), .A(n4793), .ZN(n4780) );
  AOI211_X1 U5494 ( .C1(n6280), .C2(n4782), .A(n4781), .B(n4780), .ZN(n4783)
         );
  OAI21_X1 U5495 ( .B1(n6223), .B2(n6096), .A(n4783), .ZN(U3013) );
  INV_X1 U5496 ( .A(n4784), .ZN(n4801) );
  XNOR2_X1 U5497 ( .A(n3436), .B(n4785), .ZN(n4786) );
  OAI222_X1 U5498 ( .A1(n4804), .A2(n4677), .B1(n4787), .B2(n6649), .C1(n4801), 
        .C2(n4786), .ZN(U3463) );
  AND2_X1 U5499 ( .A1(n4790), .A2(n4789), .ZN(n4791) );
  XNOR2_X1 U5500 ( .A(n4788), .B(n4791), .ZN(n6102) );
  NOR2_X1 U5501 ( .A1(n4792), .A2(n4850), .ZN(n4795) );
  INV_X1 U5502 ( .A(n4793), .ZN(n4794) );
  MUX2_X1 U5503 ( .A(n4795), .B(n4794), .S(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .Z(n4796) );
  INV_X1 U5504 ( .A(n4796), .ZN(n4798) );
  AOI22_X1 U5505 ( .A1(n6280), .A2(n6322), .B1(n6277), .B2(REIP_REG_6__SCAN_IN), .ZN(n4797) );
  OAI211_X1 U5506 ( .C1(n6102), .C2(n6223), .A(n4798), .B(n4797), .ZN(U3012)
         );
  AOI211_X1 U5507 ( .C1(n6640), .C2(n6736), .A(n6585), .B(n4801), .ZN(n4802)
         );
  AOI21_X1 U5508 ( .B1(n5953), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n4802), 
        .ZN(n4803) );
  OAI21_X1 U5509 ( .B1(n6607), .B2(n4804), .A(n4803), .ZN(U3464) );
  INV_X1 U5510 ( .A(n4805), .ZN(n4810) );
  CLKBUF_X1 U5511 ( .A(n4806), .Z(n4807) );
  INV_X1 U5512 ( .A(n4807), .ZN(n4809) );
  AOI21_X1 U5513 ( .B1(n4810), .B2(n4809), .A(n4808), .ZN(n5383) );
  INV_X1 U5514 ( .A(n5383), .ZN(n4819) );
  OR2_X1 U5515 ( .A1(n4842), .A2(n4812), .ZN(n4813) );
  AND2_X1 U5516 ( .A1(n4811), .A2(n4813), .ZN(n6203) );
  AOI22_X1 U5517 ( .A1(n6071), .A2(n6203), .B1(EBX_REG_8__SCAN_IN), .B2(n5445), 
        .ZN(n4814) );
  OAI21_X1 U5518 ( .B1(n4819), .B2(n6061), .A(n4814), .ZN(U2851) );
  AND2_X1 U5519 ( .A1(n4816), .A2(n4815), .ZN(n4817) );
  NOR2_X1 U5520 ( .A1(n4807), .A2(n4817), .ZN(n6333) );
  INV_X1 U5521 ( .A(n6333), .ZN(n4843) );
  INV_X1 U5522 ( .A(DATAI_7_), .ZN(n5601) );
  OAI222_X1 U5523 ( .A1(n4843), .A2(n5678), .B1(n5677), .B2(n5601), .C1(n6514), 
        .C2(n4730), .ZN(U2884) );
  INV_X1 U5524 ( .A(EAX_REG_8__SCAN_IN), .ZN(n5973) );
  OAI222_X1 U5525 ( .A1(n4819), .A2(n5678), .B1(n5677), .B2(n4818), .C1(n6514), 
        .C2(n5973), .ZN(U2883) );
  OR2_X1 U5526 ( .A1(n4808), .A2(n4821), .ZN(n4822) );
  NAND2_X1 U5527 ( .A1(n4857), .A2(n4822), .ZN(n4923) );
  INV_X1 U5528 ( .A(n4860), .ZN(n4823) );
  AOI21_X1 U5529 ( .B1(n4824), .B2(n4811), .A(n4823), .ZN(n6238) );
  AOI22_X1 U5530 ( .A1(n6071), .A2(n6238), .B1(EBX_REG_9__SCAN_IN), .B2(n5445), 
        .ZN(n4825) );
  OAI21_X1 U5531 ( .B1(n4923), .B2(n6061), .A(n4825), .ZN(U2850) );
  OR2_X1 U5532 ( .A1(n4835), .A2(n5238), .ZN(n4826) );
  INV_X1 U5533 ( .A(n4827), .ZN(n4831) );
  INV_X1 U5534 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4828) );
  AOI22_X1 U5535 ( .A1(n6397), .A2(n4828), .B1(n5386), .B2(REIP_REG_1__SCAN_IN), .ZN(n4830) );
  NAND2_X1 U5536 ( .A1(n6395), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4829)
         );
  OAI211_X1 U5537 ( .C1(n4831), .C2(n6390), .A(n4830), .B(n4829), .ZN(n4832)
         );
  AOI21_X1 U5538 ( .B1(n6415), .B2(EBX_REG_1__SCAN_IN), .A(n4832), .ZN(n4838)
         );
  INV_X1 U5539 ( .A(n4833), .ZN(n4834) );
  NOR2_X1 U5540 ( .A1(n4835), .A2(n4834), .ZN(n6294) );
  INV_X1 U5541 ( .A(REIP_REG_1__SCAN_IN), .ZN(n4836) );
  AOI22_X1 U5542 ( .A1(n4800), .A2(n6294), .B1(n6296), .B2(n4836), .ZN(n4837)
         );
  OAI211_X1 U5543 ( .C1(n6318), .C2(n6082), .A(n4838), .B(n4837), .ZN(U2826)
         );
  INV_X1 U5544 ( .A(DATAI_9_), .ZN(n5460) );
  INV_X1 U5545 ( .A(EAX_REG_9__SCAN_IN), .ZN(n5975) );
  OAI222_X1 U5546 ( .A1(n4923), .A2(n5678), .B1(n5677), .B2(n5460), .C1(n6514), 
        .C2(n5975), .ZN(U2882) );
  NOR2_X1 U5547 ( .A1(n4840), .A2(n4839), .ZN(n4841) );
  OR2_X1 U5548 ( .A1(n4842), .A2(n4841), .ZN(n6335) );
  INV_X1 U5549 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4844) );
  OAI222_X1 U5550 ( .A1(n6335), .A2(n6060), .B1(n4844), .B2(n6075), .C1(n4843), 
        .C2(n6061), .ZN(U2852) );
  XOR2_X1 U5551 ( .A(n4845), .B(n4846), .Z(n4988) );
  NAND2_X1 U5552 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n4847), .ZN(n4848)
         );
  NAND2_X1 U5553 ( .A1(n6277), .A2(REIP_REG_4__SCAN_IN), .ZN(n4989) );
  OAI211_X1 U5554 ( .C1(n4849), .C2(n6227), .A(n4848), .B(n4989), .ZN(n4854)
         );
  AOI211_X1 U5555 ( .C1(n4852), .C2(n4001), .A(n4851), .B(n4850), .ZN(n4853)
         );
  AOI211_X1 U5556 ( .C1(n6281), .C2(n4988), .A(n4854), .B(n4853), .ZN(n4855)
         );
  INV_X1 U5557 ( .A(n4855), .ZN(U3014) );
  NAND2_X1 U5558 ( .A1(n4857), .A2(n4856), .ZN(n4858) );
  NAND2_X1 U5559 ( .A1(n4877), .A2(n4858), .ZN(n4945) );
  AND2_X1 U5560 ( .A1(n4860), .A2(n4859), .ZN(n4861) );
  OR2_X1 U5561 ( .A1(n4861), .A2(n4879), .ZN(n6226) );
  INV_X1 U5562 ( .A(n6226), .ZN(n4862) );
  AOI22_X1 U5563 ( .A1(n6071), .A2(n4862), .B1(EBX_REG_10__SCAN_IN), .B2(n5445), .ZN(n4863) );
  OAI21_X1 U5564 ( .B1(n4945), .B2(n6061), .A(n4863), .ZN(U2849) );
  INV_X1 U5565 ( .A(DATAI_10_), .ZN(n5567) );
  INV_X1 U5566 ( .A(EAX_REG_10__SCAN_IN), .ZN(n5977) );
  OAI222_X1 U5567 ( .A1(n4945), .A2(n5678), .B1(n5677), .B2(n5567), .C1(n6514), 
        .C2(n5977), .ZN(U2881) );
  INV_X1 U5568 ( .A(n4864), .ZN(n4871) );
  AND2_X1 U5569 ( .A1(n6295), .A2(n4868), .ZN(n4865) );
  INV_X1 U5570 ( .A(n4946), .ZN(n4884) );
  NOR2_X1 U5571 ( .A1(REIP_REG_9__SCAN_IN), .A2(n4884), .ZN(n4887) );
  AOI22_X1 U5572 ( .A1(n6415), .A2(EBX_REG_9__SCAN_IN), .B1(n6418), .B2(n6238), 
        .ZN(n4866) );
  NAND2_X1 U5573 ( .A1(n6371), .A2(n6137), .ZN(n6348) );
  OAI211_X1 U5574 ( .C1(n6412), .C2(n4867), .A(n4866), .B(n6348), .ZN(n4875)
         );
  NAND2_X1 U5575 ( .A1(n6295), .A2(n6371), .ZN(n6303) );
  INV_X1 U5576 ( .A(n6303), .ZN(n4869) );
  NAND2_X1 U5577 ( .A1(n4869), .A2(n4868), .ZN(n4870) );
  AND2_X1 U5578 ( .A1(n6304), .A2(n4870), .ZN(n6337) );
  AOI21_X1 U5579 ( .B1(n6296), .B2(n4871), .A(n6337), .ZN(n5380) );
  INV_X1 U5580 ( .A(n5380), .ZN(n4872) );
  AOI22_X1 U5581 ( .A1(n4872), .A2(REIP_REG_9__SCAN_IN), .B1(n6397), .B2(n4926), .ZN(n4873) );
  OAI21_X1 U5582 ( .B1(n6391), .B2(n4923), .A(n4873), .ZN(n4874) );
  OR3_X1 U5583 ( .A1(n4887), .A2(n4875), .A3(n4874), .ZN(U2818) );
  AND2_X1 U5584 ( .A1(n4877), .A2(n4876), .ZN(n4878) );
  OR2_X1 U5585 ( .A1(n4878), .A2(n4907), .ZN(n4911) );
  INV_X1 U5586 ( .A(n4879), .ZN(n4881) );
  INV_X1 U5587 ( .A(n4909), .ZN(n4880) );
  AOI21_X1 U5588 ( .B1(n4882), .B2(n4881), .A(n4880), .ZN(n6247) );
  AOI22_X1 U5589 ( .A1(n6071), .A2(n6247), .B1(EBX_REG_11__SCAN_IN), .B2(n5445), .ZN(n4883) );
  OAI21_X1 U5590 ( .B1(n4911), .B2(n6061), .A(n4883), .ZN(U2848) );
  NAND2_X1 U5591 ( .A1(n5380), .A2(REIP_REG_10__SCAN_IN), .ZN(n4886) );
  NOR2_X1 U5592 ( .A1(n6003), .A2(n4884), .ZN(n4885) );
  OAI22_X1 U5593 ( .A1(n4887), .A2(n4886), .B1(REIP_REG_10__SCAN_IN), .B2(
        n4885), .ZN(n4892) );
  OAI21_X1 U5594 ( .B1(n6410), .B2(n4939), .A(n6348), .ZN(n4888) );
  AOI21_X1 U5595 ( .B1(PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n6395), .A(n4888), 
        .ZN(n4889) );
  OAI21_X1 U5596 ( .B1(n6390), .B2(n6226), .A(n4889), .ZN(n4890) );
  AOI21_X1 U5597 ( .B1(n6415), .B2(EBX_REG_10__SCAN_IN), .A(n4890), .ZN(n4891)
         );
  OAI211_X1 U5598 ( .C1(n4945), .C2(n6391), .A(n4892), .B(n4891), .ZN(U2817)
         );
  INV_X1 U5599 ( .A(DATAI_11_), .ZN(n5592) );
  INV_X1 U5600 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5979) );
  OAI222_X1 U5601 ( .A1(n4911), .A2(n5678), .B1(n5677), .B2(n5592), .C1(n6514), 
        .C2(n5979), .ZN(U2880) );
  NAND2_X1 U5602 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n4894), .ZN(n6146) );
  INV_X1 U5603 ( .A(n6146), .ZN(n4895) );
  AND2_X2 U5604 ( .A1(n6659), .A2(n4895), .ZN(n5804) );
  NAND2_X1 U5605 ( .A1(n6710), .A2(n4896), .ZN(n6153) );
  NAND2_X1 U5606 ( .A1(n6153), .A2(n6482), .ZN(n4897) );
  NAND2_X1 U5607 ( .A1(n6482), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4899) );
  NAND2_X1 U5608 ( .A1(n6736), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4898) );
  AND2_X1 U5609 ( .A1(n4899), .A2(n4898), .ZN(n6076) );
  OR2_X2 U5610 ( .A1(n6123), .A2(n6076), .ZN(n6122) );
  AOI21_X1 U5611 ( .B1(n6123), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n4900), 
        .ZN(n4901) );
  OAI21_X1 U5612 ( .B1(n6122), .B2(n5387), .A(n4901), .ZN(n4902) );
  AOI21_X1 U5613 ( .B1(n5804), .B2(n5392), .A(n4902), .ZN(n4903) );
  OAI21_X1 U5614 ( .B1(n4904), .B2(n6424), .A(n4903), .ZN(U2983) );
  OAI21_X1 U5615 ( .B1(n4907), .B2(n4906), .A(n4905), .ZN(n4968) );
  NAND2_X1 U5616 ( .A1(n4909), .A2(n4908), .ZN(n4910) );
  AND2_X1 U5617 ( .A1(n4979), .A2(n4910), .ZN(n4966) );
  INV_X1 U5618 ( .A(n4966), .ZN(n4948) );
  OAI222_X1 U5619 ( .A1(n4968), .A2(n6061), .B1(n6075), .B2(n3739), .C1(n4948), 
        .C2(n6060), .ZN(U2847) );
  INV_X1 U5620 ( .A(DATAI_12_), .ZN(n5487) );
  INV_X1 U5621 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5981) );
  OAI222_X1 U5622 ( .A1(n4968), .A2(n5678), .B1(n5677), .B2(n5487), .C1(n6514), 
        .C2(n5981), .ZN(U2879) );
  INV_X1 U5623 ( .A(n4911), .ZN(n4935) );
  OAI21_X1 U5624 ( .B1(n5386), .B2(n5324), .A(n6304), .ZN(n4984) );
  AOI21_X1 U5625 ( .B1(n6395), .B2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6360), 
        .ZN(n4913) );
  AOI22_X1 U5626 ( .A1(n6415), .A2(EBX_REG_11__SCAN_IN), .B1(n6418), .B2(n6247), .ZN(n4912) );
  OAI211_X1 U5627 ( .C1(n6255), .C2(n4984), .A(n4913), .B(n4912), .ZN(n4916)
         );
  NAND4_X1 U5628 ( .A1(REIP_REG_9__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        n4946), .A4(n6255), .ZN(n4914) );
  OAI21_X1 U5629 ( .B1(n6410), .B2(n4933), .A(n4914), .ZN(n4915) );
  AOI211_X1 U5630 ( .C1(n4935), .C2(n6419), .A(n4916), .B(n4915), .ZN(n4917)
         );
  INV_X1 U5631 ( .A(n4917), .ZN(U2816) );
  NAND2_X1 U5632 ( .A1(n4999), .A2(n4919), .ZN(n4922) );
  NAND2_X1 U5633 ( .A1(n4922), .A2(n4921), .ZN(n4920) );
  OAI21_X1 U5634 ( .B1(n4922), .B2(n4921), .A(n4920), .ZN(n6239) );
  INV_X1 U5635 ( .A(n6122), .ZN(n5826) );
  NAND2_X1 U5636 ( .A1(n6277), .A2(REIP_REG_9__SCAN_IN), .ZN(n6236) );
  OAI21_X1 U5637 ( .B1(n6101), .B2(n4867), .A(n6236), .ZN(n4925) );
  INV_X2 U5638 ( .A(n5804), .ZN(n7005) );
  NOR2_X1 U5639 ( .A1(n4923), .A2(n7005), .ZN(n4924) );
  AOI211_X1 U5640 ( .C1(n5826), .C2(n4926), .A(n4925), .B(n4924), .ZN(n4927)
         );
  OAI21_X1 U5641 ( .B1(n6424), .B2(n6239), .A(n4927), .ZN(U2977) );
  XNOR2_X1 U5642 ( .A(n5692), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4937)
         );
  NAND2_X1 U5643 ( .A1(n4928), .A2(n4937), .ZN(n6229) );
  OAI21_X1 U5644 ( .B1(n4100), .B2(n5692), .A(n6229), .ZN(n4931) );
  INV_X1 U5645 ( .A(n4953), .ZN(n4929) );
  AOI21_X1 U5646 ( .B1(n5692), .B2(n6250), .A(n4929), .ZN(n4930) );
  NAND2_X1 U5647 ( .A1(n4931), .A2(n4930), .ZN(n4954) );
  OAI21_X1 U5648 ( .B1(n4931), .B2(n4930), .A(n4954), .ZN(n6246) );
  AOI22_X1 U5649 ( .A1(n6123), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .B1(n6277), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n4932) );
  OAI21_X1 U5650 ( .B1(n6122), .B2(n4933), .A(n4932), .ZN(n4934) );
  AOI21_X1 U5651 ( .B1(n4935), .B2(n5804), .A(n4934), .ZN(n4936) );
  OAI21_X1 U5652 ( .B1(n6246), .B2(n6424), .A(n4936), .ZN(U2975) );
  NOR2_X1 U5653 ( .A1(n4928), .A2(n4937), .ZN(n6224) );
  INV_X1 U5654 ( .A(n6224), .ZN(n4938) );
  INV_X1 U5655 ( .A(n6424), .ZN(n6128) );
  NAND3_X1 U5656 ( .A1(n4938), .A2(n6128), .A3(n6229), .ZN(n4944) );
  INV_X1 U5657 ( .A(n4939), .ZN(n4942) );
  INV_X1 U5658 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4940) );
  OAI22_X1 U5659 ( .A1(n6101), .A2(n4940), .B1(n6269), .B2(n6225), .ZN(n4941)
         );
  AOI21_X1 U5660 ( .B1(n4942), .B2(n5826), .A(n4941), .ZN(n4943) );
  OAI211_X1 U5661 ( .C1(n7005), .C2(n4945), .A(n4944), .B(n4943), .ZN(U2976)
         );
  OAI22_X1 U5662 ( .A1(n4968), .A2(n6391), .B1(n4971), .B2(n6410), .ZN(n4952)
         );
  NAND2_X1 U5663 ( .A1(n4947), .A2(n4946), .ZN(n6384) );
  INV_X1 U5664 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6007) );
  OAI22_X1 U5665 ( .A1(n6383), .A2(n3739), .B1(n6390), .B2(n4948), .ZN(n4949)
         );
  AOI211_X1 U5666 ( .C1(n6395), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6360), 
        .B(n4949), .ZN(n4950) );
  OAI221_X1 U5667 ( .B1(REIP_REG_12__SCAN_IN), .B2(n6384), .C1(n6007), .C2(
        n4984), .A(n4950), .ZN(n4951) );
  OR2_X1 U5668 ( .A1(n4952), .A2(n4951), .ZN(U2815) );
  NAND2_X1 U5669 ( .A1(n4954), .A2(n4953), .ZN(n4956) );
  XNOR2_X1 U5670 ( .A(n5692), .B(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4955)
         );
  XNOR2_X1 U5671 ( .A(n4956), .B(n4955), .ZN(n4975) );
  NOR2_X1 U5672 ( .A1(n6269), .A2(n6007), .ZN(n4969) );
  INV_X1 U5673 ( .A(n4957), .ZN(n4958) );
  NOR2_X1 U5674 ( .A1(n5905), .A2(n4960), .ZN(n4961) );
  NOR2_X1 U5675 ( .A1(n6249), .A2(n6250), .ZN(n4964) );
  OAI21_X1 U5676 ( .B1(n4958), .B2(n6217), .A(n6196), .ZN(n4959) );
  AOI21_X1 U5677 ( .B1(n6199), .B2(n4960), .A(n4959), .ZN(n5915) );
  INV_X1 U5678 ( .A(n5915), .ZN(n6252) );
  AOI221_X1 U5679 ( .B1(n5901), .B2(n6250), .C1(n4961), .C2(n6250), .A(n6252), 
        .ZN(n4962) );
  INV_X1 U5680 ( .A(n4962), .ZN(n4963) );
  MUX2_X1 U5681 ( .A(n4964), .B(n4963), .S(INSTADDRPOINTER_REG_12__SCAN_IN), 
        .Z(n4965) );
  AOI211_X1 U5682 ( .C1(n6280), .C2(n4966), .A(n4969), .B(n4965), .ZN(n4967)
         );
  OAI21_X1 U5683 ( .B1(n4975), .B2(n6223), .A(n4967), .ZN(U3006) );
  INV_X1 U5684 ( .A(n4968), .ZN(n4973) );
  AOI21_X1 U5685 ( .B1(n6123), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n4969), 
        .ZN(n4970) );
  OAI21_X1 U5686 ( .B1(n6122), .B2(n4971), .A(n4970), .ZN(n4972) );
  AOI21_X1 U5687 ( .B1(n4973), .B2(n5804), .A(n4972), .ZN(n4974) );
  OAI21_X1 U5688 ( .B1(n4975), .B2(n6424), .A(n4974), .ZN(U2974) );
  XNOR2_X1 U5689 ( .A(n4976), .B(n4977), .ZN(n5829) );
  INV_X1 U5690 ( .A(n5367), .ZN(n4978) );
  AOI21_X1 U5691 ( .B1(n4980), .B2(n4979), .A(n4978), .ZN(n6168) );
  AOI22_X1 U5692 ( .A1(n6071), .A2(n6168), .B1(EBX_REG_13__SCAN_IN), .B2(n5445), .ZN(n4981) );
  OAI21_X1 U5693 ( .B1(n5829), .B2(n6061), .A(n4981), .ZN(U2846) );
  INV_X1 U5694 ( .A(n6384), .ZN(n5328) );
  OAI211_X1 U5695 ( .C1(REIP_REG_12__SCAN_IN), .C2(REIP_REG_13__SCAN_IN), .A(
        n5328), .B(n5371), .ZN(n4987) );
  INV_X1 U5696 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6009) );
  AOI21_X1 U5697 ( .B1(n6395), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6360), 
        .ZN(n4983) );
  AOI22_X1 U5698 ( .A1(n6415), .A2(EBX_REG_13__SCAN_IN), .B1(n6418), .B2(n6168), .ZN(n4982) );
  OAI211_X1 U5699 ( .C1(n6009), .C2(n4984), .A(n4983), .B(n4982), .ZN(n4985)
         );
  AOI21_X1 U5700 ( .B1(n6397), .B2(n5825), .A(n4985), .ZN(n4986) );
  OAI211_X1 U5701 ( .C1(n5829), .C2(n6391), .A(n4987), .B(n4986), .ZN(U2814)
         );
  INV_X1 U5702 ( .A(n4988), .ZN(n4995) );
  INV_X1 U5703 ( .A(n6300), .ZN(n4993) );
  INV_X1 U5704 ( .A(n4989), .ZN(n4990) );
  AOI21_X1 U5705 ( .B1(n6123), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n4990), 
        .ZN(n4991) );
  OAI21_X1 U5706 ( .B1(n6122), .B2(n6299), .A(n4991), .ZN(n4992) );
  AOI21_X1 U5707 ( .B1(n4993), .B2(n5804), .A(n4992), .ZN(n4994) );
  OAI21_X1 U5708 ( .B1(n4995), .B2(n6424), .A(n4994), .ZN(U2982) );
  INV_X1 U5709 ( .A(DATAI_13_), .ZN(n5590) );
  OAI222_X1 U5710 ( .A1(n6514), .A2(n5983), .B1(n5677), .B2(n5590), .C1(n5678), 
        .C2(n5829), .ZN(U2878) );
  OR2_X1 U5711 ( .A1(n4997), .A2(n4996), .ZN(n4998) );
  NAND2_X1 U5712 ( .A1(n4999), .A2(n4998), .ZN(n6206) );
  AOI22_X1 U5713 ( .A1(n6123), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6277), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n5000) );
  OAI21_X1 U5714 ( .B1(n6122), .B2(n5376), .A(n5000), .ZN(n5001) );
  AOI21_X1 U5715 ( .B1(n5383), .B2(n5804), .A(n5001), .ZN(n5002) );
  OAI21_X1 U5716 ( .B1(n6424), .B2(n6206), .A(n5002), .ZN(U2978) );
  NAND2_X1 U5717 ( .A1(n5782), .A2(n5691), .ZN(n5004) );
  XNOR2_X1 U5718 ( .A(n5006), .B(n5005), .ZN(n5164) );
  AND2_X1 U5719 ( .A1(n6277), .A2(REIP_REG_30__SCAN_IN), .ZN(n5159) );
  NOR3_X1 U5720 ( .A1(n5843), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5007), 
        .ZN(n5008) );
  AOI211_X1 U5721 ( .C1(n5009), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5159), .B(n5008), .ZN(n5015) );
  OAI22_X1 U5722 ( .A1(n5269), .A2(n3451), .B1(n5010), .B2(n5271), .ZN(n5011)
         );
  XOR2_X1 U5723 ( .A(n5012), .B(n5011), .Z(n5265) );
  INV_X1 U5724 ( .A(n5265), .ZN(n5013) );
  NAND2_X1 U5725 ( .A1(n5013), .A2(n6280), .ZN(n5014) );
  OAI211_X1 U5726 ( .C1(n5164), .C2(n6223), .A(n5015), .B(n5014), .ZN(U2988)
         );
  AOI22_X1 U5727 ( .A1(n5068), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n5085), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5019) );
  AOI22_X1 U5728 ( .A1(n5077), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n5018) );
  AOI22_X1 U5729 ( .A1(n5078), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n5017) );
  AOI22_X1 U5730 ( .A1(n5087), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5016) );
  NAND4_X1 U5731 ( .A1(n5019), .A2(n5018), .A3(n5017), .A4(n5016), .ZN(n5025)
         );
  AOI22_X1 U5732 ( .A1(n3434), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5079), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5023) );
  AOI22_X1 U5733 ( .A1(n5076), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5022) );
  AOI22_X1 U5734 ( .A1(n5075), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5021) );
  AOI22_X1 U5735 ( .A1(n5080), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4427), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5020) );
  NAND4_X1 U5736 ( .A1(n5023), .A2(n5022), .A3(n5021), .A4(n5020), .ZN(n5024)
         );
  NOR2_X1 U5737 ( .A1(n5025), .A2(n5024), .ZN(n5107) );
  AOI22_X1 U5738 ( .A1(n5075), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5079), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5029) );
  AOI22_X1 U5739 ( .A1(n5087), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n5085), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n5028) );
  AOI22_X1 U5740 ( .A1(n5051), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5027) );
  AOI22_X1 U5741 ( .A1(n3434), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5026) );
  NAND4_X1 U5742 ( .A1(n5029), .A2(n5028), .A3(n5027), .A4(n5026), .ZN(n5035)
         );
  AOI22_X1 U5743 ( .A1(n5077), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5033) );
  AOI22_X1 U5744 ( .A1(n5037), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n5056), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5032) );
  AOI22_X1 U5745 ( .A1(n5086), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n5031) );
  AOI22_X1 U5746 ( .A1(n5068), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5030) );
  NAND4_X1 U5747 ( .A1(n5033), .A2(n5032), .A3(n5031), .A4(n5030), .ZN(n5034)
         );
  NOR2_X1 U5748 ( .A1(n5035), .A2(n5034), .ZN(n5116) );
  AOI22_X1 U5749 ( .A1(n5068), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5041) );
  AOI22_X1 U5750 ( .A1(n5079), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n5040) );
  AOI22_X1 U5751 ( .A1(n5076), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5039) );
  AOI22_X1 U5752 ( .A1(n5037), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n5038) );
  NAND4_X1 U5753 ( .A1(n5041), .A2(n5040), .A3(n5039), .A4(n5038), .ZN(n5048)
         );
  AOI22_X1 U5754 ( .A1(n5087), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n5042), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n5046) );
  AOI22_X1 U5755 ( .A1(n3434), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n5045) );
  AOI22_X1 U5756 ( .A1(n5080), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n5056), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5044) );
  AOI22_X1 U5757 ( .A1(n5077), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n5043) );
  NAND4_X1 U5758 ( .A1(n5046), .A2(n5045), .A3(n5044), .A4(n5043), .ZN(n5047)
         );
  NOR2_X1 U5759 ( .A1(n5048), .A2(n5047), .ZN(n5129) );
  OR2_X1 U5760 ( .A1(n5050), .A2(n5049), .ZN(n5130) );
  NOR2_X1 U5761 ( .A1(n5129), .A2(n5130), .ZN(n5122) );
  AOI22_X1 U5762 ( .A1(n5077), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n5079), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n5055) );
  AOI22_X1 U5763 ( .A1(n5051), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n5054) );
  AOI22_X1 U5764 ( .A1(n5076), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5053) );
  AOI22_X1 U5765 ( .A1(n5087), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5052) );
  NAND4_X1 U5766 ( .A1(n5055), .A2(n5054), .A3(n5053), .A4(n5052), .ZN(n5062)
         );
  AOI22_X1 U5767 ( .A1(n5075), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5078), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5060) );
  AOI22_X1 U5768 ( .A1(n5068), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n5059) );
  AOI22_X1 U5769 ( .A1(n5085), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5058) );
  AOI22_X1 U5770 ( .A1(n3434), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5056), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5057) );
  NAND4_X1 U5771 ( .A1(n5060), .A2(n5059), .A3(n5058), .A4(n5057), .ZN(n5061)
         );
  OR2_X1 U5772 ( .A1(n5062), .A2(n5061), .ZN(n5123) );
  NAND2_X1 U5773 ( .A1(n5122), .A2(n5123), .ZN(n5117) );
  NOR2_X1 U5774 ( .A1(n5116), .A2(n5117), .ZN(n5147) );
  AOI22_X1 U5775 ( .A1(n5077), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n5079), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5067) );
  AOI22_X1 U5776 ( .A1(n5051), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n5066) );
  AOI22_X1 U5777 ( .A1(n5076), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n5088), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5065) );
  AOI22_X1 U5778 ( .A1(n5087), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5064) );
  NAND4_X1 U5779 ( .A1(n5067), .A2(n5066), .A3(n5065), .A4(n5064), .ZN(n5074)
         );
  AOI22_X1 U5780 ( .A1(n5075), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5078), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5072) );
  AOI22_X1 U5781 ( .A1(n5068), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n5071) );
  AOI22_X1 U5782 ( .A1(n5085), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5070) );
  AOI22_X1 U5783 ( .A1(n3434), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4427), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5069) );
  NAND4_X1 U5784 ( .A1(n5072), .A2(n5071), .A3(n5070), .A4(n5069), .ZN(n5073)
         );
  OR2_X1 U5785 ( .A1(n5074), .A2(n5073), .ZN(n5148) );
  NAND2_X1 U5786 ( .A1(n5147), .A2(n5148), .ZN(n5106) );
  NOR2_X1 U5787 ( .A1(n5107), .A2(n5106), .ZN(n5096) );
  AOI22_X1 U5788 ( .A1(n5075), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5051), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5084) );
  AOI22_X1 U5789 ( .A1(n5077), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5083) );
  AOI22_X1 U5790 ( .A1(n5079), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n5078), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5082) );
  AOI22_X1 U5791 ( .A1(n5080), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n5056), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5081) );
  NAND4_X1 U5792 ( .A1(n5084), .A2(n5083), .A3(n5082), .A4(n5081), .ZN(n5094)
         );
  AOI22_X1 U5793 ( .A1(n5068), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5085), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5092) );
  AOI22_X1 U5794 ( .A1(n5087), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5086), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n5091) );
  AOI22_X1 U5795 ( .A1(n3434), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n5090) );
  AOI22_X1 U5796 ( .A1(n5088), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n5063), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5089) );
  NAND4_X1 U5797 ( .A1(n5092), .A2(n5091), .A3(n5090), .A4(n5089), .ZN(n5093)
         );
  NOR2_X1 U5798 ( .A1(n5094), .A2(n5093), .ZN(n5095) );
  XNOR2_X1 U5799 ( .A(n5096), .B(n5095), .ZN(n5097) );
  NAND2_X1 U5800 ( .A1(n5097), .A2(n5149), .ZN(n5102) );
  NAND2_X1 U5801 ( .A1(n6720), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5098)
         );
  NAND2_X1 U5802 ( .A1(n5141), .A2(n5098), .ZN(n5099) );
  AOI21_X1 U5803 ( .B1(n5221), .B2(EAX_REG_30__SCAN_IN), .A(n5099), .ZN(n5101)
         );
  XNOR2_X1 U5804 ( .A(n5105), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5257)
         );
  AOI21_X1 U5805 ( .B1(n5102), .B2(n5101), .A(n5100), .ZN(n5223) );
  NAND2_X1 U5806 ( .A1(n5103), .A2(n5272), .ZN(n5104) );
  NAND2_X1 U5807 ( .A1(n5105), .A2(n5104), .ZN(n5696) );
  XNOR2_X1 U5808 ( .A(n5107), .B(n5106), .ZN(n5110) );
  AOI21_X1 U5809 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6720), .A(n5154), 
        .ZN(n5109) );
  NAND2_X1 U5810 ( .A1(n4154), .A2(EAX_REG_29__SCAN_IN), .ZN(n5108) );
  OAI211_X1 U5811 ( .C1(n5110), .C2(n5134), .A(n5109), .B(n5108), .ZN(n5111)
         );
  OAI21_X1 U5812 ( .B1(n5141), .B2(n5696), .A(n5111), .ZN(n5268) );
  INV_X1 U5813 ( .A(n5112), .ZN(n5114) );
  INV_X1 U5814 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5113) );
  NAND2_X1 U5815 ( .A1(n5114), .A2(n5113), .ZN(n5115) );
  NAND2_X1 U5816 ( .A1(n5153), .A2(n5115), .ZN(n5713) );
  XNOR2_X1 U5817 ( .A(n5117), .B(n5116), .ZN(n5120) );
  AOI21_X1 U5818 ( .B1(PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6720), .A(n5154), 
        .ZN(n5119) );
  NAND2_X1 U5819 ( .A1(n4154), .A2(EAX_REG_27__SCAN_IN), .ZN(n5118) );
  OAI211_X1 U5820 ( .C1(n5120), .C2(n5134), .A(n5119), .B(n5118), .ZN(n5121)
         );
  OAI21_X1 U5821 ( .B1(n5141), .B2(n5713), .A(n5121), .ZN(n5291) );
  INV_X1 U5822 ( .A(n5291), .ZN(n5146) );
  XOR2_X1 U5823 ( .A(n5123), .B(n5122), .Z(n5124) );
  NAND2_X1 U5824 ( .A1(n5124), .A2(n5149), .ZN(n5128) );
  INV_X1 U5825 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5125) );
  AOI21_X1 U5826 ( .B1(n5125), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n5126) );
  AOI21_X1 U5827 ( .B1(n5221), .B2(EAX_REG_26__SCAN_IN), .A(n5126), .ZN(n5127)
         );
  XNOR2_X1 U5828 ( .A(n5140), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5722)
         );
  AOI22_X1 U5829 ( .A1(n5128), .A2(n5127), .B1(n5154), .B2(n5722), .ZN(n5305)
         );
  XNOR2_X1 U5830 ( .A(n5130), .B(n5129), .ZN(n5135) );
  NAND2_X1 U5831 ( .A1(n6720), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5131)
         );
  NAND2_X1 U5832 ( .A1(n5141), .A2(n5131), .ZN(n5132) );
  AOI21_X1 U5833 ( .B1(n4154), .B2(EAX_REG_25__SCAN_IN), .A(n5132), .ZN(n5133)
         );
  OAI21_X1 U5834 ( .B1(n5135), .B2(n5134), .A(n5133), .ZN(n5143) );
  INV_X1 U5835 ( .A(n5136), .ZN(n5138) );
  INV_X1 U5836 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5137) );
  NAND2_X1 U5837 ( .A1(n5138), .A2(n5137), .ZN(n5139) );
  NAND2_X1 U5838 ( .A1(n5140), .A2(n5139), .ZN(n5732) );
  OR2_X1 U5839 ( .A1(n5732), .A2(n5141), .ZN(n5142) );
  NAND2_X1 U5840 ( .A1(n5143), .A2(n5142), .ZN(n5165) );
  NOR2_X1 U5841 ( .A1(n5165), .A2(n5144), .ZN(n5167) );
  AND2_X1 U5842 ( .A1(n5305), .A2(n5167), .ZN(n5145) );
  XOR2_X1 U5843 ( .A(n5148), .B(n5147), .Z(n5150) );
  NAND2_X1 U5844 ( .A1(n5150), .A2(n5149), .ZN(n5156) );
  NOR2_X1 U5845 ( .A1(n5151), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5152) );
  AOI211_X1 U5846 ( .C1(n5221), .C2(EAX_REG_28__SCAN_IN), .A(n5154), .B(n5152), 
        .ZN(n5155) );
  XNOR2_X1 U5847 ( .A(n5153), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5700)
         );
  AOI22_X1 U5848 ( .A1(n5156), .A2(n5155), .B1(n5154), .B2(n5700), .ZN(n5281)
         );
  INV_X1 U5849 ( .A(n5266), .ZN(n5157) );
  NOR2_X1 U5850 ( .A1(n5268), .A2(n5157), .ZN(n5158) );
  AND2_X2 U5851 ( .A1(n5158), .A2(n3439), .ZN(n5267) );
  XOR2_X2 U5852 ( .A(n5223), .B(n5267), .Z(n5447) );
  INV_X1 U5853 ( .A(n5257), .ZN(n5161) );
  AOI21_X1 U5854 ( .B1(n6123), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5159), 
        .ZN(n5160) );
  OAI21_X1 U5855 ( .B1(n6122), .B2(n5161), .A(n5160), .ZN(n5162) );
  AOI21_X1 U5856 ( .B1(n5447), .B2(n5804), .A(n5162), .ZN(n5163) );
  OAI21_X1 U5857 ( .B1(n5164), .B2(n6424), .A(n5163), .ZN(U2956) );
  INV_X1 U5858 ( .A(n5165), .ZN(n5169) );
  AOI22_X1 U5859 ( .A1(n6533), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6536), .ZN(n5173) );
  AND2_X1 U5860 ( .A1(n6914), .A2(n5170), .ZN(n5171) );
  NAND2_X1 U5861 ( .A1(n6537), .A2(DATAI_9_), .ZN(n5172) );
  OAI211_X1 U5862 ( .C1(n5735), .C2(n5678), .A(n5173), .B(n5172), .ZN(U2866)
         );
  INV_X1 U5863 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5184) );
  NOR2_X1 U5864 ( .A1(n5176), .A2(n5175), .ZN(n5177) );
  OR2_X1 U5865 ( .A1(n5174), .A2(n5177), .ZN(n5178) );
  OAI222_X1 U5866 ( .A1(n5735), .A2(n6061), .B1(n5184), .B2(n6075), .C1(n5178), 
        .C2(n6060), .ZN(U2834) );
  INV_X1 U5867 ( .A(n5178), .ZN(n6279) );
  INV_X1 U5868 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6025) );
  AOI21_X1 U5869 ( .B1(n6423), .B2(n5179), .A(n6025), .ZN(n5186) );
  INV_X1 U5870 ( .A(n5732), .ZN(n5180) );
  AOI22_X1 U5871 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n6395), .B1(n6397), 
        .B2(n5180), .ZN(n5183) );
  NOR2_X1 U5872 ( .A1(n6023), .A2(n5181), .ZN(n5244) );
  NAND3_X1 U5873 ( .A1(n6296), .A2(n5244), .A3(n6025), .ZN(n5182) );
  OAI211_X1 U5874 ( .C1(n6383), .C2(n5184), .A(n5183), .B(n5182), .ZN(n5185)
         );
  AOI211_X1 U5875 ( .C1(n6279), .C2(n6418), .A(n5186), .B(n5185), .ZN(n5187)
         );
  OAI21_X1 U5876 ( .B1(n5735), .B2(n6391), .A(n5187), .ZN(U2802) );
  INV_X1 U5877 ( .A(n5188), .ZN(n5748) );
  NOR2_X1 U5878 ( .A1(n6075), .A2(n5189), .ZN(n5190) );
  AOI21_X1 U5879 ( .B1(n5862), .B2(n6071), .A(n5190), .ZN(n5191) );
  OAI21_X1 U5880 ( .B1(n5188), .B2(n6061), .A(n5191), .ZN(U2835) );
  NOR2_X1 U5881 ( .A1(n5193), .A2(n5192), .ZN(n5194) );
  OR2_X1 U5882 ( .A1(n5195), .A2(n5194), .ZN(n5199) );
  INV_X1 U5883 ( .A(n5199), .ZN(n6182) );
  AOI22_X1 U5884 ( .A1(n6071), .A2(n6182), .B1(EBX_REG_2__SCAN_IN), .B2(n5445), 
        .ZN(n5196) );
  OAI21_X1 U5885 ( .B1(n6061), .B2(n6091), .A(n5196), .ZN(U2857) );
  INV_X1 U5886 ( .A(n4677), .ZN(n6569) );
  AOI22_X1 U5887 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6395), .B1(n5386), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n5197) );
  OAI21_X1 U5888 ( .B1(n6410), .B2(n6095), .A(n5197), .ZN(n5201) );
  OAI211_X1 U5889 ( .C1(REIP_REG_1__SCAN_IN), .C2(REIP_REG_2__SCAN_IN), .A(
        n6296), .B(n5385), .ZN(n5198) );
  OAI21_X1 U5890 ( .B1(n5199), .B2(n6390), .A(n5198), .ZN(n5200) );
  AOI211_X1 U5891 ( .C1(n6569), .C2(n6294), .A(n5201), .B(n5200), .ZN(n5203)
         );
  NAND2_X1 U5892 ( .A1(n6415), .A2(EBX_REG_2__SCAN_IN), .ZN(n5202) );
  OAI211_X1 U5893 ( .C1(n6318), .C2(n6091), .A(n5203), .B(n5202), .ZN(U2825)
         );
  INV_X1 U5894 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5210) );
  INV_X1 U5895 ( .A(n5204), .ZN(n5935) );
  AOI22_X1 U5896 ( .A1(n4153), .A2(n5939), .B1(n5935), .B2(n5210), .ZN(n6431)
         );
  INV_X1 U5897 ( .A(n6469), .ZN(n5947) );
  AOI22_X1 U5898 ( .A1(n5210), .A2(n5205), .B1(n5940), .B2(
        STATE2_REG_1__SCAN_IN), .ZN(n5206) );
  OAI21_X1 U5899 ( .B1(n6431), .B2(n5947), .A(n5206), .ZN(n5208) );
  INV_X1 U5900 ( .A(n5207), .ZN(n5937) );
  NOR2_X1 U5901 ( .A1(n5937), .A2(n5210), .ZN(n6432) );
  AOI22_X1 U5902 ( .A1(n6430), .A2(n5208), .B1(n6469), .B2(n6432), .ZN(n5209)
         );
  OAI21_X1 U5903 ( .B1(n5210), .B2(n6430), .A(n5209), .ZN(U3461) );
  INV_X1 U5904 ( .A(n5447), .ZN(n5211) );
  INV_X1 U5905 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5259) );
  OAI222_X1 U5906 ( .A1(n6061), .A2(n5211), .B1(n5259), .B2(n6075), .C1(n5265), 
        .C2(n6060), .ZN(U2829) );
  INV_X1 U5907 ( .A(n5212), .ZN(n5219) );
  INV_X1 U5908 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5213) );
  AOI22_X1 U5909 ( .A1(INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n5929), .B1(
        INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n5213), .ZN(n5945) );
  NOR3_X1 U5910 ( .A1(n6475), .A2(n5940), .A3(n5945), .ZN(n5215) );
  NOR3_X1 U5911 ( .A1(n5934), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n6478), 
        .ZN(n5214) );
  AOI211_X1 U5912 ( .C1(n5216), .C2(n6469), .A(n5215), .B(n5214), .ZN(n5217)
         );
  OAI22_X1 U5913 ( .A1(n5219), .A2(n5218), .B1(n5948), .B2(n5217), .ZN(U3459)
         );
  AOI22_X1 U5914 ( .A1(n5221), .A2(EAX_REG_31__SCAN_IN), .B1(n5220), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5222) );
  INV_X1 U5915 ( .A(n5222), .ZN(n5225) );
  NAND2_X1 U5916 ( .A1(n5267), .A2(n5223), .ZN(n5224) );
  NAND3_X1 U5917 ( .A1(n5683), .A2(n7000), .A3(n6514), .ZN(n5227) );
  AOI22_X1 U5918 ( .A1(n6533), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6536), .ZN(n5226) );
  NAND2_X1 U5919 ( .A1(n5227), .A2(n5226), .ZN(U2860) );
  INV_X1 U5920 ( .A(n5236), .ZN(n5234) );
  OR2_X1 U5921 ( .A1(n5239), .A2(n5228), .ZN(n5233) );
  NAND2_X1 U5922 ( .A1(n5230), .A2(n5229), .ZN(n5231) );
  NAND2_X1 U5923 ( .A1(n5239), .A2(n5231), .ZN(n5232) );
  OAI211_X1 U5924 ( .C1(n5235), .C2(n5234), .A(n5233), .B(n5232), .ZN(n6449)
         );
  AOI21_X1 U5925 ( .B1(n5236), .B2(n5235), .A(n4495), .ZN(n5237) );
  AOI21_X1 U5926 ( .B1(n5239), .B2(n5238), .A(n5237), .ZN(n6131) );
  OR2_X1 U5927 ( .A1(n5241), .A2(n5240), .ZN(n6139) );
  OAI21_X1 U5928 ( .B1(n6139), .B2(n5242), .A(n6500), .ZN(n6149) );
  AND2_X1 U5929 ( .A1(n6131), .A2(n6149), .ZN(n6453) );
  NOR2_X1 U5930 ( .A1(n6453), .A2(n6487), .ZN(n6425) );
  MUX2_X1 U5931 ( .A(MORE_REG_SCAN_IN), .B(n6449), .S(n6425), .Z(U3471) );
  NAND2_X1 U5932 ( .A1(n5683), .A2(n6419), .ZN(n5256) );
  AND2_X1 U5933 ( .A1(REIP_REG_25__SCAN_IN), .A2(n5244), .ZN(n5310) );
  NAND2_X1 U5934 ( .A1(REIP_REG_26__SCAN_IN), .A2(n5310), .ZN(n5248) );
  AOI21_X1 U5935 ( .B1(n6296), .B2(n5248), .A(n5386), .ZN(n5314) );
  INV_X1 U5936 ( .A(REIP_REG_28__SCAN_IN), .ZN(n5561) );
  INV_X1 U5937 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6031) );
  OR2_X1 U5938 ( .A1(n5561), .A2(n6031), .ZN(n5245) );
  NAND2_X1 U5939 ( .A1(n6304), .A2(n5245), .ZN(n5246) );
  NAND2_X1 U5940 ( .A1(n5314), .A2(n5246), .ZN(n5286) );
  AOI21_X1 U5941 ( .B1(REIP_REG_30__SCAN_IN), .B2(REIP_REG_29__SCAN_IN), .A(
        n5249), .ZN(n5247) );
  OR2_X1 U5942 ( .A1(n5286), .A2(n5247), .ZN(n5262) );
  NOR2_X1 U5943 ( .A1(n5249), .A2(n5248), .ZN(n5296) );
  NAND3_X1 U5944 ( .A1(n5296), .A2(REIP_REG_28__SCAN_IN), .A3(
        REIP_REG_27__SCAN_IN), .ZN(n5276) );
  INV_X1 U5945 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6039) );
  NAND3_X1 U5946 ( .A1(REIP_REG_30__SCAN_IN), .A2(REIP_REG_29__SCAN_IN), .A3(
        n6039), .ZN(n5253) );
  NAND2_X1 U5947 ( .A1(n6395), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5252)
         );
  NAND3_X1 U5948 ( .A1(n5250), .A2(n3818), .A3(EBX_REG_31__SCAN_IN), .ZN(n5251) );
  OAI211_X1 U5949 ( .C1(n5276), .C2(n5253), .A(n5252), .B(n5251), .ZN(n5254)
         );
  AOI21_X1 U5950 ( .B1(REIP_REG_31__SCAN_IN), .B2(n5262), .A(n5254), .ZN(n5255) );
  OAI211_X1 U5951 ( .C1(n5243), .C2(n6390), .A(n5256), .B(n5255), .ZN(U2796)
         );
  NAND2_X1 U5952 ( .A1(n5447), .A2(n6419), .ZN(n5264) );
  INV_X1 U5953 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6033) );
  OAI21_X1 U5954 ( .B1(n5276), .B2(n6033), .A(n6035), .ZN(n5261) );
  AOI22_X1 U5955 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n6395), .B1(n6397), 
        .B2(n5257), .ZN(n5258) );
  OAI21_X1 U5956 ( .B1(n6383), .B2(n5259), .A(n5258), .ZN(n5260) );
  AOI21_X1 U5957 ( .B1(n5262), .B2(n5261), .A(n5260), .ZN(n5263) );
  OAI211_X1 U5958 ( .C1(n6390), .C2(n5265), .A(n5264), .B(n5263), .ZN(U2797)
         );
  NAND2_X1 U5959 ( .A1(n3438), .A2(n5266), .ZN(n5280) );
  INV_X1 U5960 ( .A(n5698), .ZN(n5400) );
  AOI21_X1 U5961 ( .B1(n5271), .B2(n5270), .A(n5269), .ZN(n5833) );
  OAI22_X1 U5962 ( .A1(n5272), .A2(n6412), .B1(n6410), .B2(n5696), .ZN(n5273)
         );
  AOI21_X1 U5963 ( .B1(n6415), .B2(EBX_REG_29__SCAN_IN), .A(n5273), .ZN(n5275)
         );
  NAND2_X1 U5964 ( .A1(n5286), .A2(REIP_REG_29__SCAN_IN), .ZN(n5274) );
  OAI211_X1 U5965 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5276), .A(n5275), .B(n5274), .ZN(n5277) );
  AOI21_X1 U5966 ( .B1(n5833), .B2(n6418), .A(n5277), .ZN(n5278) );
  OAI21_X1 U5967 ( .B1(n5400), .B2(n6391), .A(n5278), .ZN(U2798) );
  AND2_X2 U5968 ( .A1(n5407), .A2(n5279), .ZN(n5290) );
  INV_X1 U5969 ( .A(n5454), .ZN(n5705) );
  NAND2_X1 U5970 ( .A1(n5705), .A2(n6419), .ZN(n5288) );
  NAND2_X1 U5971 ( .A1(n6415), .A2(EBX_REG_28__SCAN_IN), .ZN(n5284) );
  AOI22_X1 U5972 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n6395), .B1(n6397), 
        .B2(n5700), .ZN(n5283) );
  NAND3_X1 U5973 ( .A1(n5296), .A2(REIP_REG_27__SCAN_IN), .A3(n5561), .ZN(
        n5282) );
  NAND3_X1 U5974 ( .A1(n5284), .A2(n5283), .A3(n5282), .ZN(n5285) );
  AOI21_X1 U5975 ( .B1(REIP_REG_28__SCAN_IN), .B2(n5286), .A(n5285), .ZN(n5287) );
  OAI211_X1 U5976 ( .C1(n6390), .C2(n5401), .A(n5288), .B(n5287), .ZN(U2799)
         );
  NAND2_X1 U5977 ( .A1(n3438), .A2(n5289), .ZN(n5304) );
  AOI21_X2 U5978 ( .B1(n5291), .B2(n5304), .A(n5290), .ZN(n5715) );
  INV_X1 U5979 ( .A(n5715), .ZN(n5663) );
  OR2_X1 U5980 ( .A1(n5309), .A2(n5292), .ZN(n5294) );
  NAND2_X1 U5981 ( .A1(n5294), .A2(n5293), .ZN(n5403) );
  INV_X1 U5982 ( .A(n5403), .ZN(n5841) );
  OR2_X1 U5983 ( .A1(n5314), .A2(n6031), .ZN(n5300) );
  INV_X1 U5984 ( .A(n5713), .ZN(n5295) );
  AOI22_X1 U5985 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n6395), .B1(n6397), 
        .B2(n5295), .ZN(n5299) );
  NAND2_X1 U5986 ( .A1(n5296), .A2(n6031), .ZN(n5298) );
  NAND2_X1 U5987 ( .A1(n6415), .A2(EBX_REG_27__SCAN_IN), .ZN(n5297) );
  NAND4_X1 U5988 ( .A1(n5300), .A2(n5299), .A3(n5298), .A4(n5297), .ZN(n5301)
         );
  AOI21_X1 U5989 ( .B1(n5841), .B2(n6418), .A(n5301), .ZN(n5302) );
  OAI21_X1 U5990 ( .B1(n5663), .B2(n6391), .A(n5302), .ZN(U2800) );
  NOR2_X1 U5991 ( .A1(n5174), .A2(n5307), .ZN(n5308) );
  OR2_X1 U5992 ( .A1(n5309), .A2(n5308), .ZN(n5849) );
  INV_X1 U5993 ( .A(n5849), .ZN(n5316) );
  AOI21_X1 U5994 ( .B1(n6296), .B2(n5310), .A(REIP_REG_26__SCAN_IN), .ZN(n5313) );
  AOI22_X1 U5995 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n6395), .B1(n6397), 
        .B2(n5722), .ZN(n5312) );
  NAND2_X1 U5996 ( .A1(n6415), .A2(EBX_REG_26__SCAN_IN), .ZN(n5311) );
  OAI211_X1 U5997 ( .C1(n5314), .C2(n5313), .A(n5312), .B(n5311), .ZN(n5315)
         );
  AOI21_X1 U5998 ( .B1(n5316), .B2(n6418), .A(n5315), .ZN(n5317) );
  OAI21_X1 U5999 ( .B1(n5721), .B2(n6391), .A(n5317), .ZN(U2801) );
  AOI21_X1 U6000 ( .B1(n5335), .B2(n5321), .A(n5320), .ZN(n6520) );
  INV_X1 U6001 ( .A(n6520), .ZN(n5432) );
  NAND2_X1 U6002 ( .A1(n5342), .A2(n5322), .ZN(n5323) );
  NAND2_X1 U6003 ( .A1(n6069), .A2(n5323), .ZN(n5909) );
  INV_X1 U6004 ( .A(n5329), .ZN(n5325) );
  NOR3_X1 U6005 ( .A1(n5386), .A2(n5325), .A3(n5324), .ZN(n5355) );
  INV_X1 U6006 ( .A(n6304), .ZN(n6370) );
  AOI21_X1 U6007 ( .B1(n5355), .B2(n5330), .A(n6370), .ZN(n6363) );
  AOI22_X1 U6008 ( .A1(n5786), .A2(n6397), .B1(REIP_REG_18__SCAN_IN), .B2(
        n6363), .ZN(n5327) );
  AOI21_X1 U6009 ( .B1(n6395), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6360), 
        .ZN(n5326) );
  OAI211_X1 U6010 ( .C1(n6390), .C2(n5909), .A(n5327), .B(n5326), .ZN(n5331)
         );
  INV_X1 U6011 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U6012 ( .A1(n5329), .A2(n5328), .ZN(n6375) );
  INV_X1 U6013 ( .A(n6375), .ZN(n5353) );
  AND3_X1 U6014 ( .A1(n6016), .A2(n5330), .A3(n5353), .ZN(n6364) );
  AOI211_X1 U6015 ( .C1(n6415), .C2(EBX_REG_18__SCAN_IN), .A(n5331), .B(n6364), 
        .ZN(n5332) );
  OAI21_X1 U6016 ( .B1(n5432), .B2(n6391), .A(n5332), .ZN(U2809) );
  INV_X1 U6017 ( .A(n5335), .ZN(n5336) );
  AOI21_X1 U6018 ( .B1(n5337), .B2(n5334), .A(n5336), .ZN(n6513) );
  INV_X1 U6019 ( .A(n6513), .ZN(n5435) );
  OAI21_X1 U6020 ( .B1(n5352), .B2(n6375), .A(n6268), .ZN(n5347) );
  INV_X1 U6021 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5338) );
  OAI22_X1 U6022 ( .A1(n5338), .A2(n6412), .B1(n6121), .B2(n6410), .ZN(n5346)
         );
  INV_X1 U6023 ( .A(n5339), .ZN(n5354) );
  NAND2_X1 U6024 ( .A1(n5443), .A2(n5354), .ZN(n5341) );
  NAND2_X1 U6025 ( .A1(n5341), .A2(n5340), .ZN(n5343) );
  AND2_X1 U6026 ( .A1(n5343), .A2(n5342), .ZN(n6266) );
  INV_X1 U6027 ( .A(n6266), .ZN(n5433) );
  NAND2_X1 U6028 ( .A1(n6415), .A2(EBX_REG_17__SCAN_IN), .ZN(n5344) );
  OAI211_X1 U6029 ( .C1(n5433), .C2(n6390), .A(n5344), .B(n6348), .ZN(n5345)
         );
  AOI211_X1 U6030 ( .C1(n5347), .C2(n6363), .A(n5346), .B(n5345), .ZN(n5348)
         );
  OAI21_X1 U6031 ( .B1(n5435), .B2(n6391), .A(n5348), .ZN(U2810) );
  OAI21_X1 U6032 ( .B1(n5350), .B2(n5351), .A(n5334), .ZN(n5799) );
  OAI211_X1 U6033 ( .C1(REIP_REG_15__SCAN_IN), .C2(REIP_REG_16__SCAN_IN), .A(
        n5353), .B(n5352), .ZN(n5360) );
  XNOR2_X1 U6034 ( .A(n5443), .B(n5354), .ZN(n5436) );
  NOR2_X1 U6035 ( .A1(n6370), .A2(n5355), .ZN(n6352) );
  AOI22_X1 U6036 ( .A1(n5794), .A2(n6397), .B1(REIP_REG_16__SCAN_IN), .B2(
        n6352), .ZN(n5357) );
  AOI21_X1 U6037 ( .B1(n6395), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6360), 
        .ZN(n5356) );
  OAI211_X1 U6038 ( .C1(n6390), .C2(n5436), .A(n5357), .B(n5356), .ZN(n5358)
         );
  AOI21_X1 U6039 ( .B1(n6415), .B2(EBX_REG_16__SCAN_IN), .A(n5358), .ZN(n5359)
         );
  OAI211_X1 U6040 ( .C1(n5799), .C2(n6391), .A(n5360), .B(n5359), .ZN(U2811)
         );
  OAI21_X1 U6041 ( .B1(n5363), .B2(n5362), .A(n5438), .ZN(n5814) );
  INV_X1 U6042 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5364) );
  NOR2_X1 U6043 ( .A1(n6412), .A2(n5364), .ZN(n5365) );
  AOI211_X1 U6044 ( .C1(REIP_REG_14__SCAN_IN), .C2(n6352), .A(n6360), .B(n5365), .ZN(n5370) );
  AND2_X1 U6045 ( .A1(n5367), .A2(n5366), .ZN(n5368) );
  NOR2_X1 U6046 ( .A1(n5441), .A2(n5368), .ZN(n6176) );
  NAND2_X1 U6047 ( .A1(n6418), .A2(n6176), .ZN(n5369) );
  OAI211_X1 U6048 ( .C1(n6410), .C2(n5816), .A(n5370), .B(n5369), .ZN(n5373)
         );
  NOR3_X1 U6049 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5371), .A3(n6384), .ZN(n5372) );
  AOI211_X1 U6050 ( .C1(n6415), .C2(EBX_REG_14__SCAN_IN), .A(n5373), .B(n5372), 
        .ZN(n5374) );
  OAI21_X1 U6051 ( .B1(n5814), .B2(n6391), .A(n5374), .ZN(U2813) );
  NOR3_X1 U6052 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6338), .A3(n6340), .ZN(n5382)
         );
  NAND2_X1 U6053 ( .A1(n6395), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5375)
         );
  OAI211_X1 U6054 ( .C1(n6410), .C2(n5376), .A(n6348), .B(n5375), .ZN(n5377)
         );
  AOI21_X1 U6055 ( .B1(n6418), .B2(n6203), .A(n5377), .ZN(n5379) );
  NAND2_X1 U6056 ( .A1(n6415), .A2(EBX_REG_8__SCAN_IN), .ZN(n5378) );
  OAI211_X1 U6057 ( .C1(n5380), .C2(n6001), .A(n5379), .B(n5378), .ZN(n5381)
         );
  AOI211_X1 U6058 ( .C1(n5383), .C2(n6419), .A(n5382), .B(n5381), .ZN(n5384)
         );
  INV_X1 U6059 ( .A(n5384), .ZN(U2819) );
  AND2_X1 U6060 ( .A1(n6304), .A2(n6303), .ZN(n5391) );
  OAI21_X1 U6061 ( .B1(n5386), .B2(n5385), .A(n5993), .ZN(n5390) );
  OAI22_X1 U6062 ( .A1(n5388), .A2(n6412), .B1(n6410), .B2(n5387), .ZN(n5389)
         );
  AOI21_X1 U6063 ( .B1(n5391), .B2(n5390), .A(n5389), .ZN(n5397) );
  INV_X1 U6064 ( .A(n6318), .ZN(n5393) );
  AOI22_X1 U6065 ( .A1(n5393), .A2(n5392), .B1(n6415), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n5396) );
  AOI22_X1 U6066 ( .A1(n6294), .A2(n6630), .B1(n6418), .B2(n5394), .ZN(n5395)
         );
  NAND3_X1 U6067 ( .A1(n5397), .A2(n5396), .A3(n5395), .ZN(U2824) );
  OAI22_X1 U6068 ( .A1(n5243), .A2(n6060), .B1(n6075), .B2(n5398), .ZN(U2828)
         );
  AOI22_X1 U6069 ( .A1(n5833), .A2(n6071), .B1(EBX_REG_29__SCAN_IN), .B2(n5445), .ZN(n5399) );
  OAI21_X1 U6070 ( .B1(n5400), .B2(n6061), .A(n5399), .ZN(U2830) );
  OAI222_X1 U6071 ( .A1(n6061), .A2(n5454), .B1(n5402), .B2(n6075), .C1(n5401), 
        .C2(n6060), .ZN(U2831) );
  INV_X1 U6072 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5404) );
  OAI222_X1 U6073 ( .A1(n6061), .A2(n5663), .B1(n5404), .B2(n6075), .C1(n5403), 
        .C2(n6060), .ZN(U2832) );
  OAI222_X1 U6074 ( .A1(n5721), .A2(n6061), .B1(n5405), .B2(n6075), .C1(n5849), 
        .C2(n6060), .ZN(U2833) );
  INV_X1 U6075 ( .A(n5406), .ZN(n5408) );
  INV_X1 U6076 ( .A(n3439), .ZN(n5415) );
  INV_X1 U6077 ( .A(n6535), .ZN(n5413) );
  INV_X1 U6078 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U6079 ( .A1(n5420), .A2(n5409), .ZN(n5410) );
  NAND2_X1 U6080 ( .A1(n5411), .A2(n5410), .ZN(n6416) );
  OAI222_X1 U6081 ( .A1(n5413), .A2(n6061), .B1(n5412), .B2(n6075), .C1(n6060), 
        .C2(n6416), .ZN(U2836) );
  NAND2_X1 U6082 ( .A1(n5884), .A2(n5418), .ZN(n5419) );
  NAND2_X1 U6083 ( .A1(n5420), .A2(n5419), .ZN(n5874) );
  INV_X1 U6084 ( .A(n5874), .ZN(n6400) );
  AOI22_X1 U6085 ( .A1(n6400), .A2(n6071), .B1(EBX_REG_22__SCAN_IN), .B2(n5445), .ZN(n5421) );
  OAI21_X1 U6086 ( .B1(n6399), .B2(n6061), .A(n5421), .ZN(U2837) );
  NOR2_X1 U6087 ( .A1(n6068), .A2(n5423), .ZN(n5424) );
  OR2_X1 U6088 ( .A1(n5422), .A2(n5424), .ZN(n6377) );
  AND2_X1 U6089 ( .A1(n5427), .A2(n5428), .ZN(n5429) );
  NOR2_X1 U6090 ( .A1(n5426), .A2(n5429), .ZN(n5779) );
  INV_X1 U6091 ( .A(n5779), .ZN(n6378) );
  OAI222_X1 U6092 ( .A1(n6060), .A2(n6377), .B1(n6075), .B2(n3771), .C1(n6378), 
        .C2(n6061), .ZN(U2839) );
  INV_X1 U6093 ( .A(n5909), .ZN(n5430) );
  AOI22_X1 U6094 ( .A1(n5430), .A2(n6071), .B1(EBX_REG_18__SCAN_IN), .B2(n5445), .ZN(n5431) );
  OAI21_X1 U6095 ( .B1(n5432), .B2(n6061), .A(n5431), .ZN(U2841) );
  INV_X1 U6096 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5434) );
  OAI222_X1 U6097 ( .A1(n5435), .A2(n6061), .B1(n5434), .B2(n6075), .C1(n5433), 
        .C2(n6060), .ZN(U2842) );
  INV_X1 U6098 ( .A(n5436), .ZN(n6257) );
  AOI22_X1 U6099 ( .A1(n6257), .A2(n6071), .B1(EBX_REG_16__SCAN_IN), .B2(n5445), .ZN(n5437) );
  OAI21_X1 U6100 ( .B1(n5799), .B2(n6061), .A(n5437), .ZN(U2843) );
  AOI21_X1 U6101 ( .B1(n5439), .B2(n5438), .A(n5350), .ZN(n6354) );
  INV_X1 U6102 ( .A(n6354), .ZN(n5675) );
  INV_X1 U6103 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5444) );
  NOR2_X1 U6104 ( .A1(n5441), .A2(n5440), .ZN(n5442) );
  OR2_X1 U6105 ( .A1(n5443), .A2(n5442), .ZN(n5918) );
  OAI222_X1 U6106 ( .A1(n5675), .A2(n6061), .B1(n5444), .B2(n6075), .C1(n5918), 
        .C2(n6060), .ZN(U2844) );
  AOI22_X1 U6107 ( .A1(n6071), .A2(n6176), .B1(EBX_REG_14__SCAN_IN), .B2(n5445), .ZN(n5446) );
  OAI21_X1 U6108 ( .B1(n5814), .B2(n6061), .A(n5446), .ZN(U2845) );
  NAND2_X1 U6109 ( .A1(n5447), .A2(n6534), .ZN(n5449) );
  AOI22_X1 U6110 ( .A1(n6533), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6536), .ZN(n5448) );
  OAI211_X1 U6111 ( .C1(n6516), .C2(n5676), .A(n5449), .B(n5448), .ZN(U2861)
         );
  NAND2_X1 U6112 ( .A1(n5698), .A2(n6534), .ZN(n5451) );
  AOI22_X1 U6113 ( .A1(n6533), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6536), .ZN(n5450) );
  OAI211_X1 U6114 ( .C1(n6516), .C2(n5590), .A(n5451), .B(n5450), .ZN(U2862)
         );
  AOI22_X1 U6115 ( .A1(n6533), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6536), .ZN(n5453) );
  NAND2_X1 U6116 ( .A1(n6537), .A2(DATAI_12_), .ZN(n5452) );
  OAI211_X1 U6117 ( .C1(n5454), .C2(n5678), .A(n5453), .B(n5452), .ZN(U2863)
         );
  INV_X1 U6118 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6374) );
  INV_X1 U6119 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6402) );
  AOI22_X1 U6120 ( .A1(REIP_REG_23__SCAN_IN), .A2(keyinput_59), .B1(n6023), 
        .B2(keyinput_58), .ZN(n5455) );
  OAI221_X1 U6121 ( .B1(REIP_REG_23__SCAN_IN), .B2(keyinput_59), .C1(n6023), 
        .C2(keyinput_58), .A(n5455), .ZN(n5550) );
  INV_X1 U6122 ( .A(keyinput_57), .ZN(n5548) );
  INV_X1 U6123 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6027) );
  AOI22_X1 U6124 ( .A1(REIP_REG_28__SCAN_IN), .A2(keyinput_54), .B1(n6031), 
        .B2(keyinput_55), .ZN(n5456) );
  OAI221_X1 U6125 ( .B1(REIP_REG_28__SCAN_IN), .B2(keyinput_54), .C1(n6031), 
        .C2(keyinput_55), .A(n5456), .ZN(n5545) );
  INV_X1 U6126 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6035) );
  AOI22_X1 U6127 ( .A1(REIP_REG_31__SCAN_IN), .A2(keyinput_51), .B1(n6035), 
        .B2(keyinput_52), .ZN(n5457) );
  OAI221_X1 U6128 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_51), .C1(n6035), 
        .C2(keyinput_52), .A(n5457), .ZN(n5542) );
  INV_X1 U6129 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5645) );
  INV_X1 U6130 ( .A(keyinput_50), .ZN(n5540) );
  INV_X1 U6131 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6053) );
  INV_X1 U6132 ( .A(keyinput_49), .ZN(n5538) );
  INV_X1 U6133 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6056) );
  INV_X1 U6134 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6058) );
  INV_X1 U6135 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6141) );
  AOI22_X1 U6136 ( .A1(n6058), .A2(keyinput_47), .B1(keyinput_46), .B2(n6141), 
        .ZN(n5458) );
  OAI221_X1 U6137 ( .B1(n6058), .B2(keyinput_47), .C1(n6141), .C2(keyinput_46), 
        .A(n5458), .ZN(n5535) );
  INV_X1 U6138 ( .A(keyinput_45), .ZN(n5533) );
  INV_X1 U6139 ( .A(keyinput_44), .ZN(n5531) );
  INV_X1 U6140 ( .A(MORE_REG_SCAN_IN), .ZN(n6450) );
  XOR2_X1 U6141 ( .A(M_IO_N_REG_SCAN_IN), .B(keyinput_40), .Z(n5529) );
  INV_X1 U6142 ( .A(keyinput_39), .ZN(n5524) );
  INV_X1 U6143 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6132) );
  INV_X1 U6144 ( .A(keyinput_38), .ZN(n5522) );
  INV_X1 U6145 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5954) );
  INV_X1 U6146 ( .A(BS16_N), .ZN(n5950) );
  INV_X1 U6147 ( .A(keyinput_34), .ZN(n5516) );
  INV_X1 U6148 ( .A(keyinput_32), .ZN(n5510) );
  INV_X1 U6149 ( .A(keyinput_30), .ZN(n5504) );
  INV_X1 U6150 ( .A(keyinput_24), .ZN(n5495) );
  AOI22_X1 U6151 ( .A1(n5567), .A2(keyinput_21), .B1(keyinput_22), .B2(n5460), 
        .ZN(n5459) );
  OAI221_X1 U6152 ( .B1(n5567), .B2(keyinput_21), .C1(n5460), .C2(keyinput_22), 
        .A(n5459), .ZN(n5492) );
  OAI22_X1 U6153 ( .A1(DATAI_14_), .A2(keyinput_17), .B1(keyinput_18), .B2(
        DATAI_13_), .ZN(n5461) );
  AOI221_X1 U6154 ( .B1(DATAI_14_), .B2(keyinput_17), .C1(DATAI_13_), .C2(
        keyinput_18), .A(n5461), .ZN(n5490) );
  INV_X1 U6155 ( .A(DATAI_18_), .ZN(n6791) );
  INV_X1 U6156 ( .A(keyinput_13), .ZN(n5481) );
  INV_X1 U6157 ( .A(DATAI_28_), .ZN(n6873) );
  OAI22_X1 U6158 ( .A1(n6873), .A2(keyinput_3), .B1(DATAI_29_), .B2(keyinput_2), .ZN(n5462) );
  AOI221_X1 U6159 ( .B1(n6873), .B2(keyinput_3), .C1(keyinput_2), .C2(
        DATAI_29_), .A(n5462), .ZN(n5468) );
  AOI22_X1 U6160 ( .A1(DATAI_30_), .A2(keyinput_1), .B1(DATAI_31_), .B2(
        keyinput_0), .ZN(n5463) );
  OAI221_X1 U6161 ( .B1(DATAI_30_), .B2(keyinput_1), .C1(DATAI_31_), .C2(
        keyinput_0), .A(n5463), .ZN(n5467) );
  INV_X1 U6162 ( .A(DATAI_27_), .ZN(n5465) );
  NAND3_X1 U6163 ( .A1(n5468), .A2(n5467), .A3(n5466), .ZN(n5469) );
  AOI21_X1 U6164 ( .B1(DATAI_27_), .B2(keyinput_4), .A(n5469), .ZN(n5474) );
  AOI22_X1 U6165 ( .A1(DATAI_24_), .A2(keyinput_7), .B1(DATAI_23_), .B2(
        keyinput_8), .ZN(n5470) );
  OAI221_X1 U6166 ( .B1(DATAI_24_), .B2(keyinput_7), .C1(DATAI_23_), .C2(
        keyinput_8), .A(n5470), .ZN(n5473) );
  AOI22_X1 U6167 ( .A1(DATAI_26_), .A2(keyinput_5), .B1(DATAI_25_), .B2(
        keyinput_6), .ZN(n5471) );
  OAI221_X1 U6168 ( .B1(DATAI_26_), .B2(keyinput_5), .C1(DATAI_25_), .C2(
        keyinput_6), .A(n5471), .ZN(n5472) );
  NOR3_X1 U6169 ( .A1(n5474), .A2(n5473), .A3(n5472), .ZN(n5479) );
  INV_X1 U6170 ( .A(DATAI_21_), .ZN(n6913) );
  INV_X1 U6171 ( .A(DATAI_19_), .ZN(n6832) );
  AOI22_X1 U6172 ( .A1(n6913), .A2(keyinput_10), .B1(keyinput_12), .B2(n6832), 
        .ZN(n5475) );
  OAI221_X1 U6173 ( .B1(n6913), .B2(keyinput_10), .C1(n6832), .C2(keyinput_12), 
        .A(n5475), .ZN(n5478) );
  AOI22_X1 U6174 ( .A1(DATAI_22_), .A2(keyinput_9), .B1(DATAI_20_), .B2(
        keyinput_11), .ZN(n5476) );
  OAI221_X1 U6175 ( .B1(DATAI_22_), .B2(keyinput_9), .C1(DATAI_20_), .C2(
        keyinput_11), .A(n5476), .ZN(n5477) );
  AOI221_X1 U6176 ( .B1(DATAI_18_), .B2(keyinput_13), .C1(n6791), .C2(n5481), 
        .A(n5480), .ZN(n5484) );
  INV_X1 U6177 ( .A(DATAI_16_), .ZN(n6551) );
  AOI22_X1 U6178 ( .A1(keyinput_16), .A2(DATAI_15_), .B1(n6551), .B2(
        keyinput_15), .ZN(n5482) );
  OAI221_X1 U6179 ( .B1(keyinput_16), .B2(DATAI_15_), .C1(n6551), .C2(
        keyinput_15), .A(n5482), .ZN(n5483) );
  OAI21_X1 U6180 ( .B1(DATAI_17_), .B2(keyinput_14), .A(n5485), .ZN(n5489) );
  AOI22_X1 U6181 ( .A1(n5487), .A2(keyinput_19), .B1(keyinput_20), .B2(n5592), 
        .ZN(n5486) );
  OAI221_X1 U6182 ( .B1(n5487), .B2(keyinput_19), .C1(n5592), .C2(keyinput_20), 
        .A(n5486), .ZN(n5488) );
  AOI21_X1 U6183 ( .B1(n5490), .B2(n5489), .A(n5488), .ZN(n5491) );
  OAI22_X1 U6184 ( .A1(n5492), .A2(n5491), .B1(keyinput_23), .B2(DATAI_8_), 
        .ZN(n5493) );
  AOI221_X1 U6185 ( .B1(DATAI_7_), .B2(n5495), .C1(n5601), .C2(keyinput_24), 
        .A(n5494), .ZN(n5502) );
  XNOR2_X1 U6186 ( .A(DATAI_6_), .B(keyinput_25), .ZN(n5501) );
  OAI22_X1 U6187 ( .A1(n5497), .A2(keyinput_27), .B1(n5604), .B2(keyinput_28), 
        .ZN(n5496) );
  AOI221_X1 U6188 ( .B1(n5497), .B2(keyinput_27), .C1(keyinput_28), .C2(n5604), 
        .A(n5496), .ZN(n5500) );
  OAI22_X1 U6189 ( .A1(n5603), .A2(keyinput_29), .B1(DATAI_5_), .B2(
        keyinput_26), .ZN(n5498) );
  AOI221_X1 U6190 ( .B1(n5603), .B2(keyinput_29), .C1(keyinput_26), .C2(
        DATAI_5_), .A(n5498), .ZN(n5499) );
  OAI211_X1 U6191 ( .C1(n5502), .C2(n5501), .A(n5500), .B(n5499), .ZN(n5503)
         );
  OAI221_X1 U6192 ( .B1(DATAI_1_), .B2(keyinput_30), .C1(n5612), .C2(n5504), 
        .A(n5503), .ZN(n5508) );
  INV_X1 U6193 ( .A(keyinput_31), .ZN(n5505) );
  OAI221_X1 U6194 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_32), .C1(n6511), 
        .C2(n5510), .A(n5509), .ZN(n5514) );
  INV_X1 U6195 ( .A(NA_N), .ZN(n6503) );
  INV_X1 U6196 ( .A(keyinput_33), .ZN(n5511) );
  OAI221_X1 U6197 ( .B1(BS16_N), .B2(keyinput_34), .C1(n5950), .C2(n5516), .A(
        n5515), .ZN(n5519) );
  INV_X1 U6198 ( .A(HOLD), .ZN(n6493) );
  OAI22_X1 U6199 ( .A1(n6493), .A2(keyinput_36), .B1(READY_N), .B2(keyinput_35), .ZN(n5517) );
  AOI221_X1 U6200 ( .B1(n6493), .B2(keyinput_36), .C1(keyinput_35), .C2(
        READY_N), .A(n5517), .ZN(n5518) );
  OAI21_X1 U6201 ( .B1(keyinput_37), .B2(READREQUEST_REG_SCAN_IN), .A(n5520), 
        .ZN(n5521) );
  OAI221_X1 U6202 ( .B1(keyinput_38), .B2(ADS_N_REG_SCAN_IN), .C1(n5522), .C2(
        n5954), .A(n5521), .ZN(n5523) );
  OAI221_X1 U6203 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n5524), .C1(n6132), .C2(
        keyinput_39), .A(n5523), .ZN(n5528) );
  XOR2_X1 U6204 ( .A(D_C_N_REG_SCAN_IN), .B(keyinput_41), .Z(n5527) );
  INV_X1 U6205 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6495) );
  AOI22_X1 U6206 ( .A1(n6495), .A2(keyinput_42), .B1(n6736), .B2(keyinput_43), 
        .ZN(n5525) );
  OAI221_X1 U6207 ( .B1(n6495), .B2(keyinput_42), .C1(n6736), .C2(keyinput_43), 
        .A(n5525), .ZN(n5526) );
  AOI221_X1 U6208 ( .B1(MORE_REG_SCAN_IN), .B2(n5531), .C1(n6450), .C2(
        keyinput_44), .A(n5530), .ZN(n5532) );
  AOI221_X1 U6209 ( .B1(FLUSH_REG_SCAN_IN), .B2(n5533), .C1(n6451), .C2(
        keyinput_45), .A(n5532), .ZN(n5534) );
  OAI22_X1 U6210 ( .A1(keyinput_48), .A2(n6056), .B1(n5535), .B2(n5534), .ZN(
        n5536) );
  AOI221_X1 U6211 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_49), .C1(
        n6053), .C2(n5538), .A(n5537), .ZN(n5539) );
  AOI221_X1 U6212 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_50), .C1(
        n5645), .C2(n5540), .A(n5539), .ZN(n5541) );
  OAI22_X1 U6213 ( .A1(n5542), .A2(n5541), .B1(keyinput_53), .B2(
        REIP_REG_29__SCAN_IN), .ZN(n5543) );
  AOI21_X1 U6214 ( .B1(keyinput_53), .B2(REIP_REG_29__SCAN_IN), .A(n5543), 
        .ZN(n5544) );
  OAI22_X1 U6215 ( .A1(keyinput_56), .A2(n6027), .B1(n5545), .B2(n5544), .ZN(
        n5546) );
  AOI221_X1 U6216 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5548), .C1(n6025), .C2(
        keyinput_57), .A(n5547), .ZN(n5549) );
  OAI22_X1 U6217 ( .A1(keyinput_60), .A2(n6402), .B1(n5550), .B2(n5549), .ZN(
        n5551) );
  AOI21_X1 U6218 ( .B1(keyinput_60), .B2(n6402), .A(n5551), .ZN(n5554) );
  INV_X1 U6219 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6401) );
  AOI22_X1 U6220 ( .A1(n6157), .A2(keyinput_63), .B1(n6401), .B2(keyinput_61), 
        .ZN(n5552) );
  OAI221_X1 U6221 ( .B1(n6157), .B2(keyinput_63), .C1(n6401), .C2(keyinput_61), 
        .A(n5552), .ZN(n5553) );
  OAI21_X1 U6222 ( .B1(keyinput_62), .B2(n6374), .A(n5555), .ZN(n5660) );
  OAI22_X1 U6223 ( .A1(n6401), .A2(keyinput_125), .B1(n6157), .B2(keyinput_127), .ZN(n5558) );
  INV_X1 U6224 ( .A(keyinput_127), .ZN(n5556) );
  NOR2_X1 U6225 ( .A1(n5556), .A2(REIP_REG_19__SCAN_IN), .ZN(n5557) );
  AOI211_X1 U6226 ( .C1(keyinput_125), .C2(n6401), .A(n5558), .B(n5557), .ZN(
        n5659) );
  OAI22_X1 U6227 ( .A1(REIP_REG_24__SCAN_IN), .A2(keyinput_122), .B1(
        REIP_REG_23__SCAN_IN), .B2(keyinput_123), .ZN(n5559) );
  AOI221_X1 U6228 ( .B1(REIP_REG_24__SCAN_IN), .B2(keyinput_122), .C1(
        keyinput_123), .C2(REIP_REG_23__SCAN_IN), .A(n5559), .ZN(n5655) );
  INV_X1 U6229 ( .A(keyinput_121), .ZN(n5653) );
  OAI22_X1 U6230 ( .A1(n5561), .A2(keyinput_118), .B1(REIP_REG_27__SCAN_IN), 
        .B2(keyinput_119), .ZN(n5560) );
  AOI221_X1 U6231 ( .B1(n5561), .B2(keyinput_118), .C1(keyinput_119), .C2(
        REIP_REG_27__SCAN_IN), .A(n5560), .ZN(n5650) );
  AOI22_X1 U6232 ( .A1(n6035), .A2(keyinput_116), .B1(n6039), .B2(keyinput_115), .ZN(n5562) );
  OAI221_X1 U6233 ( .B1(n6035), .B2(keyinput_116), .C1(n6039), .C2(
        keyinput_115), .A(n5562), .ZN(n5648) );
  INV_X1 U6234 ( .A(keyinput_114), .ZN(n5644) );
  INV_X1 U6235 ( .A(keyinput_113), .ZN(n5642) );
  AOI22_X1 U6236 ( .A1(BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput_111), .B1(
        n6141), .B2(keyinput_110), .ZN(n5563) );
  OAI221_X1 U6237 ( .B1(BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_111), .C1(
        n6141), .C2(keyinput_110), .A(n5563), .ZN(n5639) );
  INV_X1 U6238 ( .A(keyinput_109), .ZN(n5637) );
  INV_X1 U6239 ( .A(keyinput_108), .ZN(n5635) );
  OAI22_X1 U6240 ( .A1(n6736), .A2(keyinput_107), .B1(keyinput_105), .B2(
        D_C_N_REG_SCAN_IN), .ZN(n5564) );
  AOI221_X1 U6241 ( .B1(n6736), .B2(keyinput_107), .C1(D_C_N_REG_SCAN_IN), 
        .C2(keyinput_105), .A(n5564), .ZN(n5632) );
  INV_X1 U6242 ( .A(keyinput_104), .ZN(n5630) );
  INV_X1 U6243 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6510) );
  INV_X1 U6244 ( .A(keyinput_103), .ZN(n5628) );
  INV_X1 U6245 ( .A(keyinput_102), .ZN(n5626) );
  AOI22_X1 U6246 ( .A1(HOLD), .A2(keyinput_100), .B1(n6500), .B2(keyinput_99), 
        .ZN(n5565) );
  OAI221_X1 U6247 ( .B1(HOLD), .B2(keyinput_100), .C1(n6500), .C2(keyinput_99), 
        .A(n5565), .ZN(n5624) );
  INV_X1 U6248 ( .A(keyinput_98), .ZN(n5621) );
  INV_X1 U6249 ( .A(keyinput_97), .ZN(n5619) );
  INV_X1 U6250 ( .A(keyinput_96), .ZN(n5617) );
  INV_X1 U6251 ( .A(keyinput_95), .ZN(n5615) );
  INV_X1 U6252 ( .A(keyinput_94), .ZN(n5611) );
  XOR2_X1 U6253 ( .A(DATAI_6_), .B(keyinput_89), .Z(n5609) );
  INV_X1 U6254 ( .A(keyinput_88), .ZN(n5600) );
  OAI22_X1 U6255 ( .A1(n5567), .A2(keyinput_85), .B1(DATAI_9_), .B2(
        keyinput_86), .ZN(n5566) );
  AOI221_X1 U6256 ( .B1(n5567), .B2(keyinput_85), .C1(keyinput_86), .C2(
        DATAI_9_), .A(n5566), .ZN(n5597) );
  INV_X1 U6257 ( .A(DATAI_17_), .ZN(n6751) );
  INV_X1 U6258 ( .A(keyinput_77), .ZN(n5584) );
  INV_X1 U6259 ( .A(DATAI_29_), .ZN(n6915) );
  OAI22_X1 U6260 ( .A1(n6915), .A2(keyinput_66), .B1(keyinput_67), .B2(
        DATAI_28_), .ZN(n5568) );
  AOI221_X1 U6261 ( .B1(n6915), .B2(keyinput_66), .C1(DATAI_28_), .C2(
        keyinput_67), .A(n5568), .ZN(n5571) );
  AOI22_X1 U6262 ( .A1(DATAI_30_), .A2(keyinput_65), .B1(DATAI_31_), .B2(
        keyinput_64), .ZN(n5569) );
  OAI221_X1 U6263 ( .B1(DATAI_30_), .B2(keyinput_65), .C1(DATAI_31_), .C2(
        keyinput_64), .A(n5569), .ZN(n5570) );
  OAI211_X1 U6264 ( .C1(DATAI_27_), .C2(keyinput_68), .A(n5571), .B(n5570), 
        .ZN(n5572) );
  AOI21_X1 U6265 ( .B1(DATAI_27_), .B2(keyinput_68), .A(n5572), .ZN(n5577) );
  INV_X1 U6266 ( .A(DATAI_23_), .ZN(n7004) );
  INV_X1 U6267 ( .A(DATAI_25_), .ZN(n6749) );
  AOI22_X1 U6268 ( .A1(n7004), .A2(keyinput_72), .B1(n6749), .B2(keyinput_70), 
        .ZN(n5573) );
  OAI221_X1 U6269 ( .B1(n7004), .B2(keyinput_72), .C1(n6749), .C2(keyinput_70), 
        .A(n5573), .ZN(n5576) );
  INV_X1 U6270 ( .A(DATAI_24_), .ZN(n6540) );
  AOI22_X1 U6271 ( .A1(DATAI_26_), .A2(keyinput_69), .B1(n6540), .B2(
        keyinput_71), .ZN(n5574) );
  OAI221_X1 U6272 ( .B1(DATAI_26_), .B2(keyinput_69), .C1(n6540), .C2(
        keyinput_71), .A(n5574), .ZN(n5575) );
  NOR3_X1 U6273 ( .A1(n5577), .A2(n5576), .A3(n5575), .ZN(n5582) );
  INV_X1 U6274 ( .A(DATAI_22_), .ZN(n6956) );
  AOI22_X1 U6275 ( .A1(n6832), .A2(keyinput_76), .B1(n6956), .B2(keyinput_73), 
        .ZN(n5578) );
  OAI221_X1 U6276 ( .B1(n6832), .B2(keyinput_76), .C1(n6956), .C2(keyinput_73), 
        .A(n5578), .ZN(n5581) );
  AOI22_X1 U6277 ( .A1(DATAI_21_), .A2(keyinput_74), .B1(DATAI_20_), .B2(
        keyinput_75), .ZN(n5579) );
  OAI221_X1 U6278 ( .B1(DATAI_21_), .B2(keyinput_74), .C1(DATAI_20_), .C2(
        keyinput_75), .A(n5579), .ZN(n5580) );
  NOR3_X1 U6279 ( .A1(n5582), .A2(n5581), .A3(n5580), .ZN(n5583) );
  AOI221_X1 U6280 ( .B1(DATAI_18_), .B2(n5584), .C1(n6791), .C2(keyinput_77), 
        .A(n5583), .ZN(n5588) );
  OAI22_X1 U6281 ( .A1(n5674), .A2(keyinput_80), .B1(n6551), .B2(keyinput_79), 
        .ZN(n5585) );
  AOI221_X1 U6282 ( .B1(n5674), .B2(keyinput_80), .C1(keyinput_79), .C2(n6551), 
        .A(n5585), .ZN(n5586) );
  OAI21_X1 U6283 ( .B1(keyinput_78), .B2(n6751), .A(n5586), .ZN(n5587) );
  AOI211_X1 U6284 ( .C1(keyinput_78), .C2(n6751), .A(n5588), .B(n5587), .ZN(
        n5595) );
  AOI22_X1 U6285 ( .A1(DATAI_14_), .A2(keyinput_81), .B1(n5590), .B2(
        keyinput_82), .ZN(n5589) );
  OAI221_X1 U6286 ( .B1(DATAI_14_), .B2(keyinput_81), .C1(n5590), .C2(
        keyinput_82), .A(n5589), .ZN(n5594) );
  OAI22_X1 U6287 ( .A1(n5592), .A2(keyinput_84), .B1(DATAI_12_), .B2(
        keyinput_83), .ZN(n5591) );
  AOI221_X1 U6288 ( .B1(n5592), .B2(keyinput_84), .C1(keyinput_83), .C2(
        DATAI_12_), .A(n5591), .ZN(n5593) );
  OAI21_X1 U6289 ( .B1(n5595), .B2(n5594), .A(n5593), .ZN(n5596) );
  AOI22_X1 U6290 ( .A1(n5597), .A2(n5596), .B1(keyinput_87), .B2(DATAI_8_), 
        .ZN(n5598) );
  OAI21_X1 U6291 ( .B1(keyinput_87), .B2(DATAI_8_), .A(n5598), .ZN(n5599) );
  OAI221_X1 U6292 ( .B1(DATAI_7_), .B2(keyinput_88), .C1(n5601), .C2(n5600), 
        .A(n5599), .ZN(n5608) );
  AOI22_X1 U6293 ( .A1(n5604), .A2(keyinput_92), .B1(n5603), .B2(keyinput_93), 
        .ZN(n5602) );
  OAI221_X1 U6294 ( .B1(n5604), .B2(keyinput_92), .C1(n5603), .C2(keyinput_93), 
        .A(n5602), .ZN(n5607) );
  AOI22_X1 U6295 ( .A1(DATAI_4_), .A2(keyinput_91), .B1(DATAI_5_), .B2(
        keyinput_90), .ZN(n5605) );
  OAI221_X1 U6296 ( .B1(DATAI_4_), .B2(keyinput_91), .C1(DATAI_5_), .C2(
        keyinput_90), .A(n5605), .ZN(n5606) );
  AOI211_X1 U6297 ( .C1(n5609), .C2(n5608), .A(n5607), .B(n5606), .ZN(n5610)
         );
  AOI221_X1 U6298 ( .B1(DATAI_1_), .B2(keyinput_94), .C1(n5612), .C2(n5611), 
        .A(n5610), .ZN(n5613) );
  AOI221_X1 U6299 ( .B1(DATAI_0_), .B2(n5615), .C1(n5614), .C2(keyinput_95), 
        .A(n5613), .ZN(n5616) );
  AOI221_X1 U6300 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n5617), .C1(n6511), .C2(
        keyinput_96), .A(n5616), .ZN(n5618) );
  AOI221_X1 U6301 ( .B1(NA_N), .B2(n5619), .C1(n6503), .C2(keyinput_97), .A(
        n5618), .ZN(n5620) );
  AOI221_X1 U6302 ( .B1(BS16_N), .B2(n5621), .C1(n5950), .C2(keyinput_98), .A(
        n5620), .ZN(n5623) );
  NAND2_X1 U6303 ( .A1(READREQUEST_REG_SCAN_IN), .A2(keyinput_101), .ZN(n5622)
         );
  OAI221_X1 U6304 ( .B1(n5624), .B2(n5623), .C1(READREQUEST_REG_SCAN_IN), .C2(
        keyinput_101), .A(n5622), .ZN(n5625) );
  OAI221_X1 U6305 ( .B1(ADS_N_REG_SCAN_IN), .B2(keyinput_102), .C1(n5954), 
        .C2(n5626), .A(n5625), .ZN(n5627) );
  OAI221_X1 U6306 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(keyinput_103), .C1(n6132), 
        .C2(n5628), .A(n5627), .ZN(n5629) );
  OAI221_X1 U6307 ( .B1(M_IO_N_REG_SCAN_IN), .B2(n5630), .C1(n6510), .C2(
        keyinput_104), .A(n5629), .ZN(n5631) );
  OAI211_X1 U6308 ( .C1(REQUESTPENDING_REG_SCAN_IN), .C2(keyinput_106), .A(
        n5632), .B(n5631), .ZN(n5633) );
  AOI21_X1 U6309 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_106), .A(
        n5633), .ZN(n5634) );
  AOI221_X1 U6310 ( .B1(MORE_REG_SCAN_IN), .B2(n5635), .C1(n6450), .C2(
        keyinput_108), .A(n5634), .ZN(n5636) );
  AOI221_X1 U6311 ( .B1(FLUSH_REG_SCAN_IN), .B2(keyinput_109), .C1(n6451), 
        .C2(n5637), .A(n5636), .ZN(n5638) );
  OAI22_X1 U6312 ( .A1(n5639), .A2(n5638), .B1(keyinput_112), .B2(
        BYTEENABLE_REG_1__SCAN_IN), .ZN(n5640) );
  AOI21_X1 U6313 ( .B1(keyinput_112), .B2(BYTEENABLE_REG_1__SCAN_IN), .A(n5640), .ZN(n5641) );
  AOI221_X1 U6314 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(n5642), .C1(n6053), 
        .C2(keyinput_113), .A(n5641), .ZN(n5643) );
  AOI221_X1 U6315 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_114), .C1(
        n5645), .C2(n5644), .A(n5643), .ZN(n5647) );
  NAND2_X1 U6316 ( .A1(n6033), .A2(keyinput_117), .ZN(n5646) );
  OAI221_X1 U6317 ( .B1(n5648), .B2(n5647), .C1(n6033), .C2(keyinput_117), .A(
        n5646), .ZN(n5649) );
  AOI22_X1 U6318 ( .A1(n5650), .A2(n5649), .B1(keyinput_120), .B2(
        REIP_REG_26__SCAN_IN), .ZN(n5651) );
  OAI21_X1 U6319 ( .B1(keyinput_120), .B2(REIP_REG_26__SCAN_IN), .A(n5651), 
        .ZN(n5652) );
  OAI221_X1 U6320 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5653), .C1(n6025), .C2(
        keyinput_121), .A(n5652), .ZN(n5654) );
  AOI22_X1 U6321 ( .A1(n5655), .A2(n5654), .B1(keyinput_124), .B2(
        REIP_REG_22__SCAN_IN), .ZN(n5656) );
  OAI21_X1 U6322 ( .B1(REIP_REG_22__SCAN_IN), .B2(keyinput_124), .A(n5656), 
        .ZN(n5658) );
  XNOR2_X1 U6323 ( .A(REIP_REG_20__SCAN_IN), .B(keyinput_126), .ZN(n5657) );
  NAND4_X1 U6324 ( .A1(n5660), .A2(n5659), .A3(n5658), .A4(n5657), .ZN(n5665)
         );
  AOI22_X1 U6325 ( .A1(n6533), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n6536), .ZN(n5662) );
  NAND2_X1 U6326 ( .A1(n6537), .A2(DATAI_11_), .ZN(n5661) );
  XNOR2_X1 U6327 ( .A(n5665), .B(n5664), .ZN(U2864) );
  AOI22_X1 U6328 ( .A1(n6533), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6536), .ZN(n5667) );
  NAND2_X1 U6329 ( .A1(n6537), .A2(DATAI_10_), .ZN(n5666) );
  OAI211_X1 U6330 ( .C1(n5721), .C2(n5678), .A(n5667), .B(n5666), .ZN(U2865)
         );
  NAND2_X1 U6331 ( .A1(n5748), .A2(n6534), .ZN(n5669) );
  AOI22_X1 U6332 ( .A1(n6533), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6536), .ZN(n5668) );
  OAI211_X1 U6333 ( .C1(n6516), .C2(n4818), .A(n5669), .B(n5668), .ZN(U2867)
         );
  AOI22_X1 U6334 ( .A1(n6533), .A2(DATAI_20_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n6536), .ZN(n5671) );
  NAND2_X1 U6335 ( .A1(n6537), .A2(DATAI_4_), .ZN(n5670) );
  OAI211_X1 U6336 ( .C1(n6378), .C2(n5678), .A(n5671), .B(n5670), .ZN(U2871)
         );
  AOI22_X1 U6337 ( .A1(n6533), .A2(DATAI_16_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n6536), .ZN(n5673) );
  NAND2_X1 U6338 ( .A1(n6537), .A2(DATAI_0_), .ZN(n5672) );
  OAI211_X1 U6339 ( .C1(n5799), .C2(n5678), .A(n5673), .B(n5672), .ZN(U2875)
         );
  INV_X1 U6340 ( .A(EAX_REG_15__SCAN_IN), .ZN(n5988) );
  OAI222_X1 U6341 ( .A1(n5675), .A2(n5678), .B1(n5677), .B2(n5674), .C1(n6514), 
        .C2(n5988), .ZN(U2876) );
  INV_X1 U6342 ( .A(EAX_REG_14__SCAN_IN), .ZN(n5985) );
  OAI222_X1 U6343 ( .A1(n5814), .A2(n5678), .B1(n5677), .B2(n5676), .C1(n6514), 
        .C2(n5985), .ZN(U2877) );
  AOI21_X1 U6344 ( .B1(n6123), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5679), 
        .ZN(n5680) );
  OAI21_X1 U6345 ( .B1(n6122), .B2(n5681), .A(n5680), .ZN(n5682) );
  AOI21_X1 U6346 ( .B1(n5683), .B2(n5804), .A(n5682), .ZN(n5684) );
  OAI21_X1 U6347 ( .B1(n5685), .B2(n6424), .A(n5684), .ZN(U2955) );
  INV_X1 U6348 ( .A(n5686), .ZN(n5687) );
  NAND2_X1 U6349 ( .A1(n5688), .A2(n5687), .ZN(n5690) );
  NAND2_X1 U6350 ( .A1(n5692), .A2(n4143), .ZN(n5689) );
  NAND2_X1 U6351 ( .A1(n5690), .A2(n5689), .ZN(n5694) );
  XNOR2_X1 U6352 ( .A(n5692), .B(n5691), .ZN(n5693) );
  XNOR2_X1 U6353 ( .A(n5694), .B(n5693), .ZN(n5838) );
  AND2_X1 U6354 ( .A1(n6277), .A2(REIP_REG_29__SCAN_IN), .ZN(n5832) );
  AOI21_X1 U6355 ( .B1(n6123), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5832), 
        .ZN(n5695) );
  OAI21_X1 U6356 ( .B1(n6122), .B2(n5696), .A(n5695), .ZN(n5697) );
  AOI21_X1 U6357 ( .B1(n5698), .B2(n5804), .A(n5697), .ZN(n5699) );
  OAI21_X1 U6358 ( .B1(n6424), .B2(n5838), .A(n5699), .ZN(U2957) );
  INV_X1 U6359 ( .A(n5700), .ZN(n5703) );
  AOI21_X1 U6360 ( .B1(n6123), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5701), 
        .ZN(n5702) );
  OAI21_X1 U6361 ( .B1(n6122), .B2(n5703), .A(n5702), .ZN(n5704) );
  AOI21_X1 U6362 ( .B1(n5705), .B2(n5804), .A(n5704), .ZN(n5706) );
  OAI21_X1 U6363 ( .B1(n5707), .B2(n6424), .A(n5706), .ZN(U2958) );
  OR2_X1 U6364 ( .A1(n5692), .A2(n5708), .ZN(n5718) );
  NAND2_X1 U6365 ( .A1(n5709), .A2(n5718), .ZN(n5711) );
  XNOR2_X1 U6366 ( .A(n4095), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5710)
         );
  XNOR2_X1 U6367 ( .A(n5711), .B(n5710), .ZN(n5847) );
  AND2_X1 U6368 ( .A1(n6277), .A2(REIP_REG_27__SCAN_IN), .ZN(n5840) );
  AOI21_X1 U6369 ( .B1(n6123), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5840), 
        .ZN(n5712) );
  OAI21_X1 U6370 ( .B1(n6122), .B2(n5713), .A(n5712), .ZN(n5714) );
  AOI21_X1 U6371 ( .B1(n5715), .B2(n5804), .A(n5714), .ZN(n5716) );
  OAI21_X1 U6372 ( .B1(n5847), .B2(n6424), .A(n5716), .ZN(U2959) );
  NAND2_X1 U6373 ( .A1(n5718), .A2(n5717), .ZN(n5720) );
  XOR2_X1 U6374 ( .A(n5720), .B(n5719), .Z(n5856) );
  INV_X1 U6375 ( .A(n5721), .ZN(n5726) );
  INV_X1 U6376 ( .A(n5722), .ZN(n5724) );
  AND2_X1 U6377 ( .A1(n6277), .A2(REIP_REG_26__SCAN_IN), .ZN(n5851) );
  AOI21_X1 U6378 ( .B1(n6123), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5851), 
        .ZN(n5723) );
  OAI21_X1 U6379 ( .B1(n6122), .B2(n5724), .A(n5723), .ZN(n5725) );
  AOI21_X1 U6380 ( .B1(n5726), .B2(n5804), .A(n5725), .ZN(n5727) );
  OAI21_X1 U6381 ( .B1(n6424), .B2(n5856), .A(n5727), .ZN(U2960) );
  XOR2_X1 U6382 ( .A(n5730), .B(n5729), .Z(n6278) );
  AOI22_X1 U6383 ( .A1(n6123), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .B1(n6277), 
        .B2(REIP_REG_25__SCAN_IN), .ZN(n5731) );
  OAI21_X1 U6384 ( .B1(n6122), .B2(n5732), .A(n5731), .ZN(n5733) );
  INV_X1 U6385 ( .A(n5733), .ZN(n5734) );
  INV_X1 U6386 ( .A(n5736), .ZN(n5737) );
  OAI21_X1 U6387 ( .B1(n6424), .B2(n6278), .A(n5737), .ZN(U2961) );
  INV_X1 U6388 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6159) );
  XNOR2_X1 U6389 ( .A(n4095), .B(n6159), .ZN(n6125) );
  OR2_X2 U6390 ( .A1(n3446), .A2(n6125), .ZN(n6126) );
  INV_X1 U6391 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5774) );
  NOR2_X1 U6392 ( .A1(n5692), .A2(n5774), .ZN(n5738) );
  OAI22_X1 U6393 ( .A1(n6126), .A2(n5738), .B1(n5782), .B2(n5893), .ZN(n5768)
         );
  INV_X1 U6394 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5890) );
  XNOR2_X1 U6395 ( .A(n4095), .B(n5890), .ZN(n5767) );
  NAND2_X1 U6396 ( .A1(n5782), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5739) );
  NAND3_X1 U6397 ( .A1(n5692), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5742) );
  INV_X1 U6398 ( .A(n6126), .ZN(n5741) );
  NAND4_X1 U6399 ( .A1(n5741), .A2(n5782), .A3(n5740), .A4(n5774), .ZN(n5751)
         );
  OAI22_X1 U6400 ( .A1(n5759), .A2(n5742), .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5751), .ZN(n5743) );
  XNOR2_X1 U6401 ( .A(n5743), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5864)
         );
  INV_X1 U6402 ( .A(n5744), .ZN(n5746) );
  AND2_X1 U6403 ( .A1(n6277), .A2(REIP_REG_24__SCAN_IN), .ZN(n5861) );
  AOI21_X1 U6404 ( .B1(n6123), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5861), 
        .ZN(n5745) );
  OAI21_X1 U6405 ( .B1(n6122), .B2(n5746), .A(n5745), .ZN(n5747) );
  AOI21_X1 U6406 ( .B1(n5748), .B2(n5804), .A(n5747), .ZN(n5749) );
  OAI21_X1 U6407 ( .B1(n5864), .B2(n6424), .A(n5749), .ZN(U2962) );
  NAND3_X1 U6408 ( .A1(n5692), .A2(n5866), .A3(n5893), .ZN(n5752) );
  OAI21_X1 U6409 ( .B1(n5750), .B2(n5752), .A(n5751), .ZN(n5753) );
  XNOR2_X1 U6410 ( .A(n5753), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5871)
         );
  NAND2_X1 U6411 ( .A1(n6277), .A2(REIP_REG_23__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U6412 ( .A1(n6123), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5754)
         );
  OAI211_X1 U6413 ( .C1(n6122), .C2(n6411), .A(n5867), .B(n5754), .ZN(n5755)
         );
  AOI21_X1 U6414 ( .B1(n6535), .B2(n5804), .A(n5755), .ZN(n5756) );
  OAI21_X1 U6415 ( .B1(n5871), .B2(n6424), .A(n5756), .ZN(U2963) );
  XNOR2_X1 U6416 ( .A(n4095), .B(n5757), .ZN(n5758) );
  XNOR2_X1 U6417 ( .A(n5759), .B(n5758), .ZN(n5880) );
  NAND2_X1 U6418 ( .A1(n6277), .A2(REIP_REG_22__SCAN_IN), .ZN(n5873) );
  OAI21_X1 U6419 ( .B1(n6101), .B2(n5760), .A(n5873), .ZN(n5762) );
  NOR2_X1 U6420 ( .A1(n6399), .A2(n7005), .ZN(n5761) );
  OAI21_X1 U6421 ( .B1(n5880), .B2(n6424), .A(n5763), .ZN(U2964) );
  NOR2_X1 U6422 ( .A1(n5426), .A2(n5764), .ZN(n5765) );
  OR2_X1 U6423 ( .A1(n5414), .A2(n5765), .ZN(n6526) );
  NAND2_X1 U6424 ( .A1(n5768), .A2(n5767), .ZN(n5881) );
  NAND3_X1 U6425 ( .A1(n5766), .A2(n6128), .A3(n5881), .ZN(n5772) );
  NAND2_X1 U6426 ( .A1(n6277), .A2(REIP_REG_21__SCAN_IN), .ZN(n5885) );
  INV_X1 U6427 ( .A(n5885), .ZN(n5770) );
  NOR2_X1 U6428 ( .A1(n6122), .A2(n6387), .ZN(n5769) );
  AOI211_X1 U6429 ( .C1(n6123), .C2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5770), 
        .B(n5769), .ZN(n5771) );
  OAI211_X1 U6430 ( .C1(n7005), .C2(n6526), .A(n5772), .B(n5771), .ZN(U2965)
         );
  NAND2_X1 U6431 ( .A1(n6126), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5773) );
  MUX2_X1 U6432 ( .A(n5773), .B(n6126), .S(n5782), .Z(n5775) );
  XNOR2_X1 U6433 ( .A(n5775), .B(n5774), .ZN(n5899) );
  INV_X1 U6434 ( .A(n6369), .ZN(n5777) );
  NAND2_X1 U6435 ( .A1(n6123), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5776)
         );
  NAND2_X1 U6436 ( .A1(n6277), .A2(REIP_REG_20__SCAN_IN), .ZN(n5892) );
  OAI211_X1 U6437 ( .C1(n6122), .C2(n5777), .A(n5776), .B(n5892), .ZN(n5778)
         );
  AOI21_X1 U6438 ( .B1(n5779), .B2(n5804), .A(n5778), .ZN(n5780) );
  OAI21_X1 U6439 ( .B1(n5899), .B2(n6424), .A(n5780), .ZN(U2966) );
  INV_X1 U6440 ( .A(n5781), .ZN(n5784) );
  NAND2_X1 U6441 ( .A1(n5692), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6115) );
  AOI21_X1 U6442 ( .B1(n5782), .B2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5781), 
        .ZN(n6114) );
  OR2_X1 U6443 ( .A1(n5692), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6113)
         );
  INV_X1 U6444 ( .A(n6113), .ZN(n5783) );
  NAND2_X1 U6445 ( .A1(n6114), .A2(n5783), .ZN(n6117) );
  OAI21_X1 U6446 ( .B1(n5784), .B2(n6115), .A(n6117), .ZN(n5785) );
  XNOR2_X1 U6447 ( .A(n5785), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5914)
         );
  INV_X1 U6448 ( .A(n5786), .ZN(n5788) );
  AOI22_X1 U6449 ( .A1(n6123), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .B1(n6277), 
        .B2(REIP_REG_18__SCAN_IN), .ZN(n5787) );
  OAI21_X1 U6450 ( .B1(n6122), .B2(n5788), .A(n5787), .ZN(n5789) );
  AOI21_X1 U6451 ( .B1(n6520), .B2(n5804), .A(n5789), .ZN(n5790) );
  OAI21_X1 U6452 ( .B1(n5914), .B2(n6424), .A(n5790), .ZN(U2968) );
  XNOR2_X1 U6453 ( .A(n4095), .B(n6262), .ZN(n5792) );
  XNOR2_X1 U6454 ( .A(n5791), .B(n5792), .ZN(n6259) );
  NAND2_X1 U6455 ( .A1(n6259), .A2(n6128), .ZN(n5798) );
  INV_X1 U6456 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5793) );
  NOR2_X1 U6457 ( .A1(n6269), .A2(n5793), .ZN(n6256) );
  INV_X1 U6458 ( .A(n5794), .ZN(n5795) );
  NOR2_X1 U6459 ( .A1(n6122), .A2(n5795), .ZN(n5796) );
  AOI211_X1 U6460 ( .C1(n6123), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6256), 
        .B(n5796), .ZN(n5797) );
  OAI211_X1 U6461 ( .C1(n7005), .C2(n5799), .A(n5798), .B(n5797), .ZN(U2970)
         );
  NAND2_X1 U6462 ( .A1(n5800), .A2(n5810), .ZN(n5803) );
  NOR2_X1 U6463 ( .A1(n5801), .A2(n3463), .ZN(n5802) );
  XNOR2_X1 U6464 ( .A(n5803), .B(n5802), .ZN(n5922) );
  NAND2_X1 U6465 ( .A1(n6354), .A2(n5804), .ZN(n5808) );
  INV_X1 U6466 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5805) );
  NOR2_X1 U6467 ( .A1(n6269), .A2(n5805), .ZN(n5919) );
  AND2_X1 U6468 ( .A1(n6123), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5806)
         );
  AOI211_X1 U6469 ( .C1(n5826), .C2(n6353), .A(n5919), .B(n5806), .ZN(n5807)
         );
  OAI211_X1 U6470 ( .C1(n5922), .C2(n6424), .A(n5808), .B(n5807), .ZN(U2971)
         );
  INV_X1 U6471 ( .A(n5810), .ZN(n5812) );
  NOR2_X1 U6472 ( .A1(n5812), .A2(n5811), .ZN(n5813) );
  XNOR2_X1 U6473 ( .A(n5809), .B(n5813), .ZN(n6175) );
  INV_X1 U6474 ( .A(n6175), .ZN(n5820) );
  INV_X1 U6475 ( .A(n5814), .ZN(n5818) );
  AOI22_X1 U6476 ( .A1(n6123), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6277), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5815) );
  OAI21_X1 U6477 ( .B1(n6122), .B2(n5816), .A(n5815), .ZN(n5817) );
  AOI21_X1 U6478 ( .B1(n5818), .B2(n5804), .A(n5817), .ZN(n5819) );
  OAI21_X1 U6479 ( .B1(n5820), .B2(n6424), .A(n5819), .ZN(U2972) );
  XNOR2_X1 U6480 ( .A(n5821), .B(n5822), .ZN(n6170) );
  NAND2_X1 U6481 ( .A1(n6170), .A2(n6128), .ZN(n5828) );
  NAND2_X1 U6482 ( .A1(n6277), .A2(REIP_REG_13__SCAN_IN), .ZN(n6166) );
  OAI21_X1 U6483 ( .B1(n6101), .B2(n5823), .A(n6166), .ZN(n5824) );
  AOI21_X1 U6484 ( .B1(n5826), .B2(n5825), .A(n5824), .ZN(n5827) );
  OAI211_X1 U6485 ( .C1(n5829), .C2(n7005), .A(n5828), .B(n5827), .ZN(U2973)
         );
  INV_X1 U6486 ( .A(n5834), .ZN(n5830) );
  NOR3_X1 U6487 ( .A1(n5843), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5830), 
        .ZN(n5831) );
  AOI211_X1 U6488 ( .C1(n5833), .C2(n6280), .A(n5832), .B(n5831), .ZN(n5837)
         );
  OAI21_X1 U6489 ( .B1(n5834), .B2(n5917), .A(n5839), .ZN(n5835) );
  NAND2_X1 U6490 ( .A1(n5835), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5836) );
  OAI211_X1 U6491 ( .C1(n5838), .C2(n6223), .A(n5837), .B(n5836), .ZN(U2989)
         );
  INV_X1 U6492 ( .A(n5839), .ZN(n5845) );
  AOI21_X1 U6493 ( .B1(n5841), .B2(n6280), .A(n5840), .ZN(n5842) );
  OAI21_X1 U6494 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5843), .A(n5842), 
        .ZN(n5844) );
  AOI21_X1 U6495 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5845), .A(n5844), 
        .ZN(n5846) );
  OAI21_X1 U6496 ( .B1(n5847), .B2(n6223), .A(n5846), .ZN(U2991) );
  AOI21_X1 U6497 ( .B1(n6285), .B2(n5708), .A(n5848), .ZN(n5853) );
  NOR2_X1 U6498 ( .A1(n5849), .A2(n6227), .ZN(n5850) );
  AOI211_X1 U6499 ( .C1(n5853), .C2(n5852), .A(n5851), .B(n5850), .ZN(n5855)
         );
  NAND2_X1 U6500 ( .A1(n5857), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5854) );
  OAI211_X1 U6501 ( .C1(n5856), .C2(n6223), .A(n5855), .B(n5854), .ZN(U2992)
         );
  NAND3_X1 U6502 ( .A1(n5887), .A2(n5866), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5858) );
  INV_X1 U6503 ( .A(n5857), .ZN(n6286) );
  AOI21_X1 U6504 ( .B1(n5859), .B2(n5858), .A(n6286), .ZN(n5860) );
  AOI211_X1 U6505 ( .C1(n6280), .C2(n5862), .A(n5861), .B(n5860), .ZN(n5863)
         );
  OAI21_X1 U6506 ( .B1(n5864), .B2(n6223), .A(n5863), .ZN(U2994) );
  NAND3_X1 U6507 ( .A1(n5887), .A2(n5866), .A3(n5865), .ZN(n5868) );
  OAI211_X1 U6508 ( .C1(n6227), .C2(n6416), .A(n5868), .B(n5867), .ZN(n5869)
         );
  AOI21_X1 U6509 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5877), .A(n5869), 
        .ZN(n5870) );
  OAI21_X1 U6510 ( .B1(n5871), .B2(n6223), .A(n5870), .ZN(U2995) );
  INV_X1 U6511 ( .A(n5872), .ZN(n5876) );
  OAI21_X1 U6512 ( .B1(n5874), .B2(n6227), .A(n5873), .ZN(n5875) );
  AOI21_X1 U6513 ( .B1(n5876), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5875), 
        .ZN(n5879) );
  NAND2_X1 U6514 ( .A1(n5877), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5878) );
  OAI211_X1 U6515 ( .C1(n5880), .C2(n6223), .A(n5879), .B(n5878), .ZN(U2996)
         );
  NAND3_X1 U6516 ( .A1(n5766), .A2(n6281), .A3(n5881), .ZN(n5889) );
  OR2_X1 U6517 ( .A1(n5422), .A2(n5882), .ZN(n5883) );
  NAND2_X1 U6518 ( .A1(n5884), .A2(n5883), .ZN(n6389) );
  OAI21_X1 U6519 ( .B1(n6389), .B2(n6227), .A(n5885), .ZN(n5886) );
  AOI21_X1 U6520 ( .B1(n5887), .B2(n5890), .A(n5886), .ZN(n5888) );
  OAI211_X1 U6521 ( .C1(n5891), .C2(n5890), .A(n5889), .B(n5888), .ZN(U2997)
         );
  INV_X1 U6522 ( .A(n6158), .ZN(n5897) );
  OAI21_X1 U6523 ( .B1(n6377), .B2(n6227), .A(n5892), .ZN(n5896) );
  NOR3_X1 U6524 ( .A1(n6164), .A2(n5894), .A3(n5893), .ZN(n5895) );
  AOI211_X1 U6525 ( .C1(INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n5897), .A(n5896), .B(n5895), .ZN(n5898) );
  OAI21_X1 U6526 ( .B1(n5899), .B2(n6223), .A(n5898), .ZN(U2998) );
  INV_X1 U6527 ( .A(n6199), .ZN(n6220) );
  INV_X1 U6528 ( .A(n5900), .ZN(n5902) );
  OAI21_X1 U6529 ( .B1(n6272), .B2(n5902), .A(n5901), .ZN(n5903) );
  OAI211_X1 U6530 ( .C1(n6220), .C2(n5904), .A(n5903), .B(n6196), .ZN(n6271)
         );
  INV_X1 U6531 ( .A(n6271), .ZN(n5906) );
  AOI221_X1 U6532 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5906), .C1(
        n5905), .C2(n5906), .A(n5908), .ZN(n5912) );
  NOR2_X1 U6533 ( .A1(n6249), .A2(n5907), .ZN(n6273) );
  AND3_X1 U6534 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6273), .A3(n5908), 
        .ZN(n5911) );
  OAI22_X1 U6535 ( .A1(n6227), .A2(n5909), .B1(n6016), .B2(n6269), .ZN(n5910)
         );
  NOR3_X1 U6536 ( .A1(n5912), .A2(n5911), .A3(n5910), .ZN(n5913) );
  OAI21_X1 U6537 ( .B1(n5914), .B2(n6223), .A(n5913), .ZN(U3000) );
  OAI21_X1 U6538 ( .B1(n5917), .B2(n5916), .A(n5915), .ZN(n6258) );
  NOR3_X1 U6539 ( .A1(n6249), .A2(n6174), .A3(n6179), .ZN(n6260) );
  AOI22_X1 U6540 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n6258), .B1(n6260), .B2(n6261), .ZN(n5921) );
  INV_X1 U6541 ( .A(n5918), .ZN(n6347) );
  AOI21_X1 U6542 ( .B1(n6280), .B2(n6347), .A(n5919), .ZN(n5920) );
  OAI211_X1 U6543 ( .C1(n5922), .C2(n6223), .A(n5921), .B(n5920), .ZN(U3003)
         );
  NAND2_X1 U6544 ( .A1(n5923), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5933)
         );
  XNOR2_X1 U6545 ( .A(n5925), .B(n5929), .ZN(n5926) );
  XNOR2_X1 U6546 ( .A(n5924), .B(n5926), .ZN(n6086) );
  OAI22_X1 U6547 ( .A1(n6223), .A2(n6086), .B1(n4836), .B2(n6269), .ZN(n5927)
         );
  AOI21_X1 U6548 ( .B1(n6280), .B2(n5928), .A(n5927), .ZN(n5932) );
  NAND3_X1 U6549 ( .A1(n6165), .A2(n5930), .A3(n5929), .ZN(n5931) );
  NAND3_X1 U6550 ( .A1(n5933), .A2(n5932), .A3(n5931), .ZN(U3017) );
  NAND3_X1 U6551 ( .A1(n5935), .A2(n5934), .A3(n5942), .ZN(n5936) );
  OAI21_X1 U6552 ( .B1(n5937), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n5936), 
        .ZN(n5938) );
  AOI21_X1 U6553 ( .B1(n4800), .B2(n5939), .A(n5938), .ZN(n6435) );
  NOR2_X1 U6554 ( .A1(n6475), .A2(n5940), .ZN(n5944) );
  INV_X1 U6555 ( .A(n5941), .ZN(n5943) );
  AOI22_X1 U6556 ( .A1(n5945), .A2(n5944), .B1(n5943), .B2(n5942), .ZN(n5946)
         );
  OAI21_X1 U6557 ( .B1(n6435), .B2(n5947), .A(n5946), .ZN(n5949) );
  MUX2_X1 U6558 ( .A(n5949), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(n5948), 
        .Z(U3460) );
  INV_X1 U6559 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5951) );
  INV_X1 U6560 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6501) );
  INV_X1 U6561 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6142) );
  AOI21_X1 U6562 ( .B1(n6142), .B2(STATE_REG_1__SCAN_IN), .A(n6501), .ZN(n5955) );
  NAND2_X1 U6563 ( .A1(n6142), .A2(n6501), .ZN(n6136) );
  AOI21_X1 U6564 ( .B1(n5950), .B2(n6136), .A(n5952), .ZN(n6490) );
  AOI21_X1 U6565 ( .B1(n5951), .B2(n5952), .A(n6490), .ZN(U3451) );
  AND2_X1 U6566 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n5952), .ZN(U3180) );
  AND2_X1 U6567 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n5952), .ZN(U3179) );
  AND2_X1 U6568 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n5952), .ZN(U3178) );
  AND2_X1 U6569 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n5952), .ZN(U3177) );
  AND2_X1 U6570 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n5952), .ZN(U3176) );
  AND2_X1 U6571 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n5952), .ZN(U3175) );
  AND2_X1 U6572 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n5952), .ZN(U3174) );
  AND2_X1 U6573 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n5952), .ZN(U3173) );
  AND2_X1 U6574 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n5952), .ZN(U3172) );
  AND2_X1 U6575 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n5952), .ZN(U3171) );
  AND2_X1 U6576 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n5952), .ZN(U3170) );
  AND2_X1 U6577 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n5952), .ZN(U3169) );
  AND2_X1 U6578 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n5952), .ZN(U3168) );
  AND2_X1 U6579 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n5952), .ZN(U3167) );
  AND2_X1 U6580 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n5952), .ZN(U3166) );
  AND2_X1 U6581 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n5952), .ZN(U3165) );
  AND2_X1 U6582 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n5952), .ZN(U3164) );
  AND2_X1 U6583 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n5952), .ZN(U3163) );
  AND2_X1 U6584 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n5952), .ZN(U3162) );
  AND2_X1 U6585 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n5952), .ZN(U3161) );
  AND2_X1 U6586 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n5952), .ZN(U3160) );
  AND2_X1 U6587 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n5952), .ZN(U3159) );
  AND2_X1 U6588 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n5952), .ZN(U3158) );
  AND2_X1 U6589 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n5952), .ZN(U3157) );
  AND2_X1 U6590 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n5952), .ZN(U3156) );
  AND2_X1 U6591 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n5952), .ZN(U3155) );
  AND2_X1 U6592 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n5952), .ZN(U3154) );
  AND2_X1 U6593 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n5952), .ZN(U3153) );
  AND2_X1 U6594 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n5952), .ZN(U3152) );
  AND2_X1 U6595 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n5952), .ZN(U3151) );
  AND2_X1 U6596 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n5953), .ZN(U3019)
         );
  AND2_X1 U6597 ( .A1(n5969), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI21_X1 U6598 ( .B1(n5955), .B2(n5954), .A(n6512), .ZN(U2789) );
  AOI22_X1 U6599 ( .A1(n6154), .A2(LWORD_REG_0__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n5957) );
  OAI21_X1 U6600 ( .B1(n5958), .B2(n5987), .A(n5957), .ZN(U2923) );
  AOI22_X1 U6601 ( .A1(n6154), .A2(LWORD_REG_1__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n5959) );
  OAI21_X1 U6602 ( .B1(n5960), .B2(n5987), .A(n5959), .ZN(U2922) );
  AOI22_X1 U6603 ( .A1(n6154), .A2(LWORD_REG_2__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n5961) );
  OAI21_X1 U6604 ( .B1(n5962), .B2(n5987), .A(n5961), .ZN(U2921) );
  AOI22_X1 U6605 ( .A1(n6154), .A2(LWORD_REG_3__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n5963) );
  OAI21_X1 U6606 ( .B1(n5964), .B2(n5987), .A(n5963), .ZN(U2920) );
  AOI22_X1 U6607 ( .A1(n6154), .A2(LWORD_REG_4__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n5965) );
  OAI21_X1 U6608 ( .B1(n5966), .B2(n5987), .A(n5965), .ZN(U2919) );
  AOI22_X1 U6609 ( .A1(n6154), .A2(LWORD_REG_5__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n5967) );
  OAI21_X1 U6610 ( .B1(n5968), .B2(n5987), .A(n5967), .ZN(U2918) );
  AOI22_X1 U6611 ( .A1(n6154), .A2(LWORD_REG_6__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n5970) );
  OAI21_X1 U6612 ( .B1(n4727), .B2(n5987), .A(n5970), .ZN(U2917) );
  AOI22_X1 U6613 ( .A1(n6154), .A2(LWORD_REG_7__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n5971) );
  OAI21_X1 U6614 ( .B1(n4730), .B2(n5987), .A(n5971), .ZN(U2916) );
  AOI22_X1 U6615 ( .A1(n6154), .A2(LWORD_REG_8__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n5972) );
  OAI21_X1 U6616 ( .B1(n5973), .B2(n5987), .A(n5972), .ZN(U2915) );
  AOI22_X1 U6617 ( .A1(n6154), .A2(LWORD_REG_9__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n5974) );
  OAI21_X1 U6618 ( .B1(n5975), .B2(n5987), .A(n5974), .ZN(U2914) );
  AOI22_X1 U6619 ( .A1(n6154), .A2(LWORD_REG_10__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n5976) );
  OAI21_X1 U6620 ( .B1(n5977), .B2(n5987), .A(n5976), .ZN(U2913) );
  AOI22_X1 U6621 ( .A1(n6154), .A2(LWORD_REG_11__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n5978) );
  OAI21_X1 U6622 ( .B1(n5979), .B2(n5987), .A(n5978), .ZN(U2912) );
  AOI22_X1 U6623 ( .A1(n6154), .A2(LWORD_REG_12__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n5980) );
  OAI21_X1 U6624 ( .B1(n5981), .B2(n5987), .A(n5980), .ZN(U2911) );
  AOI22_X1 U6625 ( .A1(n6154), .A2(LWORD_REG_13__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n5982) );
  OAI21_X1 U6626 ( .B1(n5983), .B2(n5987), .A(n5982), .ZN(U2910) );
  AOI22_X1 U6627 ( .A1(n6154), .A2(LWORD_REG_14__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n5984) );
  OAI21_X1 U6628 ( .B1(n5985), .B2(n5987), .A(n5984), .ZN(U2909) );
  AOI22_X1 U6629 ( .A1(n6154), .A2(LWORD_REG_15__SCAN_IN), .B1(n5969), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n5986) );
  OAI21_X1 U6630 ( .B1(n5988), .B2(n5987), .A(n5986), .ZN(U2908) );
  AND2_X1 U6631 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6512), .ZN(n6036) );
  INV_X2 U6632 ( .A(n6512), .ZN(n6509) );
  INV_X1 U6633 ( .A(n6038), .ZN(n6028) );
  AOI22_X1 U6634 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6509), .ZN(n5989) );
  OAI21_X1 U6635 ( .B1(n4836), .B2(n6030), .A(n5989), .ZN(U3184) );
  INV_X1 U6636 ( .A(REIP_REG_2__SCAN_IN), .ZN(n5991) );
  AOI22_X1 U6637 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6509), .ZN(n5990) );
  OAI21_X1 U6638 ( .B1(n5991), .B2(n6030), .A(n5990), .ZN(U3185) );
  AOI22_X1 U6639 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6509), .ZN(n5992) );
  OAI21_X1 U6640 ( .B1(n5993), .B2(n6030), .A(n5992), .ZN(U3186) );
  AOI22_X1 U6641 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6509), .ZN(n5994) );
  OAI21_X1 U6642 ( .B1(n6309), .B2(n6030), .A(n5994), .ZN(U3187) );
  AOI22_X1 U6643 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6509), .ZN(n5995) );
  OAI21_X1 U6644 ( .B1(n6308), .B2(n6030), .A(n5995), .ZN(U3188) );
  INV_X1 U6645 ( .A(REIP_REG_6__SCAN_IN), .ZN(n5997) );
  AOI22_X1 U6646 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6509), .ZN(n5996) );
  OAI21_X1 U6647 ( .B1(n5997), .B2(n6030), .A(n5996), .ZN(U3189) );
  INV_X1 U6648 ( .A(REIP_REG_7__SCAN_IN), .ZN(n5999) );
  AOI22_X1 U6649 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6509), .ZN(n5998) );
  OAI21_X1 U6650 ( .B1(n5999), .B2(n6030), .A(n5998), .ZN(U3190) );
  AOI22_X1 U6651 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6509), .ZN(n6000) );
  OAI21_X1 U6652 ( .B1(n6001), .B2(n6030), .A(n6000), .ZN(U3191) );
  AOI22_X1 U6653 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6509), .ZN(n6002) );
  OAI21_X1 U6654 ( .B1(n6003), .B2(n6030), .A(n6002), .ZN(U3192) );
  AOI22_X1 U6655 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6509), .ZN(n6004) );
  OAI21_X1 U6656 ( .B1(n6225), .B2(n6030), .A(n6004), .ZN(U3193) );
  AOI22_X1 U6657 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6509), .ZN(n6005) );
  OAI21_X1 U6658 ( .B1(n6255), .B2(n6030), .A(n6005), .ZN(U3194) );
  AOI22_X1 U6659 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6509), .ZN(n6006) );
  OAI21_X1 U6660 ( .B1(n6007), .B2(n6030), .A(n6006), .ZN(U3195) );
  AOI22_X1 U6661 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6509), .ZN(n6008) );
  OAI21_X1 U6662 ( .B1(n6009), .B2(n6030), .A(n6008), .ZN(U3196) );
  AOI22_X1 U6663 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6509), .ZN(n6010) );
  OAI21_X1 U6664 ( .B1(n6011), .B2(n6030), .A(n6010), .ZN(U3197) );
  AOI22_X1 U6665 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6509), .ZN(n6012) );
  OAI21_X1 U6666 ( .B1(n5805), .B2(n6030), .A(n6012), .ZN(U3198) );
  AOI22_X1 U6667 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6036), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6509), .ZN(n6013) );
  OAI21_X1 U6668 ( .B1(n6268), .B2(n6038), .A(n6013), .ZN(U3199) );
  AOI22_X1 U6669 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6509), .ZN(n6014) );
  OAI21_X1 U6670 ( .B1(n6268), .B2(n6030), .A(n6014), .ZN(U3200) );
  AOI22_X1 U6671 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6509), .ZN(n6015) );
  OAI21_X1 U6672 ( .B1(n6016), .B2(n6030), .A(n6015), .ZN(U3201) );
  AOI22_X1 U6673 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6509), .ZN(n6017) );
  OAI21_X1 U6674 ( .B1(n6157), .B2(n6030), .A(n6017), .ZN(U3202) );
  AOI22_X1 U6675 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6509), .ZN(n6018) );
  OAI21_X1 U6676 ( .B1(n6374), .B2(n6030), .A(n6018), .ZN(U3203) );
  AOI22_X1 U6677 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6036), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6509), .ZN(n6019) );
  OAI21_X1 U6678 ( .B1(n6402), .B2(n6038), .A(n6019), .ZN(U3204) );
  AOI22_X1 U6679 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6509), .ZN(n6020) );
  OAI21_X1 U6680 ( .B1(n6402), .B2(n6030), .A(n6020), .ZN(U3205) );
  AOI22_X1 U6681 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6036), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6509), .ZN(n6021) );
  OAI21_X1 U6682 ( .B1(n6023), .B2(n6038), .A(n6021), .ZN(U3206) );
  AOI22_X1 U6683 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6509), .ZN(n6022) );
  OAI21_X1 U6684 ( .B1(n6023), .B2(n6030), .A(n6022), .ZN(U3207) );
  AOI22_X1 U6685 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6509), .ZN(n6024) );
  OAI21_X1 U6686 ( .B1(n6025), .B2(n6030), .A(n6024), .ZN(U3208) );
  AOI22_X1 U6687 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6509), .ZN(n6026) );
  OAI21_X1 U6688 ( .B1(n6027), .B2(n6030), .A(n6026), .ZN(U3209) );
  AOI22_X1 U6689 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6028), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6509), .ZN(n6029) );
  OAI21_X1 U6690 ( .B1(n6031), .B2(n6030), .A(n6029), .ZN(U3210) );
  AOI22_X1 U6691 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6036), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6509), .ZN(n6032) );
  OAI21_X1 U6692 ( .B1(n6033), .B2(n6038), .A(n6032), .ZN(U3211) );
  AOI22_X1 U6693 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6036), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6509), .ZN(n6034) );
  OAI21_X1 U6694 ( .B1(n6035), .B2(n6038), .A(n6034), .ZN(U3212) );
  AOI22_X1 U6695 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6036), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6509), .ZN(n6037) );
  OAI21_X1 U6696 ( .B1(n6039), .B2(n6038), .A(n6037), .ZN(U3213) );
  MUX2_X1 U6697 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6512), .Z(U3445) );
  AOI221_X1 U6698 ( .B1(REIP_REG_0__SCAN_IN), .B2(REIP_REG_1__SCAN_IN), .C1(
        DATAWIDTH_REG_0__SCAN_IN), .C2(REIP_REG_1__SCAN_IN), .A(
        DATAWIDTH_REG_1__SCAN_IN), .ZN(n6050) );
  NOR4_X1 U6699 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(
        DATAWIDTH_REG_10__SCAN_IN), .ZN(n6043) );
  NOR4_X1 U6700 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n6042) );
  NOR4_X1 U6701 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_2__SCAN_IN), .ZN(
        n6041) );
  NOR4_X1 U6702 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(
        n6040) );
  NAND4_X1 U6703 ( .A1(n6043), .A2(n6042), .A3(n6041), .A4(n6040), .ZN(n6049)
         );
  NOR4_X1 U6704 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_27__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n6047) );
  AOI211_X1 U6705 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_31__SCAN_IN), .B(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6046) );
  NOR4_X1 U6706 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n6045) );
  NOR4_X1 U6707 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_23__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n6044) );
  NAND4_X1 U6708 ( .A1(n6047), .A2(n6046), .A3(n6045), .A4(n6044), .ZN(n6048)
         );
  NOR2_X1 U6709 ( .A1(n6049), .A2(n6048), .ZN(n6059) );
  MUX2_X1 U6710 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(n6050), .S(n6059), .Z(
        U2795) );
  MUX2_X1 U6711 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6512), .Z(U3446) );
  AOI21_X1 U6712 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6051) );
  OAI221_X1 U6713 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6051), .C1(n4836), .C2(
        REIP_REG_0__SCAN_IN), .A(n6059), .ZN(n6052) );
  OAI21_X1 U6714 ( .B1(n6059), .B2(n6053), .A(n6052), .ZN(U3468) );
  MUX2_X1 U6715 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6512), .Z(U3447) );
  NOR3_X1 U6716 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6054) );
  OAI21_X1 U6717 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6054), .A(n6059), .ZN(n6055)
         );
  OAI21_X1 U6718 ( .B1(n6059), .B2(n6056), .A(n6055), .ZN(U2794) );
  MUX2_X1 U6719 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6512), .Z(U3448) );
  OAI21_X1 U6720 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6059), .ZN(n6057) );
  OAI21_X1 U6721 ( .B1(n6059), .B2(n6058), .A(n6057), .ZN(U3469) );
  OAI22_X1 U6722 ( .A1(n6526), .A2(n6061), .B1(n6060), .B2(n6389), .ZN(n6062)
         );
  INV_X1 U6723 ( .A(n6062), .ZN(n6063) );
  OAI21_X1 U6724 ( .B1(n6075), .B2(n6064), .A(n6063), .ZN(U2838) );
  INV_X1 U6725 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U6726 ( .A1(n6066), .A2(n6065), .ZN(n6067) );
  AND2_X1 U6727 ( .A1(n5427), .A2(n6067), .ZN(n6523) );
  AOI21_X1 U6728 ( .B1(n6070), .B2(n6069), .A(n6068), .ZN(n6362) );
  AOI22_X1 U6729 ( .A1(n6523), .A2(n6072), .B1(n6071), .B2(n6362), .ZN(n6073)
         );
  OAI21_X1 U6730 ( .B1(n6075), .B2(n6074), .A(n6073), .ZN(U2840) );
  NAND2_X1 U6731 ( .A1(n6076), .A2(n6101), .ZN(n6078) );
  AOI22_X1 U6732 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n6078), .B1(n5804), 
        .B2(n6077), .ZN(n6080) );
  NAND2_X1 U6733 ( .A1(n6277), .A2(REIP_REG_0__SCAN_IN), .ZN(n6079) );
  OAI211_X1 U6734 ( .C1(n6424), .C2(n6081), .A(n6080), .B(n6079), .ZN(U2986)
         );
  NOR2_X1 U6735 ( .A1(n6269), .A2(n4836), .ZN(n6084) );
  OAI22_X1 U6736 ( .A1(n6122), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n7005), 
        .B2(n6082), .ZN(n6083) );
  AOI211_X1 U6737 ( .C1(n6123), .C2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n6084), 
        .B(n6083), .ZN(n6085) );
  OAI21_X1 U6738 ( .B1(n6424), .B2(n6086), .A(n6085), .ZN(U2985) );
  AOI22_X1 U6739 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6123), .B1(n6277), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U6740 ( .A1(n6089), .A2(n6088), .ZN(n6090) );
  XNOR2_X1 U6741 ( .A(n6087), .B(n6090), .ZN(n6187) );
  OAI22_X1 U6742 ( .A1(n6187), .A2(n6424), .B1(n7005), .B2(n6091), .ZN(n6092)
         );
  INV_X1 U6743 ( .A(n6092), .ZN(n6093) );
  OAI211_X1 U6744 ( .C1(n6122), .C2(n6095), .A(n6094), .B(n6093), .ZN(U2984)
         );
  OAI222_X1 U6745 ( .A1(n6122), .A2(n6321), .B1(n6096), .B2(n6424), .C1(n7005), 
        .C2(n6317), .ZN(n6097) );
  INV_X1 U6746 ( .A(n6097), .ZN(n6099) );
  OAI211_X1 U6747 ( .C1(n6101), .C2(n6100), .A(n6099), .B(n6098), .ZN(U2981)
         );
  AOI22_X1 U6748 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6123), .B1(n6277), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n6105) );
  OAI22_X1 U6749 ( .A1(n6102), .A2(n6424), .B1(n6326), .B2(n7005), .ZN(n6103)
         );
  INV_X1 U6750 ( .A(n6103), .ZN(n6104) );
  OAI211_X1 U6751 ( .C1(n6122), .C2(n6332), .A(n6105), .B(n6104), .ZN(U2980)
         );
  AOI22_X1 U6752 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n6123), .B1(n6277), 
        .B2(REIP_REG_7__SCAN_IN), .ZN(n6112) );
  OR2_X1 U6753 ( .A1(n6107), .A2(n6106), .ZN(n6108) );
  NAND2_X1 U6754 ( .A1(n6109), .A2(n6108), .ZN(n6211) );
  INV_X1 U6755 ( .A(n6211), .ZN(n6110) );
  AOI22_X1 U6756 ( .A1(n6110), .A2(n6128), .B1(n5804), .B2(n6333), .ZN(n6111)
         );
  OAI211_X1 U6757 ( .C1(n6122), .C2(n6346), .A(n6112), .B(n6111), .ZN(U2979)
         );
  AOI22_X1 U6758 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n6123), .B1(n6277), 
        .B2(REIP_REG_17__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U6759 ( .A1(n6113), .A2(n6115), .ZN(n6116) );
  MUX2_X1 U6760 ( .A(n6116), .B(n6115), .S(n6114), .Z(n6118) );
  NAND2_X1 U6761 ( .A1(n6118), .A2(n6117), .ZN(n6267) );
  AOI22_X1 U6762 ( .A1(n6267), .A2(n6128), .B1(n5804), .B2(n6513), .ZN(n6119)
         );
  OAI211_X1 U6763 ( .C1(n6122), .C2(n6121), .A(n6120), .B(n6119), .ZN(U2969)
         );
  AOI22_X1 U6764 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n6123), .B1(n6277), 
        .B2(REIP_REG_19__SCAN_IN), .ZN(n6130) );
  INV_X1 U6765 ( .A(n6125), .ZN(n6127) );
  OAI21_X1 U6766 ( .B1(n3447), .B2(n6127), .A(n6126), .ZN(n6161) );
  AOI22_X1 U6767 ( .A1(n6161), .A2(n6128), .B1(n5804), .B2(n6523), .ZN(n6129)
         );
  OAI211_X1 U6768 ( .C1(n6122), .C2(n6357), .A(n6130), .B(n6129), .ZN(U2967)
         );
  AND2_X1 U6769 ( .A1(n6131), .A2(n6461), .ZN(n6133) );
  OAI22_X1 U6770 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6134), .B1(n6133), .B2(
        n6132), .ZN(U2790) );
  NOR2_X1 U6771 ( .A1(n6512), .A2(D_C_N_REG_SCAN_IN), .ZN(n6135) );
  AOI22_X1 U6772 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n6512), .B1(n6136), .B2(
        n6135), .ZN(U2791) );
  AOI221_X1 U6773 ( .B1(n6152), .B2(n6139), .C1(READREQUEST_REG_SCAN_IN), .C2(
        n6138), .A(n6137), .ZN(n6140) );
  INV_X1 U6774 ( .A(n6140), .ZN(U3474) );
  AOI22_X1 U6775 ( .A1(n6512), .A2(READREQUEST_REG_SCAN_IN), .B1(n6141), .B2(
        n6509), .ZN(U3470) );
  NOR2_X1 U6776 ( .A1(n6142), .A2(n6493), .ZN(n6492) );
  NOR2_X1 U6777 ( .A1(n6501), .A2(n6495), .ZN(n6504) );
  AOI21_X1 U6778 ( .B1(HOLD), .B2(STATE_REG_1__SCAN_IN), .A(n6504), .ZN(n6144)
         );
  NAND2_X1 U6779 ( .A1(STATE_REG_1__SCAN_IN), .A2(READY_N), .ZN(n6505) );
  OAI211_X1 U6780 ( .C1(n6492), .C2(n6144), .A(n6143), .B(n6505), .ZN(U3182)
         );
  NOR2_X1 U6781 ( .A1(READY_N), .A2(n6482), .ZN(n6145) );
  AOI21_X1 U6782 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n6145), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n6147) );
  OAI21_X1 U6783 ( .B1(n6148), .B2(n6147), .A(n6146), .ZN(U3150) );
  AOI211_X1 U6784 ( .C1(n3818), .C2(n6736), .A(n6720), .B(n6149), .ZN(n6151)
         );
  INV_X1 U6785 ( .A(n6150), .ZN(n6479) );
  OAI21_X1 U6786 ( .B1(n6151), .B2(n6482), .A(n6479), .ZN(n6156) );
  AOI211_X1 U6787 ( .C1(n6154), .C2(n6500), .A(n6153), .B(n6152), .ZN(n6155)
         );
  MUX2_X1 U6788 ( .A(n6156), .B(REQUESTPENDING_REG_SCAN_IN), .S(n6155), .Z(
        U3472) );
  OAI22_X1 U6789 ( .A1(n6159), .A2(n6158), .B1(n6269), .B2(n6157), .ZN(n6160)
         );
  INV_X1 U6790 ( .A(n6160), .ZN(n6163) );
  AOI22_X1 U6791 ( .A1(n6161), .A2(n6281), .B1(n6280), .B2(n6362), .ZN(n6162)
         );
  OAI211_X1 U6792 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n6164), .A(n6163), .B(n6162), .ZN(U2999) );
  AOI21_X1 U6793 ( .B1(n6165), .B2(n6174), .A(n6252), .ZN(n6178) );
  INV_X1 U6794 ( .A(n6166), .ZN(n6167) );
  AOI21_X1 U6795 ( .B1(n6280), .B2(n6168), .A(n6167), .ZN(n6172) );
  NOR4_X1 U6796 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6249), .A3(n4099), 
        .A4(n6250), .ZN(n6169) );
  AOI21_X1 U6797 ( .B1(n6170), .B2(n6281), .A(n6169), .ZN(n6171) );
  OAI211_X1 U6798 ( .C1(n6178), .C2(n6173), .A(n6172), .B(n6171), .ZN(U3005)
         );
  OR2_X1 U6799 ( .A1(n6249), .A2(n6174), .ZN(n6180) );
  AOI222_X1 U6800 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6277), .B1(n6280), .B2(
        n6176), .C1(n6281), .C2(n6175), .ZN(n6177) );
  OAI221_X1 U6801 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n6180), .C1(
        n6179), .C2(n6178), .A(n6177), .ZN(U3004) );
  NAND2_X1 U6802 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6181), .ZN(n6194)
         );
  NAND2_X1 U6803 ( .A1(n6280), .A2(n6182), .ZN(n6191) );
  NAND2_X1 U6804 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6184) );
  OAI21_X1 U6805 ( .B1(n6184), .B2(n3700), .A(n6183), .ZN(n6185) );
  INV_X1 U6806 ( .A(n6185), .ZN(n6186) );
  OR2_X1 U6807 ( .A1(n6217), .A2(n6186), .ZN(n6190) );
  OR2_X1 U6808 ( .A1(n6223), .A2(n6187), .ZN(n6189) );
  NAND2_X1 U6809 ( .A1(n6277), .A2(REIP_REG_2__SCAN_IN), .ZN(n6188) );
  AND4_X1 U6810 ( .A1(n6191), .A2(n6190), .A3(n6189), .A4(n6188), .ZN(n6192)
         );
  OAI221_X1 U6811 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6194), .C1(n3700), .C2(n6193), .A(n6192), .ZN(U3016) );
  INV_X1 U6812 ( .A(n6195), .ZN(n6201) );
  OAI21_X1 U6813 ( .B1(n6201), .B2(n6217), .A(n6196), .ZN(n6197) );
  AOI21_X1 U6814 ( .B1(n6199), .B2(n6198), .A(n6197), .ZN(n6216) );
  NAND2_X1 U6815 ( .A1(n6201), .A2(n6200), .ZN(n6231) );
  INV_X1 U6816 ( .A(n6231), .ZN(n6202) );
  OAI211_X1 U6817 ( .C1(INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6232), .B(n6202), .ZN(n6205) );
  AOI22_X1 U6818 ( .A1(n6280), .A2(n6203), .B1(n6277), .B2(REIP_REG_8__SCAN_IN), .ZN(n6204) );
  OAI211_X1 U6819 ( .C1(n6206), .C2(n6223), .A(n6205), .B(n6204), .ZN(n6207)
         );
  INV_X1 U6820 ( .A(n6207), .ZN(n6208) );
  OAI21_X1 U6821 ( .B1(n6216), .B2(n6209), .A(n6208), .ZN(U3010) );
  INV_X1 U6822 ( .A(n6335), .ZN(n6210) );
  AOI22_X1 U6823 ( .A1(n6280), .A2(n6210), .B1(n6277), .B2(REIP_REG_7__SCAN_IN), .ZN(n6214) );
  OAI22_X1 U6824 ( .A1(n6231), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .B1(n6211), 
        .B2(n6223), .ZN(n6212) );
  INV_X1 U6825 ( .A(n6212), .ZN(n6213) );
  OAI211_X1 U6826 ( .C1(n6216), .C2(n6215), .A(n6214), .B(n6213), .ZN(U3011)
         );
  OAI22_X1 U6827 ( .A1(n6220), .A2(n6219), .B1(n6218), .B2(n6217), .ZN(n6221)
         );
  NOR2_X1 U6828 ( .A1(n6222), .A2(n6221), .ZN(n6245) );
  NOR2_X1 U6829 ( .A1(n6224), .A2(n6223), .ZN(n6230) );
  OAI22_X1 U6830 ( .A1(n6227), .A2(n6226), .B1(n6225), .B2(n6269), .ZN(n6228)
         );
  AOI21_X1 U6831 ( .B1(n6230), .B2(n6229), .A(n6228), .ZN(n6235) );
  NOR2_X1 U6832 ( .A1(n6232), .A2(n6231), .ZN(n6241) );
  NAND2_X1 U6833 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6233) );
  OAI211_X1 U6834 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A(n6241), .B(n6233), .ZN(n6234) );
  OAI211_X1 U6835 ( .C1(n6245), .C2(n4100), .A(n6235), .B(n6234), .ZN(U3008)
         );
  INV_X1 U6836 ( .A(n6236), .ZN(n6237) );
  AOI21_X1 U6837 ( .B1(n6280), .B2(n6238), .A(n6237), .ZN(n6243) );
  INV_X1 U6838 ( .A(n6239), .ZN(n6240) );
  AOI22_X1 U6839 ( .A1(n6241), .A2(n6244), .B1(n6240), .B2(n6281), .ZN(n6242)
         );
  OAI211_X1 U6840 ( .C1(n6245), .C2(n6244), .A(n6243), .B(n6242), .ZN(U3009)
         );
  INV_X1 U6841 ( .A(n6246), .ZN(n6248) );
  AOI22_X1 U6842 ( .A1(n6248), .A2(n6281), .B1(n6280), .B2(n6247), .ZN(n6254)
         );
  INV_X1 U6843 ( .A(n6249), .ZN(n6251) );
  AOI22_X1 U6844 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6252), .B1(n6251), .B2(n6250), .ZN(n6253) );
  OAI211_X1 U6845 ( .C1(n6255), .C2(n6269), .A(n6254), .B(n6253), .ZN(U3007)
         );
  AOI21_X1 U6846 ( .B1(n6280), .B2(n6257), .A(n6256), .ZN(n6265) );
  AOI22_X1 U6847 ( .A1(n6259), .A2(n6281), .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n6258), .ZN(n6264) );
  OAI221_X1 U6848 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .C1(n6262), .C2(n6261), .A(n6260), 
        .ZN(n6263) );
  NAND3_X1 U6849 ( .A1(n6265), .A2(n6264), .A3(n6263), .ZN(U3002) );
  AOI22_X1 U6850 ( .A1(n6267), .A2(n6281), .B1(n6280), .B2(n6266), .ZN(n6275)
         );
  NOR2_X1 U6851 ( .A1(n6269), .A2(n6268), .ZN(n6270) );
  AOI221_X1 U6852 ( .B1(n6273), .B2(n6272), .C1(n6271), .C2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A(n6270), .ZN(n6274) );
  NAND2_X1 U6853 ( .A1(n6275), .A2(n6274), .ZN(U3001) );
  AOI22_X1 U6854 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6277), .B1(n6276), .B2(
        n6285), .ZN(n6284) );
  INV_X1 U6855 ( .A(n6278), .ZN(n6282) );
  AOI22_X1 U6856 ( .A1(n6282), .A2(n6281), .B1(n6280), .B2(n6279), .ZN(n6283)
         );
  OAI211_X1 U6857 ( .C1(n6286), .C2(n6285), .A(n6284), .B(n6283), .ZN(U2993)
         );
  INV_X1 U6858 ( .A(n6287), .ZN(n6288) );
  AOI22_X1 U6859 ( .A1(REIP_REG_0__SCAN_IN), .A2(n6304), .B1(n6418), .B2(n6288), .ZN(n6291) );
  NAND2_X1 U6860 ( .A1(n6412), .A2(n6410), .ZN(n6289) );
  AOI222_X1 U6861 ( .A1(n6289), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .B1(n6294), 
        .B2(n4153), .C1(EBX_REG_0__SCAN_IN), .C2(n6415), .ZN(n6290) );
  OAI211_X1 U6862 ( .C1(n6318), .C2(n6292), .A(n6291), .B(n6290), .ZN(U2827)
         );
  AOI22_X1 U6863 ( .A1(n6418), .A2(n6293), .B1(n6395), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6307) );
  INV_X1 U6864 ( .A(n6426), .ZN(n6298) );
  INV_X1 U6865 ( .A(n6294), .ZN(n6297) );
  NAND2_X1 U6866 ( .A1(n6296), .A2(n6295), .ZN(n6310) );
  OAI22_X1 U6867 ( .A1(n6298), .A2(n6297), .B1(n6310), .B2(REIP_REG_4__SCAN_IN), .ZN(n6302) );
  OAI22_X1 U6868 ( .A1(n6318), .A2(n6300), .B1(n6299), .B2(n6410), .ZN(n6301)
         );
  AOI211_X1 U6869 ( .C1(EBX_REG_4__SCAN_IN), .C2(n6415), .A(n6302), .B(n6301), 
        .ZN(n6306) );
  NAND3_X1 U6870 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6304), .A3(n6303), .ZN(n6305) );
  NAND4_X1 U6871 ( .A1(n6307), .A2(n6306), .A3(n6348), .A4(n6305), .ZN(U2823)
         );
  OAI21_X1 U6872 ( .B1(n6310), .B2(n6309), .A(n6308), .ZN(n6311) );
  NAND2_X1 U6873 ( .A1(n6311), .A2(n6337), .ZN(n6316) );
  NAND2_X1 U6874 ( .A1(n6395), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6312)
         );
  OAI211_X1 U6875 ( .C1(n6390), .C2(n6313), .A(n6348), .B(n6312), .ZN(n6314)
         );
  AOI21_X1 U6876 ( .B1(n6415), .B2(EBX_REG_5__SCAN_IN), .A(n6314), .ZN(n6315)
         );
  OAI211_X1 U6877 ( .C1(n6318), .C2(n6317), .A(n6316), .B(n6315), .ZN(n6319)
         );
  INV_X1 U6878 ( .A(n6319), .ZN(n6320) );
  OAI21_X1 U6879 ( .B1(n6321), .B2(n6410), .A(n6320), .ZN(U2822) );
  OR2_X1 U6880 ( .A1(n6340), .A2(REIP_REG_6__SCAN_IN), .ZN(n6330) );
  NAND2_X1 U6881 ( .A1(n6337), .A2(REIP_REG_6__SCAN_IN), .ZN(n6329) );
  INV_X1 U6882 ( .A(n6322), .ZN(n6323) );
  OAI22_X1 U6883 ( .A1(n6324), .A2(n6383), .B1(n6323), .B2(n6390), .ZN(n6325)
         );
  AOI211_X1 U6884 ( .C1(n6395), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6360), 
        .B(n6325), .ZN(n6328) );
  OR2_X1 U6885 ( .A1(n6326), .A2(n6391), .ZN(n6327) );
  AND4_X1 U6886 ( .A1(n6330), .A2(n6329), .A3(n6328), .A4(n6327), .ZN(n6331)
         );
  OAI21_X1 U6887 ( .B1(n6332), .B2(n6410), .A(n6331), .ZN(U2821) );
  NAND2_X1 U6888 ( .A1(n6333), .A2(n6419), .ZN(n6344) );
  NAND2_X1 U6889 ( .A1(n6395), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6334)
         );
  OAI211_X1 U6890 ( .C1(n6390), .C2(n6335), .A(n6348), .B(n6334), .ZN(n6336)
         );
  AOI21_X1 U6891 ( .B1(n6415), .B2(EBX_REG_7__SCAN_IN), .A(n6336), .ZN(n6343)
         );
  NAND2_X1 U6892 ( .A1(n6337), .A2(REIP_REG_7__SCAN_IN), .ZN(n6342) );
  OAI21_X1 U6893 ( .B1(REIP_REG_6__SCAN_IN), .B2(REIP_REG_7__SCAN_IN), .A(
        n6338), .ZN(n6339) );
  OR2_X1 U6894 ( .A1(n6340), .A2(n6339), .ZN(n6341) );
  AND4_X1 U6895 ( .A1(n6344), .A2(n6343), .A3(n6342), .A4(n6341), .ZN(n6345)
         );
  OAI21_X1 U6896 ( .B1(n6346), .B2(n6410), .A(n6345), .ZN(U2820) );
  AOI22_X1 U6897 ( .A1(n6415), .A2(EBX_REG_15__SCAN_IN), .B1(n6418), .B2(n6347), .ZN(n6349) );
  OAI211_X1 U6898 ( .C1(n6412), .C2(n6350), .A(n6349), .B(n6348), .ZN(n6351)
         );
  AOI21_X1 U6899 ( .B1(REIP_REG_15__SCAN_IN), .B2(n6352), .A(n6351), .ZN(n6356) );
  AOI22_X1 U6900 ( .A1(n6354), .A2(n6419), .B1(n6397), .B2(n6353), .ZN(n6355)
         );
  OAI211_X1 U6901 ( .C1(REIP_REG_15__SCAN_IN), .C2(n6375), .A(n6356), .B(n6355), .ZN(U2812) );
  INV_X1 U6902 ( .A(n6357), .ZN(n6358) );
  AOI22_X1 U6903 ( .A1(n6358), .A2(n6397), .B1(EBX_REG_19__SCAN_IN), .B2(n6415), .ZN(n6368) );
  NOR3_X1 U6904 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6359), .A3(n6375), .ZN(n6361) );
  AOI211_X1 U6905 ( .C1(n6395), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6361), 
        .B(n6360), .ZN(n6367) );
  AOI22_X1 U6906 ( .A1(n6523), .A2(n6419), .B1(n6418), .B2(n6362), .ZN(n6366)
         );
  OAI21_X1 U6907 ( .B1(n6364), .B2(n6363), .A(REIP_REG_19__SCAN_IN), .ZN(n6365) );
  NAND4_X1 U6908 ( .A1(n6368), .A2(n6367), .A3(n6366), .A4(n6365), .ZN(U2808)
         );
  AOI22_X1 U6909 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n6395), .B1(n6369), 
        .B2(n6397), .ZN(n6382) );
  AOI21_X1 U6910 ( .B1(n6372), .B2(n6371), .A(n6370), .ZN(n6396) );
  INV_X1 U6911 ( .A(n6373), .ZN(n6376) );
  OAI21_X1 U6912 ( .B1(n6376), .B2(n6375), .A(n6374), .ZN(n6380) );
  OAI22_X1 U6913 ( .A1(n6378), .A2(n6391), .B1(n6377), .B2(n6390), .ZN(n6379)
         );
  AOI21_X1 U6914 ( .B1(n6396), .B2(n6380), .A(n6379), .ZN(n6381) );
  OAI211_X1 U6915 ( .C1(n3771), .C2(n6383), .A(n6382), .B(n6381), .ZN(U2807)
         );
  NOR2_X1 U6916 ( .A1(n6385), .A2(n6384), .ZN(n6408) );
  AOI22_X1 U6917 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n6395), .B1(
        EBX_REG_21__SCAN_IN), .B2(n6415), .ZN(n6386) );
  OAI21_X1 U6918 ( .B1(n6387), .B2(n6410), .A(n6386), .ZN(n6388) );
  AOI221_X1 U6919 ( .B1(n6396), .B2(REIP_REG_21__SCAN_IN), .C1(n6408), .C2(
        n6401), .A(n6388), .ZN(n6394) );
  OAI22_X1 U6920 ( .A1(n6526), .A2(n6391), .B1(n6390), .B2(n6389), .ZN(n6392)
         );
  INV_X1 U6921 ( .A(n6392), .ZN(n6393) );
  NAND2_X1 U6922 ( .A1(n6394), .A2(n6393), .ZN(U2806) );
  AOI22_X1 U6923 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n6395), .B1(
        EBX_REG_22__SCAN_IN), .B2(n6415), .ZN(n6407) );
  AOI22_X1 U6924 ( .A1(n6398), .A2(n6397), .B1(REIP_REG_22__SCAN_IN), .B2(
        n6396), .ZN(n6406) );
  INV_X1 U6925 ( .A(n6399), .ZN(n6530) );
  AOI22_X1 U6926 ( .A1(n6530), .A2(n6419), .B1(n6400), .B2(n6418), .ZN(n6405)
         );
  NOR2_X1 U6927 ( .A1(n6402), .A2(n6401), .ZN(n6409) );
  INV_X1 U6928 ( .A(n6409), .ZN(n6403) );
  OAI211_X1 U6929 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n6408), .B(n6403), .ZN(n6404) );
  NAND4_X1 U6930 ( .A1(n6407), .A2(n6406), .A3(n6405), .A4(n6404), .ZN(U2805)
         );
  AOI21_X1 U6931 ( .B1(n6409), .B2(n6408), .A(REIP_REG_23__SCAN_IN), .ZN(n6422) );
  INV_X1 U6932 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6413) );
  OAI22_X1 U6933 ( .A1(n6413), .A2(n6412), .B1(n6411), .B2(n6410), .ZN(n6414)
         );
  AOI21_X1 U6934 ( .B1(EBX_REG_23__SCAN_IN), .B2(n6415), .A(n6414), .ZN(n6421)
         );
  INV_X1 U6935 ( .A(n6416), .ZN(n6417) );
  AOI22_X1 U6936 ( .A1(n6535), .A2(n6419), .B1(n6418), .B2(n6417), .ZN(n6420)
         );
  OAI211_X1 U6937 ( .C1(n6423), .C2(n6422), .A(n6421), .B(n6420), .ZN(U2804)
         );
  OAI21_X1 U6938 ( .B1(n6425), .B2(n6451), .A(n6424), .ZN(U2793) );
  INV_X1 U6939 ( .A(n4135), .ZN(n6427) );
  NAND4_X1 U6940 ( .A1(n6428), .A2(n6427), .A3(n6469), .A4(n6426), .ZN(n6429)
         );
  OAI21_X1 U6941 ( .B1(n6430), .B2(n4694), .A(n6429), .ZN(U3455) );
  INV_X1 U6942 ( .A(n6431), .ZN(n6433) );
  NOR3_X1 U6943 ( .A1(n6433), .A2(n6432), .A3(n6709), .ZN(n6434) );
  NAND2_X1 U6944 ( .A1(n6434), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6438) );
  OAI22_X1 U6945 ( .A1(n6436), .A2(n6435), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6434), .ZN(n6437) );
  NAND2_X1 U6946 ( .A1(n6438), .A2(n6437), .ZN(n6441) );
  INV_X1 U6947 ( .A(n6439), .ZN(n6440) );
  AOI21_X1 U6948 ( .B1(n6441), .B2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(n6440), 
        .ZN(n6443) );
  NOR2_X1 U6949 ( .A1(n6441), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6442)
         );
  OAI22_X1 U6950 ( .A1(n6443), .A2(n6442), .B1(n3500), .B2(n6444), .ZN(n6446)
         );
  NAND2_X1 U6951 ( .A1(n6444), .A2(n3500), .ZN(n6445) );
  NAND2_X1 U6952 ( .A1(n6446), .A2(n6445), .ZN(n6460) );
  INV_X1 U6953 ( .A(n6447), .ZN(n6457) );
  NOR2_X1 U6954 ( .A1(n6449), .A2(n6448), .ZN(n6455) );
  NAND2_X1 U6955 ( .A1(n6451), .A2(n6450), .ZN(n6452) );
  NAND2_X1 U6956 ( .A1(n6453), .A2(n6452), .ZN(n6454) );
  NAND4_X1 U6957 ( .A1(n6457), .A2(n6456), .A3(n6455), .A4(n6454), .ZN(n6458)
         );
  AOI21_X1 U6958 ( .B1(n6460), .B2(n6459), .A(n6458), .ZN(n6488) );
  NAND2_X1 U6959 ( .A1(n6488), .A2(n6461), .ZN(n6463) );
  NAND2_X1 U6960 ( .A1(READY_N), .A2(n6154), .ZN(n6462) );
  NAND2_X1 U6961 ( .A1(n6463), .A2(n6462), .ZN(n6467) );
  NAND2_X1 U6962 ( .A1(n6465), .A2(n6464), .ZN(n6466) );
  OAI221_X1 U6963 ( .B1(n6468), .B2(READY_N), .C1(n6468), .C2(n6720), .A(
        STATE2_REG_0__SCAN_IN), .ZN(n6480) );
  NAND3_X1 U6964 ( .A1(n6469), .A2(STATE2_REG_0__SCAN_IN), .A3(n6500), .ZN(
        n6470) );
  NAND3_X1 U6965 ( .A1(n6470), .A2(n6487), .A3(n6477), .ZN(n6471) );
  OAI21_X1 U6966 ( .B1(n6472), .B2(n6477), .A(n6471), .ZN(n6474) );
  OAI211_X1 U6967 ( .C1(n6475), .C2(n6480), .A(n6474), .B(n6473), .ZN(U3149)
         );
  OAI221_X1 U6968 ( .B1(n6744), .B2(STATE2_REG_0__SCAN_IN), .C1(n6744), .C2(
        n6477), .A(n6476), .ZN(U3453) );
  OAI21_X1 U6969 ( .B1(n6479), .B2(n6478), .A(n6477), .ZN(n6481) );
  OAI221_X1 U6970 ( .B1(n6483), .B2(n6482), .C1(n6481), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6480), .ZN(n6484) );
  INV_X1 U6971 ( .A(n6484), .ZN(n6486) );
  OAI211_X1 U6972 ( .C1(n6488), .C2(n6487), .A(n6486), .B(n6485), .ZN(U3148)
         );
  AOI21_X1 U6973 ( .B1(n5952), .B2(STATEBS16_REG_SCAN_IN), .A(n6490), .ZN(
        n6489) );
  INV_X1 U6974 ( .A(n6489), .ZN(U2792) );
  AOI21_X1 U6975 ( .B1(n5952), .B2(DATAWIDTH_REG_1__SCAN_IN), .A(n6490), .ZN(
        n6491) );
  INV_X1 U6976 ( .A(n6491), .ZN(U3452) );
  INV_X1 U6977 ( .A(n6492), .ZN(n6498) );
  INV_X1 U6978 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6494) );
  NOR2_X1 U6979 ( .A1(n6494), .A2(n6493), .ZN(n6496) );
  AOI221_X1 U6980 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6503), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6507) );
  AOI221_X1 U6981 ( .B1(n6496), .B2(n6509), .C1(n6495), .C2(n6509), .A(n6507), 
        .ZN(n6497) );
  OAI221_X1 U6982 ( .B1(n6499), .B2(n6505), .C1(n6499), .C2(n6498), .A(n6497), 
        .ZN(U3181) );
  AOI221_X1 U6983 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6500), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6502) );
  AOI221_X1 U6984 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6502), .C2(HOLD), .A(n6501), .ZN(n6508) );
  AOI21_X1 U6985 ( .B1(n6504), .B2(n6503), .A(STATE_REG_2__SCAN_IN), .ZN(n6506) );
  OAI22_X1 U6986 ( .A1(n6508), .A2(n6507), .B1(n6506), .B2(n6505), .ZN(U3183)
         );
  AOI22_X1 U6987 ( .A1(n6512), .A2(n6511), .B1(n6510), .B2(n6509), .ZN(U3473)
         );
  AOI22_X1 U6988 ( .A1(n6513), .A2(n6534), .B1(n6533), .B2(DATAI_17_), .ZN(
        n6519) );
  OAI22_X1 U6989 ( .A1(n6516), .A2(n5612), .B1(n6515), .B2(n6514), .ZN(n6517)
         );
  INV_X1 U6990 ( .A(n6517), .ZN(n6518) );
  NAND2_X1 U6991 ( .A1(n6519), .A2(n6518), .ZN(U2874) );
  AOI22_X1 U6992 ( .A1(n6520), .A2(n6534), .B1(n6533), .B2(DATAI_18_), .ZN(
        n6522) );
  AOI22_X1 U6993 ( .A1(n6537), .A2(DATAI_2_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n6536), .ZN(n6521) );
  NAND2_X1 U6994 ( .A1(n6522), .A2(n6521), .ZN(U2873) );
  AOI22_X1 U6995 ( .A1(n6523), .A2(n6534), .B1(n6533), .B2(DATAI_19_), .ZN(
        n6525) );
  AOI22_X1 U6996 ( .A1(n6537), .A2(DATAI_3_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n6536), .ZN(n6524) );
  NAND2_X1 U6997 ( .A1(n6525), .A2(n6524), .ZN(U2872) );
  INV_X1 U6998 ( .A(n6526), .ZN(n6527) );
  AOI22_X1 U6999 ( .A1(n6527), .A2(n6534), .B1(n6533), .B2(DATAI_21_), .ZN(
        n6529) );
  AOI22_X1 U7000 ( .A1(n6537), .A2(DATAI_5_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n6536), .ZN(n6528) );
  NAND2_X1 U7001 ( .A1(n6529), .A2(n6528), .ZN(U2870) );
  AOI22_X1 U7002 ( .A1(n6530), .A2(n6534), .B1(n6533), .B2(DATAI_22_), .ZN(
        n6532) );
  AOI22_X1 U7003 ( .A1(n6537), .A2(DATAI_6_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n6536), .ZN(n6531) );
  NAND2_X1 U7004 ( .A1(n6532), .A2(n6531), .ZN(U2869) );
  AOI22_X1 U7005 ( .A1(n6535), .A2(n6534), .B1(n6533), .B2(DATAI_23_), .ZN(
        n6539) );
  AOI22_X1 U7006 ( .A1(n6537), .A2(DATAI_7_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n6536), .ZN(n6538) );
  NAND2_X1 U7007 ( .A1(n6539), .A2(n6538), .ZN(U2868) );
  INV_X1 U7008 ( .A(n6725), .ZN(n6748) );
  NAND3_X1 U7009 ( .A1(n6541), .A2(n6663), .A3(n6566), .ZN(n6552) );
  NAND2_X1 U7010 ( .A1(DATAI_0_), .A2(n6999), .ZN(n6662) );
  AND2_X1 U7011 ( .A1(n4153), .A2(n6630), .ZN(n6608) );
  NOR2_X1 U7012 ( .A1(n4677), .A2(n6607), .ZN(n6631) );
  NOR2_X1 U7013 ( .A1(n6542), .A2(n3500), .ZN(n7002) );
  AOI21_X1 U7014 ( .B1(n6608), .B2(n6631), .A(n7002), .ZN(n6549) );
  NAND3_X1 U7015 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6555) );
  OAI22_X1 U7016 ( .A1(n6549), .A2(n6710), .B1(n6555), .B2(n6720), .ZN(n7003)
         );
  NOR2_X2 U7017 ( .A1(n7001), .A2(n6545), .ZN(n6734) );
  AOI22_X1 U7018 ( .A1(n6735), .A2(n7003), .B1(n6734), .B2(n7002), .ZN(n6554)
         );
  INV_X1 U7019 ( .A(n6552), .ZN(n6547) );
  NAND2_X1 U7020 ( .A1(n6659), .A2(n6736), .ZN(n6699) );
  OAI21_X1 U7021 ( .B1(n6547), .B2(n7005), .A(n6699), .ZN(n6548) );
  AOI22_X1 U7022 ( .A1(n6549), .A2(n6548), .B1(n6710), .B2(n6555), .ZN(n6550)
         );
  NAND2_X1 U7023 ( .A1(n6685), .A2(n6550), .ZN(n7007) );
  NOR2_X1 U7024 ( .A1(n7005), .A2(n6551), .ZN(n6745) );
  AOI22_X1 U7025 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n7007), .B1(n6745), 
        .B2(n7006), .ZN(n6553) );
  OAI211_X1 U7026 ( .C1(n6748), .C2(n7010), .A(n6554), .B(n6553), .ZN(U3140)
         );
  INV_X1 U7027 ( .A(n6745), .ZN(n6728) );
  INV_X1 U7028 ( .A(n6631), .ZN(n6638) );
  NAND2_X1 U7029 ( .A1(n6630), .A2(n6659), .ZN(n6739) );
  NAND2_X1 U7030 ( .A1(n6677), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6556) );
  OR2_X1 U7031 ( .A1(n6557), .A2(n6720), .ZN(n6669) );
  OAI22_X1 U7032 ( .A1(n6638), .A2(n6739), .B1(n6556), .B2(n6669), .ZN(n7012)
         );
  NOR2_X1 U7033 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6555), .ZN(n7011)
         );
  AOI22_X1 U7034 ( .A1(n6735), .A2(n7012), .B1(n6734), .B2(n7011), .ZN(n6565)
         );
  INV_X1 U7035 ( .A(n7011), .ZN(n6558) );
  INV_X1 U7036 ( .A(n6556), .ZN(n6597) );
  NOR2_X1 U7037 ( .A1(n6597), .A2(n6720), .ZN(n6601) );
  NAND2_X1 U7038 ( .A1(n6557), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6730) );
  NAND2_X1 U7039 ( .A1(n6999), .A2(n6730), .ZN(n6674) );
  AOI211_X1 U7040 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6558), .A(n6601), .B(
        n6674), .ZN(n6563) );
  NOR2_X1 U7041 ( .A1(n6630), .A2(n6710), .ZN(n6578) );
  NOR2_X1 U7042 ( .A1(n6631), .A2(n6710), .ZN(n6642) );
  NAND2_X1 U7043 ( .A1(n6566), .A2(n6723), .ZN(n6559) );
  NOR2_X1 U7044 ( .A1(n3436), .A2(n6559), .ZN(n6560) );
  OAI21_X1 U7045 ( .B1(n7013), .B2(n7018), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6561) );
  OAI21_X1 U7046 ( .B1(n6578), .B2(n6642), .A(n6561), .ZN(n6562) );
  NAND2_X1 U7047 ( .A1(n6563), .A2(n6562), .ZN(n7014) );
  AOI22_X1 U7048 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n7014), .B1(n6725), 
        .B2(n7018), .ZN(n6564) );
  OAI211_X1 U7049 ( .C1(n6728), .C2(n7010), .A(n6565), .B(n6564), .ZN(U3132)
         );
  NAND3_X1 U7050 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6717), .ZN(n6577) );
  NOR2_X1 U7051 ( .A1(n6709), .A2(n6577), .ZN(n7019) );
  NAND2_X1 U7052 ( .A1(n6566), .A2(n6696), .ZN(n6567) );
  NOR2_X1 U7053 ( .A1(n3436), .A2(n6567), .ZN(n6568) );
  AOI22_X1 U7054 ( .A1(n6734), .A2(n7019), .B1(n7027), .B2(n6725), .ZN(n6576)
         );
  INV_X1 U7055 ( .A(n6577), .ZN(n6571) );
  NAND2_X1 U7056 ( .A1(n6569), .A2(n6607), .ZN(n6670) );
  INV_X1 U7057 ( .A(n6670), .ZN(n6650) );
  AOI21_X1 U7058 ( .B1(n6608), .B2(n6650), .A(n7019), .ZN(n6574) );
  NAND3_X1 U7059 ( .A1(n6659), .A2(n6574), .A3(n6572), .ZN(n6570) );
  OAI211_X1 U7060 ( .C1(n6659), .C2(n6571), .A(n6685), .B(n6570), .ZN(n7021)
         );
  NAND2_X1 U7061 ( .A1(n6659), .A2(n6572), .ZN(n6573) );
  OAI22_X1 U7062 ( .A1(n6574), .A2(n6573), .B1(n6720), .B2(n6577), .ZN(n7020)
         );
  AOI22_X1 U7063 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n7021), .B1(n6735), 
        .B2(n7020), .ZN(n6575) );
  OAI211_X1 U7064 ( .C1(n6728), .C2(n7017), .A(n6576), .B(n6575), .ZN(U3124)
         );
  INV_X1 U7065 ( .A(n6677), .ZN(n6667) );
  NAND2_X1 U7066 ( .A1(n6667), .A2(n6676), .ZN(n6618) );
  OAI22_X1 U7067 ( .A1(n6739), .A2(n6670), .B1(n6618), .B2(n6669), .ZN(n7026)
         );
  NOR2_X1 U7068 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6577), .ZN(n7025)
         );
  AOI22_X1 U7069 ( .A1(n6735), .A2(n7026), .B1(n6734), .B2(n7025), .ZN(n6584)
         );
  NAND2_X1 U7070 ( .A1(n6670), .A2(n6659), .ZN(n6673) );
  INV_X1 U7071 ( .A(n6579), .ZN(n6664) );
  AND2_X1 U7072 ( .A1(n6666), .A2(n6664), .ZN(n6586) );
  NAND2_X1 U7073 ( .A1(n6586), .A2(n6663), .ZN(n6592) );
  AOI21_X1 U7074 ( .B1(n7031), .B2(n7024), .A(n6736), .ZN(n6580) );
  AOI21_X1 U7075 ( .B1(n6732), .B2(n6673), .A(n6580), .ZN(n6581) );
  NOR2_X1 U7076 ( .A1(n6581), .A2(n6674), .ZN(n6582) );
  NAND2_X1 U7077 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6618), .ZN(n6622) );
  OAI211_X1 U7078 ( .C1(n7025), .C2(n6744), .A(n6582), .B(n6622), .ZN(n7028)
         );
  AOI22_X1 U7079 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n7028), .B1(n6725), 
        .B2(n7033), .ZN(n6583) );
  OAI211_X1 U7080 ( .C1(n6728), .C2(n7024), .A(n6584), .B(n6583), .ZN(U3116)
         );
  AOI21_X1 U7081 ( .B1(n6586), .B2(n6585), .A(n6710), .ZN(n6590) );
  NAND2_X1 U7082 ( .A1(n4677), .A2(n4800), .ZN(n6692) );
  NAND3_X1 U7083 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6649), .ZN(n6599) );
  INV_X1 U7084 ( .A(n6599), .ZN(n6587) );
  AND2_X1 U7085 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6587), .ZN(n7032)
         );
  AOI21_X1 U7086 ( .B1(n6608), .B2(n6697), .A(n7032), .ZN(n6589) );
  INV_X1 U7087 ( .A(n6589), .ZN(n6588) );
  AOI22_X1 U7088 ( .A1(n6590), .A2(n6588), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6587), .ZN(n7037) );
  AOI22_X1 U7089 ( .A1(n6734), .A2(n7032), .B1(n7033), .B2(n6745), .ZN(n6594)
         );
  AOI22_X1 U7090 ( .A1(n6590), .A2(n6589), .B1(n6599), .B2(n6710), .ZN(n6591)
         );
  NAND2_X1 U7091 ( .A1(n6685), .A2(n6591), .ZN(n7034) );
  NOR2_X2 U7092 ( .A1(n6592), .A2(n6723), .ZN(n7039) );
  AOI22_X1 U7093 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n7034), .B1(n7039), 
        .B2(n6725), .ZN(n6593) );
  OAI211_X1 U7094 ( .C1(n7037), .C2(n6662), .A(n6594), .B(n6593), .ZN(U3108)
         );
  INV_X1 U7095 ( .A(n7044), .ZN(n6595) );
  NAND2_X1 U7096 ( .A1(n6595), .A2(n6659), .ZN(n6596) );
  OAI21_X1 U7097 ( .B1(n6596), .B2(n7039), .A(n6699), .ZN(n6603) );
  AND2_X1 U7098 ( .A1(n6697), .A2(n6630), .ZN(n6600) );
  INV_X1 U7099 ( .A(n6730), .ZN(n6598) );
  NOR2_X1 U7100 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6599), .ZN(n7038)
         );
  AOI22_X1 U7101 ( .A1(n6734), .A2(n7038), .B1(n7044), .B2(n6725), .ZN(n6606)
         );
  INV_X1 U7102 ( .A(n6600), .ZN(n6602) );
  NAND2_X1 U7103 ( .A1(n6999), .A2(n6669), .ZN(n6740) );
  AOI211_X1 U7104 ( .C1(n6603), .C2(n6602), .A(n6740), .B(n6601), .ZN(n6604)
         );
  AOI22_X1 U7105 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n7040), .B1(n7039), 
        .B2(n6745), .ZN(n6605) );
  OAI211_X1 U7106 ( .C1(n7043), .C2(n6662), .A(n6606), .B(n6605), .ZN(U3100)
         );
  NOR3_X1 U7107 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n3500), .ZN(n6614) );
  INV_X1 U7108 ( .A(n6614), .ZN(n6619) );
  NAND2_X1 U7109 ( .A1(n4677), .A2(n6607), .ZN(n6731) );
  INV_X1 U7110 ( .A(n6731), .ZN(n6707) );
  NOR2_X1 U7111 ( .A1(n6709), .A2(n6619), .ZN(n7045) );
  AOI21_X1 U7112 ( .B1(n6608), .B2(n6707), .A(n7045), .ZN(n6611) );
  OAI21_X1 U7113 ( .B1(n6615), .B2(n6736), .A(n6659), .ZN(n6610) );
  OAI22_X1 U7114 ( .A1(n6720), .A2(n6619), .B1(n6611), .B2(n6610), .ZN(n6609)
         );
  AOI22_X1 U7115 ( .A1(n6734), .A2(n7045), .B1(n7044), .B2(n6745), .ZN(n6617)
         );
  INV_X1 U7116 ( .A(n6610), .ZN(n6612) );
  NAND2_X1 U7117 ( .A1(n6612), .A2(n6611), .ZN(n6613) );
  OAI211_X1 U7118 ( .C1(n6659), .C2(n6614), .A(n6685), .B(n6613), .ZN(n7046)
         );
  AOI22_X1 U7119 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n7046), .B1(n6725), 
        .B2(n7052), .ZN(n6616) );
  OAI211_X1 U7120 ( .C1(n7049), .C2(n6662), .A(n6617), .B(n6616), .ZN(U3092)
         );
  OAI22_X1 U7121 ( .A1(n6739), .A2(n6731), .B1(n6730), .B2(n6618), .ZN(n7051)
         );
  NOR2_X1 U7122 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6619), .ZN(n7050)
         );
  AOI22_X1 U7123 ( .A1(n6735), .A2(n7051), .B1(n6734), .B2(n7050), .ZN(n6625)
         );
  NAND2_X1 U7124 ( .A1(n6731), .A2(n6659), .ZN(n6738) );
  AND2_X1 U7125 ( .A1(n6641), .A2(n6663), .ZN(n6626) );
  AOI21_X1 U7126 ( .B1(n7061), .B2(n6974), .A(n6736), .ZN(n6620) );
  AOI21_X1 U7127 ( .B1(n6732), .B2(n6738), .A(n6620), .ZN(n6621) );
  NOR2_X1 U7128 ( .A1(n6621), .A2(n6740), .ZN(n6623) );
  AOI22_X1 U7129 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n7053), .B1(n6725), 
        .B2(n6971), .ZN(n6624) );
  OAI211_X1 U7130 ( .C1(n6728), .C2(n6974), .A(n6625), .B(n6624), .ZN(U3084)
         );
  INV_X1 U7131 ( .A(n6627), .ZN(n7056) );
  AOI22_X1 U7132 ( .A1(n6734), .A2(n7056), .B1(n6971), .B2(n6745), .ZN(n6637)
         );
  AND2_X1 U7133 ( .A1(n6628), .A2(n6659), .ZN(n6633) );
  NOR2_X1 U7134 ( .A1(n6630), .A2(n6629), .ZN(n6708) );
  AOI21_X1 U7135 ( .B1(n6708), .B2(n6631), .A(n7056), .ZN(n6634) );
  AOI22_X1 U7136 ( .A1(n6633), .A2(n6634), .B1(n6639), .B2(n6710), .ZN(n6632)
         );
  NAND2_X1 U7137 ( .A1(n6685), .A2(n6632), .ZN(n7058) );
  INV_X1 U7138 ( .A(n6633), .ZN(n6635) );
  OAI22_X1 U7139 ( .A1(n6635), .A2(n6634), .B1(n6639), .B2(n6720), .ZN(n7057)
         );
  AOI22_X1 U7140 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n7058), .B1(n6735), 
        .B2(n7057), .ZN(n6636) );
  OAI211_X1 U7141 ( .C1(n6748), .C2(n6936), .A(n6637), .B(n6636), .ZN(U3076)
         );
  NAND2_X1 U7142 ( .A1(n6677), .A2(n3500), .ZN(n6691) );
  OAI22_X1 U7143 ( .A1(n6732), .A2(n6638), .B1(n6669), .B2(n6691), .ZN(n7064)
         );
  NOR2_X1 U7144 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6639), .ZN(n7063)
         );
  AOI22_X1 U7145 ( .A1(n6735), .A2(n7064), .B1(n6734), .B2(n7063), .ZN(n6648)
         );
  OAI21_X1 U7146 ( .B1(n7072), .B2(n7065), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6645) );
  INV_X1 U7147 ( .A(n6642), .ZN(n6643) );
  NAND2_X1 U7148 ( .A1(n6643), .A2(n6739), .ZN(n6644) );
  AOI21_X1 U7149 ( .B1(n6645), .B2(n6644), .A(n6674), .ZN(n6646) );
  NAND2_X1 U7150 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6691), .ZN(n6703) );
  OAI211_X1 U7151 ( .C1(n7063), .C2(n6744), .A(n6646), .B(n6703), .ZN(n7066)
         );
  AOI22_X1 U7152 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n7066), .B1(n6725), 
        .B2(n7072), .ZN(n6647) );
  OAI211_X1 U7153 ( .C1(n6728), .C2(n6936), .A(n6648), .B(n6647), .ZN(U3068)
         );
  NOR3_X1 U7154 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6649), .ZN(n6658) );
  OAI21_X1 U7155 ( .B1(n6653), .B2(n6710), .A(n6699), .ZN(n6656) );
  NAND2_X1 U7156 ( .A1(n6708), .A2(n6650), .ZN(n6652) );
  INV_X1 U7157 ( .A(n6658), .ZN(n6671) );
  NOR2_X1 U7158 ( .A1(n6709), .A2(n6671), .ZN(n7071) );
  INV_X1 U7159 ( .A(n7071), .ZN(n6651) );
  NAND2_X1 U7160 ( .A1(n6652), .A2(n6651), .ZN(n6654) );
  AOI22_X1 U7161 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6658), .B1(n6656), .B2(
        n6654), .ZN(n7077) );
  AOI22_X1 U7162 ( .A1(n6734), .A2(n7071), .B1(n6725), .B2(n7080), .ZN(n6661)
         );
  INV_X1 U7163 ( .A(n6654), .ZN(n6655) );
  NAND2_X1 U7164 ( .A1(n6656), .A2(n6655), .ZN(n6657) );
  OAI211_X1 U7165 ( .C1(n6659), .C2(n6658), .A(n6685), .B(n6657), .ZN(n7073)
         );
  AOI22_X1 U7166 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n7073), .B1(n6745), 
        .B2(n7072), .ZN(n6660) );
  OAI211_X1 U7167 ( .C1(n7077), .C2(n6662), .A(n6661), .B(n6660), .ZN(U3060)
         );
  NAND2_X1 U7168 ( .A1(n6664), .A2(n6663), .ZN(n6665) );
  INV_X1 U7169 ( .A(n6676), .ZN(n6668) );
  NAND2_X1 U7170 ( .A1(n6668), .A2(n6667), .ZN(n6729) );
  OAI22_X1 U7171 ( .A1(n6732), .A2(n6670), .B1(n6669), .B2(n6729), .ZN(n7079)
         );
  NOR2_X1 U7172 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6671), .ZN(n7078)
         );
  AOI22_X1 U7173 ( .A1(n6735), .A2(n7079), .B1(n6734), .B2(n7078), .ZN(n6680)
         );
  AOI21_X1 U7174 ( .B1(n7084), .B2(n6984), .A(n6736), .ZN(n6672) );
  AOI21_X1 U7175 ( .B1(n6739), .B2(n6673), .A(n6672), .ZN(n6675) );
  NOR2_X1 U7176 ( .A1(n6675), .A2(n6674), .ZN(n6678) );
  OAI21_X1 U7177 ( .B1(n6677), .B2(n6676), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n6742) );
  AOI22_X1 U7178 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(n7081), .B1(n6745), 
        .B2(n7080), .ZN(n6679) );
  OAI211_X1 U7179 ( .C1(n6748), .C2(n7084), .A(n6680), .B(n6679), .ZN(U3052)
         );
  NOR2_X1 U7180 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6718) );
  INV_X1 U7181 ( .A(n6718), .ZN(n6733) );
  NOR2_X1 U7182 ( .A1(n6733), .A2(n6681), .ZN(n7086) );
  AOI22_X1 U7183 ( .A1(n6734), .A2(n7086), .B1(n7094), .B2(n6725), .ZN(n6690)
         );
  INV_X1 U7184 ( .A(n6682), .ZN(n6683) );
  AOI21_X1 U7185 ( .B1(n6683), .B2(STATEBS16_REG_SCAN_IN), .A(n6710), .ZN(
        n6686) );
  AOI21_X1 U7186 ( .B1(n6708), .B2(n6697), .A(n7086), .ZN(n6688) );
  NAND2_X1 U7187 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6718), .ZN(n6693) );
  AOI22_X1 U7188 ( .A1(n6686), .A2(n6688), .B1(n6710), .B2(n6693), .ZN(n6684)
         );
  NAND2_X1 U7189 ( .A1(n6685), .A2(n6684), .ZN(n7088) );
  INV_X1 U7190 ( .A(n6686), .ZN(n6687) );
  OAI22_X1 U7191 ( .A1(n6688), .A2(n6687), .B1(n6720), .B2(n6693), .ZN(n7087)
         );
  AOI22_X1 U7192 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n7088), .B1(n6735), 
        .B2(n7087), .ZN(n6689) );
  OAI211_X1 U7193 ( .C1(n6728), .C2(n7084), .A(n6690), .B(n6689), .ZN(U3044)
         );
  OAI22_X1 U7194 ( .A1(n6732), .A2(n6692), .B1(n6730), .B2(n6691), .ZN(n7093)
         );
  NOR2_X1 U7195 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6693), .ZN(n7092)
         );
  AOI22_X1 U7196 ( .A1(n6735), .A2(n7093), .B1(n6734), .B2(n7092), .ZN(n6706)
         );
  NAND2_X1 U7197 ( .A1(n6695), .A2(n6694), .ZN(n6724) );
  NAND2_X1 U7198 ( .A1(n7091), .A2(n7098), .ZN(n6700) );
  AOI22_X1 U7199 ( .A1(n6700), .A2(n6699), .B1(n6698), .B2(n6697), .ZN(n6701)
         );
  NOR2_X1 U7200 ( .A1(n6701), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6704) );
  INV_X1 U7201 ( .A(n6740), .ZN(n6702) );
  AOI22_X1 U7202 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n7095), .B1(n6725), 
        .B2(n7101), .ZN(n6705) );
  OAI211_X1 U7203 ( .C1(n6728), .C2(n7091), .A(n6706), .B(n6705), .ZN(U3036)
         );
  NAND2_X1 U7204 ( .A1(n6708), .A2(n6707), .ZN(n6714) );
  NOR3_X2 U7205 ( .A1(n6709), .A2(n6733), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n7099) );
  INV_X1 U7206 ( .A(n7099), .ZN(n6711) );
  AOI21_X1 U7207 ( .B1(n6714), .B2(n6711), .A(n6710), .ZN(n6713) );
  NOR3_X1 U7208 ( .A1(n6720), .A2(n6733), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6712) );
  AOI22_X1 U7209 ( .A1(n6735), .A2(n7100), .B1(n6734), .B2(n7099), .ZN(n6727)
         );
  INV_X1 U7210 ( .A(n6724), .ZN(n6716) );
  INV_X1 U7211 ( .A(n6714), .ZN(n6715) );
  AOI21_X1 U7212 ( .B1(n6716), .B2(STATEBS16_REG_SCAN_IN), .A(n6715), .ZN(
        n6721) );
  NAND2_X1 U7213 ( .A1(n6718), .A2(n6717), .ZN(n6719) );
  AOI221_X1 U7214 ( .B1(n6721), .B2(n6720), .C1(n6719), .C2(
        STATE2_REG_2__SCAN_IN), .A(STATE2_REG_3__SCAN_IN), .ZN(n6722) );
  OAI21_X1 U7215 ( .B1(n7099), .B2(n6722), .A(n6999), .ZN(n7102) );
  AOI22_X1 U7216 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n7102), .B1(n6725), 
        .B2(n7111), .ZN(n6726) );
  OAI211_X1 U7217 ( .C1(n6728), .C2(n7098), .A(n6727), .B(n6726), .ZN(U3028)
         );
  OAI22_X1 U7218 ( .A1(n6732), .A2(n6731), .B1(n6730), .B2(n6729), .ZN(n7108)
         );
  NOR3_X2 U7219 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6733), .ZN(n7106) );
  AOI22_X1 U7220 ( .A1(n6735), .A2(n7108), .B1(n6734), .B2(n7106), .ZN(n6747)
         );
  AOI21_X1 U7221 ( .B1(n7105), .B2(n7115), .A(n6736), .ZN(n6737) );
  AOI21_X1 U7222 ( .B1(n6739), .B2(n6738), .A(n6737), .ZN(n6741) );
  NOR2_X1 U7223 ( .A1(n6741), .A2(n6740), .ZN(n6743) );
  OAI211_X1 U7224 ( .C1(n7106), .C2(n6744), .A(n6743), .B(n6742), .ZN(n7112)
         );
  AOI22_X1 U7225 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n7112), .B1(n6745), 
        .B2(n7111), .ZN(n6746) );
  OAI211_X1 U7226 ( .C1(n6748), .C2(n7115), .A(n6747), .B(n6746), .ZN(U3020)
         );
  NOR2_X1 U7227 ( .A1(n7005), .A2(n6749), .ZN(n6772) );
  NAND2_X1 U7228 ( .A1(DATAI_1_), .A2(n6999), .ZN(n6775) );
  NOR2_X2 U7229 ( .A1(n7001), .A2(n6750), .ZN(n6784) );
  AOI22_X1 U7230 ( .A1(n6785), .A2(n7003), .B1(n6784), .B2(n7002), .ZN(n6753)
         );
  NOR2_X2 U7231 ( .A1(n7005), .A2(n6751), .ZN(n6786) );
  AOI22_X1 U7232 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n7007), .B1(n6786), 
        .B2(n7006), .ZN(n6752) );
  OAI211_X1 U7233 ( .C1(n6789), .C2(n7010), .A(n6753), .B(n6752), .ZN(U3141)
         );
  AOI22_X1 U7234 ( .A1(n6785), .A2(n7012), .B1(n6784), .B2(n7011), .ZN(n6755)
         );
  AOI22_X1 U7235 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n7014), .B1(n6786), 
        .B2(n7013), .ZN(n6754) );
  OAI211_X1 U7236 ( .C1(n6789), .C2(n7017), .A(n6755), .B(n6754), .ZN(U3133)
         );
  AOI22_X1 U7237 ( .A1(n6784), .A2(n7019), .B1(n7018), .B2(n6786), .ZN(n6757)
         );
  AOI22_X1 U7238 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n7021), .B1(n6785), 
        .B2(n7020), .ZN(n6756) );
  OAI211_X1 U7239 ( .C1(n6789), .C2(n7024), .A(n6757), .B(n6756), .ZN(U3125)
         );
  AOI22_X1 U7240 ( .A1(n6785), .A2(n7026), .B1(n6784), .B2(n7025), .ZN(n6759)
         );
  AOI22_X1 U7241 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n7028), .B1(n6786), 
        .B2(n7027), .ZN(n6758) );
  OAI211_X1 U7242 ( .C1(n6789), .C2(n7031), .A(n6759), .B(n6758), .ZN(U3117)
         );
  AOI22_X1 U7243 ( .A1(n6784), .A2(n7032), .B1(n7039), .B2(n6772), .ZN(n6761)
         );
  AOI22_X1 U7244 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n7034), .B1(n6786), 
        .B2(n7033), .ZN(n6760) );
  OAI211_X1 U7245 ( .C1(n7037), .C2(n6775), .A(n6761), .B(n6760), .ZN(U3109)
         );
  AOI22_X1 U7246 ( .A1(n6784), .A2(n7038), .B1(n7044), .B2(n6772), .ZN(n6763)
         );
  AOI22_X1 U7247 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n7040), .B1(n7039), 
        .B2(n6786), .ZN(n6762) );
  OAI211_X1 U7248 ( .C1(n7043), .C2(n6775), .A(n6763), .B(n6762), .ZN(U3101)
         );
  AOI22_X1 U7249 ( .A1(n6784), .A2(n7045), .B1(n7044), .B2(n6786), .ZN(n6765)
         );
  AOI22_X1 U7250 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n7046), .B1(n6772), 
        .B2(n7052), .ZN(n6764) );
  OAI211_X1 U7251 ( .C1(n7049), .C2(n6775), .A(n6765), .B(n6764), .ZN(U3093)
         );
  AOI22_X1 U7252 ( .A1(n6785), .A2(n7051), .B1(n6784), .B2(n7050), .ZN(n6767)
         );
  AOI22_X1 U7253 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(n7053), .B1(n6786), 
        .B2(n7052), .ZN(n6766) );
  OAI211_X1 U7254 ( .C1(n6789), .C2(n7061), .A(n6767), .B(n6766), .ZN(U3085)
         );
  AOI22_X1 U7255 ( .A1(n6784), .A2(n7056), .B1(n6786), .B2(n6971), .ZN(n6769)
         );
  AOI22_X1 U7256 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n7058), .B1(n6785), 
        .B2(n7057), .ZN(n6768) );
  OAI211_X1 U7257 ( .C1(n6789), .C2(n6936), .A(n6769), .B(n6768), .ZN(U3077)
         );
  AOI22_X1 U7258 ( .A1(n6785), .A2(n7064), .B1(n6784), .B2(n7063), .ZN(n6771)
         );
  AOI22_X1 U7259 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n7066), .B1(n6786), 
        .B2(n7065), .ZN(n6770) );
  OAI211_X1 U7260 ( .C1(n6789), .C2(n7069), .A(n6771), .B(n6770), .ZN(U3069)
         );
  AOI22_X1 U7261 ( .A1(n6784), .A2(n7071), .B1(n7080), .B2(n6772), .ZN(n6774)
         );
  AOI22_X1 U7262 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n7073), .B1(n6786), 
        .B2(n7072), .ZN(n6773) );
  OAI211_X1 U7263 ( .C1(n7077), .C2(n6775), .A(n6774), .B(n6773), .ZN(U3061)
         );
  AOI22_X1 U7264 ( .A1(n6785), .A2(n7079), .B1(n6784), .B2(n7078), .ZN(n6777)
         );
  AOI22_X1 U7265 ( .A1(INSTQUEUE_REG_4__1__SCAN_IN), .A2(n7081), .B1(n6786), 
        .B2(n7080), .ZN(n6776) );
  OAI211_X1 U7266 ( .C1(n6789), .C2(n7084), .A(n6777), .B(n6776), .ZN(U3053)
         );
  AOI22_X1 U7267 ( .A1(n6784), .A2(n7086), .B1(n6786), .B2(n7085), .ZN(n6779)
         );
  AOI22_X1 U7268 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n7088), .B1(n6785), 
        .B2(n7087), .ZN(n6778) );
  OAI211_X1 U7269 ( .C1(n7091), .C2(n6789), .A(n6779), .B(n6778), .ZN(U3045)
         );
  AOI22_X1 U7270 ( .A1(n6785), .A2(n7093), .B1(n6784), .B2(n7092), .ZN(n6781)
         );
  AOI22_X1 U7271 ( .A1(INSTQUEUE_REG_2__1__SCAN_IN), .A2(n7095), .B1(n7094), 
        .B2(n6786), .ZN(n6780) );
  OAI211_X1 U7272 ( .C1(n7098), .C2(n6789), .A(n6781), .B(n6780), .ZN(U3037)
         );
  AOI22_X1 U7273 ( .A1(n6785), .A2(n7100), .B1(n6784), .B2(n7099), .ZN(n6783)
         );
  AOI22_X1 U7274 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n7102), .B1(n7101), 
        .B2(n6786), .ZN(n6782) );
  OAI211_X1 U7275 ( .C1(n7105), .C2(n6789), .A(n6783), .B(n6782), .ZN(U3029)
         );
  AOI22_X1 U7276 ( .A1(n6785), .A2(n7108), .B1(n6784), .B2(n7106), .ZN(n6788)
         );
  AOI22_X1 U7277 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(n7112), .B1(n7111), 
        .B2(n6786), .ZN(n6787) );
  OAI211_X1 U7278 ( .C1(n6789), .C2(n7115), .A(n6788), .B(n6787), .ZN(U3021)
         );
  INV_X1 U7279 ( .A(n6821), .ZN(n6830) );
  NAND2_X1 U7280 ( .A1(DATAI_2_), .A2(n6999), .ZN(n6814) );
  NOR2_X2 U7281 ( .A1(n7001), .A2(n6790), .ZN(n6825) );
  AOI22_X1 U7282 ( .A1(n6826), .A2(n7003), .B1(n6825), .B2(n7002), .ZN(n6793)
         );
  NOR2_X1 U7283 ( .A1(n7005), .A2(n6791), .ZN(n6827) );
  AOI22_X1 U7284 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(n7007), .B1(n6827), 
        .B2(n7006), .ZN(n6792) );
  OAI211_X1 U7285 ( .C1(n6830), .C2(n7010), .A(n6793), .B(n6792), .ZN(U3142)
         );
  INV_X1 U7286 ( .A(n6827), .ZN(n6824) );
  AOI22_X1 U7287 ( .A1(n6826), .A2(n7012), .B1(n6825), .B2(n7011), .ZN(n6795)
         );
  AOI22_X1 U7288 ( .A1(INSTQUEUE_REG_14__2__SCAN_IN), .A2(n7014), .B1(n6821), 
        .B2(n7018), .ZN(n6794) );
  OAI211_X1 U7289 ( .C1(n6824), .C2(n7010), .A(n6795), .B(n6794), .ZN(U3134)
         );
  AOI22_X1 U7290 ( .A1(n6825), .A2(n7019), .B1(n7027), .B2(n6821), .ZN(n6797)
         );
  AOI22_X1 U7291 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n7021), .B1(n6826), 
        .B2(n7020), .ZN(n6796) );
  OAI211_X1 U7292 ( .C1(n6824), .C2(n7017), .A(n6797), .B(n6796), .ZN(U3126)
         );
  AOI22_X1 U7293 ( .A1(n6826), .A2(n7026), .B1(n6825), .B2(n7025), .ZN(n6799)
         );
  AOI22_X1 U7294 ( .A1(INSTQUEUE_REG_12__2__SCAN_IN), .A2(n7028), .B1(n6821), 
        .B2(n7033), .ZN(n6798) );
  OAI211_X1 U7295 ( .C1(n6824), .C2(n7024), .A(n6799), .B(n6798), .ZN(U3118)
         );
  AOI22_X1 U7296 ( .A1(n6825), .A2(n7032), .B1(n7039), .B2(n6821), .ZN(n6801)
         );
  AOI22_X1 U7297 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n7034), .B1(n6827), 
        .B2(n7033), .ZN(n6800) );
  OAI211_X1 U7298 ( .C1(n7037), .C2(n6814), .A(n6801), .B(n6800), .ZN(U3110)
         );
  AOI22_X1 U7299 ( .A1(n6825), .A2(n7038), .B1(n7044), .B2(n6821), .ZN(n6803)
         );
  AOI22_X1 U7300 ( .A1(INSTQUEUE_REG_10__2__SCAN_IN), .A2(n7040), .B1(n7039), 
        .B2(n6827), .ZN(n6802) );
  OAI211_X1 U7301 ( .C1(n7043), .C2(n6814), .A(n6803), .B(n6802), .ZN(U3102)
         );
  AOI22_X1 U7302 ( .A1(n6825), .A2(n7045), .B1(n6821), .B2(n7052), .ZN(n6805)
         );
  AOI22_X1 U7303 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n7046), .B1(n7044), 
        .B2(n6827), .ZN(n6804) );
  OAI211_X1 U7304 ( .C1(n7049), .C2(n6814), .A(n6805), .B(n6804), .ZN(U3094)
         );
  AOI22_X1 U7305 ( .A1(n6826), .A2(n7051), .B1(n6825), .B2(n7050), .ZN(n6807)
         );
  AOI22_X1 U7306 ( .A1(INSTQUEUE_REG_8__2__SCAN_IN), .A2(n7053), .B1(n6821), 
        .B2(n6971), .ZN(n6806) );
  OAI211_X1 U7307 ( .C1(n6824), .C2(n6974), .A(n6807), .B(n6806), .ZN(U3086)
         );
  AOI22_X1 U7308 ( .A1(n6825), .A2(n7056), .B1(n6821), .B2(n7065), .ZN(n6809)
         );
  AOI22_X1 U7309 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n7058), .B1(n6826), 
        .B2(n7057), .ZN(n6808) );
  OAI211_X1 U7310 ( .C1(n6824), .C2(n7061), .A(n6809), .B(n6808), .ZN(U3078)
         );
  AOI22_X1 U7311 ( .A1(n6826), .A2(n7064), .B1(n6825), .B2(n7063), .ZN(n6811)
         );
  AOI22_X1 U7312 ( .A1(INSTQUEUE_REG_6__2__SCAN_IN), .A2(n7066), .B1(n6821), 
        .B2(n7072), .ZN(n6810) );
  OAI211_X1 U7313 ( .C1(n6824), .C2(n6936), .A(n6811), .B(n6810), .ZN(U3070)
         );
  AOI22_X1 U7314 ( .A1(n6825), .A2(n7071), .B1(n6827), .B2(n7072), .ZN(n6813)
         );
  AOI22_X1 U7315 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n7073), .B1(n6821), 
        .B2(n7080), .ZN(n6812) );
  OAI211_X1 U7316 ( .C1(n7077), .C2(n6814), .A(n6813), .B(n6812), .ZN(U3062)
         );
  AOI22_X1 U7317 ( .A1(n6826), .A2(n7079), .B1(n6825), .B2(n7078), .ZN(n6816)
         );
  AOI22_X1 U7318 ( .A1(INSTQUEUE_REG_4__2__SCAN_IN), .A2(n7081), .B1(n6821), 
        .B2(n7085), .ZN(n6815) );
  OAI211_X1 U7319 ( .C1(n6824), .C2(n6984), .A(n6816), .B(n6815), .ZN(U3054)
         );
  AOI22_X1 U7320 ( .A1(n6825), .A2(n7086), .B1(n7085), .B2(n6827), .ZN(n6818)
         );
  AOI22_X1 U7321 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n7088), .B1(n6826), 
        .B2(n7087), .ZN(n6817) );
  OAI211_X1 U7322 ( .C1(n7091), .C2(n6830), .A(n6818), .B(n6817), .ZN(U3046)
         );
  AOI22_X1 U7323 ( .A1(n6826), .A2(n7093), .B1(n6825), .B2(n7092), .ZN(n6820)
         );
  AOI22_X1 U7324 ( .A1(INSTQUEUE_REG_2__2__SCAN_IN), .A2(n7095), .B1(n7101), 
        .B2(n6821), .ZN(n6819) );
  OAI211_X1 U7325 ( .C1(n7091), .C2(n6824), .A(n6820), .B(n6819), .ZN(U3038)
         );
  AOI22_X1 U7326 ( .A1(n6826), .A2(n7100), .B1(n6825), .B2(n7099), .ZN(n6823)
         );
  AOI22_X1 U7327 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n7102), .B1(n7111), 
        .B2(n6821), .ZN(n6822) );
  OAI211_X1 U7328 ( .C1(n7098), .C2(n6824), .A(n6823), .B(n6822), .ZN(U3030)
         );
  AOI22_X1 U7329 ( .A1(n6826), .A2(n7108), .B1(n6825), .B2(n7106), .ZN(n6829)
         );
  AOI22_X1 U7330 ( .A1(INSTQUEUE_REG_0__2__SCAN_IN), .A2(n7112), .B1(n7111), 
        .B2(n6827), .ZN(n6828) );
  OAI211_X1 U7331 ( .C1(n6830), .C2(n7115), .A(n6829), .B(n6828), .ZN(U3022)
         );
  AND2_X1 U7332 ( .A1(n5804), .A2(DATAI_27_), .ZN(n6858) );
  INV_X1 U7333 ( .A(n6858), .ZN(n6871) );
  NAND2_X1 U7334 ( .A1(DATAI_3_), .A2(n6999), .ZN(n6855) );
  NOR2_X2 U7335 ( .A1(n7001), .A2(n6831), .ZN(n6866) );
  AOI22_X1 U7336 ( .A1(n6867), .A2(n7003), .B1(n6866), .B2(n7002), .ZN(n6834)
         );
  NOR2_X1 U7337 ( .A1(n7005), .A2(n6832), .ZN(n6868) );
  AOI22_X1 U7338 ( .A1(INSTQUEUE_REG_15__3__SCAN_IN), .A2(n7007), .B1(n6868), 
        .B2(n7006), .ZN(n6833) );
  OAI211_X1 U7339 ( .C1(n6871), .C2(n7010), .A(n6834), .B(n6833), .ZN(U3143)
         );
  AOI22_X1 U7340 ( .A1(n6867), .A2(n7012), .B1(n6866), .B2(n7011), .ZN(n6836)
         );
  AOI22_X1 U7341 ( .A1(INSTQUEUE_REG_14__3__SCAN_IN), .A2(n7014), .B1(n6868), 
        .B2(n7013), .ZN(n6835) );
  OAI211_X1 U7342 ( .C1(n6871), .C2(n7017), .A(n6836), .B(n6835), .ZN(U3135)
         );
  INV_X1 U7343 ( .A(n6868), .ZN(n6861) );
  AOI22_X1 U7344 ( .A1(n6866), .A2(n7019), .B1(n7027), .B2(n6858), .ZN(n6838)
         );
  AOI22_X1 U7345 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n7021), .B1(n6867), 
        .B2(n7020), .ZN(n6837) );
  OAI211_X1 U7346 ( .C1(n6861), .C2(n7017), .A(n6838), .B(n6837), .ZN(U3127)
         );
  AOI22_X1 U7347 ( .A1(n6867), .A2(n7026), .B1(n6866), .B2(n7025), .ZN(n6840)
         );
  AOI22_X1 U7348 ( .A1(INSTQUEUE_REG_12__3__SCAN_IN), .A2(n7028), .B1(n6868), 
        .B2(n7027), .ZN(n6839) );
  OAI211_X1 U7349 ( .C1(n6871), .C2(n7031), .A(n6840), .B(n6839), .ZN(U3119)
         );
  AOI22_X1 U7350 ( .A1(n6866), .A2(n7032), .B1(n7033), .B2(n6868), .ZN(n6842)
         );
  AOI22_X1 U7351 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n7034), .B1(n7039), 
        .B2(n6858), .ZN(n6841) );
  OAI211_X1 U7352 ( .C1(n7037), .C2(n6855), .A(n6842), .B(n6841), .ZN(U3111)
         );
  AOI22_X1 U7353 ( .A1(n6866), .A2(n7038), .B1(n7044), .B2(n6858), .ZN(n6844)
         );
  AOI22_X1 U7354 ( .A1(INSTQUEUE_REG_10__3__SCAN_IN), .A2(n7040), .B1(n7039), 
        .B2(n6868), .ZN(n6843) );
  OAI211_X1 U7355 ( .C1(n7043), .C2(n6855), .A(n6844), .B(n6843), .ZN(U3103)
         );
  AOI22_X1 U7356 ( .A1(n6866), .A2(n7045), .B1(n6858), .B2(n7052), .ZN(n6846)
         );
  AOI22_X1 U7357 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n7046), .B1(n7044), 
        .B2(n6868), .ZN(n6845) );
  OAI211_X1 U7358 ( .C1(n7049), .C2(n6855), .A(n6846), .B(n6845), .ZN(U3095)
         );
  AOI22_X1 U7359 ( .A1(n6867), .A2(n7051), .B1(n6866), .B2(n7050), .ZN(n6848)
         );
  AOI22_X1 U7360 ( .A1(INSTQUEUE_REG_8__3__SCAN_IN), .A2(n7053), .B1(n6858), 
        .B2(n6971), .ZN(n6847) );
  OAI211_X1 U7361 ( .C1(n6861), .C2(n6974), .A(n6848), .B(n6847), .ZN(U3087)
         );
  AOI22_X1 U7362 ( .A1(n6866), .A2(n7056), .B1(n6858), .B2(n7065), .ZN(n6850)
         );
  AOI22_X1 U7363 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n7058), .B1(n6867), 
        .B2(n7057), .ZN(n6849) );
  OAI211_X1 U7364 ( .C1(n6861), .C2(n7061), .A(n6850), .B(n6849), .ZN(U3079)
         );
  AOI22_X1 U7365 ( .A1(n6867), .A2(n7064), .B1(n6866), .B2(n7063), .ZN(n6852)
         );
  AOI22_X1 U7366 ( .A1(INSTQUEUE_REG_6__3__SCAN_IN), .A2(n7066), .B1(n6868), 
        .B2(n7065), .ZN(n6851) );
  OAI211_X1 U7367 ( .C1(n6871), .C2(n7069), .A(n6852), .B(n6851), .ZN(U3071)
         );
  AOI22_X1 U7368 ( .A1(n6866), .A2(n7071), .B1(n7072), .B2(n6868), .ZN(n6854)
         );
  AOI22_X1 U7369 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n7073), .B1(n6858), 
        .B2(n7080), .ZN(n6853) );
  OAI211_X1 U7370 ( .C1(n7077), .C2(n6855), .A(n6854), .B(n6853), .ZN(U3063)
         );
  AOI22_X1 U7371 ( .A1(n6867), .A2(n7079), .B1(n6866), .B2(n7078), .ZN(n6857)
         );
  AOI22_X1 U7372 ( .A1(INSTQUEUE_REG_4__3__SCAN_IN), .A2(n7081), .B1(n6858), 
        .B2(n7085), .ZN(n6856) );
  OAI211_X1 U7373 ( .C1(n6861), .C2(n6984), .A(n6857), .B(n6856), .ZN(U3055)
         );
  AOI22_X1 U7374 ( .A1(n6866), .A2(n7086), .B1(n7094), .B2(n6858), .ZN(n6860)
         );
  AOI22_X1 U7375 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n7088), .B1(n6867), 
        .B2(n7087), .ZN(n6859) );
  OAI211_X1 U7376 ( .C1(n6861), .C2(n7084), .A(n6860), .B(n6859), .ZN(U3047)
         );
  AOI22_X1 U7377 ( .A1(n6867), .A2(n7093), .B1(n6866), .B2(n7092), .ZN(n6863)
         );
  AOI22_X1 U7378 ( .A1(INSTQUEUE_REG_2__3__SCAN_IN), .A2(n7095), .B1(n7094), 
        .B2(n6868), .ZN(n6862) );
  OAI211_X1 U7379 ( .C1(n7098), .C2(n6871), .A(n6863), .B(n6862), .ZN(U3039)
         );
  AOI22_X1 U7380 ( .A1(n6867), .A2(n7100), .B1(n6866), .B2(n7099), .ZN(n6865)
         );
  AOI22_X1 U7381 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n7102), .B1(n7101), 
        .B2(n6868), .ZN(n6864) );
  OAI211_X1 U7382 ( .C1(n7105), .C2(n6871), .A(n6865), .B(n6864), .ZN(U3031)
         );
  AOI22_X1 U7383 ( .A1(n6867), .A2(n7108), .B1(n6866), .B2(n7106), .ZN(n6870)
         );
  AOI22_X1 U7384 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(n7112), .B1(n7111), 
        .B2(n6868), .ZN(n6869) );
  OAI211_X1 U7385 ( .C1(n6871), .C2(n7115), .A(n6870), .B(n6869), .ZN(U3023)
         );
  AND2_X1 U7386 ( .A1(n5804), .A2(DATAI_20_), .ZN(n6909) );
  INV_X1 U7387 ( .A(n6909), .ZN(n6906) );
  NAND2_X1 U7388 ( .A1(DATAI_4_), .A2(n6999), .ZN(n6896) );
  NOR2_X2 U7389 ( .A1(n7001), .A2(n6872), .ZN(n6907) );
  AOI22_X1 U7390 ( .A1(n6908), .A2(n7003), .B1(n6907), .B2(n7002), .ZN(n6875)
         );
  NOR2_X2 U7391 ( .A1(n7005), .A2(n6873), .ZN(n6903) );
  AOI22_X1 U7392 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n7007), .B1(n6903), 
        .B2(n7013), .ZN(n6874) );
  OAI211_X1 U7393 ( .C1(n6906), .C2(n7115), .A(n6875), .B(n6874), .ZN(U3144)
         );
  AOI22_X1 U7394 ( .A1(n6908), .A2(n7012), .B1(n6907), .B2(n7011), .ZN(n6877)
         );
  AOI22_X1 U7395 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n7014), .B1(n6903), 
        .B2(n7018), .ZN(n6876) );
  OAI211_X1 U7396 ( .C1(n6906), .C2(n7010), .A(n6877), .B(n6876), .ZN(U3136)
         );
  AOI22_X1 U7397 ( .A1(n6907), .A2(n7019), .B1(n7027), .B2(n6903), .ZN(n6879)
         );
  AOI22_X1 U7398 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n7021), .B1(n6908), 
        .B2(n7020), .ZN(n6878) );
  OAI211_X1 U7399 ( .C1(n6906), .C2(n7017), .A(n6879), .B(n6878), .ZN(U3128)
         );
  AOI22_X1 U7400 ( .A1(n6908), .A2(n7026), .B1(n6907), .B2(n7025), .ZN(n6881)
         );
  AOI22_X1 U7401 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n7028), .B1(n6903), 
        .B2(n7033), .ZN(n6880) );
  OAI211_X1 U7402 ( .C1(n6906), .C2(n7024), .A(n6881), .B(n6880), .ZN(U3120)
         );
  AOI22_X1 U7403 ( .A1(n6907), .A2(n7032), .B1(n7039), .B2(n6903), .ZN(n6883)
         );
  AOI22_X1 U7404 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n7034), .B1(n6909), 
        .B2(n7033), .ZN(n6882) );
  OAI211_X1 U7405 ( .C1(n7037), .C2(n6896), .A(n6883), .B(n6882), .ZN(U3112)
         );
  AOI22_X1 U7406 ( .A1(n6907), .A2(n7038), .B1(n7044), .B2(n6903), .ZN(n6885)
         );
  AOI22_X1 U7407 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n7040), .B1(n7039), 
        .B2(n6909), .ZN(n6884) );
  OAI211_X1 U7408 ( .C1(n7043), .C2(n6896), .A(n6885), .B(n6884), .ZN(U3104)
         );
  AOI22_X1 U7409 ( .A1(n6907), .A2(n7045), .B1(n7044), .B2(n6909), .ZN(n6887)
         );
  AOI22_X1 U7410 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n7046), .B1(n6903), 
        .B2(n7052), .ZN(n6886) );
  OAI211_X1 U7411 ( .C1(n7049), .C2(n6896), .A(n6887), .B(n6886), .ZN(U3096)
         );
  AOI22_X1 U7412 ( .A1(n6908), .A2(n7051), .B1(n6907), .B2(n7050), .ZN(n6889)
         );
  AOI22_X1 U7413 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n7053), .B1(n6903), 
        .B2(n6971), .ZN(n6888) );
  OAI211_X1 U7414 ( .C1(n6906), .C2(n6974), .A(n6889), .B(n6888), .ZN(U3088)
         );
  INV_X1 U7415 ( .A(n6903), .ZN(n6912) );
  AOI22_X1 U7416 ( .A1(n6907), .A2(n7056), .B1(n6909), .B2(n6971), .ZN(n6891)
         );
  AOI22_X1 U7417 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n7058), .B1(n6908), 
        .B2(n7057), .ZN(n6890) );
  OAI211_X1 U7418 ( .C1(n6912), .C2(n6936), .A(n6891), .B(n6890), .ZN(U3080)
         );
  AOI22_X1 U7419 ( .A1(n6908), .A2(n7064), .B1(n6907), .B2(n7063), .ZN(n6893)
         );
  AOI22_X1 U7420 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n7066), .B1(n6903), 
        .B2(n7072), .ZN(n6892) );
  OAI211_X1 U7421 ( .C1(n6906), .C2(n6936), .A(n6893), .B(n6892), .ZN(U3072)
         );
  AOI22_X1 U7422 ( .A1(n6907), .A2(n7071), .B1(n6909), .B2(n7072), .ZN(n6895)
         );
  AOI22_X1 U7423 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n7073), .B1(n6903), 
        .B2(n7080), .ZN(n6894) );
  OAI211_X1 U7424 ( .C1(n7077), .C2(n6896), .A(n6895), .B(n6894), .ZN(U3064)
         );
  AOI22_X1 U7425 ( .A1(n6908), .A2(n7079), .B1(n6907), .B2(n7078), .ZN(n6898)
         );
  AOI22_X1 U7426 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n7081), .B1(n6903), 
        .B2(n7085), .ZN(n6897) );
  OAI211_X1 U7427 ( .C1(n6906), .C2(n6984), .A(n6898), .B(n6897), .ZN(U3056)
         );
  AOI22_X1 U7428 ( .A1(n6907), .A2(n7086), .B1(n7085), .B2(n6909), .ZN(n6900)
         );
  AOI22_X1 U7429 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n7088), .B1(n6908), 
        .B2(n7087), .ZN(n6899) );
  OAI211_X1 U7430 ( .C1(n7091), .C2(n6912), .A(n6900), .B(n6899), .ZN(U3048)
         );
  AOI22_X1 U7431 ( .A1(n6908), .A2(n7093), .B1(n6907), .B2(n7092), .ZN(n6902)
         );
  AOI22_X1 U7432 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n7095), .B1(n7101), 
        .B2(n6903), .ZN(n6901) );
  OAI211_X1 U7433 ( .C1(n7091), .C2(n6906), .A(n6902), .B(n6901), .ZN(U3040)
         );
  AOI22_X1 U7434 ( .A1(n6908), .A2(n7100), .B1(n6907), .B2(n7099), .ZN(n6905)
         );
  AOI22_X1 U7435 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n7102), .B1(n7111), 
        .B2(n6903), .ZN(n6904) );
  OAI211_X1 U7436 ( .C1(n7098), .C2(n6906), .A(n6905), .B(n6904), .ZN(U3032)
         );
  AOI22_X1 U7437 ( .A1(n6908), .A2(n7108), .B1(n6907), .B2(n7106), .ZN(n6911)
         );
  AOI22_X1 U7438 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n7112), .B1(n7111), 
        .B2(n6909), .ZN(n6910) );
  OAI211_X1 U7439 ( .C1(n6912), .C2(n7115), .A(n6911), .B(n6910), .ZN(U3024)
         );
  NOR2_X1 U7440 ( .A1(n7005), .A2(n6913), .ZN(n6937) );
  INV_X1 U7441 ( .A(n6937), .ZN(n6954) );
  NAND2_X1 U7442 ( .A1(DATAI_5_), .A2(n6999), .ZN(n6940) );
  NOR2_X2 U7443 ( .A1(n7001), .A2(n6914), .ZN(n6949) );
  AOI22_X1 U7444 ( .A1(n6950), .A2(n7003), .B1(n6949), .B2(n7002), .ZN(n6917)
         );
  NOR2_X2 U7445 ( .A1(n7005), .A2(n6915), .ZN(n6951) );
  AOI22_X1 U7446 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n7007), .B1(n6951), 
        .B2(n7013), .ZN(n6916) );
  OAI211_X1 U7447 ( .C1(n6954), .C2(n7115), .A(n6917), .B(n6916), .ZN(U3145)
         );
  AOI22_X1 U7448 ( .A1(n6950), .A2(n7012), .B1(n6949), .B2(n7011), .ZN(n6919)
         );
  AOI22_X1 U7449 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(n7014), .B1(n6951), 
        .B2(n7018), .ZN(n6918) );
  OAI211_X1 U7450 ( .C1(n6954), .C2(n7010), .A(n6919), .B(n6918), .ZN(U3137)
         );
  AOI22_X1 U7451 ( .A1(n6949), .A2(n7019), .B1(n7027), .B2(n6951), .ZN(n6921)
         );
  AOI22_X1 U7452 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n7021), .B1(n6950), 
        .B2(n7020), .ZN(n6920) );
  OAI211_X1 U7453 ( .C1(n6954), .C2(n7017), .A(n6921), .B(n6920), .ZN(U3129)
         );
  AOI22_X1 U7454 ( .A1(n6950), .A2(n7026), .B1(n6949), .B2(n7025), .ZN(n6923)
         );
  AOI22_X1 U7455 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n7028), .B1(n6951), 
        .B2(n7033), .ZN(n6922) );
  OAI211_X1 U7456 ( .C1(n6954), .C2(n7024), .A(n6923), .B(n6922), .ZN(U3121)
         );
  AOI22_X1 U7457 ( .A1(n6949), .A2(n7032), .B1(n7039), .B2(n6951), .ZN(n6925)
         );
  AOI22_X1 U7458 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n7034), .B1(n6937), 
        .B2(n7033), .ZN(n6924) );
  OAI211_X1 U7459 ( .C1(n7037), .C2(n6940), .A(n6925), .B(n6924), .ZN(U3113)
         );
  AOI22_X1 U7460 ( .A1(n6949), .A2(n7038), .B1(n7044), .B2(n6951), .ZN(n6927)
         );
  AOI22_X1 U7461 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n7040), .B1(n7039), 
        .B2(n6937), .ZN(n6926) );
  OAI211_X1 U7462 ( .C1(n7043), .C2(n6940), .A(n6927), .B(n6926), .ZN(U3105)
         );
  AOI22_X1 U7463 ( .A1(n6949), .A2(n7045), .B1(n6951), .B2(n7052), .ZN(n6929)
         );
  AOI22_X1 U7464 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n7046), .B1(n7044), 
        .B2(n6937), .ZN(n6928) );
  OAI211_X1 U7465 ( .C1(n7049), .C2(n6940), .A(n6929), .B(n6928), .ZN(U3097)
         );
  AOI22_X1 U7466 ( .A1(n6950), .A2(n7051), .B1(n6949), .B2(n7050), .ZN(n6931)
         );
  AOI22_X1 U7467 ( .A1(INSTQUEUE_REG_8__5__SCAN_IN), .A2(n7053), .B1(n6951), 
        .B2(n6971), .ZN(n6930) );
  OAI211_X1 U7468 ( .C1(n6954), .C2(n6974), .A(n6931), .B(n6930), .ZN(U3089)
         );
  AOI22_X1 U7469 ( .A1(n6949), .A2(n7056), .B1(n6951), .B2(n7065), .ZN(n6933)
         );
  AOI22_X1 U7470 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n7058), .B1(n6950), 
        .B2(n7057), .ZN(n6932) );
  OAI211_X1 U7471 ( .C1(n6954), .C2(n7061), .A(n6933), .B(n6932), .ZN(U3081)
         );
  AOI22_X1 U7472 ( .A1(n6950), .A2(n7064), .B1(n6949), .B2(n7063), .ZN(n6935)
         );
  AOI22_X1 U7473 ( .A1(INSTQUEUE_REG_6__5__SCAN_IN), .A2(n7066), .B1(n6951), 
        .B2(n7072), .ZN(n6934) );
  OAI211_X1 U7474 ( .C1(n6954), .C2(n6936), .A(n6935), .B(n6934), .ZN(U3073)
         );
  AOI22_X1 U7475 ( .A1(n6949), .A2(n7071), .B1(n6951), .B2(n7080), .ZN(n6939)
         );
  AOI22_X1 U7476 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n7073), .B1(n6937), 
        .B2(n7072), .ZN(n6938) );
  OAI211_X1 U7477 ( .C1(n7077), .C2(n6940), .A(n6939), .B(n6938), .ZN(U3065)
         );
  AOI22_X1 U7478 ( .A1(n6950), .A2(n7079), .B1(n6949), .B2(n7078), .ZN(n6942)
         );
  AOI22_X1 U7479 ( .A1(INSTQUEUE_REG_4__5__SCAN_IN), .A2(n7081), .B1(n6951), 
        .B2(n7085), .ZN(n6941) );
  OAI211_X1 U7480 ( .C1(n6954), .C2(n6984), .A(n6942), .B(n6941), .ZN(U3057)
         );
  AOI22_X1 U7481 ( .A1(n6949), .A2(n7086), .B1(n7094), .B2(n6951), .ZN(n6944)
         );
  AOI22_X1 U7482 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n7088), .B1(n6950), 
        .B2(n7087), .ZN(n6943) );
  OAI211_X1 U7483 ( .C1(n6954), .C2(n7084), .A(n6944), .B(n6943), .ZN(U3049)
         );
  AOI22_X1 U7484 ( .A1(n6950), .A2(n7093), .B1(n6949), .B2(n7092), .ZN(n6946)
         );
  AOI22_X1 U7485 ( .A1(INSTQUEUE_REG_2__5__SCAN_IN), .A2(n7095), .B1(n7101), 
        .B2(n6951), .ZN(n6945) );
  OAI211_X1 U7486 ( .C1(n7091), .C2(n6954), .A(n6946), .B(n6945), .ZN(U3041)
         );
  AOI22_X1 U7487 ( .A1(n6950), .A2(n7100), .B1(n6949), .B2(n7099), .ZN(n6948)
         );
  AOI22_X1 U7488 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n7102), .B1(n7111), 
        .B2(n6951), .ZN(n6947) );
  OAI211_X1 U7489 ( .C1(n7098), .C2(n6954), .A(n6948), .B(n6947), .ZN(U3033)
         );
  AOI22_X1 U7490 ( .A1(n6950), .A2(n7108), .B1(n6949), .B2(n7106), .ZN(n6953)
         );
  AOI22_X1 U7491 ( .A1(INSTQUEUE_REG_0__5__SCAN_IN), .A2(n7112), .B1(n6951), 
        .B2(n7006), .ZN(n6952) );
  OAI211_X1 U7492 ( .C1(n7105), .C2(n6954), .A(n6953), .B(n6952), .ZN(U3025)
         );
  INV_X1 U7493 ( .A(n6989), .ZN(n6998) );
  NAND2_X1 U7494 ( .A1(DATAI_6_), .A2(n6999), .ZN(n6981) );
  NOR2_X2 U7495 ( .A1(n7001), .A2(n6955), .ZN(n6993) );
  AOI22_X1 U7496 ( .A1(n6994), .A2(n7003), .B1(n6993), .B2(n7002), .ZN(n6958)
         );
  NOR2_X1 U7497 ( .A1(n7005), .A2(n6956), .ZN(n6995) );
  AOI22_X1 U7498 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n7007), .B1(n6995), 
        .B2(n7006), .ZN(n6957) );
  OAI211_X1 U7499 ( .C1(n6998), .C2(n7010), .A(n6958), .B(n6957), .ZN(U3146)
         );
  INV_X1 U7500 ( .A(n6995), .ZN(n6992) );
  AOI22_X1 U7501 ( .A1(n6994), .A2(n7012), .B1(n6993), .B2(n7011), .ZN(n6960)
         );
  AOI22_X1 U7502 ( .A1(INSTQUEUE_REG_14__6__SCAN_IN), .A2(n7014), .B1(n6989), 
        .B2(n7018), .ZN(n6959) );
  OAI211_X1 U7503 ( .C1(n6992), .C2(n7010), .A(n6960), .B(n6959), .ZN(U3138)
         );
  AOI22_X1 U7504 ( .A1(n6993), .A2(n7019), .B1(n7018), .B2(n6995), .ZN(n6962)
         );
  AOI22_X1 U7505 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n7021), .B1(n6994), 
        .B2(n7020), .ZN(n6961) );
  OAI211_X1 U7506 ( .C1(n6998), .C2(n7024), .A(n6962), .B(n6961), .ZN(U3130)
         );
  AOI22_X1 U7507 ( .A1(n6994), .A2(n7026), .B1(n6993), .B2(n7025), .ZN(n6964)
         );
  AOI22_X1 U7508 ( .A1(INSTQUEUE_REG_12__6__SCAN_IN), .A2(n7028), .B1(n6995), 
        .B2(n7027), .ZN(n6963) );
  OAI211_X1 U7509 ( .C1(n6998), .C2(n7031), .A(n6964), .B(n6963), .ZN(U3122)
         );
  AOI22_X1 U7510 ( .A1(n6993), .A2(n7032), .B1(n7039), .B2(n6989), .ZN(n6966)
         );
  AOI22_X1 U7511 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n7034), .B1(n6995), 
        .B2(n7033), .ZN(n6965) );
  OAI211_X1 U7512 ( .C1(n7037), .C2(n6981), .A(n6966), .B(n6965), .ZN(U3114)
         );
  AOI22_X1 U7513 ( .A1(n6993), .A2(n7038), .B1(n7044), .B2(n6989), .ZN(n6968)
         );
  AOI22_X1 U7514 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(n7040), .B1(n7039), 
        .B2(n6995), .ZN(n6967) );
  OAI211_X1 U7515 ( .C1(n7043), .C2(n6981), .A(n6968), .B(n6967), .ZN(U3106)
         );
  AOI22_X1 U7516 ( .A1(n6993), .A2(n7045), .B1(n6989), .B2(n7052), .ZN(n6970)
         );
  AOI22_X1 U7517 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n7046), .B1(n7044), 
        .B2(n6995), .ZN(n6969) );
  OAI211_X1 U7518 ( .C1(n7049), .C2(n6981), .A(n6970), .B(n6969), .ZN(U3098)
         );
  AOI22_X1 U7519 ( .A1(n6994), .A2(n7051), .B1(n6993), .B2(n7050), .ZN(n6973)
         );
  AOI22_X1 U7520 ( .A1(INSTQUEUE_REG_8__6__SCAN_IN), .A2(n7053), .B1(n6989), 
        .B2(n6971), .ZN(n6972) );
  OAI211_X1 U7521 ( .C1(n6992), .C2(n6974), .A(n6973), .B(n6972), .ZN(U3090)
         );
  AOI22_X1 U7522 ( .A1(n6993), .A2(n7056), .B1(n6989), .B2(n7065), .ZN(n6976)
         );
  AOI22_X1 U7523 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n7058), .B1(n6994), 
        .B2(n7057), .ZN(n6975) );
  OAI211_X1 U7524 ( .C1(n6992), .C2(n7061), .A(n6976), .B(n6975), .ZN(U3082)
         );
  AOI22_X1 U7525 ( .A1(n6994), .A2(n7064), .B1(n6993), .B2(n7063), .ZN(n6978)
         );
  AOI22_X1 U7526 ( .A1(INSTQUEUE_REG_6__6__SCAN_IN), .A2(n7066), .B1(n6995), 
        .B2(n7065), .ZN(n6977) );
  OAI211_X1 U7527 ( .C1(n6998), .C2(n7069), .A(n6978), .B(n6977), .ZN(U3074)
         );
  AOI22_X1 U7528 ( .A1(n6993), .A2(n7071), .B1(n6995), .B2(n7072), .ZN(n6980)
         );
  AOI22_X1 U7529 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n7073), .B1(n6989), 
        .B2(n7080), .ZN(n6979) );
  OAI211_X1 U7530 ( .C1(n7077), .C2(n6981), .A(n6980), .B(n6979), .ZN(U3066)
         );
  AOI22_X1 U7531 ( .A1(n6994), .A2(n7079), .B1(n6993), .B2(n7078), .ZN(n6983)
         );
  AOI22_X1 U7532 ( .A1(INSTQUEUE_REG_4__6__SCAN_IN), .A2(n7081), .B1(n6989), 
        .B2(n7085), .ZN(n6982) );
  OAI211_X1 U7533 ( .C1(n6992), .C2(n6984), .A(n6983), .B(n6982), .ZN(U3058)
         );
  AOI22_X1 U7534 ( .A1(n6993), .A2(n7086), .B1(n7094), .B2(n6989), .ZN(n6986)
         );
  AOI22_X1 U7535 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n7088), .B1(n6994), 
        .B2(n7087), .ZN(n6985) );
  OAI211_X1 U7536 ( .C1(n6992), .C2(n7084), .A(n6986), .B(n6985), .ZN(U3050)
         );
  AOI22_X1 U7537 ( .A1(n6994), .A2(n7093), .B1(n6993), .B2(n7092), .ZN(n6988)
         );
  AOI22_X1 U7538 ( .A1(INSTQUEUE_REG_2__6__SCAN_IN), .A2(n7095), .B1(n7101), 
        .B2(n6989), .ZN(n6987) );
  OAI211_X1 U7539 ( .C1(n7091), .C2(n6992), .A(n6988), .B(n6987), .ZN(U3042)
         );
  AOI22_X1 U7540 ( .A1(n6994), .A2(n7100), .B1(n6993), .B2(n7099), .ZN(n6991)
         );
  AOI22_X1 U7541 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n7102), .B1(n7111), 
        .B2(n6989), .ZN(n6990) );
  OAI211_X1 U7542 ( .C1(n7098), .C2(n6992), .A(n6991), .B(n6990), .ZN(U3034)
         );
  AOI22_X1 U7543 ( .A1(n6994), .A2(n7108), .B1(n6993), .B2(n7106), .ZN(n6997)
         );
  AOI22_X1 U7544 ( .A1(INSTQUEUE_REG_0__6__SCAN_IN), .A2(n7112), .B1(n7111), 
        .B2(n6995), .ZN(n6996) );
  OAI211_X1 U7545 ( .C1(n6998), .C2(n7115), .A(n6997), .B(n6996), .ZN(U3026)
         );
  AND2_X1 U7546 ( .A1(n5804), .A2(DATAI_31_), .ZN(n7070) );
  INV_X1 U7547 ( .A(n7070), .ZN(n7116) );
  NAND2_X1 U7548 ( .A1(DATAI_7_), .A2(n6999), .ZN(n7076) );
  NOR2_X2 U7549 ( .A1(n7001), .A2(n7000), .ZN(n7107) );
  AOI22_X1 U7550 ( .A1(n7109), .A2(n7003), .B1(n7107), .B2(n7002), .ZN(n7009)
         );
  NOR2_X2 U7551 ( .A1(n7005), .A2(n7004), .ZN(n7110) );
  AOI22_X1 U7552 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n7007), .B1(n7110), 
        .B2(n7006), .ZN(n7008) );
  OAI211_X1 U7553 ( .C1(n7116), .C2(n7010), .A(n7009), .B(n7008), .ZN(U3147)
         );
  AOI22_X1 U7554 ( .A1(n7109), .A2(n7012), .B1(n7107), .B2(n7011), .ZN(n7016)
         );
  AOI22_X1 U7555 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n7014), .B1(n7110), 
        .B2(n7013), .ZN(n7015) );
  OAI211_X1 U7556 ( .C1(n7116), .C2(n7017), .A(n7016), .B(n7015), .ZN(U3139)
         );
  AOI22_X1 U7557 ( .A1(n7107), .A2(n7019), .B1(n7018), .B2(n7110), .ZN(n7023)
         );
  AOI22_X1 U7558 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n7021), .B1(n7109), 
        .B2(n7020), .ZN(n7022) );
  OAI211_X1 U7559 ( .C1(n7116), .C2(n7024), .A(n7023), .B(n7022), .ZN(U3131)
         );
  AOI22_X1 U7560 ( .A1(n7109), .A2(n7026), .B1(n7107), .B2(n7025), .ZN(n7030)
         );
  AOI22_X1 U7561 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(n7028), .B1(n7110), 
        .B2(n7027), .ZN(n7029) );
  OAI211_X1 U7562 ( .C1(n7116), .C2(n7031), .A(n7030), .B(n7029), .ZN(U3123)
         );
  AOI22_X1 U7563 ( .A1(n7107), .A2(n7032), .B1(n7039), .B2(n7070), .ZN(n7036)
         );
  AOI22_X1 U7564 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n7034), .B1(n7110), 
        .B2(n7033), .ZN(n7035) );
  OAI211_X1 U7565 ( .C1(n7037), .C2(n7076), .A(n7036), .B(n7035), .ZN(U3115)
         );
  AOI22_X1 U7566 ( .A1(n7107), .A2(n7038), .B1(n7044), .B2(n7070), .ZN(n7042)
         );
  AOI22_X1 U7567 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n7040), .B1(n7039), 
        .B2(n7110), .ZN(n7041) );
  OAI211_X1 U7568 ( .C1(n7043), .C2(n7076), .A(n7042), .B(n7041), .ZN(U3107)
         );
  AOI22_X1 U7569 ( .A1(n7107), .A2(n7045), .B1(n7044), .B2(n7110), .ZN(n7048)
         );
  AOI22_X1 U7570 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n7046), .B1(n7070), 
        .B2(n7052), .ZN(n7047) );
  OAI211_X1 U7571 ( .C1(n7049), .C2(n7076), .A(n7048), .B(n7047), .ZN(U3099)
         );
  AOI22_X1 U7572 ( .A1(n7109), .A2(n7051), .B1(n7107), .B2(n7050), .ZN(n7055)
         );
  AOI22_X1 U7573 ( .A1(INSTQUEUE_REG_8__7__SCAN_IN), .A2(n7053), .B1(n7110), 
        .B2(n7052), .ZN(n7054) );
  OAI211_X1 U7574 ( .C1(n7116), .C2(n7061), .A(n7055), .B(n7054), .ZN(U3091)
         );
  INV_X1 U7575 ( .A(n7110), .ZN(n7062) );
  AOI22_X1 U7576 ( .A1(n7107), .A2(n7056), .B1(n7065), .B2(n7070), .ZN(n7060)
         );
  AOI22_X1 U7577 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n7058), .B1(n7109), 
        .B2(n7057), .ZN(n7059) );
  OAI211_X1 U7578 ( .C1(n7062), .C2(n7061), .A(n7060), .B(n7059), .ZN(U3083)
         );
  AOI22_X1 U7579 ( .A1(n7109), .A2(n7064), .B1(n7107), .B2(n7063), .ZN(n7068)
         );
  AOI22_X1 U7580 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(n7066), .B1(n7110), 
        .B2(n7065), .ZN(n7067) );
  OAI211_X1 U7581 ( .C1(n7116), .C2(n7069), .A(n7068), .B(n7067), .ZN(U3075)
         );
  AOI22_X1 U7582 ( .A1(n7107), .A2(n7071), .B1(n7070), .B2(n7080), .ZN(n7075)
         );
  AOI22_X1 U7583 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n7073), .B1(n7110), 
        .B2(n7072), .ZN(n7074) );
  OAI211_X1 U7584 ( .C1(n7077), .C2(n7076), .A(n7075), .B(n7074), .ZN(U3067)
         );
  AOI22_X1 U7585 ( .A1(n7109), .A2(n7079), .B1(n7107), .B2(n7078), .ZN(n7083)
         );
  AOI22_X1 U7586 ( .A1(INSTQUEUE_REG_4__7__SCAN_IN), .A2(n7081), .B1(n7110), 
        .B2(n7080), .ZN(n7082) );
  OAI211_X1 U7587 ( .C1(n7116), .C2(n7084), .A(n7083), .B(n7082), .ZN(U3059)
         );
  AOI22_X1 U7588 ( .A1(n7107), .A2(n7086), .B1(n7110), .B2(n7085), .ZN(n7090)
         );
  AOI22_X1 U7589 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n7088), .B1(n7109), 
        .B2(n7087), .ZN(n7089) );
  OAI211_X1 U7590 ( .C1(n7091), .C2(n7116), .A(n7090), .B(n7089), .ZN(U3051)
         );
  AOI22_X1 U7591 ( .A1(n7109), .A2(n7093), .B1(n7107), .B2(n7092), .ZN(n7097)
         );
  AOI22_X1 U7592 ( .A1(INSTQUEUE_REG_2__7__SCAN_IN), .A2(n7095), .B1(n7094), 
        .B2(n7110), .ZN(n7096) );
  OAI211_X1 U7593 ( .C1(n7098), .C2(n7116), .A(n7097), .B(n7096), .ZN(U3043)
         );
  AOI22_X1 U7594 ( .A1(n7109), .A2(n7100), .B1(n7107), .B2(n7099), .ZN(n7104)
         );
  AOI22_X1 U7595 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n7102), .B1(n7101), 
        .B2(n7110), .ZN(n7103) );
  OAI211_X1 U7596 ( .C1(n7105), .C2(n7116), .A(n7104), .B(n7103), .ZN(U3035)
         );
  AOI22_X1 U7597 ( .A1(n7109), .A2(n7108), .B1(n7107), .B2(n7106), .ZN(n7114)
         );
  AOI22_X1 U7598 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n7112), .B1(n7111), 
        .B2(n7110), .ZN(n7113) );
  OAI211_X1 U7599 ( .C1(n7116), .C2(n7115), .A(n7114), .B(n7113), .ZN(U3027)
         );
  AND2_X2 U3997 ( .A1(n3487), .A2(n4592), .ZN(n4229) );
  BUF_X2 U3540 ( .A(n3622), .Z(n5037) );
  AND4_X1 U3977 ( .A1(n3473), .A2(n3472), .A3(n3471), .A4(n3470), .ZN(n3495)
         );
  CLKBUF_X2 U3477 ( .A(n3897), .Z(n5086) );
  NOR2_X2 U3967 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3487) );
  NAND2_X2 U3597 ( .A1(n3448), .A2(n3925), .ZN(n3820) );
  CLKBUF_X3 U3580 ( .A(n3820), .Z(n3451) );
  CLKBUF_X1 U34680 ( .A(n3637), .Z(n3651) );
  CLKBUF_X1 U3482 ( .A(n3938), .Z(n3939) );
  AND2_X1 U3544 ( .A1(n3485), .A2(n4592), .ZN(n3897) );
  CLKBUF_X1 U3634 ( .A(n4820), .Z(n4857) );
  CLKBUF_X1 U3695 ( .A(n4593), .Z(n6630) );
endmodule

