

module b14_C_AntiSAT_k_256_2 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4989, n4990, n4991, n4992;

  CLKBUF_X2 U2463 ( .A(n2502), .Z(n2222) );
  AND2_X1 U2464 ( .A1(n2466), .A2(n2468), .ZN(n2492) );
  NAND2_X1 U2465 ( .A1(n3336), .A2(IR_REG_31__SCAN_IN), .ZN(n2462) );
  NOR2_X1 U2466 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2488)
         );
  NAND2_X1 U2467 ( .A1(n2771), .A2(n2821), .ZN(n2973) );
  INV_X2 U2468 ( .A(n3443), .ZN(n3511) );
  NAND2_X1 U2469 ( .A1(n4283), .A2(n2468), .ZN(n2502) );
  INV_X1 U2470 ( .A(IR_REG_31__SCAN_IN), .ZN(n2794) );
  AND4_X1 U2471 ( .A1(n2514), .A2(n2513), .A3(n2512), .A4(n2511), .ZN(n3067)
         );
  AND2_X1 U2472 ( .A1(n4544), .A2(n2821), .ZN(n4585) );
  INV_X2 U2473 ( .A(n4519), .ZN(n4337) );
  NOR2_X2 U2474 ( .A1(n4064), .A2(n4052), .ZN(n4048) );
  XNOR2_X2 U2475 ( .A(n2745), .B(n2744), .ZN(n2821) );
  INV_X2 U2476 ( .A(n2835), .ZN(n2499) );
  AOI22_X2 U2477 ( .A1(n3166), .A2(n2570), .B1(n3268), .B2(n3820), .ZN(n3241)
         );
  MUX2_X1 U2478 ( .A(REG1_REG_28__SCAN_IN), .B(n2825), .S(n4610), .Z(n2819) );
  MUX2_X1 U2479 ( .A(REG0_REG_28__SCAN_IN), .B(n2825), .S(n4596), .Z(n2826) );
  NAND2_X1 U2480 ( .A1(n3389), .A2(n3388), .ZN(n4322) );
  NAND2_X1 U2481 ( .A1(n2381), .A2(n2379), .ZN(n3386) );
  NAND2_X1 U2482 ( .A1(n3223), .A2(n3222), .ZN(n3259) );
  NOR3_X2 U2483 ( .A1(n4502), .A2(n2270), .A3(n3278), .ZN(n3329) );
  NAND2_X1 U2484 ( .A1(n3091), .A2(n3069), .ZN(n2526) );
  INV_X1 U2485 ( .A(n3033), .ZN(n3455) );
  INV_X1 U2486 ( .A(n3199), .ZN(n3044) );
  AND4_X1 U2487 ( .A1(n2534), .A2(n2533), .A3(n2532), .A4(n2531), .ZN(n3199)
         );
  INV_X2 U2488 ( .A(n2975), .ZN(n3509) );
  NAND2_X2 U2489 ( .A1(n2809), .A2(n2808), .ZN(n2950) );
  INV_X1 U2490 ( .A(n2491), .ZN(n2979) );
  INV_X1 U2491 ( .A(n4545), .ZN(n3011) );
  INV_X1 U2492 ( .A(n3090), .ZN(n3098) );
  NAND2_X1 U2493 ( .A1(n2743), .A2(IR_REG_31__SCAN_IN), .ZN(n2745) );
  INV_X1 U2494 ( .A(n2779), .ZN(n2771) );
  XNOR2_X1 U2495 ( .A(n2742), .B(n2741), .ZN(n3905) );
  NAND2_X1 U2496 ( .A1(n2464), .A2(IR_REG_31__SCAN_IN), .ZN(n2465) );
  XNOR2_X1 U2497 ( .A(n2795), .B(IR_REG_26__SCAN_IN), .ZN(n2859) );
  NAND2_X1 U2498 ( .A1(n2736), .A2(IR_REG_31__SCAN_IN), .ZN(n2742) );
  OR2_X1 U2499 ( .A1(n2646), .A2(n2239), .ZN(n2389) );
  NOR3_X1 U2500 ( .A1(n2432), .A2(n2235), .A3(n2431), .ZN(n2430) );
  AND2_X1 U2501 ( .A1(n2427), .A2(n2384), .ZN(n2451) );
  AND2_X1 U2502 ( .A1(n2474), .A2(n2386), .ZN(n2384) );
  AND2_X1 U2503 ( .A1(n2429), .A2(n2428), .ZN(n2427) );
  AND2_X1 U2504 ( .A1(n2385), .A2(n2428), .ZN(n2291) );
  NAND2_X1 U2505 ( .A1(n2263), .A2(n2262), .ZN(n2432) );
  AND2_X1 U2506 ( .A1(n2385), .A2(n2265), .ZN(n2264) );
  AND3_X1 U2507 ( .A1(n2438), .A2(n2488), .A3(n2399), .ZN(n2474) );
  AND2_X1 U2508 ( .A1(n2386), .A2(n2450), .ZN(n2385) );
  AND2_X1 U2509 ( .A1(n2567), .A2(n2444), .ZN(n2445) );
  AND2_X1 U2510 ( .A1(n2443), .A2(n2448), .ZN(n2386) );
  AND2_X1 U2511 ( .A1(n4793), .A2(n2523), .ZN(n2438) );
  NOR2_X1 U2512 ( .A1(n2437), .A2(IR_REG_18__SCAN_IN), .ZN(n2388) );
  NOR2_X1 U2513 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2450)
         );
  NOR2_X1 U2514 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2453)
         );
  NOR2_X1 U2515 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2452)
         );
  INV_X1 U2516 ( .A(IR_REG_25__SCAN_IN), .ZN(n2262) );
  NOR2_X1 U2517 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2567)
         );
  XNOR2_X2 U2519 ( .A(n2792), .B(IR_REG_24__SCAN_IN), .ZN(n2809) );
  OAI21_X2 U2520 ( .B1(n4084), .B2(n3735), .A(n3734), .ZN(n4067) );
  NAND2_X2 U2521 ( .A1(n4112), .A2(n2660), .ZN(n4084) );
  AOI21_X2 U2522 ( .B1(n3988), .B2(n2706), .A(n2705), .ZN(n3966) );
  OAI21_X2 U2523 ( .B1(n4010), .B2(n3729), .A(n3730), .ZN(n3988) );
  NAND2_X1 U2524 ( .A1(n2460), .A2(n2459), .ZN(n2223) );
  NAND2_X1 U2525 ( .A1(n2460), .A2(n2459), .ZN(n2224) );
  NOR2_X2 U2526 ( .A1(n3478), .A2(n2367), .ZN(n2364) );
  NOR2_X2 U2527 ( .A1(n3479), .A2(n3436), .ZN(n3478) );
  AOI21_X2 U2528 ( .B1(n3277), .B2(n2608), .A(n2607), .ZN(n3291) );
  AOI21_X2 U2529 ( .B1(n4487), .B2(n4489), .A(n2435), .ZN(n3277) );
  AOI21_X2 U2530 ( .B1(n3118), .B2(n3757), .A(n2441), .ZN(n3157) );
  OAI211_X2 U2531 ( .C1(n2403), .C2(n2405), .A(n2538), .B(n2401), .ZN(n3118)
         );
  OAI22_X2 U2532 ( .A1(n3087), .A2(n2516), .B1(n3067), .B2(n3098), .ZN(n3042)
         );
  NOR2_X1 U2533 ( .A1(n4283), .A2(n2468), .ZN(n2501) );
  XNOR2_X2 U2534 ( .A(n2465), .B(IR_REG_29__SCAN_IN), .ZN(n2468) );
  INV_X1 U2535 ( .A(n3702), .ZN(n2306) );
  OR2_X1 U2536 ( .A1(n4397), .A2(n2886), .ZN(n2887) );
  INV_X1 U2537 ( .A(IR_REG_13__SCAN_IN), .ZN(n2428) );
  NOR2_X1 U2538 ( .A1(n2629), .A2(n2397), .ZN(n2396) );
  INV_X1 U2539 ( .A(n2398), .ZN(n2397) );
  NAND2_X1 U2540 ( .A1(n3738), .A2(n3737), .ZN(n2421) );
  INV_X1 U2541 ( .A(n2456), .ZN(n2263) );
  OAI21_X1 U2542 ( .B1(n3635), .B2(n3631), .A(n3632), .ZN(n3501) );
  NAND2_X1 U2543 ( .A1(n2344), .A2(n2917), .ZN(n2342) );
  INV_X1 U2544 ( .A(n2887), .ZN(n2344) );
  NAND2_X1 U2545 ( .A1(n2383), .A2(n3469), .ZN(n2382) );
  NAND2_X1 U2546 ( .A1(n3130), .A2(n2378), .ZN(n2377) );
  INV_X1 U2547 ( .A(n3107), .ZN(n2378) );
  NAND2_X1 U2548 ( .A1(n2370), .A2(n2368), .ZN(n2367) );
  NAND2_X1 U2549 ( .A1(n3441), .A2(n2369), .ZN(n2368) );
  INV_X1 U2550 ( .A(n3576), .ZN(n2369) );
  NAND2_X1 U2551 ( .A1(n3844), .A2(n2899), .ZN(n2900) );
  NOR2_X1 U2552 ( .A1(n4448), .A2(n2352), .ZN(n3881) );
  AND2_X1 U2553 ( .A1(n4457), .A2(REG1_REG_15__SCAN_IN), .ZN(n2352) );
  NAND2_X1 U2554 ( .A1(n3931), .A2(n2281), .ZN(n2280) );
  NAND2_X1 U2555 ( .A1(n2284), .A2(n3714), .ZN(n2282) );
  NOR2_X1 U2556 ( .A1(n3773), .A2(n2285), .ZN(n2281) );
  NAND2_X1 U2557 ( .A1(n2290), .A2(n2287), .ZN(n2286) );
  INV_X1 U2558 ( .A(n3798), .ZN(n2287) );
  NOR2_X1 U2559 ( .A1(n3744), .A2(n2289), .ZN(n2288) );
  NAND2_X1 U2560 ( .A1(n2274), .A2(n2273), .ZN(n2769) );
  AND2_X1 U2561 ( .A1(n3789), .A2(n3709), .ZN(n2273) );
  NOR2_X1 U2562 ( .A1(n4123), .A2(n3733), .ZN(n4086) );
  AND2_X1 U2563 ( .A1(n2306), .A2(n3701), .ZN(n2300) );
  NAND2_X1 U2564 ( .A1(n2251), .A2(n2306), .ZN(n2303) );
  AND2_X1 U2565 ( .A1(n3695), .A2(n3701), .ZN(n2305) );
  NAND2_X1 U2566 ( .A1(n4488), .A2(n2300), .ZN(n2302) );
  OR2_X1 U2567 ( .A1(n3136), .A2(n3197), .ZN(n2407) );
  AOI21_X1 U2568 ( .B1(n2419), .B2(n2417), .A(n2416), .ZN(n2415) );
  INV_X1 U2569 ( .A(n2422), .ZN(n2417) );
  INV_X1 U2570 ( .A(n3919), .ZN(n2416) );
  NAND2_X1 U2571 ( .A1(n4142), .A2(n4124), .ZN(n2648) );
  NAND2_X1 U2572 ( .A1(n2537), .A2(n2526), .ZN(n2402) );
  INV_X1 U2573 ( .A(n2230), .ZN(n2405) );
  AND2_X1 U2574 ( .A1(n2796), .A2(n2859), .ZN(n2845) );
  INV_X1 U2575 ( .A(IR_REG_2__SCAN_IN), .ZN(n2442) );
  INV_X1 U2576 ( .A(IR_REG_1__SCAN_IN), .ZN(n2330) );
  NAND2_X1 U2577 ( .A1(n2360), .A2(n2249), .ZN(n2359) );
  NAND2_X1 U2578 ( .A1(n2361), .A2(n3641), .ZN(n2360) );
  INV_X1 U2579 ( .A(n2367), .ZN(n2355) );
  NAND2_X1 U2580 ( .A1(n2249), .A2(n2363), .ZN(n2362) );
  NAND2_X1 U2581 ( .A1(n3501), .A2(n3502), .ZN(n3500) );
  NAND2_X1 U2582 ( .A1(n3413), .A2(n3412), .ZN(n3414) );
  INV_X1 U2583 ( .A(n3410), .ZN(n3413) );
  NAND2_X1 U2584 ( .A1(n3393), .A2(n3395), .ZN(n3396) );
  INV_X1 U2585 ( .A(n3442), .ZN(n2370) );
  NOR2_X1 U2586 ( .A1(n2242), .A2(n2226), .ZN(n2363) );
  NAND2_X1 U2587 ( .A1(n2942), .A2(n3905), .ZN(n2974) );
  AND2_X1 U2588 ( .A1(n2861), .A2(n2859), .ZN(n2808) );
  AOI21_X1 U2589 ( .B1(n3651), .B2(REG2_REG_2__SCAN_IN), .A(n2426), .ZN(n2425)
         );
  NAND2_X1 U2590 ( .A1(n4285), .A2(REG1_REG_2__SCAN_IN), .ZN(n2336) );
  NAND2_X1 U2591 ( .A1(n3850), .A2(n2873), .ZN(n2875) );
  NAND2_X1 U2592 ( .A1(n4293), .A2(REG2_REG_3__SCAN_IN), .ZN(n4292) );
  NAND2_X1 U2593 ( .A1(n4371), .A2(n2907), .ZN(n4381) );
  NAND2_X1 U2594 ( .A1(n4381), .A2(n4382), .ZN(n4380) );
  NAND2_X1 U2595 ( .A1(n2341), .A2(n2339), .ZN(n4407) );
  NAND2_X1 U2596 ( .A1(n3874), .A2(n2343), .ZN(n2341) );
  NOR2_X1 U2597 ( .A1(n4408), .A2(n4832), .ZN(n2340) );
  OAI21_X1 U2598 ( .B1(n4434), .B2(n4432), .A(n2257), .ZN(n3864) );
  XNOR2_X1 U2599 ( .A(n3881), .B(n2332), .ZN(n4467) );
  NAND2_X1 U2600 ( .A1(n4467), .A2(n4855), .ZN(n4466) );
  NOR2_X1 U2601 ( .A1(n4452), .A2(n2333), .ZN(n3867) );
  AND2_X1 U2602 ( .A1(n4457), .A2(REG2_REG_15__SCAN_IN), .ZN(n2333) );
  NOR2_X1 U2603 ( .A1(n2729), .A2(n2423), .ZN(n2422) );
  INV_X1 U2604 ( .A(n3738), .ZN(n2423) );
  AND2_X1 U2605 ( .A1(n3739), .A2(n3738), .ZN(n3949) );
  AND4_X1 U2606 ( .A1(n2728), .A2(n2727), .A3(n2726), .A4(n2725), .ZN(n3952)
         );
  AOI21_X1 U2607 ( .B1(n2396), .B2(n2394), .A(n2250), .ZN(n2393) );
  INV_X1 U2608 ( .A(n2396), .ZN(n2395) );
  NAND2_X1 U2609 ( .A1(n4989), .A2(n3472), .ZN(n2398) );
  INV_X1 U2610 ( .A(n3322), .ZN(n3763) );
  NAND2_X1 U2611 ( .A1(n3376), .A2(n2618), .ZN(n2619) );
  OR2_X1 U2612 ( .A1(n2561), .A2(n2560), .ZN(n2571) );
  NAND2_X1 U2613 ( .A1(n2936), .A2(n4287), .ZN(n4491) );
  NAND2_X1 U2614 ( .A1(n2950), .A2(n4522), .ZN(n2956) );
  AND2_X1 U2615 ( .A1(n2780), .A2(n2779), .ZN(n4544) );
  INV_X1 U2616 ( .A(n2450), .ZN(n2431) );
  INV_X1 U2617 ( .A(n2432), .ZN(n2261) );
  INV_X1 U2618 ( .A(IR_REG_23__SCAN_IN), .ZN(n2811) );
  XNOR2_X1 U2619 ( .A(n2810), .B(n2811), .ZN(n3026) );
  NAND2_X1 U2620 ( .A1(n2668), .A2(n2667), .ZN(n2736) );
  INV_X1 U2621 ( .A(IR_REG_19__SCAN_IN), .ZN(n2741) );
  INV_X1 U2622 ( .A(n2488), .ZN(n2489) );
  INV_X1 U2623 ( .A(n4318), .ZN(n3638) );
  AND3_X1 U2624 ( .A1(n2342), .A2(n3872), .A3(REG1_REG_10__SCAN_IN), .ZN(n3873) );
  AND2_X1 U2625 ( .A1(n2546), .A2(n2427), .ZN(n2449) );
  XNOR2_X1 U2626 ( .A(n3864), .B(n4529), .ZN(n4441) );
  NOR2_X1 U2627 ( .A1(n4441), .A2(n3318), .ZN(n4440) );
  XNOR2_X1 U2628 ( .A(n3867), .B(n2332), .ZN(n4465) );
  NAND2_X1 U2629 ( .A1(n4465), .A2(n4464), .ZN(n4463) );
  INV_X1 U2630 ( .A(n2668), .ZN(n2656) );
  AND2_X1 U2631 ( .A1(n4341), .A2(n3837), .ZN(n4483) );
  AOI21_X1 U2632 ( .B1(n3885), .B2(n3884), .A(n4447), .ZN(n3890) );
  AND2_X1 U2633 ( .A1(n2818), .A2(n2817), .ZN(n2866) );
  INV_X1 U2634 ( .A(n2286), .ZN(n2285) );
  NAND2_X1 U2635 ( .A1(n4086), .A2(n2241), .ZN(n2274) );
  NOR2_X1 U2636 ( .A1(n2753), .A2(n2314), .ZN(n2313) );
  INV_X1 U2637 ( .A(n3667), .ZN(n2314) );
  NAND2_X1 U2638 ( .A1(n3468), .A2(n2380), .ZN(n2379) );
  NAND2_X1 U2639 ( .A1(n3467), .A2(n2382), .ZN(n2381) );
  INV_X1 U2640 ( .A(n3469), .ZN(n2380) );
  NAND2_X1 U2641 ( .A1(n4357), .A2(n2244), .ZN(n2906) );
  AOI21_X1 U2642 ( .B1(REG1_REG_11__SCAN_IN), .B2(n3875), .A(n4407), .ZN(n3876) );
  INV_X1 U2643 ( .A(n2327), .ZN(n2324) );
  AND2_X1 U2644 ( .A1(n3364), .A2(n4503), .ZN(n3695) );
  AND3_X1 U2645 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2477) );
  INV_X1 U2646 ( .A(n2313), .ZN(n2308) );
  AOI21_X1 U2647 ( .B1(n2312), .B2(n2313), .A(n2311), .ZN(n2310) );
  INV_X1 U2648 ( .A(n3670), .ZN(n2311) );
  NAND2_X1 U2649 ( .A1(n3206), .A2(n2266), .ZN(n3171) );
  AND2_X1 U2650 ( .A1(n2267), .A2(n3256), .ZN(n2266) );
  NOR2_X1 U2651 ( .A1(n3232), .A2(n3190), .ZN(n2267) );
  AND2_X1 U2652 ( .A1(n2428), .A2(n2457), .ZN(n2265) );
  INV_X1 U2653 ( .A(IR_REG_11__SCAN_IN), .ZN(n2593) );
  INV_X1 U2654 ( .A(IR_REG_6__SCAN_IN), .ZN(n2443) );
  OAI22_X1 U2655 ( .A1(n4989), .A2(n3448), .B1(n3472), .B2(n3447), .ZN(n3469)
         );
  OAI22_X1 U2656 ( .A1(n3567), .A2(n3401), .B1(n3400), .B2(n3568), .ZN(n3635)
         );
  NAND2_X1 U2657 ( .A1(n2375), .A2(n2234), .ZN(n3178) );
  NAND2_X1 U2658 ( .A1(n3064), .A2(n2376), .ZN(n2375) );
  OR2_X1 U2659 ( .A1(n2890), .A2(IR_REG_27__SCAN_IN), .ZN(n2460) );
  INV_X1 U2660 ( .A(n3559), .ZN(n2361) );
  NAND2_X1 U2661 ( .A1(n3386), .A2(n3387), .ZN(n4323) );
  NAND2_X1 U2662 ( .A1(n2483), .A2(REG3_REG_0__SCAN_IN), .ZN(n2496) );
  NAND2_X1 U2663 ( .A1(n2898), .A2(n2897), .ZN(n3844) );
  XNOR2_X1 U2664 ( .A(n2900), .B(n2874), .ZN(n4293) );
  OAI22_X1 U2665 ( .A1(n4348), .A2(n2905), .B1(n2904), .B2(n2903), .ZN(n4358)
         );
  NAND2_X1 U2666 ( .A1(n4358), .A2(n4359), .ZN(n4357) );
  XNOR2_X1 U2667 ( .A(n2906), .B(n2880), .ZN(n4372) );
  NAND2_X1 U2668 ( .A1(n4363), .A2(n2233), .ZN(n2881) );
  NAND2_X1 U2669 ( .A1(n4380), .A2(n2908), .ZN(n2910) );
  XNOR2_X1 U2670 ( .A(n3876), .B(n4427), .ZN(n4418) );
  OAI21_X1 U2671 ( .B1(n4418), .B2(n2350), .A(n2349), .ZN(n4428) );
  NAND2_X1 U2672 ( .A1(n2351), .A2(REG1_REG_12__SCAN_IN), .ZN(n2350) );
  NAND2_X1 U2673 ( .A1(n3877), .A2(n2351), .ZN(n2349) );
  INV_X1 U2674 ( .A(n4429), .ZN(n2351) );
  NOR2_X1 U2675 ( .A1(n4418), .A2(n4419), .ZN(n4417) );
  NAND2_X1 U2676 ( .A1(n4412), .A2(n2315), .ZN(n3862) );
  NAND2_X1 U2677 ( .A1(n3875), .A2(REG2_REG_11__SCAN_IN), .ZN(n2315) );
  AOI21_X1 U2678 ( .B1(n3878), .B2(REG1_REG_13__SCAN_IN), .A(n4428), .ZN(n3879) );
  NAND2_X1 U2679 ( .A1(n4466), .A2(n3882), .ZN(n4478) );
  NOR2_X1 U2680 ( .A1(n2328), .A2(n3893), .ZN(n2327) );
  NAND2_X1 U2681 ( .A1(n2326), .A2(n2324), .ZN(n2321) );
  NAND2_X1 U2682 ( .A1(n3902), .A2(n2323), .ZN(n2322) );
  NAND2_X1 U2683 ( .A1(n3870), .A2(n2324), .ZN(n2323) );
  AND2_X1 U2684 ( .A1(n3713), .A2(DATAI_27_), .ZN(n3932) );
  AND2_X1 U2685 ( .A1(n2279), .A2(n2277), .ZN(n3929) );
  NAND2_X1 U2686 ( .A1(n2278), .A2(n3931), .ZN(n2277) );
  INV_X1 U2687 ( .A(n2282), .ZN(n2278) );
  NAND2_X1 U2688 ( .A1(n2275), .A2(n2282), .ZN(n3930) );
  OR2_X1 U2689 ( .A1(n3991), .A2(n2276), .ZN(n2275) );
  INV_X1 U2690 ( .A(n2281), .ZN(n2276) );
  NAND2_X1 U2691 ( .A1(n2283), .A2(n2286), .ZN(n3950) );
  NAND2_X1 U2692 ( .A1(n3991), .A2(n2288), .ZN(n2283) );
  OR2_X1 U2693 ( .A1(n2707), .A2(n3561), .ZN(n2723) );
  INV_X1 U2694 ( .A(n3979), .ZN(n3972) );
  NAND2_X1 U2695 ( .A1(n3991), .A2(n3787), .ZN(n3968) );
  AND2_X1 U2696 ( .A1(n2693), .A2(REG3_REG_23__SCAN_IN), .ZN(n2699) );
  NOR2_X1 U2697 ( .A1(n2686), .A2(n3612), .ZN(n2693) );
  AND2_X1 U2698 ( .A1(n3713), .A2(DATAI_22_), .ZN(n4041) );
  NOR2_X1 U2699 ( .A1(n2685), .A2(n2411), .ZN(n2410) );
  INV_X1 U2700 ( .A(n2677), .ZN(n2411) );
  NAND2_X1 U2701 ( .A1(n2409), .A2(n2408), .ZN(n4030) );
  AND2_X1 U2702 ( .A1(n2692), .A2(n2243), .ZN(n2408) );
  AND4_X1 U2703 ( .A1(n2691), .A2(n2690), .A3(n2689), .A4(n2688), .ZN(n4056)
         );
  INV_X1 U2704 ( .A(n3544), .ZN(n4052) );
  AND2_X1 U2705 ( .A1(n3728), .A2(n4015), .ZN(n4051) );
  NOR2_X1 U2706 ( .A1(n2661), .A2(n3504), .ZN(n2670) );
  AND2_X1 U2707 ( .A1(REG3_REG_17__SCAN_IN), .A2(n2650), .ZN(n2651) );
  OAI21_X1 U2708 ( .B1(n4141), .B2(n4153), .A(n2757), .ZN(n4123) );
  NAND2_X1 U2709 ( .A1(n2392), .A2(n2390), .ZN(n4152) );
  AOI21_X1 U2710 ( .B1(n2393), .B2(n2395), .A(n2391), .ZN(n2390) );
  NAND2_X1 U2711 ( .A1(n2298), .A2(n2297), .ZN(n3324) );
  NAND2_X1 U2712 ( .A1(n2301), .A2(n3698), .ZN(n2297) );
  NAND2_X1 U2713 ( .A1(n4488), .A2(n2247), .ZN(n2298) );
  AND2_X1 U2714 ( .A1(n2302), .A2(n2299), .ZN(n3312) );
  AND2_X1 U2715 ( .A1(n4494), .A2(n3278), .ZN(n2607) );
  AND2_X1 U2716 ( .A1(n2598), .A2(REG3_REG_12__SCAN_IN), .ZN(n2609) );
  AND2_X1 U2717 ( .A1(n2609), .A2(REG3_REG_13__SCAN_IN), .ZN(n2611) );
  NAND2_X1 U2718 ( .A1(n2304), .A2(n3701), .ZN(n3295) );
  OR2_X1 U2719 ( .A1(n4488), .A2(n3695), .ZN(n2304) );
  INV_X1 U2720 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2584) );
  INV_X1 U2721 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2914) );
  OR2_X1 U2722 ( .A1(n2571), .A2(n2914), .ZN(n2585) );
  NAND2_X1 U2723 ( .A1(n3136), .A2(n3197), .ZN(n2538) );
  OAI21_X1 U2724 ( .B1(n3089), .B2(n2308), .A(n2310), .ZN(n3019) );
  INV_X1 U2725 ( .A(n4491), .ZN(n4126) );
  NAND2_X1 U2726 ( .A1(n4555), .A2(n3098), .ZN(n3097) );
  OR2_X1 U2727 ( .A1(n3097), .A2(n3069), .ZN(n3049) );
  NAND2_X1 U2728 ( .A1(n3088), .A2(n3667), .ZN(n3043) );
  OAI21_X1 U2729 ( .B1(n2829), .B2(n2752), .A(n3662), .ZN(n3089) );
  NAND2_X1 U2730 ( .A1(n3089), .A2(n3760), .ZN(n3088) );
  INV_X1 U2731 ( .A(n2930), .ZN(n3093) );
  INV_X1 U2732 ( .A(n3005), .ZN(n2996) );
  INV_X1 U2733 ( .A(n3825), .ZN(n3078) );
  AND2_X1 U2734 ( .A1(n3825), .A2(n4545), .ZN(n3074) );
  NAND2_X1 U2735 ( .A1(n3759), .A2(n3074), .ZN(n3076) );
  INV_X1 U2736 ( .A(n4145), .ZN(n4497) );
  AND2_X1 U2737 ( .A1(n4544), .A2(n4284), .ZN(n4162) );
  AOI21_X1 U2738 ( .B1(n2415), .B2(n2420), .A(n2248), .ZN(n2413) );
  NAND2_X1 U2739 ( .A1(n3957), .A2(n3941), .ZN(n3940) );
  OR2_X1 U2740 ( .A1(n3940), .A2(n3921), .ZN(n3924) );
  AND2_X1 U2741 ( .A1(n3977), .A2(n3959), .ZN(n3957) );
  NOR2_X1 U2742 ( .A1(n4000), .A2(n3972), .ZN(n3977) );
  NAND2_X1 U2743 ( .A1(n2272), .A2(n4001), .ZN(n4000) );
  INV_X1 U2744 ( .A(n3484), .ZN(n4020) );
  OR2_X1 U2745 ( .A1(n4096), .A2(n4074), .ZN(n4064) );
  AND2_X1 U2746 ( .A1(n4131), .A2(n3405), .ZN(n4098) );
  NAND2_X1 U2747 ( .A1(n4098), .A2(n4097), .ZN(n4096) );
  OR2_X1 U2748 ( .A1(n4148), .A2(n4147), .ZN(n4150) );
  NOR2_X1 U2749 ( .A1(n4150), .A2(n4124), .ZN(n4131) );
  NAND2_X1 U2750 ( .A1(n3376), .A2(n3472), .ZN(n2270) );
  INV_X1 U2751 ( .A(n3551), .ZN(n3278) );
  NOR2_X1 U2752 ( .A1(n3171), .A2(n3496), .ZN(n4504) );
  NAND2_X1 U2753 ( .A1(n3206), .A2(n3181), .ZN(n3158) );
  NOR2_X1 U2754 ( .A1(n3049), .A2(n3114), .ZN(n3204) );
  AND2_X1 U2755 ( .A1(n3204), .A2(n3203), .ZN(n3206) );
  NAND2_X1 U2756 ( .A1(n2402), .A2(n2230), .ZN(n2404) );
  INV_X1 U2757 ( .A(n4577), .ZN(n4580) );
  OAI21_X1 U2758 ( .B1(n2224), .B2(n2498), .A(n2497), .ZN(n4545) );
  NAND2_X1 U2759 ( .A1(n2223), .A2(DATAI_0_), .ZN(n2497) );
  INV_X1 U2760 ( .A(n2845), .ZN(n2865) );
  INV_X1 U2761 ( .A(n2956), .ZN(n2945) );
  NAND2_X1 U2762 ( .A1(n2789), .A2(n2788), .ZN(n2814) );
  INV_X1 U2763 ( .A(n2787), .ZN(n2788) );
  INV_X1 U2764 ( .A(n2786), .ZN(n2789) );
  XNOR2_X1 U2765 ( .A(n2747), .B(n2746), .ZN(n2780) );
  NAND2_X1 U2766 ( .A1(n2790), .A2(IR_REG_31__SCAN_IN), .ZN(n2747) );
  NAND2_X1 U2767 ( .A1(n2740), .A2(n2790), .ZN(n2779) );
  MUX2_X1 U2768 ( .A(IR_REG_31__SCAN_IN), .B(n2737), .S(IR_REG_21__SCAN_IN), 
        .Z(n2740) );
  INV_X1 U2769 ( .A(IR_REG_20__SCAN_IN), .ZN(n2744) );
  XNOR2_X1 U2770 ( .A(n2647), .B(IR_REG_17__SCAN_IN), .ZN(n3883) );
  INV_X1 U2771 ( .A(IR_REG_16__SCAN_IN), .ZN(n4698) );
  INV_X1 U2772 ( .A(IR_REG_10__SCAN_IN), .ZN(n2579) );
  NOR2_X1 U2773 ( .A1(IR_REG_2__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2399)
         );
  INV_X1 U2774 ( .A(n2515), .ZN(n2400) );
  INV_X1 U2775 ( .A(IR_REG_3__SCAN_IN), .ZN(n4793) );
  INV_X1 U2776 ( .A(IR_REG_4__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U2777 ( .A1(n2237), .A2(IR_REG_0__SCAN_IN), .ZN(n2331) );
  NAND2_X1 U2778 ( .A1(n2330), .A2(n2794), .ZN(n2329) );
  INV_X1 U2779 ( .A(n3932), .ZN(n3941) );
  INV_X1 U2780 ( .A(n2353), .ZN(n3517) );
  INV_X1 U2781 ( .A(n2362), .ZN(n2356) );
  OAI21_X1 U2782 ( .B1(n2362), .B2(n2355), .A(n2359), .ZN(n2354) );
  AND4_X1 U2783 ( .A1(n2590), .A2(n2589), .A3(n2588), .A4(n2587), .ZN(n3552)
         );
  NAND2_X1 U2784 ( .A1(n3357), .A2(n3356), .ZN(n3490) );
  AND4_X1 U2785 ( .A1(n2566), .A2(n2565), .A3(n2564), .A4(n2563), .ZN(n3493)
         );
  INV_X1 U2786 ( .A(n3227), .ZN(n3232) );
  INV_X1 U2787 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3543) );
  NAND2_X1 U2788 ( .A1(n2371), .A2(n2372), .ZN(n3541) );
  INV_X1 U2789 ( .A(n2373), .ZN(n2372) );
  NAND2_X1 U2790 ( .A1(n3501), .A2(n2227), .ZN(n2371) );
  OAI21_X1 U2791 ( .B1(n3414), .B2(n2374), .A(n3586), .ZN(n2373) );
  NAND2_X1 U2792 ( .A1(n3108), .A2(n3107), .ZN(n3131) );
  NAND2_X1 U2793 ( .A1(n2370), .A2(n2366), .ZN(n2365) );
  INV_X1 U2794 ( .A(n3061), .ZN(n3069) );
  NAND2_X1 U2795 ( .A1(n3538), .A2(n3587), .ZN(n3584) );
  INV_X1 U2796 ( .A(n4041), .ZN(n4037) );
  OAI21_X1 U2797 ( .B1(n3541), .B2(n3535), .A(n3536), .ZN(n3610) );
  INV_X1 U2798 ( .A(n2596), .ZN(n4503) );
  OAI21_X1 U2799 ( .B1(n3713), .B2(n2507), .A(n2506), .ZN(n3005) );
  INV_X1 U2800 ( .A(n4285), .ZN(n2507) );
  NAND2_X1 U2801 ( .A1(n2223), .A2(DATAI_2_), .ZN(n2506) );
  AND4_X1 U2802 ( .A1(n2545), .A2(n2544), .A3(n2543), .A4(n2542), .ZN(n3230)
         );
  INV_X1 U2803 ( .A(n2357), .ZN(n3643) );
  OAI21_X1 U2804 ( .B1(n2364), .B2(n2358), .A(n2361), .ZN(n2357) );
  INV_X1 U2805 ( .A(n2363), .ZN(n2358) );
  INV_X1 U2806 ( .A(n4331), .ZN(n3648) );
  INV_X1 U2807 ( .A(n3326), .ZN(n4317) );
  AND2_X1 U2808 ( .A1(n2948), .A2(n4151), .ZN(n4318) );
  NOR2_X1 U2809 ( .A1(n3447), .A2(n2944), .ZN(n3811) );
  INV_X1 U2810 ( .A(n3230), .ZN(n3823) );
  OR2_X1 U2811 ( .A1(n2828), .A2(n2950), .ZN(n3822) );
  INV_X1 U2812 ( .A(n4522), .ZN(n2828) );
  CLKBUF_X1 U2813 ( .A(n2930), .Z(n2995) );
  AND2_X1 U2814 ( .A1(n2889), .A2(n2888), .ZN(n4341) );
  NAND2_X1 U2815 ( .A1(n3828), .A2(n3838), .ZN(n3843) );
  NAND2_X1 U2816 ( .A1(n2337), .A2(n2334), .ZN(n3850) );
  XNOR2_X1 U2817 ( .A(n2875), .B(n2874), .ZN(n4291) );
  NAND2_X1 U2818 ( .A1(n4364), .A2(n4365), .ZN(n4363) );
  XNOR2_X1 U2819 ( .A(n2881), .B(n2880), .ZN(n4370) );
  NAND2_X1 U2820 ( .A1(n4370), .A2(REG1_REG_6__SCAN_IN), .ZN(n4369) );
  XNOR2_X1 U2821 ( .A(n2910), .B(n4537), .ZN(n4394) );
  XNOR2_X1 U2822 ( .A(n2345), .B(n2909), .ZN(n4389) );
  NOR2_X1 U2823 ( .A1(n4389), .A2(n4390), .ZN(n4388) );
  OAI21_X1 U2824 ( .B1(n4389), .B2(n2347), .A(n2346), .ZN(n4397) );
  NAND2_X1 U2825 ( .A1(n2348), .A2(REG1_REG_8__SCAN_IN), .ZN(n2347) );
  NAND2_X1 U2826 ( .A1(n2884), .A2(n2348), .ZN(n2346) );
  INV_X1 U2827 ( .A(n4398), .ZN(n2348) );
  NAND2_X1 U2828 ( .A1(n2342), .A2(n3872), .ZN(n2891) );
  NAND2_X1 U2829 ( .A1(n3859), .A2(n3860), .ZN(n4413) );
  NAND2_X1 U2830 ( .A1(n4413), .A2(n4414), .ZN(n4412) );
  INV_X1 U2831 ( .A(n3873), .ZN(n2338) );
  XNOR2_X1 U2832 ( .A(n3862), .B(n4427), .ZN(n4424) );
  XNOR2_X1 U2833 ( .A(n2638), .B(IR_REG_15__SCAN_IN), .ZN(n4457) );
  NOR2_X1 U2834 ( .A1(n4440), .A2(n3865), .ZN(n4454) );
  AND2_X1 U2835 ( .A1(n4341), .A2(n2981), .ZN(n4458) );
  NAND2_X1 U2836 ( .A1(n4463), .A2(n3868), .ZN(n4475) );
  AND2_X1 U2837 ( .A1(n4341), .A2(n3833), .ZN(n4481) );
  NOR2_X1 U2838 ( .A1(n2326), .A2(n2327), .ZN(n2320) );
  NOR2_X1 U2839 ( .A1(n3906), .A2(n2229), .ZN(n2318) );
  NAND2_X1 U2840 ( .A1(n4483), .A2(n2258), .ZN(n2319) );
  INV_X1 U2841 ( .A(n3870), .ZN(n2325) );
  INV_X1 U2842 ( .A(n4481), .ZN(n4447) );
  NAND2_X1 U2843 ( .A1(n2296), .A2(n2294), .ZN(n4174) );
  XNOR2_X1 U2844 ( .A(n3924), .B(n3741), .ZN(n4175) );
  NAND2_X1 U2845 ( .A1(n2414), .A2(n2419), .ZN(n3920) );
  NAND2_X1 U2846 ( .A1(n2418), .A2(n3738), .ZN(n3938) );
  NAND2_X1 U2847 ( .A1(n4048), .A2(n4037), .ZN(n4194) );
  NAND2_X1 U2848 ( .A1(n3311), .A2(n2398), .ZN(n3323) );
  AND2_X1 U2850 ( .A1(n4337), .A2(n3018), .ZN(n4068) );
  AND2_X1 U2851 ( .A1(n2406), .A2(n2526), .ZN(n3016) );
  INV_X1 U2852 ( .A(n3905), .ZN(n3897) );
  NOR2_X1 U2853 ( .A1(n2849), .A2(n3005), .ZN(n4555) );
  OR2_X2 U2854 ( .A1(n2956), .A2(n2847), .ZN(n4151) );
  AND2_X2 U2855 ( .A1(n2823), .A2(n2935), .ZN(n4610) );
  NAND2_X1 U2856 ( .A1(n4165), .A2(n2269), .ZN(n4335) );
  OR2_X1 U2857 ( .A1(n4166), .A2(n4169), .ZN(n2269) );
  AND2_X2 U2858 ( .A1(n2824), .A2(n2823), .ZN(n4596) );
  XNOR2_X1 U2859 ( .A(n2774), .B(IR_REG_28__SCAN_IN), .ZN(n4287) );
  OR2_X1 U2860 ( .A1(n2787), .A2(n2794), .ZN(n2795) );
  NAND2_X1 U2861 ( .A1(n2791), .A2(IR_REG_31__SCAN_IN), .ZN(n2792) );
  AND2_X1 U2862 ( .A1(n3026), .A2(STATE_REG_SCAN_IN), .ZN(n4522) );
  INV_X1 U2863 ( .A(n3878), .ZN(n4530) );
  INV_X1 U2864 ( .A(DATAI_13_), .ZN(n4884) );
  INV_X1 U2865 ( .A(n2893), .ZN(n4542) );
  INV_X2 U2866 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  AOI21_X1 U2867 ( .B1(n3890), .B2(n3889), .A(n3888), .ZN(n3891) );
  OAI21_X1 U2868 ( .B1(n4335), .B2(n4135), .A(n2268), .ZN(U3261) );
  AOI22_X1 U2869 ( .A1(n4519), .A2(REG2_REG_30__SCAN_IN), .B1(n4337), .B2(
        n4336), .ZN(n2268) );
  INV_X1 U2870 ( .A(n2492), .ZN(n2510) );
  INV_X2 U2871 ( .A(n2510), .ZN(n2573) );
  AND2_X1 U2872 ( .A1(n4173), .A2(n4577), .ZN(n2225) );
  AND2_X1 U2873 ( .A1(n2409), .A2(n2243), .ZN(n4029) );
  INV_X1 U2874 ( .A(n3744), .ZN(n2290) );
  INV_X1 U2875 ( .A(n2420), .ZN(n2419) );
  OAI22_X1 U2876 ( .A1(n2729), .A2(n2421), .B1(n3941), .B2(n3952), .ZN(n2420)
         );
  NAND2_X1 U2877 ( .A1(n2400), .A2(n2438), .ZN(n2535) );
  AND2_X1 U2878 ( .A1(n2366), .A2(n3576), .ZN(n2226) );
  INV_X1 U2879 ( .A(n3762), .ZN(n2394) );
  AND2_X1 U2880 ( .A1(n3502), .A2(n3587), .ZN(n2227) );
  INV_X1 U2881 ( .A(n4408), .ZN(n2343) );
  AND4_X1 U2882 ( .A1(n2645), .A2(n2644), .A3(n2643), .A4(n2642), .ZN(n4300)
         );
  OR3_X1 U2883 ( .A1(n4502), .A2(n3278), .A3(n3606), .ZN(n2228) );
  INV_X1 U2884 ( .A(n3875), .ZN(n4534) );
  AND2_X1 U2885 ( .A1(n2595), .A2(n2604), .ZN(n3875) );
  AND2_X1 U2886 ( .A1(n4483), .A2(n2259), .ZN(n2229) );
  CLKBUF_X3 U2887 ( .A(n2501), .Z(n2720) );
  OR2_X1 U2888 ( .A1(n3044), .A2(n3114), .ZN(n2230) );
  AND2_X1 U2889 ( .A1(n2467), .A2(n4283), .ZN(n2231) );
  NOR2_X1 U2890 ( .A1(n2646), .A2(n2432), .ZN(n2787) );
  AND2_X1 U2891 ( .A1(n2474), .A2(n2443), .ZN(n2546) );
  NAND2_X1 U2892 ( .A1(n2678), .A2(n2677), .ZN(n4046) );
  OR2_X1 U2893 ( .A1(n3478), .A2(n2365), .ZN(n2232) );
  INV_X1 U2894 ( .A(n3190), .ZN(n3181) );
  OR2_X1 U2895 ( .A1(n4542), .A2(n4896), .ZN(n2233) );
  AND2_X1 U2896 ( .A1(n2377), .A2(n3135), .ZN(n2234) );
  OR2_X1 U2897 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2235)
         );
  NAND2_X1 U2898 ( .A1(n2236), .A2(n2489), .ZN(n2894) );
  INV_X1 U2899 ( .A(IR_REG_18__SCAN_IN), .ZN(n2667) );
  NAND2_X1 U2900 ( .A1(n2488), .A2(n2442), .ZN(n2515) );
  OAI21_X1 U2901 ( .B1(n2288), .B2(n2285), .A(n3656), .ZN(n2284) );
  NAND2_X1 U2902 ( .A1(n3500), .A2(n3414), .ZN(n3538) );
  AND2_X1 U2903 ( .A1(n2331), .A2(n2329), .ZN(n2236) );
  AND2_X1 U2904 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2237)
         );
  AND3_X1 U2905 ( .A1(n2446), .A2(n2579), .A3(n2593), .ZN(n2238) );
  INV_X1 U2906 ( .A(IR_REG_28__SCAN_IN), .ZN(n2463) );
  NAND2_X1 U2907 ( .A1(n2388), .A2(n2387), .ZN(n2239) );
  INV_X1 U2908 ( .A(n3787), .ZN(n2289) );
  NAND2_X1 U2909 ( .A1(n3044), .A2(n3110), .ZN(n2240) );
  NAND2_X1 U2910 ( .A1(n2546), .A2(n2445), .ZN(n2578) );
  OAI21_X1 U2911 ( .B1(n3549), .B2(n3383), .A(n3382), .ZN(n3467) );
  INV_X1 U2912 ( .A(n3317), .ZN(n3472) );
  AND2_X1 U2913 ( .A1(n4011), .A2(n4013), .ZN(n2241) );
  NOR2_X1 U2914 ( .A1(n3450), .A2(n3449), .ZN(n2242) );
  NAND2_X1 U2915 ( .A1(n3309), .A2(n3762), .ZN(n3311) );
  OR2_X1 U2916 ( .A1(n4075), .A2(n4052), .ZN(n2243) );
  INV_X1 U2917 ( .A(n3468), .ZN(n2383) );
  INV_X1 U2918 ( .A(n2909), .ZN(n4537) );
  OR2_X1 U2919 ( .A1(n4542), .A2(n4869), .ZN(n2244) );
  NOR2_X1 U2920 ( .A1(n4417), .A2(n3877), .ZN(n2245) );
  INV_X1 U2921 ( .A(n3587), .ZN(n2374) );
  INV_X1 U2922 ( .A(n2272), .ZN(n4009) );
  NOR2_X1 U2923 ( .A1(n4194), .A2(n4020), .ZN(n2272) );
  OR2_X1 U2924 ( .A1(n4056), .A2(n4037), .ZN(n2246) );
  AND2_X1 U2925 ( .A1(n2300), .A2(n3698), .ZN(n2247) );
  AND2_X1 U2926 ( .A1(n3933), .A2(n3921), .ZN(n2248) );
  NAND2_X1 U2927 ( .A1(n3459), .A2(n3458), .ZN(n2249) );
  INV_X1 U2928 ( .A(n2295), .ZN(n2294) );
  OAI21_X1 U2929 ( .B1(n3917), .B2(n4491), .A(n3916), .ZN(n2295) );
  NOR2_X1 U2930 ( .A1(n4299), .A2(n4317), .ZN(n2250) );
  INV_X1 U2931 ( .A(n2301), .ZN(n2299) );
  NAND2_X1 U2932 ( .A1(n2303), .A2(n2394), .ZN(n2301) );
  OR2_X1 U2933 ( .A1(n3700), .A2(n2305), .ZN(n2251) );
  OR2_X1 U2934 ( .A1(n4142), .A2(n4124), .ZN(n2252) );
  AND2_X1 U2935 ( .A1(n2546), .A2(n2429), .ZN(n2253) );
  OAI21_X1 U2936 ( .B1(n2790), .B2(IR_REG_22__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2810) );
  INV_X1 U2937 ( .A(n4153), .ZN(n2391) );
  NAND2_X1 U2938 ( .A1(n3206), .A2(n2267), .ZN(n2254) );
  AND2_X2 U2939 ( .A1(n2848), .A2(n4151), .ZN(n4519) );
  INV_X1 U2940 ( .A(n2780), .ZN(n2942) );
  AND2_X1 U2941 ( .A1(n4118), .A2(n4585), .ZN(n4513) );
  INV_X1 U2942 ( .A(n4303), .ZN(n4147) );
  AND2_X1 U2943 ( .A1(n3667), .A2(n3664), .ZN(n3760) );
  INV_X1 U2944 ( .A(n3760), .ZN(n2312) );
  NOR2_X1 U2945 ( .A1(n4388), .A2(n2884), .ZN(n2255) );
  INV_X1 U2946 ( .A(n2271), .ZN(n3302) );
  NOR2_X1 U2947 ( .A1(n4502), .A2(n3278), .ZN(n2271) );
  AND2_X1 U2948 ( .A1(n2338), .A2(n3872), .ZN(n2256) );
  INV_X1 U2949 ( .A(n4527), .ZN(n2332) );
  NAND2_X1 U2950 ( .A1(n2458), .A2(IR_REG_31__SCAN_IN), .ZN(n2890) );
  INV_X1 U2951 ( .A(n3741), .ZN(n3925) );
  OR2_X1 U2952 ( .A1(n3878), .A2(REG2_REG_13__SCAN_IN), .ZN(n2257) );
  INV_X1 U2953 ( .A(n4001), .ZN(n3995) );
  AND2_X1 U2954 ( .A1(n2325), .A2(n2326), .ZN(n2258) );
  AND2_X1 U2955 ( .A1(n2322), .A2(n2321), .ZN(n2259) );
  AND2_X1 U2956 ( .A1(n4483), .A2(n2320), .ZN(n2260) );
  INV_X1 U2957 ( .A(n3902), .ZN(n2326) );
  INV_X1 U2958 ( .A(IR_REG_12__SCAN_IN), .ZN(n2446) );
  INV_X1 U2959 ( .A(IR_REG_14__SCAN_IN), .ZN(n2448) );
  INV_X1 U2960 ( .A(IR_REG_17__SCAN_IN), .ZN(n2387) );
  INV_X1 U2961 ( .A(REG2_REG_18__SCAN_IN), .ZN(n2328) );
  NAND4_X1 U2962 ( .A1(n2264), .A2(n2261), .A3(n2474), .A4(n2429), .ZN(n2458)
         );
  AND2_X2 U2963 ( .A1(n2445), .A2(n2238), .ZN(n2429) );
  OR2_X1 U2965 ( .A1(n3991), .A2(n2280), .ZN(n2279) );
  NAND3_X1 U2966 ( .A1(n2429), .A2(n2474), .A3(n2291), .ZN(n2646) );
  NAND2_X1 U2967 ( .A1(n4175), .A2(n4585), .ZN(n2292) );
  NAND3_X1 U2968 ( .A1(n2296), .A2(n2293), .A3(n2292), .ZN(n4243) );
  NOR2_X2 U2969 ( .A1(n2225), .A2(n2295), .ZN(n2293) );
  NOR2_X1 U2970 ( .A1(n3924), .A2(n3925), .ZN(n4166) );
  NAND2_X1 U2971 ( .A1(n3914), .A2(n4145), .ZN(n2296) );
  NAND2_X1 U2972 ( .A1(n2302), .A2(n2303), .ZN(n3777) );
  NAND3_X1 U2973 ( .A1(n2309), .A2(n2307), .A3(n3684), .ZN(n3196) );
  NAND3_X1 U2974 ( .A1(n2240), .A2(n2310), .A3(n2308), .ZN(n2307) );
  NAND3_X1 U2975 ( .A1(n2240), .A2(n2310), .A3(n3089), .ZN(n2309) );
  NAND2_X1 U2976 ( .A1(n3869), .A2(n2260), .ZN(n2317) );
  INV_X1 U2977 ( .A(n2316), .ZN(n3907) );
  OAI211_X1 U2978 ( .C1(n3869), .C2(n2319), .A(n2318), .B(n2317), .ZN(n2316)
         );
  NOR2_X1 U2979 ( .A1(n3869), .A2(n3870), .ZN(n3900) );
  MUX2_X1 U2980 ( .A(n2895), .B(REG2_REG_1__SCAN_IN), .S(n2894), .Z(n3828) );
  NAND2_X1 U2981 ( .A1(n2489), .A2(IR_REG_31__SCAN_IN), .ZN(n2505) );
  INV_X1 U2982 ( .A(n2335), .ZN(n2334) );
  OAI21_X1 U2983 ( .B1(n4285), .B2(REG1_REG_2__SCAN_IN), .A(n2336), .ZN(n2335)
         );
  NAND2_X1 U2984 ( .A1(n3847), .A2(n3848), .ZN(n2337) );
  NAND3_X1 U2985 ( .A1(n2342), .A2(n3872), .A3(n2340), .ZN(n2339) );
  INV_X1 U2986 ( .A(n2883), .ZN(n2345) );
  NAND2_X4 U2987 ( .A1(n2950), .A2(n2973), .ZN(n3508) );
  AOI21_X1 U2988 ( .B1(n3478), .B2(n2356), .A(n2354), .ZN(n2353) );
  NOR2_X1 U2989 ( .A1(n2364), .A2(n2226), .ZN(n3558) );
  OAI21_X1 U2990 ( .B1(n3478), .B2(n3442), .A(n3441), .ZN(n3575) );
  INV_X1 U2991 ( .A(n3441), .ZN(n2366) );
  AND2_X1 U2992 ( .A1(n3063), .A2(n3130), .ZN(n2376) );
  NAND2_X1 U2993 ( .A1(n3064), .A2(n3063), .ZN(n3108) );
  INV_X1 U2994 ( .A(n2451), .ZN(n2628) );
  NOR2_X1 U2995 ( .A1(n2646), .A2(IR_REG_17__SCAN_IN), .ZN(n2668) );
  NAND2_X1 U2996 ( .A1(n2389), .A2(IR_REG_31__SCAN_IN), .ZN(n2737) );
  INV_X1 U2997 ( .A(n2389), .ZN(n2739) );
  NAND3_X1 U2998 ( .A1(n3261), .A2(n3263), .A3(n3260), .ZN(n3357) );
  NAND2_X1 U2999 ( .A1(n3261), .A2(n3260), .ZN(n3262) );
  OAI21_X1 U3000 ( .B1(n3309), .B2(n2395), .A(n2393), .ZN(n4154) );
  NAND2_X1 U3001 ( .A1(n3309), .A2(n2393), .ZN(n2392) );
  NAND3_X1 U3002 ( .A1(n2407), .A2(n2230), .A3(n2402), .ZN(n2401) );
  OAI21_X1 U3003 ( .B1(n2405), .B2(n2406), .A(n2404), .ZN(n3194) );
  NAND2_X1 U3004 ( .A1(n3042), .A2(n3758), .ZN(n2406) );
  NAND3_X1 U3005 ( .A1(n3042), .A2(n3758), .A3(n2407), .ZN(n2403) );
  NAND2_X1 U3006 ( .A1(n2678), .A2(n2410), .ZN(n2409) );
  NAND2_X1 U3007 ( .A1(n2412), .A2(n2413), .ZN(n3923) );
  NAND2_X1 U3008 ( .A1(n3948), .A2(n2415), .ZN(n2412) );
  NAND2_X1 U3009 ( .A1(n3948), .A2(n2422), .ZN(n2414) );
  OR2_X1 U3010 ( .A1(n3948), .A2(n3737), .ZN(n2418) );
  NAND2_X1 U3011 ( .A1(n2492), .A2(REG1_REG_2__SCAN_IN), .ZN(n2424) );
  NAND2_X1 U3012 ( .A1(n2503), .A2(n2504), .ZN(n2426) );
  NAND2_X1 U3013 ( .A1(n2930), .A2(n2996), .ZN(n3665) );
  NAND2_X1 U3014 ( .A1(n2425), .A2(n2424), .ZN(n2930) );
  AND2_X2 U3015 ( .A1(n2451), .A2(n2430), .ZN(n2773) );
  NOR2_X1 U3016 ( .A1(n2646), .A2(n2456), .ZN(n2784) );
  BUF_X4 U3017 ( .A(n3033), .Z(n3448) );
  NAND2_X1 U3018 ( .A1(n2950), .A2(n2941), .ZN(n3179) );
  INV_X1 U3019 ( .A(n2949), .ZN(n3031) );
  OR2_X1 U3020 ( .A1(n2950), .A2(n2951), .ZN(n2433) );
  AND2_X1 U3021 ( .A1(n2585), .A2(n2584), .ZN(n2434) );
  AND2_X1 U3022 ( .A1(n3552), .A2(n4503), .ZN(n2435) );
  AND2_X1 U3023 ( .A1(n2463), .A2(IR_REG_27__SCAN_IN), .ZN(n2436) );
  INV_X1 U3024 ( .A(IR_REG_9__SCAN_IN), .ZN(n2444) );
  AND2_X1 U3025 ( .A1(n4016), .A2(n2765), .ZN(n4033) );
  OR2_X1 U3026 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2437)
         );
  INV_X2 U3027 ( .A(n3822), .ZN(U4043) );
  OR2_X1 U3028 ( .A1(n3340), .A2(n4281), .ZN(n2439) );
  OR2_X1 U3029 ( .A1(n3340), .A2(n4237), .ZN(n2440) );
  AND2_X1 U3030 ( .A1(n3823), .A2(n3190), .ZN(n2441) );
  INV_X1 U3031 ( .A(IR_REG_0__SCAN_IN), .ZN(n2498) );
  OR2_X2 U3032 ( .A1(n3508), .A2(n4585), .ZN(n3033) );
  INV_X1 U3033 ( .A(n4125), .ZN(n2659) );
  INV_X1 U3034 ( .A(n3818), .ZN(n2618) );
  OR2_X1 U3035 ( .A1(n2618), .A2(n3376), .ZN(n2617) );
  INV_X1 U3036 ( .A(n3411), .ZN(n3412) );
  INV_X1 U3037 ( .A(n3394), .ZN(n3395) );
  OR2_X1 U3038 ( .A1(n4092), .A2(n4074), .ZN(n2676) );
  INV_X1 U3039 ( .A(IR_REG_21__SCAN_IN), .ZN(n2738) );
  OAI22_X1 U3040 ( .A1(n2835), .A2(n3033), .B1(n2979), .B2(n3031), .ZN(n2990)
         );
  NAND2_X1 U3041 ( .A1(n3405), .A2(n2659), .ZN(n2660) );
  OR2_X1 U3042 ( .A1(n3480), .A2(n3481), .ZN(n3436) );
  INV_X1 U3043 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2560) );
  NAND2_X1 U3044 ( .A1(n2224), .A2(DATAI_1_), .ZN(n2490) );
  NAND2_X1 U3045 ( .A1(n4127), .A2(n4147), .ZN(n2641) );
  AND2_X1 U3046 ( .A1(n3697), .A2(n3683), .ZN(n3322) );
  AND2_X1 U3047 ( .A1(n2942), .A2(n2771), .ZN(n2936) );
  AND2_X1 U3048 ( .A1(n3713), .A2(DATAI_28_), .ZN(n3921) );
  INV_X1 U3049 ( .A(IR_REG_22__SCAN_IN), .ZN(n2746) );
  INV_X1 U3050 ( .A(n3183), .ZN(n3184) );
  INV_X1 U3051 ( .A(REG3_REG_19__SCAN_IN), .ZN(n3504) );
  INV_X1 U3052 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3612) );
  INV_X1 U3053 ( .A(n4294), .ZN(n2874) );
  INV_X1 U3054 ( .A(n4540), .ZN(n2880) );
  INV_X1 U3055 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4301) );
  INV_X1 U3056 ( .A(n4287), .ZN(n2981) );
  AND4_X1 U3057 ( .A1(n2735), .A2(n2734), .A3(n2733), .A4(n2732), .ZN(n3917)
         );
  INV_X1 U3058 ( .A(n3973), .ZN(n3935) );
  INV_X1 U3059 ( .A(n4034), .ZN(n3999) );
  INV_X1 U3060 ( .A(n4033), .ZN(n2692) );
  AND4_X1 U3061 ( .A1(n2473), .A2(n2472), .A3(n2471), .A4(n2470), .ZN(n4989)
         );
  NOR2_X1 U3062 ( .A1(n2585), .A2(n2584), .ZN(n2598) );
  OR2_X1 U3063 ( .A1(n2771), .A2(n4562), .ZN(n2847) );
  INV_X1 U3064 ( .A(n4162), .ZN(n4490) );
  INV_X1 U3065 ( .A(n4065), .ZN(n4074) );
  OR2_X1 U3066 ( .A1(n3783), .A2(n3776), .ZN(n4153) );
  INV_X1 U3067 ( .A(n4055), .ZN(n4495) );
  INV_X1 U3068 ( .A(n3351), .ZN(n3496) );
  AND2_X1 U3069 ( .A1(n3525), .A2(n3521), .ZN(n3522) );
  OR2_X1 U3070 ( .A1(n2679), .A2(n3543), .ZN(n2686) );
  NOR2_X1 U3071 ( .A1(n4301), .A2(n2630), .ZN(n2650) );
  INV_X1 U3072 ( .A(n3376), .ZN(n3606) );
  INV_X1 U3073 ( .A(n4315), .ZN(n3619) );
  INV_X1 U3074 ( .A(n4324), .ZN(n4309) );
  INV_X1 U3075 ( .A(n2622), .ZN(n2623) );
  AND4_X1 U3076 ( .A1(n2627), .A2(n2626), .A3(n2625), .A4(n2624), .ZN(n4299)
         );
  INV_X1 U3077 ( .A(n3552), .ZN(n3364) );
  INV_X1 U3078 ( .A(n3887), .ZN(n3888) );
  NAND2_X1 U3079 ( .A1(n2772), .A2(n3805), .ZN(n4145) );
  OR2_X1 U3080 ( .A1(n2846), .A2(n2935), .ZN(n2848) );
  INV_X1 U3081 ( .A(n3308), .ZN(n4514) );
  AOI21_X1 U3082 ( .B1(n2845), .B2(n4866), .A(n2866), .ZN(n2935) );
  NAND2_X1 U3083 ( .A1(n2780), .A2(n2749), .ZN(n4562) );
  NAND2_X1 U3084 ( .A1(n3301), .A2(n4562), .ZN(n4577) );
  AND2_X1 U3085 ( .A1(n2816), .A2(n2815), .ZN(n2823) );
  INV_X1 U3086 ( .A(IR_REG_30__SCAN_IN), .ZN(n3337) );
  AND2_X1 U3087 ( .A1(n2889), .A2(n2869), .ZN(n4473) );
  OR3_X1 U3088 ( .A1(n2957), .A2(n2956), .A3(n2955), .ZN(n4324) );
  AND2_X1 U3089 ( .A1(n3030), .A2(n3029), .ZN(n4331) );
  INV_X1 U3090 ( .A(n3493), .ZN(n3820) );
  INV_X1 U3091 ( .A(n4531), .ZN(n4427) );
  INV_X1 U3092 ( .A(n4513), .ZN(n4135) );
  INV_X1 U3093 ( .A(n4068), .ZN(n4155) );
  NAND2_X1 U3094 ( .A1(n4610), .A2(n4585), .ZN(n4237) );
  INV_X1 U3095 ( .A(n4610), .ZN(n4607) );
  NAND2_X1 U3096 ( .A1(n4596), .A2(n4585), .ZN(n4281) );
  INV_X1 U3097 ( .A(n4596), .ZN(n4594) );
  INV_X1 U3098 ( .A(n4521), .ZN(n4520) );
  NAND2_X1 U3099 ( .A1(n2865), .A2(n2945), .ZN(n4521) );
  XNOR2_X1 U3100 ( .A(n2640), .B(n4698), .ZN(n4527) );
  OR2_X1 U3101 ( .A1(n2449), .A2(n2794), .ZN(n2447) );
  XNOR2_X1 U3102 ( .A(n2447), .B(IR_REG_14__SCAN_IN), .ZN(n4444) );
  NOR2_X1 U3103 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2455)
         );
  NOR2_X1 U3104 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2454)
         );
  NAND4_X1 U3105 ( .A1(n2455), .A2(n2454), .A3(n2453), .A4(n2452), .ZN(n2456)
         );
  INV_X1 U3106 ( .A(IR_REG_26__SCAN_IN), .ZN(n2457) );
  AOI21_X1 U3107 ( .B1(n2890), .B2(IR_REG_28__SCAN_IN), .A(n2436), .ZN(n2459)
         );
  NAND2_X4 U3108 ( .A1(n2460), .A2(n2459), .ZN(n3713) );
  MUX2_X1 U3109 ( .A(n4444), .B(DATAI_14_), .S(n3713), .Z(n3317) );
  NOR2_X1 U3110 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_29__SCAN_IN), .ZN(n2461)
         );
  NAND2_X1 U3111 ( .A1(n2773), .A2(n2461), .ZN(n3336) );
  XNOR2_X2 U3112 ( .A(n2462), .B(IR_REG_30__SCAN_IN), .ZN(n4283) );
  INV_X1 U3113 ( .A(n4283), .ZN(n2466) );
  NAND2_X1 U3114 ( .A1(n2773), .A2(n2463), .ZN(n2464) );
  NAND2_X1 U3115 ( .A1(n2573), .A2(REG1_REG_14__SCAN_IN), .ZN(n2473) );
  NAND2_X1 U3116 ( .A1(n2720), .A2(REG0_REG_14__SCAN_IN), .ZN(n2472) );
  INV_X1 U3117 ( .A(n2468), .ZN(n2467) );
  BUF_X4 U3118 ( .A(n2231), .Z(n3651) );
  NAND2_X1 U3119 ( .A1(n3651), .A2(REG2_REG_14__SCAN_IN), .ZN(n2471) );
  NAND2_X1 U3120 ( .A1(n2477), .A2(REG3_REG_6__SCAN_IN), .ZN(n2540) );
  INV_X1 U3121 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2539) );
  NOR2_X1 U3122 ( .A1(n2540), .A2(n2539), .ZN(n2548) );
  NAND2_X1 U3123 ( .A1(n2548), .A2(REG3_REG_8__SCAN_IN), .ZN(n2561) );
  OR2_X1 U3124 ( .A1(n2611), .A2(REG3_REG_14__SCAN_IN), .ZN(n2469) );
  NAND2_X1 U3125 ( .A1(n2611), .A2(REG3_REG_14__SCAN_IN), .ZN(n2622) );
  NAND2_X1 U3126 ( .A1(n2469), .A2(n2622), .ZN(n3471) );
  OR2_X1 U3127 ( .A1(n2222), .A2(n3471), .ZN(n2470) );
  INV_X1 U3128 ( .A(n4989), .ZN(n2621) );
  OR2_X1 U3129 ( .A1(n2474), .A2(n2794), .ZN(n2475) );
  XNOR2_X1 U3130 ( .A(n2475), .B(IR_REG_6__SCAN_IN), .ZN(n4540) );
  INV_X1 U3131 ( .A(DATAI_6_), .ZN(n2476) );
  MUX2_X1 U3132 ( .A(n2880), .B(n2476), .S(n3713), .Z(n3203) );
  INV_X1 U3133 ( .A(n3203), .ZN(n3197) );
  INV_X1 U3134 ( .A(n2477), .ZN(n2530) );
  INV_X1 U3135 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3147) );
  NAND2_X1 U3136 ( .A1(n2530), .A2(n3147), .ZN(n2478) );
  AND2_X1 U3137 ( .A1(n2478), .A2(n2540), .ZN(n4509) );
  INV_X1 U3138 ( .A(n4509), .ZN(n3151) );
  OR2_X1 U3139 ( .A1(n2222), .A2(n3151), .ZN(n2482) );
  NAND2_X1 U3140 ( .A1(n2720), .A2(REG0_REG_6__SCAN_IN), .ZN(n2481) );
  NAND2_X1 U3141 ( .A1(n3651), .A2(REG2_REG_6__SCAN_IN), .ZN(n2480) );
  NAND2_X1 U3142 ( .A1(n2573), .A2(REG1_REG_6__SCAN_IN), .ZN(n2479) );
  NAND4_X1 U3143 ( .A1(n2482), .A2(n2481), .A3(n2480), .A4(n2479), .ZN(n3136)
         );
  NAND2_X1 U3144 ( .A1(n2492), .A2(REG1_REG_1__SCAN_IN), .ZN(n2487) );
  NAND2_X1 U3145 ( .A1(n2231), .A2(REG2_REG_1__SCAN_IN), .ZN(n2486) );
  INV_X1 U3146 ( .A(n2502), .ZN(n2483) );
  NAND2_X1 U3147 ( .A1(n2483), .A2(REG3_REG_1__SCAN_IN), .ZN(n2485) );
  NAND2_X1 U31480 ( .A1(n2501), .A2(REG0_REG_1__SCAN_IN), .ZN(n2484) );
  AND4_X2 U31490 ( .A1(n2487), .A2(n2486), .A3(n2485), .A4(n2484), .ZN(n2835)
         );
  INV_X1 U3150 ( .A(n2894), .ZN(n4286) );
  OAI21_X1 U3151 ( .B1(n2224), .B2(n2894), .A(n2490), .ZN(n2491) );
  NAND2_X1 U3152 ( .A1(n2499), .A2(n2979), .ZN(n3659) );
  NAND2_X1 U3153 ( .A1(n2835), .A2(n2491), .ZN(n2750) );
  NAND2_X1 U3154 ( .A1(n2501), .A2(REG0_REG_0__SCAN_IN), .ZN(n2495) );
  NAND2_X1 U3155 ( .A1(n2492), .A2(REG1_REG_0__SCAN_IN), .ZN(n2494) );
  NAND2_X1 U3156 ( .A1(n2231), .A2(REG2_REG_0__SCAN_IN), .ZN(n2493) );
  NAND4_X1 U3157 ( .A1(n2496), .A2(n2495), .A3(n2494), .A4(n2493), .ZN(n3825)
         );
  NAND2_X1 U3158 ( .A1(n2499), .A2(n2491), .ZN(n2500) );
  NAND2_X1 U3159 ( .A1(n3076), .A2(n2500), .ZN(n2833) );
  INV_X1 U3160 ( .A(n2833), .ZN(n2508) );
  NAND2_X1 U3161 ( .A1(n2501), .A2(REG0_REG_2__SCAN_IN), .ZN(n2504) );
  INV_X1 U3162 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2851) );
  OR2_X1 U3163 ( .A1(n2502), .A2(n2851), .ZN(n2503) );
  XNOR2_X2 U3164 ( .A(n2505), .B(IR_REG_2__SCAN_IN), .ZN(n4285) );
  NAND2_X1 U3165 ( .A1(n3093), .A2(n3005), .ZN(n3662) );
  NAND2_X1 U3166 ( .A1(n3665), .A2(n3662), .ZN(n2752) );
  NAND2_X1 U3167 ( .A1(n2508), .A2(n2752), .ZN(n2831) );
  NAND2_X1 U3168 ( .A1(n3093), .A2(n2996), .ZN(n2509) );
  NAND2_X1 U3169 ( .A1(n2831), .A2(n2509), .ZN(n3087) );
  NAND2_X1 U3170 ( .A1(n2720), .A2(REG0_REG_3__SCAN_IN), .ZN(n2514) );
  NAND2_X1 U3171 ( .A1(n3651), .A2(REG2_REG_3__SCAN_IN), .ZN(n2513) );
  NAND2_X1 U3172 ( .A1(n2573), .A2(REG1_REG_3__SCAN_IN), .ZN(n2512) );
  OR2_X1 U3173 ( .A1(n2222), .A2(REG3_REG_3__SCAN_IN), .ZN(n2511) );
  INV_X1 U3174 ( .A(n3067), .ZN(n3824) );
  NAND2_X1 U3175 ( .A1(n2515), .A2(IR_REG_31__SCAN_IN), .ZN(n2521) );
  XNOR2_X1 U3176 ( .A(n2521), .B(IR_REG_3__SCAN_IN), .ZN(n4294) );
  MUX2_X1 U3177 ( .A(n4294), .B(DATAI_3_), .S(n3713), .Z(n3090) );
  NOR2_X1 U3178 ( .A1(n3824), .A2(n3090), .ZN(n2516) );
  XNOR2_X1 U3179 ( .A(REG3_REG_4__SCAN_IN), .B(REG3_REG_3__SCAN_IN), .ZN(n3072) );
  OR2_X1 U3180 ( .A1(n2222), .A2(n3072), .ZN(n2520) );
  NAND2_X1 U3181 ( .A1(n2573), .A2(REG1_REG_4__SCAN_IN), .ZN(n2519) );
  NAND2_X1 U3182 ( .A1(n2720), .A2(REG0_REG_4__SCAN_IN), .ZN(n2518) );
  NAND2_X1 U3183 ( .A1(n3651), .A2(REG2_REG_4__SCAN_IN), .ZN(n2517) );
  NAND4_X1 U3184 ( .A1(n2520), .A2(n2519), .A3(n2518), .A4(n2517), .ZN(n3091)
         );
  NAND2_X1 U3185 ( .A1(n2521), .A2(n4793), .ZN(n2522) );
  NAND2_X1 U3186 ( .A1(n2522), .A2(IR_REG_31__SCAN_IN), .ZN(n2524) );
  XNOR2_X1 U3187 ( .A(n2524), .B(n2523), .ZN(n2903) );
  INV_X1 U3188 ( .A(DATAI_4_), .ZN(n2525) );
  MUX2_X1 U3189 ( .A(n2903), .B(n2525), .S(n3713), .Z(n3061) );
  NOR2_X1 U3190 ( .A1(n3091), .A2(n3061), .ZN(n2753) );
  INV_X1 U3191 ( .A(n2753), .ZN(n3668) );
  NAND2_X1 U3192 ( .A1(n3091), .A2(n3061), .ZN(n3670) );
  NAND2_X1 U3193 ( .A1(n3668), .A2(n3670), .ZN(n3758) );
  NAND2_X1 U3194 ( .A1(n2573), .A2(REG1_REG_5__SCAN_IN), .ZN(n2534) );
  NAND2_X1 U3195 ( .A1(n2720), .A2(REG0_REG_5__SCAN_IN), .ZN(n2533) );
  NAND2_X1 U3196 ( .A1(n3651), .A2(REG2_REG_5__SCAN_IN), .ZN(n2532) );
  INV_X1 U3197 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2528) );
  NAND2_X1 U3198 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2527) );
  NAND2_X1 U3199 ( .A1(n2528), .A2(n2527), .ZN(n2529) );
  NAND2_X1 U3200 ( .A1(n2530), .A2(n2529), .ZN(n3117) );
  OR2_X1 U3201 ( .A1(n2222), .A2(n3117), .ZN(n2531) );
  NAND2_X1 U3202 ( .A1(n2535), .A2(IR_REG_31__SCAN_IN), .ZN(n2536) );
  XNOR2_X1 U3203 ( .A(n2536), .B(IR_REG_5__SCAN_IN), .ZN(n2893) );
  MUX2_X1 U3204 ( .A(n2893), .B(DATAI_5_), .S(n3713), .Z(n3114) );
  NAND2_X1 U3205 ( .A1(n3044), .A2(n3114), .ZN(n2537) );
  INV_X1 U3206 ( .A(n3136), .ZN(n3187) );
  NAND2_X1 U3207 ( .A1(n2573), .A2(REG1_REG_7__SCAN_IN), .ZN(n2545) );
  NAND2_X1 U3208 ( .A1(n2720), .A2(REG0_REG_7__SCAN_IN), .ZN(n2544) );
  NAND2_X1 U3209 ( .A1(n3651), .A2(REG2_REG_7__SCAN_IN), .ZN(n2543) );
  AND2_X1 U32100 ( .A1(n2540), .A2(n2539), .ZN(n2541) );
  OR2_X1 U32110 ( .A1(n2541), .A2(n2548), .ZN(n3193) );
  OR2_X1 U32120 ( .A1(n2222), .A2(n3193), .ZN(n2542) );
  OR2_X1 U32130 ( .A1(n2546), .A2(n2794), .ZN(n2555) );
  XNOR2_X1 U32140 ( .A(n2555), .B(IR_REG_7__SCAN_IN), .ZN(n2892) );
  MUX2_X1 U32150 ( .A(n2892), .B(DATAI_7_), .S(n3713), .Z(n3190) );
  NAND2_X1 U32160 ( .A1(n3230), .A2(n3190), .ZN(n2754) );
  AND2_X1 U32170 ( .A1(n3823), .A2(n3181), .ZN(n3676) );
  INV_X1 U32180 ( .A(n3676), .ZN(n2547) );
  NAND2_X1 U32190 ( .A1(n2754), .A2(n2547), .ZN(n3757) );
  OR2_X1 U32200 ( .A1(n2548), .A2(REG3_REG_8__SCAN_IN), .ZN(n2549) );
  NAND2_X1 U32210 ( .A1(n2561), .A2(n2549), .ZN(n3235) );
  OR2_X1 U32220 ( .A1(n2222), .A2(n3235), .ZN(n2553) );
  NAND2_X1 U32230 ( .A1(n2573), .A2(REG1_REG_8__SCAN_IN), .ZN(n2552) );
  NAND2_X1 U32240 ( .A1(n2720), .A2(REG0_REG_8__SCAN_IN), .ZN(n2551) );
  NAND2_X1 U32250 ( .A1(n3651), .A2(REG2_REG_8__SCAN_IN), .ZN(n2550) );
  NAND4_X1 U32260 ( .A1(n2553), .A2(n2552), .A3(n2551), .A4(n2550), .ZN(n3821)
         );
  INV_X1 U32270 ( .A(IR_REG_7__SCAN_IN), .ZN(n2554) );
  NAND2_X1 U32280 ( .A1(n2555), .A2(n2554), .ZN(n2556) );
  NAND2_X1 U32290 ( .A1(n2556), .A2(IR_REG_31__SCAN_IN), .ZN(n2557) );
  XNOR2_X1 U32300 ( .A(n2557), .B(IR_REG_8__SCAN_IN), .ZN(n2909) );
  INV_X1 U32310 ( .A(DATAI_8_), .ZN(n2558) );
  MUX2_X1 U32320 ( .A(n4537), .B(n2558), .S(n3713), .Z(n3227) );
  NAND2_X1 U32330 ( .A1(n3821), .A2(n3232), .ZN(n2559) );
  INV_X1 U32340 ( .A(n3821), .ZN(n3266) );
  AOI22_X2 U32350 ( .A1(n3157), .A2(n2559), .B1(n3266), .B2(n3227), .ZN(n3166)
         );
  NAND2_X1 U32360 ( .A1(n2573), .A2(REG1_REG_9__SCAN_IN), .ZN(n2566) );
  NAND2_X1 U32370 ( .A1(n2720), .A2(REG0_REG_9__SCAN_IN), .ZN(n2565) );
  NAND2_X1 U32380 ( .A1(n3651), .A2(REG2_REG_9__SCAN_IN), .ZN(n2564) );
  NAND2_X1 U32390 ( .A1(n2561), .A2(n2560), .ZN(n2562) );
  NAND2_X1 U32400 ( .A1(n2571), .A2(n2562), .ZN(n3269) );
  OR2_X1 U32410 ( .A1(n2222), .A2(n3269), .ZN(n2563) );
  NAND2_X1 U32420 ( .A1(n2546), .A2(n2567), .ZN(n2568) );
  NAND2_X1 U32430 ( .A1(n2568), .A2(IR_REG_31__SCAN_IN), .ZN(n2569) );
  XNOR2_X1 U32440 ( .A(n2569), .B(IR_REG_9__SCAN_IN), .ZN(n4535) );
  MUX2_X1 U32450 ( .A(n4535), .B(DATAI_9_), .S(n3713), .Z(n3268) );
  INV_X1 U32460 ( .A(n3268), .ZN(n3256) );
  NAND2_X1 U32470 ( .A1(n3493), .A2(n3256), .ZN(n2570) );
  NAND2_X1 U32480 ( .A1(n2571), .A2(n2914), .ZN(n2572) );
  NAND2_X1 U32490 ( .A1(n2585), .A2(n2572), .ZN(n3499) );
  OR2_X1 U32500 ( .A1(n2222), .A2(n3499), .ZN(n2577) );
  NAND2_X1 U32510 ( .A1(n2573), .A2(REG1_REG_10__SCAN_IN), .ZN(n2576) );
  NAND2_X1 U32520 ( .A1(n2720), .A2(REG0_REG_10__SCAN_IN), .ZN(n2575) );
  NAND2_X1 U32530 ( .A1(n3651), .A2(REG2_REG_10__SCAN_IN), .ZN(n2574) );
  NAND4_X1 U32540 ( .A1(n2577), .A2(n2576), .A3(n2575), .A4(n2574), .ZN(n3819)
         );
  INV_X1 U32550 ( .A(n3819), .ZN(n4492) );
  NAND2_X1 U32560 ( .A1(n2578), .A2(IR_REG_31__SCAN_IN), .ZN(n2580) );
  XNOR2_X1 U32570 ( .A(n2580), .B(n2579), .ZN(n2917) );
  INV_X1 U32580 ( .A(DATAI_10_), .ZN(n4881) );
  MUX2_X1 U32590 ( .A(n2917), .B(n4881), .S(n3713), .Z(n3351) );
  NAND2_X1 U32600 ( .A1(n3819), .A2(n3496), .ZN(n2581) );
  NAND2_X1 U32610 ( .A1(n3241), .A2(n2581), .ZN(n2583) );
  NAND2_X1 U32620 ( .A1(n3351), .A2(n4492), .ZN(n2582) );
  NAND2_X1 U32630 ( .A1(n2583), .A2(n2582), .ZN(n4487) );
  NAND2_X1 U32640 ( .A1(n2573), .A2(REG1_REG_11__SCAN_IN), .ZN(n2590) );
  NAND2_X1 U32650 ( .A1(n2720), .A2(REG0_REG_11__SCAN_IN), .ZN(n2589) );
  NAND2_X1 U32660 ( .A1(n3651), .A2(REG2_REG_11__SCAN_IN), .ZN(n2588) );
  NOR2_X1 U32670 ( .A1(n2598), .A2(n2434), .ZN(n4501) );
  INV_X1 U32680 ( .A(n4501), .ZN(n2586) );
  OR2_X1 U32690 ( .A1(n2222), .A2(n2586), .ZN(n2587) );
  OR2_X1 U32700 ( .A1(n2578), .A2(IR_REG_10__SCAN_IN), .ZN(n2591) );
  NAND2_X1 U32710 ( .A1(n2591), .A2(IR_REG_31__SCAN_IN), .ZN(n2594) );
  INV_X1 U32720 ( .A(n2594), .ZN(n2592) );
  NAND2_X1 U32730 ( .A1(n2592), .A2(IR_REG_11__SCAN_IN), .ZN(n2595) );
  NAND2_X1 U32740 ( .A1(n2594), .A2(n2593), .ZN(n2604) );
  MUX2_X1 U32750 ( .A(n3875), .B(DATAI_11_), .S(n3713), .Z(n2596) );
  NAND2_X1 U32760 ( .A1(n3552), .A2(n2596), .ZN(n3701) );
  INV_X1 U32770 ( .A(n3695), .ZN(n2597) );
  NAND2_X1 U32780 ( .A1(n3701), .A2(n2597), .ZN(n4489) );
  NOR2_X1 U32790 ( .A1(n2598), .A2(REG3_REG_12__SCAN_IN), .ZN(n2599) );
  OR2_X1 U32800 ( .A1(n2609), .A2(n2599), .ZN(n3280) );
  OR2_X1 U32810 ( .A1(n2222), .A2(n3280), .ZN(n2603) );
  NAND2_X1 U32820 ( .A1(n2573), .A2(REG1_REG_12__SCAN_IN), .ZN(n2602) );
  NAND2_X1 U32830 ( .A1(n2720), .A2(REG0_REG_12__SCAN_IN), .ZN(n2601) );
  NAND2_X1 U32840 ( .A1(n3651), .A2(REG2_REG_12__SCAN_IN), .ZN(n2600) );
  NAND4_X1 U32850 ( .A1(n2603), .A2(n2602), .A3(n2601), .A4(n2600), .ZN(n4494)
         );
  INV_X1 U32860 ( .A(n4494), .ZN(n3604) );
  NAND2_X1 U32870 ( .A1(n2604), .A2(IR_REG_31__SCAN_IN), .ZN(n2605) );
  XNOR2_X1 U32880 ( .A(n2605), .B(IR_REG_12__SCAN_IN), .ZN(n4531) );
  INV_X1 U32890 ( .A(DATAI_12_), .ZN(n2606) );
  MUX2_X1 U32900 ( .A(n4427), .B(n2606), .S(n3713), .Z(n3551) );
  NAND2_X1 U32910 ( .A1(n3604), .A2(n3551), .ZN(n2608) );
  NOR2_X1 U32920 ( .A1(n2609), .A2(REG3_REG_13__SCAN_IN), .ZN(n2610) );
  OR2_X1 U32930 ( .A1(n2611), .A2(n2610), .ZN(n3609) );
  OR2_X1 U32940 ( .A1(n2222), .A2(n3609), .ZN(n2615) );
  NAND2_X1 U32950 ( .A1(n2573), .A2(REG1_REG_13__SCAN_IN), .ZN(n2614) );
  NAND2_X1 U32960 ( .A1(n2720), .A2(REG0_REG_13__SCAN_IN), .ZN(n2613) );
  NAND2_X1 U32970 ( .A1(n3651), .A2(REG2_REG_13__SCAN_IN), .ZN(n2612) );
  NAND4_X1 U32980 ( .A1(n2615), .A2(n2614), .A3(n2613), .A4(n2612), .ZN(n3818)
         );
  OR2_X1 U32990 ( .A1(n2253), .A2(n2794), .ZN(n2616) );
  XNOR2_X1 U33000 ( .A(n2616), .B(IR_REG_13__SCAN_IN), .ZN(n3878) );
  MUX2_X1 U33010 ( .A(n4530), .B(n4884), .S(n3713), .Z(n3376) );
  NAND2_X1 U33020 ( .A1(n3291), .A2(n2617), .ZN(n2620) );
  NAND2_X1 U33030 ( .A1(n2620), .A2(n2619), .ZN(n3309) );
  NAND2_X1 U33040 ( .A1(n4989), .A2(n3317), .ZN(n3698) );
  NAND2_X1 U33050 ( .A1(n2621), .A2(n3472), .ZN(n3682) );
  NAND2_X1 U33060 ( .A1(n3698), .A2(n3682), .ZN(n3762) );
  NAND2_X1 U33070 ( .A1(n2720), .A2(REG0_REG_15__SCAN_IN), .ZN(n2627) );
  NAND2_X1 U33080 ( .A1(n3651), .A2(REG2_REG_15__SCAN_IN), .ZN(n2626) );
  NAND2_X1 U33090 ( .A1(n2573), .A2(REG1_REG_15__SCAN_IN), .ZN(n2625) );
  NAND2_X1 U33100 ( .A1(REG3_REG_15__SCAN_IN), .A2(n2623), .ZN(n2630) );
  OAI21_X1 U33110 ( .B1(REG3_REG_15__SCAN_IN), .B2(n2623), .A(n2630), .ZN(
        n4330) );
  OR2_X1 U33120 ( .A1(n2222), .A2(n4330), .ZN(n2624) );
  INV_X1 U33130 ( .A(n4299), .ZN(n3817) );
  NAND2_X1 U33140 ( .A1(n2628), .A2(IR_REG_31__SCAN_IN), .ZN(n2638) );
  MUX2_X1 U33150 ( .A(n4457), .B(DATAI_15_), .S(n3713), .Z(n3326) );
  NOR2_X1 U33160 ( .A1(n3817), .A2(n3326), .ZN(n2629) );
  INV_X1 U33170 ( .A(n2630), .ZN(n2632) );
  INV_X1 U33180 ( .A(n2650), .ZN(n2631) );
  OAI21_X1 U33190 ( .B1(REG3_REG_16__SCAN_IN), .B2(n2632), .A(n2631), .ZN(
        n4313) );
  OR2_X1 U33200 ( .A1(n2222), .A2(n4313), .ZN(n2636) );
  NAND2_X1 U33210 ( .A1(n2720), .A2(REG0_REG_16__SCAN_IN), .ZN(n2635) );
  NAND2_X1 U33220 ( .A1(n3651), .A2(REG2_REG_16__SCAN_IN), .ZN(n2634) );
  NAND2_X1 U33230 ( .A1(n2573), .A2(REG1_REG_16__SCAN_IN), .ZN(n2633) );
  NAND4_X1 U33240 ( .A1(n2636), .A2(n2635), .A3(n2634), .A4(n2633), .ZN(n4127)
         );
  INV_X1 U33250 ( .A(IR_REG_15__SCAN_IN), .ZN(n2637) );
  NAND2_X1 U33260 ( .A1(n2638), .A2(n2637), .ZN(n2639) );
  NAND2_X1 U33270 ( .A1(n2639), .A2(IR_REG_31__SCAN_IN), .ZN(n2640) );
  INV_X1 U33280 ( .A(DATAI_16_), .ZN(n4526) );
  MUX2_X1 U33290 ( .A(n4527), .B(n4526), .S(n3713), .Z(n4303) );
  AND2_X1 U33300 ( .A1(n4127), .A2(n4303), .ZN(n3783) );
  NOR2_X1 U33310 ( .A1(n4127), .A2(n4303), .ZN(n3776) );
  INV_X1 U33320 ( .A(n4127), .ZN(n4314) );
  NAND2_X1 U33330 ( .A1(n4152), .A2(n2641), .ZN(n4121) );
  NAND2_X1 U33340 ( .A1(n2720), .A2(REG0_REG_17__SCAN_IN), .ZN(n2645) );
  NAND2_X1 U33350 ( .A1(n3651), .A2(REG2_REG_17__SCAN_IN), .ZN(n2644) );
  NAND2_X1 U33360 ( .A1(n2573), .A2(REG1_REG_17__SCAN_IN), .ZN(n2643) );
  XNOR2_X1 U33370 ( .A(REG3_REG_17__SCAN_IN), .B(n2650), .ZN(n4136) );
  OR2_X1 U33380 ( .A1(n2222), .A2(n4136), .ZN(n2642) );
  INV_X1 U33390 ( .A(n4300), .ZN(n4142) );
  NAND2_X1 U33400 ( .A1(n2646), .A2(IR_REG_31__SCAN_IN), .ZN(n2647) );
  MUX2_X1 U33410 ( .A(n3883), .B(DATAI_17_), .S(n3713), .Z(n4124) );
  NAND2_X1 U33420 ( .A1(n4121), .A2(n2252), .ZN(n2649) );
  INV_X1 U33430 ( .A(n4124), .ZN(n4133) );
  NAND2_X1 U33440 ( .A1(n2649), .A2(n2648), .ZN(n4114) );
  NAND2_X1 U33450 ( .A1(n2651), .A2(REG3_REG_18__SCAN_IN), .ZN(n2661) );
  OAI21_X1 U33460 ( .B1(n2651), .B2(REG3_REG_18__SCAN_IN), .A(n2661), .ZN(
        n4111) );
  OR2_X1 U33470 ( .A1(n2222), .A2(n4111), .ZN(n2655) );
  NAND2_X1 U33480 ( .A1(n2573), .A2(REG1_REG_18__SCAN_IN), .ZN(n2654) );
  NAND2_X1 U33490 ( .A1(n2720), .A2(REG0_REG_18__SCAN_IN), .ZN(n2653) );
  NAND2_X1 U33500 ( .A1(n3651), .A2(REG2_REG_18__SCAN_IN), .ZN(n2652) );
  NAND4_X1 U33510 ( .A1(n2655), .A2(n2654), .A3(n2653), .A4(n2652), .ZN(n4125)
         );
  NAND2_X1 U33520 ( .A1(n2656), .A2(IR_REG_31__SCAN_IN), .ZN(n2657) );
  XNOR2_X1 U3353 ( .A(n2657), .B(n2667), .ZN(n3893) );
  INV_X1 U33540 ( .A(DATAI_18_), .ZN(n2658) );
  MUX2_X1 U3355 ( .A(n3893), .B(n2658), .S(n3713), .Z(n3405) );
  NOR2_X1 U3356 ( .A1(n4125), .A2(n3405), .ZN(n2760) );
  AND2_X1 U3357 ( .A1(n4125), .A2(n3405), .ZN(n4087) );
  NOR2_X1 U3358 ( .A1(n2760), .A2(n4087), .ZN(n4115) );
  OR2_X2 U3359 ( .A1(n4114), .A2(n4115), .ZN(n4112) );
  INV_X1 U3360 ( .A(n3405), .ZN(n4109) );
  AND2_X1 U3361 ( .A1(n2661), .A2(n3504), .ZN(n2662) );
  OR2_X1 U3362 ( .A1(n2662), .A2(n2670), .ZN(n4099) );
  OR2_X1 U3363 ( .A1(n2222), .A2(n4099), .ZN(n2666) );
  NAND2_X1 U3364 ( .A1(n2573), .A2(REG1_REG_19__SCAN_IN), .ZN(n2665) );
  NAND2_X1 U3365 ( .A1(n2720), .A2(REG0_REG_19__SCAN_IN), .ZN(n2664) );
  NAND2_X1 U3366 ( .A1(n3651), .A2(REG2_REG_19__SCAN_IN), .ZN(n2663) );
  NAND4_X1 U3367 ( .A1(n2666), .A2(n2665), .A3(n2664), .A4(n2663), .ZN(n4105)
         );
  INV_X1 U3368 ( .A(DATAI_19_), .ZN(n2669) );
  MUX2_X1 U3369 ( .A(n3905), .B(n2669), .S(n3713), .Z(n4097) );
  INV_X1 U3370 ( .A(n4097), .ZN(n4091) );
  NOR2_X1 U3371 ( .A1(n4105), .A2(n4091), .ZN(n3735) );
  NAND2_X1 U3372 ( .A1(n4105), .A2(n4091), .ZN(n3734) );
  NAND2_X1 U3373 ( .A1(n2670), .A2(REG3_REG_20__SCAN_IN), .ZN(n2679) );
  OR2_X1 U3374 ( .A1(n2670), .A2(REG3_REG_20__SCAN_IN), .ZN(n2671) );
  NAND2_X1 U3375 ( .A1(n2679), .A2(n2671), .ZN(n4079) );
  OR2_X1 U3376 ( .A1(n2222), .A2(n4079), .ZN(n2675) );
  NAND2_X1 U3377 ( .A1(n2573), .A2(REG1_REG_20__SCAN_IN), .ZN(n2674) );
  NAND2_X1 U3378 ( .A1(n2720), .A2(REG0_REG_20__SCAN_IN), .ZN(n2673) );
  NAND2_X1 U3379 ( .A1(n3651), .A2(REG2_REG_20__SCAN_IN), .ZN(n2672) );
  NAND4_X1 U3380 ( .A1(n2675), .A2(n2674), .A3(n2673), .A4(n2672), .ZN(n4092)
         );
  NAND2_X1 U3381 ( .A1(n3713), .A2(DATAI_20_), .ZN(n4065) );
  NAND2_X1 U3382 ( .A1(n4067), .A2(n2676), .ZN(n2678) );
  NAND2_X1 U3383 ( .A1(n4092), .A2(n4074), .ZN(n2677) );
  NAND2_X1 U3384 ( .A1(n2679), .A2(n3543), .ZN(n2680) );
  NAND2_X1 U3385 ( .A1(n2686), .A2(n2680), .ZN(n4059) );
  OR2_X1 U3386 ( .A1(n2222), .A2(n4059), .ZN(n2684) );
  NAND2_X1 U3387 ( .A1(n2573), .A2(REG1_REG_21__SCAN_IN), .ZN(n2683) );
  NAND2_X1 U3388 ( .A1(n2720), .A2(REG0_REG_21__SCAN_IN), .ZN(n2682) );
  NAND2_X1 U3389 ( .A1(n3651), .A2(REG2_REG_21__SCAN_IN), .ZN(n2681) );
  NAND4_X1 U3390 ( .A1(n2684), .A2(n2683), .A3(n2682), .A4(n2681), .ZN(n4075)
         );
  INV_X1 U3391 ( .A(n4075), .ZN(n3613) );
  NAND2_X1 U3392 ( .A1(n3713), .A2(DATAI_21_), .ZN(n3544) );
  NOR2_X1 U3393 ( .A1(n3613), .A2(n3544), .ZN(n2685) );
  NAND2_X1 U3394 ( .A1(n2573), .A2(REG1_REG_22__SCAN_IN), .ZN(n2691) );
  NAND2_X1 U3395 ( .A1(n2720), .A2(REG0_REG_22__SCAN_IN), .ZN(n2690) );
  NAND2_X1 U3396 ( .A1(n3651), .A2(REG2_REG_22__SCAN_IN), .ZN(n2689) );
  AND2_X1 U3397 ( .A1(n2686), .A2(n3612), .ZN(n2687) );
  OR2_X1 U3398 ( .A1(n2687), .A2(n2693), .ZN(n4040) );
  OR2_X1 U3399 ( .A1(n2222), .A2(n4040), .ZN(n2688) );
  NAND2_X1 U3400 ( .A1(n4056), .A2(n4041), .ZN(n4016) );
  INV_X1 U3401 ( .A(n4056), .ZN(n2922) );
  NAND2_X1 U3402 ( .A1(n2922), .A2(n4037), .ZN(n2765) );
  NAND2_X1 U3403 ( .A1(n4030), .A2(n2246), .ZN(n4010) );
  NOR2_X1 U3404 ( .A1(n2693), .A2(REG3_REG_23__SCAN_IN), .ZN(n2694) );
  OR2_X1 U3405 ( .A1(n2699), .A2(n2694), .ZN(n4024) );
  OR2_X1 U3406 ( .A1(n2222), .A2(n4024), .ZN(n2698) );
  NAND2_X1 U3407 ( .A1(n2573), .A2(REG1_REG_23__SCAN_IN), .ZN(n2697) );
  NAND2_X1 U3408 ( .A1(n2720), .A2(REG0_REG_23__SCAN_IN), .ZN(n2696) );
  NAND2_X1 U3409 ( .A1(n3651), .A2(REG2_REG_23__SCAN_IN), .ZN(n2695) );
  NAND4_X1 U3410 ( .A1(n2698), .A2(n2697), .A3(n2696), .A4(n2695), .ZN(n4034)
         );
  NAND2_X1 U3411 ( .A1(n3713), .A2(DATAI_23_), .ZN(n3484) );
  AND2_X1 U3412 ( .A1(n4034), .A2(n4020), .ZN(n3729) );
  NAND2_X1 U3413 ( .A1(n3999), .A2(n3484), .ZN(n3730) );
  NAND2_X1 U3414 ( .A1(n2699), .A2(REG3_REG_24__SCAN_IN), .ZN(n2707) );
  OR2_X1 U3415 ( .A1(n2699), .A2(REG3_REG_24__SCAN_IN), .ZN(n2700) );
  NAND2_X1 U3416 ( .A1(n2707), .A2(n2700), .ZN(n4002) );
  OR2_X1 U3417 ( .A1(n2222), .A2(n4002), .ZN(n2704) );
  NAND2_X1 U3418 ( .A1(n2573), .A2(REG1_REG_24__SCAN_IN), .ZN(n2703) );
  NAND2_X1 U3419 ( .A1(n2720), .A2(REG0_REG_24__SCAN_IN), .ZN(n2702) );
  NAND2_X1 U3420 ( .A1(n3651), .A2(REG2_REG_24__SCAN_IN), .ZN(n2701) );
  NAND4_X1 U3421 ( .A1(n2704), .A2(n2703), .A3(n2702), .A4(n2701), .ZN(n4021)
         );
  NAND2_X1 U3422 ( .A1(n3713), .A2(DATAI_24_), .ZN(n4001) );
  NAND2_X1 U3423 ( .A1(n4021), .A2(n3995), .ZN(n2706) );
  NOR2_X1 U3424 ( .A1(n4021), .A2(n3995), .ZN(n2705) );
  INV_X1 U3425 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3561) );
  NAND2_X1 U3426 ( .A1(n2707), .A2(n3561), .ZN(n2708) );
  NAND2_X1 U3427 ( .A1(n2723), .A2(n2708), .ZN(n3981) );
  OR2_X1 U3428 ( .A1(n2222), .A2(n3981), .ZN(n2712) );
  NAND2_X1 U3429 ( .A1(n2573), .A2(REG1_REG_25__SCAN_IN), .ZN(n2711) );
  NAND2_X1 U3430 ( .A1(n2720), .A2(REG0_REG_25__SCAN_IN), .ZN(n2710) );
  NAND2_X1 U3431 ( .A1(n3651), .A2(REG2_REG_25__SCAN_IN), .ZN(n2709) );
  NAND4_X1 U3432 ( .A1(n2712), .A2(n2711), .A3(n2710), .A4(n2709), .ZN(n3996)
         );
  INV_X1 U3433 ( .A(n3996), .ZN(n3956) );
  NAND2_X1 U3434 ( .A1(n3713), .A2(DATAI_25_), .ZN(n3979) );
  NAND2_X1 U3435 ( .A1(n3956), .A2(n3979), .ZN(n2713) );
  NAND2_X1 U3436 ( .A1(n3966), .A2(n2713), .ZN(n2715) );
  NAND2_X1 U3437 ( .A1(n3996), .A2(n3972), .ZN(n2714) );
  NAND2_X1 U3438 ( .A1(n2715), .A2(n2714), .ZN(n3948) );
  INV_X1 U3439 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3644) );
  XNOR2_X1 U3440 ( .A(n2723), .B(n3644), .ZN(n3960) );
  OR2_X1 U3441 ( .A1(n2222), .A2(n3960), .ZN(n2719) );
  NAND2_X1 U3442 ( .A1(n2573), .A2(REG1_REG_26__SCAN_IN), .ZN(n2718) );
  NAND2_X1 U3443 ( .A1(n2720), .A2(REG0_REG_26__SCAN_IN), .ZN(n2717) );
  NAND2_X1 U3444 ( .A1(n3651), .A2(REG2_REG_26__SCAN_IN), .ZN(n2716) );
  NAND4_X1 U3445 ( .A1(n2719), .A2(n2718), .A3(n2717), .A4(n2716), .ZN(n3973)
         );
  NAND2_X1 U3446 ( .A1(n3713), .A2(DATAI_26_), .ZN(n3959) );
  INV_X1 U3447 ( .A(n3959), .ZN(n2770) );
  AND2_X1 U3448 ( .A1(n3973), .A2(n2770), .ZN(n3737) );
  NAND2_X1 U3449 ( .A1(n3935), .A2(n3959), .ZN(n3738) );
  NAND2_X1 U3450 ( .A1(n2573), .A2(REG1_REG_27__SCAN_IN), .ZN(n2728) );
  NAND2_X1 U3451 ( .A1(n2720), .A2(REG0_REG_27__SCAN_IN), .ZN(n2727) );
  NAND2_X1 U3452 ( .A1(n3651), .A2(REG2_REG_27__SCAN_IN), .ZN(n2726) );
  INV_X1 U3453 ( .A(n2723), .ZN(n2721) );
  AOI21_X1 U3454 ( .B1(n2721), .B2(REG3_REG_26__SCAN_IN), .A(
        REG3_REG_27__SCAN_IN), .ZN(n2724) );
  NAND2_X1 U3455 ( .A1(REG3_REG_26__SCAN_IN), .A2(REG3_REG_27__SCAN_IN), .ZN(
        n2722) );
  NOR2_X1 U3456 ( .A1(n2723), .A2(n2722), .ZN(n2730) );
  OR2_X1 U3457 ( .A1(n2724), .A2(n2730), .ZN(n3942) );
  OR2_X1 U34580 ( .A1(n2222), .A2(n3942), .ZN(n2725) );
  INV_X1 U34590 ( .A(n3952), .ZN(n2924) );
  NOR2_X1 U3460 ( .A1(n2924), .A2(n3932), .ZN(n2729) );
  NAND2_X1 U3461 ( .A1(n2573), .A2(REG1_REG_28__SCAN_IN), .ZN(n2735) );
  NAND2_X1 U3462 ( .A1(n2720), .A2(REG0_REG_28__SCAN_IN), .ZN(n2734) );
  NAND2_X1 U3463 ( .A1(n3651), .A2(REG2_REG_28__SCAN_IN), .ZN(n2733) );
  NAND2_X1 U3464 ( .A1(n2730), .A2(REG3_REG_28__SCAN_IN), .ZN(n3909) );
  OR2_X1 U3465 ( .A1(n2730), .A2(REG3_REG_28__SCAN_IN), .ZN(n2731) );
  NAND2_X1 U3466 ( .A1(n3909), .A2(n2731), .ZN(n3523) );
  OR2_X1 U34670 ( .A1(n2222), .A2(n3523), .ZN(n2732) );
  OR2_X1 U3468 ( .A1(n3917), .A2(n3921), .ZN(n3911) );
  NAND2_X1 U34690 ( .A1(n3917), .A2(n3921), .ZN(n3792) );
  NAND2_X1 U3470 ( .A1(n3911), .A2(n3792), .ZN(n3919) );
  XNOR2_X1 U34710 ( .A(n3920), .B(n3919), .ZN(n3347) );
  NAND2_X1 U3472 ( .A1(n2739), .A2(n2738), .ZN(n2790) );
  NAND2_X1 U34730 ( .A1(n2742), .A2(n2741), .ZN(n2743) );
  XNOR2_X1 U3474 ( .A(n2973), .B(n2942), .ZN(n2748) );
  NAND2_X1 U34750 ( .A1(n2748), .A2(n3905), .ZN(n3301) );
  AND2_X1 U3476 ( .A1(n2821), .A2(n3897), .ZN(n2749) );
  NAND2_X1 U34770 ( .A1(n3078), .A2(n4545), .ZN(n3658) );
  OR2_X1 U3478 ( .A1(n3759), .A2(n3658), .ZN(n2751) );
  AND2_X1 U34790 ( .A1(n2751), .A2(n2750), .ZN(n2829) );
  NAND2_X1 U3480 ( .A1(n3067), .A2(n3090), .ZN(n3667) );
  NAND2_X1 U34810 ( .A1(n3824), .A2(n3098), .ZN(n3664) );
  INV_X1 U3482 ( .A(n3114), .ZN(n3110) );
  NAND2_X1 U34830 ( .A1(n3199), .A2(n3114), .ZN(n3684) );
  NAND2_X1 U3484 ( .A1(n3136), .A2(n3203), .ZN(n3685) );
  NOR2_X1 U34850 ( .A1(n3136), .A2(n3203), .ZN(n3672) );
  AOI21_X1 U3486 ( .B1(n3196), .B2(n3685), .A(n3672), .ZN(n3119) );
  AOI21_X1 U34870 ( .B1(n3119), .B2(n2754), .A(n3676), .ZN(n3153) );
  NOR2_X1 U3488 ( .A1(n3821), .A2(n3227), .ZN(n3679) );
  NAND2_X1 U34890 ( .A1(n3821), .A2(n3227), .ZN(n3152) );
  OAI21_X1 U3490 ( .B1(n3153), .B2(n3679), .A(n3152), .ZN(n3167) );
  AND2_X1 U34910 ( .A1(n3820), .A2(n3256), .ZN(n3165) );
  NAND2_X1 U3492 ( .A1(n3493), .A2(n3268), .ZN(n3678) );
  OAI21_X1 U34930 ( .B1(n3167), .B2(n3165), .A(n3678), .ZN(n3237) );
  NAND2_X1 U3494 ( .A1(n3819), .A2(n3351), .ZN(n3236) );
  NOR2_X1 U34950 ( .A1(n3819), .A2(n3351), .ZN(n3691) );
  AOI21_X1 U3496 ( .B1(n3237), .B2(n3236), .A(n3691), .ZN(n4488) );
  NAND2_X1 U34970 ( .A1(n4494), .A2(n3551), .ZN(n3293) );
  NAND2_X1 U3498 ( .A1(n3818), .A2(n3376), .ZN(n2755) );
  NAND2_X1 U34990 ( .A1(n3293), .A2(n2755), .ZN(n3700) );
  NAND2_X1 U3500 ( .A1(n3604), .A2(n3278), .ZN(n3292) );
  OAI22_X1 U35010 ( .A1(n3700), .A2(n3292), .B1(n3818), .B2(n3376), .ZN(n3702)
         );
  NAND2_X1 U3502 ( .A1(n4299), .A2(n3326), .ZN(n3697) );
  NAND2_X1 U35030 ( .A1(n3817), .A2(n4317), .ZN(n3683) );
  INV_X1 U3504 ( .A(n3683), .ZN(n2756) );
  AOI21_X1 U35050 ( .B1(n3324), .B2(n3322), .A(n2756), .ZN(n4141) );
  INV_X1 U35060 ( .A(n3783), .ZN(n2757) );
  NOR2_X1 U35070 ( .A1(n4300), .A2(n4124), .ZN(n3733) );
  AND2_X1 U35080 ( .A1(n4105), .A2(n4097), .ZN(n2758) );
  NOR2_X1 U35090 ( .A1(n4087), .A2(n2758), .ZN(n4011) );
  NAND2_X1 U35100 ( .A1(n4092), .A2(n4065), .ZN(n4013) );
  NAND2_X1 U35110 ( .A1(n3613), .A2(n4052), .ZN(n4015) );
  INV_X1 U35120 ( .A(n4015), .ZN(n2759) );
  INV_X1 U35130 ( .A(n4016), .ZN(n2767) );
  NOR2_X1 U35140 ( .A1(n2759), .A2(n2767), .ZN(n3789) );
  INV_X1 U35150 ( .A(n2760), .ZN(n4088) );
  NAND2_X1 U35160 ( .A1(n4300), .A2(n4124), .ZN(n3732) );
  NAND2_X1 U35170 ( .A1(n4088), .A2(n3732), .ZN(n2761) );
  NAND2_X1 U35180 ( .A1(n4011), .A2(n2761), .ZN(n2763) );
  INV_X1 U35190 ( .A(n4105), .ZN(n4078) );
  NAND2_X1 U35200 ( .A1(n4078), .A2(n4091), .ZN(n2762) );
  NAND2_X1 U35210 ( .A1(n2763), .A2(n2762), .ZN(n4070) );
  NOR2_X1 U35220 ( .A1(n4092), .A2(n4065), .ZN(n2764) );
  OR2_X1 U35230 ( .A1(n4070), .A2(n2764), .ZN(n4012) );
  NAND2_X1 U35240 ( .A1(n4012), .A2(n4013), .ZN(n3709) );
  AND2_X1 U35250 ( .A1(n4075), .A2(n3544), .ZN(n3710) );
  INV_X1 U35260 ( .A(n3710), .ZN(n3728) );
  INV_X1 U35270 ( .A(n2765), .ZN(n2766) );
  AOI21_X1 U35280 ( .B1(n4034), .B2(n3484), .A(n2766), .ZN(n3712) );
  OAI21_X1 U35290 ( .B1(n2767), .B2(n3728), .A(n3712), .ZN(n3790) );
  INV_X1 U35300 ( .A(n3790), .ZN(n2768) );
  NAND2_X1 U35310 ( .A1(n2769), .A2(n2768), .ZN(n3991) );
  NOR2_X1 U35320 ( .A1(n4021), .A2(n4001), .ZN(n3745) );
  NOR2_X1 U35330 ( .A1(n4034), .A2(n3484), .ZN(n3989) );
  NOR2_X1 U35340 ( .A1(n3745), .A2(n3989), .ZN(n3787) );
  NAND2_X1 U35350 ( .A1(n4021), .A2(n4001), .ZN(n3967) );
  NAND2_X1 U35360 ( .A1(n3996), .A2(n3979), .ZN(n3742) );
  AND2_X1 U35370 ( .A1(n3967), .A2(n3742), .ZN(n3798) );
  NOR2_X1 U35380 ( .A1(n3996), .A2(n3979), .ZN(n3744) );
  NAND2_X1 U35390 ( .A1(n3935), .A2(n2770), .ZN(n3656) );
  NAND2_X1 U35400 ( .A1(n3973), .A2(n3959), .ZN(n3714) );
  INV_X1 U35410 ( .A(n3714), .ZN(n3773) );
  NAND2_X1 U35420 ( .A1(n2924), .A2(n3941), .ZN(n3715) );
  NAND2_X1 U35430 ( .A1(n3952), .A2(n3932), .ZN(n3791) );
  NAND2_X1 U35440 ( .A1(n3715), .A2(n3791), .ZN(n3939) );
  INV_X1 U35450 ( .A(n3939), .ZN(n3931) );
  NAND2_X1 U35460 ( .A1(n3929), .A2(n3791), .ZN(n3912) );
  XOR2_X1 U35470 ( .A(n3919), .B(n3912), .Z(n2783) );
  NAND2_X1 U35480 ( .A1(n2942), .A2(n3897), .ZN(n2772) );
  INV_X1 U35490 ( .A(n2821), .ZN(n4284) );
  NAND2_X1 U35500 ( .A1(n2771), .A2(n4284), .ZN(n3805) );
  OR2_X1 U35510 ( .A1(n2773), .A2(n2794), .ZN(n2774) );
  OR2_X1 U35520 ( .A1(n2222), .A2(n3909), .ZN(n2778) );
  NAND2_X1 U35530 ( .A1(n2573), .A2(REG1_REG_29__SCAN_IN), .ZN(n2777) );
  NAND2_X1 U35540 ( .A1(n2501), .A2(REG0_REG_29__SCAN_IN), .ZN(n2776) );
  NAND2_X1 U35550 ( .A1(n3651), .A2(REG2_REG_29__SCAN_IN), .ZN(n2775) );
  NAND4_X1 U35560 ( .A1(n2778), .A2(n2777), .A3(n2776), .A4(n2775), .ZN(n3816)
         );
  NAND2_X1 U35570 ( .A1(n2936), .A2(n2981), .ZN(n4055) );
  AOI22_X1 U35580 ( .A1(n3816), .A2(n4495), .B1(n4162), .B2(n3921), .ZN(n2781)
         );
  OAI21_X1 U35590 ( .B1(n3952), .B2(n4491), .A(n2781), .ZN(n2782) );
  AOI21_X1 U35600 ( .B1(n2783), .B2(n4145), .A(n2782), .ZN(n3342) );
  OAI21_X1 U35610 ( .B1(n3347), .B2(n4580), .A(n3342), .ZN(n2825) );
  NOR2_X1 U35620 ( .A1(n2784), .A2(n2794), .ZN(n2785) );
  MUX2_X1 U35630 ( .A(n2794), .B(n2785), .S(IR_REG_25__SCAN_IN), .Z(n2786) );
  NAND2_X1 U35640 ( .A1(n2814), .A2(B_REG_SCAN_IN), .ZN(n2793) );
  NAND2_X1 U35650 ( .A1(n2810), .A2(n2811), .ZN(n2791) );
  MUX2_X1 U35660 ( .A(n2793), .B(B_REG_SCAN_IN), .S(n2809), .Z(n2796) );
  NOR2_X1 U35670 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_26__SCAN_IN), .ZN(n2800)
         );
  NOR4_X1 U35680 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_31__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2799) );
  NOR4_X1 U35690 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2798) );
  NOR4_X1 U35700 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2797) );
  AND4_X1 U35710 ( .A1(n2800), .A2(n2799), .A3(n2798), .A4(n2797), .ZN(n2806)
         );
  NOR4_X1 U35720 ( .A1(D_REG_9__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n2804) );
  NOR4_X1 U35730 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_11__SCAN_IN), .ZN(n2803) );
  NOR4_X1 U35740 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n2802) );
  NOR4_X1 U35750 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_19__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2801) );
  AND4_X1 U35760 ( .A1(n2804), .A2(n2803), .A3(n2802), .A4(n2801), .ZN(n2805)
         );
  NAND2_X1 U35770 ( .A1(n2806), .A2(n2805), .ZN(n2841) );
  NAND2_X1 U35780 ( .A1(n2821), .A2(n3905), .ZN(n2807) );
  NAND2_X1 U35790 ( .A1(n2936), .A2(n2807), .ZN(n2939) );
  NAND2_X1 U35800 ( .A1(n2939), .A2(n2847), .ZN(n2812) );
  INV_X1 U35810 ( .A(n2814), .ZN(n2861) );
  OR2_X1 U3582 ( .A1(n2812), .A2(n2956), .ZN(n2813) );
  AOI21_X1 U3583 ( .B1(n2845), .B2(n2841), .A(n2813), .ZN(n2816) );
  INV_X1 U3584 ( .A(n2859), .ZN(n2817) );
  NAND2_X1 U3585 ( .A1(n2817), .A2(n2814), .ZN(n2843) );
  OAI21_X1 U3586 ( .B1(n2865), .B2(D_REG_1__SCAN_IN), .A(n2843), .ZN(n2815) );
  INV_X1 U3587 ( .A(D_REG_0__SCAN_IN), .ZN(n4866) );
  INV_X1 U3588 ( .A(n2809), .ZN(n2818) );
  INV_X1 U3589 ( .A(n2819), .ZN(n2822) );
  NAND2_X1 U3590 ( .A1(n2979), .A2(n3011), .ZN(n2849) );
  NAND2_X1 U3591 ( .A1(n4504), .A2(n4503), .ZN(n4502) );
  NAND2_X1 U3592 ( .A1(n3329), .A2(n4317), .ZN(n4148) );
  NAND2_X1 U3593 ( .A1(n3940), .A2(n3921), .ZN(n2820) );
  NAND2_X1 U3594 ( .A1(n3924), .A2(n2820), .ZN(n3340) );
  NAND2_X1 U3595 ( .A1(n2822), .A2(n2440), .ZN(U3546) );
  INV_X1 U3596 ( .A(n2935), .ZN(n2824) );
  INV_X1 U3597 ( .A(n2826), .ZN(n2827) );
  NAND2_X1 U3598 ( .A1(n2827), .A2(n2439), .ZN(U3514) );
  XNOR2_X1 U3599 ( .A(n2752), .B(n2829), .ZN(n2830) );
  NAND2_X1 U3600 ( .A1(n2830), .A2(n4145), .ZN(n2840) );
  INV_X1 U3601 ( .A(n2752), .ZN(n2832) );
  NAND2_X1 U3602 ( .A1(n2833), .A2(n2832), .ZN(n2834) );
  NAND2_X1 U3603 ( .A1(n2831), .A2(n2834), .ZN(n4559) );
  INV_X1 U3604 ( .A(n3301), .ZN(n4500) );
  NAND2_X1 U3605 ( .A1(n4559), .A2(n4500), .ZN(n2839) );
  OAI22_X1 U3606 ( .A1(n3067), .A2(n4055), .B1(n4490), .B2(n2996), .ZN(n2837)
         );
  NOR2_X1 U3607 ( .A1(n2835), .A2(n4491), .ZN(n2836) );
  NOR2_X1 U3608 ( .A1(n2837), .A2(n2836), .ZN(n2838) );
  NAND3_X1 U3609 ( .A1(n2840), .A2(n2839), .A3(n2838), .ZN(n4557) );
  INV_X1 U3610 ( .A(n2841), .ZN(n2842) );
  NAND2_X1 U3611 ( .A1(n2842), .A2(D_REG_1__SCAN_IN), .ZN(n2844) );
  INV_X1 U3612 ( .A(n2843), .ZN(n2867) );
  AOI21_X1 U3613 ( .B1(n2845), .B2(n2844), .A(n2867), .ZN(n2934) );
  NAND3_X1 U3614 ( .A1(n2934), .A2(n2945), .A3(n2939), .ZN(n2846) );
  MUX2_X1 U3615 ( .A(n4557), .B(REG2_REG_2__SCAN_IN), .S(n4519), .Z(n2855) );
  AND2_X1 U3616 ( .A1(n4337), .A2(n3905), .ZN(n4118) );
  INV_X1 U3617 ( .A(n2849), .ZN(n3073) );
  NOR2_X1 U3618 ( .A1(n3073), .A2(n2996), .ZN(n4556) );
  NOR3_X1 U3619 ( .A1(n4135), .A2(n4555), .A3(n4556), .ZN(n2854) );
  INV_X1 U3620 ( .A(n4559), .ZN(n2852) );
  INV_X1 U3621 ( .A(n2973), .ZN(n2941) );
  NAND2_X1 U3622 ( .A1(n2941), .A2(n3897), .ZN(n3017) );
  INV_X1 U3623 ( .A(n3017), .ZN(n2850) );
  NAND2_X1 U3624 ( .A1(n4337), .A2(n2850), .ZN(n3308) );
  OAI22_X1 U3625 ( .A1(n2852), .A2(n3308), .B1(n2851), .B2(n4151), .ZN(n2853)
         );
  OR3_X1 U3626 ( .A1(n2855), .A2(n2854), .A3(n2853), .ZN(U3288) );
  MUX2_X1 U3627 ( .A(n2525), .B(n2903), .S(STATE_REG_SCAN_IN), .Z(n2856) );
  INV_X1 U3628 ( .A(n2856), .ZN(U3348) );
  MUX2_X1 U3629 ( .A(n2917), .B(n4881), .S(U3149), .Z(n2857) );
  INV_X1 U3630 ( .A(n2857), .ZN(U3342) );
  INV_X1 U3631 ( .A(n3893), .ZN(n3901) );
  NAND2_X1 U3632 ( .A1(n3901), .A2(STATE_REG_SCAN_IN), .ZN(n2858) );
  OAI21_X1 U3633 ( .B1(STATE_REG_SCAN_IN), .B2(n2658), .A(n2858), .ZN(U3334)
         );
  INV_X1 U3634 ( .A(DATAI_26_), .ZN(n4673) );
  NAND2_X1 U3635 ( .A1(n2859), .A2(STATE_REG_SCAN_IN), .ZN(n2860) );
  OAI21_X1 U3636 ( .B1(STATE_REG_SCAN_IN), .B2(n4673), .A(n2860), .ZN(U3326)
         );
  INV_X1 U3637 ( .A(DATAI_25_), .ZN(n2863) );
  NAND2_X1 U3638 ( .A1(n2861), .A2(STATE_REG_SCAN_IN), .ZN(n2862) );
  OAI21_X1 U3639 ( .B1(STATE_REG_SCAN_IN), .B2(n2863), .A(n2862), .ZN(U3327)
         );
  MUX2_X1 U3640 ( .A(n2669), .B(n3905), .S(STATE_REG_SCAN_IN), .Z(n2864) );
  INV_X1 U3641 ( .A(n2864), .ZN(U3333) );
  AOI22_X1 U3642 ( .A1(n4521), .A2(n4866), .B1(n2866), .B2(n4522), .ZN(U3458)
         );
  INV_X1 U3643 ( .A(D_REG_1__SCAN_IN), .ZN(n4821) );
  AOI22_X1 U3644 ( .A1(n4521), .A2(n4821), .B1(n2867), .B2(n4522), .ZN(U3459)
         );
  OR2_X1 U3645 ( .A1(n3026), .A2(U3149), .ZN(n3814) );
  NAND2_X1 U3646 ( .A1(n2956), .A2(n3814), .ZN(n2889) );
  INV_X1 U3647 ( .A(n3713), .ZN(n2868) );
  AOI21_X1 U3648 ( .B1(n2936), .B2(n3026), .A(n2868), .ZN(n2888) );
  INV_X1 U3649 ( .A(n2888), .ZN(n2869) );
  NOR2_X1 U3650 ( .A1(n4473), .A2(U4043), .ZN(U3148) );
  INV_X1 U3651 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n2871) );
  NAND2_X1 U3652 ( .A1(U4043), .A2(n3091), .ZN(n2870) );
  OAI21_X1 U3653 ( .B1(U4043), .B2(n2871), .A(n2870), .ZN(U3554) );
  INV_X1 U3654 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4832) );
  INV_X1 U3655 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4604) );
  INV_X1 U3656 ( .A(n2892), .ZN(n4539) );
  NOR2_X1 U3657 ( .A1(n4604), .A2(n4539), .ZN(n4377) );
  INV_X1 U3658 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4896) );
  AOI22_X1 U3659 ( .A1(n2893), .A2(REG1_REG_5__SCAN_IN), .B1(n4896), .B2(n4542), .ZN(n4365) );
  INV_X1 U3660 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2872) );
  MUX2_X1 U3661 ( .A(n2872), .B(REG1_REG_1__SCAN_IN), .S(n2894), .Z(n3826) );
  AND2_X1 U3662 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3827)
         );
  NAND2_X1 U3663 ( .A1(n3826), .A2(n3827), .ZN(n3847) );
  NAND2_X1 U3664 ( .A1(n4286), .A2(REG1_REG_1__SCAN_IN), .ZN(n3848) );
  INV_X1 U3665 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4852) );
  NAND2_X1 U3666 ( .A1(n4285), .A2(REG1_REG_2__SCAN_IN), .ZN(n2873) );
  NAND2_X1 U3667 ( .A1(n2875), .A2(n4294), .ZN(n2876) );
  NAND2_X1 U3668 ( .A1(REG1_REG_3__SCAN_IN), .A2(n4291), .ZN(n4290) );
  NAND2_X1 U3669 ( .A1(n2876), .A2(n4290), .ZN(n2877) );
  INV_X1 U3670 ( .A(n2903), .ZN(n4345) );
  XNOR2_X1 U3671 ( .A(n2877), .B(n4345), .ZN(n4346) );
  INV_X1 U3672 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2879) );
  INV_X1 U3673 ( .A(n2877), .ZN(n2878) );
  OAI22_X1 U3674 ( .A1(n4346), .A2(n2879), .B1(n2878), .B2(n2903), .ZN(n4364)
         );
  NAND2_X1 U3675 ( .A1(n4540), .A2(n2881), .ZN(n2882) );
  NAND2_X1 U3676 ( .A1(n2882), .A2(n4369), .ZN(n4378) );
  OAI22_X1 U3677 ( .A1(n4377), .A2(n4378), .B1(REG1_REG_7__SCAN_IN), .B2(n2892), .ZN(n2883) );
  NOR2_X1 U3678 ( .A1(n4537), .A2(n2883), .ZN(n2884) );
  INV_X1 U3679 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4390) );
  NAND2_X1 U3680 ( .A1(n4535), .A2(REG1_REG_9__SCAN_IN), .ZN(n2885) );
  OAI21_X1 U3681 ( .B1(n4535), .B2(REG1_REG_9__SCAN_IN), .A(n2885), .ZN(n4398)
         );
  AND2_X1 U3682 ( .A1(n4535), .A2(REG1_REG_9__SCAN_IN), .ZN(n2886) );
  INV_X1 U3683 ( .A(n2917), .ZN(n3857) );
  NAND2_X1 U3684 ( .A1(n2887), .A2(n3857), .ZN(n3872) );
  XNOR2_X1 U3685 ( .A(n2890), .B(IR_REG_27__SCAN_IN), .ZN(n4339) );
  INV_X1 U3686 ( .A(n4339), .ZN(n3833) );
  AOI211_X1 U3687 ( .C1(n4832), .C2(n2891), .A(n3873), .B(n4447), .ZN(n2919)
         );
  INV_X1 U3688 ( .A(n4458), .ZN(n4486) );
  NAND2_X1 U3689 ( .A1(n4535), .A2(REG2_REG_9__SCAN_IN), .ZN(n2912) );
  INV_X1 U3690 ( .A(n4535), .ZN(n4406) );
  AOI22_X1 U3691 ( .A1(n4535), .A2(REG2_REG_9__SCAN_IN), .B1(n3172), .B2(n4406), .ZN(n4403) );
  NAND2_X1 U3692 ( .A1(REG2_REG_7__SCAN_IN), .A2(n2892), .ZN(n2908) );
  INV_X1 U3693 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3125) );
  AOI22_X1 U3694 ( .A1(REG2_REG_7__SCAN_IN), .A2(n2892), .B1(n4539), .B2(n3125), .ZN(n4382) );
  INV_X1 U3695 ( .A(REG2_REG_5__SCAN_IN), .ZN(n4869) );
  AOI22_X1 U3696 ( .A1(n2893), .A2(REG2_REG_5__SCAN_IN), .B1(n4869), .B2(n4542), .ZN(n4359) );
  INV_X1 U3697 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2895) );
  AND2_X1 U3698 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3838)
         );
  NAND2_X1 U3699 ( .A1(n4286), .A2(REG2_REG_1__SCAN_IN), .ZN(n3842) );
  NAND2_X1 U3700 ( .A1(n3843), .A2(n3842), .ZN(n2898) );
  INV_X1 U3701 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2896) );
  MUX2_X1 U3702 ( .A(REG2_REG_2__SCAN_IN), .B(n2896), .S(n4285), .Z(n2897) );
  NAND2_X1 U3703 ( .A1(n4285), .A2(REG2_REG_2__SCAN_IN), .ZN(n2899) );
  NAND2_X1 U3704 ( .A1(n2900), .A2(n4294), .ZN(n2901) );
  NAND2_X1 U3705 ( .A1(n2901), .A2(n4292), .ZN(n2902) );
  XNOR2_X1 U3706 ( .A(n2902), .B(n4345), .ZN(n4348) );
  INV_X1 U3707 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2905) );
  INV_X1 U3708 ( .A(n2902), .ZN(n2904) );
  NAND2_X1 U3709 ( .A1(n4540), .A2(n2906), .ZN(n2907) );
  NAND2_X1 U3710 ( .A1(REG2_REG_6__SCAN_IN), .A2(n4372), .ZN(n4371) );
  NAND2_X1 U3711 ( .A1(n2909), .A2(n2910), .ZN(n2911) );
  NAND2_X1 U3712 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4394), .ZN(n4393) );
  NAND2_X1 U3713 ( .A1(n2911), .A2(n4393), .ZN(n4402) );
  NAND2_X1 U3714 ( .A1(n4403), .A2(n4402), .ZN(n4401) );
  NAND2_X1 U3715 ( .A1(n2912), .A2(n4401), .ZN(n3858) );
  XNOR2_X1 U3716 ( .A(n3858), .B(n2917), .ZN(n2913) );
  AND2_X1 U3717 ( .A1(n4287), .A2(n4339), .ZN(n3837) );
  NAND2_X1 U3718 ( .A1(REG2_REG_10__SCAN_IN), .A2(n2913), .ZN(n3859) );
  OAI211_X1 U3719 ( .C1(n2913), .C2(REG2_REG_10__SCAN_IN), .A(n4483), .B(n3859), .ZN(n2916) );
  NOR2_X1 U3720 ( .A1(STATE_REG_SCAN_IN), .A2(n2914), .ZN(n3495) );
  AOI21_X1 U3721 ( .B1(n4473), .B2(ADDR_REG_10__SCAN_IN), .A(n3495), .ZN(n2915) );
  OAI211_X1 U3722 ( .C1(n4486), .C2(n2917), .A(n2916), .B(n2915), .ZN(n2918)
         );
  OR2_X1 U3723 ( .A1(n2919), .A2(n2918), .ZN(U3250) );
  INV_X1 U3724 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n2921) );
  NAND2_X1 U3725 ( .A1(n4142), .A2(U4043), .ZN(n2920) );
  OAI21_X1 U3726 ( .B1(U4043), .B2(n2921), .A(n2920), .ZN(U3567) );
  INV_X1 U3727 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4803) );
  NAND2_X1 U3728 ( .A1(n2922), .A2(U4043), .ZN(n2923) );
  OAI21_X1 U3729 ( .B1(U4043), .B2(n4803), .A(n2923), .ZN(U3572) );
  INV_X1 U3730 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n2926) );
  NAND2_X1 U3731 ( .A1(n2924), .A2(U4043), .ZN(n2925) );
  OAI21_X1 U3732 ( .B1(U4043), .B2(n2926), .A(n2925), .ZN(U3577) );
  INV_X1 U3733 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n4817) );
  INV_X1 U3734 ( .A(n3917), .ZN(n3933) );
  NAND2_X1 U3735 ( .A1(n3933), .A2(U4043), .ZN(n2927) );
  OAI21_X1 U3736 ( .B1(U4043), .B2(n4817), .A(n2927), .ZN(U3578) );
  INV_X1 U3737 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n2929) );
  NAND2_X1 U3738 ( .A1(n3364), .A2(U4043), .ZN(n2928) );
  OAI21_X1 U3739 ( .B1(U4043), .B2(n2929), .A(n2928), .ZN(U3561) );
  INV_X1 U3740 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n4764) );
  NAND2_X1 U3741 ( .A1(n2995), .A2(U4043), .ZN(n2931) );
  OAI21_X1 U3742 ( .B1(U4043), .B2(n4764), .A(n2931), .ZN(U3552) );
  INV_X1 U3743 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n4772) );
  NAND2_X1 U3744 ( .A1(U4043), .A2(n4034), .ZN(n2932) );
  OAI21_X1 U3745 ( .B1(U4043), .B2(n4772), .A(n2932), .ZN(U3573) );
  INV_X1 U3746 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n4792) );
  NAND2_X1 U3747 ( .A1(n3044), .A2(U4043), .ZN(n2933) );
  OAI21_X1 U3748 ( .B1(U4043), .B2(n4792), .A(n2933), .ZN(U3555) );
  NAND2_X1 U3749 ( .A1(n2935), .A2(n2934), .ZN(n2957) );
  AOI21_X1 U3750 ( .B1(n4544), .B2(n3897), .A(n2936), .ZN(n2937) );
  NAND2_X1 U3751 ( .A1(n4490), .A2(n2937), .ZN(n2955) );
  NAND2_X1 U3752 ( .A1(n2955), .A2(n4490), .ZN(n2938) );
  NAND2_X1 U3753 ( .A1(n2957), .A2(n2938), .ZN(n2940) );
  NAND2_X1 U3754 ( .A1(n2940), .A2(n2939), .ZN(n3028) );
  INV_X1 U3755 ( .A(n3028), .ZN(n2946) );
  INV_X1 U3756 ( .A(n2974), .ZN(n2943) );
  NAND2_X1 U3757 ( .A1(n4522), .A2(n2943), .ZN(n2944) );
  NAND2_X1 U3758 ( .A1(n2957), .A2(n3811), .ZN(n3029) );
  NAND3_X1 U3759 ( .A1(n2946), .A2(n2945), .A3(n3029), .ZN(n3006) );
  INV_X1 U3760 ( .A(n3006), .ZN(n2961) );
  INV_X1 U3761 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2960) );
  INV_X1 U3762 ( .A(n3811), .ZN(n2947) );
  OR2_X1 U3763 ( .A1(n2957), .A2(n2947), .ZN(n2982) );
  OR2_X2 U3764 ( .A1(n2982), .A2(n4287), .ZN(n4315) );
  OR3_X1 U3765 ( .A1(n2957), .A2(n4490), .A3(n2956), .ZN(n2948) );
  INV_X1 U3766 ( .A(n3179), .ZN(n2949) );
  OAI22_X1 U3767 ( .A1(n3078), .A2(n3031), .B1(n3011), .B2(n3508), .ZN(n2976)
         );
  INV_X1 U3768 ( .A(n2976), .ZN(n2952) );
  INV_X1 U3769 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2951) );
  NAND2_X1 U3770 ( .A1(n2952), .A2(n2433), .ZN(n2972) );
  INV_X1 U3771 ( .A(n2950), .ZN(n2953) );
  AOI22_X1 U3772 ( .A1(n2949), .A2(n4545), .B1(n2953), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2954) );
  OAI21_X1 U3773 ( .B1(n3078), .B2(n3033), .A(n2954), .ZN(n2971) );
  XNOR2_X1 U3774 ( .A(n2972), .B(n2971), .ZN(n3834) );
  OAI22_X1 U3775 ( .A1(n4318), .A2(n3011), .B1(n3834), .B2(n4324), .ZN(n2958)
         );
  AOI21_X1 U3776 ( .B1(n3619), .B2(n2499), .A(n2958), .ZN(n2959) );
  OAI21_X1 U3777 ( .B1(n2961), .B2(n2960), .A(n2959), .ZN(U3229) );
  INV_X1 U3778 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n2963) );
  NAND2_X1 U3779 ( .A1(U4043), .A2(n4127), .ZN(n2962) );
  OAI21_X1 U3780 ( .B1(U4043), .B2(n2963), .A(n2962), .ZN(U3566) );
  INV_X1 U3781 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4823) );
  NAND2_X1 U3782 ( .A1(n2573), .A2(REG1_REG_30__SCAN_IN), .ZN(n2966) );
  NAND2_X1 U3783 ( .A1(n3651), .A2(REG2_REG_30__SCAN_IN), .ZN(n2965) );
  NAND2_X1 U3784 ( .A1(n2720), .A2(REG0_REG_30__SCAN_IN), .ZN(n2964) );
  NAND3_X1 U3785 ( .A1(n2966), .A2(n2965), .A3(n2964), .ZN(n3915) );
  NAND2_X1 U3786 ( .A1(U4043), .A2(n3915), .ZN(n2967) );
  OAI21_X1 U3787 ( .B1(U4043), .B2(n4823), .A(n2967), .ZN(U3580) );
  INV_X1 U3788 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n4766) );
  NAND2_X1 U3789 ( .A1(U4043), .A2(n4105), .ZN(n2968) );
  OAI21_X1 U3790 ( .B1(U4043), .B2(n4766), .A(n2968), .ZN(U3569) );
  INV_X1 U3791 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n2970) );
  NAND2_X1 U3792 ( .A1(U4043), .A2(n3136), .ZN(n2969) );
  OAI21_X1 U3793 ( .B1(U4043), .B2(n2970), .A(n2969), .ZN(U3556) );
  NAND2_X1 U3794 ( .A1(n2972), .A2(n2971), .ZN(n2978) );
  NAND2_X2 U3795 ( .A1(n2974), .A2(n2973), .ZN(n2975) );
  OR2_X1 U3796 ( .A1(n2976), .A2(n2975), .ZN(n2977) );
  NAND2_X1 U3797 ( .A1(n2978), .A2(n2977), .ZN(n2987) );
  OAI22_X1 U3798 ( .A1(n2835), .A2(n3179), .B1(n2979), .B2(n3508), .ZN(n2980)
         );
  XNOR2_X1 U3799 ( .A(n2980), .B(n3509), .ZN(n2989) );
  XNOR2_X1 U3800 ( .A(n2989), .B(n2990), .ZN(n2988) );
  XNOR2_X1 U3801 ( .A(n2987), .B(n2988), .ZN(n2985) );
  OR2_X2 U3802 ( .A1(n2982), .A2(n2981), .ZN(n4316) );
  INV_X1 U3803 ( .A(n4316), .ZN(n3620) );
  AOI22_X1 U3804 ( .A1(n3006), .A2(REG3_REG_1__SCAN_IN), .B1(n3620), .B2(n3825), .ZN(n2984) );
  AOI22_X1 U3805 ( .A1(n2491), .A2(n3638), .B1(n3619), .B2(n2995), .ZN(n2983)
         );
  OAI211_X1 U3806 ( .C1(n2985), .C2(n4324), .A(n2984), .B(n2983), .ZN(U3219)
         );
  INV_X1 U3807 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n4899) );
  NAND2_X1 U3808 ( .A1(n2499), .A2(U4043), .ZN(n2986) );
  OAI21_X1 U3809 ( .B1(U4043), .B2(n4899), .A(n2986), .ZN(U3551) );
  NAND2_X1 U3810 ( .A1(n2988), .A2(n2987), .ZN(n2993) );
  INV_X1 U3811 ( .A(n2989), .ZN(n2991) );
  NAND2_X1 U3812 ( .A1(n2991), .A2(n2990), .ZN(n2992) );
  NAND2_X1 U3813 ( .A1(n2993), .A2(n2992), .ZN(n3000) );
  NOR2_X1 U3814 ( .A1(n3031), .A2(n2996), .ZN(n2994) );
  AOI21_X1 U3815 ( .B1(n2995), .B2(n3455), .A(n2994), .ZN(n2999) );
  OAI22_X1 U3816 ( .A1(n3093), .A2(n3031), .B1(n2996), .B2(n3508), .ZN(n2997)
         );
  XNOR2_X1 U3817 ( .A(n2997), .B(n3509), .ZN(n2998) );
  NAND2_X1 U3818 ( .A1(n2998), .A2(n2999), .ZN(n3034) );
  OAI21_X1 U3819 ( .B1(n2999), .B2(n2998), .A(n3034), .ZN(n3004) );
  INV_X1 U3820 ( .A(n3000), .ZN(n3002) );
  INV_X1 U3821 ( .A(n3004), .ZN(n3001) );
  NAND2_X1 U3822 ( .A1(n3002), .A2(n3001), .ZN(n3035) );
  INV_X1 U3823 ( .A(n3035), .ZN(n3003) );
  AOI21_X1 U3824 ( .B1(n3000), .B2(n3004), .A(n3003), .ZN(n3009) );
  AOI22_X1 U3825 ( .A1(n3005), .A2(n3638), .B1(n3619), .B2(n3824), .ZN(n3008)
         );
  AOI22_X1 U3826 ( .A1(n3006), .A2(REG3_REG_2__SCAN_IN), .B1(n3620), .B2(n2499), .ZN(n3007) );
  OAI211_X1 U3827 ( .C1(n3009), .C2(n4324), .A(n3008), .B(n3007), .ZN(U3234)
         );
  INV_X1 U3828 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3835) );
  OR2_X1 U3829 ( .A1(n3078), .A2(n4545), .ZN(n3660) );
  NAND2_X1 U3830 ( .A1(n3660), .A2(n3658), .ZN(n4546) );
  NAND2_X1 U3831 ( .A1(n4514), .A2(n4546), .ZN(n3015) );
  AOI21_X1 U3832 ( .B1(n4544), .B2(n3905), .A(n4162), .ZN(n3012) );
  NAND2_X1 U3833 ( .A1(n3301), .A2(n4497), .ZN(n3010) );
  AOI22_X1 U3834 ( .A1(n4546), .A2(n3010), .B1(n4495), .B2(n2499), .ZN(n4548)
         );
  OAI21_X1 U3835 ( .B1(n3012), .B2(n3011), .A(n4548), .ZN(n3013) );
  INV_X1 U3836 ( .A(n4151), .ZN(n4508) );
  AOI22_X1 U3837 ( .A1(n3013), .A2(n4337), .B1(REG3_REG_0__SCAN_IN), .B2(n4508), .ZN(n3014) );
  OAI211_X1 U3838 ( .C1(n4337), .C2(n3835), .A(n3015), .B(n3014), .ZN(U3290)
         );
  NAND2_X1 U3839 ( .A1(n2240), .A2(n3684), .ZN(n3751) );
  XOR2_X1 U3840 ( .A(n3751), .B(n3016), .Z(n4570) );
  NAND2_X1 U3841 ( .A1(n3301), .A2(n3017), .ZN(n3018) );
  XOR2_X1 U3842 ( .A(n3751), .B(n3019), .Z(n3022) );
  OAI22_X1 U3843 ( .A1(n3187), .A2(n4055), .B1(n4490), .B2(n3110), .ZN(n3020)
         );
  AOI21_X1 U3844 ( .B1(n4126), .B2(n3091), .A(n3020), .ZN(n3021) );
  OAI21_X1 U3845 ( .B1(n3022), .B2(n4497), .A(n3021), .ZN(n4572) );
  NAND2_X1 U3846 ( .A1(n4572), .A2(n4337), .ZN(n3025) );
  AOI21_X1 U3847 ( .B1(n3114), .B2(n3049), .A(n3204), .ZN(n4573) );
  OAI22_X1 U3848 ( .A1(n4337), .A2(n4869), .B1(n3117), .B2(n4151), .ZN(n3023)
         );
  AOI21_X1 U3849 ( .B1(n4513), .B2(n4573), .A(n3023), .ZN(n3024) );
  OAI211_X1 U3850 ( .C1(n4570), .C2(n4155), .A(n3025), .B(n3024), .ZN(U3285)
         );
  NAND2_X1 U3851 ( .A1(n2950), .A2(n3026), .ZN(n3027) );
  OAI21_X1 U3852 ( .B1(n3028), .B2(n3027), .A(STATE_REG_SCAN_IN), .ZN(n3030)
         );
  OAI22_X1 U3853 ( .A1(n3067), .A2(n3447), .B1(n3098), .B2(n3508), .ZN(n3032)
         );
  XNOR2_X1 U3854 ( .A(n3032), .B(n3509), .ZN(n3057) );
  INV_X2 U3855 ( .A(n2949), .ZN(n3447) );
  OAI22_X1 U3856 ( .A1(n3067), .A2(n3448), .B1(n3098), .B2(n3447), .ZN(n3055)
         );
  XNOR2_X1 U3857 ( .A(n3057), .B(n3055), .ZN(n3037) );
  NAND2_X1 U3858 ( .A1(n3035), .A2(n3034), .ZN(n3036) );
  NAND2_X1 U3859 ( .A1(n3036), .A2(n3037), .ZN(n3064) );
  OAI21_X1 U3860 ( .B1(n3037), .B2(n3036), .A(n3064), .ZN(n3038) );
  NAND2_X1 U3861 ( .A1(n3038), .A2(n4309), .ZN(n3041) );
  INV_X1 U3862 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4811) );
  NOR2_X1 U3863 ( .A1(STATE_REG_SCAN_IN), .A2(n4811), .ZN(n4289) );
  INV_X1 U3864 ( .A(n3091), .ZN(n3112) );
  OAI22_X1 U3865 ( .A1(n3112), .A2(n4315), .B1(n4316), .B2(n3093), .ZN(n3039)
         );
  AOI211_X1 U3866 ( .C1(n3090), .C2(n3638), .A(n4289), .B(n3039), .ZN(n3040)
         );
  OAI211_X1 U3867 ( .C1(REG3_REG_3__SCAN_IN), .C2(n4331), .A(n3041), .B(n3040), 
        .ZN(U3215) );
  XNOR2_X1 U3868 ( .A(n3042), .B(n3758), .ZN(n3052) );
  XOR2_X1 U3869 ( .A(n3758), .B(n3043), .Z(n3047) );
  AOI22_X1 U3870 ( .A1(n3044), .A2(n4495), .B1(n4162), .B2(n3069), .ZN(n3045)
         );
  OAI21_X1 U3871 ( .B1(n3067), .B2(n4491), .A(n3045), .ZN(n3046) );
  AOI21_X1 U3872 ( .B1(n3047), .B2(n4145), .A(n3046), .ZN(n3048) );
  OAI21_X1 U3873 ( .B1(n3301), .B2(n3052), .A(n3048), .ZN(n4567) );
  INV_X1 U3874 ( .A(n3097), .ZN(n3050) );
  OAI211_X1 U3875 ( .C1(n3050), .C2(n3061), .A(n4585), .B(n3049), .ZN(n4566)
         );
  OAI22_X1 U3876 ( .A1(n4566), .A2(n3897), .B1(n4151), .B2(n3072), .ZN(n3051)
         );
  OAI21_X1 U3877 ( .B1(n4567), .B2(n3051), .A(n4337), .ZN(n3054) );
  INV_X1 U3878 ( .A(n3052), .ZN(n4569) );
  AOI22_X1 U3879 ( .A1(n4569), .A2(n4514), .B1(REG2_REG_4__SCAN_IN), .B2(n4519), .ZN(n3053) );
  NAND2_X1 U3880 ( .A1(n3054), .A2(n3053), .ZN(U3286) );
  INV_X1 U3881 ( .A(n3055), .ZN(n3056) );
  NAND2_X1 U3882 ( .A1(n3057), .A2(n3056), .ZN(n3062) );
  AND2_X1 U3883 ( .A1(n3064), .A2(n3062), .ZN(n3066) );
  NAND2_X1 U3884 ( .A1(n3091), .A2(n2949), .ZN(n3059) );
  OR2_X1 U3885 ( .A1(n3061), .A2(n3508), .ZN(n3058) );
  NAND2_X1 U3886 ( .A1(n3059), .A2(n3058), .ZN(n3060) );
  XNOR2_X1 U3887 ( .A(n3060), .B(n3509), .ZN(n3104) );
  OAI22_X1 U3888 ( .A1(n3112), .A2(n3448), .B1(n3031), .B2(n3061), .ZN(n3105)
         );
  XNOR2_X1 U3889 ( .A(n3104), .B(n3105), .ZN(n3065) );
  AND2_X1 U3890 ( .A1(n3065), .A2(n3062), .ZN(n3063) );
  OAI211_X1 U3891 ( .C1(n3066), .C2(n3065), .A(n4309), .B(n3108), .ZN(n3071)
         );
  INV_X1 U3892 ( .A(REG3_REG_4__SCAN_IN), .ZN(n4867) );
  NOR2_X1 U3893 ( .A1(STATE_REG_SCAN_IN), .A2(n4867), .ZN(n4350) );
  OAI22_X1 U3894 ( .A1(n3067), .A2(n4316), .B1(n4315), .B2(n3199), .ZN(n3068)
         );
  AOI211_X1 U3895 ( .C1(n3069), .C2(n3638), .A(n4350), .B(n3068), .ZN(n3070)
         );
  OAI211_X1 U3896 ( .C1(n4331), .C2(n3072), .A(n3071), .B(n3070), .ZN(U3227)
         );
  AOI21_X1 U3897 ( .B1(n4545), .B2(n2491), .A(n3073), .ZN(n4553) );
  OR2_X1 U3898 ( .A1(n3759), .A2(n3074), .ZN(n3075) );
  NAND2_X1 U3899 ( .A1(n3076), .A2(n3075), .ZN(n4550) );
  INV_X1 U3900 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3077) );
  OAI22_X1 U3901 ( .A1(n3308), .A2(n4550), .B1(n3077), .B2(n4151), .ZN(n3085)
         );
  OAI22_X1 U3902 ( .A1(n3093), .A2(n4055), .B1(n4490), .B2(n2979), .ZN(n3080)
         );
  NOR2_X1 U3903 ( .A1(n3078), .A2(n4491), .ZN(n3079) );
  NOR2_X1 U3904 ( .A1(n3080), .A2(n3079), .ZN(n3083) );
  XNOR2_X1 U3905 ( .A(n3759), .B(n3658), .ZN(n3081) );
  NAND2_X1 U3906 ( .A1(n3081), .A2(n4145), .ZN(n3082) );
  OAI211_X1 U3907 ( .C1(n4550), .C2(n3301), .A(n3083), .B(n3082), .ZN(n4551)
         );
  MUX2_X1 U3908 ( .A(REG2_REG_1__SCAN_IN), .B(n4551), .S(n4337), .Z(n3084) );
  AOI211_X1 U3909 ( .C1(n4513), .C2(n4553), .A(n3085), .B(n3084), .ZN(n3086)
         );
  INV_X1 U3910 ( .A(n3086), .ZN(U3289) );
  XNOR2_X1 U3911 ( .A(n3087), .B(n3760), .ZN(n4563) );
  OAI21_X1 U3912 ( .B1(n3760), .B2(n3089), .A(n3088), .ZN(n3095) );
  AOI22_X1 U3913 ( .A1(n3091), .A2(n4495), .B1(n3090), .B2(n4162), .ZN(n3092)
         );
  OAI21_X1 U3914 ( .B1(n3093), .B2(n4491), .A(n3092), .ZN(n3094) );
  AOI21_X1 U3915 ( .B1(n3095), .B2(n4145), .A(n3094), .ZN(n3096) );
  OAI21_X1 U3916 ( .B1(n4563), .B2(n3301), .A(n3096), .ZN(n4565) );
  INV_X1 U3917 ( .A(n4565), .ZN(n3103) );
  INV_X1 U3918 ( .A(n4563), .ZN(n3101) );
  OAI21_X1 U3919 ( .B1(n4555), .B2(n3098), .A(n3097), .ZN(n4561) );
  AOI22_X1 U3920 ( .A1(n4519), .A2(REG2_REG_3__SCAN_IN), .B1(n4508), .B2(n4811), .ZN(n3099) );
  OAI21_X1 U3921 ( .B1(n4135), .B2(n4561), .A(n3099), .ZN(n3100) );
  AOI21_X1 U3922 ( .B1(n4514), .B2(n3101), .A(n3100), .ZN(n3102) );
  OAI21_X1 U3923 ( .B1(n4519), .B2(n3103), .A(n3102), .ZN(U3287) );
  INV_X1 U3924 ( .A(n3104), .ZN(n3106) );
  NAND2_X1 U3925 ( .A1(n3106), .A2(n3105), .ZN(n3107) );
  OAI22_X1 U3926 ( .A1(n3199), .A2(n3447), .B1(n3110), .B2(n3508), .ZN(n3109)
         );
  XNOR2_X1 U3927 ( .A(n3109), .B(n3509), .ZN(n3132) );
  OAI22_X1 U3928 ( .A1(n3199), .A2(n3448), .B1(n3110), .B2(n3447), .ZN(n3133)
         );
  XNOR2_X1 U3929 ( .A(n3132), .B(n3133), .ZN(n3130) );
  XOR2_X1 U3930 ( .A(n3131), .B(n3130), .Z(n3111) );
  NAND2_X1 U3931 ( .A1(n3111), .A2(n4309), .ZN(n3116) );
  AND2_X1 U3932 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n4362) );
  OAI22_X1 U3933 ( .A1(n3112), .A2(n4316), .B1(n4315), .B2(n3187), .ZN(n3113)
         );
  AOI211_X1 U3934 ( .C1(n3114), .C2(n3638), .A(n4362), .B(n3113), .ZN(n3115)
         );
  OAI211_X1 U3935 ( .C1(n4331), .C2(n3117), .A(n3116), .B(n3115), .ZN(U3224)
         );
  XOR2_X1 U3936 ( .A(n3118), .B(n3757), .Z(n4578) );
  INV_X1 U3937 ( .A(n4578), .ZN(n3129) );
  XOR2_X1 U3938 ( .A(n3757), .B(n3119), .Z(n3122) );
  OAI22_X1 U3939 ( .A1(n3266), .A2(n4055), .B1(n4490), .B2(n3181), .ZN(n3120)
         );
  AOI21_X1 U3940 ( .B1(n4126), .B2(n3136), .A(n3120), .ZN(n3121) );
  OAI21_X1 U3941 ( .B1(n3122), .B2(n4497), .A(n3121), .ZN(n4575) );
  NAND2_X1 U3942 ( .A1(n4575), .A2(n4337), .ZN(n3128) );
  INV_X1 U3943 ( .A(n3206), .ZN(n3124) );
  INV_X1 U3944 ( .A(n4585), .ZN(n4587) );
  INV_X1 U3945 ( .A(n3158), .ZN(n3123) );
  AOI211_X1 U3946 ( .C1(n3190), .C2(n3124), .A(n4587), .B(n3123), .ZN(n4576)
         );
  OAI22_X1 U3947 ( .A1(n4337), .A2(n3125), .B1(n3193), .B2(n4151), .ZN(n3126)
         );
  AOI21_X1 U3948 ( .B1(n4576), .B2(n4118), .A(n3126), .ZN(n3127) );
  OAI211_X1 U3949 ( .C1(n3129), .C2(n4155), .A(n3128), .B(n3127), .ZN(U3283)
         );
  INV_X1 U3950 ( .A(n3132), .ZN(n3134) );
  NAND2_X1 U3951 ( .A1(n3134), .A2(n3133), .ZN(n3135) );
  NAND2_X1 U3952 ( .A1(n3136), .A2(n3443), .ZN(n3138) );
  OR2_X1 U3953 ( .A1(n3203), .A2(n3508), .ZN(n3137) );
  NAND2_X1 U3954 ( .A1(n3138), .A2(n3137), .ZN(n3139) );
  XNOR2_X1 U3955 ( .A(n3139), .B(n2975), .ZN(n3140) );
  OAI22_X1 U3956 ( .A1(n3187), .A2(n3448), .B1(n3203), .B2(n3447), .ZN(n3141)
         );
  AND2_X1 U3957 ( .A1(n3140), .A2(n3141), .ZN(n3177) );
  INV_X1 U3958 ( .A(n3177), .ZN(n3144) );
  INV_X1 U3959 ( .A(n3140), .ZN(n3143) );
  INV_X1 U3960 ( .A(n3141), .ZN(n3142) );
  NAND2_X1 U3961 ( .A1(n3143), .A2(n3142), .ZN(n3176) );
  NAND2_X1 U3962 ( .A1(n3144), .A2(n3176), .ZN(n3145) );
  XNOR2_X1 U3963 ( .A(n3178), .B(n3145), .ZN(n3146) );
  NAND2_X1 U3964 ( .A1(n3146), .A2(n4309), .ZN(n3150) );
  NOR2_X1 U3965 ( .A1(STATE_REG_SCAN_IN), .A2(n3147), .ZN(n4368) );
  OAI22_X1 U3966 ( .A1(n3199), .A2(n4316), .B1(n4315), .B2(n3230), .ZN(n3148)
         );
  AOI211_X1 U3967 ( .C1(n3197), .C2(n3638), .A(n4368), .B(n3148), .ZN(n3149)
         );
  OAI211_X1 U3968 ( .C1(n4331), .C2(n3151), .A(n3150), .B(n3149), .ZN(U3236)
         );
  INV_X1 U3969 ( .A(n3152), .ZN(n3677) );
  OR2_X1 U3970 ( .A1(n3677), .A2(n3679), .ZN(n3753) );
  XNOR2_X1 U3971 ( .A(n3153), .B(n3753), .ZN(n3156) );
  OAI22_X1 U3972 ( .A1(n3493), .A2(n4055), .B1(n4490), .B2(n3227), .ZN(n3154)
         );
  AOI21_X1 U3973 ( .B1(n4126), .B2(n3823), .A(n3154), .ZN(n3155) );
  OAI21_X1 U3974 ( .B1(n3156), .B2(n4497), .A(n3155), .ZN(n3213) );
  INV_X1 U3975 ( .A(n3213), .ZN(n3164) );
  XNOR2_X1 U3976 ( .A(n3157), .B(n3753), .ZN(n3214) );
  NAND2_X1 U3977 ( .A1(n3158), .A2(n3232), .ZN(n3159) );
  NAND2_X1 U3978 ( .A1(n2254), .A2(n3159), .ZN(n3219) );
  NOR2_X1 U3979 ( .A1(n4135), .A2(n3219), .ZN(n3162) );
  INV_X1 U3980 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3160) );
  OAI22_X1 U3981 ( .A1(n4337), .A2(n3160), .B1(n3235), .B2(n4151), .ZN(n3161)
         );
  AOI211_X1 U3982 ( .C1(n3214), .C2(n4068), .A(n3162), .B(n3161), .ZN(n3163)
         );
  OAI21_X1 U3983 ( .B1(n3164), .B2(n4519), .A(n3163), .ZN(U3282) );
  INV_X1 U3984 ( .A(n3165), .ZN(n3692) );
  NAND2_X1 U3985 ( .A1(n3692), .A2(n3678), .ZN(n3752) );
  XNOR2_X1 U3986 ( .A(n3166), .B(n3752), .ZN(n4581) );
  XOR2_X1 U3987 ( .A(n3752), .B(n3167), .Z(n3170) );
  OAI22_X1 U3988 ( .A1(n4492), .A2(n4055), .B1(n4490), .B2(n3256), .ZN(n3168)
         );
  AOI21_X1 U3989 ( .B1(n4126), .B2(n3821), .A(n3168), .ZN(n3169) );
  OAI21_X1 U3990 ( .B1(n3170), .B2(n4497), .A(n3169), .ZN(n4582) );
  NAND2_X1 U3991 ( .A1(n4582), .A2(n4337), .ZN(n3175) );
  INV_X1 U3992 ( .A(n3171), .ZN(n3243) );
  AOI21_X1 U3993 ( .B1(n3268), .B2(n2254), .A(n3243), .ZN(n4584) );
  INV_X1 U3994 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3172) );
  OAI22_X1 U3995 ( .A1(n4337), .A2(n3172), .B1(n3269), .B2(n4151), .ZN(n3173)
         );
  AOI21_X1 U3996 ( .B1(n4584), .B2(n4513), .A(n3173), .ZN(n3174) );
  OAI211_X1 U3997 ( .C1(n4581), .C2(n4155), .A(n3175), .B(n3174), .ZN(U3281)
         );
  OAI21_X1 U3998 ( .B1(n3178), .B2(n3177), .A(n3176), .ZN(n3182) );
  OAI22_X1 U3999 ( .A1(n3230), .A2(n3511), .B1(n3508), .B2(n3181), .ZN(n3180)
         );
  XNOR2_X1 U4000 ( .A(n3180), .B(n2975), .ZN(n3221) );
  OAI22_X1 U4001 ( .A1(n3230), .A2(n3448), .B1(n3511), .B2(n3181), .ZN(n3220)
         );
  XNOR2_X1 U4002 ( .A(n3221), .B(n3220), .ZN(n3183) );
  AOI21_X1 U4003 ( .B1(n3182), .B2(n3183), .A(n4324), .ZN(n3186) );
  INV_X1 U4004 ( .A(n3182), .ZN(n3185) );
  NAND2_X1 U4005 ( .A1(n3185), .A2(n3184), .ZN(n3223) );
  NAND2_X1 U4006 ( .A1(n3186), .A2(n3223), .ZN(n3192) );
  NAND2_X1 U4007 ( .A1(REG3_REG_7__SCAN_IN), .A2(U3149), .ZN(n4384) );
  INV_X1 U4008 ( .A(n4384), .ZN(n3189) );
  OAI22_X1 U4009 ( .A1(n3187), .A2(n4316), .B1(n4315), .B2(n3266), .ZN(n3188)
         );
  AOI211_X1 U4010 ( .C1(n3190), .C2(n3638), .A(n3189), .B(n3188), .ZN(n3191)
         );
  OAI211_X1 U4011 ( .C1(n4331), .C2(n3193), .A(n3192), .B(n3191), .ZN(U3210)
         );
  INV_X1 U4012 ( .A(n3685), .ZN(n3195) );
  OR2_X1 U4013 ( .A1(n3195), .A2(n3672), .ZN(n3761) );
  XNOR2_X1 U4014 ( .A(n3194), .B(n3761), .ZN(n4510) );
  XOR2_X1 U4015 ( .A(n3761), .B(n3196), .Z(n3202) );
  AOI22_X1 U4016 ( .A1(n3823), .A2(n4495), .B1(n4162), .B2(n3197), .ZN(n3198)
         );
  OAI21_X1 U4017 ( .B1(n3199), .B2(n4491), .A(n3198), .ZN(n3201) );
  NOR2_X1 U4018 ( .A1(n4510), .A2(n3301), .ZN(n3200) );
  AOI211_X1 U4019 ( .C1(n3202), .C2(n4145), .A(n3201), .B(n3200), .ZN(n4518)
         );
  OAI21_X1 U4020 ( .B1(n4510), .B2(n4562), .A(n4518), .ZN(n3211) );
  NOR2_X1 U4021 ( .A1(n3204), .A2(n3203), .ZN(n3205) );
  OR2_X1 U4022 ( .A1(n3206), .A2(n3205), .ZN(n4511) );
  INV_X1 U4023 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3207) );
  OAI22_X1 U4024 ( .A1(n4511), .A2(n4281), .B1(n4596), .B2(n3207), .ZN(n3208)
         );
  AOI21_X1 U4025 ( .B1(n3211), .B2(n4596), .A(n3208), .ZN(n3209) );
  INV_X1 U4026 ( .A(n3209), .ZN(U3479) );
  INV_X1 U4027 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4840) );
  OAI22_X1 U4028 ( .A1(n4511), .A2(n4237), .B1(n4610), .B2(n4840), .ZN(n3210)
         );
  AOI21_X1 U4029 ( .B1(n3211), .B2(n4610), .A(n3210), .ZN(n3212) );
  INV_X1 U4030 ( .A(n3212), .ZN(U3524) );
  AOI21_X1 U4031 ( .B1(n3214), .B2(n4577), .A(n3213), .ZN(n3216) );
  MUX2_X1 U4032 ( .A(n4390), .B(n3216), .S(n4610), .Z(n3215) );
  OAI21_X1 U4033 ( .B1(n3219), .B2(n4237), .A(n3215), .ZN(U3526) );
  INV_X1 U4034 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3217) );
  MUX2_X1 U4035 ( .A(n3217), .B(n3216), .S(n4596), .Z(n3218) );
  OAI21_X1 U4036 ( .B1(n3219), .B2(n4281), .A(n3218), .ZN(U3483) );
  NAND2_X1 U4037 ( .A1(n3221), .A2(n3220), .ZN(n3222) );
  NAND2_X1 U4038 ( .A1(n3821), .A2(n3443), .ZN(n3225) );
  OR2_X1 U4039 ( .A1(n3227), .A2(n3508), .ZN(n3224) );
  NAND2_X1 U4040 ( .A1(n3225), .A2(n3224), .ZN(n3226) );
  XNOR2_X1 U4041 ( .A(n3226), .B(n2975), .ZN(n3257) );
  OAI22_X1 U4042 ( .A1(n3266), .A2(n3448), .B1(n3227), .B2(n3447), .ZN(n3258)
         );
  XNOR2_X1 U40430 ( .A(n3257), .B(n3258), .ZN(n3228) );
  XNOR2_X1 U4044 ( .A(n3259), .B(n3228), .ZN(n3229) );
  NAND2_X1 U4045 ( .A1(n3229), .A2(n4309), .ZN(n3234) );
  INV_X1 U4046 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4833) );
  NOR2_X1 U4047 ( .A1(STATE_REG_SCAN_IN), .A2(n4833), .ZN(n4391) );
  OAI22_X1 U4048 ( .A1(n3230), .A2(n4316), .B1(n4315), .B2(n3493), .ZN(n3231)
         );
  AOI211_X1 U4049 ( .C1(n3232), .C2(n3638), .A(n4391), .B(n3231), .ZN(n3233)
         );
  OAI211_X1 U4050 ( .C1(n4331), .C2(n3235), .A(n3234), .B(n3233), .ZN(U3218)
         );
  INV_X1 U4051 ( .A(n3236), .ZN(n3694) );
  OR2_X1 U4052 ( .A1(n3694), .A2(n3691), .ZN(n3754) );
  XNOR2_X1 U4053 ( .A(n3237), .B(n3754), .ZN(n3240) );
  OAI22_X1 U4054 ( .A1(n3552), .A2(n4055), .B1(n4490), .B2(n3351), .ZN(n3238)
         );
  AOI21_X1 U4055 ( .B1(n4126), .B2(n3820), .A(n3238), .ZN(n3239) );
  OAI21_X1 U4056 ( .B1(n3240), .B2(n4497), .A(n3239), .ZN(n3249) );
  INV_X1 U4057 ( .A(n3249), .ZN(n3248) );
  XNOR2_X1 U4058 ( .A(n3241), .B(n3754), .ZN(n3250) );
  INV_X1 U4059 ( .A(n4504), .ZN(n3242) );
  OAI21_X1 U4060 ( .B1(n3243), .B2(n3351), .A(n3242), .ZN(n3254) );
  NOR2_X1 U4061 ( .A1(n3254), .A2(n4135), .ZN(n3246) );
  INV_X1 U4062 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3244) );
  OAI22_X1 U4063 ( .A1(n4337), .A2(n3244), .B1(n3499), .B2(n4151), .ZN(n3245)
         );
  AOI211_X1 U4064 ( .C1(n3250), .C2(n4068), .A(n3246), .B(n3245), .ZN(n3247)
         );
  OAI21_X1 U4065 ( .B1(n3248), .B2(n4519), .A(n3247), .ZN(U3280) );
  AOI21_X1 U4066 ( .B1(n3250), .B2(n4577), .A(n3249), .ZN(n3252) );
  MUX2_X1 U4067 ( .A(n4832), .B(n3252), .S(n4610), .Z(n3251) );
  OAI21_X1 U4068 ( .B1(n3254), .B2(n4237), .A(n3251), .ZN(U3528) );
  INV_X1 U4069 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4714) );
  MUX2_X1 U4070 ( .A(n4714), .B(n3252), .S(n4596), .Z(n3253) );
  OAI21_X1 U4071 ( .B1(n3254), .B2(n4281), .A(n3253), .ZN(U3487) );
  OAI22_X1 U4072 ( .A1(n3493), .A2(n3511), .B1(n3256), .B2(n3508), .ZN(n3255)
         );
  XNOR2_X1 U4073 ( .A(n3255), .B(n2975), .ZN(n3352) );
  OAI22_X1 U4074 ( .A1(n3493), .A2(n3448), .B1(n3256), .B2(n3447), .ZN(n3353)
         );
  XNOR2_X1 U4075 ( .A(n3352), .B(n3353), .ZN(n3265) );
  OAI21_X1 U4076 ( .B1(n3259), .B2(n3258), .A(n3257), .ZN(n3261) );
  NAND2_X1 U4077 ( .A1(n3259), .A2(n3258), .ZN(n3260) );
  INV_X1 U4078 ( .A(n3265), .ZN(n3263) );
  INV_X1 U4079 ( .A(n3357), .ZN(n3264) );
  AOI21_X1 U4080 ( .B1(n3265), .B2(n3262), .A(n3264), .ZN(n3273) );
  AND2_X1 U4081 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4399) );
  OAI22_X1 U4082 ( .A1(n3266), .A2(n4316), .B1(n4315), .B2(n4492), .ZN(n3267)
         );
  AOI211_X1 U4083 ( .C1(n3268), .C2(n3638), .A(n4399), .B(n3267), .ZN(n3272)
         );
  INV_X1 U4084 ( .A(n3269), .ZN(n3270) );
  NAND2_X1 U4085 ( .A1(n3648), .A2(n3270), .ZN(n3271) );
  OAI211_X1 U4086 ( .C1(n3273), .C2(n4324), .A(n3272), .B(n3271), .ZN(U3228)
         );
  NAND2_X1 U4087 ( .A1(n3292), .A2(n3293), .ZN(n3755) );
  XNOR2_X1 U4088 ( .A(n3295), .B(n3755), .ZN(n3276) );
  OAI22_X1 U4089 ( .A1(n2618), .A2(n4055), .B1(n4490), .B2(n3551), .ZN(n3274)
         );
  AOI21_X1 U4090 ( .B1(n4126), .B2(n3364), .A(n3274), .ZN(n3275) );
  OAI21_X1 U4091 ( .B1(n3276), .B2(n4497), .A(n3275), .ZN(n3285) );
  INV_X1 U4092 ( .A(n3285), .ZN(n3284) );
  XOR2_X1 U4093 ( .A(n3755), .B(n3277), .Z(n3286) );
  NAND2_X1 U4094 ( .A1(n4502), .A2(n3278), .ZN(n3279) );
  NAND2_X1 U4095 ( .A1(n3302), .A2(n3279), .ZN(n3290) );
  INV_X1 U4096 ( .A(n3280), .ZN(n3555) );
  AOI22_X1 U4097 ( .A1(n4519), .A2(REG2_REG_12__SCAN_IN), .B1(n3555), .B2(
        n4508), .ZN(n3281) );
  OAI21_X1 U4098 ( .B1(n3290), .B2(n4135), .A(n3281), .ZN(n3282) );
  AOI21_X1 U4099 ( .B1(n3286), .B2(n4068), .A(n3282), .ZN(n3283) );
  OAI21_X1 U4100 ( .B1(n4519), .B2(n3284), .A(n3283), .ZN(U3278) );
  INV_X1 U4101 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4419) );
  AOI21_X1 U4102 ( .B1(n3286), .B2(n4577), .A(n3285), .ZN(n3288) );
  MUX2_X1 U4103 ( .A(n4419), .B(n3288), .S(n4610), .Z(n3287) );
  OAI21_X1 U4104 ( .B1(n3290), .B2(n4237), .A(n3287), .ZN(U3530) );
  INV_X1 U4105 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4713) );
  MUX2_X1 U4106 ( .A(n4713), .B(n3288), .S(n4596), .Z(n3289) );
  OAI21_X1 U4107 ( .B1(n3290), .B2(n4281), .A(n3289), .ZN(U3491) );
  XNOR2_X1 U4108 ( .A(n3818), .B(n3606), .ZN(n3764) );
  XNOR2_X1 U4109 ( .A(n3291), .B(n3764), .ZN(n4232) );
  OAI22_X1 U4110 ( .A1(n4989), .A2(n4055), .B1(n4490), .B2(n3376), .ZN(n3299)
         );
  INV_X1 U4111 ( .A(n3292), .ZN(n3294) );
  OAI21_X1 U4112 ( .B1(n3295), .B2(n3294), .A(n3293), .ZN(n3296) );
  XNOR2_X1 U4113 ( .A(n3296), .B(n3764), .ZN(n3297) );
  NOR2_X1 U4114 ( .A1(n3297), .A2(n4497), .ZN(n3298) );
  AOI211_X1 U4115 ( .C1(n4126), .C2(n4494), .A(n3299), .B(n3298), .ZN(n3300)
         );
  OAI21_X1 U4116 ( .B1(n3301), .B2(n4232), .A(n3300), .ZN(n4233) );
  NAND2_X1 U4117 ( .A1(n4233), .A2(n4337), .ZN(n3307) );
  OAI21_X1 U4118 ( .B1(n2271), .B2(n3376), .A(n2228), .ZN(n4282) );
  INV_X1 U4119 ( .A(n4282), .ZN(n3305) );
  INV_X1 U4120 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3303) );
  OAI22_X1 U4121 ( .A1(n4337), .A2(n3303), .B1(n3609), .B2(n4151), .ZN(n3304)
         );
  AOI21_X1 U4122 ( .B1(n3305), .B2(n4513), .A(n3304), .ZN(n3306) );
  OAI211_X1 U4123 ( .C1(n4232), .C2(n3308), .A(n3307), .B(n3306), .ZN(U3277)
         );
  OAI21_X1 U4124 ( .B1(n3309), .B2(n3762), .A(n3311), .ZN(n4226) );
  AOI21_X1 U4125 ( .B1(n3777), .B2(n3762), .A(n3312), .ZN(n3315) );
  OAI22_X1 U4126 ( .A1(n4299), .A2(n4055), .B1(n4490), .B2(n3472), .ZN(n3313)
         );
  AOI21_X1 U4127 ( .B1(n4126), .B2(n3818), .A(n3313), .ZN(n3314) );
  OAI21_X1 U4128 ( .B1(n3315), .B2(n4497), .A(n3314), .ZN(n3316) );
  AOI21_X1 U4129 ( .B1(n4500), .B2(n4226), .A(n3316), .ZN(n4230) );
  INV_X1 U4130 ( .A(n3329), .ZN(n4228) );
  NAND2_X1 U4131 ( .A1(n2228), .A2(n3317), .ZN(n4227) );
  AND3_X1 U4132 ( .A1(n4228), .A2(n4513), .A3(n4227), .ZN(n3320) );
  INV_X1 U4133 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3318) );
  OAI22_X1 U4134 ( .A1(n4337), .A2(n3318), .B1(n3471), .B2(n4151), .ZN(n3319)
         );
  AOI211_X1 U4135 ( .C1(n4226), .C2(n4514), .A(n3320), .B(n3319), .ZN(n3321)
         );
  OAI21_X1 U4136 ( .B1(n4230), .B2(n4519), .A(n3321), .ZN(U3276) );
  XNOR2_X1 U4137 ( .A(n3323), .B(n3763), .ZN(n4223) );
  INV_X1 U4138 ( .A(n4223), .ZN(n3335) );
  XNOR2_X1 U4139 ( .A(n3324), .B(n3763), .ZN(n3325) );
  NAND2_X1 U4140 ( .A1(n3325), .A2(n4145), .ZN(n3328) );
  AOI22_X1 U4141 ( .A1(n4127), .A2(n4495), .B1(n4162), .B2(n3326), .ZN(n3327)
         );
  OAI211_X1 U4142 ( .C1(n4989), .C2(n4491), .A(n3328), .B(n3327), .ZN(n4222)
         );
  OR2_X1 U4143 ( .A1(n3329), .A2(n4317), .ZN(n3330) );
  NAND2_X1 U4144 ( .A1(n4148), .A2(n3330), .ZN(n4276) );
  NOR2_X1 U4145 ( .A1(n4276), .A2(n4135), .ZN(n3333) );
  INV_X1 U4146 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3331) );
  OAI22_X1 U4147 ( .A1(n4337), .A2(n3331), .B1(n4330), .B2(n4151), .ZN(n3332)
         );
  AOI211_X1 U4148 ( .C1(n4222), .C2(n4337), .A(n3333), .B(n3332), .ZN(n3334)
         );
  OAI21_X1 U4149 ( .B1(n3335), .B2(n4155), .A(n3334), .ZN(U3275) );
  NAND3_X1 U4150 ( .A1(n3337), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3339) );
  INV_X1 U4151 ( .A(DATAI_31_), .ZN(n3338) );
  OAI22_X1 U4152 ( .A1(n3336), .A2(n3339), .B1(STATE_REG_SCAN_IN), .B2(n3338), 
        .ZN(U3321) );
  INV_X1 U4153 ( .A(n3340), .ZN(n3345) );
  INV_X1 U4154 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3341) );
  OAI22_X1 U4155 ( .A1(n4337), .A2(n3341), .B1(n3523), .B2(n4151), .ZN(n3344)
         );
  NOR2_X1 U4156 ( .A1(n3342), .A2(n4519), .ZN(n3343) );
  AOI211_X1 U4157 ( .C1(n4513), .C2(n3345), .A(n3344), .B(n3343), .ZN(n3346)
         );
  OAI21_X1 U4158 ( .B1(n3347), .B2(n4155), .A(n3346), .ZN(U3262) );
  NAND2_X1 U4159 ( .A1(n3819), .A2(n3443), .ZN(n3349) );
  OR2_X1 U4160 ( .A1(n3351), .A2(n3508), .ZN(n3348) );
  NAND2_X1 U4161 ( .A1(n3349), .A2(n3348), .ZN(n3350) );
  XNOR2_X1 U4162 ( .A(n3350), .B(n3509), .ZN(n3358) );
  OAI22_X1 U4163 ( .A1(n4492), .A2(n3448), .B1(n3511), .B2(n3351), .ZN(n3359)
         );
  XNOR2_X1 U4164 ( .A(n3358), .B(n3359), .ZN(n3491) );
  INV_X1 U4165 ( .A(n3352), .ZN(n3355) );
  INV_X1 U4166 ( .A(n3353), .ZN(n3354) );
  NAND2_X1 U4167 ( .A1(n3355), .A2(n3354), .ZN(n3489) );
  AND2_X1 U4168 ( .A1(n3491), .A2(n3489), .ZN(n3356) );
  INV_X1 U4169 ( .A(n3358), .ZN(n3360) );
  NAND2_X1 U4170 ( .A1(n3360), .A2(n3359), .ZN(n3361) );
  NAND2_X1 U4171 ( .A1(n3490), .A2(n3361), .ZN(n3623) );
  OAI22_X1 U4172 ( .A1(n3552), .A2(n3511), .B1(n4503), .B2(n3508), .ZN(n3362)
         );
  XNOR2_X1 U4173 ( .A(n3362), .B(n3509), .ZN(n3365) );
  NOR2_X1 U4174 ( .A1(n3511), .A2(n4503), .ZN(n3363) );
  AOI21_X1 U4175 ( .B1(n3364), .B2(n3455), .A(n3363), .ZN(n3366) );
  NAND2_X1 U4176 ( .A1(n3365), .A2(n3366), .ZN(n3624) );
  NAND2_X1 U4177 ( .A1(n3623), .A2(n3624), .ZN(n3622) );
  INV_X1 U4178 ( .A(n3365), .ZN(n3368) );
  INV_X1 U4179 ( .A(n3366), .ZN(n3367) );
  NAND2_X1 U4180 ( .A1(n3368), .A2(n3367), .ZN(n3626) );
  NAND2_X1 U4181 ( .A1(n3622), .A2(n3626), .ZN(n3549) );
  NAND2_X1 U4182 ( .A1(n4494), .A2(n3443), .ZN(n3370) );
  OR2_X1 U4183 ( .A1(n3551), .A2(n3508), .ZN(n3369) );
  NAND2_X1 U4184 ( .A1(n3370), .A2(n3369), .ZN(n3371) );
  XNOR2_X1 U4185 ( .A(n3371), .B(n3509), .ZN(n3595) );
  NOR2_X1 U4186 ( .A1(n3511), .A2(n3551), .ZN(n3372) );
  AOI21_X1 U4187 ( .B1(n3455), .B2(n4494), .A(n3372), .ZN(n3597) );
  INV_X2 U4188 ( .A(n3447), .ZN(n3443) );
  NAND2_X1 U4189 ( .A1(n3818), .A2(n3443), .ZN(n3374) );
  OR2_X1 U4190 ( .A1(n3376), .A2(n3508), .ZN(n3373) );
  NAND2_X1 U4191 ( .A1(n3374), .A2(n3373), .ZN(n3375) );
  XNOR2_X1 U4192 ( .A(n3375), .B(n2975), .ZN(n3377) );
  OAI22_X1 U4193 ( .A1(n2618), .A2(n3448), .B1(n3511), .B2(n3376), .ZN(n3378)
         );
  NAND2_X1 U4194 ( .A1(n3377), .A2(n3378), .ZN(n3599) );
  OAI21_X1 U4195 ( .B1(n3595), .B2(n3597), .A(n3599), .ZN(n3383) );
  NAND3_X1 U4196 ( .A1(n3599), .A2(n3597), .A3(n3595), .ZN(n3381) );
  INV_X1 U4197 ( .A(n3377), .ZN(n3380) );
  INV_X1 U4198 ( .A(n3378), .ZN(n3379) );
  NAND2_X1 U4199 ( .A1(n3380), .A2(n3379), .ZN(n3600) );
  AND2_X1 U4200 ( .A1(n3381), .A2(n3600), .ZN(n3382) );
  OAI22_X1 U4201 ( .A1(n4989), .A2(n3511), .B1(n3472), .B2(n3508), .ZN(n3384)
         );
  XNOR2_X1 U4202 ( .A(n3384), .B(n3509), .ZN(n3468) );
  OAI22_X1 U4203 ( .A1(n4299), .A2(n3511), .B1(n3508), .B2(n4317), .ZN(n3385)
         );
  XNOR2_X1 U4204 ( .A(n3385), .B(n3509), .ZN(n3387) );
  OAI22_X1 U4205 ( .A1(n4299), .A2(n3448), .B1(n3511), .B2(n4317), .ZN(n4321)
         );
  NAND2_X1 U4206 ( .A1(n4323), .A2(n4321), .ZN(n4306) );
  INV_X1 U4207 ( .A(n3386), .ZN(n3389) );
  INV_X1 U4208 ( .A(n3387), .ZN(n3388) );
  NAND2_X1 U4209 ( .A1(n4127), .A2(n3443), .ZN(n3391) );
  OR2_X1 U4210 ( .A1(n4303), .A2(n3508), .ZN(n3390) );
  NAND2_X1 U4211 ( .A1(n3391), .A2(n3390), .ZN(n3392) );
  XNOR2_X1 U4212 ( .A(n3392), .B(n3509), .ZN(n3393) );
  OAI22_X1 U4213 ( .A1(n4314), .A2(n3448), .B1(n3511), .B2(n4303), .ZN(n3394)
         );
  XNOR2_X1 U4214 ( .A(n3393), .B(n3394), .ZN(n4308) );
  NAND3_X1 U4215 ( .A1(n4306), .A2(n4322), .A3(n4308), .ZN(n3397) );
  NAND2_X1 U4216 ( .A1(n3397), .A2(n3396), .ZN(n3567) );
  OAI22_X1 U4217 ( .A1(n4300), .A2(n3447), .B1(n4133), .B2(n3508), .ZN(n3398)
         );
  XNOR2_X1 U4218 ( .A(n3398), .B(n2975), .ZN(n3569) );
  OAI22_X1 U4219 ( .A1(n4300), .A2(n3448), .B1(n4133), .B2(n3447), .ZN(n3399)
         );
  NOR2_X1 U4220 ( .A1(n3569), .A2(n3399), .ZN(n3401) );
  INV_X1 U4221 ( .A(n3569), .ZN(n3400) );
  INV_X1 U4222 ( .A(n3399), .ZN(n3568) );
  NAND2_X1 U4223 ( .A1(n4125), .A2(n3443), .ZN(n3403) );
  OR2_X1 U4224 ( .A1(n3405), .A2(n3508), .ZN(n3402) );
  NAND2_X1 U4225 ( .A1(n3403), .A2(n3402), .ZN(n3404) );
  XNOR2_X1 U4226 ( .A(n3404), .B(n3509), .ZN(n3408) );
  NOR2_X1 U4227 ( .A1(n3447), .A2(n3405), .ZN(n3406) );
  AOI21_X1 U4228 ( .B1(n3455), .B2(n4125), .A(n3406), .ZN(n3407) );
  NOR2_X1 U4229 ( .A1(n3408), .A2(n3407), .ZN(n3631) );
  NAND2_X1 U4230 ( .A1(n3408), .A2(n3407), .ZN(n3632) );
  OAI22_X1 U4231 ( .A1(n4078), .A2(n3448), .B1(n4097), .B2(n3511), .ZN(n3411)
         );
  OAI22_X1 U4232 ( .A1(n4078), .A2(n3511), .B1(n4097), .B2(n3508), .ZN(n3409)
         );
  XNOR2_X1 U4233 ( .A(n3409), .B(n2975), .ZN(n3410) );
  XOR2_X1 U4234 ( .A(n3411), .B(n3410), .Z(n3502) );
  NAND2_X1 U4235 ( .A1(n4092), .A2(n3443), .ZN(n3416) );
  OR2_X1 U4236 ( .A1(n3508), .A2(n4065), .ZN(n3415) );
  NAND2_X1 U4237 ( .A1(n3416), .A2(n3415), .ZN(n3417) );
  XNOR2_X1 U4238 ( .A(n3417), .B(n2975), .ZN(n3418) );
  INV_X1 U4239 ( .A(n4092), .ZN(n3542) );
  OAI22_X1 U4240 ( .A1(n3542), .A2(n3448), .B1(n3511), .B2(n4065), .ZN(n3419)
         );
  NAND2_X1 U4241 ( .A1(n3418), .A2(n3419), .ZN(n3587) );
  INV_X1 U4242 ( .A(n3418), .ZN(n3421) );
  INV_X1 U4243 ( .A(n3419), .ZN(n3420) );
  NAND2_X1 U4244 ( .A1(n3421), .A2(n3420), .ZN(n3586) );
  NAND2_X1 U4245 ( .A1(n4075), .A2(n3443), .ZN(n3423) );
  OR2_X1 U4246 ( .A1(n3508), .A2(n3544), .ZN(n3422) );
  NAND2_X1 U4247 ( .A1(n3423), .A2(n3422), .ZN(n3424) );
  XNOR2_X1 U4248 ( .A(n3424), .B(n3509), .ZN(n3426) );
  NOR2_X1 U4249 ( .A1(n3031), .A2(n3544), .ZN(n3425) );
  AOI21_X1 U4250 ( .B1(n3455), .B2(n4075), .A(n3425), .ZN(n3427) );
  AND2_X1 U4251 ( .A1(n3426), .A2(n3427), .ZN(n3535) );
  INV_X1 U4252 ( .A(n3426), .ZN(n3429) );
  INV_X1 U4253 ( .A(n3427), .ZN(n3428) );
  NAND2_X1 U4254 ( .A1(n3429), .A2(n3428), .ZN(n3536) );
  OAI22_X1 U4255 ( .A1(n4056), .A2(n3447), .B1(n4037), .B2(n3508), .ZN(n3430)
         );
  XNOR2_X1 U4256 ( .A(n3430), .B(n2975), .ZN(n3435) );
  OAI22_X1 U4257 ( .A1(n4056), .A2(n3448), .B1(n4037), .B2(n3447), .ZN(n3434)
         );
  XNOR2_X1 U4258 ( .A(n3435), .B(n3434), .ZN(n3611) );
  NOR2_X2 U4259 ( .A1(n3610), .A2(n3611), .ZN(n3479) );
  NAND2_X1 U4260 ( .A1(n4034), .A2(n3443), .ZN(n3432) );
  OR2_X1 U4261 ( .A1(n3508), .A2(n3484), .ZN(n3431) );
  NAND2_X1 U4262 ( .A1(n3432), .A2(n3431), .ZN(n3433) );
  XNOR2_X1 U4263 ( .A(n3433), .B(n2975), .ZN(n3438) );
  OAI22_X1 U4264 ( .A1(n3999), .A2(n3448), .B1(n3511), .B2(n3484), .ZN(n3437)
         );
  XNOR2_X1 U4265 ( .A(n3438), .B(n3437), .ZN(n3480) );
  NOR2_X1 U4266 ( .A1(n3435), .A2(n3434), .ZN(n3481) );
  AND2_X1 U4267 ( .A1(n3438), .A2(n3437), .ZN(n3442) );
  INV_X1 U4268 ( .A(n4021), .ZN(n3976) );
  OAI22_X1 U4269 ( .A1(n3976), .A2(n3448), .B1(n4001), .B2(n3511), .ZN(n3441)
         );
  INV_X1 U4270 ( .A(n3508), .ZN(n3439) );
  AOI22_X1 U4271 ( .A1(n3443), .A2(n4021), .B1(n3439), .B2(n3995), .ZN(n3440)
         );
  XNOR2_X1 U4272 ( .A(n3440), .B(n2975), .ZN(n3576) );
  NAND2_X1 U4273 ( .A1(n3996), .A2(n3443), .ZN(n3445) );
  OR2_X1 U4274 ( .A1(n3508), .A2(n3979), .ZN(n3444) );
  NAND2_X1 U4275 ( .A1(n3445), .A2(n3444), .ZN(n3446) );
  XNOR2_X1 U4276 ( .A(n3446), .B(n2975), .ZN(n3450) );
  OAI22_X1 U4277 ( .A1(n3956), .A2(n3448), .B1(n3979), .B2(n3447), .ZN(n3449)
         );
  AND2_X1 U4278 ( .A1(n3450), .A2(n3449), .ZN(n3559) );
  NAND2_X1 U4279 ( .A1(n3973), .A2(n3443), .ZN(n3452) );
  OR2_X1 U4280 ( .A1(n3508), .A2(n3959), .ZN(n3451) );
  NAND2_X1 U4281 ( .A1(n3452), .A2(n3451), .ZN(n3453) );
  XNOR2_X1 U4282 ( .A(n3453), .B(n3509), .ZN(n3459) );
  INV_X1 U4283 ( .A(n3459), .ZN(n3457) );
  NOR2_X1 U4284 ( .A1(n3511), .A2(n3959), .ZN(n3454) );
  AOI21_X1 U4285 ( .B1(n3455), .B2(n3973), .A(n3454), .ZN(n3458) );
  INV_X1 U4286 ( .A(n3458), .ZN(n3456) );
  NAND2_X1 U4287 ( .A1(n3457), .A2(n3456), .ZN(n3641) );
  OAI22_X1 U4288 ( .A1(n3952), .A2(n3033), .B1(n3511), .B2(n3941), .ZN(n3518)
         );
  OAI22_X1 U4289 ( .A1(n3952), .A2(n3447), .B1(n3508), .B2(n3941), .ZN(n3460)
         );
  XNOR2_X1 U4290 ( .A(n3460), .B(n2975), .ZN(n3519) );
  XOR2_X1 U4291 ( .A(n3518), .B(n3519), .Z(n3516) );
  XNOR2_X1 U4292 ( .A(n3517), .B(n3516), .ZN(n3466) );
  INV_X1 U4293 ( .A(n3942), .ZN(n3464) );
  INV_X1 U4294 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3461) );
  OAI22_X1 U4295 ( .A1(n4318), .A2(n3941), .B1(STATE_REG_SCAN_IN), .B2(n3461), 
        .ZN(n3463) );
  OAI22_X1 U4296 ( .A1(n3935), .A2(n4316), .B1(n4315), .B2(n3917), .ZN(n3462)
         );
  AOI211_X1 U4297 ( .C1(n3648), .C2(n3464), .A(n3463), .B(n3462), .ZN(n3465)
         );
  OAI21_X1 U4298 ( .B1(n3466), .B2(n4324), .A(n3465), .ZN(U3211) );
  XOR2_X1 U4299 ( .A(n3469), .B(n3468), .Z(n3470) );
  XNOR2_X1 U4300 ( .A(n3467), .B(n3470), .ZN(n3477) );
  INV_X1 U4301 ( .A(n3471), .ZN(n3475) );
  NAND2_X1 U4302 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4445) );
  OAI21_X1 U4303 ( .B1(n4318), .B2(n3472), .A(n4445), .ZN(n3474) );
  OAI22_X1 U4304 ( .A1(n2618), .A2(n4316), .B1(n4315), .B2(n4299), .ZN(n3473)
         );
  AOI211_X1 U4305 ( .C1(n3648), .C2(n3475), .A(n3474), .B(n3473), .ZN(n3476)
         );
  OAI21_X1 U4306 ( .B1(n3477), .B2(n4324), .A(n3476), .ZN(U3212) );
  INV_X1 U4307 ( .A(n3478), .ZN(n3483) );
  OAI21_X1 U4308 ( .B1(n3479), .B2(n3481), .A(n3480), .ZN(n3482) );
  NAND3_X1 U4309 ( .A1(n3483), .A2(n4309), .A3(n3482), .ZN(n3488) );
  NOR2_X1 U4310 ( .A1(n4318), .A2(n3484), .ZN(n3486) );
  OAI22_X1 U4311 ( .A1(n3976), .A2(n4315), .B1(n4316), .B2(n4056), .ZN(n3485)
         );
  AOI211_X1 U4312 ( .C1(REG3_REG_23__SCAN_IN), .C2(U3149), .A(n3486), .B(n3485), .ZN(n3487) );
  OAI211_X1 U4313 ( .C1(n4331), .C2(n4024), .A(n3488), .B(n3487), .ZN(U3213)
         );
  AND2_X1 U4314 ( .A1(n3357), .A2(n3489), .ZN(n3492) );
  OAI211_X1 U4315 ( .C1(n3492), .C2(n3491), .A(n4309), .B(n3490), .ZN(n3498)
         );
  OAI22_X1 U4316 ( .A1(n3493), .A2(n4316), .B1(n4315), .B2(n3552), .ZN(n3494)
         );
  AOI211_X1 U4317 ( .C1(n3496), .C2(n3638), .A(n3495), .B(n3494), .ZN(n3497)
         );
  OAI211_X1 U4318 ( .C1(n4331), .C2(n3499), .A(n3498), .B(n3497), .ZN(U3214)
         );
  OAI21_X1 U4319 ( .B1(n3502), .B2(n3501), .A(n3500), .ZN(n3503) );
  NAND2_X1 U4320 ( .A1(n3503), .A2(n4309), .ZN(n3507) );
  NOR2_X1 U4321 ( .A1(STATE_REG_SCAN_IN), .A2(n3504), .ZN(n3903) );
  OAI22_X1 U4322 ( .A1(n3542), .A2(n4315), .B1(n4316), .B2(n2659), .ZN(n3505)
         );
  AOI211_X1 U4323 ( .C1(n4091), .C2(n3638), .A(n3903), .B(n3505), .ZN(n3506)
         );
  OAI211_X1 U4324 ( .C1(n4331), .C2(n4099), .A(n3507), .B(n3506), .ZN(U3216)
         );
  INV_X1 U4325 ( .A(n3921), .ZN(n3512) );
  OAI22_X1 U4326 ( .A1(n3917), .A2(n3447), .B1(n3512), .B2(n3508), .ZN(n3510)
         );
  XNOR2_X1 U4327 ( .A(n3510), .B(n3509), .ZN(n3514) );
  OAI22_X1 U4328 ( .A1(n3917), .A2(n3448), .B1(n3512), .B2(n3511), .ZN(n3513)
         );
  XNOR2_X1 U4329 ( .A(n3514), .B(n3513), .ZN(n3525) );
  INV_X1 U4330 ( .A(n3525), .ZN(n3515) );
  NAND2_X1 U4331 ( .A1(n3515), .A2(n4309), .ZN(n3534) );
  NAND2_X1 U4332 ( .A1(n3517), .A2(n3516), .ZN(n3533) );
  NAND2_X1 U4333 ( .A1(n3519), .A2(n3518), .ZN(n3524) );
  INV_X1 U4334 ( .A(n3524), .ZN(n3520) );
  NOR2_X1 U4335 ( .A1(n3520), .A2(n4324), .ZN(n3521) );
  NAND2_X1 U4336 ( .A1(n3533), .A2(n3522), .ZN(n3532) );
  INV_X1 U4337 ( .A(n3523), .ZN(n3530) );
  NOR3_X1 U4338 ( .A1(n3525), .A2(n4324), .A3(n3524), .ZN(n3529) );
  AOI22_X1 U4339 ( .A1(n3638), .A2(n3921), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3527) );
  NAND2_X1 U4340 ( .A1(n3619), .A2(n3816), .ZN(n3526) );
  OAI211_X1 U4341 ( .C1(n3952), .C2(n4316), .A(n3527), .B(n3526), .ZN(n3528)
         );
  AOI211_X1 U4342 ( .C1(n3530), .C2(n3648), .A(n3529), .B(n3528), .ZN(n3531)
         );
  OAI211_X1 U4343 ( .C1(n3534), .C2(n3533), .A(n3532), .B(n3531), .ZN(U3217)
         );
  INV_X1 U4344 ( .A(n3535), .ZN(n3537) );
  NAND2_X1 U4345 ( .A1(n3537), .A2(n3536), .ZN(n3540) );
  INV_X1 U4346 ( .A(n3586), .ZN(n3585) );
  OAI211_X1 U4347 ( .C1(n3538), .C2(n3585), .A(n3587), .B(n3540), .ZN(n3539)
         );
  OAI211_X1 U4348 ( .C1(n3541), .C2(n3540), .A(n4309), .B(n3539), .ZN(n3548)
         );
  OAI22_X1 U4349 ( .A1(n3542), .A2(n4316), .B1(n4315), .B2(n4056), .ZN(n3546)
         );
  OAI22_X1 U4350 ( .A1(n4318), .A2(n3544), .B1(STATE_REG_SCAN_IN), .B2(n3543), 
        .ZN(n3545) );
  NOR2_X1 U4351 ( .A1(n3546), .A2(n3545), .ZN(n3547) );
  OAI211_X1 U4352 ( .C1(n4331), .C2(n4059), .A(n3548), .B(n3547), .ZN(U3220)
         );
  INV_X1 U4353 ( .A(n3595), .ZN(n3594) );
  XNOR2_X1 U4354 ( .A(n3594), .B(n3597), .ZN(n3550) );
  XNOR2_X1 U4355 ( .A(n3549), .B(n3550), .ZN(n3557) );
  NAND2_X1 U4356 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4420) );
  OAI21_X1 U4357 ( .B1(n4318), .B2(n3551), .A(n4420), .ZN(n3554) );
  OAI22_X1 U4358 ( .A1(n3552), .A2(n4316), .B1(n4315), .B2(n2618), .ZN(n3553)
         );
  AOI211_X1 U4359 ( .C1(n3648), .C2(n3555), .A(n3554), .B(n3553), .ZN(n3556)
         );
  OAI21_X1 U4360 ( .B1(n3557), .B2(n4324), .A(n3556), .ZN(U3221) );
  NOR2_X1 U4361 ( .A1(n2242), .A2(n3559), .ZN(n3560) );
  XNOR2_X1 U4362 ( .A(n3558), .B(n3560), .ZN(n3566) );
  INV_X1 U4363 ( .A(n3981), .ZN(n3564) );
  OAI22_X1 U4364 ( .A1(n4318), .A2(n3979), .B1(STATE_REG_SCAN_IN), .B2(n3561), 
        .ZN(n3563) );
  OAI22_X1 U4365 ( .A1(n3976), .A2(n4316), .B1(n4315), .B2(n3935), .ZN(n3562)
         );
  AOI211_X1 U4366 ( .C1(n3648), .C2(n3564), .A(n3563), .B(n3562), .ZN(n3565)
         );
  OAI21_X1 U4367 ( .B1(n3566), .B2(n4324), .A(n3565), .ZN(U3222) );
  XNOR2_X1 U4368 ( .A(n3569), .B(n3568), .ZN(n3570) );
  XNOR2_X1 U4369 ( .A(n3567), .B(n3570), .ZN(n3571) );
  NAND2_X1 U4370 ( .A1(n3571), .A2(n4309), .ZN(n3574) );
  AND2_X1 U4371 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4472) );
  OAI22_X1 U4372 ( .A1(n4314), .A2(n4316), .B1(n4315), .B2(n2659), .ZN(n3572)
         );
  AOI211_X1 U4373 ( .C1(n4124), .C2(n3638), .A(n4472), .B(n3572), .ZN(n3573)
         );
  OAI211_X1 U4374 ( .C1(n4331), .C2(n4136), .A(n3574), .B(n3573), .ZN(U3225)
         );
  NAND2_X1 U4375 ( .A1(n2232), .A2(n3575), .ZN(n3577) );
  XNOR2_X1 U4376 ( .A(n3577), .B(n3576), .ZN(n3583) );
  INV_X1 U4377 ( .A(n4002), .ZN(n3581) );
  INV_X1 U4378 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3578) );
  OAI22_X1 U4379 ( .A1(n4318), .A2(n4001), .B1(STATE_REG_SCAN_IN), .B2(n3578), 
        .ZN(n3580) );
  OAI22_X1 U4380 ( .A1(n3999), .A2(n4316), .B1(n4315), .B2(n3956), .ZN(n3579)
         );
  AOI211_X1 U4381 ( .C1(n3648), .C2(n3581), .A(n3580), .B(n3579), .ZN(n3582)
         );
  OAI21_X1 U4382 ( .B1(n3583), .B2(n4324), .A(n3582), .ZN(U3226) );
  NOR2_X1 U4383 ( .A1(n3584), .A2(n3585), .ZN(n3589) );
  AOI21_X1 U4384 ( .B1(n3587), .B2(n3586), .A(n3538), .ZN(n3588) );
  OAI21_X1 U4385 ( .B1(n3589), .B2(n3588), .A(n4309), .ZN(n3593) );
  NOR2_X1 U4386 ( .A1(n4318), .A2(n4065), .ZN(n3591) );
  OAI22_X1 U4387 ( .A1(n4078), .A2(n4316), .B1(n4315), .B2(n3613), .ZN(n3590)
         );
  AOI211_X1 U4388 ( .C1(REG3_REG_20__SCAN_IN), .C2(U3149), .A(n3591), .B(n3590), .ZN(n3592) );
  OAI211_X1 U4389 ( .C1(n4331), .C2(n4079), .A(n3593), .B(n3592), .ZN(U3230)
         );
  NOR2_X1 U4390 ( .A1(n3549), .A2(n3594), .ZN(n3598) );
  INV_X1 U4391 ( .A(n3549), .ZN(n3596) );
  OAI22_X1 U4392 ( .A1(n3598), .A2(n3597), .B1(n3596), .B2(n3595), .ZN(n3602)
         );
  NAND2_X1 U4393 ( .A1(n3600), .A2(n3599), .ZN(n3601) );
  XNOR2_X1 U4394 ( .A(n3602), .B(n3601), .ZN(n3603) );
  NAND2_X1 U4395 ( .A1(n3603), .A2(n4309), .ZN(n3608) );
  INV_X1 U4396 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4688) );
  NOR2_X1 U4397 ( .A1(STATE_REG_SCAN_IN), .A2(n4688), .ZN(n4431) );
  OAI22_X1 U4398 ( .A1(n3604), .A2(n4316), .B1(n4315), .B2(n4989), .ZN(n3605)
         );
  AOI211_X1 U4399 ( .C1(n3606), .C2(n3638), .A(n4431), .B(n3605), .ZN(n3607)
         );
  OAI211_X1 U4400 ( .C1(n4331), .C2(n3609), .A(n3608), .B(n3607), .ZN(U3231)
         );
  AOI21_X1 U4401 ( .B1(n3611), .B2(n3610), .A(n3479), .ZN(n3618) );
  INV_X1 U4402 ( .A(n4040), .ZN(n3616) );
  OAI22_X1 U4403 ( .A1(n4318), .A2(n4037), .B1(STATE_REG_SCAN_IN), .B2(n3612), 
        .ZN(n3615) );
  OAI22_X1 U4404 ( .A1(n3613), .A2(n4316), .B1(n4315), .B2(n3999), .ZN(n3614)
         );
  AOI211_X1 U4405 ( .C1(n3648), .C2(n3616), .A(n3615), .B(n3614), .ZN(n3617)
         );
  OAI21_X1 U4406 ( .B1(n3618), .B2(n4324), .A(n3617), .ZN(U3232) );
  AOI22_X1 U4407 ( .A1(n3620), .A2(n3819), .B1(n3619), .B2(n4494), .ZN(n3621)
         );
  NAND2_X1 U4408 ( .A1(REG3_REG_11__SCAN_IN), .A2(U3149), .ZN(n4409) );
  OAI211_X1 U4409 ( .C1(n4318), .C2(n4503), .A(n3621), .B(n4409), .ZN(n3629)
         );
  INV_X1 U4410 ( .A(n3622), .ZN(n3627) );
  AOI21_X1 U4411 ( .B1(n3626), .B2(n3624), .A(n3623), .ZN(n3625) );
  AOI211_X1 U4412 ( .C1(n3627), .C2(n3626), .A(n4324), .B(n3625), .ZN(n3628)
         );
  AOI211_X1 U4413 ( .C1(n4501), .C2(n3648), .A(n3629), .B(n3628), .ZN(n3630)
         );
  INV_X1 U4414 ( .A(n3630), .ZN(U3233) );
  INV_X1 U4415 ( .A(n3631), .ZN(n3633) );
  NAND2_X1 U4416 ( .A1(n3633), .A2(n3632), .ZN(n3634) );
  XNOR2_X1 U4417 ( .A(n3635), .B(n3634), .ZN(n3636) );
  NAND2_X1 U4418 ( .A1(n3636), .A2(n4309), .ZN(n3640) );
  AND2_X1 U4419 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n3886) );
  OAI22_X1 U4420 ( .A1(n4300), .A2(n4316), .B1(n4315), .B2(n4078), .ZN(n3637)
         );
  AOI211_X1 U4421 ( .C1(n4109), .C2(n3638), .A(n3886), .B(n3637), .ZN(n3639)
         );
  OAI211_X1 U4422 ( .C1(n4331), .C2(n4111), .A(n3640), .B(n3639), .ZN(U3235)
         );
  NAND2_X1 U4423 ( .A1(n2249), .A2(n3641), .ZN(n3642) );
  XNOR2_X1 U4424 ( .A(n3643), .B(n3642), .ZN(n3650) );
  INV_X1 U4425 ( .A(n3960), .ZN(n3647) );
  OAI22_X1 U4426 ( .A1(n4318), .A2(n3959), .B1(STATE_REG_SCAN_IN), .B2(n3644), 
        .ZN(n3646) );
  OAI22_X1 U4427 ( .A1(n3956), .A2(n4316), .B1(n4315), .B2(n3952), .ZN(n3645)
         );
  AOI211_X1 U4428 ( .C1(n3648), .C2(n3647), .A(n3646), .B(n3645), .ZN(n3649)
         );
  OAI21_X1 U4429 ( .B1(n3650), .B2(n4324), .A(n3649), .ZN(U3237) );
  NAND2_X1 U4430 ( .A1(n3713), .A2(DATAI_30_), .ZN(n4169) );
  NAND2_X1 U4431 ( .A1(n3915), .A2(n4169), .ZN(n3802) );
  NAND2_X1 U4432 ( .A1(n2492), .A2(REG1_REG_31__SCAN_IN), .ZN(n3654) );
  NAND2_X1 U4433 ( .A1(n2720), .A2(REG0_REG_31__SCAN_IN), .ZN(n3653) );
  NAND2_X1 U4434 ( .A1(n3651), .A2(REG2_REG_31__SCAN_IN), .ZN(n3652) );
  NAND3_X1 U4435 ( .A1(n3654), .A2(n3653), .A3(n3652), .ZN(n4160) );
  NAND2_X1 U4436 ( .A1(n3713), .A2(DATAI_31_), .ZN(n4159) );
  OR2_X1 U4437 ( .A1(n4160), .A2(n4159), .ZN(n3655) );
  NAND2_X1 U4438 ( .A1(n3802), .A2(n3655), .ZN(n3740) );
  INV_X1 U4439 ( .A(n3740), .ZN(n3727) );
  INV_X1 U4440 ( .A(n3656), .ZN(n3657) );
  NOR2_X1 U4441 ( .A1(n3657), .A2(n3744), .ZN(n3794) );
  INV_X1 U4442 ( .A(n3658), .ZN(n3661) );
  OAI211_X1 U4443 ( .C1(n3661), .C2(n2771), .A(n3660), .B(n3659), .ZN(n3663)
         );
  NAND3_X1 U4444 ( .A1(n3663), .A2(n3662), .A3(n2750), .ZN(n3666) );
  NAND3_X1 U4445 ( .A1(n3666), .A2(n3665), .A3(n3664), .ZN(n3669) );
  NAND3_X1 U4446 ( .A1(n3669), .A2(n3668), .A3(n3667), .ZN(n3671) );
  NAND4_X1 U4447 ( .A1(n3671), .A2(n3670), .A3(n2240), .A4(n3685), .ZN(n3675)
         );
  INV_X1 U4448 ( .A(n3757), .ZN(n3674) );
  INV_X1 U4449 ( .A(n3672), .ZN(n3673) );
  NAND3_X1 U4450 ( .A1(n3675), .A2(n3674), .A3(n3673), .ZN(n3681) );
  NOR2_X1 U4451 ( .A1(n3677), .A2(n3676), .ZN(n3687) );
  INV_X1 U4452 ( .A(n3678), .ZN(n3680) );
  AOI211_X1 U4453 ( .C1(n3681), .C2(n3687), .A(n3680), .B(n3679), .ZN(n3690)
         );
  NAND2_X1 U4454 ( .A1(n3683), .A2(n3682), .ZN(n3689) );
  INV_X1 U4455 ( .A(n3684), .ZN(n3686) );
  NAND2_X1 U4456 ( .A1(n3689), .A2(n3697), .ZN(n3778) );
  NAND4_X1 U4457 ( .A1(n3687), .A2(n3686), .A3(n3778), .A4(n3685), .ZN(n3688)
         );
  OAI21_X1 U4458 ( .B1(n3690), .B2(n3689), .A(n3688), .ZN(n3693) );
  AOI22_X1 U4459 ( .A1(n3693), .A2(n3692), .B1(n3691), .B2(n3778), .ZN(n3696)
         );
  OR4_X1 U4460 ( .A1(n3696), .A2(n3695), .A3(n3694), .A4(n3700), .ZN(n3705) );
  NAND2_X1 U4461 ( .A1(n3698), .A2(n3697), .ZN(n3779) );
  INV_X1 U4462 ( .A(n3779), .ZN(n3699) );
  OAI21_X1 U4463 ( .B1(n3701), .B2(n3700), .A(n3699), .ZN(n3703) );
  OAI21_X1 U4464 ( .B1(n3703), .B2(n3702), .A(n3778), .ZN(n3704) );
  AOI21_X1 U4465 ( .B1(n3705), .B2(n3704), .A(n3783), .ZN(n3707) );
  INV_X1 U4466 ( .A(n4011), .ZN(n3706) );
  NOR2_X1 U4467 ( .A1(n3706), .A2(n3733), .ZN(n3781) );
  OAI211_X1 U4468 ( .C1(n3776), .C2(n3707), .A(n3781), .B(n4013), .ZN(n3708)
         );
  OAI221_X1 U4469 ( .B1(n3710), .B2(n3709), .C1(n3710), .C2(n3708), .A(n3789), 
        .ZN(n3711) );
  OAI221_X1 U4470 ( .B1(n2289), .B2(n3712), .C1(n2289), .C2(n3711), .A(n3798), 
        .ZN(n3717) );
  NAND2_X1 U4471 ( .A1(n3713), .A2(DATAI_29_), .ZN(n3741) );
  NAND2_X1 U4472 ( .A1(n3816), .A2(n3741), .ZN(n3719) );
  NAND4_X1 U4473 ( .A1(n3719), .A2(n3911), .A3(n3715), .A4(n3714), .ZN(n3716)
         );
  AOI21_X1 U4474 ( .B1(n3794), .B2(n3717), .A(n3716), .ZN(n3724) );
  INV_X1 U4475 ( .A(n3792), .ZN(n3910) );
  INV_X1 U4476 ( .A(n3791), .ZN(n3718) );
  NOR2_X1 U4477 ( .A1(n3910), .A2(n3718), .ZN(n3723) );
  NAND2_X1 U4478 ( .A1(n3719), .A2(n3911), .ZN(n3772) );
  INV_X1 U4479 ( .A(n4169), .ZN(n3721) );
  INV_X1 U4480 ( .A(n3915), .ZN(n3720) );
  INV_X1 U4481 ( .A(n4160), .ZN(n3803) );
  INV_X1 U4482 ( .A(n4159), .ZN(n4163) );
  NOR2_X1 U4483 ( .A1(n3803), .A2(n4163), .ZN(n3725) );
  AOI21_X1 U4484 ( .B1(n3721), .B2(n3720), .A(n3725), .ZN(n3795) );
  INV_X1 U4485 ( .A(n3816), .ZN(n3722) );
  NAND2_X1 U4486 ( .A1(n3722), .A2(n3925), .ZN(n3793) );
  OAI211_X1 U4487 ( .C1(n3723), .C2(n3772), .A(n3795), .B(n3793), .ZN(n3775)
         );
  OR2_X1 U4488 ( .A1(n3724), .A2(n3775), .ZN(n3726) );
  AOI21_X1 U4489 ( .B1(n3727), .B2(n3726), .A(n3725), .ZN(n3771) );
  INV_X1 U4490 ( .A(n3729), .ZN(n3731) );
  NAND2_X1 U4491 ( .A1(n3731), .A2(n3730), .ZN(n4018) );
  XNOR2_X1 U4492 ( .A(n4092), .B(n4074), .ZN(n4072) );
  NAND4_X1 U4493 ( .A1(n4033), .A2(n4051), .A3(n4018), .A4(n4072), .ZN(n3750)
         );
  INV_X1 U4494 ( .A(n3732), .ZN(n4085) );
  NOR2_X1 U4495 ( .A1(n3733), .A2(n4085), .ZN(n4122) );
  INV_X1 U4496 ( .A(n3734), .ZN(n3736) );
  OR2_X1 U4497 ( .A1(n3736), .A2(n3735), .ZN(n4090) );
  NAND4_X1 U4498 ( .A1(n4115), .A2(n2391), .A3(n4122), .A4(n4090), .ZN(n3749)
         );
  INV_X1 U4499 ( .A(n3737), .ZN(n3739) );
  OR4_X1 U4500 ( .A1(n3949), .A2(n3939), .A3(n3919), .A4(n3740), .ZN(n3748) );
  XOR2_X1 U4501 ( .A(n3741), .B(n3816), .Z(n3922) );
  INV_X1 U4502 ( .A(n3742), .ZN(n3743) );
  NOR2_X1 U4503 ( .A1(n3744), .A2(n3743), .ZN(n3970) );
  INV_X1 U4504 ( .A(n3967), .ZN(n3746) );
  OR2_X1 U4505 ( .A1(n3746), .A2(n3745), .ZN(n3987) );
  INV_X1 U4506 ( .A(n3987), .ZN(n3992) );
  NAND4_X1 U4507 ( .A1(n3922), .A2(n3970), .A3(n3992), .A4(n3795), .ZN(n3747)
         );
  NOR4_X1 U4508 ( .A1(n3750), .A2(n3749), .A3(n3748), .A4(n3747), .ZN(n3769)
         );
  OR4_X1 U4509 ( .A1(n3753), .A2(n3752), .A3(n3751), .A4(n4489), .ZN(n3756) );
  NOR4_X1 U4510 ( .A1(n3756), .A2(n4546), .A3(n3755), .A4(n3754), .ZN(n3767)
         );
  NOR4_X1 U4511 ( .A1(n2752), .A2(n3759), .A3(n3758), .A4(n3757), .ZN(n3766)
         );
  NOR4_X1 U4512 ( .A1(n2312), .A2(n3763), .A3(n3762), .A4(n3761), .ZN(n3765)
         );
  AND4_X1 U4513 ( .A1(n3767), .A2(n3766), .A3(n3765), .A4(n3764), .ZN(n3768)
         );
  AOI21_X1 U4514 ( .B1(n3769), .B2(n3768), .A(n2771), .ZN(n3770) );
  MUX2_X1 U4515 ( .A(n3771), .B(n3770), .S(n4284), .Z(n3809) );
  NOR3_X1 U4516 ( .A1(n3939), .A2(n3773), .A3(n3772), .ZN(n3774) );
  NOR2_X1 U4517 ( .A1(n3775), .A2(n3774), .ZN(n3801) );
  INV_X1 U4518 ( .A(n3776), .ZN(n3785) );
  INV_X1 U4519 ( .A(n3777), .ZN(n3780) );
  OAI21_X1 U4520 ( .B1(n3780), .B2(n3779), .A(n3778), .ZN(n3784) );
  INV_X1 U4521 ( .A(n3781), .ZN(n3782) );
  AOI211_X1 U4522 ( .C1(n3785), .C2(n3784), .A(n3783), .B(n3782), .ZN(n3786)
         );
  OAI21_X1 U4523 ( .B1(n3786), .B2(n4012), .A(n4013), .ZN(n3788) );
  OAI221_X1 U4524 ( .B1(n3790), .B2(n3789), .C1(n3790), .C2(n3788), .A(n3787), 
        .ZN(n3799) );
  NAND4_X1 U4525 ( .A1(n3794), .A2(n3793), .A3(n3792), .A4(n3791), .ZN(n3797)
         );
  INV_X1 U4526 ( .A(n3795), .ZN(n3796) );
  AOI211_X1 U4527 ( .C1(n3799), .C2(n3798), .A(n3797), .B(n3796), .ZN(n3800)
         );
  OAI22_X1 U4528 ( .A1(n3801), .A2(n3800), .B1(n4160), .B2(n4169), .ZN(n3807)
         );
  INV_X1 U4529 ( .A(n3802), .ZN(n3804) );
  OAI21_X1 U4530 ( .B1(n3804), .B2(n3803), .A(n4163), .ZN(n3806) );
  AOI21_X1 U4531 ( .B1(n3807), .B2(n3806), .A(n3805), .ZN(n3808) );
  NOR2_X1 U4532 ( .A1(n3809), .A2(n3808), .ZN(n3810) );
  XNOR2_X1 U4533 ( .A(n3810), .B(n3897), .ZN(n3815) );
  NAND2_X1 U4534 ( .A1(n3811), .A2(n3837), .ZN(n3812) );
  OAI211_X1 U4535 ( .C1(n2942), .C2(n3814), .A(n3812), .B(B_REG_SCAN_IN), .ZN(
        n3813) );
  OAI21_X1 U4536 ( .B1(n3815), .B2(n3814), .A(n3813), .ZN(U3239) );
  MUX2_X1 U4537 ( .A(n4160), .B(DATAO_REG_31__SCAN_IN), .S(n3822), .Z(U3581)
         );
  MUX2_X1 U4538 ( .A(n3816), .B(DATAO_REG_29__SCAN_IN), .S(n3822), .Z(U3579)
         );
  MUX2_X1 U4539 ( .A(n3973), .B(DATAO_REG_26__SCAN_IN), .S(n3822), .Z(U3576)
         );
  MUX2_X1 U4540 ( .A(n3996), .B(DATAO_REG_25__SCAN_IN), .S(n3822), .Z(U3575)
         );
  MUX2_X1 U4541 ( .A(n4021), .B(DATAO_REG_24__SCAN_IN), .S(n3822), .Z(U3574)
         );
  MUX2_X1 U4542 ( .A(n4075), .B(DATAO_REG_21__SCAN_IN), .S(n3822), .Z(U3571)
         );
  MUX2_X1 U4543 ( .A(n4092), .B(DATAO_REG_20__SCAN_IN), .S(n3822), .Z(U3570)
         );
  MUX2_X1 U4544 ( .A(n4125), .B(DATAO_REG_18__SCAN_IN), .S(n3822), .Z(U3568)
         );
  MUX2_X1 U4545 ( .A(DATAO_REG_15__SCAN_IN), .B(n3817), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4546 ( .A(n3818), .B(DATAO_REG_13__SCAN_IN), .S(n3822), .Z(U3563)
         );
  MUX2_X1 U4547 ( .A(n4494), .B(DATAO_REG_12__SCAN_IN), .S(n3822), .Z(U3562)
         );
  MUX2_X1 U4548 ( .A(n3819), .B(DATAO_REG_10__SCAN_IN), .S(n3822), .Z(U3560)
         );
  MUX2_X1 U4549 ( .A(n3820), .B(DATAO_REG_9__SCAN_IN), .S(n3822), .Z(U3559) );
  MUX2_X1 U4550 ( .A(n3821), .B(DATAO_REG_8__SCAN_IN), .S(n3822), .Z(U3558) );
  MUX2_X1 U4551 ( .A(n3823), .B(DATAO_REG_7__SCAN_IN), .S(n3822), .Z(U3557) );
  MUX2_X1 U4552 ( .A(DATAO_REG_3__SCAN_IN), .B(n3824), .S(U4043), .Z(U3553) );
  MUX2_X1 U4553 ( .A(DATAO_REG_0__SCAN_IN), .B(n3825), .S(U4043), .Z(U3550) );
  OAI211_X1 U4554 ( .C1(n3827), .C2(n3826), .A(n4481), .B(n3847), .ZN(n3832)
         );
  OAI211_X1 U4555 ( .C1(n3838), .C2(n3828), .A(n4483), .B(n3843), .ZN(n3831)
         );
  AOI22_X1 U4556 ( .A1(n4473), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3830) );
  NAND2_X1 U4557 ( .A1(n4458), .A2(n4286), .ZN(n3829) );
  NAND4_X1 U4558 ( .A1(n3832), .A2(n3831), .A3(n3830), .A4(n3829), .ZN(U3241)
         );
  NAND3_X1 U4559 ( .A1(n3834), .A2(n4287), .A3(n3833), .ZN(n3840) );
  NAND2_X1 U4560 ( .A1(n4339), .A2(n3835), .ZN(n3836) );
  NAND2_X1 U4561 ( .A1(n4287), .A2(n3836), .ZN(n4340) );
  AOI22_X1 U4562 ( .A1(n3838), .A2(n3837), .B1(n4340), .B2(n2498), .ZN(n3839)
         );
  NAND3_X1 U4563 ( .A1(n3840), .A2(U4043), .A3(n3839), .ZN(n4355) );
  AOI22_X1 U4564 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4473), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3855) );
  MUX2_X1 U4565 ( .A(n2896), .B(REG2_REG_2__SCAN_IN), .S(n4285), .Z(n3841) );
  NAND3_X1 U4566 ( .A1(n3843), .A2(n3842), .A3(n3841), .ZN(n3845) );
  AND3_X1 U4567 ( .A1(n4483), .A2(n3845), .A3(n3844), .ZN(n3846) );
  AOI21_X1 U4568 ( .B1(n4458), .B2(n4285), .A(n3846), .ZN(n3854) );
  INV_X1 U4569 ( .A(n3847), .ZN(n3852) );
  MUX2_X1 U4570 ( .A(n4852), .B(REG1_REG_2__SCAN_IN), .S(n4285), .Z(n3849) );
  NAND2_X1 U4571 ( .A1(n3849), .A2(n3848), .ZN(n3851) );
  OAI211_X1 U4572 ( .C1(n3852), .C2(n3851), .A(n4481), .B(n3850), .ZN(n3853)
         );
  NAND4_X1 U4573 ( .A1(n4355), .A2(n3855), .A3(n3854), .A4(n3853), .ZN(U3242)
         );
  XNOR2_X1 U4574 ( .A(n3901), .B(REG2_REG_18__SCAN_IN), .ZN(n3870) );
  NOR2_X1 U4575 ( .A1(n3883), .A2(REG2_REG_17__SCAN_IN), .ZN(n3856) );
  AOI21_X1 U4576 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3883), .A(n3856), .ZN(n4476) );
  INV_X1 U4577 ( .A(n4444), .ZN(n4529) );
  NOR2_X1 U4578 ( .A1(n3303), .A2(n4530), .ZN(n4432) );
  INV_X1 U4579 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4580 ( .A1(n3875), .A2(REG2_REG_11__SCAN_IN), .B1(n3861), .B2(
        n4534), .ZN(n4414) );
  NAND2_X1 U4581 ( .A1(n3858), .A2(n3857), .ZN(n3860) );
  NAND2_X1 U4582 ( .A1(n4531), .A2(n3862), .ZN(n3863) );
  NAND2_X1 U4583 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4424), .ZN(n4423) );
  NAND2_X1 U4584 ( .A1(n3863), .A2(n4423), .ZN(n4434) );
  NOR2_X1 U4585 ( .A1(n4529), .A2(n3864), .ZN(n3865) );
  NAND2_X1 U4586 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4457), .ZN(n3866) );
  OAI21_X1 U4587 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4457), .A(n3866), .ZN(n4453) );
  NOR2_X1 U4588 ( .A1(n4454), .A2(n4453), .ZN(n4452) );
  NAND2_X1 U4589 ( .A1(n3867), .A2(n4527), .ZN(n3868) );
  INV_X1 U4590 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4464) );
  NAND2_X1 U4591 ( .A1(n4476), .A2(n4475), .ZN(n4474) );
  OAI21_X1 U4592 ( .B1(n3883), .B2(REG2_REG_17__SCAN_IN), .A(n4474), .ZN(n3869) );
  AOI21_X1 U4593 ( .B1(n3870), .B2(n3869), .A(n3900), .ZN(n3871) );
  NAND2_X1 U4594 ( .A1(n4483), .A2(n3871), .ZN(n3892) );
  INV_X1 U4595 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4216) );
  INV_X1 U4596 ( .A(n3883), .ZN(n4525) );
  AOI22_X1 U4597 ( .A1(n3883), .A2(REG1_REG_17__SCAN_IN), .B1(n4216), .B2(
        n4525), .ZN(n4479) );
  INV_X1 U4598 ( .A(n3872), .ZN(n3874) );
  INV_X1 U4599 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4608) );
  AOI22_X1 U4600 ( .A1(n3875), .A2(n4608), .B1(REG1_REG_11__SCAN_IN), .B2(
        n4534), .ZN(n4408) );
  NOR2_X1 U4601 ( .A1(n3876), .A2(n4427), .ZN(n3877) );
  INV_X1 U4602 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4235) );
  AOI22_X1 U4603 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4530), .B1(n3878), .B2(
        n4235), .ZN(n4429) );
  NOR2_X1 U4604 ( .A1(n3879), .A2(n4529), .ZN(n3880) );
  INV_X1 U4605 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4873) );
  XOR2_X1 U4606 ( .A(n4444), .B(n3879), .Z(n4439) );
  NOR2_X1 U4607 ( .A1(n4873), .A2(n4439), .ZN(n4438) );
  NOR2_X1 U4608 ( .A1(n3880), .A2(n4438), .ZN(n4450) );
  INV_X1 U4609 ( .A(n4457), .ZN(n4528) );
  INV_X1 U4610 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4224) );
  AOI22_X1 U4611 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4528), .B1(n4457), .B2(
        n4224), .ZN(n4449) );
  NOR2_X1 U4612 ( .A1(n4450), .A2(n4449), .ZN(n4448) );
  NAND2_X1 U4613 ( .A1(n3881), .A2(n4527), .ZN(n3882) );
  INV_X1 U4614 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4855) );
  NAND2_X1 U4615 ( .A1(n4479), .A2(n4478), .ZN(n4477) );
  OAI21_X1 U4616 ( .B1(n3883), .B2(REG1_REG_17__SCAN_IN), .A(n4477), .ZN(n3885) );
  INV_X1 U4617 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4729) );
  OR2_X1 U4618 ( .A1(n3893), .A2(n4729), .ZN(n3894) );
  OAI21_X1 U4619 ( .B1(n3901), .B2(REG1_REG_18__SCAN_IN), .A(n3894), .ZN(n3884) );
  NOR2_X1 U4620 ( .A1(n3885), .A2(n3884), .ZN(n3896) );
  INV_X1 U4621 ( .A(n3896), .ZN(n3889) );
  AOI21_X1 U4622 ( .B1(n4473), .B2(ADDR_REG_18__SCAN_IN), .A(n3886), .ZN(n3887) );
  OAI211_X1 U4623 ( .C1(n3893), .C2(n4486), .A(n3892), .B(n3891), .ZN(U3258)
         );
  INV_X1 U4624 ( .A(n3894), .ZN(n3895) );
  NOR2_X1 U4625 ( .A1(n3896), .A2(n3895), .ZN(n3899) );
  XNOR2_X1 U4626 ( .A(n3897), .B(REG1_REG_19__SCAN_IN), .ZN(n3898) );
  XNOR2_X1 U4627 ( .A(n3899), .B(n3898), .ZN(n3908) );
  INV_X1 U4628 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4897) );
  MUX2_X1 U4629 ( .A(n4897), .B(REG2_REG_19__SCAN_IN), .S(n3905), .Z(n3902) );
  AOI21_X1 U4630 ( .B1(n4473), .B2(ADDR_REG_19__SCAN_IN), .A(n3903), .ZN(n3904) );
  OAI21_X1 U4631 ( .B1(n4486), .B2(n3905), .A(n3904), .ZN(n3906) );
  OAI21_X1 U4632 ( .B1(n3908), .B2(n4447), .A(n3907), .ZN(U3259) );
  INV_X1 U4633 ( .A(n3909), .ZN(n3918) );
  AOI21_X1 U4634 ( .B1(n3912), .B2(n3911), .A(n3910), .ZN(n3913) );
  XOR2_X1 U4635 ( .A(n3922), .B(n3913), .Z(n3914) );
  AOI21_X1 U4636 ( .B1(B_REG_SCAN_IN), .B2(n4339), .A(n4055), .ZN(n4161) );
  AOI22_X1 U4637 ( .A1(n4161), .A2(n3915), .B1(n3925), .B2(n4162), .ZN(n3916)
         );
  AOI21_X1 U4638 ( .B1(n3918), .B2(n4508), .A(n4174), .ZN(n3928) );
  XNOR2_X1 U4639 ( .A(n3923), .B(n3922), .ZN(n4173) );
  NAND2_X1 U4640 ( .A1(n4173), .A2(n4068), .ZN(n3927) );
  AOI22_X1 U4641 ( .A1(n4175), .A2(n4513), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4519), .ZN(n3926) );
  OAI211_X1 U4642 ( .C1(n4519), .C2(n3928), .A(n3927), .B(n3926), .ZN(U3354)
         );
  OAI21_X1 U4643 ( .B1(n3931), .B2(n3930), .A(n3929), .ZN(n3937) );
  AOI22_X1 U4644 ( .A1(n3933), .A2(n4495), .B1(n4162), .B2(n3932), .ZN(n3934)
         );
  OAI21_X1 U4645 ( .B1(n3935), .B2(n4491), .A(n3934), .ZN(n3936) );
  AOI21_X1 U4646 ( .B1(n3937), .B2(n4145), .A(n3936), .ZN(n4177) );
  XNOR2_X1 U4647 ( .A(n3938), .B(n3939), .ZN(n4176) );
  NAND2_X1 U4648 ( .A1(n4176), .A2(n4068), .ZN(n3947) );
  OAI21_X1 U4649 ( .B1(n3957), .B2(n3941), .A(n3940), .ZN(n4179) );
  INV_X1 U4650 ( .A(n4179), .ZN(n3945) );
  INV_X1 U4651 ( .A(REG2_REG_27__SCAN_IN), .ZN(n3943) );
  OAI22_X1 U4652 ( .A1(n4337), .A2(n3943), .B1(n3942), .B2(n4151), .ZN(n3944)
         );
  AOI21_X1 U4653 ( .B1(n3945), .B2(n4513), .A(n3944), .ZN(n3946) );
  OAI211_X1 U4654 ( .C1(n4177), .C2(n4519), .A(n3947), .B(n3946), .ZN(U3263)
         );
  XOR2_X1 U4655 ( .A(n3949), .B(n3948), .Z(n4181) );
  INV_X1 U4656 ( .A(n4181), .ZN(n3965) );
  XNOR2_X1 U4657 ( .A(n3950), .B(n3949), .ZN(n3951) );
  NAND2_X1 U4658 ( .A1(n3951), .A2(n4145), .ZN(n3955) );
  OAI22_X1 U4659 ( .A1(n3952), .A2(n4055), .B1(n4490), .B2(n3959), .ZN(n3953)
         );
  INV_X1 U4660 ( .A(n3953), .ZN(n3954) );
  OAI211_X1 U4661 ( .C1(n3956), .C2(n4491), .A(n3955), .B(n3954), .ZN(n4180)
         );
  INV_X1 U4662 ( .A(n3957), .ZN(n3958) );
  OAI21_X1 U4663 ( .B1(n3977), .B2(n3959), .A(n3958), .ZN(n4248) );
  NOR2_X1 U4664 ( .A1(n4248), .A2(n4135), .ZN(n3963) );
  INV_X1 U4665 ( .A(REG2_REG_26__SCAN_IN), .ZN(n3961) );
  OAI22_X1 U4666 ( .A1(n4337), .A2(n3961), .B1(n3960), .B2(n4151), .ZN(n3962)
         );
  AOI211_X1 U4667 ( .C1(n4180), .C2(n4337), .A(n3963), .B(n3962), .ZN(n3964)
         );
  OAI21_X1 U4668 ( .B1(n3965), .B2(n4155), .A(n3964), .ZN(U3264) );
  XNOR2_X1 U4669 ( .A(n3966), .B(n3970), .ZN(n4185) );
  INV_X1 U4670 ( .A(n4185), .ZN(n3986) );
  NAND2_X1 U4671 ( .A1(n3968), .A2(n3967), .ZN(n3969) );
  XOR2_X1 U4672 ( .A(n3970), .B(n3969), .Z(n3971) );
  NAND2_X1 U4673 ( .A1(n3971), .A2(n4145), .ZN(n3975) );
  AOI22_X1 U4674 ( .A1(n3973), .A2(n4495), .B1(n4162), .B2(n3972), .ZN(n3974)
         );
  OAI211_X1 U4675 ( .C1(n3976), .C2(n4491), .A(n3975), .B(n3974), .ZN(n4184)
         );
  INV_X1 U4676 ( .A(n4000), .ZN(n3980) );
  INV_X1 U4677 ( .A(n3977), .ZN(n3978) );
  OAI21_X1 U4678 ( .B1(n3980), .B2(n3979), .A(n3978), .ZN(n4251) );
  NOR2_X1 U4679 ( .A1(n4251), .A2(n4135), .ZN(n3984) );
  INV_X1 U4680 ( .A(REG2_REG_25__SCAN_IN), .ZN(n3982) );
  OAI22_X1 U4681 ( .A1(n4337), .A2(n3982), .B1(n3981), .B2(n4151), .ZN(n3983)
         );
  AOI211_X1 U4682 ( .C1(n4184), .C2(n4337), .A(n3984), .B(n3983), .ZN(n3985)
         );
  OAI21_X1 U4683 ( .B1(n3986), .B2(n4155), .A(n3985), .ZN(U3265) );
  XNOR2_X1 U4684 ( .A(n3988), .B(n3987), .ZN(n4188) );
  INV_X1 U4685 ( .A(n4188), .ZN(n4007) );
  INV_X1 U4686 ( .A(n3989), .ZN(n3990) );
  NAND2_X1 U4687 ( .A1(n3991), .A2(n3990), .ZN(n3993) );
  XNOR2_X1 U4688 ( .A(n3993), .B(n3992), .ZN(n3994) );
  NAND2_X1 U4689 ( .A1(n3994), .A2(n4145), .ZN(n3998) );
  AOI22_X1 U4690 ( .A1(n3996), .A2(n4495), .B1(n4162), .B2(n3995), .ZN(n3997)
         );
  OAI211_X1 U4691 ( .C1(n3999), .C2(n4491), .A(n3998), .B(n3997), .ZN(n4187)
         );
  OAI21_X1 U4692 ( .B1(n2272), .B2(n4001), .A(n4000), .ZN(n4255) );
  NOR2_X1 U4693 ( .A1(n4255), .A2(n4135), .ZN(n4005) );
  INV_X1 U4694 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4003) );
  OAI22_X1 U4695 ( .A1(n4337), .A2(n4003), .B1(n4002), .B2(n4151), .ZN(n4004)
         );
  AOI211_X1 U4696 ( .C1(n4187), .C2(n4337), .A(n4005), .B(n4004), .ZN(n4006)
         );
  OAI21_X1 U4697 ( .B1(n4007), .B2(n4155), .A(n4006), .ZN(U3266) );
  NAND2_X1 U4698 ( .A1(n4194), .A2(n4020), .ZN(n4008) );
  NAND2_X1 U4699 ( .A1(n4009), .A2(n4008), .ZN(n4258) );
  XNOR2_X1 U4700 ( .A(n4010), .B(n4018), .ZN(n4191) );
  NAND2_X1 U4701 ( .A1(n4191), .A2(n4068), .ZN(n4028) );
  AND2_X1 U4702 ( .A1(n4011), .A2(n4086), .ZN(n4069) );
  OR2_X1 U4703 ( .A1(n4012), .A2(n4069), .ZN(n4014) );
  AND2_X1 U4704 ( .A1(n4014), .A2(n4013), .ZN(n4050) );
  NAND2_X1 U4705 ( .A1(n4050), .A2(n4051), .ZN(n4049) );
  NAND2_X1 U4706 ( .A1(n4015), .A2(n4049), .ZN(n4032) );
  NAND2_X1 U4707 ( .A1(n4033), .A2(n4032), .ZN(n4031) );
  NAND2_X1 U4708 ( .A1(n4016), .A2(n4031), .ZN(n4017) );
  XNOR2_X1 U4709 ( .A(n4018), .B(n4017), .ZN(n4019) );
  NAND2_X1 U4710 ( .A1(n4019), .A2(n4145), .ZN(n4023) );
  AOI22_X1 U4711 ( .A1(n4021), .A2(n4495), .B1(n4020), .B2(n4162), .ZN(n4022)
         );
  OAI211_X1 U4712 ( .C1(n4056), .C2(n4491), .A(n4023), .B(n4022), .ZN(n4190)
         );
  INV_X1 U4713 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4025) );
  OAI22_X1 U4714 ( .A1(n4337), .A2(n4025), .B1(n4024), .B2(n4151), .ZN(n4026)
         );
  AOI21_X1 U4715 ( .B1(n4337), .B2(n4190), .A(n4026), .ZN(n4027) );
  OAI211_X1 U4716 ( .C1(n4258), .C2(n4135), .A(n4028), .B(n4027), .ZN(U3267)
         );
  OAI21_X1 U4717 ( .B1(n4029), .B2(n2692), .A(n4030), .ZN(n4198) );
  OAI21_X1 U4718 ( .B1(n4033), .B2(n4032), .A(n4031), .ZN(n4039) );
  NAND2_X1 U4719 ( .A1(n4075), .A2(n4126), .ZN(n4036) );
  NAND2_X1 U4720 ( .A1(n4034), .A2(n4495), .ZN(n4035) );
  OAI211_X1 U4721 ( .C1(n4490), .C2(n4037), .A(n4036), .B(n4035), .ZN(n4038)
         );
  AOI21_X1 U4722 ( .B1(n4039), .B2(n4145), .A(n4038), .ZN(n4197) );
  OAI22_X1 U4723 ( .A1(n4197), .A2(n4519), .B1(n4040), .B2(n4151), .ZN(n4044)
         );
  INV_X1 U4724 ( .A(n4048), .ZN(n4042) );
  NAND2_X1 U4725 ( .A1(n4042), .A2(n4041), .ZN(n4195) );
  AND3_X1 U4726 ( .A1(n4195), .A2(n4513), .A3(n4194), .ZN(n4043) );
  AOI211_X1 U4727 ( .C1(n4519), .C2(REG2_REG_22__SCAN_IN), .A(n4044), .B(n4043), .ZN(n4045) );
  OAI21_X1 U4728 ( .B1(n4198), .B2(n4155), .A(n4045), .ZN(U3268) );
  XOR2_X1 U4729 ( .A(n4051), .B(n4046), .Z(n4202) );
  AND2_X1 U4730 ( .A1(n4064), .A2(n4052), .ZN(n4047) );
  NOR2_X1 U4731 ( .A1(n4048), .A2(n4047), .ZN(n4199) );
  OAI21_X1 U4732 ( .B1(n4051), .B2(n4050), .A(n4049), .ZN(n4058) );
  NAND2_X1 U4733 ( .A1(n4162), .A2(n4052), .ZN(n4054) );
  NAND2_X1 U4734 ( .A1(n4092), .A2(n4126), .ZN(n4053) );
  OAI211_X1 U4735 ( .C1(n4056), .C2(n4055), .A(n4054), .B(n4053), .ZN(n4057)
         );
  AOI21_X1 U4736 ( .B1(n4058), .B2(n4145), .A(n4057), .ZN(n4201) );
  NOR2_X1 U4737 ( .A1(n4201), .A2(n4519), .ZN(n4062) );
  INV_X1 U4738 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4060) );
  OAI22_X1 U4739 ( .A1(n4337), .A2(n4060), .B1(n4059), .B2(n4151), .ZN(n4061)
         );
  AOI211_X1 U4740 ( .C1(n4199), .C2(n4513), .A(n4062), .B(n4061), .ZN(n4063)
         );
  OAI21_X1 U4741 ( .B1(n4202), .B2(n4155), .A(n4063), .ZN(U3269) );
  INV_X1 U4742 ( .A(n4096), .ZN(n4066) );
  OAI21_X1 U4743 ( .B1(n4066), .B2(n4065), .A(n4064), .ZN(n4263) );
  XNOR2_X1 U4744 ( .A(n4067), .B(n4072), .ZN(n4204) );
  NAND2_X1 U4745 ( .A1(n4204), .A2(n4068), .ZN(n4083) );
  NOR2_X1 U4746 ( .A1(n4070), .A2(n4069), .ZN(n4071) );
  XOR2_X1 U4747 ( .A(n4072), .B(n4071), .Z(n4073) );
  NAND2_X1 U4748 ( .A1(n4073), .A2(n4145), .ZN(n4077) );
  AOI22_X1 U4749 ( .A1(n4075), .A2(n4495), .B1(n4162), .B2(n4074), .ZN(n4076)
         );
  OAI211_X1 U4750 ( .C1(n4078), .C2(n4491), .A(n4077), .B(n4076), .ZN(n4203)
         );
  INV_X1 U4751 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4080) );
  OAI22_X1 U4752 ( .A1(n4337), .A2(n4080), .B1(n4079), .B2(n4151), .ZN(n4081)
         );
  AOI21_X1 U4753 ( .B1(n4203), .B2(n4337), .A(n4081), .ZN(n4082) );
  OAI211_X1 U4754 ( .C1(n4263), .C2(n4135), .A(n4083), .B(n4082), .ZN(U3270)
         );
  XOR2_X1 U4755 ( .A(n4090), .B(n4084), .Z(n4208) );
  INV_X1 U4756 ( .A(n4208), .ZN(n4103) );
  NOR2_X1 U4757 ( .A1(n4086), .A2(n4085), .ZN(n4104) );
  AOI21_X1 U4758 ( .B1(n4104), .B2(n4088), .A(n4087), .ZN(n4089) );
  XOR2_X1 U4759 ( .A(n4090), .B(n4089), .Z(n4095) );
  AOI22_X1 U4760 ( .A1(n4092), .A2(n4495), .B1(n4091), .B2(n4162), .ZN(n4094)
         );
  NAND2_X1 U4761 ( .A1(n4125), .A2(n4126), .ZN(n4093) );
  OAI211_X1 U4762 ( .C1(n4095), .C2(n4497), .A(n4094), .B(n4093), .ZN(n4207)
         );
  OAI21_X1 U4763 ( .B1(n4098), .B2(n4097), .A(n4096), .ZN(n4266) );
  NOR2_X1 U4764 ( .A1(n4266), .A2(n4135), .ZN(n4101) );
  OAI22_X1 U4765 ( .A1(n4337), .A2(n4897), .B1(n4099), .B2(n4151), .ZN(n4100)
         );
  AOI211_X1 U4766 ( .C1(n4207), .C2(n4337), .A(n4101), .B(n4100), .ZN(n4102)
         );
  OAI21_X1 U4767 ( .B1(n4155), .B2(n4103), .A(n4102), .ZN(U3271) );
  XOR2_X1 U4768 ( .A(n4115), .B(n4104), .Z(n4108) );
  AOI22_X1 U4769 ( .A1(n4105), .A2(n4495), .B1(n4162), .B2(n4109), .ZN(n4106)
         );
  OAI21_X1 U4770 ( .B1(n4300), .B2(n4491), .A(n4106), .ZN(n4107) );
  AOI21_X1 U4771 ( .B1(n4108), .B2(n4145), .A(n4107), .ZN(n4212) );
  XNOR2_X1 U4772 ( .A(n4131), .B(n4109), .ZN(n4110) );
  NAND2_X1 U4773 ( .A1(n4110), .A2(n4585), .ZN(n4211) );
  INV_X1 U4774 ( .A(n4211), .ZN(n4119) );
  OAI22_X1 U4775 ( .A1(n4337), .A2(n2328), .B1(n4111), .B2(n4151), .ZN(n4117)
         );
  INV_X1 U4776 ( .A(n4112), .ZN(n4113) );
  AOI21_X1 U4777 ( .B1(n4115), .B2(n4114), .A(n4113), .ZN(n4213) );
  NOR2_X1 U4778 ( .A1(n4213), .A2(n4155), .ZN(n4116) );
  AOI211_X1 U4779 ( .C1(n4119), .C2(n4118), .A(n4117), .B(n4116), .ZN(n4120)
         );
  OAI21_X1 U4780 ( .B1(n4519), .B2(n4212), .A(n4120), .ZN(U3272) );
  XNOR2_X1 U4781 ( .A(n4121), .B(n4122), .ZN(n4215) );
  INV_X1 U4782 ( .A(n4215), .ZN(n4140) );
  XNOR2_X1 U4783 ( .A(n4123), .B(n4122), .ZN(n4130) );
  AOI22_X1 U4784 ( .A1(n4125), .A2(n4495), .B1(n4162), .B2(n4124), .ZN(n4129)
         );
  NAND2_X1 U4785 ( .A1(n4127), .A2(n4126), .ZN(n4128) );
  OAI211_X1 U4786 ( .C1(n4130), .C2(n4497), .A(n4129), .B(n4128), .ZN(n4214)
         );
  INV_X1 U4787 ( .A(n4150), .ZN(n4134) );
  INV_X1 U4788 ( .A(n4131), .ZN(n4132) );
  OAI21_X1 U4789 ( .B1(n4134), .B2(n4133), .A(n4132), .ZN(n4271) );
  NOR2_X1 U4790 ( .A1(n4271), .A2(n4135), .ZN(n4138) );
  OAI22_X1 U4791 ( .A1(n4337), .A2(n4824), .B1(n4136), .B2(n4151), .ZN(n4137)
         );
  AOI211_X1 U4792 ( .C1(n4214), .C2(n4337), .A(n4138), .B(n4137), .ZN(n4139)
         );
  OAI21_X1 U4793 ( .B1(n4155), .B2(n4140), .A(n4139), .ZN(U3273) );
  XNOR2_X1 U4794 ( .A(n4141), .B(n2391), .ZN(n4146) );
  AOI22_X1 U4795 ( .A1(n4142), .A2(n4495), .B1(n4147), .B2(n4162), .ZN(n4143)
         );
  OAI21_X1 U4796 ( .B1(n4299), .B2(n4491), .A(n4143), .ZN(n4144) );
  AOI21_X1 U4797 ( .B1(n4146), .B2(n4145), .A(n4144), .ZN(n4220) );
  NAND2_X1 U4798 ( .A1(n4148), .A2(n4147), .ZN(n4149) );
  AND2_X1 U4799 ( .A1(n4150), .A2(n4149), .ZN(n4218) );
  OAI22_X1 U4800 ( .A1(n4337), .A2(n4464), .B1(n4313), .B2(n4151), .ZN(n4157)
         );
  OAI21_X1 U4801 ( .B1(n4154), .B2(n4153), .A(n4152), .ZN(n4221) );
  NOR2_X1 U4802 ( .A1(n4221), .A2(n4155), .ZN(n4156) );
  AOI211_X1 U4803 ( .C1(n4218), .C2(n4513), .A(n4157), .B(n4156), .ZN(n4158)
         );
  OAI21_X1 U4804 ( .B1(n4519), .B2(n4220), .A(n4158), .ZN(U3274) );
  NAND2_X1 U4805 ( .A1(n4166), .A2(n4169), .ZN(n4165) );
  XNOR2_X1 U4806 ( .A(n4165), .B(n4159), .ZN(n4332) );
  INV_X1 U4807 ( .A(n4332), .ZN(n4239) );
  INV_X1 U4808 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4742) );
  AND2_X1 U4809 ( .A1(n4161), .A2(n4160), .ZN(n4167) );
  AOI21_X1 U4810 ( .B1(n4163), .B2(n4162), .A(n4167), .ZN(n4334) );
  MUX2_X1 U4811 ( .A(n4742), .B(n4334), .S(n4610), .Z(n4164) );
  OAI21_X1 U4812 ( .B1(n4239), .B2(n4237), .A(n4164), .ZN(U3549) );
  INV_X1 U4813 ( .A(n4167), .ZN(n4168) );
  OAI21_X1 U4814 ( .B1(n4169), .B2(n4490), .A(n4168), .ZN(n4336) );
  INV_X1 U4815 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4170) );
  NOR2_X1 U4816 ( .A1(n4610), .A2(n4170), .ZN(n4171) );
  AOI21_X1 U4817 ( .B1(n4610), .B2(n4336), .A(n4171), .ZN(n4172) );
  OAI21_X1 U4818 ( .B1(n4335), .B2(n4237), .A(n4172), .ZN(U3548) );
  MUX2_X1 U4819 ( .A(REG1_REG_29__SCAN_IN), .B(n4243), .S(n4610), .Z(U3547) );
  NAND2_X1 U4820 ( .A1(n4176), .A2(n4577), .ZN(n4178) );
  OAI211_X1 U4821 ( .C1(n4587), .C2(n4179), .A(n4178), .B(n4177), .ZN(n4244)
         );
  MUX2_X1 U4822 ( .A(REG1_REG_27__SCAN_IN), .B(n4244), .S(n4610), .Z(U3545) );
  INV_X1 U4823 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4182) );
  AOI21_X1 U4824 ( .B1(n4181), .B2(n4577), .A(n4180), .ZN(n4245) );
  MUX2_X1 U4825 ( .A(n4182), .B(n4245), .S(n4610), .Z(n4183) );
  OAI21_X1 U4826 ( .B1(n4237), .B2(n4248), .A(n4183), .ZN(U3544) );
  INV_X1 U4827 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4857) );
  AOI21_X1 U4828 ( .B1(n4185), .B2(n4577), .A(n4184), .ZN(n4249) );
  MUX2_X1 U4829 ( .A(n4857), .B(n4249), .S(n4610), .Z(n4186) );
  OAI21_X1 U4830 ( .B1(n4237), .B2(n4251), .A(n4186), .ZN(U3543) );
  INV_X1 U4831 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4880) );
  AOI21_X1 U4832 ( .B1(n4188), .B2(n4577), .A(n4187), .ZN(n4252) );
  MUX2_X1 U4833 ( .A(n4880), .B(n4252), .S(n4610), .Z(n4189) );
  OAI21_X1 U4834 ( .B1(n4237), .B2(n4255), .A(n4189), .ZN(U3542) );
  INV_X1 U4835 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4192) );
  AOI21_X1 U4836 ( .B1(n4191), .B2(n4577), .A(n4190), .ZN(n4256) );
  MUX2_X1 U4837 ( .A(n4192), .B(n4256), .S(n4610), .Z(n4193) );
  OAI21_X1 U4838 ( .B1(n4237), .B2(n4258), .A(n4193), .ZN(U3541) );
  NAND3_X1 U4839 ( .A1(n4195), .A2(n4585), .A3(n4194), .ZN(n4196) );
  OAI211_X1 U4840 ( .C1(n4198), .C2(n4580), .A(n4197), .B(n4196), .ZN(n4259)
         );
  MUX2_X1 U4841 ( .A(REG1_REG_22__SCAN_IN), .B(n4259), .S(n4610), .Z(U3540) );
  NAND2_X1 U4842 ( .A1(n4199), .A2(n4585), .ZN(n4200) );
  OAI211_X1 U4843 ( .C1(n4202), .C2(n4580), .A(n4201), .B(n4200), .ZN(n4260)
         );
  MUX2_X1 U4844 ( .A(REG1_REG_21__SCAN_IN), .B(n4260), .S(n4610), .Z(U3539) );
  INV_X1 U4845 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4205) );
  AOI21_X1 U4846 ( .B1(n4204), .B2(n4577), .A(n4203), .ZN(n4261) );
  MUX2_X1 U4847 ( .A(n4205), .B(n4261), .S(n4610), .Z(n4206) );
  OAI21_X1 U4848 ( .B1(n4237), .B2(n4263), .A(n4206), .ZN(U3538) );
  INV_X1 U4849 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4209) );
  AOI21_X1 U4850 ( .B1(n4208), .B2(n4577), .A(n4207), .ZN(n4264) );
  MUX2_X1 U4851 ( .A(n4209), .B(n4264), .S(n4610), .Z(n4210) );
  OAI21_X1 U4852 ( .B1(n4237), .B2(n4266), .A(n4210), .ZN(U3537) );
  OAI211_X1 U4853 ( .C1(n4213), .C2(n4580), .A(n4212), .B(n4211), .ZN(n4267)
         );
  MUX2_X1 U4854 ( .A(REG1_REG_18__SCAN_IN), .B(n4267), .S(n4610), .Z(U3536) );
  AOI21_X1 U4855 ( .B1(n4215), .B2(n4577), .A(n4214), .ZN(n4268) );
  MUX2_X1 U4856 ( .A(n4216), .B(n4268), .S(n4610), .Z(n4217) );
  OAI21_X1 U4857 ( .B1(n4237), .B2(n4271), .A(n4217), .ZN(U3535) );
  NAND2_X1 U4858 ( .A1(n4218), .A2(n4585), .ZN(n4219) );
  OAI211_X1 U4859 ( .C1(n4221), .C2(n4580), .A(n4220), .B(n4219), .ZN(n4272)
         );
  MUX2_X1 U4860 ( .A(REG1_REG_16__SCAN_IN), .B(n4272), .S(n4610), .Z(U3534) );
  AOI21_X1 U4861 ( .B1(n4577), .B2(n4223), .A(n4222), .ZN(n4273) );
  MUX2_X1 U4862 ( .A(n4224), .B(n4273), .S(n4610), .Z(n4225) );
  OAI21_X1 U4863 ( .B1(n4237), .B2(n4276), .A(n4225), .ZN(U3533) );
  INV_X1 U4864 ( .A(n4226), .ZN(n4231) );
  NAND3_X1 U4865 ( .A1(n4228), .A2(n4585), .A3(n4227), .ZN(n4229) );
  OAI211_X1 U4866 ( .C1(n4231), .C2(n4562), .A(n4230), .B(n4229), .ZN(n4277)
         );
  MUX2_X1 U4867 ( .A(REG1_REG_14__SCAN_IN), .B(n4277), .S(n4610), .Z(U3532) );
  INV_X1 U4868 ( .A(n4562), .ZN(n4593) );
  INV_X1 U4869 ( .A(n4232), .ZN(n4234) );
  AOI21_X1 U4870 ( .B1(n4593), .B2(n4234), .A(n4233), .ZN(n4278) );
  MUX2_X1 U4871 ( .A(n4235), .B(n4278), .S(n4610), .Z(n4236) );
  OAI21_X1 U4872 ( .B1(n4237), .B2(n4282), .A(n4236), .ZN(U3531) );
  INV_X1 U4873 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4726) );
  MUX2_X1 U4874 ( .A(n4726), .B(n4334), .S(n4596), .Z(n4238) );
  OAI21_X1 U4875 ( .B1(n4239), .B2(n4281), .A(n4238), .ZN(U3517) );
  INV_X1 U4876 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4240) );
  NOR2_X1 U4877 ( .A1(n4596), .A2(n4240), .ZN(n4241) );
  AOI21_X1 U4878 ( .B1(n4596), .B2(n4336), .A(n4241), .ZN(n4242) );
  OAI21_X1 U4879 ( .B1(n4335), .B2(n4281), .A(n4242), .ZN(U3516) );
  MUX2_X1 U4880 ( .A(REG0_REG_29__SCAN_IN), .B(n4243), .S(n4596), .Z(U3515) );
  MUX2_X1 U4881 ( .A(REG0_REG_27__SCAN_IN), .B(n4244), .S(n4596), .Z(U3513) );
  INV_X1 U4882 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4246) );
  MUX2_X1 U4883 ( .A(n4246), .B(n4245), .S(n4596), .Z(n4247) );
  OAI21_X1 U4884 ( .B1(n4248), .B2(n4281), .A(n4247), .ZN(U3512) );
  INV_X1 U4885 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4727) );
  MUX2_X1 U4886 ( .A(n4727), .B(n4249), .S(n4596), .Z(n4250) );
  OAI21_X1 U4887 ( .B1(n4251), .B2(n4281), .A(n4250), .ZN(U3511) );
  INV_X1 U4888 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4253) );
  MUX2_X1 U4889 ( .A(n4253), .B(n4252), .S(n4596), .Z(n4254) );
  OAI21_X1 U4890 ( .B1(n4255), .B2(n4281), .A(n4254), .ZN(U3510) );
  INV_X1 U4891 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4723) );
  MUX2_X1 U4892 ( .A(n4723), .B(n4256), .S(n4596), .Z(n4257) );
  OAI21_X1 U4893 ( .B1(n4258), .B2(n4281), .A(n4257), .ZN(U3509) );
  MUX2_X1 U4894 ( .A(REG0_REG_22__SCAN_IN), .B(n4259), .S(n4596), .Z(U3508) );
  MUX2_X1 U4895 ( .A(REG0_REG_21__SCAN_IN), .B(n4260), .S(n4596), .Z(U3507) );
  INV_X1 U4896 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4720) );
  MUX2_X1 U4897 ( .A(n4720), .B(n4261), .S(n4596), .Z(n4262) );
  OAI21_X1 U4898 ( .B1(n4263), .B2(n4281), .A(n4262), .ZN(U3506) );
  INV_X1 U4899 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4721) );
  MUX2_X1 U4900 ( .A(n4721), .B(n4264), .S(n4596), .Z(n4265) );
  OAI21_X1 U4901 ( .B1(n4266), .B2(n4281), .A(n4265), .ZN(U3505) );
  MUX2_X1 U4902 ( .A(REG0_REG_18__SCAN_IN), .B(n4267), .S(n4596), .Z(U3503) );
  INV_X1 U4903 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4269) );
  MUX2_X1 U4904 ( .A(n4269), .B(n4268), .S(n4596), .Z(n4270) );
  OAI21_X1 U4905 ( .B1(n4271), .B2(n4281), .A(n4270), .ZN(U3501) );
  MUX2_X1 U4906 ( .A(REG0_REG_16__SCAN_IN), .B(n4272), .S(n4596), .Z(U3499) );
  INV_X1 U4907 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4274) );
  MUX2_X1 U4908 ( .A(n4274), .B(n4273), .S(n4596), .Z(n4275) );
  OAI21_X1 U4909 ( .B1(n4276), .B2(n4281), .A(n4275), .ZN(U3497) );
  MUX2_X1 U4910 ( .A(REG0_REG_14__SCAN_IN), .B(n4277), .S(n4596), .Z(U3495) );
  INV_X1 U4911 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4279) );
  MUX2_X1 U4912 ( .A(n4279), .B(n4278), .S(n4596), .Z(n4280) );
  OAI21_X1 U4913 ( .B1(n4282), .B2(n4281), .A(n4280), .ZN(U3493) );
  MUX2_X1 U4914 ( .A(DATAI_30_), .B(n4283), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4915 ( .A(n2468), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U4916 ( .A(n4339), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U4917 ( .A(n2809), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U4918 ( .A(n2942), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U4919 ( .A(n2771), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U4920 ( .A(DATAI_20_), .B(n4284), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4921 ( .A(DATAI_3_), .B(n4294), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U4922 ( .A(n4285), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4923 ( .A(n4286), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  OAI22_X1 U4924 ( .A1(U3149), .A2(n4287), .B1(DATAI_28_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4288) );
  INV_X1 U4925 ( .A(n4288), .ZN(U3324) );
  AOI21_X1 U4926 ( .B1(n4473), .B2(ADDR_REG_3__SCAN_IN), .A(n4289), .ZN(n4298)
         );
  OAI211_X1 U4927 ( .C1(REG1_REG_3__SCAN_IN), .C2(n4291), .A(n4481), .B(n4290), 
        .ZN(n4297) );
  OAI211_X1 U4928 ( .C1(REG2_REG_3__SCAN_IN), .C2(n4293), .A(n4483), .B(n4292), 
        .ZN(n4296) );
  NAND2_X1 U4929 ( .A1(n4458), .A2(n4294), .ZN(n4295) );
  NAND4_X1 U4930 ( .A1(n4298), .A2(n4297), .A3(n4296), .A4(n4295), .ZN(U3243)
         );
  OAI22_X1 U4931 ( .A1(n4300), .A2(n4315), .B1(n4316), .B2(n4299), .ZN(n4305)
         );
  NOR2_X1 U4932 ( .A1(STATE_REG_SCAN_IN), .A2(n4301), .ZN(n4462) );
  INV_X1 U4933 ( .A(n4462), .ZN(n4302) );
  OAI21_X1 U4934 ( .B1(n4318), .B2(n4303), .A(n4302), .ZN(n4304) );
  NOR2_X1 U4935 ( .A1(n4305), .A2(n4304), .ZN(n4312) );
  NAND2_X1 U4936 ( .A1(n4306), .A2(n4322), .ZN(n4307) );
  XOR2_X1 U4937 ( .A(n4308), .B(n4307), .Z(n4310) );
  NAND2_X1 U4938 ( .A1(n4310), .A2(n4309), .ZN(n4311) );
  OAI211_X1 U4939 ( .C1(n4331), .C2(n4313), .A(n4312), .B(n4311), .ZN(U3223)
         );
  OAI22_X1 U4940 ( .A1(n4989), .A2(n4316), .B1(n4315), .B2(n4314), .ZN(n4320)
         );
  INV_X1 U4941 ( .A(REG3_REG_15__SCAN_IN), .ZN(n4839) );
  OR2_X1 U4942 ( .A1(STATE_REG_SCAN_IN), .A2(n4839), .ZN(n4459) );
  OAI21_X1 U4943 ( .B1(n4318), .B2(n4317), .A(n4459), .ZN(n4319) );
  NOR2_X1 U4944 ( .A1(n4320), .A2(n4319), .ZN(n4329) );
  INV_X1 U4945 ( .A(n4322), .ZN(n4327) );
  AOI21_X1 U4946 ( .B1(n4323), .B2(n4322), .A(n4321), .ZN(n4325) );
  NOR2_X1 U4947 ( .A1(n4325), .A2(n4324), .ZN(n4326) );
  OAI21_X1 U4948 ( .B1(n4327), .B2(n4306), .A(n4326), .ZN(n4328) );
  OAI211_X1 U4949 ( .C1(n4331), .C2(n4330), .A(n4329), .B(n4328), .ZN(U3238)
         );
  AOI22_X1 U4950 ( .A1(n4332), .A2(n4513), .B1(n4519), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4333) );
  OAI21_X1 U4951 ( .B1(n4519), .B2(n4334), .A(n4333), .ZN(U3260) );
  INV_X1 U4952 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4751) );
  INV_X1 U4953 ( .A(n4340), .ZN(n4338) );
  OAI211_X1 U4954 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4339), .A(n4341), .B(n4338), 
        .ZN(n4344) );
  AOI22_X1 U4955 ( .A1(n4341), .A2(n4340), .B1(n4481), .B2(n2951), .ZN(n4343)
         );
  AOI22_X1 U4956 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4473), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4342) );
  OAI221_X1 U4957 ( .B1(IR_REG_0__SCAN_IN), .B2(n4344), .C1(n2498), .C2(n4343), 
        .A(n4342), .ZN(U3240) );
  NAND2_X1 U4958 ( .A1(n4458), .A2(n4345), .ZN(n4354) );
  XNOR2_X1 U4959 ( .A(n4346), .B(REG1_REG_4__SCAN_IN), .ZN(n4347) );
  NAND2_X1 U4960 ( .A1(n4481), .A2(n4347), .ZN(n4353) );
  XNOR2_X1 U4961 ( .A(n4348), .B(REG2_REG_4__SCAN_IN), .ZN(n4349) );
  NAND2_X1 U4962 ( .A1(n4483), .A2(n4349), .ZN(n4352) );
  AOI21_X1 U4963 ( .B1(n4473), .B2(ADDR_REG_4__SCAN_IN), .A(n4350), .ZN(n4351)
         );
  AND4_X1 U4964 ( .A1(n4354), .A2(n4353), .A3(n4352), .A4(n4351), .ZN(n4356)
         );
  NAND2_X1 U4965 ( .A1(n4356), .A2(n4355), .ZN(U3244) );
  INV_X1 U4966 ( .A(n4473), .ZN(n4461) );
  INV_X1 U4967 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n4893) );
  OAI211_X1 U4968 ( .C1(n4359), .C2(n4358), .A(n4483), .B(n4357), .ZN(n4360)
         );
  OAI21_X1 U4969 ( .B1(n4461), .B2(n4893), .A(n4360), .ZN(n4361) );
  NOR2_X1 U4970 ( .A1(n4362), .A2(n4361), .ZN(n4367) );
  OAI211_X1 U4971 ( .C1(n4365), .C2(n4364), .A(n4481), .B(n4363), .ZN(n4366)
         );
  OAI211_X1 U4972 ( .C1(n4486), .C2(n4542), .A(n4367), .B(n4366), .ZN(U3245)
         );
  AOI21_X1 U4973 ( .B1(n4473), .B2(ADDR_REG_6__SCAN_IN), .A(n4368), .ZN(n4376)
         );
  OAI211_X1 U4974 ( .C1(REG1_REG_6__SCAN_IN), .C2(n4370), .A(n4481), .B(n4369), 
        .ZN(n4375) );
  OAI211_X1 U4975 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4372), .A(n4483), .B(n4371), 
        .ZN(n4374) );
  NAND2_X1 U4976 ( .A1(n4540), .A2(n4458), .ZN(n4373) );
  NAND4_X1 U4977 ( .A1(n4376), .A2(n4375), .A3(n4374), .A4(n4373), .ZN(U3246)
         );
  AOI21_X1 U4978 ( .B1(n4604), .B2(n4539), .A(n4377), .ZN(n4379) );
  XOR2_X1 U4979 ( .A(n4379), .B(n4378), .Z(n4386) );
  INV_X1 U4980 ( .A(ADDR_REG_7__SCAN_IN), .ZN(n4753) );
  OAI211_X1 U4981 ( .C1(n4382), .C2(n4381), .A(n4483), .B(n4380), .ZN(n4383)
         );
  OAI211_X1 U4982 ( .C1(n4461), .C2(n4753), .A(n4384), .B(n4383), .ZN(n4385)
         );
  AOI21_X1 U4983 ( .B1(n4386), .B2(n4481), .A(n4385), .ZN(n4387) );
  OAI21_X1 U4984 ( .B1(n4539), .B2(n4486), .A(n4387), .ZN(U3247) );
  AOI211_X1 U4985 ( .C1(n4390), .C2(n4389), .A(n4388), .B(n4447), .ZN(n4392)
         );
  AOI211_X1 U4986 ( .C1(n4473), .C2(ADDR_REG_8__SCAN_IN), .A(n4392), .B(n4391), 
        .ZN(n4396) );
  OAI211_X1 U4987 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4394), .A(n4483), .B(n4393), 
        .ZN(n4395) );
  OAI211_X1 U4988 ( .C1(n4486), .C2(n4537), .A(n4396), .B(n4395), .ZN(U3248)
         );
  AOI211_X1 U4989 ( .C1(n2255), .C2(n4398), .A(n4397), .B(n4447), .ZN(n4400)
         );
  AOI211_X1 U4990 ( .C1(n4473), .C2(ADDR_REG_9__SCAN_IN), .A(n4400), .B(n4399), 
        .ZN(n4405) );
  OAI211_X1 U4991 ( .C1(n4403), .C2(n4402), .A(n4483), .B(n4401), .ZN(n4404)
         );
  OAI211_X1 U4992 ( .C1(n4486), .C2(n4406), .A(n4405), .B(n4404), .ZN(U3249)
         );
  AOI211_X1 U4993 ( .C1(n2256), .C2(n4408), .A(n4407), .B(n4447), .ZN(n4411)
         );
  INV_X1 U4994 ( .A(n4409), .ZN(n4410) );
  AOI211_X1 U4995 ( .C1(n4473), .C2(ADDR_REG_11__SCAN_IN), .A(n4411), .B(n4410), .ZN(n4416) );
  OAI211_X1 U4996 ( .C1(n4414), .C2(n4413), .A(n4483), .B(n4412), .ZN(n4415)
         );
  OAI211_X1 U4997 ( .C1(n4486), .C2(n4534), .A(n4416), .B(n4415), .ZN(U3251)
         );
  AOI211_X1 U4998 ( .C1(n4419), .C2(n4418), .A(n4417), .B(n4447), .ZN(n4422)
         );
  INV_X1 U4999 ( .A(n4420), .ZN(n4421) );
  AOI211_X1 U5000 ( .C1(n4473), .C2(ADDR_REG_12__SCAN_IN), .A(n4422), .B(n4421), .ZN(n4426) );
  OAI211_X1 U5001 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4424), .A(n4483), .B(n4423), .ZN(n4425) );
  OAI211_X1 U5002 ( .C1(n4486), .C2(n4427), .A(n4426), .B(n4425), .ZN(U3252)
         );
  AOI211_X1 U5003 ( .C1(n2245), .C2(n4429), .A(n4428), .B(n4447), .ZN(n4430)
         );
  AOI211_X1 U5004 ( .C1(n4473), .C2(ADDR_REG_13__SCAN_IN), .A(n4431), .B(n4430), .ZN(n4437) );
  AOI21_X1 U5005 ( .B1(n3303), .B2(n4530), .A(n4432), .ZN(n4435) );
  INV_X1 U5006 ( .A(n4483), .ZN(n4451) );
  AOI21_X1 U5007 ( .B1(n4435), .B2(n4434), .A(n4451), .ZN(n4433) );
  OAI21_X1 U5008 ( .B1(n4435), .B2(n4434), .A(n4433), .ZN(n4436) );
  OAI211_X1 U5009 ( .C1(n4486), .C2(n4530), .A(n4437), .B(n4436), .ZN(U3253)
         );
  INV_X1 U5010 ( .A(ADDR_REG_14__SCAN_IN), .ZN(n4754) );
  AOI211_X1 U5011 ( .C1(n4873), .C2(n4439), .A(n4438), .B(n4447), .ZN(n4443)
         );
  AOI211_X1 U5012 ( .C1(n3318), .C2(n4441), .A(n4440), .B(n4451), .ZN(n4442)
         );
  AOI211_X1 U5013 ( .C1(n4458), .C2(n4444), .A(n4443), .B(n4442), .ZN(n4446)
         );
  OAI211_X1 U5014 ( .C1(n4461), .C2(n4754), .A(n4446), .B(n4445), .ZN(U3254)
         );
  INV_X1 U5015 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n4806) );
  AOI211_X1 U5016 ( .C1(n4450), .C2(n4449), .A(n4448), .B(n4447), .ZN(n4456)
         );
  AOI211_X1 U5017 ( .C1(n4454), .C2(n4453), .A(n4452), .B(n4451), .ZN(n4455)
         );
  AOI211_X1 U5018 ( .C1(n4458), .C2(n4457), .A(n4456), .B(n4455), .ZN(n4460)
         );
  OAI211_X1 U5019 ( .C1(n4461), .C2(n4806), .A(n4460), .B(n4459), .ZN(U3255)
         );
  AOI21_X1 U5020 ( .B1(n4473), .B2(ADDR_REG_16__SCAN_IN), .A(n4462), .ZN(n4471) );
  OAI21_X1 U5021 ( .B1(n4465), .B2(n4464), .A(n4463), .ZN(n4469) );
  OAI21_X1 U5022 ( .B1(n4467), .B2(n4855), .A(n4466), .ZN(n4468) );
  AOI22_X1 U5023 ( .A1(n4483), .A2(n4469), .B1(n4481), .B2(n4468), .ZN(n4470)
         );
  OAI211_X1 U5024 ( .C1(n4527), .C2(n4486), .A(n4471), .B(n4470), .ZN(U3256)
         );
  AOI21_X1 U5025 ( .B1(n4473), .B2(ADDR_REG_17__SCAN_IN), .A(n4472), .ZN(n4485) );
  OAI21_X1 U5026 ( .B1(n4476), .B2(n4475), .A(n4474), .ZN(n4482) );
  OAI21_X1 U5027 ( .B1(n4479), .B2(n4478), .A(n4477), .ZN(n4480) );
  AOI22_X1 U5028 ( .A1(n4483), .A2(n4482), .B1(n4481), .B2(n4480), .ZN(n4484)
         );
  OAI211_X1 U5029 ( .C1(n4525), .C2(n4486), .A(n4485), .B(n4484), .ZN(U3257)
         );
  XNOR2_X1 U5030 ( .A(n4487), .B(n4489), .ZN(n4592) );
  XOR2_X1 U5031 ( .A(n4489), .B(n4488), .Z(n4498) );
  OAI22_X1 U5032 ( .A1(n4492), .A2(n4491), .B1(n4503), .B2(n4490), .ZN(n4493)
         );
  AOI21_X1 U5033 ( .B1(n4495), .B2(n4494), .A(n4493), .ZN(n4496) );
  OAI21_X1 U5034 ( .B1(n4498), .B2(n4497), .A(n4496), .ZN(n4499) );
  AOI21_X1 U5035 ( .B1(n4500), .B2(n4592), .A(n4499), .ZN(n4589) );
  AOI22_X1 U5036 ( .A1(n4501), .A2(n4508), .B1(REG2_REG_11__SCAN_IN), .B2(
        n4519), .ZN(n4507) );
  OAI21_X1 U5037 ( .B1(n4504), .B2(n4503), .A(n4502), .ZN(n4588) );
  INV_X1 U5038 ( .A(n4588), .ZN(n4505) );
  AOI22_X1 U5039 ( .A1(n4592), .A2(n4514), .B1(n4513), .B2(n4505), .ZN(n4506)
         );
  OAI211_X1 U5040 ( .C1(n4519), .C2(n4589), .A(n4507), .B(n4506), .ZN(U3279)
         );
  AOI22_X1 U5041 ( .A1(n4509), .A2(n4508), .B1(REG2_REG_6__SCAN_IN), .B2(n4519), .ZN(n4517) );
  INV_X1 U5042 ( .A(n4510), .ZN(n4515) );
  INV_X1 U5043 ( .A(n4511), .ZN(n4512) );
  AOI22_X1 U5044 ( .A1(n4515), .A2(n4514), .B1(n4513), .B2(n4512), .ZN(n4516)
         );
  OAI211_X1 U5045 ( .C1(n4519), .C2(n4518), .A(n4517), .B(n4516), .ZN(U3284)
         );
  AND2_X1 U5046 ( .A1(D_REG_31__SCAN_IN), .A2(n4521), .ZN(U3291) );
  AND2_X1 U5047 ( .A1(n4521), .A2(D_REG_30__SCAN_IN), .ZN(U3292) );
  AND2_X1 U5048 ( .A1(D_REG_29__SCAN_IN), .A2(n4521), .ZN(U3293) );
  AND2_X1 U5049 ( .A1(D_REG_28__SCAN_IN), .A2(n4521), .ZN(U3294) );
  AND2_X1 U5050 ( .A1(D_REG_27__SCAN_IN), .A2(n4521), .ZN(U3295) );
  AND2_X1 U5051 ( .A1(n4521), .A2(D_REG_26__SCAN_IN), .ZN(U3296) );
  INV_X1 U5052 ( .A(D_REG_25__SCAN_IN), .ZN(n4835) );
  NOR2_X1 U5053 ( .A1(n4520), .A2(n4835), .ZN(U3297) );
  AND2_X1 U5054 ( .A1(D_REG_24__SCAN_IN), .A2(n4521), .ZN(U3298) );
  INV_X1 U5055 ( .A(D_REG_23__SCAN_IN), .ZN(n4854) );
  NOR2_X1 U5056 ( .A1(n4520), .A2(n4854), .ZN(U3299) );
  AND2_X1 U5057 ( .A1(D_REG_22__SCAN_IN), .A2(n4521), .ZN(U3300) );
  INV_X1 U5058 ( .A(D_REG_21__SCAN_IN), .ZN(n4858) );
  NOR2_X1 U5059 ( .A1(n4520), .A2(n4858), .ZN(U3301) );
  AND2_X1 U5060 ( .A1(D_REG_20__SCAN_IN), .A2(n4521), .ZN(U3302) );
  AND2_X1 U5061 ( .A1(D_REG_19__SCAN_IN), .A2(n4521), .ZN(U3303) );
  AND2_X1 U5062 ( .A1(D_REG_18__SCAN_IN), .A2(n4521), .ZN(U3304) );
  AND2_X1 U5063 ( .A1(D_REG_17__SCAN_IN), .A2(n4521), .ZN(U3305) );
  INV_X1 U5064 ( .A(D_REG_16__SCAN_IN), .ZN(n4709) );
  NOR2_X1 U5065 ( .A1(n4520), .A2(n4709), .ZN(U3306) );
  AND2_X1 U5066 ( .A1(n4521), .A2(D_REG_15__SCAN_IN), .ZN(U3307) );
  AND2_X1 U5067 ( .A1(D_REG_14__SCAN_IN), .A2(n4521), .ZN(U3308) );
  INV_X1 U5068 ( .A(D_REG_13__SCAN_IN), .ZN(n4805) );
  NOR2_X1 U5069 ( .A1(n4520), .A2(n4805), .ZN(U3309) );
  AND2_X1 U5070 ( .A1(D_REG_12__SCAN_IN), .A2(n4521), .ZN(U3310) );
  AND2_X1 U5071 ( .A1(D_REG_11__SCAN_IN), .A2(n4521), .ZN(U3311) );
  AND2_X1 U5072 ( .A1(D_REG_10__SCAN_IN), .A2(n4521), .ZN(U3312) );
  AND2_X1 U5073 ( .A1(D_REG_9__SCAN_IN), .A2(n4521), .ZN(U3313) );
  AND2_X1 U5074 ( .A1(n4521), .A2(D_REG_8__SCAN_IN), .ZN(U3314) );
  AND2_X1 U5075 ( .A1(D_REG_7__SCAN_IN), .A2(n4521), .ZN(U3315) );
  AND2_X1 U5076 ( .A1(D_REG_6__SCAN_IN), .A2(n4521), .ZN(U3316) );
  INV_X1 U5077 ( .A(D_REG_5__SCAN_IN), .ZN(n4820) );
  NOR2_X1 U5078 ( .A1(n4520), .A2(n4820), .ZN(U3317) );
  AND2_X1 U5079 ( .A1(D_REG_4__SCAN_IN), .A2(n4521), .ZN(U3318) );
  AND2_X1 U5080 ( .A1(D_REG_3__SCAN_IN), .A2(n4521), .ZN(U3319) );
  AND2_X1 U5081 ( .A1(n4521), .A2(D_REG_2__SCAN_IN), .ZN(U3320) );
  INV_X1 U5082 ( .A(DATAI_23_), .ZN(n4523) );
  AOI21_X1 U5083 ( .B1(U3149), .B2(n4523), .A(n4522), .ZN(U3329) );
  INV_X1 U5084 ( .A(DATAI_17_), .ZN(n4524) );
  AOI22_X1 U5085 ( .A1(STATE_REG_SCAN_IN), .A2(n4525), .B1(n4524), .B2(U3149), 
        .ZN(U3335) );
  AOI22_X1 U5086 ( .A1(STATE_REG_SCAN_IN), .A2(n4527), .B1(n4526), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5087 ( .A(DATAI_15_), .ZN(n4808) );
  AOI22_X1 U5088 ( .A1(STATE_REG_SCAN_IN), .A2(n4528), .B1(n4808), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5089 ( .A(DATAI_14_), .ZN(n4678) );
  AOI22_X1 U5090 ( .A1(STATE_REG_SCAN_IN), .A2(n4529), .B1(n4678), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U5091 ( .A1(STATE_REG_SCAN_IN), .A2(n4530), .B1(n4884), .B2(U3149), 
        .ZN(U3339) );
  OAI22_X1 U5092 ( .A1(U3149), .A2(n4531), .B1(DATAI_12_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4532) );
  INV_X1 U5093 ( .A(n4532), .ZN(U3340) );
  INV_X1 U5094 ( .A(DATAI_11_), .ZN(n4533) );
  AOI22_X1 U5095 ( .A1(STATE_REG_SCAN_IN), .A2(n4534), .B1(n4533), .B2(U3149), 
        .ZN(U3341) );
  OAI22_X1 U5096 ( .A1(U3149), .A2(n4535), .B1(DATAI_9_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4536) );
  INV_X1 U5097 ( .A(n4536), .ZN(U3343) );
  AOI22_X1 U5098 ( .A1(STATE_REG_SCAN_IN), .A2(n4537), .B1(n2558), .B2(U3149), 
        .ZN(U3344) );
  INV_X1 U5099 ( .A(DATAI_7_), .ZN(n4538) );
  AOI22_X1 U5100 ( .A1(STATE_REG_SCAN_IN), .A2(n4539), .B1(n4538), .B2(U3149), 
        .ZN(U3345) );
  OAI22_X1 U5101 ( .A1(U3149), .A2(n4540), .B1(DATAI_6_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4541) );
  INV_X1 U5102 ( .A(n4541), .ZN(U3346) );
  INV_X1 U5103 ( .A(DATAI_5_), .ZN(n4677) );
  AOI22_X1 U5104 ( .A1(STATE_REG_SCAN_IN), .A2(n4542), .B1(n4677), .B2(U3149), 
        .ZN(U3347) );
  INV_X1 U5105 ( .A(DATAI_0_), .ZN(n4543) );
  AOI22_X1 U5106 ( .A1(STATE_REG_SCAN_IN), .A2(n2498), .B1(n4543), .B2(U3149), 
        .ZN(U3352) );
  AOI22_X1 U5107 ( .A1(n4546), .A2(n4593), .B1(n4545), .B2(n4544), .ZN(n4547)
         );
  AND2_X1 U5108 ( .A1(n4548), .A2(n4547), .ZN(n4597) );
  INV_X1 U5109 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4549) );
  AOI22_X1 U5110 ( .A1(n4596), .A2(n4597), .B1(n4549), .B2(n4594), .ZN(U3467)
         );
  NOR2_X1 U5111 ( .A1(n4550), .A2(n4562), .ZN(n4552) );
  AOI211_X1 U5112 ( .C1(n4585), .C2(n4553), .A(n4552), .B(n4551), .ZN(n4598)
         );
  INV_X1 U5113 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4554) );
  AOI22_X1 U5114 ( .A1(n4596), .A2(n4598), .B1(n4554), .B2(n4594), .ZN(U3469)
         );
  NOR3_X1 U5115 ( .A1(n4556), .A2(n4555), .A3(n4587), .ZN(n4558) );
  AOI211_X1 U5116 ( .C1(n4593), .C2(n4559), .A(n4558), .B(n4557), .ZN(n4599)
         );
  INV_X1 U5117 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4560) );
  AOI22_X1 U5118 ( .A1(n4596), .A2(n4599), .B1(n4560), .B2(n4594), .ZN(U3471)
         );
  OAI22_X1 U5119 ( .A1(n4563), .A2(n4562), .B1(n4587), .B2(n4561), .ZN(n4564)
         );
  NOR2_X1 U5120 ( .A1(n4565), .A2(n4564), .ZN(n4601) );
  INV_X1 U5121 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4836) );
  AOI22_X1 U5122 ( .A1(n4596), .A2(n4601), .B1(n4836), .B2(n4594), .ZN(U3473)
         );
  INV_X1 U5123 ( .A(n4566), .ZN(n4568) );
  AOI211_X1 U5124 ( .C1(n4569), .C2(n4593), .A(n4568), .B(n4567), .ZN(n4602)
         );
  INV_X1 U5125 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4711) );
  AOI22_X1 U5126 ( .A1(n4596), .A2(n4602), .B1(n4711), .B2(n4594), .ZN(U3475)
         );
  NOR2_X1 U5127 ( .A1(n4570), .A2(n4580), .ZN(n4571) );
  AOI211_X1 U5128 ( .C1(n4585), .C2(n4573), .A(n4572), .B(n4571), .ZN(n4603)
         );
  INV_X1 U5129 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4574) );
  AOI22_X1 U5130 ( .A1(n4596), .A2(n4603), .B1(n4574), .B2(n4594), .ZN(U3477)
         );
  AOI211_X1 U5131 ( .C1(n4578), .C2(n4577), .A(n4576), .B(n4575), .ZN(n4605)
         );
  INV_X1 U5132 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4579) );
  AOI22_X1 U5133 ( .A1(n4596), .A2(n4605), .B1(n4579), .B2(n4594), .ZN(U3481)
         );
  NOR2_X1 U5134 ( .A1(n4581), .A2(n4580), .ZN(n4583) );
  AOI211_X1 U5135 ( .C1(n4585), .C2(n4584), .A(n4583), .B(n4582), .ZN(n4606)
         );
  INV_X1 U5136 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4586) );
  AOI22_X1 U5137 ( .A1(n4596), .A2(n4606), .B1(n4586), .B2(n4594), .ZN(U3485)
         );
  NOR2_X1 U5138 ( .A1(n4588), .A2(n4587), .ZN(n4591) );
  INV_X1 U5139 ( .A(n4589), .ZN(n4590) );
  AOI211_X1 U5140 ( .C1(n4593), .C2(n4592), .A(n4591), .B(n4590), .ZN(n4609)
         );
  INV_X1 U5141 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4595) );
  AOI22_X1 U5142 ( .A1(n4596), .A2(n4609), .B1(n4595), .B2(n4594), .ZN(U3489)
         );
  AOI22_X1 U5143 ( .A1(n4610), .A2(n4597), .B1(n2951), .B2(n4607), .ZN(U3518)
         );
  AOI22_X1 U5144 ( .A1(n4610), .A2(n4598), .B1(n2872), .B2(n4607), .ZN(U3519)
         );
  AOI22_X1 U5145 ( .A1(n4610), .A2(n4599), .B1(n4852), .B2(n4607), .ZN(U3520)
         );
  INV_X1 U5146 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4600) );
  AOI22_X1 U5147 ( .A1(n4610), .A2(n4601), .B1(n4600), .B2(n4607), .ZN(U3521)
         );
  AOI22_X1 U5148 ( .A1(n4610), .A2(n4602), .B1(n2879), .B2(n4607), .ZN(U3522)
         );
  AOI22_X1 U5149 ( .A1(n4610), .A2(n4603), .B1(n4896), .B2(n4607), .ZN(U3523)
         );
  AOI22_X1 U5150 ( .A1(n4610), .A2(n4605), .B1(n4604), .B2(n4607), .ZN(U3525)
         );
  INV_X1 U5151 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4810) );
  AOI22_X1 U5152 ( .A1(n4610), .A2(n4606), .B1(n4810), .B2(n4607), .ZN(U3527)
         );
  AOI22_X1 U5153 ( .A1(n4610), .A2(n4609), .B1(n4608), .B2(n4607), .ZN(U3529)
         );
  AOI22_X1 U5154 ( .A1(DATAI_18_), .A2(keyinput197), .B1(DATAI_28_), .B2(
        keyinput202), .ZN(n4611) );
  OAI221_X1 U5155 ( .B1(DATAI_18_), .B2(keyinput197), .C1(DATAI_28_), .C2(
        keyinput202), .A(n4611), .ZN(n4618) );
  AOI22_X1 U5156 ( .A1(DATAI_10_), .A2(keyinput150), .B1(DATAI_15_), .B2(
        keyinput188), .ZN(n4612) );
  OAI221_X1 U5157 ( .B1(DATAI_10_), .B2(keyinput150), .C1(DATAI_15_), .C2(
        keyinput188), .A(n4612), .ZN(n4617) );
  AOI22_X1 U5158 ( .A1(DATAI_4_), .A2(keyinput171), .B1(DATAI_3_), .B2(
        keyinput145), .ZN(n4613) );
  OAI221_X1 U5159 ( .B1(DATAI_4_), .B2(keyinput171), .C1(DATAI_3_), .C2(
        keyinput145), .A(n4613), .ZN(n4616) );
  AOI22_X1 U5160 ( .A1(REG3_REG_7__SCAN_IN), .A2(keyinput130), .B1(
        STATE_REG_SCAN_IN), .B2(keyinput165), .ZN(n4614) );
  OAI221_X1 U5161 ( .B1(REG3_REG_7__SCAN_IN), .B2(keyinput130), .C1(
        STATE_REG_SCAN_IN), .C2(keyinput165), .A(n4614), .ZN(n4615) );
  NOR4_X1 U5162 ( .A1(n4618), .A2(n4617), .A3(n4616), .A4(n4615), .ZN(n4646)
         );
  AOI22_X1 U5163 ( .A1(REG3_REG_23__SCAN_IN), .A2(keyinput233), .B1(
        REG3_REG_28__SCAN_IN), .B2(keyinput203), .ZN(n4619) );
  OAI221_X1 U5164 ( .B1(REG3_REG_23__SCAN_IN), .B2(keyinput233), .C1(
        REG3_REG_28__SCAN_IN), .C2(keyinput203), .A(n4619), .ZN(n4626) );
  AOI22_X1 U5165 ( .A1(REG3_REG_12__SCAN_IN), .A2(keyinput154), .B1(
        REG3_REG_16__SCAN_IN), .B2(keyinput177), .ZN(n4620) );
  OAI221_X1 U5166 ( .B1(REG3_REG_12__SCAN_IN), .B2(keyinput154), .C1(
        REG3_REG_16__SCAN_IN), .C2(keyinput177), .A(n4620), .ZN(n4625) );
  AOI22_X1 U5167 ( .A1(IR_REG_6__SCAN_IN), .A2(keyinput160), .B1(
        IR_REG_7__SCAN_IN), .B2(keyinput191), .ZN(n4621) );
  OAI221_X1 U5168 ( .B1(IR_REG_6__SCAN_IN), .B2(keyinput160), .C1(
        IR_REG_7__SCAN_IN), .C2(keyinput191), .A(n4621), .ZN(n4624) );
  AOI22_X1 U5169 ( .A1(IR_REG_8__SCAN_IN), .A2(keyinput139), .B1(
        IR_REG_14__SCAN_IN), .B2(keyinput254), .ZN(n4622) );
  OAI221_X1 U5170 ( .B1(IR_REG_8__SCAN_IN), .B2(keyinput139), .C1(
        IR_REG_14__SCAN_IN), .C2(keyinput254), .A(n4622), .ZN(n4623) );
  NOR4_X1 U5171 ( .A1(n4626), .A2(n4625), .A3(n4624), .A4(n4623), .ZN(n4645)
         );
  AOI22_X1 U5172 ( .A1(IR_REG_28__SCAN_IN), .A2(keyinput137), .B1(
        IR_REG_25__SCAN_IN), .B2(keyinput209), .ZN(n4627) );
  OAI221_X1 U5173 ( .B1(IR_REG_28__SCAN_IN), .B2(keyinput137), .C1(
        IR_REG_25__SCAN_IN), .C2(keyinput209), .A(n4627), .ZN(n4634) );
  AOI22_X1 U5174 ( .A1(D_REG_0__SCAN_IN), .A2(keyinput170), .B1(
        IR_REG_31__SCAN_IN), .B2(keyinput243), .ZN(n4628) );
  OAI221_X1 U5175 ( .B1(D_REG_0__SCAN_IN), .B2(keyinput170), .C1(
        IR_REG_31__SCAN_IN), .C2(keyinput243), .A(n4628), .ZN(n4633) );
  AOI22_X1 U5176 ( .A1(D_REG_5__SCAN_IN), .A2(keyinput224), .B1(
        D_REG_2__SCAN_IN), .B2(keyinput128), .ZN(n4629) );
  OAI221_X1 U5177 ( .B1(D_REG_5__SCAN_IN), .B2(keyinput224), .C1(
        D_REG_2__SCAN_IN), .C2(keyinput128), .A(n4629), .ZN(n4632) );
  AOI22_X1 U5178 ( .A1(D_REG_23__SCAN_IN), .A2(keyinput186), .B1(
        D_REG_15__SCAN_IN), .B2(keyinput178), .ZN(n4630) );
  OAI221_X1 U5179 ( .B1(D_REG_23__SCAN_IN), .B2(keyinput186), .C1(
        D_REG_15__SCAN_IN), .C2(keyinput178), .A(n4630), .ZN(n4631) );
  NOR4_X1 U5180 ( .A1(n4634), .A2(n4633), .A3(n4632), .A4(n4631), .ZN(n4644)
         );
  AOI22_X1 U5181 ( .A1(D_REG_21__SCAN_IN), .A2(keyinput206), .B1(
        D_REG_26__SCAN_IN), .B2(keyinput201), .ZN(n4635) );
  OAI221_X1 U5182 ( .B1(D_REG_21__SCAN_IN), .B2(keyinput206), .C1(
        D_REG_26__SCAN_IN), .C2(keyinput201), .A(n4635), .ZN(n4642) );
  AOI22_X1 U5183 ( .A1(REG0_REG_0__SCAN_IN), .A2(keyinput227), .B1(
        D_REG_30__SCAN_IN), .B2(keyinput208), .ZN(n4636) );
  OAI221_X1 U5184 ( .B1(REG0_REG_0__SCAN_IN), .B2(keyinput227), .C1(
        D_REG_30__SCAN_IN), .C2(keyinput208), .A(n4636), .ZN(n4641) );
  AOI22_X1 U5185 ( .A1(REG0_REG_1__SCAN_IN), .A2(keyinput249), .B1(
        REG0_REG_5__SCAN_IN), .B2(keyinput168), .ZN(n4637) );
  OAI221_X1 U5186 ( .B1(REG0_REG_1__SCAN_IN), .B2(keyinput249), .C1(
        REG0_REG_5__SCAN_IN), .C2(keyinput168), .A(n4637), .ZN(n4640) );
  AOI22_X1 U5187 ( .A1(REG0_REG_18__SCAN_IN), .A2(keyinput158), .B1(
        REG0_REG_13__SCAN_IN), .B2(keyinput235), .ZN(n4638) );
  OAI221_X1 U5188 ( .B1(REG0_REG_18__SCAN_IN), .B2(keyinput158), .C1(
        REG0_REG_13__SCAN_IN), .C2(keyinput235), .A(n4638), .ZN(n4639) );
  NOR4_X1 U5189 ( .A1(n4642), .A2(n4641), .A3(n4640), .A4(n4639), .ZN(n4643)
         );
  NAND4_X1 U5190 ( .A1(n4646), .A2(n4645), .A3(n4644), .A4(n4643), .ZN(n4788)
         );
  AOI22_X1 U5191 ( .A1(REG1_REG_0__SCAN_IN), .A2(keyinput195), .B1(
        REG1_REG_2__SCAN_IN), .B2(keyinput183), .ZN(n4647) );
  OAI221_X1 U5192 ( .B1(REG1_REG_0__SCAN_IN), .B2(keyinput195), .C1(
        REG1_REG_2__SCAN_IN), .C2(keyinput183), .A(n4647), .ZN(n4654) );
  AOI22_X1 U5193 ( .A1(REG1_REG_4__SCAN_IN), .A2(keyinput135), .B1(
        REG1_REG_3__SCAN_IN), .B2(keyinput250), .ZN(n4648) );
  OAI221_X1 U5194 ( .B1(REG1_REG_4__SCAN_IN), .B2(keyinput135), .C1(
        REG1_REG_3__SCAN_IN), .C2(keyinput250), .A(n4648), .ZN(n4653) );
  AOI22_X1 U5195 ( .A1(REG1_REG_5__SCAN_IN), .A2(keyinput153), .B1(
        REG1_REG_6__SCAN_IN), .B2(keyinput222), .ZN(n4649) );
  OAI221_X1 U5196 ( .B1(REG1_REG_5__SCAN_IN), .B2(keyinput153), .C1(
        REG1_REG_6__SCAN_IN), .C2(keyinput222), .A(n4649), .ZN(n4652) );
  AOI22_X1 U5197 ( .A1(REG1_REG_9__SCAN_IN), .A2(keyinput232), .B1(
        REG1_REG_10__SCAN_IN), .B2(keyinput215), .ZN(n4650) );
  OAI221_X1 U5198 ( .B1(REG1_REG_9__SCAN_IN), .B2(keyinput232), .C1(
        REG1_REG_10__SCAN_IN), .C2(keyinput215), .A(n4650), .ZN(n4651) );
  NOR4_X1 U5199 ( .A1(n4654), .A2(n4653), .A3(n4652), .A4(n4651), .ZN(n4686)
         );
  AOI22_X1 U5200 ( .A1(REG2_REG_9__SCAN_IN), .A2(keyinput163), .B1(
        REG1_REG_14__SCAN_IN), .B2(keyinput159), .ZN(n4655) );
  OAI221_X1 U5201 ( .B1(REG2_REG_9__SCAN_IN), .B2(keyinput163), .C1(
        REG1_REG_14__SCAN_IN), .C2(keyinput159), .A(n4655), .ZN(n4662) );
  AOI22_X1 U5202 ( .A1(REG2_REG_19__SCAN_IN), .A2(keyinput169), .B1(
        REG2_REG_25__SCAN_IN), .B2(keyinput142), .ZN(n4656) );
  OAI221_X1 U5203 ( .B1(REG2_REG_19__SCAN_IN), .B2(keyinput169), .C1(
        REG2_REG_25__SCAN_IN), .C2(keyinput142), .A(n4656), .ZN(n4661) );
  AOI22_X1 U5204 ( .A1(ADDR_REG_15__SCAN_IN), .A2(keyinput156), .B1(
        ADDR_REG_17__SCAN_IN), .B2(keyinput133), .ZN(n4657) );
  OAI221_X1 U5205 ( .B1(ADDR_REG_15__SCAN_IN), .B2(keyinput156), .C1(
        ADDR_REG_17__SCAN_IN), .C2(keyinput133), .A(n4657), .ZN(n4660) );
  AOI22_X1 U5206 ( .A1(ADDR_REG_3__SCAN_IN), .A2(keyinput205), .B1(
        ADDR_REG_12__SCAN_IN), .B2(keyinput230), .ZN(n4658) );
  OAI221_X1 U5207 ( .B1(ADDR_REG_3__SCAN_IN), .B2(keyinput205), .C1(
        ADDR_REG_12__SCAN_IN), .C2(keyinput230), .A(n4658), .ZN(n4659) );
  NOR4_X1 U5208 ( .A1(n4662), .A2(n4661), .A3(n4660), .A4(n4659), .ZN(n4685)
         );
  AOI22_X1 U5209 ( .A1(DATAO_REG_6__SCAN_IN), .A2(keyinput176), .B1(
        DATAO_REG_4__SCAN_IN), .B2(keyinput172), .ZN(n4663) );
  OAI221_X1 U5210 ( .B1(DATAO_REG_6__SCAN_IN), .B2(keyinput176), .C1(
        DATAO_REG_4__SCAN_IN), .C2(keyinput172), .A(n4663), .ZN(n4670) );
  AOI22_X1 U5211 ( .A1(DATAO_REG_11__SCAN_IN), .A2(keyinput213), .B1(
        DATAO_REG_5__SCAN_IN), .B2(keyinput245), .ZN(n4664) );
  OAI221_X1 U5212 ( .B1(DATAO_REG_11__SCAN_IN), .B2(keyinput213), .C1(
        DATAO_REG_5__SCAN_IN), .C2(keyinput245), .A(n4664), .ZN(n4669) );
  AOI22_X1 U5213 ( .A1(DATAO_REG_17__SCAN_IN), .A2(keyinput134), .B1(
        DATAO_REG_16__SCAN_IN), .B2(keyinput212), .ZN(n4665) );
  OAI221_X1 U5214 ( .B1(DATAO_REG_17__SCAN_IN), .B2(keyinput134), .C1(
        DATAO_REG_16__SCAN_IN), .C2(keyinput212), .A(n4665), .ZN(n4668) );
  AOI22_X1 U5215 ( .A1(DATAO_REG_27__SCAN_IN), .A2(keyinput231), .B1(
        REG3_REG_18__SCAN_IN), .B2(keyinput148), .ZN(n4666) );
  OAI221_X1 U5216 ( .B1(DATAO_REG_27__SCAN_IN), .B2(keyinput231), .C1(
        REG3_REG_18__SCAN_IN), .C2(keyinput148), .A(n4666), .ZN(n4667) );
  NOR4_X1 U5217 ( .A1(n4670), .A2(n4669), .A3(n4668), .A4(n4667), .ZN(n4684)
         );
  AOI22_X1 U5218 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput132), .B1(
        D_REG_8__SCAN_IN), .B2(keyinput175), .ZN(n4671) );
  OAI221_X1 U5219 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput132), .C1(
        D_REG_8__SCAN_IN), .C2(keyinput175), .A(n4671), .ZN(n4682) );
  AOI22_X1 U5220 ( .A1(n4673), .A2(keyinput237), .B1(keyinput200), .B2(n2669), 
        .ZN(n4672) );
  OAI221_X1 U5221 ( .B1(n4673), .B2(keyinput237), .C1(n2669), .C2(keyinput200), 
        .A(n4672), .ZN(n4681) );
  INV_X1 U5222 ( .A(DATAI_21_), .ZN(n4675) );
  AOI22_X1 U5223 ( .A1(n4675), .A2(keyinput140), .B1(keyinput155), .B2(n4884), 
        .ZN(n4674) );
  OAI221_X1 U5224 ( .B1(n4675), .B2(keyinput140), .C1(n4884), .C2(keyinput155), 
        .A(n4674), .ZN(n4680) );
  AOI22_X1 U5225 ( .A1(n4678), .A2(keyinput216), .B1(keyinput255), .B2(n4677), 
        .ZN(n4676) );
  OAI221_X1 U5226 ( .B1(n4678), .B2(keyinput216), .C1(n4677), .C2(keyinput255), 
        .A(n4676), .ZN(n4679) );
  NOR4_X1 U5227 ( .A1(n4682), .A2(n4681), .A3(n4680), .A4(n4679), .ZN(n4683)
         );
  NAND4_X1 U5228 ( .A1(n4686), .A2(n4685), .A3(n4684), .A4(n4683), .ZN(n4787)
         );
  AOI22_X1 U5229 ( .A1(n4867), .A2(keyinput174), .B1(n4688), .B2(keyinput221), 
        .ZN(n4687) );
  OAI221_X1 U5230 ( .B1(n4867), .B2(keyinput174), .C1(n4688), .C2(keyinput221), 
        .A(n4687), .ZN(n4696) );
  AOI22_X1 U5231 ( .A1(n4811), .A2(keyinput204), .B1(n4833), .B2(keyinput219), 
        .ZN(n4689) );
  OAI221_X1 U5232 ( .B1(n4811), .B2(keyinput204), .C1(n4833), .C2(keyinput219), 
        .A(n4689), .ZN(n4695) );
  XNOR2_X1 U5233 ( .A(DATAI_2_), .B(keyinput242), .ZN(n4693) );
  XNOR2_X1 U5234 ( .A(DATAI_1_), .B(keyinput236), .ZN(n4692) );
  XNOR2_X1 U5235 ( .A(IR_REG_3__SCAN_IN), .B(keyinput229), .ZN(n4691) );
  XNOR2_X1 U5236 ( .A(IR_REG_0__SCAN_IN), .B(keyinput184), .ZN(n4690) );
  NAND4_X1 U5237 ( .A1(n4693), .A2(n4692), .A3(n4691), .A4(n4690), .ZN(n4694)
         );
  NOR3_X1 U5238 ( .A1(n4696), .A2(n4695), .A3(n4694), .ZN(n4737) );
  AOI22_X1 U5239 ( .A1(n2446), .A2(keyinput182), .B1(keyinput246), .B2(n4698), 
        .ZN(n4697) );
  OAI221_X1 U5240 ( .B1(n2446), .B2(keyinput182), .C1(n4698), .C2(keyinput246), 
        .A(n4697), .ZN(n4706) );
  XNOR2_X1 U5241 ( .A(keyinput194), .B(n2444), .ZN(n4705) );
  XNOR2_X1 U5242 ( .A(keyinput240), .B(n2387), .ZN(n4704) );
  XNOR2_X1 U5243 ( .A(IR_REG_5__SCAN_IN), .B(keyinput214), .ZN(n4702) );
  XNOR2_X1 U5244 ( .A(IR_REG_4__SCAN_IN), .B(keyinput192), .ZN(n4701) );
  XNOR2_X1 U5245 ( .A(IR_REG_26__SCAN_IN), .B(keyinput226), .ZN(n4700) );
  XNOR2_X1 U5246 ( .A(IR_REG_13__SCAN_IN), .B(keyinput252), .ZN(n4699) );
  NAND4_X1 U5247 ( .A1(n4702), .A2(n4701), .A3(n4700), .A4(n4699), .ZN(n4703)
         );
  NOR4_X1 U5248 ( .A1(n4706), .A2(n4705), .A3(n4704), .A4(n4703), .ZN(n4736)
         );
  AOI22_X1 U5249 ( .A1(n4821), .A2(keyinput220), .B1(keyinput196), .B2(n4805), 
        .ZN(n4707) );
  OAI221_X1 U5250 ( .B1(n4821), .B2(keyinput220), .C1(n4805), .C2(keyinput196), 
        .A(n4707), .ZN(n4718) );
  AOI22_X1 U5251 ( .A1(n4709), .A2(keyinput207), .B1(keyinput218), .B2(n4835), 
        .ZN(n4708) );
  OAI221_X1 U5252 ( .B1(n4709), .B2(keyinput207), .C1(n4835), .C2(keyinput218), 
        .A(n4708), .ZN(n4717) );
  AOI22_X1 U5253 ( .A1(n4836), .A2(keyinput223), .B1(keyinput199), .B2(n4711), 
        .ZN(n4710) );
  OAI221_X1 U5254 ( .B1(n4836), .B2(keyinput223), .C1(n4711), .C2(keyinput199), 
        .A(n4710), .ZN(n4716) );
  AOI22_X1 U5255 ( .A1(n4714), .A2(keyinput193), .B1(n4713), .B2(keyinput138), 
        .ZN(n4712) );
  OAI221_X1 U5256 ( .B1(n4714), .B2(keyinput193), .C1(n4713), .C2(keyinput138), 
        .A(n4712), .ZN(n4715) );
  NOR4_X1 U5257 ( .A1(n4718), .A2(n4717), .A3(n4716), .A4(n4715), .ZN(n4735)
         );
  AOI22_X1 U5258 ( .A1(n4721), .A2(keyinput198), .B1(n4720), .B2(keyinput151), 
        .ZN(n4719) );
  OAI221_X1 U5259 ( .B1(n4721), .B2(keyinput198), .C1(n4720), .C2(keyinput151), 
        .A(n4719), .ZN(n4733) );
  INV_X1 U5260 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4724) );
  AOI22_X1 U5261 ( .A1(n4724), .A2(keyinput161), .B1(n4723), .B2(keyinput234), 
        .ZN(n4722) );
  OAI221_X1 U5262 ( .B1(n4724), .B2(keyinput161), .C1(n4723), .C2(keyinput234), 
        .A(n4722), .ZN(n4732) );
  AOI22_X1 U5263 ( .A1(n4727), .A2(keyinput211), .B1(keyinput144), .B2(n4726), 
        .ZN(n4725) );
  OAI221_X1 U5264 ( .B1(n4727), .B2(keyinput211), .C1(n4726), .C2(keyinput144), 
        .A(n4725), .ZN(n4731) );
  AOI22_X1 U5265 ( .A1(n4855), .A2(keyinput190), .B1(keyinput143), .B2(n4729), 
        .ZN(n4728) );
  OAI221_X1 U5266 ( .B1(n4855), .B2(keyinput190), .C1(n4729), .C2(keyinput143), 
        .A(n4728), .ZN(n4730) );
  NOR4_X1 U5267 ( .A1(n4733), .A2(n4732), .A3(n4731), .A4(n4730), .ZN(n4734)
         );
  NAND4_X1 U5268 ( .A1(n4737), .A2(n4736), .A3(n4735), .A4(n4734), .ZN(n4786)
         );
  INV_X1 U5269 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4739) );
  AOI22_X1 U5270 ( .A1(n4739), .A2(keyinput181), .B1(keyinput146), .B2(n4880), 
        .ZN(n4738) );
  OAI221_X1 U5271 ( .B1(n4739), .B2(keyinput181), .C1(n4880), .C2(keyinput146), 
        .A(n4738), .ZN(n4747) );
  AOI22_X1 U5272 ( .A1(n4857), .A2(keyinput210), .B1(keyinput248), .B2(n2896), 
        .ZN(n4740) );
  OAI221_X1 U5273 ( .B1(n4857), .B2(keyinput210), .C1(n2896), .C2(keyinput248), 
        .A(n4740), .ZN(n4746) );
  AOI22_X1 U5274 ( .A1(n4742), .A2(keyinput189), .B1(n2905), .B2(keyinput157), 
        .ZN(n4741) );
  OAI221_X1 U5275 ( .B1(n4742), .B2(keyinput189), .C1(n2905), .C2(keyinput157), 
        .A(n4741), .ZN(n4745) );
  AOI22_X1 U5276 ( .A1(n4869), .A2(keyinput167), .B1(n3318), .B2(keyinput141), 
        .ZN(n4743) );
  OAI221_X1 U5277 ( .B1(n4869), .B2(keyinput167), .C1(n3318), .C2(keyinput141), 
        .A(n4743), .ZN(n4744) );
  NOR4_X1 U5278 ( .A1(n4747), .A2(n4746), .A3(n4745), .A4(n4744), .ZN(n4784)
         );
  INV_X1 U5279 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4824) );
  AOI22_X1 U5280 ( .A1(n4824), .A2(keyinput251), .B1(keyinput180), .B2(n3331), 
        .ZN(n4748) );
  OAI221_X1 U5281 ( .B1(n4824), .B2(keyinput251), .C1(n3331), .C2(keyinput180), 
        .A(n4748), .ZN(n4758) );
  AOI22_X1 U5282 ( .A1(n4060), .A2(keyinput166), .B1(keyinput241), .B2(n4003), 
        .ZN(n4749) );
  OAI221_X1 U5283 ( .B1(n4060), .B2(keyinput166), .C1(n4003), .C2(keyinput241), 
        .A(n4749), .ZN(n4757) );
  INV_X1 U5284 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4790) );
  AOI22_X1 U5285 ( .A1(n4751), .A2(keyinput228), .B1(keyinput217), .B2(n4790), 
        .ZN(n4750) );
  OAI221_X1 U5286 ( .B1(n4751), .B2(keyinput228), .C1(n4790), .C2(keyinput217), 
        .A(n4750), .ZN(n4756) );
  AOI22_X1 U5287 ( .A1(n4754), .A2(keyinput173), .B1(keyinput152), .B2(n4753), 
        .ZN(n4752) );
  OAI221_X1 U5288 ( .B1(n4754), .B2(keyinput173), .C1(n4753), .C2(keyinput152), 
        .A(n4752), .ZN(n4755) );
  NOR4_X1 U5289 ( .A1(n4758), .A2(n4757), .A3(n4756), .A4(n4755), .ZN(n4783)
         );
  INV_X1 U5290 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n4802) );
  AOI22_X1 U5291 ( .A1(n4893), .A2(keyinput149), .B1(n4802), .B2(keyinput164), 
        .ZN(n4759) );
  OAI221_X1 U5292 ( .B1(n4893), .B2(keyinput149), .C1(n4802), .C2(keyinput164), 
        .A(n4759), .ZN(n4770) );
  INV_X1 U5293 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n4761) );
  AOI22_X1 U5294 ( .A1(n4761), .A2(keyinput225), .B1(keyinput185), .B2(n4899), 
        .ZN(n4760) );
  OAI221_X1 U5295 ( .B1(n4761), .B2(keyinput225), .C1(n4899), .C2(keyinput185), 
        .A(n4760), .ZN(n4769) );
  INV_X1 U5296 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n4763) );
  AOI22_X1 U5297 ( .A1(n4764), .A2(keyinput187), .B1(keyinput131), .B2(n4763), 
        .ZN(n4762) );
  OAI221_X1 U5298 ( .B1(n4764), .B2(keyinput187), .C1(n4763), .C2(keyinput131), 
        .A(n4762), .ZN(n4768) );
  AOI22_X1 U5299 ( .A1(n4766), .A2(keyinput179), .B1(keyinput136), .B2(n4803), 
        .ZN(n4765) );
  OAI221_X1 U5300 ( .B1(n4766), .B2(keyinput179), .C1(n4803), .C2(keyinput136), 
        .A(n4765), .ZN(n4767) );
  NOR4_X1 U5301 ( .A1(n4770), .A2(n4769), .A3(n4768), .A4(n4767), .ZN(n4782)
         );
  AOI22_X1 U5302 ( .A1(n4772), .A2(keyinput147), .B1(keyinput238), .B2(n4817), 
        .ZN(n4771) );
  OAI221_X1 U5303 ( .B1(n4772), .B2(keyinput147), .C1(n4817), .C2(keyinput238), 
        .A(n4771), .ZN(n4780) );
  INV_X1 U5304 ( .A(B_REG_SCAN_IN), .ZN(n4774) );
  AOI22_X1 U5305 ( .A1(n4823), .A2(keyinput244), .B1(n4774), .B2(keyinput129), 
        .ZN(n4773) );
  OAI221_X1 U5306 ( .B1(n4823), .B2(keyinput244), .C1(n4774), .C2(keyinput129), 
        .A(n4773), .ZN(n4779) );
  AOI22_X1 U5307 ( .A1(n4839), .A2(keyinput239), .B1(keyinput253), .B2(n2851), 
        .ZN(n4775) );
  OAI221_X1 U5308 ( .B1(n4839), .B2(keyinput239), .C1(n2851), .C2(keyinput253), 
        .A(n4775), .ZN(n4778) );
  INV_X1 U5309 ( .A(ADDR_REG_19__SCAN_IN), .ZN(n4818) );
  INV_X1 U5310 ( .A(IR_REG_29__SCAN_IN), .ZN(n4871) );
  AOI22_X1 U5311 ( .A1(n4818), .A2(keyinput247), .B1(n4871), .B2(keyinput162), 
        .ZN(n4776) );
  OAI221_X1 U5312 ( .B1(n4818), .B2(keyinput247), .C1(n4871), .C2(keyinput162), 
        .A(n4776), .ZN(n4777) );
  NOR4_X1 U5313 ( .A1(n4780), .A2(n4779), .A3(n4778), .A4(n4777), .ZN(n4781)
         );
  NAND4_X1 U5314 ( .A1(n4784), .A2(n4783), .A3(n4782), .A4(n4781), .ZN(n4785)
         );
  NOR4_X1 U5315 ( .A1(n4788), .A2(n4787), .A3(n4786), .A4(n4785), .ZN(n4987)
         );
  AOI22_X1 U5316 ( .A1(DATAO_REG_19__SCAN_IN), .A2(keyinput51), .B1(n4790), 
        .B2(keyinput89), .ZN(n4789) );
  OAI221_X1 U5317 ( .B1(DATAO_REG_19__SCAN_IN), .B2(keyinput51), .C1(n4790), 
        .C2(keyinput89), .A(n4789), .ZN(n4800) );
  AOI22_X1 U5318 ( .A1(DATAO_REG_23__SCAN_IN), .A2(keyinput19), .B1(
        DATAO_REG_2__SCAN_IN), .B2(keyinput59), .ZN(n4791) );
  OAI221_X1 U5319 ( .B1(DATAO_REG_23__SCAN_IN), .B2(keyinput19), .C1(
        DATAO_REG_2__SCAN_IN), .C2(keyinput59), .A(n4791), .ZN(n4796) );
  XNOR2_X1 U5320 ( .A(n4792), .B(keyinput117), .ZN(n4795) );
  XNOR2_X1 U5321 ( .A(n4793), .B(keyinput101), .ZN(n4794) );
  OR3_X1 U5322 ( .A1(n4796), .A2(n4795), .A3(n4794), .ZN(n4799) );
  AOI22_X1 U5323 ( .A1(DATAO_REG_14__SCAN_IN), .A2(keyinput3), .B1(
        REG0_REG_20__SCAN_IN), .B2(keyinput23), .ZN(n4797) );
  OAI221_X1 U5324 ( .B1(DATAO_REG_14__SCAN_IN), .B2(keyinput3), .C1(
        REG0_REG_20__SCAN_IN), .C2(keyinput23), .A(n4797), .ZN(n4798) );
  NOR3_X1 U5325 ( .A1(n4800), .A2(n4799), .A3(n4798), .ZN(n4850) );
  AOI22_X1 U5326 ( .A1(n4803), .A2(keyinput8), .B1(n4802), .B2(keyinput36), 
        .ZN(n4801) );
  OAI221_X1 U5327 ( .B1(n4803), .B2(keyinput8), .C1(n4802), .C2(keyinput36), 
        .A(n4801), .ZN(n4815) );
  AOI22_X1 U5328 ( .A1(n4806), .A2(keyinput28), .B1(n4805), .B2(keyinput68), 
        .ZN(n4804) );
  OAI221_X1 U5329 ( .B1(n4806), .B2(keyinput28), .C1(n4805), .C2(keyinput68), 
        .A(n4804), .ZN(n4814) );
  AOI22_X1 U5330 ( .A1(n4808), .A2(keyinput60), .B1(n2669), .B2(keyinput72), 
        .ZN(n4807) );
  OAI221_X1 U5331 ( .B1(n4808), .B2(keyinput60), .C1(n2669), .C2(keyinput72), 
        .A(n4807), .ZN(n4813) );
  AOI22_X1 U5332 ( .A1(n4811), .A2(keyinput76), .B1(keyinput104), .B2(n4810), 
        .ZN(n4809) );
  OAI221_X1 U5333 ( .B1(n4811), .B2(keyinput76), .C1(n4810), .C2(keyinput104), 
        .A(n4809), .ZN(n4812) );
  NOR4_X1 U5334 ( .A1(n4815), .A2(n4814), .A3(n4813), .A4(n4812), .ZN(n4849)
         );
  AOI22_X1 U5335 ( .A1(n4818), .A2(keyinput119), .B1(keyinput110), .B2(n4817), 
        .ZN(n4816) );
  OAI221_X1 U5336 ( .B1(n4818), .B2(keyinput119), .C1(n4817), .C2(keyinput110), 
        .A(n4816), .ZN(n4830) );
  AOI22_X1 U5337 ( .A1(n4821), .A2(keyinput92), .B1(keyinput96), .B2(n4820), 
        .ZN(n4819) );
  OAI221_X1 U5338 ( .B1(n4821), .B2(keyinput92), .C1(n4820), .C2(keyinput96), 
        .A(n4819), .ZN(n4829) );
  AOI22_X1 U5339 ( .A1(n4823), .A2(keyinput116), .B1(n2448), .B2(keyinput126), 
        .ZN(n4822) );
  OAI221_X1 U5340 ( .B1(n4823), .B2(keyinput116), .C1(n2448), .C2(keyinput126), 
        .A(n4822), .ZN(n4828) );
  XOR2_X1 U5341 ( .A(n4824), .B(keyinput123), .Z(n4826) );
  XNOR2_X1 U5342 ( .A(IR_REG_4__SCAN_IN), .B(keyinput64), .ZN(n4825) );
  NAND2_X1 U5343 ( .A1(n4826), .A2(n4825), .ZN(n4827) );
  NOR4_X1 U5344 ( .A1(n4830), .A2(n4829), .A3(n4828), .A4(n4827), .ZN(n4848)
         );
  AOI22_X1 U5345 ( .A1(n4833), .A2(keyinput91), .B1(keyinput87), .B2(n4832), 
        .ZN(n4831) );
  OAI221_X1 U5346 ( .B1(n4833), .B2(keyinput91), .C1(n4832), .C2(keyinput87), 
        .A(n4831), .ZN(n4846) );
  AOI22_X1 U5347 ( .A1(n4836), .A2(keyinput95), .B1(n4835), .B2(keyinput90), 
        .ZN(n4834) );
  OAI221_X1 U5348 ( .B1(n4836), .B2(keyinput95), .C1(n4835), .C2(keyinput90), 
        .A(n4834), .ZN(n4845) );
  INV_X1 U5349 ( .A(ADDR_REG_12__SCAN_IN), .ZN(n4838) );
  AOI22_X1 U5350 ( .A1(n4839), .A2(keyinput111), .B1(keyinput102), .B2(n4838), 
        .ZN(n4837) );
  OAI221_X1 U5351 ( .B1(n4839), .B2(keyinput111), .C1(n4838), .C2(keyinput102), 
        .A(n4837), .ZN(n4844) );
  XOR2_X1 U5352 ( .A(n4840), .B(keyinput94), .Z(n4842) );
  XNOR2_X1 U5353 ( .A(IR_REG_26__SCAN_IN), .B(keyinput98), .ZN(n4841) );
  NAND2_X1 U5354 ( .A1(n4842), .A2(n4841), .ZN(n4843) );
  NOR4_X1 U5355 ( .A1(n4846), .A2(n4845), .A3(n4844), .A4(n4843), .ZN(n4847)
         );
  NAND4_X1 U5356 ( .A1(n4850), .A2(n4849), .A3(n4848), .A4(n4847), .ZN(n4986)
         );
  AOI22_X1 U5357 ( .A1(n2446), .A2(keyinput54), .B1(keyinput55), .B2(n4852), 
        .ZN(n4851) );
  OAI221_X1 U5358 ( .B1(n2446), .B2(keyinput54), .C1(n4852), .C2(keyinput55), 
        .A(n4851), .ZN(n4864) );
  AOI22_X1 U5359 ( .A1(n4855), .A2(keyinput62), .B1(n4854), .B2(keyinput58), 
        .ZN(n4853) );
  OAI221_X1 U5360 ( .B1(n4855), .B2(keyinput62), .C1(n4854), .C2(keyinput58), 
        .A(n4853), .ZN(n4863) );
  AOI22_X1 U5361 ( .A1(n4858), .A2(keyinput78), .B1(keyinput82), .B2(n4857), 
        .ZN(n4856) );
  OAI221_X1 U5362 ( .B1(n4858), .B2(keyinput78), .C1(n4857), .C2(keyinput82), 
        .A(n4856), .ZN(n4862) );
  XNOR2_X1 U5363 ( .A(IR_REG_7__SCAN_IN), .B(keyinput63), .ZN(n4860) );
  XNOR2_X1 U5364 ( .A(REG3_REG_28__SCAN_IN), .B(keyinput75), .ZN(n4859) );
  NAND2_X1 U5365 ( .A1(n4860), .A2(n4859), .ZN(n4861) );
  NOR4_X1 U5366 ( .A1(n4864), .A2(n4863), .A3(n4862), .A4(n4861), .ZN(n4909)
         );
  AOI22_X1 U5367 ( .A1(n4867), .A2(keyinput46), .B1(n4866), .B2(keyinput42), 
        .ZN(n4865) );
  OAI221_X1 U5368 ( .B1(n4867), .B2(keyinput46), .C1(n4866), .C2(keyinput42), 
        .A(n4865), .ZN(n4878) );
  AOI22_X1 U5369 ( .A1(n2525), .A2(keyinput43), .B1(n4869), .B2(keyinput39), 
        .ZN(n4868) );
  OAI221_X1 U5370 ( .B1(n2525), .B2(keyinput43), .C1(n4869), .C2(keyinput39), 
        .A(n4868), .ZN(n4877) );
  AOI22_X1 U5371 ( .A1(n4871), .A2(keyinput34), .B1(keyinput35), .B2(n3172), 
        .ZN(n4870) );
  OAI221_X1 U5372 ( .B1(n4871), .B2(keyinput34), .C1(n3172), .C2(keyinput35), 
        .A(n4870), .ZN(n4876) );
  INV_X1 U5373 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4874) );
  AOI22_X1 U5374 ( .A1(n4874), .A2(keyinput30), .B1(n4873), .B2(keyinput31), 
        .ZN(n4872) );
  OAI221_X1 U5375 ( .B1(n4874), .B2(keyinput30), .C1(n4873), .C2(keyinput31), 
        .A(n4872), .ZN(n4875) );
  NOR4_X1 U5376 ( .A1(n4878), .A2(n4877), .A3(n4876), .A4(n4875), .ZN(n4908)
         );
  AOI22_X1 U5377 ( .A1(n4881), .A2(keyinput22), .B1(keyinput18), .B2(n4880), 
        .ZN(n4879) );
  OAI221_X1 U5378 ( .B1(n4881), .B2(keyinput22), .C1(n4880), .C2(keyinput18), 
        .A(n4879), .ZN(n4891) );
  AOI22_X1 U5379 ( .A1(n2879), .A2(keyinput7), .B1(n2539), .B2(keyinput2), 
        .ZN(n4882) );
  OAI221_X1 U5380 ( .B1(n2879), .B2(keyinput7), .C1(n2539), .C2(keyinput2), 
        .A(n4882), .ZN(n4890) );
  INV_X1 U5381 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4885) );
  AOI22_X1 U5382 ( .A1(n4885), .A2(keyinput26), .B1(keyinput27), .B2(n4884), 
        .ZN(n4883) );
  OAI221_X1 U5383 ( .B1(n4885), .B2(keyinput26), .C1(n4884), .C2(keyinput27), 
        .A(n4883), .ZN(n4889) );
  XNOR2_X1 U5384 ( .A(REG1_REG_18__SCAN_IN), .B(keyinput15), .ZN(n4887) );
  XNOR2_X1 U5385 ( .A(IR_REG_8__SCAN_IN), .B(keyinput11), .ZN(n4886) );
  NAND2_X1 U5386 ( .A1(n4887), .A2(n4886), .ZN(n4888) );
  NOR4_X1 U5387 ( .A1(n4891), .A2(n4890), .A3(n4889), .A4(n4888), .ZN(n4907)
         );
  INV_X1 U5388 ( .A(DATAI_3_), .ZN(n4894) );
  AOI22_X1 U5389 ( .A1(n4894), .A2(keyinput17), .B1(keyinput21), .B2(n4893), 
        .ZN(n4892) );
  OAI221_X1 U5390 ( .B1(n4894), .B2(keyinput17), .C1(n4893), .C2(keyinput21), 
        .A(n4892), .ZN(n4905) );
  AOI22_X1 U5391 ( .A1(n4897), .A2(keyinput41), .B1(keyinput25), .B2(n4896), 
        .ZN(n4895) );
  OAI221_X1 U5392 ( .B1(n4897), .B2(keyinput41), .C1(n4896), .C2(keyinput25), 
        .A(n4895), .ZN(n4904) );
  AOI22_X1 U5393 ( .A1(n3318), .A2(keyinput13), .B1(keyinput57), .B2(n4899), 
        .ZN(n4898) );
  OAI221_X1 U5394 ( .B1(n3318), .B2(keyinput13), .C1(n4899), .C2(keyinput57), 
        .A(n4898), .ZN(n4903) );
  XOR2_X1 U5395 ( .A(n2658), .B(keyinput69), .Z(n4901) );
  XNOR2_X1 U5396 ( .A(IR_REG_28__SCAN_IN), .B(keyinput9), .ZN(n4900) );
  NAND2_X1 U5397 ( .A1(n4901), .A2(n4900), .ZN(n4902) );
  NOR4_X1 U5398 ( .A1(n4905), .A2(n4904), .A3(n4903), .A4(n4902), .ZN(n4906)
         );
  NAND4_X1 U5399 ( .A1(n4909), .A2(n4908), .A3(n4907), .A4(n4906), .ZN(n4985)
         );
  OAI22_X1 U5400 ( .A1(REG3_REG_16__SCAN_IN), .A2(keyinput49), .B1(
        REG1_REG_31__SCAN_IN), .B2(keyinput61), .ZN(n4910) );
  AOI221_X1 U5401 ( .B1(REG3_REG_16__SCAN_IN), .B2(keyinput49), .C1(keyinput61), .C2(REG1_REG_31__SCAN_IN), .A(n4910), .ZN(n4917) );
  OAI22_X1 U5402 ( .A1(REG0_REG_22__SCAN_IN), .A2(keyinput33), .B1(keyinput53), 
        .B2(REG1_REG_21__SCAN_IN), .ZN(n4911) );
  AOI221_X1 U5403 ( .B1(REG0_REG_22__SCAN_IN), .B2(keyinput33), .C1(
        REG1_REG_21__SCAN_IN), .C2(keyinput53), .A(n4911), .ZN(n4916) );
  OAI22_X1 U5404 ( .A1(IR_REG_31__SCAN_IN), .A2(keyinput115), .B1(
        REG0_REG_0__SCAN_IN), .B2(keyinput99), .ZN(n4912) );
  AOI221_X1 U5405 ( .B1(IR_REG_31__SCAN_IN), .B2(keyinput115), .C1(keyinput99), 
        .C2(REG0_REG_0__SCAN_IN), .A(n4912), .ZN(n4915) );
  OAI22_X1 U5406 ( .A1(D_REG_2__SCAN_IN), .A2(keyinput0), .B1(keyinput45), 
        .B2(ADDR_REG_14__SCAN_IN), .ZN(n4913) );
  AOI221_X1 U5407 ( .B1(D_REG_2__SCAN_IN), .B2(keyinput0), .C1(
        ADDR_REG_14__SCAN_IN), .C2(keyinput45), .A(n4913), .ZN(n4914) );
  NAND4_X1 U5408 ( .A1(n4917), .A2(n4916), .A3(n4915), .A4(n4914), .ZN(n4945)
         );
  OAI22_X1 U5409 ( .A1(REG3_REG_13__SCAN_IN), .A2(keyinput93), .B1(
        ADDR_REG_0__SCAN_IN), .B2(keyinput97), .ZN(n4918) );
  AOI221_X1 U5410 ( .B1(REG3_REG_13__SCAN_IN), .B2(keyinput93), .C1(keyinput97), .C2(ADDR_REG_0__SCAN_IN), .A(n4918), .ZN(n4925) );
  OAI22_X1 U5411 ( .A1(REG3_REG_23__SCAN_IN), .A2(keyinput105), .B1(keyinput65), .B2(REG0_REG_10__SCAN_IN), .ZN(n4919) );
  AOI221_X1 U5412 ( .B1(REG3_REG_23__SCAN_IN), .B2(keyinput105), .C1(
        REG0_REG_10__SCAN_IN), .C2(keyinput65), .A(n4919), .ZN(n4924) );
  OAI22_X1 U5413 ( .A1(B_REG_SCAN_IN), .A2(keyinput1), .B1(
        ADDR_REG_17__SCAN_IN), .B2(keyinput5), .ZN(n4920) );
  AOI221_X1 U5414 ( .B1(B_REG_SCAN_IN), .B2(keyinput1), .C1(keyinput5), .C2(
        ADDR_REG_17__SCAN_IN), .A(n4920), .ZN(n4923) );
  OAI22_X1 U5415 ( .A1(IR_REG_25__SCAN_IN), .A2(keyinput81), .B1(
        STATE_REG_SCAN_IN), .B2(keyinput37), .ZN(n4921) );
  AOI221_X1 U5416 ( .B1(IR_REG_25__SCAN_IN), .B2(keyinput81), .C1(keyinput37), 
        .C2(STATE_REG_SCAN_IN), .A(n4921), .ZN(n4922) );
  NAND4_X1 U5417 ( .A1(n4925), .A2(n4924), .A3(n4923), .A4(n4922), .ZN(n4944)
         );
  OAI22_X1 U5418 ( .A1(IR_REG_17__SCAN_IN), .A2(keyinput112), .B1(keyinput108), 
        .B2(DATAI_1_), .ZN(n4926) );
  AOI221_X1 U5419 ( .B1(IR_REG_17__SCAN_IN), .B2(keyinput112), .C1(DATAI_1_), 
        .C2(keyinput108), .A(n4926), .ZN(n4933) );
  OAI22_X1 U5420 ( .A1(IR_REG_13__SCAN_IN), .A2(keyinput124), .B1(keyinput84), 
        .B2(DATAO_REG_16__SCAN_IN), .ZN(n4927) );
  AOI221_X1 U5421 ( .B1(IR_REG_13__SCAN_IN), .B2(keyinput124), .C1(
        DATAO_REG_16__SCAN_IN), .C2(keyinput84), .A(n4927), .ZN(n4932) );
  OAI22_X1 U5422 ( .A1(D_REG_8__SCAN_IN), .A2(keyinput47), .B1(
        REG0_REG_4__SCAN_IN), .B2(keyinput71), .ZN(n4928) );
  AOI221_X1 U5423 ( .B1(D_REG_8__SCAN_IN), .B2(keyinput47), .C1(keyinput71), 
        .C2(REG0_REG_4__SCAN_IN), .A(n4928), .ZN(n4931) );
  OAI22_X1 U5424 ( .A1(DATAI_14_), .A2(keyinput88), .B1(REG1_REG_0__SCAN_IN), 
        .B2(keyinput67), .ZN(n4929) );
  AOI221_X1 U5425 ( .B1(DATAI_14_), .B2(keyinput88), .C1(keyinput67), .C2(
        REG1_REG_0__SCAN_IN), .A(n4929), .ZN(n4930) );
  NAND4_X1 U5426 ( .A1(n4933), .A2(n4932), .A3(n4931), .A4(n4930), .ZN(n4943)
         );
  OAI22_X1 U5427 ( .A1(REG0_REG_25__SCAN_IN), .A2(keyinput83), .B1(
        DATAO_REG_27__SCAN_IN), .B2(keyinput103), .ZN(n4934) );
  AOI221_X1 U5428 ( .B1(REG0_REG_25__SCAN_IN), .B2(keyinput83), .C1(
        keyinput103), .C2(DATAO_REG_27__SCAN_IN), .A(n4934), .ZN(n4941) );
  OAI22_X1 U5429 ( .A1(D_REG_16__SCAN_IN), .A2(keyinput79), .B1(keyinput107), 
        .B2(REG0_REG_13__SCAN_IN), .ZN(n4935) );
  AOI221_X1 U5430 ( .B1(D_REG_16__SCAN_IN), .B2(keyinput79), .C1(
        REG0_REG_13__SCAN_IN), .C2(keyinput107), .A(n4935), .ZN(n4940) );
  OAI22_X1 U5431 ( .A1(D_REG_30__SCAN_IN), .A2(keyinput80), .B1(keyinput120), 
        .B2(REG2_REG_2__SCAN_IN), .ZN(n4936) );
  AOI221_X1 U5432 ( .B1(D_REG_30__SCAN_IN), .B2(keyinput80), .C1(
        REG2_REG_2__SCAN_IN), .C2(keyinput120), .A(n4936), .ZN(n4939) );
  OAI22_X1 U5433 ( .A1(DATAI_5_), .A2(keyinput127), .B1(REG2_REG_30__SCAN_IN), 
        .B2(keyinput100), .ZN(n4937) );
  AOI221_X1 U5434 ( .B1(DATAI_5_), .B2(keyinput127), .C1(keyinput100), .C2(
        REG2_REG_30__SCAN_IN), .A(n4937), .ZN(n4938) );
  NAND4_X1 U5435 ( .A1(n4941), .A2(n4940), .A3(n4939), .A4(n4938), .ZN(n4942)
         );
  NOR4_X1 U5436 ( .A1(n4945), .A2(n4944), .A3(n4943), .A4(n4942), .ZN(n4983)
         );
  OAI22_X1 U5437 ( .A1(REG2_REG_25__SCAN_IN), .A2(keyinput14), .B1(
        REG0_REG_12__SCAN_IN), .B2(keyinput10), .ZN(n4946) );
  AOI221_X1 U5438 ( .B1(REG2_REG_25__SCAN_IN), .B2(keyinput14), .C1(keyinput10), .C2(REG0_REG_12__SCAN_IN), .A(n4946), .ZN(n4953) );
  OAI22_X1 U5439 ( .A1(D_REG_15__SCAN_IN), .A2(keyinput50), .B1(
        REG2_REG_21__SCAN_IN), .B2(keyinput38), .ZN(n4947) );
  AOI221_X1 U5440 ( .B1(D_REG_15__SCAN_IN), .B2(keyinput50), .C1(keyinput38), 
        .C2(REG2_REG_21__SCAN_IN), .A(n4947), .ZN(n4952) );
  OAI22_X1 U5441 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput4), .B1(
        REG3_REG_2__SCAN_IN), .B2(keyinput125), .ZN(n4948) );
  AOI221_X1 U5442 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput4), .C1(keyinput125), .C2(REG3_REG_2__SCAN_IN), .A(n4948), .ZN(n4951) );
  OAI22_X1 U5443 ( .A1(REG2_REG_4__SCAN_IN), .A2(keyinput29), .B1(keyinput6), 
        .B2(DATAO_REG_17__SCAN_IN), .ZN(n4949) );
  AOI221_X1 U5444 ( .B1(REG2_REG_4__SCAN_IN), .B2(keyinput29), .C1(
        DATAO_REG_17__SCAN_IN), .C2(keyinput6), .A(n4949), .ZN(n4950) );
  NAND4_X1 U5445 ( .A1(n4953), .A2(n4952), .A3(n4951), .A4(n4950), .ZN(n4981)
         );
  OAI22_X1 U5446 ( .A1(IR_REG_16__SCAN_IN), .A2(keyinput118), .B1(
        REG1_REG_3__SCAN_IN), .B2(keyinput122), .ZN(n4954) );
  AOI221_X1 U5447 ( .B1(IR_REG_16__SCAN_IN), .B2(keyinput118), .C1(keyinput122), .C2(REG1_REG_3__SCAN_IN), .A(n4954), .ZN(n4961) );
  OAI22_X1 U5448 ( .A1(REG0_REG_23__SCAN_IN), .A2(keyinput106), .B1(
        keyinput114), .B2(DATAI_2_), .ZN(n4955) );
  AOI221_X1 U5449 ( .B1(REG0_REG_23__SCAN_IN), .B2(keyinput106), .C1(DATAI_2_), 
        .C2(keyinput114), .A(n4955), .ZN(n4960) );
  OAI22_X1 U5450 ( .A1(IR_REG_9__SCAN_IN), .A2(keyinput66), .B1(keyinput70), 
        .B2(REG0_REG_19__SCAN_IN), .ZN(n4956) );
  AOI221_X1 U5451 ( .B1(IR_REG_9__SCAN_IN), .B2(keyinput66), .C1(
        REG0_REG_19__SCAN_IN), .C2(keyinput70), .A(n4956), .ZN(n4959) );
  OAI22_X1 U5452 ( .A1(IR_REG_5__SCAN_IN), .A2(keyinput86), .B1(DATAI_28_), 
        .B2(keyinput74), .ZN(n4957) );
  AOI221_X1 U5453 ( .B1(IR_REG_5__SCAN_IN), .B2(keyinput86), .C1(keyinput74), 
        .C2(DATAI_28_), .A(n4957), .ZN(n4958) );
  NAND4_X1 U5454 ( .A1(n4961), .A2(n4960), .A3(n4959), .A4(n4958), .ZN(n4980)
         );
  OAI22_X1 U5455 ( .A1(IR_REG_6__SCAN_IN), .A2(keyinput32), .B1(keyinput40), 
        .B2(REG0_REG_5__SCAN_IN), .ZN(n4962) );
  AOI221_X1 U5456 ( .B1(IR_REG_6__SCAN_IN), .B2(keyinput32), .C1(
        REG0_REG_5__SCAN_IN), .C2(keyinput40), .A(n4962), .ZN(n4969) );
  OAI22_X1 U5457 ( .A1(REG2_REG_15__SCAN_IN), .A2(keyinput52), .B1(keyinput24), 
        .B2(ADDR_REG_7__SCAN_IN), .ZN(n4963) );
  AOI221_X1 U5458 ( .B1(REG2_REG_15__SCAN_IN), .B2(keyinput52), .C1(
        ADDR_REG_7__SCAN_IN), .C2(keyinput24), .A(n4963), .ZN(n4968) );
  OAI22_X1 U5459 ( .A1(D_REG_26__SCAN_IN), .A2(keyinput73), .B1(keyinput85), 
        .B2(DATAO_REG_11__SCAN_IN), .ZN(n4964) );
  AOI221_X1 U5460 ( .B1(D_REG_26__SCAN_IN), .B2(keyinput73), .C1(
        DATAO_REG_11__SCAN_IN), .C2(keyinput85), .A(n4964), .ZN(n4967) );
  OAI22_X1 U5461 ( .A1(REG0_REG_31__SCAN_IN), .A2(keyinput16), .B1(
        ADDR_REG_3__SCAN_IN), .B2(keyinput77), .ZN(n4965) );
  AOI221_X1 U5462 ( .B1(REG0_REG_31__SCAN_IN), .B2(keyinput16), .C1(keyinput77), .C2(ADDR_REG_3__SCAN_IN), .A(n4965), .ZN(n4966) );
  NAND4_X1 U5463 ( .A1(n4969), .A2(n4968), .A3(n4967), .A4(n4966), .ZN(n4979)
         );
  OAI22_X1 U5464 ( .A1(DATAI_21_), .A2(keyinput12), .B1(keyinput113), .B2(
        REG2_REG_24__SCAN_IN), .ZN(n4970) );
  AOI221_X1 U5465 ( .B1(DATAI_21_), .B2(keyinput12), .C1(REG2_REG_24__SCAN_IN), 
        .C2(keyinput113), .A(n4970), .ZN(n4977) );
  OAI22_X1 U5466 ( .A1(REG3_REG_18__SCAN_IN), .A2(keyinput20), .B1(
        REG0_REG_1__SCAN_IN), .B2(keyinput121), .ZN(n4971) );
  AOI221_X1 U5467 ( .B1(REG3_REG_18__SCAN_IN), .B2(keyinput20), .C1(
        keyinput121), .C2(REG0_REG_1__SCAN_IN), .A(n4971), .ZN(n4976) );
  OAI22_X1 U5468 ( .A1(IR_REG_0__SCAN_IN), .A2(keyinput56), .B1(keyinput48), 
        .B2(DATAO_REG_6__SCAN_IN), .ZN(n4972) );
  AOI221_X1 U5469 ( .B1(IR_REG_0__SCAN_IN), .B2(keyinput56), .C1(
        DATAO_REG_6__SCAN_IN), .C2(keyinput48), .A(n4972), .ZN(n4975) );
  OAI22_X1 U5470 ( .A1(DATAI_26_), .A2(keyinput109), .B1(DATAO_REG_4__SCAN_IN), 
        .B2(keyinput44), .ZN(n4973) );
  AOI221_X1 U5471 ( .B1(DATAI_26_), .B2(keyinput109), .C1(keyinput44), .C2(
        DATAO_REG_4__SCAN_IN), .A(n4973), .ZN(n4974) );
  NAND4_X1 U5472 ( .A1(n4977), .A2(n4976), .A3(n4975), .A4(n4974), .ZN(n4978)
         );
  NOR4_X1 U5473 ( .A1(n4981), .A2(n4980), .A3(n4979), .A4(n4978), .ZN(n4982)
         );
  NAND2_X1 U5474 ( .A1(n4983), .A2(n4982), .ZN(n4984) );
  NOR4_X1 U5475 ( .A1(n4987), .A2(n4986), .A3(n4985), .A4(n4984), .ZN(n4992)
         );
  NAND2_X1 U5476 ( .A1(n4989), .A2(U4043), .ZN(n4990) );
  OAI21_X1 U5477 ( .B1(U4043), .B2(DATAO_REG_14__SCAN_IN), .A(n4990), .ZN(
        n4991) );
  XNOR2_X1 U5478 ( .A(n4992), .B(n4991), .ZN(U3564) );
  NAND2_X1 U2518 ( .A1(n2750), .A2(n3659), .ZN(n3759) );
endmodule

