

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput0, keyinput1, keyinput2, 
        keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, 
        keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, 
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, 
        keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, 
        keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, 
        keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, 
        keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, 
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, 
        keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, 
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, 
        keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, 
        keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, 
        keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, 
        keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, 
        keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, 
        keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, 
        keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, 
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, 
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, 
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, 
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, 
        keyinput124, keyinput125, keyinput126, keyinput127 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084;

  INV_X1 U3548 ( .A(n6144), .ZN(n6237) );
  CLKBUF_X1 U3549 ( .A(n4660), .Z(n3104) );
  NAND2_X1 U3550 ( .A1(n5579), .A2(n5580), .ZN(n5568) );
  NAND2_X1 U3551 ( .A1(n4206), .A2(n4205), .ZN(n4207) );
  INV_X1 U3552 ( .A(n6518), .ZN(n3601) );
  NAND2_X1 U3553 ( .A1(n4308), .A2(n4462), .ZN(n4468) );
  CLKBUF_X2 U3554 ( .A(n3446), .Z(n4019) );
  INV_X2 U3555 ( .A(n4294), .ZN(n4348) );
  CLKBUF_X2 U3556 ( .A(n4039), .Z(n3118) );
  CLKBUF_X2 U3557 ( .A(n3463), .Z(n4057) );
  CLKBUF_X2 U3558 ( .A(n3294), .Z(n3115) );
  CLKBUF_X2 U3559 ( .A(n3509), .Z(n4054) );
  INV_X2 U3560 ( .A(n3362), .ZN(n4041) );
  CLKBUF_X2 U3561 ( .A(n3413), .Z(n4620) );
  INV_X1 U3562 ( .A(n3585), .ZN(n5374) );
  AND2_X2 U3563 ( .A1(n3277), .A2(n4788), .ZN(n3509) );
  CLKBUF_X1 U3564 ( .A(n6166), .Z(n3100) );
  NOR2_X1 U3565 ( .A1(n4526), .A2(n4505), .ZN(n6166) );
  AND4_X1 U3566 ( .A1(n3274), .A2(n3273), .A3(n3272), .A4(n3271), .ZN(n3283)
         );
  NAND2_X1 U3567 ( .A1(n3522), .A2(n3521), .ZN(n3525) );
  INV_X1 U3568 ( .A(n4537), .ZN(n4538) );
  AND4_X1 U3569 ( .A1(n3383), .A2(n3382), .A3(n3381), .A4(n3380), .ZN(n3389)
         );
  INV_X1 U3570 ( .A(n3659), .ZN(n4080) );
  OR2_X1 U3571 ( .A1(n5963), .A2(n4419), .ZN(n5944) );
  NAND2_X1 U3573 ( .A1(n3740), .A2(n3739), .ZN(n3752) );
  NAND2_X1 U3574 ( .A1(n5735), .A2(n5916), .ZN(n3144) );
  OR2_X1 U3575 ( .A1(n5965), .A2(n5897), .ZN(n5953) );
  CLKBUF_X3 U3576 ( .A(n6076), .Z(n3106) );
  INV_X1 U3577 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6603) );
  BUF_X1 U3578 ( .A(n4167), .Z(n5029) );
  XNOR2_X1 U3579 ( .A(n3262), .B(n4082), .ZN(n5376) );
  INV_X1 U3580 ( .A(n6175), .ZN(n6258) );
  OR2_X1 U3581 ( .A1(n3137), .A2(n4427), .ZN(n5692) );
  INV_X1 U3582 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3269) );
  NAND2_X2 U3583 ( .A1(n3389), .A2(n3388), .ZN(n3413) );
  AND4_X4 U3584 ( .A1(n3339), .A2(n3338), .A3(n3337), .A4(n3336), .ZN(n3445)
         );
  AND4_X2 U3585 ( .A1(n3331), .A2(n3330), .A3(n3329), .A4(n3328), .ZN(n3337)
         );
  AND4_X2 U3586 ( .A1(n3335), .A2(n3334), .A3(n3333), .A4(n3332), .ZN(n3336)
         );
  NOR2_X1 U3587 ( .A1(n3431), .A2(n4381), .ZN(n4140) );
  AND2_X4 U3588 ( .A1(n3306), .A2(n3305), .ZN(n3410) );
  XNOR2_X2 U3589 ( .A(n4207), .B(n6401), .ZN(n6337) );
  AND2_X1 U3590 ( .A1(n3278), .A2(n3326), .ZN(n3101) );
  AND2_X1 U3591 ( .A1(n3278), .A2(n3326), .ZN(n3117) );
  INV_X1 U3592 ( .A(n6337), .ZN(n3164) );
  INV_X1 U3593 ( .A(n3610), .ZN(n3526) );
  NAND2_X1 U3594 ( .A1(n6266), .A2(n5374), .ZN(n5672) );
  NAND2_X1 U3595 ( .A1(n4348), .A2(n4462), .ZN(n4499) );
  INV_X4 U3596 ( .A(n4364), .ZN(n4462) );
  INV_X2 U3598 ( .A(n3412), .ZN(n3102) );
  INV_X2 U3599 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3268) );
  AOI21_X1 U3600 ( .B1(n5916), .B2(n5742), .A(n5741), .ZN(n5931) );
  XNOR2_X1 U3601 ( .A(n4438), .B(n4437), .ZN(n4484) );
  AOI21_X1 U3602 ( .B1(n5802), .B2(n5801), .A(n3212), .ZN(n5794) );
  NAND2_X1 U3603 ( .A1(n3207), .A2(n3205), .ZN(n5786) );
  AOI21_X1 U3604 ( .B1(n5747), .B2(n6349), .A(n5746), .ZN(n5748) );
  AOI21_X1 U3605 ( .B1(n5376), .B2(n6349), .A(n4149), .ZN(n3236) );
  AND2_X1 U3606 ( .A1(n4452), .A2(n4451), .ZN(n5733) );
  AOI21_X1 U3607 ( .B1(n5429), .B2(n5440), .A(n5428), .ZN(n5765) );
  OAI21_X1 U3608 ( .B1(n5692), .B2(n5888), .A(n4430), .ZN(n4431) );
  OR2_X1 U3609 ( .A1(n5402), .A2(n5403), .ZN(n5404) );
  NAND2_X1 U3610 ( .A1(n3214), .A2(n3134), .ZN(n5783) );
  XNOR2_X1 U3611 ( .A(n4534), .B(n4533), .ZN(n5726) );
  AND2_X1 U3612 ( .A1(n3988), .A2(n3178), .ZN(n4534) );
  NAND2_X1 U3613 ( .A1(n3148), .A2(n3215), .ZN(n3147) );
  NAND2_X1 U3614 ( .A1(n3240), .A2(n3238), .ZN(n4236) );
  CLKBUF_X1 U3615 ( .A(n5427), .Z(n5440) );
  INV_X1 U3616 ( .A(n5381), .ZN(n5911) );
  AOI21_X1 U3617 ( .B1(n3239), .B2(n3215), .A(n3150), .ZN(n3149) );
  INV_X1 U3618 ( .A(n3204), .ZN(n3203) );
  AND2_X1 U3619 ( .A1(n3136), .A2(n4235), .ZN(n3215) );
  INV_X1 U3620 ( .A(n4240), .ZN(n3245) );
  OR2_X1 U3621 ( .A1(n3740), .A2(n3739), .ZN(n3157) );
  OR2_X1 U3622 ( .A1(n5848), .A2(n4239), .ZN(n4240) );
  AND2_X1 U3623 ( .A1(n5503), .A2(REIP_REG_20__SCAN_IN), .ZN(n5478) );
  AND2_X1 U3624 ( .A1(n4173), .A2(n4172), .ZN(n4864) );
  NAND2_X1 U3625 ( .A1(n3155), .A2(n3652), .ZN(n4868) );
  INV_X1 U3626 ( .A(n5483), .ZN(n3222) );
  NAND2_X1 U3627 ( .A1(n3645), .A2(n3644), .ZN(n4825) );
  AND2_X1 U3628 ( .A1(n6452), .A2(n5028), .ZN(n6593) );
  NOR2_X2 U3629 ( .A1(n4940), .A2(n5218), .ZN(n7076) );
  NAND2_X1 U3630 ( .A1(n6063), .A2(n6045), .ZN(n6079) );
  NAND2_X1 U3631 ( .A1(n4369), .A2(n4368), .ZN(n5483) );
  NAND2_X1 U3632 ( .A1(n3612), .A2(n3801), .ZN(n4827) );
  OR2_X1 U3633 ( .A1(n6392), .A2(n4817), .ZN(n5983) );
  OR2_X1 U3634 ( .A1(n5628), .A2(n4508), .ZN(n6144) );
  AND2_X2 U3635 ( .A1(n3526), .A2(n3611), .ZN(n3602) );
  AND2_X1 U3636 ( .A1(n6044), .A2(n4405), .ZN(n6392) );
  NAND2_X1 U3637 ( .A1(n6184), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5628) );
  NAND2_X2 U3638 ( .A1(n6741), .A2(n4503), .ZN(n6184) );
  CLKBUF_X1 U3639 ( .A(n4887), .Z(n4888) );
  NAND2_X1 U3640 ( .A1(n4278), .A2(n4277), .ZN(n4404) );
  OAI21_X1 U3641 ( .B1(n4157), .B2(n4219), .A(n4161), .ZN(n4691) );
  NAND2_X1 U3642 ( .A1(n3633), .A2(n3632), .ZN(n4157) );
  NAND2_X1 U3643 ( .A1(n3193), .A2(n3528), .ZN(n4630) );
  AOI21_X1 U3644 ( .B1(n3235), .B2(n3631), .A(n4218), .ZN(n3620) );
  AND2_X1 U3645 ( .A1(n4855), .A2(n4885), .ZN(n4884) );
  NOR2_X1 U3646 ( .A1(n4661), .A2(n4390), .ZN(n4394) );
  AND2_X1 U3647 ( .A1(n4314), .A2(n4313), .ZN(n4885) );
  NAND3_X1 U3648 ( .A1(n3419), .A2(n3434), .A3(n4140), .ZN(n3438) );
  INV_X1 U3649 ( .A(n3492), .ZN(n3630) );
  MUX2_X1 U3650 ( .A(n3491), .B(n4218), .S(n3490), .Z(n3492) );
  INV_X1 U3651 ( .A(n3402), .ZN(n4839) );
  NOR2_X1 U3652 ( .A1(n4381), .A2(n4089), .ZN(n3351) );
  OR2_X1 U3653 ( .A1(n3534), .A2(n4222), .ZN(n3479) );
  NAND2_X1 U3654 ( .A1(n3533), .A2(n3534), .ZN(n4127) );
  NAND2_X1 U3655 ( .A1(n4158), .A2(n3413), .ZN(n4336) );
  OR2_X1 U3656 ( .A1(n3119), .A2(n4872), .ZN(n3533) );
  AND3_X2 U3657 ( .A1(n3397), .A2(STATE2_REG_0__SCAN_IN), .A3(n3102), .ZN(
        n3461) );
  OR2_X1 U3658 ( .A1(n3489), .A2(n3488), .ZN(n4159) );
  OR2_X1 U3659 ( .A1(n3474), .A2(n3473), .ZN(n4222) );
  INV_X2 U3660 ( .A(n3412), .ZN(n4287) );
  INV_X2 U3661 ( .A(n3445), .ZN(n3397) );
  OR2_X2 U3662 ( .A1(n3350), .A2(n3349), .ZN(n3585) );
  AND4_X2 U3663 ( .A1(n3375), .A2(n3374), .A3(n3373), .A4(n3372), .ZN(n3412)
         );
  AND4_X1 U3664 ( .A1(n3387), .A2(n3386), .A3(n3385), .A4(n3384), .ZN(n3388)
         );
  AND4_X1 U3665 ( .A1(n3355), .A2(n3354), .A3(n3353), .A4(n3352), .ZN(n3375)
         );
  AND4_X1 U3666 ( .A1(n3298), .A2(n3297), .A3(n3296), .A4(n3295), .ZN(n3306)
         );
  AND2_X1 U3667 ( .A1(n3300), .A2(n3299), .ZN(n3304) );
  AND4_X1 U3668 ( .A1(n3321), .A2(n3320), .A3(n3319), .A4(n3318), .ZN(n3339)
         );
  AND4_X1 U3669 ( .A1(n3325), .A2(n3324), .A3(n3323), .A4(n3322), .ZN(n3338)
         );
  AND4_X1 U3670 ( .A1(n3366), .A2(n3365), .A3(n3364), .A4(n3363), .ZN(n3373)
         );
  AND4_X1 U3671 ( .A1(n3359), .A2(n3358), .A3(n3357), .A4(n3356), .ZN(n3374)
         );
  AND4_X1 U3672 ( .A1(n3371), .A2(n3370), .A3(n3369), .A4(n3368), .ZN(n3372)
         );
  OR2_X1 U3673 ( .A1(n4750), .A2(n3367), .ZN(n3368) );
  AOI21_X1 U3674 ( .B1(n3360), .B2(INSTQUEUE_REG_8__1__SCAN_IN), .A(n3377), 
        .ZN(n3383) );
  BUF_X2 U3675 ( .A(n3991), .Z(n4032) );
  BUF_X2 U3676 ( .A(n4033), .Z(n4053) );
  BUF_X2 U3677 ( .A(n4055), .Z(n4014) );
  BUF_X2 U3678 ( .A(n3462), .Z(n4058) );
  NAND2_X2 U3679 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6752), .ZN(n4576) );
  BUF_X2 U3680 ( .A(n3360), .Z(n4056) );
  BUF_X2 U3681 ( .A(n3378), .Z(n3907) );
  AND2_X1 U3682 ( .A1(n4040), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3377) );
  AND2_X2 U3683 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4677) );
  INV_X2 U3684 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3246) );
  NOR2_X2 U3685 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4744) );
  CLKBUF_X1 U3686 ( .A(n5205), .Z(n3103) );
  NAND2_X2 U3687 ( .A1(n3316), .A2(n3315), .ZN(n3396) );
  AND4_X1 U3688 ( .A1(n3314), .A2(n3313), .A3(n3312), .A4(n3311), .ZN(n3315)
         );
  OR2_X1 U3689 ( .A1(n3362), .A2(n3317), .ZN(n3319) );
  AND2_X2 U3690 ( .A1(n4788), .A2(n4744), .ZN(n3294) );
  NAND2_X1 U3691 ( .A1(n3445), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3534) );
  OAI211_X1 U3692 ( .C1(n3442), .C2(n3441), .A(n3440), .B(n3439), .ZN(n3478)
         );
  XNOR2_X1 U3693 ( .A(n3527), .B(n3528), .ZN(n4660) );
  OR2_X2 U3694 ( .A1(n3409), .A2(n4336), .ZN(n3426) );
  NAND2_X2 U3695 ( .A1(n3396), .A2(n3410), .ZN(n4453) );
  INV_X2 U3696 ( .A(n3396), .ZN(n3634) );
  NAND2_X2 U3697 ( .A1(n3460), .A2(n3459), .ZN(n3622) );
  AOI21_X2 U3698 ( .B1(n5029), .B2(n4209), .A(n4170), .ZN(n6356) );
  NOR2_X2 U3699 ( .A1(n4881), .A2(n4856), .ZN(n4855) );
  BUF_X4 U3701 ( .A(n6076), .Z(n3107) );
  INV_X2 U3702 ( .A(n4229), .ZN(n6076) );
  NAND2_X2 U3703 ( .A1(n3151), .A2(n3241), .ZN(n5736) );
  AND2_X1 U3704 ( .A1(n3326), .A2(n4745), .ZN(n3108) );
  AND2_X4 U3706 ( .A1(n3246), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3277)
         );
  AND2_X4 U3707 ( .A1(n4744), .A2(n3326), .ZN(n4039) );
  AND2_X1 U3708 ( .A1(n3277), .A2(n3276), .ZN(n3109) );
  INV_X1 U3709 ( .A(n3413), .ZN(n3110) );
  INV_X1 U3710 ( .A(n3413), .ZN(n3111) );
  AOI21_X2 U3711 ( .B1(n6344), .B2(n3153), .A(n3135), .ZN(n3152) );
  XNOR2_X2 U3712 ( .A(n4189), .B(n6420), .ZN(n6344) );
  AND2_X1 U3713 ( .A1(n3326), .A2(n4745), .ZN(n3112) );
  AND2_X1 U3714 ( .A1(n3326), .A2(n4745), .ZN(n3113) );
  AND2_X1 U3715 ( .A1(n3326), .A2(n4745), .ZN(n3116) );
  NAND2_X2 U3716 ( .A1(n4851), .A2(n4868), .ZN(n5024) );
  AND4_X2 U3717 ( .A1(n3646), .A2(n4825), .A3(n4852), .A4(n4853), .ZN(n4851)
         );
  XNOR2_X2 U3718 ( .A(n4181), .B(n6430), .ZN(n4863) );
  NAND2_X2 U3719 ( .A1(n4180), .A2(n4179), .ZN(n4181) );
  NOR2_X4 U3720 ( .A1(n5024), .A2(n5025), .ZN(n5068) );
  NAND2_X2 U3721 ( .A1(n6163), .A2(n5608), .ZN(n5144) );
  NOR3_X4 U3722 ( .A1(n5022), .A2(n5136), .A3(n3227), .ZN(n6163) );
  NAND2_X2 U3723 ( .A1(n4258), .A2(n3404), .ZN(n4283) );
  NOR2_X2 U3724 ( .A1(n4439), .A2(n3258), .ZN(n4425) );
  AOI21_X2 U3725 ( .B1(n3200), .B2(n3203), .A(n3198), .ZN(n3197) );
  OAI21_X2 U3726 ( .B1(n4865), .B2(n3154), .A(n3152), .ZN(n5093) );
  NAND2_X2 U3727 ( .A1(n4864), .A2(n4863), .ZN(n4865) );
  AOI22_X2 U3728 ( .A1(n5792), .A2(n4252), .B1(n5794), .B2(n4251), .ZN(n4253)
         );
  NOR2_X4 U3729 ( .A1(n5760), .A2(n5758), .ZN(n5735) );
  NAND2_X2 U3730 ( .A1(n5736), .A2(n4245), .ZN(n5760) );
  AOI21_X2 U3731 ( .B1(n5769), .B2(n5808), .A(n3120), .ZN(n5802) );
  NAND2_X2 U3732 ( .A1(n5783), .A2(n4240), .ZN(n5769) );
  NOR2_X2 U3733 ( .A1(n5568), .A2(n3216), .ZN(n5493) );
  XNOR2_X2 U3734 ( .A(n3525), .B(n3524), .ZN(n3611) );
  XNOR2_X1 U3735 ( .A(n3478), .B(n3477), .ZN(n3636) );
  XNOR2_X1 U3736 ( .A(n4301), .B(n4692), .ZN(n4819) );
  NAND2_X1 U3737 ( .A1(n3503), .A2(n3502), .ZN(n3527) );
  INV_X1 U3738 ( .A(n3412), .ZN(n3119) );
  NAND2_X1 U3739 ( .A1(n3403), .A2(n3634), .ZN(n3423) );
  AOI21_X1 U3740 ( .B1(n3423), .B2(n4158), .A(n5374), .ZN(n3401) );
  NAND2_X1 U3741 ( .A1(n4772), .A2(n6717), .ZN(n4711) );
  AND2_X2 U3742 ( .A1(n3268), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3276)
         );
  AND2_X1 U3743 ( .A1(n3942), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3943)
         );
  AND2_X1 U3744 ( .A1(n3243), .A2(n3149), .ZN(n3146) );
  INV_X1 U3745 ( .A(n3240), .ZN(n3148) );
  NOR2_X2 U3746 ( .A1(n4232), .A2(n3196), .ZN(n3204) );
  INV_X1 U3747 ( .A(n4227), .ZN(n3196) );
  AND4_X1 U3748 ( .A1(n3430), .A2(n3426), .A3(n3429), .A4(n4749), .ZN(n3436)
         );
  AND2_X1 U3749 ( .A1(n3390), .A2(n4274), .ZN(n3391) );
  OR2_X1 U3750 ( .A1(n4279), .A2(n3409), .ZN(n4780) );
  NAND2_X1 U3751 ( .A1(n4236), .A2(n3215), .ZN(n3214) );
  CLKBUF_X1 U3752 ( .A(n4742), .Z(n4743) );
  INV_X1 U3753 ( .A(n4157), .ZN(n5218) );
  NOR2_X1 U3754 ( .A1(n4135), .A2(n4267), .ZN(n4136) );
  INV_X1 U3755 ( .A(n4028), .ZN(n4502) );
  INV_X1 U3756 ( .A(n4605), .ZN(n4610) );
  NAND2_X1 U3757 ( .A1(n3558), .A2(n3557), .ZN(n3591) );
  INV_X1 U3758 ( .A(n3248), .ZN(n3181) );
  BUF_X1 U3759 ( .A(n4040), .Z(n3973) );
  AOI22_X1 U3760 ( .A1(n3996), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3379), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3291) );
  NAND2_X1 U3761 ( .A1(n3259), .A2(n3266), .ZN(n3258) );
  INV_X1 U3762 ( .A(n5460), .ZN(n3259) );
  NAND2_X1 U3763 ( .A1(n3251), .A2(n5582), .ZN(n3250) );
  INV_X1 U3764 ( .A(n5566), .ZN(n3251) );
  NOR2_X1 U3765 ( .A1(n7047), .A2(n3184), .ZN(n3183) );
  INV_X1 U3766 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3184) );
  NOR2_X2 U3767 ( .A1(n3396), .A2(n6603), .ZN(n3778) );
  INV_X1 U3768 ( .A(n5432), .ZN(n3231) );
  NOR2_X1 U3769 ( .A1(n5482), .A2(n3224), .ZN(n3223) );
  INV_X1 U3770 ( .A(n4486), .ZN(n3224) );
  INV_X1 U3771 ( .A(n5801), .ZN(n3211) );
  INV_X1 U3772 ( .A(n3209), .ZN(n3208) );
  OAI21_X1 U3773 ( .B1(n5808), .B2(n3120), .A(n3213), .ZN(n3209) );
  NAND2_X1 U3774 ( .A1(n3208), .A2(n3120), .ZN(n3206) );
  NAND2_X1 U3775 ( .A1(n4347), .A2(n3218), .ZN(n3217) );
  INV_X1 U3776 ( .A(n5552), .ZN(n3218) );
  INV_X1 U3777 ( .A(n4237), .ZN(n3150) );
  INV_X1 U3778 ( .A(n5890), .ZN(n3202) );
  OR2_X1 U3779 ( .A1(n3226), .A2(n4340), .ZN(n3225) );
  OR2_X1 U3780 ( .A1(n5147), .A2(n5364), .ZN(n3226) );
  NAND2_X1 U3781 ( .A1(n4884), .A2(n5023), .ZN(n5022) );
  NAND2_X1 U3782 ( .A1(n4925), .A2(n4158), .ZN(n4168) );
  NAND2_X1 U3783 ( .A1(n3476), .A2(n3478), .ZN(n3501) );
  AND2_X1 U3784 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4976) );
  NAND2_X1 U3785 ( .A1(n6603), .A2(n6129), .ZN(n4028) );
  CLKBUF_X1 U3786 ( .A(n4272), .Z(n4273) );
  INV_X1 U3787 ( .A(n4151), .ZN(n6746) );
  AND2_X1 U3788 ( .A1(n4460), .A2(n4459), .ZN(n5442) );
  INV_X1 U3789 ( .A(n4767), .ZN(n4713) );
  INV_X1 U3790 ( .A(n3801), .ZN(n4079) );
  AND2_X1 U3791 ( .A1(n3260), .A2(n3179), .ZN(n3178) );
  NAND2_X1 U3792 ( .A1(n4009), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4076)
         );
  NAND2_X1 U3793 ( .A1(n3869), .A2(n3128), .ZN(n3941) );
  NAND2_X1 U3794 ( .A1(n3781), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3818)
         );
  NAND2_X1 U3795 ( .A1(n3705), .A2(n3182), .ZN(n3764) );
  AND2_X1 U3796 ( .A1(n3126), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3182)
         );
  INV_X1 U3797 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n7047) );
  NOR2_X1 U3798 ( .A1(n3690), .A2(n6159), .ZN(n3705) );
  NAND3_X1 U3799 ( .A1(n3649), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .A3(n3125), 
        .ZN(n3690) );
  INV_X1 U3800 ( .A(n4198), .ZN(n3234) );
  INV_X1 U3801 ( .A(n4827), .ZN(n3645) );
  AND2_X1 U3802 ( .A1(n4830), .A2(n4829), .ZN(n4859) );
  AND2_X1 U3803 ( .A1(n4473), .A2(n4472), .ZN(n5407) );
  NOR2_X1 U3804 ( .A1(n4367), .A2(n5510), .ZN(n4368) );
  INV_X1 U3805 ( .A(n5509), .ZN(n4369) );
  AND2_X1 U3806 ( .A1(n4355), .A2(n4354), .ZN(n5538) );
  NAND2_X1 U3807 ( .A1(n3200), .A2(n5891), .ZN(n3199) );
  INV_X1 U3808 ( .A(n5857), .ZN(n3198) );
  INV_X1 U3809 ( .A(n4182), .ZN(n3153) );
  NAND2_X1 U3810 ( .A1(n5093), .A2(n5092), .ZN(n5091) );
  XNOR2_X1 U3811 ( .A(n3623), .B(n3622), .ZN(n4887) );
  XNOR2_X1 U3812 ( .A(n3620), .B(n3496), .ZN(n3623) );
  AND2_X1 U3813 ( .A1(n6449), .A2(n5212), .ZN(n5032) );
  AND2_X1 U3814 ( .A1(n5032), .A2(n5218), .ZN(n5097) );
  OR2_X1 U3815 ( .A1(n3104), .A2(n4786), .ZN(n6560) );
  NAND2_X1 U3816 ( .A1(n4900), .A2(n4872), .ZN(n5100) );
  INV_X1 U3817 ( .A(n4888), .ZN(n5212) );
  AND2_X1 U3818 ( .A1(n4891), .A2(n4931), .ZN(n4894) );
  AND2_X1 U3819 ( .A1(n4976), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5255)
         );
  AOI21_X1 U3820 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6651), .A(n5100), .ZN(
        n6523) );
  AOI21_X1 U3821 ( .B1(n6175), .B2(n5751), .A(n3194), .ZN(n5420) );
  AND2_X1 U3822 ( .A1(n6241), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3194)
         );
  INV_X1 U3823 ( .A(n6210), .ZN(n6249) );
  AND3_X1 U3824 ( .A1(n6423), .A2(n6720), .A3(n4971), .ZN(n4503) );
  INV_X1 U3825 ( .A(n5733), .ZN(n5679) );
  NAND2_X1 U3826 ( .A1(n4843), .A2(n6717), .ZN(n4844) );
  XNOR2_X1 U3827 ( .A(n4146), .B(n4145), .ZN(n5389) );
  NAND2_X1 U3828 ( .A1(n4009), .A2(n3185), .ZN(n4144) );
  INV_X1 U3829 ( .A(n5789), .ZN(n3160) );
  NAND2_X1 U3830 ( .A1(n6334), .A2(n4141), .ZN(n5884) );
  INV_X1 U3831 ( .A(n5884), .ZN(n6354) );
  OR2_X1 U3832 ( .A1(n4711), .A2(n4780), .ZN(n6334) );
  XNOR2_X1 U3833 ( .A(n3237), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5895)
         );
  OAI21_X1 U3834 ( .B1(n5786), .B2(n5785), .A(n5784), .ZN(n5787) );
  NAND2_X1 U3835 ( .A1(n5786), .A2(n4435), .ZN(n4438) );
  INV_X1 U3836 ( .A(n6423), .ZN(n6433) );
  NAND2_X1 U3837 ( .A1(n3629), .A2(n3630), .ZN(n3633) );
  INV_X1 U3838 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6651) );
  INV_X1 U3839 ( .A(n6655), .ZN(n6594) );
  INV_X1 U3840 ( .A(n5029), .ZN(n6452) );
  OR2_X1 U3841 ( .A1(n6655), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6109) );
  NAND2_X1 U3842 ( .A1(n5255), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4931) );
  AND2_X1 U3843 ( .A1(n4138), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6717) );
  AOI22_X1 U3844 ( .A1(n3446), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3465) );
  NAND2_X1 U3845 ( .A1(n3110), .A2(n4261), .ZN(n3411) );
  INV_X1 U3846 ( .A(n3533), .ZN(n3523) );
  OR2_X1 U3847 ( .A1(n3938), .A2(n3937), .ZN(n3949) );
  AND2_X1 U3848 ( .A1(n6518), .A2(n3591), .ZN(n3252) );
  OR2_X1 U3849 ( .A1(n3581), .A2(n3580), .ZN(n4211) );
  OR2_X1 U3850 ( .A1(n3568), .A2(n3567), .ZN(n4202) );
  AND2_X1 U3851 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        STATE2_REG_0__SCAN_IN), .ZN(n3437) );
  OAI21_X1 U3852 ( .B1(n3788), .B2(n3424), .A(n3267), .ZN(n3425) );
  NAND2_X1 U3853 ( .A1(n3420), .A2(n4839), .ZN(n3442) );
  OR2_X1 U3854 ( .A1(n3458), .A2(n3457), .ZN(n4150) );
  INV_X1 U3855 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U3856 ( .A1(n3446), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3378), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3382) );
  AOI21_X1 U3857 ( .B1(n3378), .B2(INSTQUEUE_REG_12__2__SCAN_IN), .A(n3270), 
        .ZN(n3273) );
  AND2_X1 U3858 ( .A1(n3109), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3270) );
  AOI22_X1 U3859 ( .A1(n3447), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3311) );
  AOI22_X1 U3860 ( .A1(n3996), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3379), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U3861 ( .A1(n3360), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3310) );
  OR2_X1 U3862 ( .A1(n4124), .A2(n4125), .ZN(n4130) );
  AOI21_X1 U3863 ( .B1(n3378), .B2(INSTQUEUE_REG_12__7__SCAN_IN), .A(n3340), 
        .ZN(n3344) );
  AND2_X1 U3864 ( .A1(n3446), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3340) );
  XNOR2_X1 U3865 ( .A(n3174), .B(n3591), .ZN(n4183) );
  NOR2_X1 U3866 ( .A1(n4450), .A2(n3261), .ZN(n3260) );
  INV_X1 U3867 ( .A(n5403), .ZN(n3261) );
  AND2_X1 U3868 ( .A1(n3180), .A2(n3987), .ZN(n3179) );
  INV_X1 U3869 ( .A(n5416), .ZN(n3180) );
  INV_X1 U3870 ( .A(n5429), .ZN(n3987) );
  NOR2_X1 U3871 ( .A1(n6906), .A2(n3189), .ZN(n3188) );
  NAND2_X1 U3872 ( .A1(n3257), .A2(n4426), .ZN(n3256) );
  INV_X1 U3873 ( .A(n3258), .ZN(n3257) );
  NOR2_X1 U3874 ( .A1(n6983), .A2(n3187), .ZN(n3186) );
  INV_X1 U3875 ( .A(n3870), .ZN(n3869) );
  NAND2_X1 U3876 ( .A1(n5491), .A2(n3177), .ZN(n3176) );
  INV_X1 U3877 ( .A(n5508), .ZN(n3177) );
  NOR2_X1 U3878 ( .A1(n5834), .A2(n3782), .ZN(n3192) );
  INV_X1 U3879 ( .A(n4050), .ZN(n4074) );
  NAND2_X1 U3880 ( .A1(n3175), .A2(n3156), .ZN(n5523) );
  AOI21_X1 U3881 ( .B1(n3752), .B2(n5664), .A(n3127), .ZN(n3175) );
  NAND2_X1 U3882 ( .A1(n5663), .A2(n3752), .ZN(n3156) );
  NOR2_X1 U3883 ( .A1(n3249), .A2(n3250), .ZN(n3248) );
  INV_X1 U3884 ( .A(n5551), .ZN(n3249) );
  INV_X1 U3885 ( .A(n3783), .ZN(n3781) );
  AND2_X1 U3886 ( .A1(n3704), .A2(n3255), .ZN(n3254) );
  INV_X1 U3887 ( .A(n5142), .ZN(n3255) );
  NOR2_X1 U3888 ( .A1(n3614), .A2(n4860), .ZN(n3592) );
  OR2_X1 U3889 ( .A1(n3519), .A2(n3518), .ZN(n4174) );
  NAND2_X1 U3890 ( .A1(n3628), .A2(n3630), .ZN(n3235) );
  OR2_X1 U3891 ( .A1(n3788), .A2(n3789), .ZN(n4792) );
  OAI21_X1 U3892 ( .B1(n3504), .B2(n3275), .A(n3508), .ZN(n3528) );
  OAI21_X1 U3893 ( .B1(n3504), .B2(n3246), .A(n3532), .ZN(n4937) );
  AOI22_X1 U3894 ( .A1(n3360), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3290) );
  NAND2_X1 U3895 ( .A1(n3378), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3299)
         );
  NAND2_X1 U3896 ( .A1(n3109), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3300) );
  XNOR2_X1 U3897 ( .A(n4630), .B(n4937), .ZN(n4742) );
  OR2_X1 U3898 ( .A1(n3544), .A2(n3543), .ZN(n4184) );
  INV_X1 U3899 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4785) );
  INV_X1 U3900 ( .A(n4134), .ZN(n4267) );
  NAND2_X1 U3901 ( .A1(n4307), .A2(n4306), .ZN(n4881) );
  INV_X1 U3902 ( .A(n4879), .ZN(n4307) );
  INV_X1 U3903 ( .A(n4832), .ZN(n4306) );
  OR2_X1 U3904 ( .A1(n4772), .A2(n4773), .ZN(n4626) );
  NOR2_X1 U3905 ( .A1(n5731), .A2(n5405), .ZN(n3185) );
  AND2_X1 U3906 ( .A1(n4008), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4009)
         );
  NAND2_X1 U3907 ( .A1(n3943), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3963)
         );
  NAND2_X1 U3908 ( .A1(n3943), .A2(n3188), .ZN(n3984) );
  NAND2_X1 U3909 ( .A1(n3161), .A2(n3266), .ZN(n4441) );
  INV_X1 U3910 ( .A(n4439), .ZN(n3161) );
  INV_X1 U3911 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6983) );
  NAND2_X1 U3912 ( .A1(n3869), .A2(n3186), .ZN(n3900) );
  NAND2_X1 U3913 ( .A1(n3869), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3873)
         );
  OR2_X1 U3914 ( .A1(n3852), .A2(n7008), .ZN(n3870) );
  NAND2_X1 U3915 ( .A1(n3781), .A2(n3190), .ZN(n3852) );
  AND2_X1 U3916 ( .A1(n3192), .A2(n3191), .ZN(n3190) );
  NOR2_X1 U3917 ( .A1(n5817), .A2(n5828), .ZN(n3191) );
  NAND2_X1 U3918 ( .A1(n3781), .A2(n3192), .ZN(n3821) );
  AND3_X1 U3919 ( .A1(n3787), .A2(n3786), .A3(n3785), .ZN(n5566) );
  INV_X1 U3920 ( .A(n5581), .ZN(n3247) );
  NAND2_X1 U3921 ( .A1(n3763), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3783)
         );
  INV_X1 U3922 ( .A(n3764), .ZN(n3763) );
  AND2_X1 U3923 ( .A1(n3125), .A2(n3649), .ZN(n3685) );
  NAND2_X1 U3924 ( .A1(n3145), .A2(n3133), .ZN(n5205) );
  NAND2_X1 U3925 ( .A1(n5091), .A2(n3233), .ZN(n3145) );
  NAND2_X1 U3926 ( .A1(n3649), .A2(n3124), .ZN(n3658) );
  AND2_X1 U3927 ( .A1(n3649), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3655)
         );
  AND2_X1 U3928 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3592), .ZN(n3649)
         );
  NAND2_X1 U3929 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3614) );
  NAND2_X1 U3930 ( .A1(n3627), .A2(n3626), .ZN(n4735) );
  NOR2_X1 U3931 ( .A1(n3230), .A2(n5407), .ZN(n3228) );
  NAND2_X1 U3932 ( .A1(n5430), .A2(n3229), .ZN(n5419) );
  NAND2_X1 U3933 ( .A1(n5430), .A2(n5432), .ZN(n5431) );
  AOI21_X1 U3934 ( .B1(n3243), .B2(n3245), .A(n3242), .ZN(n3241) );
  NAND2_X1 U3935 ( .A1(n3147), .A2(n3146), .ZN(n3151) );
  INV_X1 U3936 ( .A(n4244), .ZN(n3242) );
  AND2_X1 U3937 ( .A1(n4291), .A2(n4290), .ZN(n4377) );
  NOR2_X1 U3938 ( .A1(n5462), .A2(n3221), .ZN(n3220) );
  INV_X1 U3939 ( .A(n3223), .ZN(n3221) );
  AND2_X1 U3940 ( .A1(n3206), .A2(n3210), .ZN(n3205) );
  NAND2_X1 U3941 ( .A1(n5769), .A2(n3208), .ZN(n3207) );
  AOI21_X1 U3942 ( .B1(n3211), .B2(n3213), .A(n5793), .ZN(n3210) );
  NOR2_X1 U3943 ( .A1(n5483), .A2(n5482), .ZN(n5481) );
  INV_X1 U3944 ( .A(n5786), .ZN(n5792) );
  AND2_X1 U3945 ( .A1(n4366), .A2(n4365), .ZN(n5510) );
  OR2_X1 U3946 ( .A1(n3217), .A2(n3219), .ZN(n3216) );
  INV_X1 U3947 ( .A(n5538), .ZN(n3219) );
  INV_X1 U3948 ( .A(n5833), .ZN(n5814) );
  NAND2_X1 U3949 ( .A1(n3147), .A2(n3149), .ZN(n5833) );
  OR2_X1 U3950 ( .A1(n5568), .A2(n5571), .ZN(n5569) );
  NAND2_X1 U3951 ( .A1(n3204), .A2(n3202), .ZN(n3201) );
  CLKBUF_X1 U3952 ( .A(n5579), .Z(n5668) );
  AND2_X1 U3953 ( .A1(n4338), .A2(n4337), .ZN(n5364) );
  OR2_X1 U3954 ( .A1(n5202), .A2(n6165), .ZN(n3227) );
  OR3_X1 U3955 ( .A1(n5022), .A2(n5136), .A3(n5202), .ZN(n6164) );
  NAND2_X1 U3956 ( .A1(n5891), .A2(n5890), .ZN(n5889) );
  CLKBUF_X1 U3957 ( .A(n5022), .Z(n5135) );
  NAND2_X1 U3958 ( .A1(n6119), .A2(n4872), .ZN(n4147) );
  NAND2_X1 U3959 ( .A1(n3393), .A2(n3392), .ZN(n4378) );
  INV_X1 U3960 ( .A(n3501), .ZN(n3443) );
  NOR2_X1 U3961 ( .A1(n5028), .A2(n5029), .ZN(n6449) );
  OR2_X1 U3962 ( .A1(n6104), .A2(n4888), .ZN(n4940) );
  AND3_X1 U3963 ( .A1(n6781), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6526) );
  INV_X1 U3964 ( .A(n5219), .ZN(n5217) );
  AOI21_X1 U3965 ( .B1(n5217), .B2(n6594), .A(n6659), .ZN(n6567) );
  AND2_X1 U3966 ( .A1(n5314), .A2(n4743), .ZN(n6598) );
  AND2_X1 U3967 ( .A1(n4888), .A2(n5218), .ZN(n6589) );
  AND2_X1 U3968 ( .A1(n5029), .A2(n4980), .ZN(n4984) );
  INV_X1 U3969 ( .A(n6109), .ZN(n6659) );
  AND2_X1 U3970 ( .A1(n4984), .A2(n5218), .ZN(n5252) );
  INV_X1 U3971 ( .A(n4158), .ZN(n4909) );
  NAND2_X1 U3972 ( .A1(n4900), .A2(n4899), .ZN(n4930) );
  INV_X1 U3973 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6781) );
  AND2_X1 U3974 ( .A1(n5369), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4138) );
  AND2_X1 U3975 ( .A1(n4872), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4715) );
  INV_X1 U3976 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n4872) );
  AND2_X1 U3977 ( .A1(n5389), .A2(n3195), .ZN(n6175) );
  AND2_X1 U3978 ( .A1(n6184), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3195) );
  AND2_X1 U3979 ( .A1(n6184), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6241) );
  INV_X1 U3980 ( .A(n6190), .ZN(n6227) );
  OR2_X1 U3981 ( .A1(n5628), .A2(n5385), .ZN(n6210) );
  AND2_X1 U3982 ( .A1(n5621), .A2(n6193), .ZN(n6214) );
  INV_X1 U3983 ( .A(n6241), .ZN(n6259) );
  INV_X1 U3984 ( .A(n6214), .ZN(n6255) );
  NOR2_X1 U3985 ( .A1(n5381), .A2(n5672), .ZN(n4544) );
  INV_X1 U3986 ( .A(n5672), .ZN(n6261) );
  INV_X1 U3987 ( .A(n6266), .ZN(n5659) );
  INV_X1 U3988 ( .A(n5715), .ZN(n5718) );
  OR2_X1 U3989 ( .A1(n5711), .A2(n5712), .ZN(n5719) );
  OR2_X1 U3990 ( .A1(n4851), .A2(n4854), .ZN(n6232) );
  INV_X1 U3991 ( .A(n5719), .ZN(n5716) );
  NAND2_X2 U3992 ( .A1(n5715), .A2(n4847), .ZN(n5721) );
  NAND2_X1 U3993 ( .A1(n6310), .A2(n4712), .ZN(n4714) );
  OR2_X1 U3994 ( .A1(n4711), .A2(n4710), .ZN(n4712) );
  INV_X1 U3995 ( .A(n6285), .ZN(n6295) );
  NAND2_X1 U3996 ( .A1(n4610), .A2(n4609), .ZN(n6308) );
  AND2_X1 U3997 ( .A1(n4608), .A2(n6310), .ZN(n6319) );
  INV_X1 U3998 ( .A(n6308), .ZN(n6304) );
  INV_X1 U3999 ( .A(n4532), .ZN(n4533) );
  INV_X1 U4000 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6906) );
  INV_X1 U4001 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5828) );
  AND2_X1 U4002 ( .A1(n3705), .A2(n3126), .ZN(n3736) );
  NAND2_X1 U4003 ( .A1(n3705), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3706)
         );
  INV_X1 U4004 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4860) );
  INV_X1 U4005 ( .A(n6334), .ZN(n6358) );
  NAND2_X1 U4006 ( .A1(n3167), .A2(n3168), .ZN(n3170) );
  AOI21_X1 U4007 ( .B1(n5738), .B2(n3173), .A(n5722), .ZN(n3167) );
  NAND2_X1 U4008 ( .A1(n3144), .A2(n3172), .ZN(n3171) );
  AND2_X1 U4009 ( .A1(n5722), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3172)
         );
  NAND2_X1 U4010 ( .A1(n5738), .A2(n3166), .ZN(n3169) );
  AND2_X1 U4011 ( .A1(n5722), .A2(n3173), .ZN(n3166) );
  INV_X1 U4012 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6913) );
  INV_X1 U4013 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6022) );
  NAND2_X1 U4014 ( .A1(n4236), .A2(n4235), .ZN(n5841) );
  NAND2_X1 U4015 ( .A1(n6338), .A2(n6337), .ZN(n6336) );
  NAND2_X1 U4016 ( .A1(n5091), .A2(n4198), .ZN(n6338) );
  OR2_X1 U4017 ( .A1(n4147), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6423) );
  INV_X1 U4019 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5369) );
  CLKBUF_X1 U4020 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n6756) );
  INV_X1 U4021 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4634) );
  NOR2_X1 U4022 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6119) );
  INV_X1 U4023 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5082) );
  INV_X1 U4024 ( .A(n5075), .ZN(n5307) );
  NOR4_X1 U4025 ( .A1(n5074), .A2(n6647), .A3(n5073), .A4(n6493), .ZN(n5290)
         );
  INV_X1 U4026 ( .A(n5310), .ZN(n5060) );
  OAI21_X1 U4027 ( .B1(n5102), .B2(n5105), .A(n5158), .ZN(n5127) );
  INV_X1 U4028 ( .A(n5357), .ZN(n5244) );
  NOR2_X2 U4029 ( .A1(n5217), .A2(n5218), .ZN(n6584) );
  AND2_X1 U4030 ( .A1(n5219), .A2(n5218), .ZN(n5357) );
  NOR2_X1 U4031 ( .A1(n4924), .A2(n5100), .ZN(n6654) );
  NOR2_X1 U4032 ( .A1(n4913), .A2(n5100), .ZN(n6671) );
  NOR2_X1 U4033 ( .A1(n6822), .A2(n5100), .ZN(n6677) );
  NOR2_X1 U4034 ( .A1(n4904), .A2(n5100), .ZN(n6689) );
  NOR2_X1 U4035 ( .A1(n4898), .A2(n5100), .ZN(n6695) );
  NOR2_X1 U4036 ( .A1(n4920), .A2(n5100), .ZN(n6701) );
  OAI211_X1 U4037 ( .C1(n6594), .C2(n6652), .A(n4988), .B(n6523), .ZN(n5018)
         );
  AND2_X1 U4038 ( .A1(n4984), .A2(n4157), .ZN(n6710) );
  AOI21_X1 U4039 ( .B1(n6652), .B2(STATE2_REG_2__SCAN_IN), .A(n4979), .ZN(
        n5021) );
  AND2_X1 U4040 ( .A1(n5260), .A2(n5259), .ZN(n5284) );
  INV_X1 U4041 ( .A(n5252), .ZN(n5289) );
  INV_X1 U4042 ( .A(n6654), .ZN(n5348) );
  OR2_X1 U4043 ( .A1(n4930), .A2(n4925), .ZN(n6590) );
  INV_X1 U4044 ( .A(n6671), .ZN(n5353) );
  INV_X1 U4045 ( .A(n6677), .ZN(n5338) );
  OR2_X1 U4046 ( .A1(n4930), .A2(n4274), .ZN(n6613) );
  INV_X1 U4047 ( .A(n6683), .ZN(n5343) );
  OR2_X1 U4048 ( .A1(n4930), .A2(n4909), .ZN(n6618) );
  NAND2_X1 U4049 ( .A1(n6349), .A2(DATAI_20_), .ZN(n6624) );
  INV_X1 U4050 ( .A(n6695), .ZN(n5325) );
  OR2_X1 U4051 ( .A1(n4930), .A2(n3410), .ZN(n6628) );
  NAND2_X1 U4052 ( .A1(n6349), .A2(DATAI_21_), .ZN(n6632) );
  OR2_X1 U4053 ( .A1(n4930), .A2(n3634), .ZN(n7072) );
  INV_X1 U4054 ( .A(n6701), .ZN(n7081) );
  NAND2_X1 U4055 ( .A1(n6349), .A2(DATAI_22_), .ZN(n7073) );
  INV_X1 U4056 ( .A(n6708), .ZN(n5333) );
  AND2_X1 U4057 ( .A1(n4897), .A2(n4896), .ZN(n4932) );
  OR2_X1 U4058 ( .A1(n4930), .A2(n5374), .ZN(n6637) );
  OAI211_X1 U4059 ( .C1(n5255), .C2(n6594), .A(n4893), .B(n6523), .ZN(n4929)
         );
  AND3_X1 U4060 ( .A1(n5029), .A2(n5311), .A3(n6518), .ZN(n5286) );
  NAND2_X1 U4061 ( .A1(n4772), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6121) );
  AND2_X1 U4062 ( .A1(n4815), .A2(n4814), .ZN(n6722) );
  NOR2_X1 U4063 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6747) );
  INV_X1 U4064 ( .A(n6722), .ZN(n4967) );
  AND2_X1 U4065 ( .A1(n4574), .A2(n4598), .ZN(n6730) );
  OR2_X1 U4066 ( .A1(n4261), .A2(STATE_REG_0__SCAN_IN), .ZN(n4767) );
  INV_X1 U4067 ( .A(STATE_REG_1__SCAN_IN), .ZN(n4573) );
  OR2_X1 U4068 ( .A1(n5914), .A2(n5672), .ZN(n4482) );
  OAI21_X1 U4069 ( .B1(n5895), .B2(n6334), .A(n3236), .ZN(U2955) );
  AOI21_X1 U4070 ( .B1(n5733), .B2(n6349), .A(n5732), .ZN(n5734) );
  OAI211_X1 U4071 ( .C1(n5969), .C2(n6334), .A(n3159), .B(n3158), .ZN(U2963)
         );
  AOI21_X1 U4072 ( .B1(n6330), .B2(n5791), .A(n5790), .ZN(n3158) );
  NAND2_X1 U4073 ( .A1(n3160), .A2(n6349), .ZN(n3159) );
  OAI21_X1 U4074 ( .B1(n5653), .B2(n6397), .A(n4493), .ZN(n4494) );
  AND2_X2 U4075 ( .A1(n3277), .A2(n3326), .ZN(n3462) );
  OR2_X1 U4076 ( .A1(n5506), .A2(n3122), .ZN(n5427) );
  AND2_X1 U4077 ( .A1(n4229), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3120)
         );
  NAND2_X1 U4078 ( .A1(n5581), .A2(n3248), .ZN(n5535) );
  NOR2_X1 U4079 ( .A1(n5144), .A2(n3226), .ZN(n5363) );
  OAI21_X1 U4080 ( .B1(n3423), .B2(n3397), .A(n3418), .ZN(n3431) );
  OR2_X1 U4081 ( .A1(n3256), .A2(n3176), .ZN(n3121) );
  OAI211_X1 U4082 ( .C1(n5082), .C2(n4122), .A(n3479), .B(n3475), .ZN(n3621)
         );
  NAND2_X1 U4083 ( .A1(n5662), .A2(n3752), .ZN(n5581) );
  OR2_X1 U4084 ( .A1(n5663), .A2(n5664), .ZN(n5662) );
  OR2_X1 U4085 ( .A1(n3121), .A2(n3966), .ZN(n3122) );
  AND2_X1 U4086 ( .A1(n3254), .A2(n3253), .ZN(n3123) );
  AND2_X1 U4087 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3124) );
  AND2_X1 U4088 ( .A1(n3124), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3125)
         );
  AND2_X1 U4089 ( .A1(n3183), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3126)
         );
  OR2_X1 U4090 ( .A1(n3181), .A2(n5537), .ZN(n3127) );
  INV_X2 U4091 ( .A(n5888), .ZN(n6349) );
  AND2_X1 U4092 ( .A1(n3186), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3128)
         );
  AND2_X1 U4093 ( .A1(n3188), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3129)
         );
  NAND2_X1 U4094 ( .A1(n5889), .A2(n4227), .ZN(n5861) );
  NAND2_X1 U4095 ( .A1(n5848), .A2(n4238), .ZN(n3130) );
  NOR2_X1 U4096 ( .A1(n3247), .A2(n3250), .ZN(n5550) );
  NAND2_X1 U4097 ( .A1(n3107), .A2(n4234), .ZN(n3131) );
  AND2_X1 U4098 ( .A1(n4207), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3132)
         );
  OAI21_X1 U4099 ( .B1(n5891), .B2(n3203), .A(n3200), .ZN(n5856) );
  NAND2_X1 U4100 ( .A1(n3240), .A2(n4233), .ZN(n5847) );
  INV_X1 U4102 ( .A(n3442), .ZN(n4380) );
  NAND2_X1 U4103 ( .A1(n3417), .A2(n4151), .ZN(n3434) );
  XNOR2_X1 U4104 ( .A(n4199), .B(n3584), .ZN(n4208) );
  AND2_X1 U4105 ( .A1(n5206), .A2(n3162), .ZN(n3133) );
  NAND2_X1 U4106 ( .A1(n3752), .A2(n3157), .ZN(n5663) );
  AND2_X1 U4107 ( .A1(n3130), .A2(n4237), .ZN(n3134) );
  AND2_X1 U4108 ( .A1(n4189), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3135)
         );
  AND2_X1 U4109 ( .A1(n4089), .A2(n4620), .ZN(n4209) );
  INV_X1 U4110 ( .A(n4209), .ZN(n4219) );
  OR2_X1 U4111 ( .A1(n5506), .A2(n3176), .ZN(n4439) );
  AND2_X2 U4112 ( .A1(n4788), .A2(n4745), .ZN(n3378) );
  AND2_X1 U4113 ( .A1(n4461), .A2(n5442), .ZN(n5430) );
  OR2_X1 U4114 ( .A1(n3106), .A2(n6035), .ZN(n3136) );
  INV_X1 U4115 ( .A(n3213), .ZN(n3212) );
  NAND2_X1 U4116 ( .A1(n3106), .A2(n4250), .ZN(n3213) );
  NOR2_X1 U4117 ( .A1(n5506), .A2(n3121), .ZN(n3137) );
  INV_X1 U4118 ( .A(n3239), .ZN(n3238) );
  NAND2_X1 U4119 ( .A1(n3131), .A2(n4233), .ZN(n3239) );
  NOR2_X1 U4120 ( .A1(n5506), .A2(n5508), .ZN(n5490) );
  INV_X1 U4121 ( .A(n3244), .ZN(n3243) );
  OAI21_X1 U4122 ( .B1(n3130), .B2(n3245), .A(n4241), .ZN(n3244) );
  NAND2_X1 U4123 ( .A1(n3326), .A2(n4745), .ZN(n4750) );
  INV_X1 U4124 ( .A(n3833), .ZN(n3659) );
  NAND2_X1 U4125 ( .A1(n3546), .A2(n3545), .ZN(n6518) );
  AND2_X1 U4126 ( .A1(n3705), .A2(n3183), .ZN(n3138) );
  NOR2_X1 U4127 ( .A1(n5568), .A2(n3217), .ZN(n3139) );
  OR2_X1 U4128 ( .A1(n5022), .A2(n5136), .ZN(n5137) );
  NAND2_X1 U4129 ( .A1(n3222), .A2(n3223), .ZN(n4485) );
  NAND2_X1 U4130 ( .A1(n4529), .A2(n6184), .ZN(n6193) );
  INV_X1 U4131 ( .A(n6193), .ZN(n6204) );
  OR2_X1 U4132 ( .A1(n5144), .A2(n5147), .ZN(n5145) );
  AND2_X1 U4133 ( .A1(n3647), .A2(n3582), .ZN(n3140) );
  INV_X1 U4134 ( .A(n3230), .ZN(n3229) );
  OR2_X1 U4135 ( .A1(n5417), .A2(n3231), .ZN(n3230) );
  INV_X1 U4136 ( .A(n3966), .ZN(n5441) );
  AND2_X1 U4137 ( .A1(n4532), .A2(n3260), .ZN(n3141) );
  AND2_X1 U4138 ( .A1(n3721), .A2(n3720), .ZN(n5142) );
  AOI21_X1 U4139 ( .B1(n5870), .B2(n4502), .A(n3735), .ZN(n5250) );
  INV_X1 U4140 ( .A(n5250), .ZN(n3253) );
  INV_X1 U4141 ( .A(n5525), .ZN(n3837) );
  INV_X1 U4142 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3189) );
  INV_X1 U4143 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3187) );
  INV_X1 U4144 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6853) );
  AND2_X1 U4145 ( .A1(n3185), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n3142)
         );
  OAI33_X1 U4146 ( .A1(n4743), .A2(n6657), .A3(n6655), .B1(n6563), .B2(n6490), 
        .B3(n6645), .ZN(n3143) );
  XNOR2_X1 U4147 ( .A(n6651), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6645)
         );
  AND2_X1 U4148 ( .A1(n3529), .A2(n4931), .ZN(n6563) );
  NAND2_X1 U4149 ( .A1(n3144), .A2(n5738), .ZN(n5728) );
  NAND2_X1 U4150 ( .A1(n3144), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3168) );
  OAI22_X2 U4151 ( .A1(n3144), .A2(n4248), .B1(n5738), .B2(n4247), .ZN(n3237)
         );
  NAND2_X2 U4152 ( .A1(n5205), .A2(n4217), .ZN(n5891) );
  INV_X1 U4153 ( .A(n6344), .ZN(n3154) );
  NAND2_X1 U4154 ( .A1(n6345), .A2(n6344), .ZN(n6347) );
  NAND2_X1 U4155 ( .A1(n4865), .A2(n4182), .ZN(n6345) );
  NAND2_X1 U4156 ( .A1(n4190), .A2(n3778), .ZN(n3155) );
  OR2_X2 U4157 ( .A1(n5461), .A2(n4425), .ZN(n5789) );
  INV_X2 U4158 ( .A(n3648), .ZN(n3571) );
  NAND2_X1 U4159 ( .A1(n3602), .A2(n3252), .ZN(n3648) );
  NAND2_X1 U4160 ( .A1(n3164), .A2(n3163), .ZN(n3162) );
  INV_X1 U4161 ( .A(n3132), .ZN(n3163) );
  NAND2_X2 U4162 ( .A1(n3571), .A2(n3140), .ZN(n4199) );
  NAND2_X1 U4163 ( .A1(n3165), .A2(n5912), .ZN(U2988) );
  NAND4_X1 U4164 ( .A1(n3170), .A2(n3171), .A3(n6440), .A4(n3169), .ZN(n3165)
         );
  NAND3_X1 U4165 ( .A1(n3170), .A2(n3171), .A3(n3169), .ZN(n5913) );
  INV_X1 U4166 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3173) );
  NAND3_X1 U4167 ( .A1(n3526), .A2(n6518), .A3(n3611), .ZN(n3174) );
  NAND2_X1 U4168 ( .A1(n4183), .A2(n3778), .ZN(n3600) );
  NAND2_X1 U4169 ( .A1(n3988), .A2(n3987), .ZN(n5415) );
  AND2_X2 U4170 ( .A1(n3988), .A2(n3179), .ZN(n5402) );
  INV_X1 U4171 ( .A(n5523), .ZN(n3838) );
  NAND2_X1 U4172 ( .A1(n4009), .A2(n3142), .ZN(n4146) );
  NAND2_X1 U4173 ( .A1(n3943), .A2(n3129), .ZN(n4007) );
  INV_X1 U4174 ( .A(n3527), .ZN(n3193) );
  OAI21_X2 U4175 ( .B1(n3438), .B2(n4380), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3504) );
  AND2_X2 U4176 ( .A1(n3201), .A2(n4231), .ZN(n3200) );
  NAND2_X2 U4177 ( .A1(n3199), .A2(n3197), .ZN(n3240) );
  NAND2_X1 U4178 ( .A1(n3222), .A2(n3220), .ZN(n4376) );
  NOR2_X2 U4179 ( .A1(n5144), .A2(n3225), .ZN(n5579) );
  AND2_X4 U4181 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4745) );
  NOR2_X4 U4182 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4788) );
  OAI21_X1 U4183 ( .B1(n5091), .B2(n3164), .A(n3232), .ZN(n5207) );
  AOI21_X1 U4184 ( .B1(n6337), .B2(n3234), .A(n3132), .ZN(n3232) );
  NOR2_X1 U4185 ( .A1(n3132), .A2(n3234), .ZN(n3233) );
  NAND2_X1 U4186 ( .A1(n3571), .A2(n3647), .ZN(n3654) );
  NAND2_X1 U4187 ( .A1(n5581), .A2(n5582), .ZN(n5565) );
  AND3_X2 U4188 ( .A1(n5067), .A2(n3123), .A3(n5068), .ZN(n3740) );
  NAND3_X1 U4189 ( .A1(n5067), .A2(n5068), .A3(n3254), .ZN(n5140) );
  NAND3_X1 U4190 ( .A1(n5067), .A2(n5068), .A3(n3704), .ZN(n5141) );
  NAND2_X1 U4191 ( .A1(n5402), .A2(n5403), .ZN(n4449) );
  NAND2_X1 U4192 ( .A1(n5402), .A2(n3141), .ZN(n3262) );
  NAND2_X1 U4193 ( .A1(n3628), .A2(n3631), .ZN(n3629) );
  NAND2_X1 U4194 ( .A1(n4449), .A2(n4450), .ZN(n4452) );
  INV_X1 U4195 ( .A(READY_N), .ZN(n4811) );
  INV_X1 U4196 ( .A(n4826), .ZN(n3644) );
  AND2_X2 U4197 ( .A1(n4715), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6744) );
  INV_X1 U4198 ( .A(n5670), .ZN(n6262) );
  OR2_X1 U4199 ( .A1(n3407), .A2(n6756), .ZN(n3263) );
  AND4_X1 U4200 ( .A1(n3282), .A2(n3281), .A3(n3280), .A4(n3279), .ZN(n3264)
         );
  NAND2_X1 U4201 ( .A1(n5072), .A2(n6603), .ZN(n6655) );
  INV_X1 U4202 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5090) );
  NOR2_X1 U4203 ( .A1(n3585), .A2(n6603), .ZN(n3833) );
  INV_X1 U4204 ( .A(n4598), .ZN(n6752) );
  INV_X1 U4205 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6159) );
  AND3_X1 U4206 ( .A1(n3703), .A2(n3702), .A3(n3701), .ZN(n3265) );
  AND2_X1 U4207 ( .A1(n5480), .A2(n4442), .ZN(n3266) );
  INV_X1 U4208 ( .A(n4845), .ZN(n3392) );
  AND2_X1 U4209 ( .A1(n6119), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3267) );
  INV_X1 U4210 ( .A(n3411), .ZN(n3405) );
  OR2_X1 U4211 ( .A1(n3556), .A2(n3555), .ZN(n4191) );
  OR2_X1 U4212 ( .A1(n4750), .A2(n3327), .ZN(n3328) );
  NOR2_X1 U4213 ( .A1(n3493), .A2(n4872), .ZN(n4218) );
  INV_X1 U4214 ( .A(n3437), .ZN(n3441) );
  OR2_X1 U4215 ( .A1(n3362), .A2(n3361), .ZN(n3365) );
  OR2_X1 U4216 ( .A1(n4124), .A2(n4123), .ZN(n4126) );
  BUF_X1 U4217 ( .A(n3403), .Z(n4089) );
  NAND2_X1 U4218 ( .A1(n4839), .A2(n3391), .ZN(n4662) );
  INV_X1 U4219 ( .A(n3461), .ZN(n4122) );
  AND2_X1 U4220 ( .A1(n4126), .A2(n4125), .ZN(n4134) );
  INV_X1 U4221 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n7008) );
  NAND2_X1 U4222 ( .A1(n6603), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3801) );
  INV_X1 U4223 ( .A(n5571), .ZN(n4347) );
  NOR2_X1 U4224 ( .A1(n4220), .A2(n4219), .ZN(n4221) );
  INV_X1 U4225 ( .A(n4662), .ZN(n3393) );
  NAND2_X1 U4226 ( .A1(n3461), .A2(n4209), .ZN(n4135) );
  OAI211_X1 U4227 ( .C1(n4122), .C2(n5090), .A(n3494), .B(n3493), .ZN(n3631)
         );
  INV_X1 U4228 ( .A(n5136), .ZN(n4323) );
  NOR2_X1 U4229 ( .A1(n4792), .A2(n4872), .ZN(n4050) );
  NAND2_X1 U4230 ( .A1(n3403), .A2(n3445), .ZN(n3409) );
  NAND2_X1 U4231 ( .A1(n4249), .A2(n4434), .ZN(n4435) );
  AND2_X1 U4232 ( .A1(n4352), .A2(n4351), .ZN(n5552) );
  AND2_X1 U4233 ( .A1(n4785), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6456)
         );
  OR2_X1 U4234 ( .A1(n5100), .A2(n5099), .ZN(n5254) );
  INV_X1 U4235 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6847) );
  AND2_X1 U4236 ( .A1(n6144), .A2(n6184), .ZN(n6253) );
  AND2_X1 U4237 ( .A1(n4326), .A2(n4325), .ZN(n5202) );
  INV_X1 U4238 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5817) );
  NAND3_X1 U4240 ( .A1(n5760), .A2(n4246), .A3(n5757), .ZN(n5738) );
  INV_X1 U4241 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6035) );
  INV_X1 U4242 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6858) );
  OR2_X1 U4243 ( .A1(n4711), .A2(n4276), .ZN(n4277) );
  NAND2_X1 U4244 ( .A1(n6121), .A2(n4871), .ZN(n4900) );
  AND2_X1 U4245 ( .A1(n6455), .A2(n6483), .ZN(n6461) );
  OR2_X1 U4246 ( .A1(n6460), .A2(n6651), .ZN(n6483) );
  NOR2_X1 U4247 ( .A1(n5254), .A2(n5101), .ZN(n5158) );
  OR2_X1 U4248 ( .A1(n6104), .A2(n5154), .ZN(n6551) );
  AND2_X1 U4249 ( .A1(n6593), .A2(n5212), .ZN(n5219) );
  INV_X1 U4250 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4975) );
  OR2_X1 U4251 ( .A1(n4930), .A2(n3111), .ZN(n6608) );
  AND2_X1 U4252 ( .A1(n4761), .A2(n4760), .ZN(n4870) );
  OR2_X1 U4253 ( .A1(n4711), .A2(n4281), .ZN(n4605) );
  OR2_X1 U4254 ( .A1(n5467), .A2(n4521), .ZN(n5436) );
  NOR2_X1 U4255 ( .A1(n5389), .A2(n5369), .ZN(n4529) );
  INV_X1 U4256 ( .A(n6253), .ZN(n6186) );
  NOR2_X1 U4257 ( .A1(n6266), .A2(n5393), .ZN(n4543) );
  NAND2_X1 U4258 ( .A1(n4626), .A2(n4455), .ZN(n4456) );
  AND2_X1 U4259 ( .A1(n5715), .A2(n4848), .ZN(n5712) );
  AND2_X1 U4260 ( .A1(n6288), .A2(n4287), .ZN(n6272) );
  AND2_X1 U4261 ( .A1(n4714), .A2(n4713), .ZN(n6288) );
  AND2_X1 U4262 ( .A1(n4620), .A2(n4811), .ZN(n4609) );
  OR2_X1 U4263 ( .A1(n4273), .A2(n6746), .ZN(n4813) );
  INV_X1 U4264 ( .A(n6310), .ZN(n6323) );
  OAI21_X1 U4265 ( .B1(n5697), .B2(n5888), .A(n4445), .ZN(n4446) );
  INV_X1 U4266 ( .A(n6363), .ZN(n6330) );
  AND2_X1 U4267 ( .A1(n4703), .A2(n4702), .ZN(n6256) );
  AND2_X1 U4268 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5916) );
  INV_X1 U4269 ( .A(n5983), .ZN(n6443) );
  INV_X1 U4270 ( .A(n6412), .ZN(n6440) );
  AND2_X2 U4271 ( .A1(n4404), .A2(n4379), .ZN(n6435) );
  NOR2_X1 U4272 ( .A1(n4775), .A2(n3111), .ZN(n5367) );
  AND2_X1 U4273 ( .A1(n5076), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6647) );
  OAI211_X1 U4274 ( .C1(n6594), .C2(n5037), .A(n5036), .B(n6523), .ZN(n5061)
         );
  INV_X1 U4275 ( .A(n6489), .ZN(n5131) );
  OAI21_X1 U4276 ( .B1(n6497), .B2(n6496), .A(n6495), .ZN(n6514) );
  OAI211_X1 U4277 ( .C1(n6594), .C2(n6491), .A(n4944), .B(n6523), .ZN(n7078)
         );
  INV_X1 U4278 ( .A(n6551), .ZN(n5188) );
  OAI21_X1 U4279 ( .B1(n6567), .B2(n6566), .A(n6565), .ZN(n6585) );
  OAI211_X1 U4280 ( .C1(n6567), .C2(n5222), .A(n6523), .B(n5221), .ZN(n5246)
         );
  OAI211_X1 U4281 ( .C1(n5322), .C2(n6598), .A(n5321), .B(n5320), .ZN(n5358)
         );
  AND2_X1 U4282 ( .A1(n4888), .A2(n4157), .ZN(n5311) );
  INV_X1 U4283 ( .A(n6663), .ZN(n6706) );
  NOR2_X1 U4284 ( .A1(n4908), .A2(n5100), .ZN(n6683) );
  NOR2_X1 U4285 ( .A1(n5069), .A2(n5100), .ZN(n6708) );
  INV_X1 U4286 ( .A(n6619), .ZN(n6684) );
  INV_X1 U4287 ( .A(n6638), .ZN(n6711) );
  INV_X1 U4288 ( .A(n6681), .ZN(n5335) );
  INV_X1 U4289 ( .A(n6705), .ZN(n7077) );
  INV_X1 U4290 ( .A(STATE_REG_0__SCAN_IN), .ZN(n4555) );
  INV_X1 U4291 ( .A(STATE_REG_2__SCAN_IN), .ZN(n4563) );
  AND2_X1 U4292 ( .A1(n4605), .A2(n4606), .ZN(n6741) );
  INV_X1 U4293 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6129) );
  INV_X1 U4294 ( .A(n6166), .ZN(n6244) );
  AND4_X1 U4295 ( .A1(n5632), .A2(n5631), .A3(n5630), .A4(n5629), .ZN(n5633)
         );
  AND2_X1 U4296 ( .A1(n4482), .A2(n4481), .ZN(n4483) );
  AND2_X2 U4297 ( .A1(n4456), .A2(n6717), .ZN(n6266) );
  INV_X1 U4298 ( .A(n5210), .ZN(n6194) );
  NAND2_X1 U4299 ( .A1(n6308), .A2(n4844), .ZN(n5715) );
  INV_X1 U4300 ( .A(n6272), .ZN(n4729) );
  OR2_X1 U4301 ( .A1(n6288), .A2(n6744), .ZN(n6285) );
  INV_X1 U4302 ( .A(n6288), .ZN(n6297) );
  INV_X1 U4303 ( .A(DATAI_0_), .ZN(n4924) );
  OR2_X1 U4304 ( .A1(n4711), .A2(n4813), .ZN(n6310) );
  INV_X1 U4305 ( .A(n6319), .ZN(n6325) );
  INV_X1 U4306 ( .A(n4431), .ZN(n4432) );
  OR2_X1 U4307 ( .A1(n6724), .A2(n6655), .ZN(n5888) );
  NAND2_X1 U4308 ( .A1(n5884), .A2(n4704), .ZN(n6363) );
  INV_X1 U4309 ( .A(n4494), .ZN(n4495) );
  INV_X1 U4310 ( .A(n6435), .ZN(n6397) );
  INV_X1 U4311 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6389) );
  NAND2_X1 U4312 ( .A1(n4404), .A2(n4286), .ZN(n6412) );
  OAI21_X1 U4313 ( .B1(n4873), .B2(n6723), .A(n5100), .ZN(n6448) );
  NOR2_X1 U4314 ( .A1(n4632), .A2(n4899), .ZN(n6125) );
  NAND2_X1 U4315 ( .A1(n5032), .A2(n4157), .ZN(n5310) );
  AOI22_X1 U4316 ( .A1(n5035), .A2(n5031), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5037), .ZN(n5064) );
  INV_X1 U4317 ( .A(n5097), .ZN(n5134) );
  NAND2_X1 U4318 ( .A1(n6449), .A2(n5311), .ZN(n6489) );
  NAND2_X1 U4319 ( .A1(n6449), .A2(n6589), .ZN(n6517) );
  AOI22_X1 U4320 ( .A1(n4943), .A2(n4939), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6491), .ZN(n7082) );
  INV_X1 U4321 ( .A(n5155), .ZN(n7074) );
  OR2_X1 U4322 ( .A1(n6519), .A2(n6518), .ZN(n6588) );
  AOI22_X1 U4323 ( .A1(n5216), .A2(n5222), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5215), .ZN(n5249) );
  AOI22_X1 U4324 ( .A1(n5317), .A2(n6598), .B1(n6645), .B2(n5316), .ZN(n5362)
         );
  NAND2_X1 U4325 ( .A1(n6593), .A2(n5311), .ZN(n6644) );
  NAND2_X1 U4326 ( .A1(n6593), .A2(n6589), .ZN(n6715) );
  INV_X1 U4327 ( .A(n6689), .ZN(n5361) );
  NAND2_X1 U4328 ( .A1(n6349), .A2(DATAI_25_), .ZN(n6675) );
  NAND2_X1 U4329 ( .A1(n6349), .A2(DATAI_30_), .ZN(n6705) );
  NAND2_X1 U4330 ( .A1(n6349), .A2(DATAI_18_), .ZN(n6617) );
  NAND2_X1 U4331 ( .A1(n6349), .A2(DATAI_23_), .ZN(n6638) );
  INV_X1 U4332 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n5072) );
  INV_X1 U4333 ( .A(n6730), .ZN(n6726) );
  INV_X1 U4334 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6395) );
  INV_X1 U4335 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6158) );
  OAI21_X1 U4336 ( .B1(n5679), .B2(n5670), .A(n4483), .ZN(U2830) );
  AND2_X2 U4337 ( .A1(n3276), .A2(n4744), .ZN(n3991) );
  AND2_X4 U4338 ( .A1(n3269), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3326)
         );
  AOI22_X1 U4339 ( .A1(n3991), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3274) );
  AND2_X4 U4340 ( .A1(n3277), .A2(n3276), .ZN(n3446) );
  AND2_X2 U4341 ( .A1(n3276), .A2(n4745), .ZN(n4055) );
  AOI22_X1 U4342 ( .A1(n4055), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3272) );
  AND2_X2 U4343 ( .A1(n4744), .A2(n4677), .ZN(n3463) );
  AND2_X4 U4344 ( .A1(n4677), .A2(n4745), .ZN(n4040) );
  AOI22_X1 U4345 ( .A1(n3463), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3271) );
  INV_X1 U4346 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3275) );
  AND2_X2 U4347 ( .A1(n3275), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3278)
         );
  AND2_X2 U4348 ( .A1(n3276), .A2(n3278), .ZN(n4033) );
  AND2_X4 U4349 ( .A1(n3326), .A2(n4745), .ZN(n3452) );
  AOI22_X1 U4350 ( .A1(n4033), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3282) );
  AND2_X2 U4351 ( .A1(n3278), .A2(n4788), .ZN(n3360) );
  AOI22_X1 U4352 ( .A1(n3360), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3281) );
  AND2_X4 U4353 ( .A1(n3278), .A2(n3326), .ZN(n3996) );
  INV_X2 U4354 ( .A(n3362), .ZN(n3379) );
  AOI22_X1 U4355 ( .A1(n3996), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3379), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3280) );
  AND2_X2 U4356 ( .A1(n3278), .A2(n4677), .ZN(n3447) );
  AOI22_X1 U4357 ( .A1(n3447), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3279) );
  NAND2_X2 U4358 ( .A1(n3283), .A2(n3264), .ZN(n3394) );
  INV_X2 U4359 ( .A(n3394), .ZN(n4274) );
  AOI22_X1 U4360 ( .A1(n3447), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3287) );
  AOI22_X1 U4361 ( .A1(n4033), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4362 ( .A1(n3991), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3285) );
  AOI22_X1 U4363 ( .A1(n4055), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3284) );
  NAND4_X1 U4364 ( .A1(n3287), .A2(n3286), .A3(n3285), .A4(n3284), .ZN(n3293)
         );
  AOI22_X1 U4365 ( .A1(n3446), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3378), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3289) );
  AOI22_X1 U4366 ( .A1(n3462), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3463), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3288) );
  NAND4_X1 U4367 ( .A1(n3291), .A2(n3290), .A3(n3289), .A4(n3288), .ZN(n3292)
         );
  OR2_X2 U4368 ( .A1(n3293), .A2(n3292), .ZN(n4158) );
  NAND2_X2 U4369 ( .A1(n4274), .A2(n4158), .ZN(n4381) );
  AOI22_X1 U4370 ( .A1(n3360), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4371 ( .A1(n3991), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3108), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3297) );
  AOI22_X1 U4372 ( .A1(n3462), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3463), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3296) );
  AOI22_X1 U4373 ( .A1(n3509), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3295) );
  AOI22_X1 U4374 ( .A1(n4033), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3303) );
  AOI22_X1 U4375 ( .A1(n4055), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3302) );
  AOI22_X1 U4376 ( .A1(n3379), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3301) );
  INV_X2 U4378 ( .A(n3410), .ZN(n3403) );
  AOI22_X1 U4379 ( .A1(n3446), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3378), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3308) );
  AOI22_X1 U4380 ( .A1(n3462), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3463), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3307) );
  AND4_X2 U4381 ( .A1(n3310), .A2(n3309), .A3(n3308), .A4(n3307), .ZN(n3316)
         );
  AOI22_X1 U4382 ( .A1(n3991), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4383 ( .A1(n4033), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3112), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4384 ( .A1(n4055), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3312) );
  NAND2_X1 U4385 ( .A1(n3996), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3321)
         );
  NAND2_X1 U4386 ( .A1(n3360), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3320) );
  INV_X1 U4387 ( .A(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3317) );
  NAND2_X1 U4388 ( .A1(n4040), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3318)
         );
  NAND2_X1 U4389 ( .A1(n3446), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3325) );
  NAND2_X1 U4390 ( .A1(n3462), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3324) );
  NAND2_X1 U4391 ( .A1(n3463), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3323) );
  NAND2_X1 U4392 ( .A1(n3378), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3322)
         );
  NAND2_X1 U4393 ( .A1(n3991), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3331) );
  NAND2_X1 U4394 ( .A1(n4033), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3330) );
  NAND2_X1 U4395 ( .A1(n4039), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3329) );
  INV_X1 U4396 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3327) );
  NAND2_X1 U4397 ( .A1(n3447), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3335)
         );
  NAND2_X1 U4398 ( .A1(n4055), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3334)
         );
  NAND2_X1 U4399 ( .A1(n3509), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3333) );
  NAND2_X1 U4400 ( .A1(n3294), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3332) );
  NAND2_X1 U4401 ( .A1(n4453), .A2(n3445), .ZN(n3395) );
  AOI22_X1 U4402 ( .A1(n3360), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3343) );
  AOI22_X1 U4403 ( .A1(n3462), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3463), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3342) );
  AOI22_X1 U4404 ( .A1(n3996), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3379), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3341) );
  NAND4_X1 U4405 ( .A1(n3344), .A2(n3343), .A3(n3342), .A4(n3341), .ZN(n3350)
         );
  AOI22_X1 U4406 ( .A1(n3991), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3348) );
  AOI22_X1 U4407 ( .A1(n4033), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3347) );
  AOI22_X1 U4408 ( .A1(n4055), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3346) );
  AOI22_X1 U4409 ( .A1(n3447), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3345) );
  NAND4_X1 U4410 ( .A1(n3348), .A2(n3347), .A3(n3346), .A4(n3345), .ZN(n3349)
         );
  NOR2_X2 U4411 ( .A1(n3395), .A2(n5374), .ZN(n4254) );
  NAND2_X1 U4412 ( .A1(n3351), .A2(n4254), .ZN(n4272) );
  INV_X1 U4413 ( .A(n4272), .ZN(n3376) );
  NAND2_X1 U4414 ( .A1(n4039), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3355) );
  NAND2_X1 U4415 ( .A1(n3991), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3354) );
  NAND2_X1 U4416 ( .A1(n3509), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3353) );
  NAND2_X1 U4417 ( .A1(n3294), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3352) );
  NAND2_X1 U4418 ( .A1(n3446), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3359) );
  NAND2_X1 U4419 ( .A1(n3996), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3358)
         );
  NAND2_X1 U4420 ( .A1(n3462), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3357) );
  NAND2_X1 U4421 ( .A1(n3463), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3356) );
  NAND2_X1 U4422 ( .A1(n3360), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3366) );
  INV_X1 U4423 ( .A(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3361) );
  NAND2_X1 U4424 ( .A1(n4040), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3364)
         );
  NAND2_X1 U4425 ( .A1(n3378), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3363)
         );
  NAND2_X1 U4426 ( .A1(n4033), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3371) );
  NAND2_X1 U4427 ( .A1(n4055), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3370)
         );
  NAND2_X1 U4428 ( .A1(n3447), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3369)
         );
  NAND2_X1 U4429 ( .A1(n3376), .A2(n4287), .ZN(n4281) );
  AOI22_X1 U4430 ( .A1(n3462), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3463), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3381) );
  AOI22_X1 U4431 ( .A1(n3996), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3379), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3380) );
  AOI22_X1 U4432 ( .A1(n3991), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3387) );
  AOI22_X1 U4433 ( .A1(n4033), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3386) );
  AOI22_X1 U4434 ( .A1(n4055), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3385) );
  AOI22_X1 U4435 ( .A1(n3447), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3384) );
  NAND2_X1 U4436 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), .ZN(
        n4551) );
  OAI21_X1 U4437 ( .B1(STATE_REG_2__SCAN_IN), .B2(STATE_REG_1__SCAN_IN), .A(
        n4551), .ZN(n4261) );
  NAND2_X2 U4438 ( .A1(n3111), .A2(n3412), .ZN(n3402) );
  NOR2_X1 U4439 ( .A1(n3403), .A2(n4158), .ZN(n3390) );
  NAND2_X1 U4440 ( .A1(n3396), .A2(n3585), .ZN(n4845) );
  NAND2_X1 U4441 ( .A1(n3395), .A2(n3394), .ZN(n3400) );
  NAND2_X1 U4442 ( .A1(n3397), .A2(n3634), .ZN(n3398) );
  OAI211_X1 U4443 ( .C1(n3634), .C2(n4274), .A(n3398), .B(n4453), .ZN(n3399)
         );
  NAND3_X1 U4444 ( .A1(n3401), .A2(n3400), .A3(n3399), .ZN(n3420) );
  INV_X1 U4445 ( .A(n3420), .ZN(n4258) );
  NOR2_X1 U4446 ( .A1(n3402), .A2(n3409), .ZN(n3404) );
  OAI211_X1 U4447 ( .C1(n4281), .C2(n3405), .A(n4378), .B(n4283), .ZN(n3406)
         );
  NAND2_X1 U4448 ( .A1(n3406), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3422) );
  INV_X1 U4449 ( .A(n3422), .ZN(n3408) );
  INV_X1 U4450 ( .A(n4147), .ZN(n3531) );
  INV_X1 U4451 ( .A(n4138), .ZN(n3530) );
  AOI22_X1 U4452 ( .A1(n3531), .A2(n6645), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n3530), .ZN(n3421) );
  INV_X1 U4453 ( .A(n3421), .ZN(n3407) );
  NAND2_X1 U4454 ( .A1(n3408), .A2(n3263), .ZN(n3500) );
  NAND2_X1 U4455 ( .A1(n3423), .A2(n3461), .ZN(n3416) );
  NAND2_X1 U4456 ( .A1(n3411), .A2(n3410), .ZN(n3415) );
  NAND2_X1 U4457 ( .A1(n3523), .A2(n4620), .ZN(n3414) );
  AND4_X2 U4458 ( .A1(n3426), .A2(n3416), .A3(n3415), .A4(n3414), .ZN(n3419)
         );
  INV_X1 U4459 ( .A(n4254), .ZN(n3417) );
  AND2_X2 U4460 ( .A1(n3110), .A2(n3102), .ZN(n4151) );
  AND2_X1 U4461 ( .A1(n4453), .A2(n3585), .ZN(n3418) );
  OAI211_X1 U4462 ( .C1(n3504), .C2(n3268), .A(n3422), .B(n3421), .ZN(n3502)
         );
  NAND2_X1 U4463 ( .A1(n3500), .A2(n3502), .ZN(n3444) );
  INV_X1 U4464 ( .A(n4151), .ZN(n3424) );
  INV_X1 U4465 ( .A(n3425), .ZN(n3430) );
  NAND2_X1 U4466 ( .A1(n4381), .A2(n4287), .ZN(n3429) );
  NOR2_X1 U4467 ( .A1(n3394), .A2(n4287), .ZN(n4621) );
  NAND2_X1 U4468 ( .A1(n3397), .A2(n3585), .ZN(n3789) );
  INV_X1 U4469 ( .A(n3789), .ZN(n3428) );
  NOR2_X1 U4470 ( .A1(n3396), .A2(n4158), .ZN(n3427) );
  NAND3_X1 U4471 ( .A1(n4621), .A2(n3428), .A3(n3427), .ZN(n4749) );
  NAND2_X1 U4472 ( .A1(n3788), .A2(n3397), .ZN(n3432) );
  NAND2_X1 U4473 ( .A1(n3432), .A2(n4287), .ZN(n3433) );
  OAI21_X1 U4474 ( .B1(n3431), .B2(n3433), .A(n4620), .ZN(n3435) );
  NAND4_X1 U4475 ( .A1(n3436), .A2(n3442), .A3(n3435), .A4(n3434), .ZN(n3476)
         );
  MUX2_X1 U4476 ( .A(n4147), .B(n4138), .S(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .Z(n3440) );
  NAND2_X1 U4477 ( .A1(n3438), .A2(n3437), .ZN(n3439) );
  XNOR2_X2 U4478 ( .A(n3444), .B(n3443), .ZN(n4786) );
  NAND2_X1 U4479 ( .A1(n4786), .A2(n4872), .ZN(n3460) );
  INV_X1 U4480 ( .A(n3534), .ZN(n3520) );
  AOI22_X1 U4481 ( .A1(n4032), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4482 ( .A1(n3446), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3450) );
  INV_X1 U4483 ( .A(n3447), .ZN(n3468) );
  AOI22_X1 U4484 ( .A1(n4034), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4485 ( .A1(n4056), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3448) );
  NAND4_X1 U4486 ( .A1(n3451), .A2(n3450), .A3(n3449), .A4(n3448), .ZN(n3458)
         );
  AOI22_X1 U4487 ( .A1(n4053), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3456) );
  AOI22_X1 U4488 ( .A1(n3996), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3455) );
  AOI22_X1 U4489 ( .A1(n4014), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4490 ( .A1(n3907), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3453) );
  NAND4_X1 U4491 ( .A1(n3456), .A2(n3455), .A3(n3454), .A4(n3453), .ZN(n3457)
         );
  NAND2_X1 U4492 ( .A1(n3520), .A2(n4150), .ZN(n3459) );
  AOI22_X1 U4493 ( .A1(n3101), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3467) );
  AOI22_X1 U4494 ( .A1(n4058), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3466) );
  AOI22_X1 U4495 ( .A1(n4056), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3464) );
  NAND4_X1 U4496 ( .A1(n3467), .A2(n3466), .A3(n3465), .A4(n3464), .ZN(n3474)
         );
  AOI22_X1 U4497 ( .A1(n4032), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4039), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3472) );
  AOI22_X1 U4498 ( .A1(n4053), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3471) );
  AOI22_X1 U4499 ( .A1(n4014), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3470) );
  INV_X2 U4500 ( .A(n3468), .ZN(n4034) );
  AOI22_X1 U4501 ( .A1(n4034), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3469) );
  NAND4_X1 U4502 ( .A1(n3472), .A2(n3471), .A3(n3470), .A4(n3469), .ZN(n3473)
         );
  NAND2_X1 U4503 ( .A1(n3523), .A2(n4150), .ZN(n3475) );
  NAND2_X1 U4504 ( .A1(n3622), .A2(n3621), .ZN(n3495) );
  INV_X1 U4505 ( .A(n3476), .ZN(n3477) );
  NAND2_X1 U4506 ( .A1(n3636), .A2(n4872), .ZN(n3628) );
  INV_X1 U4507 ( .A(n3479), .ZN(n3491) );
  NAND2_X1 U4508 ( .A1(n3445), .A2(n4222), .ZN(n3493) );
  AOI22_X1 U4509 ( .A1(n4053), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4032), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3483) );
  AOI22_X1 U4510 ( .A1(n4034), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3482) );
  AOI22_X1 U4511 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n3996), .B1(n4041), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3481) );
  AOI22_X1 U4512 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n3446), .B1(n3907), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3480) );
  NAND4_X1 U4513 ( .A1(n3483), .A2(n3482), .A3(n3481), .A4(n3480), .ZN(n3489)
         );
  AOI22_X1 U4514 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n4014), .B1(n4054), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3487) );
  AOI22_X1 U4515 ( .A1(n3118), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3486) );
  AOI22_X1 U4516 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n4058), .B1(n4057), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3485) );
  AOI22_X1 U4517 ( .A1(n4056), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3973), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3484) );
  NAND4_X1 U4518 ( .A1(n3487), .A2(n3486), .A3(n3485), .A4(n3484), .ZN(n3488)
         );
  INV_X1 U4519 ( .A(n4159), .ZN(n3490) );
  AOI21_X1 U4520 ( .B1(n4925), .B2(n4159), .A(n4872), .ZN(n3494) );
  NAND2_X1 U4521 ( .A1(n3495), .A2(n3620), .ZN(n3499) );
  INV_X1 U4522 ( .A(n3622), .ZN(n3497) );
  INV_X1 U4523 ( .A(n3621), .ZN(n3496) );
  NAND2_X1 U4524 ( .A1(n3497), .A2(n3496), .ZN(n3498) );
  NAND2_X1 U4525 ( .A1(n3499), .A2(n3498), .ZN(n3610) );
  NAND2_X1 U4526 ( .A1(n3501), .A2(n3500), .ZN(n3503) );
  NAND2_X1 U4527 ( .A1(n6456), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3507) );
  NAND2_X1 U4528 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3505) );
  NAND2_X1 U4529 ( .A1(n3505), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3506) );
  NAND2_X1 U4530 ( .A1(n3507), .A2(n3506), .ZN(n5076) );
  AOI22_X1 U4531 ( .A1(n5076), .A2(n3531), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3530), .ZN(n3508) );
  NAND2_X1 U4532 ( .A1(n4660), .A2(n4872), .ZN(n3522) );
  AOI22_X1 U4533 ( .A1(n4032), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3513) );
  AOI22_X1 U4534 ( .A1(n4053), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3512) );
  AOI22_X1 U4535 ( .A1(n4014), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3511) );
  AOI22_X1 U4536 ( .A1(n4034), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3510) );
  NAND4_X1 U4537 ( .A1(n3513), .A2(n3512), .A3(n3511), .A4(n3510), .ZN(n3519)
         );
  AOI22_X1 U4538 ( .A1(n3996), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3517) );
  AOI22_X1 U4539 ( .A1(n4058), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3516) );
  AOI22_X1 U4540 ( .A1(n3446), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3515) );
  AOI22_X1 U4541 ( .A1(n4056), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3973), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3514) );
  NAND4_X1 U4542 ( .A1(n3517), .A2(n3516), .A3(n3515), .A4(n3514), .ZN(n3518)
         );
  NAND2_X1 U4543 ( .A1(n3520), .A2(n4174), .ZN(n3521) );
  AOI22_X1 U4544 ( .A1(n3523), .A2(n4174), .B1(n3461), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3524) );
  NAND2_X1 U4545 ( .A1(n6526), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6550) );
  NAND2_X1 U4546 ( .A1(n6550), .A2(n6781), .ZN(n3529) );
  AOI22_X1 U4547 ( .A1(n6563), .A2(n3531), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3530), .ZN(n3532) );
  NAND2_X1 U4548 ( .A1(n4742), .A2(n4872), .ZN(n3546) );
  AOI22_X1 U4549 ( .A1(n4053), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3538) );
  AOI22_X1 U4550 ( .A1(n4041), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4551 ( .A1(n4056), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3973), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3536) );
  AOI22_X1 U4552 ( .A1(n3446), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3535) );
  NAND4_X1 U4553 ( .A1(n3538), .A2(n3537), .A3(n3536), .A4(n3535), .ZN(n3544)
         );
  AOI22_X1 U4554 ( .A1(n4014), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3996), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3542) );
  AOI22_X1 U4555 ( .A1(n4032), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4556 ( .A1(n3452), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4557 ( .A1(n4058), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3539) );
  NAND4_X1 U4558 ( .A1(n3542), .A2(n3541), .A3(n3540), .A4(n3539), .ZN(n3543)
         );
  AOI22_X1 U4559 ( .A1(n4127), .A2(n4184), .B1(INSTQUEUE_REG_0__3__SCAN_IN), 
        .B2(n3461), .ZN(n3545) );
  AOI22_X1 U4560 ( .A1(n4032), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3550) );
  AOI22_X1 U4561 ( .A1(n4053), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3549) );
  AOI22_X1 U4562 ( .A1(n4014), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3548) );
  AOI22_X1 U4563 ( .A1(n4034), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3547) );
  NAND4_X1 U4564 ( .A1(n3550), .A2(n3549), .A3(n3548), .A4(n3547), .ZN(n3556)
         );
  INV_X1 U4565 ( .A(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n6770) );
  AOI22_X1 U4566 ( .A1(n3101), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4567 ( .A1(n4058), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3553) );
  AOI22_X1 U4568 ( .A1(n3446), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3552) );
  AOI22_X1 U4569 ( .A1(n4056), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3973), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3551) );
  NAND4_X1 U4570 ( .A1(n3554), .A2(n3553), .A3(n3552), .A4(n3551), .ZN(n3555)
         );
  NAND2_X1 U4571 ( .A1(n4127), .A2(n4191), .ZN(n3558) );
  NAND2_X1 U4572 ( .A1(n3461), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3557) );
  AOI22_X1 U4573 ( .A1(n4034), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4574 ( .A1(n4014), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4575 ( .A1(n3101), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3560) );
  AOI22_X1 U4576 ( .A1(n4058), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3973), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3559) );
  NAND4_X1 U4577 ( .A1(n3562), .A2(n3561), .A3(n3560), .A4(n3559), .ZN(n3568)
         );
  AOI22_X1 U4578 ( .A1(n4053), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4032), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3566) );
  AOI22_X1 U4579 ( .A1(n3452), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4580 ( .A1(n4056), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4581 ( .A1(n4019), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3563) );
  NAND4_X1 U4582 ( .A1(n3566), .A2(n3565), .A3(n3564), .A4(n3563), .ZN(n3567)
         );
  NAND2_X1 U4583 ( .A1(n4127), .A2(n4202), .ZN(n3570) );
  NAND2_X1 U4584 ( .A1(n3461), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3569) );
  NAND2_X1 U4585 ( .A1(n3570), .A2(n3569), .ZN(n3647) );
  AOI22_X1 U4586 ( .A1(n4032), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3575) );
  AOI22_X1 U4587 ( .A1(n4053), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3574) );
  AOI22_X1 U4588 ( .A1(n4014), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3573) );
  AOI22_X1 U4589 ( .A1(n4034), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3572) );
  NAND4_X1 U4590 ( .A1(n3575), .A2(n3574), .A3(n3573), .A4(n3572), .ZN(n3581)
         );
  AOI22_X1 U4591 ( .A1(n3996), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3579) );
  AOI22_X1 U4592 ( .A1(n4058), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3578) );
  AOI22_X1 U4593 ( .A1(n3446), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3577) );
  AOI22_X1 U4594 ( .A1(n4056), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3973), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3576) );
  NAND4_X1 U4595 ( .A1(n3579), .A2(n3578), .A3(n3577), .A4(n3576), .ZN(n3580)
         );
  AOI22_X1 U4596 ( .A1(n4127), .A2(n4211), .B1(n3461), .B2(
        INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3653) );
  INV_X1 U4597 ( .A(n3653), .ZN(n3582) );
  INV_X1 U4598 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5086) );
  NAND2_X1 U4599 ( .A1(n4127), .A2(n4222), .ZN(n3583) );
  OAI21_X1 U4600 ( .B1(n5086), .B2(n4122), .A(n3583), .ZN(n3584) );
  NAND2_X1 U4601 ( .A1(n4208), .A2(n3778), .ZN(n3590) );
  AND2_X1 U4602 ( .A1(n3658), .A2(n6847), .ZN(n3586) );
  OR2_X1 U4603 ( .A1(n3586), .A2(n3685), .ZN(n6192) );
  NAND2_X1 U4604 ( .A1(n6192), .A2(n4502), .ZN(n3587) );
  OAI21_X1 U4605 ( .B1(n6847), .B2(n3801), .A(n3587), .ZN(n3588) );
  AOI21_X1 U4606 ( .B1(n3833), .B2(EAX_REG_7__SCAN_IN), .A(n3588), .ZN(n3589)
         );
  NAND2_X1 U4607 ( .A1(n3590), .A2(n3589), .ZN(n5067) );
  INV_X1 U4608 ( .A(n3649), .ZN(n3595) );
  INV_X1 U4609 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3593) );
  INV_X1 U4610 ( .A(n3592), .ZN(n3603) );
  NAND2_X1 U4611 ( .A1(n3593), .A2(n3603), .ZN(n3594) );
  NAND2_X1 U4612 ( .A1(n3595), .A2(n3594), .ZN(n6353) );
  NAND2_X1 U4613 ( .A1(n3392), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3613) );
  OAI21_X1 U4614 ( .B1(n6129), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6603), 
        .ZN(n3597) );
  NAND2_X1 U4615 ( .A1(n4080), .A2(EAX_REG_4__SCAN_IN), .ZN(n3596) );
  OAI211_X1 U4616 ( .C1(n3613), .C2(n4634), .A(n3597), .B(n3596), .ZN(n3598)
         );
  OAI21_X1 U4617 ( .B1(n4028), .B2(n6353), .A(n3598), .ZN(n3599) );
  NAND2_X1 U4618 ( .A1(n3600), .A2(n3599), .ZN(n4853) );
  XNOR2_X2 U4619 ( .A(n3602), .B(n3601), .ZN(n5027) );
  NAND2_X1 U4620 ( .A1(n5027), .A2(n3778), .ZN(n3609) );
  INV_X1 U4621 ( .A(n3614), .ZN(n3604) );
  OAI21_X1 U4622 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3604), .A(n3603), 
        .ZN(n5624) );
  AOI22_X1 U4623 ( .A1(n4502), .A2(n5624), .B1(n4079), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3606) );
  NAND2_X1 U4624 ( .A1(n3833), .A2(EAX_REG_3__SCAN_IN), .ZN(n3605) );
  OAI211_X1 U4625 ( .C1(n3613), .C2(n3246), .A(n3606), .B(n3605), .ZN(n3607)
         );
  INV_X1 U4626 ( .A(n3607), .ZN(n3608) );
  NAND2_X1 U4627 ( .A1(n3609), .A2(n3608), .ZN(n4852) );
  XNOR2_X1 U4628 ( .A(n3611), .B(n3610), .ZN(n4167) );
  NAND2_X1 U4629 ( .A1(n4167), .A2(n3778), .ZN(n3612) );
  INV_X1 U4630 ( .A(n3613), .ZN(n3637) );
  NAND2_X1 U4631 ( .A1(n3637), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3619) );
  INV_X1 U4632 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3616) );
  OAI21_X1 U4633 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3614), .ZN(n6362) );
  NAND2_X1 U4634 ( .A1(n4502), .A2(n6362), .ZN(n3615) );
  OAI21_X1 U4635 ( .B1(n3801), .B2(n3616), .A(n3615), .ZN(n3617) );
  AOI21_X1 U4636 ( .B1(n4080), .B2(EAX_REG_2__SCAN_IN), .A(n3617), .ZN(n3618)
         );
  NAND2_X1 U4637 ( .A1(n3619), .A2(n3618), .ZN(n4826) );
  NAND2_X1 U4638 ( .A1(n4827), .A2(n4826), .ZN(n3643) );
  NAND2_X1 U4639 ( .A1(n4887), .A2(n3778), .ZN(n3627) );
  AOI22_X1 U4640 ( .A1(n4080), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6603), .ZN(n3625) );
  NAND2_X1 U4641 ( .A1(n3637), .A2(n6756), .ZN(n3624) );
  AND2_X1 U4642 ( .A1(n3625), .A2(n3624), .ZN(n3626) );
  NAND2_X1 U4643 ( .A1(n3492), .A2(n3631), .ZN(n3632) );
  AND2_X1 U4644 ( .A1(n3634), .A2(n3585), .ZN(n3635) );
  AOI21_X1 U4645 ( .B1(n4157), .B2(n3635), .A(n6603), .ZN(n4701) );
  NAND2_X1 U4646 ( .A1(n3114), .A2(n3778), .ZN(n3641) );
  AOI22_X1 U4647 ( .A1(n4080), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6603), .ZN(n3639) );
  NAND2_X1 U4648 ( .A1(n3637), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3638) );
  AND2_X1 U4649 ( .A1(n3639), .A2(n3638), .ZN(n3640) );
  NAND2_X1 U4650 ( .A1(n3641), .A2(n3640), .ZN(n4700) );
  NAND2_X1 U4651 ( .A1(n4701), .A2(n4700), .ZN(n4703) );
  OR2_X1 U4652 ( .A1(n4700), .A2(n4028), .ZN(n3642) );
  NAND2_X1 U4653 ( .A1(n4703), .A2(n3642), .ZN(n4734) );
  NAND2_X1 U4654 ( .A1(n4735), .A2(n4734), .ZN(n4733) );
  NAND2_X1 U4655 ( .A1(n3643), .A2(n4733), .ZN(n3646) );
  XNOR2_X1 U4656 ( .A(n3648), .B(n3647), .ZN(n4190) );
  NOR2_X1 U4657 ( .A1(n3649), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3650)
         );
  NOR2_X1 U4658 ( .A1(n3655), .A2(n3650), .ZN(n6212) );
  INV_X1 U4659 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6960) );
  OAI22_X1 U4660 ( .A1(n6212), .A2(n4028), .B1(n3801), .B2(n6960), .ZN(n3651)
         );
  AOI21_X1 U4661 ( .B1(n3833), .B2(EAX_REG_5__SCAN_IN), .A(n3651), .ZN(n3652)
         );
  NAND2_X1 U4662 ( .A1(n3654), .A2(n3653), .ZN(n4200) );
  INV_X1 U4663 ( .A(n3655), .ZN(n3656) );
  INV_X1 U4664 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6199) );
  NAND2_X1 U4665 ( .A1(n3656), .A2(n6199), .ZN(n3657) );
  NAND2_X1 U4666 ( .A1(n3658), .A2(n3657), .ZN(n6343) );
  INV_X1 U4667 ( .A(EAX_REG_6__SCAN_IN), .ZN(n5066) );
  OAI22_X1 U4668 ( .A1(n3659), .A2(n5066), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6199), .ZN(n3660) );
  MUX2_X1 U4669 ( .A(n6343), .B(n3660), .S(n4028), .Z(n3661) );
  AOI21_X1 U4670 ( .B1(n4200), .B2(n3778), .A(n3661), .ZN(n5025) );
  AOI22_X1 U4671 ( .A1(n4053), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3665) );
  AOI22_X1 U4672 ( .A1(n4014), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3664) );
  AOI22_X1 U4673 ( .A1(n4034), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4674 ( .A1(n3907), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3973), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3662) );
  NAND4_X1 U4675 ( .A1(n3665), .A2(n3664), .A3(n3663), .A4(n3662), .ZN(n3671)
         );
  AOI22_X1 U4676 ( .A1(n4056), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4677 ( .A1(n4032), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4678 ( .A1(n4041), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4679 ( .A1(n4019), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3666) );
  NAND4_X1 U4680 ( .A1(n3669), .A2(n3668), .A3(n3667), .A4(n3666), .ZN(n3670)
         );
  NOR2_X1 U4681 ( .A1(n3671), .A2(n3670), .ZN(n3674) );
  INV_X1 U4682 ( .A(n3778), .ZN(n3769) );
  XNOR2_X1 U4683 ( .A(n3705), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5875)
         );
  NAND2_X1 U4684 ( .A1(n5875), .A2(n4502), .ZN(n3673) );
  AOI22_X1 U4685 ( .A1(n4080), .A2(EAX_REG_10__SCAN_IN), .B1(n4079), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3672) );
  OAI211_X1 U4686 ( .C1(n3674), .C2(n3769), .A(n3673), .B(n3672), .ZN(n5152)
         );
  AOI22_X1 U4687 ( .A1(n4014), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3678) );
  AOI22_X1 U4688 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n4019), .B1(n4058), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3677) );
  AOI22_X1 U4689 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n3117), .B1(n4041), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3676) );
  AOI22_X1 U4690 ( .A1(n3116), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3675) );
  NAND4_X1 U4691 ( .A1(n3678), .A2(n3677), .A3(n3676), .A4(n3675), .ZN(n3684)
         );
  AOI22_X1 U4692 ( .A1(n4053), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3682) );
  AOI22_X1 U4693 ( .A1(n4032), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3681) );
  AOI22_X1 U4694 ( .A1(n4056), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3973), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3680) );
  AOI22_X1 U4695 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n3907), .B1(n4057), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3679) );
  NAND4_X1 U4696 ( .A1(n3682), .A2(n3681), .A3(n3680), .A4(n3679), .ZN(n3683)
         );
  OAI21_X1 U4697 ( .B1(n3684), .B2(n3683), .A(n3778), .ZN(n3689) );
  NAND2_X1 U4698 ( .A1(n4080), .A2(EAX_REG_8__SCAN_IN), .ZN(n3688) );
  XNOR2_X1 U4699 ( .A(n3685), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U4700 ( .A1(n6174), .A2(n4502), .ZN(n3687) );
  NAND2_X1 U4701 ( .A1(n4079), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3686)
         );
  NAND4_X1 U4702 ( .A1(n3689), .A2(n3688), .A3(n3687), .A4(n3686), .ZN(n5196)
         );
  XOR2_X1 U4703 ( .A(n6159), .B(n3690), .Z(n6162) );
  AOI22_X1 U4704 ( .A1(n4053), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3694) );
  AOI22_X1 U4705 ( .A1(n3117), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3693) );
  AOI22_X1 U4706 ( .A1(n4041), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3973), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3692) );
  AOI22_X1 U4707 ( .A1(n4058), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3691) );
  NAND4_X1 U4708 ( .A1(n3694), .A2(n3693), .A3(n3692), .A4(n3691), .ZN(n3700)
         );
  AOI22_X1 U4709 ( .A1(n4014), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4056), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3698) );
  AOI22_X1 U4710 ( .A1(n4032), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3697) );
  AOI22_X1 U4711 ( .A1(n3452), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3696) );
  AOI22_X1 U4712 ( .A1(n4019), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3695) );
  NAND4_X1 U4713 ( .A1(n3698), .A2(n3697), .A3(n3696), .A4(n3695), .ZN(n3699)
         );
  OAI21_X1 U4714 ( .B1(n3700), .B2(n3699), .A(n3778), .ZN(n3703) );
  NAND2_X1 U4715 ( .A1(n4080), .A2(EAX_REG_9__SCAN_IN), .ZN(n3702) );
  NAND2_X1 U4716 ( .A1(n4079), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3701)
         );
  OAI21_X1 U4717 ( .B1(n6162), .B2(n4028), .A(n3265), .ZN(n5194) );
  AND3_X1 U4718 ( .A1(n5152), .A2(n5196), .A3(n5194), .ZN(n3704) );
  AOI21_X1 U4719 ( .B1(n7047), .B2(n3706), .A(n3138), .ZN(n6329) );
  OR2_X1 U4720 ( .A1(n6329), .A2(n4028), .ZN(n3721) );
  AOI22_X1 U4721 ( .A1(n4032), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3710) );
  AOI22_X1 U4722 ( .A1(n4053), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4014), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3709) );
  AOI22_X1 U4723 ( .A1(n4056), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3708) );
  AOI22_X1 U4724 ( .A1(n4058), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3707) );
  NAND4_X1 U4725 ( .A1(n3710), .A2(n3709), .A3(n3708), .A4(n3707), .ZN(n3716)
         );
  AOI22_X1 U4726 ( .A1(n4034), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3714) );
  AOI22_X1 U4727 ( .A1(n3452), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3713) );
  AOI22_X1 U4728 ( .A1(n4019), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3712) );
  AOI22_X1 U4729 ( .A1(n3117), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3973), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3711) );
  NAND4_X1 U4730 ( .A1(n3714), .A2(n3713), .A3(n3712), .A4(n3711), .ZN(n3715)
         );
  OAI21_X1 U4731 ( .B1(n3716), .B2(n3715), .A(n3778), .ZN(n3719) );
  NAND2_X1 U4732 ( .A1(n4080), .A2(EAX_REG_11__SCAN_IN), .ZN(n3718) );
  NAND2_X1 U4733 ( .A1(n4079), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3717)
         );
  AND3_X1 U4734 ( .A1(n3719), .A2(n3718), .A3(n3717), .ZN(n3720) );
  XNOR2_X1 U4735 ( .A(n3138), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5870)
         );
  AOI22_X1 U4736 ( .A1(n4053), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4032), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3725) );
  AOI22_X1 U4737 ( .A1(n4034), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4738 ( .A1(n4054), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3973), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4739 ( .A1(n4058), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3722) );
  NAND4_X1 U4740 ( .A1(n3725), .A2(n3724), .A3(n3723), .A4(n3722), .ZN(n3731)
         );
  AOI22_X1 U4741 ( .A1(n4014), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3729) );
  AOI22_X1 U4742 ( .A1(n4056), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3728) );
  AOI22_X1 U4743 ( .A1(n3118), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3727) );
  AOI22_X1 U4744 ( .A1(n4019), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3726) );
  NAND4_X1 U4745 ( .A1(n3729), .A2(n3728), .A3(n3727), .A4(n3726), .ZN(n3730)
         );
  OAI21_X1 U4746 ( .B1(n3731), .B2(n3730), .A(n3778), .ZN(n3734) );
  NAND2_X1 U4747 ( .A1(n3833), .A2(EAX_REG_12__SCAN_IN), .ZN(n3733) );
  NAND2_X1 U4748 ( .A1(n4079), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3732)
         );
  NAND3_X1 U4749 ( .A1(n3734), .A2(n3733), .A3(n3732), .ZN(n3735) );
  NAND2_X1 U4750 ( .A1(n3833), .A2(EAX_REG_13__SCAN_IN), .ZN(n3738) );
  OAI21_X1 U4751 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3736), .A(n3764), 
        .ZN(n6157) );
  AOI22_X1 U4752 ( .A1(n4502), .A2(n6157), .B1(n4079), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3737) );
  NAND2_X1 U4753 ( .A1(n3738), .A2(n3737), .ZN(n3739) );
  AOI22_X1 U4754 ( .A1(n4032), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3744) );
  AOI22_X1 U4755 ( .A1(n4053), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3743) );
  AOI22_X1 U4756 ( .A1(n3117), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3742) );
  AOI22_X1 U4757 ( .A1(n4058), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3741) );
  NAND4_X1 U4758 ( .A1(n3744), .A2(n3743), .A3(n3742), .A4(n3741), .ZN(n3750)
         );
  AOI22_X1 U4759 ( .A1(n4014), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4760 ( .A1(n3112), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4761 ( .A1(n4056), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3746) );
  AOI22_X1 U4762 ( .A1(n4019), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3745) );
  NAND4_X1 U4763 ( .A1(n3748), .A2(n3747), .A3(n3746), .A4(n3745), .ZN(n3749)
         );
  OR2_X1 U4764 ( .A1(n3750), .A2(n3749), .ZN(n3751) );
  NAND2_X1 U4765 ( .A1(n3778), .A2(n3751), .ZN(n5664) );
  AOI22_X1 U4766 ( .A1(n4014), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4767 ( .A1(n4056), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4768 ( .A1(n3116), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3754) );
  AOI22_X1 U4769 ( .A1(n4041), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3753) );
  NAND4_X1 U4770 ( .A1(n3756), .A2(n3755), .A3(n3754), .A4(n3753), .ZN(n3762)
         );
  AOI22_X1 U4771 ( .A1(n4032), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4772 ( .A1(n4053), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3759) );
  AOI22_X1 U4773 ( .A1(n4034), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3758) );
  AOI22_X1 U4774 ( .A1(n4019), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3757) );
  NAND4_X1 U4775 ( .A1(n3760), .A2(n3759), .A3(n3758), .A4(n3757), .ZN(n3761)
         );
  NOR2_X1 U4776 ( .A1(n3762), .A2(n3761), .ZN(n3768) );
  INV_X1 U4777 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6811) );
  NAND2_X1 U4778 ( .A1(n3764), .A2(n6811), .ZN(n3765) );
  NAND2_X1 U4779 ( .A1(n3783), .A2(n3765), .ZN(n5851) );
  AOI22_X1 U4780 ( .A1(n5851), .A2(n4502), .B1(PHYADDRPOINTER_REG_14__SCAN_IN), 
        .B2(n4079), .ZN(n3767) );
  NAND2_X1 U4781 ( .A1(n3833), .A2(EAX_REG_14__SCAN_IN), .ZN(n3766) );
  OAI211_X1 U4782 ( .C1(n3769), .C2(n3768), .A(n3767), .B(n3766), .ZN(n5582)
         );
  AOI22_X1 U4783 ( .A1(n4056), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4784 ( .A1(n4032), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4785 ( .A1(n4034), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4786 ( .A1(n4019), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3770) );
  NAND4_X1 U4787 ( .A1(n3773), .A2(n3772), .A3(n3771), .A4(n3770), .ZN(n3780)
         );
  AOI22_X1 U4788 ( .A1(n4014), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4789 ( .A1(n4053), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4790 ( .A1(n4054), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4791 ( .A1(n4041), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3774) );
  NAND4_X1 U4792 ( .A1(n3777), .A2(n3776), .A3(n3775), .A4(n3774), .ZN(n3779)
         );
  OAI21_X1 U4793 ( .B1(n3780), .B2(n3779), .A(n3778), .ZN(n3787) );
  NAND2_X1 U4794 ( .A1(n3833), .A2(EAX_REG_15__SCAN_IN), .ZN(n3786) );
  INV_X1 U4795 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3782) );
  NAND2_X1 U4796 ( .A1(n3783), .A2(n3782), .ZN(n3784) );
  NAND2_X1 U4797 ( .A1(n3818), .A2(n3784), .ZN(n5842) );
  AOI22_X1 U4798 ( .A1(n5842), .A2(n4502), .B1(PHYADDRPOINTER_REG_15__SCAN_IN), 
        .B2(n4079), .ZN(n3785) );
  AOI22_X1 U4799 ( .A1(n4053), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4800 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n4034), .B1(n3452), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4801 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n3117), .B1(n4054), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4802 ( .A1(n4019), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3790) );
  NAND4_X1 U4803 ( .A1(n3793), .A2(n3792), .A3(n3791), .A4(n3790), .ZN(n3799)
         );
  AOI22_X1 U4804 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n4056), .B1(n4058), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4805 ( .A1(n4014), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4806 ( .A1(n3118), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4807 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n3907), .B1(n4057), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3794) );
  NAND4_X1 U4808 ( .A1(n3797), .A2(n3796), .A3(n3795), .A4(n3794), .ZN(n3798)
         );
  OR2_X1 U4809 ( .A1(n3799), .A2(n3798), .ZN(n3800) );
  NAND2_X1 U4810 ( .A1(n4050), .A2(n3800), .ZN(n3804) );
  XNOR2_X1 U4811 ( .A(n3818), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5838)
         );
  INV_X1 U4812 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5834) );
  OAI22_X1 U4813 ( .A1(n5838), .A2(n4028), .B1(n5834), .B2(n3801), .ZN(n3802)
         );
  AOI21_X1 U4814 ( .B1(n3833), .B2(EAX_REG_16__SCAN_IN), .A(n3802), .ZN(n3803)
         );
  NAND2_X1 U4815 ( .A1(n3804), .A2(n3803), .ZN(n5551) );
  AOI22_X1 U4816 ( .A1(n4032), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4817 ( .A1(n4053), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4818 ( .A1(n4014), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4819 ( .A1(n4034), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3805) );
  NAND4_X1 U4820 ( .A1(n3808), .A2(n3807), .A3(n3806), .A4(n3805), .ZN(n3814)
         );
  AOI22_X1 U4821 ( .A1(n3117), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4822 ( .A1(n4058), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4823 ( .A1(n4019), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4824 ( .A1(n4056), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3809) );
  NAND4_X1 U4825 ( .A1(n3812), .A2(n3811), .A3(n3810), .A4(n3809), .ZN(n3813)
         );
  NOR2_X1 U4826 ( .A1(n3814), .A2(n3813), .ZN(n3817) );
  AOI21_X1 U4827 ( .B1(n5828), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3815) );
  AOI21_X1 U4828 ( .B1(n3833), .B2(EAX_REG_17__SCAN_IN), .A(n3815), .ZN(n3816)
         );
  OAI21_X1 U4829 ( .B1(n4074), .B2(n3817), .A(n3816), .ZN(n3820) );
  XNOR2_X1 U4830 ( .A(n3821), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5826)
         );
  NAND2_X1 U4831 ( .A1(n5826), .A2(n4502), .ZN(n3819) );
  NAND2_X1 U4832 ( .A1(n3820), .A2(n3819), .ZN(n5537) );
  OAI21_X1 U4833 ( .B1(n3821), .B2(n5828), .A(n5817), .ZN(n3822) );
  AND2_X1 U4834 ( .A1(n3822), .A2(n3852), .ZN(n5819) );
  AOI22_X1 U4835 ( .A1(n4032), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4836 ( .A1(n3117), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4837 ( .A1(n3509), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4838 ( .A1(n4056), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3823) );
  NAND4_X1 U4839 ( .A1(n3826), .A2(n3825), .A3(n3824), .A4(n3823), .ZN(n3832)
         );
  AOI22_X1 U4840 ( .A1(n4014), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3830) );
  AOI22_X1 U4841 ( .A1(n4053), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4842 ( .A1(n4058), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4843 ( .A1(n4019), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3827) );
  NAND4_X1 U4844 ( .A1(n3830), .A2(n3829), .A3(n3828), .A4(n3827), .ZN(n3831)
         );
  OR2_X1 U4845 ( .A1(n3832), .A2(n3831), .ZN(n3835) );
  INV_X1 U4846 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4638) );
  OAI22_X1 U4847 ( .A1(n3659), .A2(n4638), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5817), .ZN(n3834) );
  AOI21_X1 U4848 ( .B1(n4050), .B2(n3835), .A(n3834), .ZN(n3836) );
  MUX2_X1 U4849 ( .A(n5819), .B(n3836), .S(n4028), .Z(n5525) );
  NAND2_X1 U4850 ( .A1(n3838), .A2(n3837), .ZN(n5506) );
  AOI22_X1 U4851 ( .A1(n4032), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4852 ( .A1(n4053), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4853 ( .A1(n4014), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4854 ( .A1(n4034), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3839) );
  NAND4_X1 U4855 ( .A1(n3842), .A2(n3841), .A3(n3840), .A4(n3839), .ZN(n3848)
         );
  AOI22_X1 U4856 ( .A1(n3117), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4857 ( .A1(n4058), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4858 ( .A1(n4019), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4859 ( .A1(n4056), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3843) );
  NAND4_X1 U4860 ( .A1(n3846), .A2(n3845), .A3(n3844), .A4(n3843), .ZN(n3847)
         );
  NOR2_X1 U4861 ( .A1(n3848), .A2(n3847), .ZN(n3851) );
  AOI21_X1 U4862 ( .B1(n7008), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3849) );
  AOI21_X1 U4863 ( .B1(n3833), .B2(EAX_REG_19__SCAN_IN), .A(n3849), .ZN(n3850)
         );
  OAI21_X1 U4864 ( .B1(n4074), .B2(n3851), .A(n3850), .ZN(n3856) );
  NAND2_X1 U4865 ( .A1(n3852), .A2(n7008), .ZN(n3853) );
  NAND2_X1 U4866 ( .A1(n3870), .A2(n3853), .ZN(n5810) );
  INV_X1 U4867 ( .A(n5810), .ZN(n3854) );
  NAND2_X1 U4868 ( .A1(n3854), .A2(n4502), .ZN(n3855) );
  NAND2_X1 U4869 ( .A1(n3856), .A2(n3855), .ZN(n5508) );
  AOI22_X1 U4870 ( .A1(n4032), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4871 ( .A1(n3117), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4872 ( .A1(n4054), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4873 ( .A1(n4019), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3857) );
  NAND4_X1 U4874 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(n3866)
         );
  AOI22_X1 U4875 ( .A1(n4014), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4034), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4876 ( .A1(n4053), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4877 ( .A1(n4056), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4878 ( .A1(n4058), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3861) );
  NAND4_X1 U4879 ( .A1(n3864), .A2(n3863), .A3(n3862), .A4(n3861), .ZN(n3865)
         );
  NOR2_X1 U4880 ( .A1(n3866), .A2(n3865), .ZN(n3868) );
  AOI22_X1 U4881 ( .A1(n4080), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6603), .ZN(n3867) );
  OAI21_X1 U4882 ( .B1(n4074), .B2(n3868), .A(n3867), .ZN(n3872) );
  NAND2_X1 U4883 ( .A1(n3870), .A2(n3187), .ZN(n3871) );
  NAND2_X1 U4884 ( .A1(n3873), .A2(n3871), .ZN(n5803) );
  MUX2_X1 U4885 ( .A(n3872), .B(n5803), .S(n4502), .Z(n5491) );
  NAND2_X1 U4886 ( .A1(n3873), .A2(n6983), .ZN(n3874) );
  NAND2_X1 U4887 ( .A1(n3900), .A2(n3874), .ZN(n5797) );
  AOI22_X1 U4888 ( .A1(n4053), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4032), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4889 ( .A1(n4014), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4890 ( .A1(n3116), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4891 ( .A1(n4058), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3875) );
  NAND4_X1 U4892 ( .A1(n3878), .A2(n3877), .A3(n3876), .A4(n3875), .ZN(n3884)
         );
  AOI22_X1 U4893 ( .A1(n4034), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4894 ( .A1(n3118), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4895 ( .A1(n4019), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4896 ( .A1(n4056), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3879) );
  NAND4_X1 U4897 ( .A1(n3882), .A2(n3881), .A3(n3880), .A4(n3879), .ZN(n3883)
         );
  NOR2_X1 U4898 ( .A1(n3884), .A2(n3883), .ZN(n3886) );
  AOI22_X1 U4899 ( .A1(n4080), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6603), .ZN(n3885) );
  OAI21_X1 U4900 ( .B1(n4074), .B2(n3886), .A(n3885), .ZN(n3887) );
  MUX2_X1 U4901 ( .A(n5797), .B(n3887), .S(n4028), .Z(n5480) );
  AOI22_X1 U4902 ( .A1(n4053), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4903 ( .A1(n4055), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4904 ( .A1(n3117), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3973), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4905 ( .A1(n4056), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3888) );
  NAND4_X1 U4906 ( .A1(n3891), .A2(n3890), .A3(n3889), .A4(n3888), .ZN(n3897)
         );
  AOI22_X1 U4907 ( .A1(n4034), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4908 ( .A1(n4058), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4909 ( .A1(n4032), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4910 ( .A1(n4019), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3892) );
  NAND4_X1 U4911 ( .A1(n3895), .A2(n3894), .A3(n3893), .A4(n3892), .ZN(n3896)
         );
  NOR2_X1 U4912 ( .A1(n3897), .A2(n3896), .ZN(n3899) );
  AOI22_X1 U4913 ( .A1(n4080), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6603), .ZN(n3898) );
  OAI21_X1 U4914 ( .B1(n4074), .B2(n3899), .A(n3898), .ZN(n3902) );
  INV_X1 U4915 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6988) );
  NAND2_X1 U4916 ( .A1(n3900), .A2(n6988), .ZN(n3901) );
  NAND2_X1 U4917 ( .A1(n3941), .A2(n3901), .ZN(n5471) );
  MUX2_X1 U4918 ( .A(n3902), .B(n5471), .S(n4502), .Z(n4442) );
  AOI22_X1 U4919 ( .A1(n4032), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4920 ( .A1(n4053), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4921 ( .A1(n4014), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4922 ( .A1(n4034), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3903) );
  NAND4_X1 U4923 ( .A1(n3906), .A2(n3905), .A3(n3904), .A4(n3903), .ZN(n3913)
         );
  AOI22_X1 U4924 ( .A1(n3117), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4925 ( .A1(n4058), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4926 ( .A1(n4019), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4927 ( .A1(n4056), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3908) );
  NAND4_X1 U4928 ( .A1(n3911), .A2(n3910), .A3(n3909), .A4(n3908), .ZN(n3912)
         );
  NOR2_X1 U4929 ( .A1(n3913), .A2(n3912), .ZN(n3928) );
  AOI22_X1 U4930 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n4056), .B1(n4058), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4931 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n3117), .B1(n4041), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4932 ( .A1(n4014), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4933 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n4057), .B1(n3907), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3914) );
  NAND4_X1 U4934 ( .A1(n3917), .A2(n3916), .A3(n3915), .A4(n3914), .ZN(n3923)
         );
  AOI22_X1 U4935 ( .A1(n4032), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3921) );
  AOI22_X1 U4936 ( .A1(n4053), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4937 ( .A1(n4034), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4938 ( .A1(n4019), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3973), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3918) );
  NAND4_X1 U4939 ( .A1(n3921), .A2(n3920), .A3(n3919), .A4(n3918), .ZN(n3922)
         );
  NOR2_X1 U4940 ( .A1(n3923), .A2(n3922), .ZN(n3927) );
  XOR2_X1 U4941 ( .A(n3928), .B(n3927), .Z(n3925) );
  INV_X1 U4942 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4643) );
  INV_X1 U4943 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5788) );
  OAI22_X1 U4944 ( .A1(n3659), .A2(n4643), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5788), .ZN(n3924) );
  AOI21_X1 U4945 ( .B1(n4050), .B2(n3925), .A(n3924), .ZN(n3926) );
  XNOR2_X1 U4946 ( .A(n3941), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5791)
         );
  MUX2_X1 U4947 ( .A(n3926), .B(n5791), .S(n4502), .Z(n5460) );
  NOR2_X1 U4948 ( .A1(n3928), .A2(n3927), .ZN(n3950) );
  AOI22_X1 U4949 ( .A1(n4032), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4950 ( .A1(n4053), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4951 ( .A1(n4014), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4952 ( .A1(n4034), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3929) );
  NAND4_X1 U4953 ( .A1(n3932), .A2(n3931), .A3(n3930), .A4(n3929), .ZN(n3938)
         );
  AOI22_X1 U4954 ( .A1(n3117), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3936) );
  AOI22_X1 U4955 ( .A1(n4058), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4956 ( .A1(n4019), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4957 ( .A1(n4056), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3973), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3933) );
  NAND4_X1 U4958 ( .A1(n3936), .A2(n3935), .A3(n3934), .A4(n3933), .ZN(n3937)
         );
  INV_X1 U4959 ( .A(n3949), .ZN(n3939) );
  XNOR2_X1 U4960 ( .A(n3950), .B(n3939), .ZN(n3940) );
  NAND2_X1 U4961 ( .A1(n3940), .A2(n4050), .ZN(n3948) );
  AOI22_X1 U4962 ( .A1(n4080), .A2(EAX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n4079), .ZN(n3947) );
  INV_X1 U4963 ( .A(n3941), .ZN(n3942) );
  INV_X1 U4964 ( .A(n3943), .ZN(n3944) );
  NAND2_X1 U4965 ( .A1(n3944), .A2(n3189), .ZN(n3945) );
  NAND2_X1 U4966 ( .A1(n3963), .A2(n3945), .ZN(n5451) );
  NAND2_X1 U4967 ( .A1(n5451), .A2(n4502), .ZN(n3946) );
  NAND3_X1 U4968 ( .A1(n3948), .A2(n3947), .A3(n3946), .ZN(n4426) );
  NAND2_X1 U4969 ( .A1(n3950), .A2(n3949), .ZN(n3967) );
  AOI22_X1 U4970 ( .A1(n3113), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4971 ( .A1(n3117), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3953) );
  AOI22_X1 U4972 ( .A1(n4019), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3952) );
  AOI22_X1 U4973 ( .A1(n4057), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3973), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3951) );
  NAND4_X1 U4974 ( .A1(n3954), .A2(n3953), .A3(n3952), .A4(n3951), .ZN(n3960)
         );
  AOI22_X1 U4975 ( .A1(n4053), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4032), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4976 ( .A1(n4034), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4977 ( .A1(n4056), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4978 ( .A1(n4014), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3955) );
  NAND4_X1 U4979 ( .A1(n3958), .A2(n3957), .A3(n3956), .A4(n3955), .ZN(n3959)
         );
  NOR2_X1 U4980 ( .A1(n3960), .A2(n3959), .ZN(n3968) );
  XOR2_X1 U4981 ( .A(n3967), .B(n3968), .Z(n3962) );
  INV_X1 U4982 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4725) );
  OAI22_X1 U4983 ( .A1(n3659), .A2(n4725), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6906), .ZN(n3961) );
  AOI21_X1 U4984 ( .B1(n3962), .B2(n4050), .A(n3961), .ZN(n3965) );
  NAND2_X1 U4985 ( .A1(n3963), .A2(n6906), .ZN(n3964) );
  AND2_X1 U4986 ( .A1(n3984), .A2(n3964), .ZN(n5768) );
  MUX2_X1 U4987 ( .A(n3965), .B(n5768), .S(n4502), .Z(n3966) );
  INV_X1 U4988 ( .A(n5427), .ZN(n3988) );
  NOR2_X1 U4989 ( .A1(n3968), .A2(n3967), .ZN(n3990) );
  AOI22_X1 U4990 ( .A1(n4032), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4991 ( .A1(n4053), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3971) );
  AOI22_X1 U4992 ( .A1(n4014), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3970) );
  AOI22_X1 U4993 ( .A1(n4034), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3969) );
  NAND4_X1 U4994 ( .A1(n3972), .A2(n3971), .A3(n3970), .A4(n3969), .ZN(n3979)
         );
  AOI22_X1 U4995 ( .A1(n3117), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4996 ( .A1(n4058), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4997 ( .A1(n4019), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U4998 ( .A1(n4056), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3973), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3974) );
  NAND4_X1 U4999 ( .A1(n3977), .A2(n3976), .A3(n3975), .A4(n3974), .ZN(n3978)
         );
  OR2_X1 U5000 ( .A1(n3979), .A2(n3978), .ZN(n3989) );
  INV_X1 U5001 ( .A(n3989), .ZN(n3980) );
  XNOR2_X1 U5002 ( .A(n3990), .B(n3980), .ZN(n3983) );
  INV_X1 U5003 ( .A(EAX_REG_26__SCAN_IN), .ZN(n3981) );
  OAI22_X1 U5004 ( .A1(n3659), .A2(n3981), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6853), .ZN(n3982) );
  AOI21_X1 U5005 ( .B1(n3983), .B2(n4050), .A(n3982), .ZN(n3986) );
  NAND2_X1 U5006 ( .A1(n3984), .A2(n6853), .ZN(n3985) );
  AND2_X1 U5007 ( .A1(n4007), .A2(n3985), .ZN(n5762) );
  MUX2_X1 U5008 ( .A(n3986), .B(n5762), .S(n4502), .Z(n5429) );
  NAND2_X1 U5009 ( .A1(n3990), .A2(n3989), .ZN(n4012) );
  AOI22_X1 U5010 ( .A1(n4033), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3991), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U5011 ( .A1(n3116), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U5012 ( .A1(n4014), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U5013 ( .A1(n4058), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3992) );
  NAND4_X1 U5014 ( .A1(n3995), .A2(n3994), .A3(n3993), .A4(n3992), .ZN(n4002)
         );
  AOI22_X1 U5015 ( .A1(n4034), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U5016 ( .A1(n3118), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U5017 ( .A1(n4019), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U5018 ( .A1(n4056), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3997) );
  NAND4_X1 U5019 ( .A1(n4000), .A2(n3999), .A3(n3998), .A4(n3997), .ZN(n4001)
         );
  NOR2_X1 U5020 ( .A1(n4002), .A2(n4001), .ZN(n4013) );
  XOR2_X1 U5021 ( .A(n4012), .B(n4013), .Z(n4005) );
  INV_X1 U5022 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4003) );
  INV_X1 U5023 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5753) );
  OAI22_X1 U5024 ( .A1(n3659), .A2(n4003), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5753), .ZN(n4004) );
  AOI21_X1 U5025 ( .B1(n4005), .B2(n4050), .A(n4004), .ZN(n4006) );
  XNOR2_X1 U5026 ( .A(n4007), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5751)
         );
  MUX2_X1 U5027 ( .A(n4006), .B(n5751), .S(n4502), .Z(n5416) );
  INV_X1 U5028 ( .A(n4007), .ZN(n4008) );
  INV_X1 U5029 ( .A(n4009), .ZN(n4010) );
  INV_X1 U5030 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U5031 ( .A1(n4010), .A2(n5405), .ZN(n4011) );
  NAND2_X1 U5032 ( .A1(n4076), .A2(n4011), .ZN(n5745) );
  NOR2_X1 U5033 ( .A1(n4013), .A2(n4012), .ZN(n4031) );
  AOI22_X1 U5034 ( .A1(n4032), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U5035 ( .A1(n4033), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3452), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U5036 ( .A1(n4014), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U5037 ( .A1(n4034), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4015) );
  NAND4_X1 U5038 ( .A1(n4018), .A2(n4017), .A3(n4016), .A4(n4015), .ZN(n4025)
         );
  AOI22_X1 U5039 ( .A1(n3117), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U5040 ( .A1(n4058), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U5041 ( .A1(n4019), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U5042 ( .A1(n3360), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4020) );
  NAND4_X1 U5043 ( .A1(n4023), .A2(n4022), .A3(n4021), .A4(n4020), .ZN(n4024)
         );
  OR2_X1 U5044 ( .A1(n4025), .A2(n4024), .ZN(n4030) );
  XNOR2_X1 U5045 ( .A(n4031), .B(n4030), .ZN(n4027) );
  AOI22_X1 U5046 ( .A1(n4080), .A2(EAX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6603), .ZN(n4026) );
  OAI21_X1 U5047 ( .B1(n4027), .B2(n4074), .A(n4026), .ZN(n4029) );
  MUX2_X1 U5048 ( .A(n5745), .B(n4029), .S(n4028), .Z(n5403) );
  NAND2_X1 U5049 ( .A1(n4031), .A2(n4030), .ZN(n4069) );
  AOI22_X1 U5050 ( .A1(n4033), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4032), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4038) );
  AOI22_X1 U5051 ( .A1(n4055), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4056), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U5052 ( .A1(n4034), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4054), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U5053 ( .A1(n4058), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4035) );
  NAND4_X1 U5054 ( .A1(n4038), .A2(n4037), .A3(n4036), .A4(n4035), .ZN(n4047)
         );
  AOI22_X1 U5055 ( .A1(n3452), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U5056 ( .A1(n3117), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U5057 ( .A1(n4019), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U5058 ( .A1(n4041), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4042) );
  NAND4_X1 U5059 ( .A1(n4045), .A2(n4044), .A3(n4043), .A4(n4042), .ZN(n4046)
         );
  NOR2_X1 U5060 ( .A1(n4047), .A2(n4046), .ZN(n4070) );
  XOR2_X1 U5061 ( .A(n4069), .B(n4070), .Z(n4051) );
  INV_X1 U5062 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4048) );
  INV_X1 U5063 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5731) );
  OAI22_X1 U5064 ( .A1(n3659), .A2(n4048), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5731), .ZN(n4049) );
  AOI21_X1 U5065 ( .B1(n4051), .B2(n4050), .A(n4049), .ZN(n4052) );
  XNOR2_X1 U5066 ( .A(n4076), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5729)
         );
  MUX2_X1 U5067 ( .A(n4052), .B(n5729), .S(n4502), .Z(n4450) );
  AOI22_X1 U5068 ( .A1(n4053), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4062) );
  AOI22_X1 U5069 ( .A1(n4055), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3509), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U5070 ( .A1(n4056), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4041), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U5071 ( .A1(n4058), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4059) );
  NAND4_X1 U5072 ( .A1(n4062), .A2(n4061), .A3(n4060), .A4(n4059), .ZN(n4068)
         );
  AOI22_X1 U5073 ( .A1(n4032), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4066) );
  AOI22_X1 U5074 ( .A1(n4034), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U5075 ( .A1(n4019), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3907), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U5076 ( .A1(n3117), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4040), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4063) );
  NAND4_X1 U5077 ( .A1(n4066), .A2(n4065), .A3(n4064), .A4(n4063), .ZN(n4067)
         );
  NOR2_X1 U5078 ( .A1(n4068), .A2(n4067), .ZN(n4072) );
  NOR2_X1 U5079 ( .A1(n4070), .A2(n4069), .ZN(n4071) );
  XOR2_X1 U5080 ( .A(n4072), .B(n4071), .Z(n4075) );
  AOI22_X1 U5081 ( .A1(n4080), .A2(EAX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6603), .ZN(n4073) );
  OAI21_X1 U5082 ( .B1(n4075), .B2(n4074), .A(n4073), .ZN(n4078) );
  INV_X1 U5083 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4077) );
  XNOR2_X1 U5084 ( .A(n4144), .B(n4077), .ZN(n5724) );
  MUX2_X1 U5085 ( .A(n4078), .B(n5724), .S(n4502), .Z(n4532) );
  AOI22_X1 U5086 ( .A1(n4080), .A2(EAX_REG_31__SCAN_IN), .B1(n4079), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4081) );
  INV_X1 U5087 ( .A(n4081), .ZN(n4082) );
  NAND2_X1 U5088 ( .A1(n4715), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6724) );
  XNOR2_X1 U5089 ( .A(n6756), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4091)
         );
  NAND2_X1 U5090 ( .A1(n6651), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4093) );
  INV_X1 U5091 ( .A(n4093), .ZN(n4083) );
  NAND2_X1 U5092 ( .A1(n4091), .A2(n4083), .ZN(n4085) );
  NAND2_X1 U5093 ( .A1(n4975), .A2(n6756), .ZN(n4084) );
  NAND2_X1 U5094 ( .A1(n4085), .A2(n4084), .ZN(n4108) );
  XNOR2_X1 U5095 ( .A(n4785), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4107)
         );
  INV_X1 U5096 ( .A(n4107), .ZN(n4086) );
  NAND2_X1 U5097 ( .A1(n4108), .A2(n4086), .ZN(n4088) );
  NAND2_X1 U5098 ( .A1(n4785), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4087) );
  NAND2_X1 U5099 ( .A1(n4088), .A2(n4087), .ZN(n4118) );
  XNOR2_X1 U5100 ( .A(n6781), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4116)
         );
  XNOR2_X1 U5101 ( .A(n4118), .B(n4116), .ZN(n4121) );
  NAND2_X1 U5102 ( .A1(n4127), .A2(n4620), .ZN(n4090) );
  NAND2_X1 U5103 ( .A1(n4090), .A2(n4089), .ZN(n4101) );
  XNOR2_X1 U5104 ( .A(n4091), .B(n4093), .ZN(n4262) );
  NAND2_X1 U5105 ( .A1(n3269), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4092) );
  AND2_X1 U5106 ( .A1(n4093), .A2(n4092), .ZN(n4094) );
  AND2_X1 U5107 ( .A1(n4127), .A2(n4094), .ZN(n4098) );
  NAND2_X1 U5108 ( .A1(n3409), .A2(n4094), .ZN(n4095) );
  NAND2_X1 U5109 ( .A1(n4095), .A2(n4287), .ZN(n4097) );
  NAND2_X1 U5110 ( .A1(n3410), .A2(n4287), .ZN(n4096) );
  NAND2_X1 U5111 ( .A1(n4096), .A2(n3110), .ZN(n4111) );
  NAND2_X1 U5112 ( .A1(n4097), .A2(n4111), .ZN(n4102) );
  OAI211_X1 U5113 ( .C1(n4101), .C2(n4262), .A(n4098), .B(n4102), .ZN(n4100)
         );
  NAND3_X1 U5114 ( .A1(n4101), .A2(STATE2_REG_0__SCAN_IN), .A3(n4262), .ZN(
        n4099) );
  NAND3_X1 U5115 ( .A1(n4100), .A2(n4135), .A3(n4099), .ZN(n4106) );
  INV_X1 U5116 ( .A(n4101), .ZN(n4104) );
  INV_X1 U5117 ( .A(n4102), .ZN(n4103) );
  NAND3_X1 U5118 ( .A1(n4104), .A2(n4103), .A3(n4262), .ZN(n4105) );
  NAND2_X1 U5119 ( .A1(n4106), .A2(n4105), .ZN(n4110) );
  NAND2_X1 U5120 ( .A1(n4110), .A2(n4111), .ZN(n4109) );
  XNOR2_X1 U5121 ( .A(n4108), .B(n4107), .ZN(n4263) );
  NAND3_X1 U5122 ( .A1(n4109), .A2(n4263), .A3(n4127), .ZN(n4115) );
  INV_X1 U5123 ( .A(n4110), .ZN(n4113) );
  OAI21_X1 U5124 ( .B1(n4263), .B2(n4122), .A(n4111), .ZN(n4112) );
  NAND2_X1 U5125 ( .A1(n4113), .A2(n4112), .ZN(n4114) );
  OAI211_X1 U5126 ( .C1(n4121), .C2(n4219), .A(n4115), .B(n4114), .ZN(n4133)
         );
  INV_X1 U5127 ( .A(n4116), .ZN(n4117) );
  NAND2_X1 U5128 ( .A1(n4118), .A2(n4117), .ZN(n4120) );
  NAND2_X1 U5129 ( .A1(n6781), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4119) );
  NAND2_X1 U5130 ( .A1(n4120), .A2(n4119), .ZN(n4124) );
  NAND2_X1 U5131 ( .A1(n4634), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4125) );
  NAND2_X1 U5132 ( .A1(n4130), .A2(n4121), .ZN(n4265) );
  NAND2_X1 U5133 ( .A1(n4122), .A2(n4265), .ZN(n4132) );
  NOR2_X1 U5134 ( .A1(n4634), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4123)
         );
  NAND2_X1 U5135 ( .A1(n4127), .A2(n4134), .ZN(n4129) );
  NAND2_X1 U5136 ( .A1(n4872), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4128) );
  OAI211_X1 U5137 ( .C1(n4135), .C2(n4130), .A(n4129), .B(n4128), .ZN(n4131)
         );
  AOI21_X1 U5138 ( .B1(n4133), .B2(n4132), .A(n4131), .ZN(n4137) );
  OR2_X2 U5139 ( .A1(n4137), .A2(n4136), .ZN(n4772) );
  NAND2_X1 U5140 ( .A1(n4792), .A2(n4925), .ZN(n4139) );
  NAND2_X1 U5141 ( .A1(n4140), .A2(n4139), .ZN(n4279) );
  NAND2_X1 U5142 ( .A1(n4147), .A2(n6655), .ZN(n6743) );
  NAND2_X1 U5143 ( .A1(n6743), .A2(n4872), .ZN(n4141) );
  NAND2_X1 U5144 ( .A1(n4872), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4143) );
  NAND2_X1 U5145 ( .A1(n6129), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4142) );
  NAND2_X1 U5146 ( .A1(n4143), .A2(n4142), .ZN(n4704) );
  INV_X1 U5147 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4145) );
  NAND2_X1 U5148 ( .A1(n6433), .A2(REIP_REG_31__SCAN_IN), .ZN(n5901) );
  NAND2_X1 U5149 ( .A1(n6354), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4148)
         );
  OAI211_X1 U5150 ( .C1(n6363), .C2(n5389), .A(n5901), .B(n4148), .ZN(n4149)
         );
  NAND2_X1 U5151 ( .A1(n4887), .A2(n4209), .ZN(n4156) );
  NAND2_X1 U5152 ( .A1(n4150), .A2(n4159), .ZN(n4176) );
  OAI21_X1 U5153 ( .B1(n4159), .B2(n4150), .A(n4176), .ZN(n4153) );
  INV_X1 U5154 ( .A(n4381), .ZN(n4152) );
  OAI211_X1 U5155 ( .C1(n4153), .C2(n6746), .A(n4152), .B(n4089), .ZN(n4154)
         );
  INV_X1 U5156 ( .A(n4154), .ZN(n4155) );
  NAND2_X1 U5157 ( .A1(n4156), .A2(n4155), .ZN(n4731) );
  OAI21_X1 U5158 ( .B1(n6746), .B2(n4159), .A(n4168), .ZN(n4160) );
  INV_X1 U5159 ( .A(n4160), .ZN(n4161) );
  NAND2_X1 U5160 ( .A1(n4691), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4162)
         );
  INV_X1 U5161 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4673) );
  NAND2_X1 U5162 ( .A1(n4162), .A2(n4673), .ZN(n4164) );
  AND2_X1 U5163 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4163) );
  NAND2_X1 U5164 ( .A1(n4691), .A2(n4163), .ZN(n4165) );
  AND2_X1 U5165 ( .A1(n4164), .A2(n4165), .ZN(n4732) );
  NAND2_X1 U5166 ( .A1(n4731), .A2(n4732), .ZN(n4166) );
  NAND2_X1 U5167 ( .A1(n4166), .A2(n4165), .ZN(n6355) );
  NAND2_X1 U5168 ( .A1(n6355), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4171)
         );
  XNOR2_X1 U5169 ( .A(n4176), .B(n4174), .ZN(n4169) );
  OAI21_X1 U5170 ( .B1(n4169), .B2(n6746), .A(n4168), .ZN(n4170) );
  NAND2_X1 U5171 ( .A1(n4171), .A2(n6356), .ZN(n4173) );
  OR2_X1 U5172 ( .A1(n6355), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4172)
         );
  NAND2_X1 U5173 ( .A1(n5027), .A2(n4209), .ZN(n4180) );
  INV_X1 U5174 ( .A(n4174), .ZN(n4175) );
  NAND2_X1 U5175 ( .A1(n4176), .A2(n4175), .ZN(n4185) );
  INV_X1 U5176 ( .A(n4184), .ZN(n4177) );
  XNOR2_X1 U5177 ( .A(n4185), .B(n4177), .ZN(n4178) );
  NAND2_X1 U5178 ( .A1(n4178), .A2(n4151), .ZN(n4179) );
  INV_X1 U5179 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6430) );
  NAND2_X1 U5180 ( .A1(n4181), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4182)
         );
  NAND2_X1 U5181 ( .A1(n4183), .A2(n4209), .ZN(n4188) );
  NAND2_X1 U5182 ( .A1(n4185), .A2(n4184), .ZN(n4193) );
  XNOR2_X1 U5183 ( .A(n4193), .B(n4191), .ZN(n4186) );
  NAND2_X1 U5184 ( .A1(n4186), .A2(n4151), .ZN(n4187) );
  NAND2_X1 U5185 ( .A1(n4188), .A2(n4187), .ZN(n4189) );
  INV_X1 U5186 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6420) );
  NAND2_X1 U5187 ( .A1(n4190), .A2(n4209), .ZN(n4196) );
  INV_X1 U5188 ( .A(n4191), .ZN(n4192) );
  OR2_X1 U5189 ( .A1(n4193), .A2(n4192), .ZN(n4201) );
  XNOR2_X1 U5190 ( .A(n4201), .B(n4202), .ZN(n4194) );
  NAND2_X1 U5191 ( .A1(n4194), .A2(n4151), .ZN(n4195) );
  NAND2_X1 U5192 ( .A1(n4196), .A2(n4195), .ZN(n4197) );
  INV_X1 U5193 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6879) );
  XNOR2_X1 U5194 ( .A(n4197), .B(n6879), .ZN(n5092) );
  NAND2_X1 U5195 ( .A1(n4197), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4198)
         );
  NAND3_X1 U5196 ( .A1(n4199), .A2(n4209), .A3(n4200), .ZN(n4206) );
  INV_X1 U5197 ( .A(n4201), .ZN(n4203) );
  NAND2_X1 U5198 ( .A1(n4203), .A2(n4202), .ZN(n4210) );
  XNOR2_X1 U5199 ( .A(n4210), .B(n4211), .ZN(n4204) );
  NAND2_X1 U5200 ( .A1(n4204), .A2(n4151), .ZN(n4205) );
  INV_X1 U5201 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6401) );
  NAND2_X1 U5202 ( .A1(n4208), .A2(n4209), .ZN(n4215) );
  INV_X1 U5203 ( .A(n4210), .ZN(n4212) );
  NAND2_X1 U5204 ( .A1(n4212), .A2(n4211), .ZN(n4224) );
  XNOR2_X1 U5205 ( .A(n4224), .B(n4222), .ZN(n4213) );
  NAND2_X1 U5206 ( .A1(n4213), .A2(n4151), .ZN(n4214) );
  NAND2_X1 U5207 ( .A1(n4215), .A2(n4214), .ZN(n4216) );
  XNOR2_X1 U5208 ( .A(n4216), .B(n6389), .ZN(n5206) );
  NAND2_X1 U5209 ( .A1(n4216), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4217)
         );
  INV_X1 U5210 ( .A(n4218), .ZN(n4220) );
  NAND2_X2 U5211 ( .A1(n4199), .A2(n4221), .ZN(n4249) );
  NAND2_X1 U5212 ( .A1(n4151), .A2(n4222), .ZN(n4223) );
  OR2_X1 U5213 ( .A1(n4224), .A2(n4223), .ZN(n4225) );
  NAND2_X1 U5214 ( .A1(n4249), .A2(n4225), .ZN(n4226) );
  XNOR2_X1 U5215 ( .A(n4226), .B(n6858), .ZN(n5890) );
  NAND2_X1 U5216 ( .A1(n4226), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4227)
         );
  INV_X2 U5217 ( .A(n4249), .ZN(n4229) );
  INV_X1 U5218 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6364) );
  INV_X1 U5219 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5862) );
  INV_X1 U5220 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4334) );
  INV_X1 U5221 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6081) );
  AND4_X1 U5222 ( .A1(n6364), .A2(n5862), .A3(n4334), .A4(n6081), .ZN(n4228)
         );
  NOR2_X1 U5223 ( .A1(n3105), .A2(n4228), .ZN(n4232) );
  INV_X4 U5224 ( .A(n4229), .ZN(n5848) );
  NAND2_X1 U5225 ( .A1(n5848), .A2(n6364), .ZN(n5880) );
  NAND2_X1 U5226 ( .A1(n3107), .A2(n4334), .ZN(n5865) );
  NAND2_X1 U5227 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5864) );
  NAND2_X1 U5228 ( .A1(n3106), .A2(n5864), .ZN(n4230) );
  AND3_X1 U5229 ( .A1(n5880), .A2(n5865), .A3(n4230), .ZN(n4231) );
  XNOR2_X1 U5230 ( .A(n5848), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5857)
         );
  INV_X1 U5231 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6046) );
  NAND2_X1 U5232 ( .A1(n3107), .A2(n6046), .ZN(n4233) );
  INV_X1 U5233 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4234) );
  OR2_X1 U5234 ( .A1(n3107), .A2(n4234), .ZN(n4235) );
  NAND2_X1 U5235 ( .A1(n3106), .A2(n6035), .ZN(n4237) );
  AND2_X1 U5236 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4403) );
  NAND2_X1 U5237 ( .A1(n4403), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4238) );
  INV_X1 U5238 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6010) );
  INV_X1 U5239 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6907) );
  AND3_X1 U5240 ( .A1(n6010), .A2(n6022), .A3(n6907), .ZN(n4239) );
  AND2_X1 U5241 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5985) );
  AND2_X1 U5242 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4490) );
  AND2_X1 U5243 ( .A1(n5985), .A2(n4490), .ZN(n5781) );
  AND2_X1 U5244 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U5245 ( .A1(n5781), .A2(n5896), .ZN(n5772) );
  NAND2_X1 U5246 ( .A1(n3107), .A2(n5772), .ZN(n4241) );
  NOR2_X1 U5247 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5771) );
  NOR2_X1 U5248 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5770) );
  NOR2_X1 U5249 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5986) );
  NAND4_X1 U5250 ( .A1(n5771), .A2(n5770), .A3(n5986), .A4(n6913), .ZN(n4243)
         );
  NAND2_X1 U5251 ( .A1(n5848), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4242) );
  OAI21_X1 U5252 ( .B1(n3106), .B2(n4243), .A(n4242), .ZN(n4244) );
  NAND2_X1 U5253 ( .A1(n5848), .A2(n6913), .ZN(n4245) );
  NAND2_X1 U5254 ( .A1(n5848), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U5255 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4248) );
  NOR2_X1 U5256 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4246) );
  NOR2_X1 U5257 ( .A1(n3106), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5757)
         );
  INV_X1 U5258 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5722) );
  NAND2_X1 U5259 ( .A1(n5722), .A2(n3173), .ZN(n4247) );
  XNOR2_X1 U5260 ( .A(n5848), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5808)
         );
  XNOR2_X1 U5261 ( .A(n5848), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5801)
         );
  INV_X1 U5262 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4250) );
  XOR2_X1 U5263 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .B(n5848), .Z(n5793) );
  INV_X1 U5264 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4436) );
  NAND2_X1 U5265 ( .A1(n4229), .A2(n4436), .ZN(n5785) );
  NOR2_X1 U5266 ( .A1(n5785), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4252)
         );
  INV_X1 U5267 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6889) );
  INV_X1 U5268 ( .A(n4490), .ZN(n4416) );
  NOR3_X1 U5269 ( .A1(n4229), .A2(n6889), .A3(n4416), .ZN(n4251) );
  XNOR2_X1 U5270 ( .A(n4253), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4424)
         );
  NOR2_X1 U5271 ( .A1(n4792), .A2(n3110), .ZN(n4393) );
  INV_X1 U5272 ( .A(n4393), .ZN(n4270) );
  INV_X1 U5273 ( .A(n4279), .ZN(n4257) );
  OR2_X1 U5274 ( .A1(n4254), .A2(n4925), .ZN(n4256) );
  INV_X1 U5275 ( .A(n3788), .ZN(n4255) );
  MUX2_X1 U5276 ( .A(n4256), .B(n6746), .S(n4255), .Z(n4388) );
  NAND2_X1 U5277 ( .A1(n4257), .A2(n4388), .ZN(n4260) );
  NOR2_X1 U5278 ( .A1(n3409), .A2(n4287), .ZN(n4259) );
  NAND2_X1 U5279 ( .A1(n4258), .A2(n4259), .ZN(n4775) );
  NAND2_X1 U5280 ( .A1(n4260), .A2(n4775), .ZN(n4623) );
  NAND2_X1 U5281 ( .A1(n4620), .A2(n4767), .ZN(n4268) );
  NAND2_X1 U5282 ( .A1(n4263), .A2(n4262), .ZN(n4264) );
  OR2_X1 U5283 ( .A1(n4265), .A2(n4264), .ZN(n4266) );
  NAND2_X1 U5284 ( .A1(n4267), .A2(n4266), .ZN(n4776) );
  NOR2_X1 U5285 ( .A1(READY_N), .A2(n4776), .ZN(n4615) );
  NAND3_X1 U5286 ( .A1(n4268), .A2(n4615), .A3(n3394), .ZN(n4269) );
  OAI211_X1 U5287 ( .C1(n4772), .C2(n4270), .A(n4623), .B(n4269), .ZN(n4271)
         );
  NAND2_X1 U5288 ( .A1(n4271), .A2(n6717), .ZN(n4278) );
  OAI21_X1 U5289 ( .B1(n4620), .B2(n4713), .A(n4811), .ZN(n4618) );
  OAI211_X1 U5290 ( .C1(n4273), .C2(n4618), .A(n4287), .B(n4845), .ZN(n4275)
         );
  NAND2_X1 U5291 ( .A1(n4275), .A2(n4274), .ZN(n4276) );
  INV_X1 U5292 ( .A(n4780), .ZN(n4280) );
  NOR2_X1 U5293 ( .A1(n4279), .A2(n3402), .ZN(n4665) );
  OR2_X1 U5294 ( .A1(n4280), .A2(n4665), .ZN(n4771) );
  INV_X1 U5295 ( .A(n4771), .ZN(n4285) );
  OAI22_X1 U5296 ( .A1(n4281), .A2(n3111), .B1(n3445), .B2(n4378), .ZN(n4282)
         );
  INV_X1 U5297 ( .A(n4282), .ZN(n4284) );
  NAND3_X1 U5298 ( .A1(n4285), .A2(n4284), .A3(n4283), .ZN(n4286) );
  NAND2_X1 U5299 ( .A1(n4424), .A2(n6440), .ZN(n4423) );
  NAND2_X2 U5300 ( .A1(n3413), .A2(n3102), .ZN(n4316) );
  NAND2_X1 U5301 ( .A1(n4909), .A2(n4287), .ZN(n4300) );
  INV_X1 U5302 ( .A(n4300), .ZN(n4294) );
  INV_X1 U5303 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4420) );
  NAND2_X1 U5304 ( .A1(n4348), .A2(n4420), .ZN(n4288) );
  INV_X2 U5305 ( .A(n4336), .ZN(n4364) );
  OAI211_X1 U5306 ( .C1(EBX_REG_24__SCAN_IN), .C2(n4316), .A(n4288), .B(n4462), 
        .ZN(n4291) );
  INV_X1 U5307 ( .A(EBX_REG_24__SCAN_IN), .ZN(n4289) );
  NAND2_X1 U5308 ( .A1(n4364), .A2(n4289), .ZN(n4290) );
  INV_X2 U5309 ( .A(n4316), .ZN(n4308) );
  NAND2_X1 U5310 ( .A1(n4462), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4292)
         );
  OAI211_X1 U5311 ( .C1(n4316), .C2(EBX_REG_3__SCAN_IN), .A(n4348), .B(n4292), 
        .ZN(n4293) );
  OAI21_X1 U5312 ( .B1(n4468), .B2(EBX_REG_3__SCAN_IN), .A(n4293), .ZN(n4879)
         );
  NAND2_X1 U5313 ( .A1(n4336), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4295)
         );
  NAND2_X1 U5314 ( .A1(n4300), .A2(n4295), .ZN(n4297) );
  INV_X1 U5315 ( .A(EBX_REG_1__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U5316 ( .A1(n4308), .A2(n5638), .ZN(n4296) );
  NAND2_X1 U5317 ( .A1(n4297), .A2(n4296), .ZN(n4299) );
  NAND2_X1 U5318 ( .A1(n4364), .A2(n5638), .ZN(n4298) );
  NAND2_X1 U5319 ( .A1(n4299), .A2(n4298), .ZN(n4301) );
  MUX2_X1 U5320 ( .A(n4336), .B(n4300), .S(EBX_REG_0__SCAN_IN), .Z(n4692) );
  INV_X1 U5321 ( .A(n4301), .ZN(n4302) );
  AOI21_X2 U5322 ( .B1(n4819), .B2(n4308), .A(n4302), .ZN(n4834) );
  INV_X1 U5323 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6442) );
  NAND2_X1 U5324 ( .A1(n4348), .A2(n6442), .ZN(n4303) );
  OAI211_X1 U5325 ( .C1(EBX_REG_2__SCAN_IN), .C2(n4316), .A(n4303), .B(n4462), 
        .ZN(n4305) );
  INV_X1 U5326 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4835) );
  NAND2_X1 U5327 ( .A1(n4364), .A2(n4835), .ZN(n4304) );
  NAND2_X1 U5328 ( .A1(n4305), .A2(n4304), .ZN(n4833) );
  NAND2_X1 U5329 ( .A1(n4834), .A2(n4833), .ZN(n4832) );
  NAND2_X1 U5330 ( .A1(n4348), .A2(n6420), .ZN(n4309) );
  OAI211_X1 U5331 ( .C1(EBX_REG_4__SCAN_IN), .C2(n4316), .A(n4309), .B(n4462), 
        .ZN(n4311) );
  INV_X1 U5332 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4858) );
  NAND2_X1 U5333 ( .A1(n4364), .A2(n4858), .ZN(n4310) );
  AND2_X1 U5334 ( .A1(n4311), .A2(n4310), .ZN(n4856) );
  INV_X1 U5335 ( .A(n4468), .ZN(n4457) );
  INV_X1 U5336 ( .A(EBX_REG_5__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U5337 ( .A1(n4457), .A2(n6209), .ZN(n4314) );
  NAND2_X1 U5338 ( .A1(n4462), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4312)
         );
  OAI211_X1 U5339 ( .C1(n4316), .C2(EBX_REG_5__SCAN_IN), .A(n4348), .B(n4312), 
        .ZN(n4313) );
  NAND2_X1 U5340 ( .A1(n4462), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4315)
         );
  NAND2_X1 U5341 ( .A1(n4348), .A2(n4315), .ZN(n4318) );
  INV_X1 U5342 ( .A(n4316), .ZN(n4329) );
  INV_X1 U5343 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5026) );
  NAND2_X1 U5344 ( .A1(n4329), .A2(n5026), .ZN(n4317) );
  NAND2_X1 U5345 ( .A1(n4318), .A2(n4317), .ZN(n4320) );
  NAND2_X1 U5346 ( .A1(n4364), .A2(n5026), .ZN(n4319) );
  NAND2_X1 U5347 ( .A1(n4320), .A2(n4319), .ZN(n5023) );
  NAND2_X1 U5348 ( .A1(n4462), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4321)
         );
  OAI211_X1 U5349 ( .C1(n4316), .C2(EBX_REG_7__SCAN_IN), .A(n4348), .B(n4321), 
        .ZN(n4322) );
  OAI21_X1 U5350 ( .B1(n4468), .B2(EBX_REG_7__SCAN_IN), .A(n4322), .ZN(n5136)
         );
  NAND2_X1 U5351 ( .A1(n4348), .A2(n6858), .ZN(n4324) );
  OAI211_X1 U5352 ( .C1(EBX_REG_8__SCAN_IN), .C2(n4316), .A(n4324), .B(n4462), 
        .ZN(n4326) );
  INV_X1 U5353 ( .A(EBX_REG_8__SCAN_IN), .ZN(n7048) );
  NAND2_X1 U5354 ( .A1(n4364), .A2(n7048), .ZN(n4325) );
  NAND2_X1 U5355 ( .A1(n4462), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4327)
         );
  OAI211_X1 U5356 ( .C1(n4316), .C2(EBX_REG_9__SCAN_IN), .A(n4348), .B(n4327), 
        .ZN(n4328) );
  OAI21_X1 U5357 ( .B1(n4468), .B2(EBX_REG_9__SCAN_IN), .A(n4328), .ZN(n6165)
         );
  NAND2_X1 U5358 ( .A1(n4348), .A2(n5862), .ZN(n4330) );
  OAI211_X1 U5359 ( .C1(EBX_REG_10__SCAN_IN), .C2(n4316), .A(n4330), .B(n4462), 
        .ZN(n4332) );
  INV_X1 U5360 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U5361 ( .A1(n4364), .A2(n5671), .ZN(n4331) );
  NAND2_X1 U5362 ( .A1(n4332), .A2(n4331), .ZN(n5608) );
  MUX2_X1 U5363 ( .A(n4468), .B(n4462), .S(EBX_REG_11__SCAN_IN), .Z(n4333) );
  OAI21_X1 U5364 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n4499), .A(n4333), 
        .ZN(n5147) );
  NAND2_X1 U5365 ( .A1(n4348), .A2(n4334), .ZN(n4335) );
  OAI211_X1 U5366 ( .C1(EBX_REG_12__SCAN_IN), .C2(n4316), .A(n4335), .B(n4462), 
        .ZN(n4338) );
  INV_X1 U5367 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5365) );
  NAND2_X1 U5368 ( .A1(n4364), .A2(n5365), .ZN(n4337) );
  MUX2_X1 U5369 ( .A(n4468), .B(n4462), .S(EBX_REG_13__SCAN_IN), .Z(n4339) );
  OAI21_X1 U5370 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n4499), .A(n4339), 
        .ZN(n4340) );
  INV_X1 U5371 ( .A(n4340), .ZN(n5666) );
  NAND2_X1 U5372 ( .A1(n4462), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4341) );
  NAND2_X1 U5373 ( .A1(n4348), .A2(n4341), .ZN(n4343) );
  INV_X1 U5374 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U5375 ( .A1(n4329), .A2(n5661), .ZN(n4342) );
  NAND2_X1 U5376 ( .A1(n4343), .A2(n4342), .ZN(n4345) );
  NAND2_X1 U5377 ( .A1(n4364), .A2(n5661), .ZN(n4344) );
  NAND2_X1 U5378 ( .A1(n4345), .A2(n4344), .ZN(n5580) );
  MUX2_X1 U5379 ( .A(n4468), .B(n4462), .S(EBX_REG_15__SCAN_IN), .Z(n4346) );
  OAI21_X1 U5380 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n4499), .A(n4346), 
        .ZN(n5571) );
  NAND2_X1 U5381 ( .A1(n4348), .A2(n6022), .ZN(n4349) );
  OAI211_X1 U5382 ( .C1(EBX_REG_16__SCAN_IN), .C2(n4316), .A(n4349), .B(n4462), 
        .ZN(n4352) );
  INV_X1 U5383 ( .A(EBX_REG_16__SCAN_IN), .ZN(n4350) );
  NAND2_X1 U5384 ( .A1(n4364), .A2(n4350), .ZN(n4351) );
  INV_X1 U5385 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U5386 ( .A1(n4457), .A2(n5657), .ZN(n4355) );
  NAND2_X1 U5387 ( .A1(n4462), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4353) );
  OAI211_X1 U5388 ( .C1(n4316), .C2(EBX_REG_17__SCAN_IN), .A(n4348), .B(n4353), 
        .ZN(n4354) );
  NOR2_X1 U5389 ( .A1(n4499), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5492)
         );
  MUX2_X1 U5390 ( .A(EBX_REG_18__SCAN_IN), .B(n5492), .S(n4462), .Z(n4357) );
  NOR2_X1 U5391 ( .A1(n4468), .A2(EBX_REG_18__SCAN_IN), .ZN(n4356) );
  NOR2_X1 U5392 ( .A1(n4357), .A2(n4356), .ZN(n5526) );
  NAND2_X1 U5393 ( .A1(n5493), .A2(n5526), .ZN(n5509) );
  INV_X1 U5394 ( .A(EBX_REG_20__SCAN_IN), .ZN(n6881) );
  NAND2_X1 U5395 ( .A1(n4329), .A2(n6881), .ZN(n4359) );
  OR2_X1 U5396 ( .A1(n4499), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4358)
         );
  NAND2_X1 U5397 ( .A1(n4358), .A2(n4359), .ZN(n5498) );
  MUX2_X1 U5398 ( .A(n4359), .B(n5498), .S(n4462), .Z(n4367) );
  INV_X1 U5399 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4360) );
  NAND2_X1 U5400 ( .A1(n4348), .A2(n4360), .ZN(n4362) );
  INV_X1 U5401 ( .A(EBX_REG_19__SCAN_IN), .ZN(n4363) );
  NAND2_X1 U5402 ( .A1(n4329), .A2(n4363), .ZN(n4361) );
  NAND3_X1 U5403 ( .A1(n4362), .A2(n4462), .A3(n4361), .ZN(n4366) );
  NAND2_X1 U5404 ( .A1(n4364), .A2(n4363), .ZN(n4365) );
  NAND2_X1 U5405 ( .A1(n4462), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4370) );
  OAI211_X1 U5406 ( .C1(n4316), .C2(EBX_REG_21__SCAN_IN), .A(n4348), .B(n4370), 
        .ZN(n4371) );
  OAI21_X1 U5407 ( .B1(n4468), .B2(EBX_REG_21__SCAN_IN), .A(n4371), .ZN(n5482)
         );
  NAND2_X1 U5408 ( .A1(n4348), .A2(n4436), .ZN(n4372) );
  OAI211_X1 U5409 ( .C1(EBX_REG_22__SCAN_IN), .C2(n4316), .A(n4372), .B(n4462), 
        .ZN(n4374) );
  INV_X1 U5410 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U5411 ( .A1(n4364), .A2(n5654), .ZN(n4373) );
  NAND2_X1 U5412 ( .A1(n4374), .A2(n4373), .ZN(n4486) );
  MUX2_X1 U5413 ( .A(n4468), .B(n4462), .S(EBX_REG_23__SCAN_IN), .Z(n4375) );
  OAI21_X1 U5414 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n4499), .A(n4375), 
        .ZN(n5462) );
  NOR2_X2 U5415 ( .A1(n4376), .A2(n4377), .ZN(n4461) );
  AOI21_X1 U5416 ( .B1(n4377), .B2(n4376), .A(n4461), .ZN(n5650) );
  OAI21_X1 U5417 ( .B1(n4378), .B2(n3397), .A(n4813), .ZN(n4379) );
  INV_X1 U5418 ( .A(REIP_REG_24__SCAN_IN), .ZN(n5454) );
  NOR2_X1 U5419 ( .A1(n6423), .A2(n5454), .ZN(n4429) );
  NAND2_X1 U5420 ( .A1(n4404), .A2(n5367), .ZN(n6044) );
  NAND2_X1 U5421 ( .A1(n3431), .A2(n4364), .ZN(n4386) );
  AND2_X1 U5422 ( .A1(n4274), .A2(n4620), .ZN(n4382) );
  OAI21_X1 U5423 ( .B1(n4499), .B2(n4382), .A(n4381), .ZN(n4385) );
  AND2_X1 U5424 ( .A1(n4925), .A2(n4620), .ZN(n5626) );
  NAND2_X1 U5425 ( .A1(n5626), .A2(n3409), .ZN(n4384) );
  OAI21_X1 U5426 ( .B1(n4845), .B2(n4287), .A(n3394), .ZN(n4383) );
  NAND4_X1 U5427 ( .A1(n4386), .A2(n4385), .A3(n4384), .A4(n4383), .ZN(n4387)
         );
  NOR2_X1 U5428 ( .A1(n4380), .A2(n4387), .ZN(n4389) );
  NAND2_X1 U5429 ( .A1(n4389), .A2(n4388), .ZN(n4661) );
  OAI21_X1 U5430 ( .B1(n3426), .B2(n4287), .A(n4749), .ZN(n4390) );
  INV_X1 U5431 ( .A(n4394), .ZN(n4391) );
  NAND2_X1 U5432 ( .A1(n4404), .A2(n4391), .ZN(n4405) );
  INV_X1 U5433 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4392) );
  AND2_X1 U5434 ( .A1(n6044), .A2(n4392), .ZN(n4817) );
  NOR2_X1 U5435 ( .A1(n6389), .A2(n6858), .ZN(n6367) );
  NAND3_X1 U5436 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6367), .ZN(n4396) );
  NOR3_X1 U5437 ( .A1(n6430), .A2(n6420), .A3(n6879), .ZN(n6087) );
  NOR2_X1 U5438 ( .A1(n6442), .A2(n4673), .ZN(n6437) );
  NAND3_X1 U5439 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6087), .A3(n6437), 
        .ZN(n6088) );
  NOR2_X1 U5440 ( .A1(n4396), .A2(n6088), .ZN(n6018) );
  NAND2_X1 U5441 ( .A1(n6443), .A2(n6018), .ZN(n6063) );
  NAND2_X1 U5442 ( .A1(n4394), .A2(n4393), .ZN(n4773) );
  INV_X1 U5443 ( .A(n4773), .ZN(n4395) );
  AND2_X2 U5444 ( .A1(n4404), .A2(n4395), .ZN(n6436) );
  AOI21_X1 U5445 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6438) );
  INV_X1 U5446 ( .A(n6438), .ZN(n6086) );
  NAND2_X1 U5447 ( .A1(n6086), .A2(n6087), .ZN(n6393) );
  OR2_X1 U5448 ( .A1(n6401), .A2(n6393), .ZN(n6091) );
  NOR2_X1 U5449 ( .A1(n6091), .A2(n4396), .ZN(n4397) );
  NAND2_X1 U5450 ( .A1(n6436), .A2(n4397), .ZN(n6045) );
  NAND2_X1 U5451 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U5452 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4398) );
  NOR2_X1 U5453 ( .A1(n6064), .A2(n4398), .ZN(n6023) );
  AND2_X1 U5454 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4399) );
  NAND2_X1 U5455 ( .A1(n6023), .A2(n4399), .ZN(n4409) );
  INV_X1 U5456 ( .A(n4409), .ZN(n4400) );
  NAND2_X1 U5457 ( .A1(n6079), .A2(n4400), .ZN(n6008) );
  INV_X1 U5458 ( .A(n4403), .ZN(n4401) );
  OR2_X2 U5459 ( .A1(n6008), .A2(n4401), .ZN(n5995) );
  INV_X1 U5460 ( .A(n5985), .ZN(n4402) );
  NOR2_X1 U5461 ( .A1(n5995), .A2(n4402), .ZN(n4489) );
  NAND2_X1 U5462 ( .A1(n4489), .A2(n4490), .ZN(n5965) );
  OR2_X1 U5463 ( .A1(n6045), .A2(n4409), .ZN(n5980) );
  AND2_X1 U5464 ( .A1(n5985), .A2(n4403), .ZN(n4410) );
  INV_X1 U5465 ( .A(n4410), .ZN(n4407) );
  NOR2_X1 U5466 ( .A1(n4404), .A2(n6433), .ZN(n4697) );
  INV_X1 U5467 ( .A(n4405), .ZN(n6047) );
  OR2_X1 U5468 ( .A1(n6436), .A2(n6047), .ZN(n4414) );
  AND2_X1 U5469 ( .A1(n4414), .A2(n4392), .ZN(n4695) );
  NOR2_X1 U5470 ( .A1(n4697), .A2(n4695), .ZN(n6391) );
  INV_X1 U5471 ( .A(n6391), .ZN(n4406) );
  OR2_X1 U5472 ( .A1(n6436), .A2(n4406), .ZN(n6017) );
  OAI21_X1 U5473 ( .B1(n5980), .B2(n4407), .A(n6017), .ZN(n4413) );
  INV_X1 U5474 ( .A(n6018), .ZN(n4408) );
  NOR2_X1 U5475 ( .A1(n4409), .A2(n4408), .ZN(n5979) );
  AOI21_X1 U5476 ( .B1(n4410), .B2(n5979), .A(n6392), .ZN(n4411) );
  INV_X1 U5477 ( .A(n4411), .ZN(n4412) );
  AND2_X1 U5478 ( .A1(n4413), .A2(n4412), .ZN(n4488) );
  INV_X1 U5479 ( .A(n4414), .ZN(n4415) );
  NAND2_X1 U5480 ( .A1(n4415), .A2(n6044), .ZN(n6394) );
  NAND2_X1 U5481 ( .A1(n6394), .A2(n4416), .ZN(n4417) );
  NAND2_X1 U5482 ( .A1(n4488), .A2(n4417), .ZN(n5963) );
  INV_X1 U5483 ( .A(n6436), .ZN(n4418) );
  AOI21_X1 U5484 ( .B1(n5983), .B2(n4418), .A(n5896), .ZN(n4419) );
  INV_X1 U5485 ( .A(n5944), .ZN(n5955) );
  AOI211_X1 U5486 ( .C1(n5965), .C2(n4420), .A(n5955), .B(n5771), .ZN(n4421)
         );
  AOI211_X1 U5487 ( .C1(n5650), .C2(n6435), .A(n4429), .B(n4421), .ZN(n4422)
         );
  NAND2_X1 U5488 ( .A1(n4423), .A2(n4422), .ZN(U2994) );
  NAND2_X1 U5489 ( .A1(n4424), .A2(n6358), .ZN(n4433) );
  NOR2_X1 U5490 ( .A1(n4425), .A2(n4426), .ZN(n4427) );
  NOR2_X1 U5491 ( .A1(n6363), .A2(n5451), .ZN(n4428) );
  AOI211_X1 U5492 ( .C1(n6354), .C2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n4429), 
        .B(n4428), .ZN(n4430) );
  NAND2_X1 U5493 ( .A1(n4433), .A2(n4432), .ZN(U2962) );
  INV_X1 U5494 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4434) );
  OAI21_X1 U5495 ( .B1(n4229), .B2(n4436), .A(n5785), .ZN(n4437) );
  NAND2_X1 U5496 ( .A1(n4484), .A2(n6358), .ZN(n4448) );
  INV_X1 U5497 ( .A(n5480), .ZN(n4440) );
  NOR2_X1 U5498 ( .A1(n4439), .A2(n4440), .ZN(n4443) );
  OAI21_X1 U5499 ( .B1(n4443), .B2(n4442), .A(n4441), .ZN(n5697) );
  INV_X1 U5500 ( .A(REIP_REG_22__SCAN_IN), .ZN(n5472) );
  NOR2_X1 U5501 ( .A1(n6423), .A2(n5472), .ZN(n4492) );
  NOR2_X1 U5502 ( .A1(n6363), .A2(n5471), .ZN(n4444) );
  AOI211_X1 U5503 ( .C1(n6354), .C2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n4492), 
        .B(n4444), .ZN(n4445) );
  INV_X1 U5504 ( .A(n4446), .ZN(n4447) );
  NAND2_X1 U5505 ( .A1(n4448), .A2(n4447), .ZN(U2964) );
  INV_X1 U5506 ( .A(n4534), .ZN(n4451) );
  NAND3_X1 U5507 ( .A1(n4274), .A2(n5374), .A3(n3445), .ZN(n4454) );
  NOR2_X1 U5508 ( .A1(n4454), .A2(n4453), .ZN(n4840) );
  NAND3_X1 U5509 ( .A1(n4840), .A2(n4294), .A3(n4620), .ZN(n4455) );
  NAND2_X2 U5510 ( .A1(n6266), .A2(n3585), .ZN(n5670) );
  INV_X1 U5511 ( .A(EBX_REG_25__SCAN_IN), .ZN(n6959) );
  NAND2_X1 U5512 ( .A1(n4457), .A2(n6959), .ZN(n4460) );
  NAND2_X1 U5513 ( .A1(n4462), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4458) );
  OAI211_X1 U5514 ( .C1(n4316), .C2(EBX_REG_25__SCAN_IN), .A(n4348), .B(n4458), 
        .ZN(n4459) );
  NAND2_X1 U5515 ( .A1(n4462), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4463) );
  NAND2_X1 U5516 ( .A1(n4348), .A2(n4463), .ZN(n4465) );
  INV_X1 U5517 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U5518 ( .A1(n4329), .A2(n5648), .ZN(n4464) );
  NAND2_X1 U5519 ( .A1(n4465), .A2(n4464), .ZN(n4467) );
  NAND2_X1 U5520 ( .A1(n4364), .A2(n5648), .ZN(n4466) );
  NAND2_X1 U5521 ( .A1(n4467), .A2(n4466), .ZN(n5432) );
  MUX2_X1 U5522 ( .A(n4468), .B(n4462), .S(EBX_REG_27__SCAN_IN), .Z(n4469) );
  OAI21_X1 U5523 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n4499), .A(n4469), 
        .ZN(n5417) );
  INV_X1 U5524 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6878) );
  NAND2_X1 U5525 ( .A1(n4348), .A2(n6878), .ZN(n4470) );
  OAI211_X1 U5526 ( .C1(EBX_REG_28__SCAN_IN), .C2(n4316), .A(n4470), .B(n4462), 
        .ZN(n4473) );
  INV_X1 U5527 ( .A(EBX_REG_28__SCAN_IN), .ZN(n4471) );
  NAND2_X1 U5528 ( .A1(n4364), .A2(n4471), .ZN(n4472) );
  INV_X1 U5529 ( .A(n4499), .ZN(n4694) );
  NOR2_X1 U5530 ( .A1(n4316), .A2(EBX_REG_29__SCAN_IN), .ZN(n4474) );
  AOI21_X1 U5531 ( .B1(n4694), .B2(n3173), .A(n4474), .ZN(n4475) );
  NAND2_X2 U5532 ( .A1(n5406), .A2(n4475), .ZN(n4537) );
  INV_X1 U5533 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4480) );
  NAND2_X1 U5534 ( .A1(n4364), .A2(n4480), .ZN(n4476) );
  INV_X1 U5535 ( .A(n5406), .ZN(n4540) );
  OAI22_X1 U5536 ( .A1(n4537), .A2(n4364), .B1(n4476), .B2(n4540), .ZN(n4498)
         );
  NAND2_X1 U5537 ( .A1(n4475), .A2(n4462), .ZN(n4477) );
  NAND2_X1 U5538 ( .A1(n4477), .A2(n4476), .ZN(n4478) );
  NOR2_X1 U5539 ( .A1(n5406), .A2(n4478), .ZN(n4479) );
  OR2_X1 U5540 ( .A1(n4498), .A2(n4479), .ZN(n5914) );
  OR2_X1 U5541 ( .A1(n6266), .A2(n4480), .ZN(n4481) );
  NAND2_X1 U5542 ( .A1(n4484), .A2(n6440), .ZN(n4496) );
  OR2_X1 U5543 ( .A1(n5481), .A2(n4486), .ZN(n4487) );
  NAND2_X1 U5544 ( .A1(n4485), .A2(n4487), .ZN(n5653) );
  INV_X1 U5545 ( .A(n4488), .ZN(n5971) );
  INV_X1 U5546 ( .A(n4489), .ZN(n5973) );
  NOR3_X1 U5547 ( .A1(n5973), .A2(n5770), .A3(n4490), .ZN(n4491) );
  AOI211_X1 U5548 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5971), .A(n4492), .B(n4491), .ZN(n4493) );
  NAND2_X1 U5549 ( .A1(n4496), .A2(n4495), .ZN(U2996) );
  AND2_X1 U5550 ( .A1(n4316), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4497)
         );
  AOI21_X1 U5551 ( .B1(n4499), .B2(EBX_REG_30__SCAN_IN), .A(n4497), .ZN(n4539)
         );
  AND2_X2 U5552 ( .A1(n4537), .A2(n4462), .ZN(n4535) );
  AOI21_X1 U5553 ( .B1(n4539), .B2(n4498), .A(n4535), .ZN(n4501) );
  OAI22_X1 U5554 ( .A1(n4499), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4316), .ZN(n4500) );
  XNOR2_X1 U5555 ( .A(n4501), .B(n4500), .ZN(n5904) );
  NOR2_X1 U5556 ( .A1(n4775), .A2(n4776), .ZN(n4602) );
  NAND2_X1 U5557 ( .A1(n4602), .A2(n6717), .ZN(n4606) );
  NAND2_X1 U5558 ( .A1(n4502), .A2(n4715), .ZN(n6720) );
  NAND3_X1 U5559 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_0__SCAN_IN), 
        .A3(n6747), .ZN(n4971) );
  INV_X1 U5560 ( .A(n5628), .ZN(n4504) );
  NAND2_X1 U5561 ( .A1(n4504), .A2(EBX_REG_31__SCAN_IN), .ZN(n4526) );
  NOR2_X1 U5562 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4510) );
  INV_X1 U5563 ( .A(n4510), .ZN(n5382) );
  NAND2_X1 U5564 ( .A1(n4329), .A2(n5382), .ZN(n4505) );
  NAND2_X1 U5565 ( .A1(n4287), .A2(n4713), .ZN(n4506) );
  NAND2_X1 U5566 ( .A1(n4316), .A2(n4506), .ZN(n4507) );
  NAND2_X1 U5567 ( .A1(n4507), .A2(n4510), .ZN(n4508) );
  INV_X1 U5568 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5850) );
  INV_X1 U5569 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6151) );
  INV_X1 U5570 ( .A(REIP_REG_11__SCAN_IN), .ZN(n5601) );
  INV_X1 U5571 ( .A(REIP_REG_10__SCAN_IN), .ZN(n5614) );
  INV_X1 U5572 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5636) );
  INV_X1 U5573 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6422) );
  INV_X1 U5574 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6235) );
  NOR3_X1 U5575 ( .A1(n5636), .A2(n6422), .A3(n6235), .ZN(n6187) );
  NAND3_X1 U5576 ( .A1(REIP_REG_4__SCAN_IN), .A2(REIP_REG_5__SCAN_IN), .A3(
        n6187), .ZN(n6182) );
  NOR2_X1 U5577 ( .A1(n6395), .A2(n6182), .ZN(n6171) );
  NAND3_X1 U5578 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        n6171), .ZN(n5612) );
  NOR4_X1 U5579 ( .A1(n5601), .A2(n5614), .A3(n6158), .A4(n5612), .ZN(n5593)
         );
  NAND2_X1 U5580 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5593), .ZN(n5585) );
  NOR3_X1 U5581 ( .A1(n5850), .A2(n6151), .A3(n5585), .ZN(n5554) );
  NAND2_X1 U5582 ( .A1(n6237), .A2(n5554), .ZN(n5575) );
  NAND2_X1 U5583 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n4511) );
  NOR2_X1 U5584 ( .A1(n5575), .A2(n4511), .ZN(n5541) );
  NAND2_X1 U5585 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5541), .ZN(n5530) );
  NAND2_X1 U5586 ( .A1(REIP_REG_18__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .ZN(
        n4509) );
  NOR2_X1 U5587 ( .A1(n5530), .A2(n4509), .ZN(n5503) );
  AND3_X1 U5588 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4516) );
  NAND2_X1 U5589 ( .A1(n5478), .A2(n4516), .ZN(n5456) );
  NAND3_X1 U5590 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4519) );
  NOR2_X1 U5591 ( .A1(n5456), .A2(n4519), .ZN(n5425) );
  NAND3_X1 U5592 ( .A1(n5425), .A2(REIP_REG_27__SCAN_IN), .A3(
        REIP_REG_28__SCAN_IN), .ZN(n5399) );
  INV_X1 U5593 ( .A(REIP_REG_30__SCAN_IN), .ZN(n4601) );
  INV_X1 U5594 ( .A(REIP_REG_29__SCAN_IN), .ZN(n5386) );
  NOR4_X1 U5595 ( .A1(n5399), .A2(REIP_REG_31__SCAN_IN), .A3(n4601), .A4(n5386), .ZN(n4528) );
  NAND2_X1 U5596 ( .A1(n4713), .A2(n4510), .ZN(n4812) );
  NAND2_X1 U5597 ( .A1(n4151), .A2(n4812), .ZN(n5384) );
  INV_X1 U5598 ( .A(n5554), .ZN(n4512) );
  NOR2_X1 U5599 ( .A1(n4512), .A2(n4511), .ZN(n4513) );
  AND2_X1 U5600 ( .A1(REIP_REG_17__SCAN_IN), .A2(n4513), .ZN(n4514) );
  AND2_X1 U5601 ( .A1(n6184), .A2(n4514), .ZN(n5527) );
  NAND4_X1 U5602 ( .A1(n5527), .A2(REIP_REG_20__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .A4(REIP_REG_19__SCAN_IN), .ZN(n4515) );
  NAND2_X1 U5603 ( .A1(n6186), .A2(n4515), .ZN(n5501) );
  INV_X1 U5604 ( .A(n4516), .ZN(n4517) );
  NAND2_X1 U5605 ( .A1(n6237), .A2(n4517), .ZN(n4518) );
  NAND2_X1 U5606 ( .A1(n5501), .A2(n4518), .ZN(n5467) );
  INV_X1 U5607 ( .A(n4519), .ZN(n4520) );
  NOR2_X1 U5608 ( .A1(n6253), .A2(n4520), .ZN(n4521) );
  AND2_X1 U5609 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4522) );
  NOR2_X1 U5610 ( .A1(n6144), .A2(n4522), .ZN(n4523) );
  NOR2_X1 U5611 ( .A1(n5436), .A2(n4523), .ZN(n5411) );
  OAI211_X1 U5612 ( .C1(REIP_REG_29__SCAN_IN), .C2(n6144), .A(n5411), .B(
        REIP_REG_30__SCAN_IN), .ZN(n5387) );
  NAND3_X1 U5613 ( .A1(n5387), .A2(REIP_REG_31__SCAN_IN), .A3(n6186), .ZN(
        n4525) );
  NAND2_X1 U5614 ( .A1(n6241), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4524)
         );
  OAI211_X1 U5615 ( .C1(n4526), .C2(n5384), .A(n4525), .B(n4524), .ZN(n4527)
         );
  AOI211_X1 U5616 ( .C1(n5904), .C2(n3100), .A(n4528), .B(n4527), .ZN(n4531)
         );
  NAND2_X1 U5617 ( .A1(n5376), .A2(n6204), .ZN(n4530) );
  NAND2_X1 U5618 ( .A1(n4531), .A2(n4530), .ZN(U2796) );
  NAND2_X1 U5619 ( .A1(n5726), .A2(n6262), .ZN(n4546) );
  INV_X1 U5620 ( .A(n4539), .ZN(n4536) );
  AOI211_X2 U5621 ( .C1(n5406), .C2(n4537), .A(n4536), .B(n4535), .ZN(n4542)
         );
  AOI211_X1 U5622 ( .C1(n4364), .C2(n4540), .A(n4539), .B(n4538), .ZN(n4541)
         );
  NOR2_X1 U5623 ( .A1(n4542), .A2(n4541), .ZN(n5381) );
  INV_X1 U5624 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5393) );
  NOR2_X1 U5625 ( .A1(n4544), .A2(n4543), .ZN(n4545) );
  NAND2_X1 U5626 ( .A1(n4546), .A2(n4545), .ZN(U2829) );
  INV_X1 U5627 ( .A(HOLD), .ZN(n6936) );
  NOR2_X1 U5628 ( .A1(n6936), .A2(n4573), .ZN(n4550) );
  INV_X1 U5629 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n4549) );
  NOR2_X1 U5630 ( .A1(n4555), .A2(n4549), .ZN(n4558) );
  NAND2_X1 U5631 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n4547) );
  OAI21_X1 U5632 ( .B1(n4550), .B2(n4558), .A(n4547), .ZN(n4548) );
  OAI211_X1 U5633 ( .C1(n4811), .C2(n4573), .A(n4548), .B(n4767), .ZN(U3182)
         );
  INV_X1 U5634 ( .A(n4551), .ZN(n4557) );
  AOI22_X1 U5635 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n4560) );
  NAND2_X2 U5636 ( .A1(n4555), .A2(STATE_REG_1__SCAN_IN), .ZN(n4598) );
  OAI21_X1 U5637 ( .B1(n4550), .B2(n4549), .A(n4598), .ZN(n4554) );
  INV_X1 U5638 ( .A(NA_N), .ZN(n6844) );
  NAND2_X1 U5639 ( .A1(n4551), .A2(n4555), .ZN(n4552) );
  AOI21_X1 U5640 ( .B1(n6844), .B2(STATE_REG_2__SCAN_IN), .A(n4552), .ZN(n4561) );
  INV_X1 U5641 ( .A(n4561), .ZN(n4553) );
  OAI211_X1 U5642 ( .C1(n4557), .C2(n4560), .A(n4554), .B(n4553), .ZN(U3181)
         );
  AOI221_X1 U5643 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n4811), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n4556) );
  AOI221_X1 U5644 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n4556), .C2(HOLD), .A(n4555), .ZN(n4562) );
  AOI21_X1 U5645 ( .B1(n6844), .B2(n4558), .A(n4557), .ZN(n4559) );
  OAI22_X1 U5646 ( .A1(n4562), .A2(n4561), .B1(n4560), .B2(n4559), .ZN(U3183)
         );
  INV_X1 U5647 ( .A(REIP_REG_4__SCAN_IN), .ZN(n7024) );
  NAND2_X1 U5648 ( .A1(n4563), .A2(n6752), .ZN(n4570) );
  INV_X1 U5649 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6882) );
  INV_X1 U5650 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n6862) );
  OAI222_X1 U5651 ( .A1(n4576), .A2(n7024), .B1(n4570), .B2(n6882), .C1(n6862), 
        .C2(n6752), .ZN(U3187) );
  INV_X1 U5652 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5512) );
  INV_X1 U5653 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n6861) );
  INV_X1 U5654 ( .A(REIP_REG_20__SCAN_IN), .ZN(n4588) );
  OAI222_X1 U5655 ( .A1(n4576), .A2(n5512), .B1(n6752), .B2(n6861), .C1(n4570), 
        .C2(n4588), .ZN(U3202) );
  INV_X1 U5656 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5596) );
  INV_X1 U5657 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n6873) );
  OAI222_X1 U5658 ( .A1(n4576), .A2(n5596), .B1(n4570), .B2(n6151), .C1(n6873), 
        .C2(n6752), .ZN(U3195) );
  INV_X1 U5659 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5562) );
  INV_X1 U5660 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6910) );
  INV_X1 U5661 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5574) );
  OAI222_X1 U5662 ( .A1(n4570), .A2(n5562), .B1(n6752), .B2(n6910), .C1(n4576), 
        .C2(n5574), .ZN(U3198) );
  INV_X2 U5663 ( .A(n4570), .ZN(n4599) );
  AOI22_X1 U5664 ( .A1(n4599), .A2(REIP_REG_10__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_8__SCAN_IN), .ZN(n4564) );
  OAI21_X1 U5665 ( .B1(n6158), .B2(n4576), .A(n4564), .ZN(U3192) );
  AOI22_X1 U5666 ( .A1(n4599), .A2(REIP_REG_14__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_12__SCAN_IN), .ZN(n4565) );
  OAI21_X1 U5667 ( .B1(n6151), .B2(n4576), .A(n4565), .ZN(U3196) );
  AOI22_X1 U5668 ( .A1(n4599), .A2(REIP_REG_12__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_10__SCAN_IN), .ZN(n4566) );
  OAI21_X1 U5669 ( .B1(n5601), .B2(n4576), .A(n4566), .ZN(U3194) );
  INV_X1 U5670 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6974) );
  AOI22_X1 U5671 ( .A1(n4599), .A2(REIP_REG_9__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_7__SCAN_IN), .ZN(n4567) );
  OAI21_X1 U5672 ( .B1(n6974), .B2(n4576), .A(n4567), .ZN(U3191) );
  AOI22_X1 U5673 ( .A1(n4599), .A2(REIP_REG_6__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_4__SCAN_IN), .ZN(n4568) );
  OAI21_X1 U5674 ( .B1(n6882), .B2(n4576), .A(n4568), .ZN(U3188) );
  INV_X1 U5675 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6198) );
  AOI22_X1 U5676 ( .A1(n4599), .A2(REIP_REG_8__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_6__SCAN_IN), .ZN(n4569) );
  OAI21_X1 U5677 ( .B1(n6198), .B2(n4576), .A(n4569), .ZN(U3190) );
  INV_X1 U5678 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5435) );
  INV_X1 U5679 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6940) );
  OAI222_X1 U5680 ( .A1(n4570), .A2(n5435), .B1(n6752), .B2(n6940), .C1(n5454), 
        .C2(n4576), .ZN(U3207) );
  AOI22_X1 U5681 ( .A1(n4599), .A2(REIP_REG_4__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_2__SCAN_IN), .ZN(n4571) );
  OAI21_X1 U5682 ( .B1(n6422), .B2(n4576), .A(n4571), .ZN(U3186) );
  AOI22_X1 U5683 ( .A1(n4599), .A2(REIP_REG_3__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_1__SCAN_IN), .ZN(n4572) );
  OAI21_X1 U5684 ( .B1(n6235), .B2(n4576), .A(n4572), .ZN(U3185) );
  INV_X1 U5685 ( .A(ADS_N_REG_SCAN_IN), .ZN(n4575) );
  OAI21_X1 U5686 ( .B1(n4573), .B2(STATE_REG_2__SCAN_IN), .A(
        STATE_REG_0__SCAN_IN), .ZN(n4574) );
  OAI21_X1 U5687 ( .B1(n6752), .B2(n4575), .A(n6726), .ZN(U2789) );
  AOI22_X1 U5688 ( .A1(n4599), .A2(REIP_REG_11__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_9__SCAN_IN), .ZN(n4577) );
  OAI21_X1 U5689 ( .B1(n5614), .B2(n4576), .A(n4577), .ZN(U3193) );
  AOI22_X1 U5690 ( .A1(n4599), .A2(REIP_REG_2__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_0__SCAN_IN), .ZN(n4578) );
  OAI21_X1 U5691 ( .B1(n5636), .B2(n4576), .A(n4578), .ZN(U3184) );
  AOI22_X1 U5692 ( .A1(n4599), .A2(REIP_REG_7__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_5__SCAN_IN), .ZN(n4579) );
  OAI21_X1 U5693 ( .B1(n6395), .B2(n4576), .A(n4579), .ZN(U3189) );
  INV_X1 U5694 ( .A(REIP_REG_23__SCAN_IN), .ZN(n4581) );
  AOI22_X1 U5695 ( .A1(n4599), .A2(REIP_REG_24__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_22__SCAN_IN), .ZN(n4580) );
  OAI21_X1 U5696 ( .B1(n4581), .B2(n4576), .A(n4580), .ZN(U3206) );
  AOI22_X1 U5697 ( .A1(n4599), .A2(REIP_REG_15__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_13__SCAN_IN), .ZN(n4582) );
  OAI21_X1 U5698 ( .B1(n5850), .B2(n4576), .A(n4582), .ZN(U3197) );
  AOI22_X1 U5699 ( .A1(n4599), .A2(REIP_REG_17__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_15__SCAN_IN), .ZN(n4583) );
  OAI21_X1 U5700 ( .B1(n5562), .B2(n4576), .A(n4583), .ZN(U3199) );
  INV_X1 U5701 ( .A(REIP_REG_17__SCAN_IN), .ZN(n4585) );
  AOI22_X1 U5702 ( .A1(n4599), .A2(REIP_REG_18__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_16__SCAN_IN), .ZN(n4584) );
  OAI21_X1 U5703 ( .B1(n4585), .B2(n4576), .A(n4584), .ZN(U3200) );
  INV_X1 U5704 ( .A(REIP_REG_18__SCAN_IN), .ZN(n5816) );
  AOI22_X1 U5705 ( .A1(n4599), .A2(REIP_REG_19__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_17__SCAN_IN), .ZN(n4586) );
  OAI21_X1 U5706 ( .B1(n5816), .B2(n4576), .A(n4586), .ZN(U3201) );
  AOI22_X1 U5707 ( .A1(n4599), .A2(REIP_REG_21__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_19__SCAN_IN), .ZN(n4587) );
  OAI21_X1 U5708 ( .B1(n4588), .B2(n4576), .A(n4587), .ZN(U3203) );
  INV_X1 U5709 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5795) );
  AOI22_X1 U5710 ( .A1(n4599), .A2(REIP_REG_22__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_20__SCAN_IN), .ZN(n4589) );
  OAI21_X1 U5711 ( .B1(n5795), .B2(n4576), .A(n4589), .ZN(U3204) );
  AOI22_X1 U5712 ( .A1(n4599), .A2(REIP_REG_23__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_21__SCAN_IN), .ZN(n4590) );
  OAI21_X1 U5713 ( .B1(n5472), .B2(n4576), .A(n4590), .ZN(U3205) );
  INV_X1 U5714 ( .A(REIP_REG_27__SCAN_IN), .ZN(n5424) );
  AOI22_X1 U5715 ( .A1(n4599), .A2(REIP_REG_28__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_26__SCAN_IN), .ZN(n4591) );
  OAI21_X1 U5716 ( .B1(n5424), .B2(n4576), .A(n4591), .ZN(U3210) );
  AOI22_X1 U5717 ( .A1(n4599), .A2(REIP_REG_26__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_24__SCAN_IN), .ZN(n4592) );
  OAI21_X1 U5718 ( .B1(n5435), .B2(n4576), .A(n4592), .ZN(U3208) );
  INV_X1 U5719 ( .A(REIP_REG_26__SCAN_IN), .ZN(n4594) );
  AOI22_X1 U5720 ( .A1(n4599), .A2(REIP_REG_27__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_25__SCAN_IN), .ZN(n4593) );
  OAI21_X1 U5721 ( .B1(n4594), .B2(n4576), .A(n4593), .ZN(U3209) );
  AOI22_X1 U5722 ( .A1(n4599), .A2(REIP_REG_30__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_28__SCAN_IN), .ZN(n4595) );
  OAI21_X1 U5723 ( .B1(n5386), .B2(n4576), .A(n4595), .ZN(U3212) );
  INV_X1 U5724 ( .A(REIP_REG_28__SCAN_IN), .ZN(n4597) );
  AOI22_X1 U5725 ( .A1(n4599), .A2(REIP_REG_29__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_27__SCAN_IN), .ZN(n4596) );
  OAI21_X1 U5726 ( .B1(n4597), .B2(n4576), .A(n4596), .ZN(U3211) );
  AOI22_X1 U5727 ( .A1(n4599), .A2(REIP_REG_31__SCAN_IN), .B1(n4598), .B2(
        ADDRESS_REG_29__SCAN_IN), .ZN(n4600) );
  OAI21_X1 U5728 ( .B1(n4601), .B2(n4576), .A(n4600), .ZN(U3213) );
  NOR2_X1 U5729 ( .A1(n6655), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5513) );
  INV_X1 U5730 ( .A(n5513), .ZN(n4604) );
  INV_X1 U5731 ( .A(n4281), .ZN(n4770) );
  OAI22_X1 U5732 ( .A1(n4772), .A2(n4839), .B1(n4770), .B2(n4602), .ZN(n4769)
         );
  INV_X1 U5733 ( .A(n6717), .ZN(n4973) );
  OAI21_X1 U5734 ( .B1(n4769), .B2(n4973), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n4603) );
  OAI21_X1 U5735 ( .B1(n4604), .B2(n4872), .A(n4603), .ZN(U2790) );
  AOI211_X1 U5736 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4606), .A(n5513), .B(
        n4610), .ZN(n4607) );
  INV_X1 U5737 ( .A(n4607), .ZN(U2788) );
  INV_X1 U5738 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4612) );
  NAND2_X1 U5739 ( .A1(n4610), .A2(n4811), .ZN(n4608) );
  NAND2_X1 U5740 ( .A1(n6319), .A2(UWORD_REG_6__SCAN_IN), .ZN(n4611) );
  INV_X1 U5741 ( .A(DATAI_6_), .ZN(n4920) );
  OR2_X1 U5742 ( .A1(n6308), .A2(n4920), .ZN(n4613) );
  OAI211_X1 U5743 ( .C1(n6310), .C2(n4612), .A(n4611), .B(n4613), .ZN(U2930)
         );
  NAND2_X1 U5744 ( .A1(n6319), .A2(LWORD_REG_6__SCAN_IN), .ZN(n4614) );
  OAI211_X1 U5745 ( .C1(n6310), .C2(n5066), .A(n4614), .B(n4613), .ZN(U2945)
         );
  INV_X1 U5746 ( .A(n4615), .ZN(n4616) );
  NOR2_X1 U5747 ( .A1(n4283), .A2(n4616), .ZN(n4617) );
  AOI21_X1 U5748 ( .B1(n4772), .B2(n4665), .A(n4617), .ZN(n4842) );
  NAND2_X1 U5749 ( .A1(n5367), .A2(n4713), .ZN(n4619) );
  AOI21_X1 U5750 ( .B1(n4619), .B2(n4281), .A(n4618), .ZN(n4625) );
  NAND2_X1 U5751 ( .A1(n4621), .A2(n4620), .ZN(n4622) );
  NAND2_X1 U5752 ( .A1(n4623), .A2(n4622), .ZN(n4624) );
  AOI21_X1 U5753 ( .B1(n4772), .B2(n4625), .A(n4624), .ZN(n4627) );
  NAND3_X1 U5754 ( .A1(n4842), .A2(n4627), .A3(n4626), .ZN(n4797) );
  INV_X1 U5755 ( .A(n4797), .ZN(n4629) );
  INV_X1 U5756 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6872) );
  NAND2_X1 U5757 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .ZN(n4874) );
  INV_X1 U5758 ( .A(n4874), .ZN(n4628) );
  NAND2_X1 U5759 ( .A1(n4628), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6723) );
  OAI22_X1 U5760 ( .A1(n4629), .A2(n4973), .B1(n6872), .B2(n6723), .ZN(n4632)
         );
  NAND2_X1 U5761 ( .A1(n4872), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4816) );
  INV_X1 U5762 ( .A(n4816), .ZN(n4899) );
  INV_X1 U5763 ( .A(n6125), .ZN(n4635) );
  INV_X1 U5764 ( .A(n4283), .ZN(n4764) );
  INV_X1 U5765 ( .A(n4937), .ZN(n6658) );
  NOR2_X1 U5766 ( .A1(n4630), .A2(n6658), .ZN(n4631) );
  XNOR2_X1 U5767 ( .A(n4631), .B(n4634), .ZN(n6221) );
  NAND4_X1 U5768 ( .A1(n4632), .A2(n4764), .A3(n6119), .A4(n6221), .ZN(n4633)
         );
  OAI21_X1 U5769 ( .B1(n4635), .B2(n4634), .A(n4633), .ZN(U3455) );
  AOI222_X1 U5770 ( .A1(n6319), .A2(LWORD_REG_15__SCAN_IN), .B1(n6304), .B2(
        DATAI_15_), .C1(EAX_REG_15__SCAN_IN), .C2(n6323), .ZN(n4636) );
  INV_X1 U5771 ( .A(n4636), .ZN(U2954) );
  NAND2_X1 U5772 ( .A1(n6319), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4637) );
  NAND2_X1 U5773 ( .A1(n6304), .A2(DATAI_2_), .ZN(n4644) );
  OAI211_X1 U5774 ( .C1(n6310), .C2(n4638), .A(n4637), .B(n4644), .ZN(U2926)
         );
  INV_X1 U5775 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4640) );
  NAND2_X1 U5776 ( .A1(n6319), .A2(LWORD_REG_7__SCAN_IN), .ZN(n4639) );
  NAND2_X1 U5777 ( .A1(n6304), .A2(DATAI_7_), .ZN(n4641) );
  OAI211_X1 U5778 ( .C1(n6310), .C2(n4640), .A(n4639), .B(n4641), .ZN(U2946)
         );
  NAND2_X1 U5779 ( .A1(n6319), .A2(UWORD_REG_7__SCAN_IN), .ZN(n4642) );
  OAI211_X1 U5780 ( .C1(n6310), .C2(n4643), .A(n4642), .B(n4641), .ZN(U2931)
         );
  INV_X1 U5781 ( .A(EAX_REG_2__SCAN_IN), .ZN(n4646) );
  NAND2_X1 U5782 ( .A1(n6319), .A2(LWORD_REG_2__SCAN_IN), .ZN(n4645) );
  OAI211_X1 U5783 ( .C1(n6310), .C2(n4646), .A(n4645), .B(n4644), .ZN(U2941)
         );
  INV_X1 U5784 ( .A(LWORD_REG_1__SCAN_IN), .ZN(n4648) );
  INV_X1 U5785 ( .A(DATAI_1_), .ZN(n4913) );
  NOR2_X1 U5786 ( .A1(n6308), .A2(n4913), .ZN(n4680) );
  AOI21_X1 U5787 ( .B1(n6323), .B2(EAX_REG_1__SCAN_IN), .A(n4680), .ZN(n4647)
         );
  OAI21_X1 U5788 ( .B1(n6325), .B2(n4648), .A(n4647), .ZN(U2940) );
  INV_X1 U5789 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n4650) );
  INV_X1 U5790 ( .A(DATAI_4_), .ZN(n4904) );
  NOR2_X1 U5791 ( .A1(n6308), .A2(n4904), .ZN(n4682) );
  AOI21_X1 U5792 ( .B1(n6323), .B2(EAX_REG_4__SCAN_IN), .A(n4682), .ZN(n4649)
         );
  OAI21_X1 U5793 ( .B1(n6325), .B2(n4650), .A(n4649), .ZN(U2943) );
  INV_X1 U5794 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n4652) );
  INV_X1 U5795 ( .A(DATAI_5_), .ZN(n4898) );
  NOR2_X1 U5796 ( .A1(n6308), .A2(n4898), .ZN(n4686) );
  AOI21_X1 U5797 ( .B1(n6323), .B2(EAX_REG_5__SCAN_IN), .A(n4686), .ZN(n4651)
         );
  OAI21_X1 U5798 ( .B1(n6325), .B2(n4652), .A(n4651), .ZN(U2944) );
  INV_X1 U5799 ( .A(LWORD_REG_9__SCAN_IN), .ZN(n4654) );
  INV_X1 U5800 ( .A(DATAI_9_), .ZN(n6892) );
  NOR2_X1 U5801 ( .A1(n6308), .A2(n6892), .ZN(n4684) );
  AOI21_X1 U5802 ( .B1(n6323), .B2(EAX_REG_9__SCAN_IN), .A(n4684), .ZN(n4653)
         );
  OAI21_X1 U5803 ( .B1(n6325), .B2(n4654), .A(n4653), .ZN(U2948) );
  INV_X1 U5804 ( .A(LWORD_REG_3__SCAN_IN), .ZN(n4656) );
  INV_X1 U5805 ( .A(DATAI_3_), .ZN(n4908) );
  NOR2_X1 U5806 ( .A1(n6308), .A2(n4908), .ZN(n4657) );
  AOI21_X1 U5807 ( .B1(n6323), .B2(EAX_REG_3__SCAN_IN), .A(n4657), .ZN(n4655)
         );
  OAI21_X1 U5808 ( .B1(n6325), .B2(n4656), .A(n4655), .ZN(U2942) );
  INV_X1 U5809 ( .A(UWORD_REG_3__SCAN_IN), .ZN(n4659) );
  AOI21_X1 U5810 ( .B1(n6323), .B2(EAX_REG_19__SCAN_IN), .A(n4657), .ZN(n4658)
         );
  OAI21_X1 U5811 ( .B1(n6325), .B2(n4659), .A(n4658), .ZN(U2927) );
  INV_X1 U5812 ( .A(n4661), .ZN(n4664) );
  AND4_X1 U5813 ( .A1(n3426), .A2(n4283), .A3(n4662), .A4(n4273), .ZN(n4663)
         );
  NAND2_X1 U5814 ( .A1(n4664), .A2(n4663), .ZN(n4787) );
  NAND2_X1 U5815 ( .A1(n3104), .A2(n4787), .ZN(n4672) );
  INV_X1 U5816 ( .A(n4665), .ZN(n4666) );
  NAND2_X1 U5817 ( .A1(n4773), .A2(n4666), .ZN(n4747) );
  XNOR2_X1 U5818 ( .A(n4677), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4670)
         );
  XNOR2_X1 U5819 ( .A(n3268), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4667)
         );
  NAND2_X1 U5820 ( .A1(n5367), .A2(n4667), .ZN(n4668) );
  OAI21_X1 U5821 ( .B1(n4670), .B2(n4749), .A(n4668), .ZN(n4669) );
  AOI21_X1 U5822 ( .B1(n4747), .B2(n4670), .A(n4669), .ZN(n4671) );
  NAND2_X1 U5823 ( .A1(n4672), .A2(n4671), .ZN(n4758) );
  INV_X1 U5824 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n7051) );
  OAI22_X1 U5825 ( .A1(n4673), .A2(n7051), .B1(INSTADDRPOINTER_REG_31__SCAN_IN), .B2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6112) );
  INV_X1 U5826 ( .A(n6112), .ZN(n4674) );
  AND3_X1 U5827 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n4674), .A3(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4676) );
  INV_X1 U5828 ( .A(n4677), .ZN(n4789) );
  NOR3_X1 U5829 ( .A1(n6121), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n4789), 
        .ZN(n4675) );
  AOI211_X1 U5830 ( .C1(n6119), .C2(n4758), .A(n4676), .B(n4675), .ZN(n4679)
         );
  NOR2_X1 U5831 ( .A1(n6121), .A2(n4677), .ZN(n6111) );
  OAI21_X1 U5832 ( .B1(n6125), .B2(n6111), .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .ZN(n4678) );
  OAI21_X1 U5833 ( .B1(n6125), .B2(n4679), .A(n4678), .ZN(U3459) );
  INV_X1 U5834 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n4727) );
  AOI21_X1 U5835 ( .B1(n6323), .B2(EAX_REG_17__SCAN_IN), .A(n4680), .ZN(n4681)
         );
  OAI21_X1 U5836 ( .B1(n4727), .B2(n6325), .A(n4681), .ZN(U2925) );
  INV_X1 U5837 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n4721) );
  AOI21_X1 U5838 ( .B1(n6323), .B2(EAX_REG_20__SCAN_IN), .A(n4682), .ZN(n4683)
         );
  OAI21_X1 U5839 ( .B1(n4721), .B2(n6325), .A(n4683), .ZN(U2928) );
  INV_X1 U5840 ( .A(UWORD_REG_9__SCAN_IN), .ZN(n4724) );
  AOI21_X1 U5841 ( .B1(n6323), .B2(EAX_REG_25__SCAN_IN), .A(n4684), .ZN(n4685)
         );
  OAI21_X1 U5842 ( .B1(n4724), .B2(n6325), .A(n4685), .ZN(U2933) );
  INV_X1 U5843 ( .A(UWORD_REG_5__SCAN_IN), .ZN(n4688) );
  AOI21_X1 U5844 ( .B1(n6323), .B2(EAX_REG_21__SCAN_IN), .A(n4686), .ZN(n4687)
         );
  OAI21_X1 U5845 ( .B1(n4688), .B2(n6325), .A(n4687), .ZN(U2929) );
  INV_X1 U5846 ( .A(LWORD_REG_0__SCAN_IN), .ZN(n4690) );
  INV_X1 U5847 ( .A(EAX_REG_0__SCAN_IN), .ZN(n4689) );
  OAI222_X1 U5848 ( .A1(n4690), .A2(n6325), .B1(n6308), .B2(n4924), .C1(n4689), 
        .C2(n6310), .ZN(U2939) );
  XNOR2_X1 U5849 ( .A(n4691), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4709)
         );
  INV_X1 U5850 ( .A(n4692), .ZN(n4693) );
  AOI21_X1 U5851 ( .B1(n4694), .B2(n4392), .A(n4693), .ZN(n6250) );
  INV_X1 U5852 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6891) );
  NOR2_X1 U5853 ( .A1(n6423), .A2(n6891), .ZN(n4707) );
  AOI211_X1 U5854 ( .C1(n6435), .C2(n6250), .A(n4707), .B(n4695), .ZN(n4699)
         );
  INV_X1 U5855 ( .A(n6044), .ZN(n4696) );
  OAI21_X1 U5856 ( .B1(n4697), .B2(n4696), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4698) );
  OAI211_X1 U5857 ( .C1(n4709), .C2(n6412), .A(n4699), .B(n4698), .ZN(U3018)
         );
  OR2_X1 U5858 ( .A1(n4701), .A2(n4700), .ZN(n4702) );
  OAI21_X1 U5859 ( .B1(n6354), .B2(n4704), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4705) );
  INV_X1 U5860 ( .A(n4705), .ZN(n4706) );
  AOI211_X1 U5861 ( .C1(n6256), .C2(n6349), .A(n4707), .B(n4706), .ZN(n4708)
         );
  OAI21_X1 U5862 ( .B1(n4709), .B2(n6334), .A(n4708), .ZN(U2986) );
  INV_X1 U5863 ( .A(n5367), .ZN(n4710) );
  NAND2_X1 U5864 ( .A1(n6295), .A2(DATAO_REG_26__SCAN_IN), .ZN(n4717) );
  NAND2_X1 U5865 ( .A1(n6744), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4716) );
  OAI211_X1 U5866 ( .C1(n4729), .C2(n3981), .A(n4717), .B(n4716), .ZN(U2897)
         );
  INV_X1 U5867 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4720) );
  NAND2_X1 U5868 ( .A1(n6295), .A2(DATAO_REG_28__SCAN_IN), .ZN(n4719) );
  NAND2_X1 U5869 ( .A1(n6744), .A2(UWORD_REG_12__SCAN_IN), .ZN(n4718) );
  OAI211_X1 U5870 ( .C1(n4729), .C2(n4720), .A(n4719), .B(n4718), .ZN(U2895)
         );
  INV_X1 U5871 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n4723) );
  INV_X1 U5872 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4722) );
  INV_X1 U5873 ( .A(n6744), .ZN(n6280) );
  OAI222_X1 U5874 ( .A1(n4723), .A2(n6285), .B1(n4729), .B2(n4722), .C1(n6280), 
        .C2(n4721), .ZN(U2903) );
  INV_X1 U5875 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n4726) );
  OAI222_X1 U5876 ( .A1(n4726), .A2(n6285), .B1(n4729), .B2(n4725), .C1(n6280), 
        .C2(n4724), .ZN(U2898) );
  INV_X1 U5877 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4730) );
  INV_X1 U5878 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4728) );
  OAI222_X1 U5879 ( .A1(n4730), .A2(n6285), .B1(n4729), .B2(n4728), .C1(n6280), 
        .C2(n4727), .ZN(U2906) );
  XNOR2_X1 U5880 ( .A(n4731), .B(n4732), .ZN(n4822) );
  OAI21_X1 U5881 ( .B1(n4735), .B2(n4734), .A(n4733), .ZN(n5642) );
  INV_X1 U5882 ( .A(n5642), .ZN(n4738) );
  AOI22_X1 U5883 ( .A1(n6354), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6433), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4736) );
  OAI21_X1 U5884 ( .B1(n6363), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4736), 
        .ZN(n4737) );
  AOI21_X1 U5885 ( .B1(n4738), .B2(n6349), .A(n4737), .ZN(n4739) );
  OAI21_X1 U5886 ( .B1(n4822), .B2(n6334), .A(n4739), .ZN(U2985) );
  INV_X1 U5887 ( .A(n6256), .ZN(n4849) );
  AOI22_X1 U5888 ( .A1(n6261), .A2(n6250), .B1(EBX_REG_0__SCAN_IN), .B2(n5659), 
        .ZN(n4740) );
  OAI21_X1 U5889 ( .B1(n4849), .B2(n5670), .A(n4740), .ZN(U2859) );
  AOI222_X1 U5890 ( .A1(n6295), .A2(DATAO_REG_30__SCAN_IN), .B1(n6272), .B2(
        EAX_REG_30__SCAN_IN), .C1(n6744), .C2(UWORD_REG_14__SCAN_IN), .ZN(
        n4741) );
  INV_X1 U5891 ( .A(n4741), .ZN(U2893) );
  NAND2_X1 U5892 ( .A1(n4743), .A2(n4787), .ZN(n4757) );
  AOI21_X1 U5893 ( .B1(n4789), .B2(n4744), .A(n4745), .ZN(n4746) );
  NAND3_X1 U5894 ( .A1(n4747), .A2(n4746), .A3(n3468), .ZN(n4755) );
  NAND2_X1 U5895 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n6756), .ZN(n4748) );
  INV_X1 U5896 ( .A(n4748), .ZN(n4751) );
  MUX2_X1 U5897 ( .A(n4751), .B(n4748), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4753) );
  INV_X1 U5898 ( .A(n4749), .ZN(n4752) );
  OAI211_X1 U5899 ( .C1(n4751), .C2(n3246), .A(n3362), .B(n4750), .ZN(n6120)
         );
  AOI22_X1 U5900 ( .A1(n5367), .A2(n4753), .B1(n4752), .B2(n6120), .ZN(n4754)
         );
  AND2_X1 U5901 ( .A1(n4755), .A2(n4754), .ZN(n4756) );
  NAND2_X1 U5902 ( .A1(n4757), .A2(n4756), .ZN(n6118) );
  MUX2_X1 U5903 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6118), .S(n4797), 
        .Z(n4807) );
  MUX2_X1 U5904 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n4758), .S(n4797), 
        .Z(n4802) );
  NAND3_X1 U5905 ( .A1(n4807), .A2(n5369), .A3(n4802), .ZN(n4761) );
  NAND2_X1 U5906 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6872), .ZN(n4762) );
  INV_X1 U5907 ( .A(n4762), .ZN(n4759) );
  NAND2_X1 U5908 ( .A1(n4745), .A2(n4759), .ZN(n4760) );
  OAI21_X1 U5909 ( .B1(n4797), .B2(STATE2_REG_1__SCAN_IN), .A(n4762), .ZN(
        n4763) );
  NAND2_X1 U5910 ( .A1(n4763), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4766) );
  NAND3_X1 U5911 ( .A1(n6221), .A2(n4764), .A3(n5369), .ZN(n4765) );
  NAND2_X1 U5912 ( .A1(n4766), .A2(n4765), .ZN(n4875) );
  NAND3_X1 U5913 ( .A1(n3402), .A2(n4767), .A3(n4316), .ZN(n4768) );
  AND2_X1 U5914 ( .A1(n4768), .A2(n4811), .ZN(n6745) );
  OR2_X1 U5915 ( .A1(n4769), .A2(n6745), .ZN(n6130) );
  NOR2_X1 U5916 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n4781) );
  NOR2_X1 U5917 ( .A1(n4771), .A2(n4770), .ZN(n4774) );
  MUX2_X1 U5918 ( .A(n4774), .B(n4773), .S(n4772), .Z(n4779) );
  INV_X1 U5919 ( .A(n4775), .ZN(n4777) );
  NAND2_X1 U5920 ( .A1(n4777), .A2(n4776), .ZN(n4778) );
  AND2_X1 U5921 ( .A1(n4779), .A2(n4778), .ZN(n6739) );
  OAI211_X1 U5922 ( .C1(n6130), .C2(n4781), .A(n6739), .B(n4780), .ZN(n4782)
         );
  NOR2_X1 U5923 ( .A1(n4875), .A2(n4782), .ZN(n4810) );
  NOR2_X1 U5924 ( .A1(n4792), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4783)
         );
  AOI21_X1 U5925 ( .B1(n3114), .B2(n4787), .A(n4783), .ZN(n5368) );
  AOI21_X1 U5926 ( .B1(n5367), .B2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(n6651), 
        .ZN(n4784) );
  AND2_X1 U5927 ( .A1(n5368), .A2(n4784), .ZN(n4800) );
  NAND2_X1 U5928 ( .A1(n4802), .A2(n4785), .ZN(n4799) );
  NAND2_X1 U5929 ( .A1(n4786), .A2(n4787), .ZN(n4795) );
  INV_X1 U5930 ( .A(n4788), .ZN(n4790) );
  NAND2_X1 U5931 ( .A1(n4790), .A2(n4789), .ZN(n4791) );
  NOR2_X1 U5932 ( .A1(n4792), .A2(n4791), .ZN(n4793) );
  AOI21_X1 U5933 ( .B1(n5367), .B2(n3268), .A(n4793), .ZN(n4794) );
  NAND2_X1 U5934 ( .A1(n4795), .A2(n4794), .ZN(n6113) );
  NAND2_X1 U5935 ( .A1(n4800), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4796) );
  NAND3_X1 U5936 ( .A1(n4797), .A2(n6113), .A3(n4796), .ZN(n4798) );
  OAI211_X1 U5937 ( .C1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n4800), .A(n4799), .B(n4798), .ZN(n4806) );
  INV_X1 U5938 ( .A(n4807), .ZN(n4801) );
  NAND2_X1 U5939 ( .A1(n4801), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4805) );
  INV_X1 U5940 ( .A(n4802), .ZN(n4803) );
  AOI21_X1 U5941 ( .B1(n4803), .B2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4804) );
  NAND3_X1 U5942 ( .A1(n4806), .A2(n4805), .A3(n4804), .ZN(n4809) );
  INV_X1 U5943 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n7040) );
  NAND3_X1 U5944 ( .A1(n4807), .A2(n7040), .A3(n6781), .ZN(n4808) );
  NAND4_X1 U5945 ( .A1(n4870), .A2(n4810), .A3(n4809), .A4(n4808), .ZN(n4965)
         );
  OAI22_X1 U5946 ( .A1(n4965), .A2(n4973), .B1(n4811), .B2(n6280), .ZN(n4815)
         );
  OR2_X1 U5947 ( .A1(n4813), .A2(n4812), .ZN(n4814) );
  OAI211_X1 U5948 ( .C1(n4967), .C2(n5072), .A(n4816), .B(n6723), .ZN(U3453)
         );
  INV_X1 U5949 ( .A(n6394), .ZN(n6368) );
  OR2_X1 U5950 ( .A1(n6368), .A2(n4817), .ZN(n4818) );
  MUX2_X1 U5951 ( .A(n4818), .B(n6391), .S(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .Z(n4821) );
  XNOR2_X1 U5952 ( .A(n4819), .B(n4329), .ZN(n4823) );
  AOI22_X1 U5953 ( .A1(n6435), .A2(n4823), .B1(n6433), .B2(REIP_REG_1__SCAN_IN), .ZN(n4820) );
  OAI211_X1 U5954 ( .C1(n4822), .C2(n6412), .A(n4821), .B(n4820), .ZN(U3017)
         );
  INV_X1 U5955 ( .A(n4823), .ZN(n4824) );
  OAI222_X1 U5956 ( .A1(n4824), .A2(n5672), .B1(n5638), .B2(n6266), .C1(n5642), 
        .C2(n5670), .ZN(U2858) );
  INV_X1 U5957 ( .A(n4825), .ZN(n4831) );
  NOR2_X1 U5958 ( .A1(n4733), .A2(n3644), .ZN(n4828) );
  OR2_X1 U5959 ( .A1(n4828), .A2(n4827), .ZN(n4830) );
  NAND2_X1 U5960 ( .A1(n4733), .A2(n3644), .ZN(n4829) );
  AOI21_X1 U5961 ( .B1(n4831), .B2(n4733), .A(n4859), .ZN(n6359) );
  INV_X1 U5962 ( .A(n6359), .ZN(n4850) );
  OAI21_X1 U5963 ( .B1(n4834), .B2(n4833), .A(n4832), .ZN(n6432) );
  OAI222_X1 U5964 ( .A1(n4850), .A2(n5670), .B1(n4835), .B2(n6266), .C1(n5672), 
        .C2(n6432), .ZN(U2857) );
  AOI222_X1 U5965 ( .A1(EAX_REG_21__SCAN_IN), .A2(n6272), .B1(n6295), .B2(
        DATAO_REG_21__SCAN_IN), .C1(n6744), .C2(UWORD_REG_5__SCAN_IN), .ZN(
        n4836) );
  INV_X1 U5966 ( .A(n4836), .ZN(U2902) );
  AOI222_X1 U5967 ( .A1(EAX_REG_29__SCAN_IN), .A2(n6272), .B1(n6295), .B2(
        DATAO_REG_29__SCAN_IN), .C1(n6744), .C2(UWORD_REG_13__SCAN_IN), .ZN(
        n4837) );
  INV_X1 U5968 ( .A(n4837), .ZN(U2894) );
  AOI222_X1 U5969 ( .A1(EAX_REG_27__SCAN_IN), .A2(n6272), .B1(n6295), .B2(
        DATAO_REG_27__SCAN_IN), .C1(n6744), .C2(UWORD_REG_11__SCAN_IN), .ZN(
        n4838) );
  INV_X1 U5970 ( .A(n4838), .ZN(U2896) );
  NAND3_X1 U5971 ( .A1(n4840), .A2(n4909), .A3(n4839), .ZN(n4841) );
  NAND2_X1 U5972 ( .A1(n4842), .A2(n4841), .ZN(n4843) );
  AND2_X1 U5973 ( .A1(n3410), .A2(n3585), .ZN(n4848) );
  INV_X1 U5974 ( .A(n4848), .ZN(n4846) );
  AND2_X1 U5975 ( .A1(n4846), .A2(n4845), .ZN(n4847) );
  AND2_X1 U5976 ( .A1(n5715), .A2(n3392), .ZN(n5711) );
  INV_X1 U5977 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6855) );
  OAI222_X1 U5978 ( .A1(n5642), .A2(n5721), .B1(n5716), .B2(n4913), .C1(n5715), 
        .C2(n6855), .ZN(U2890) );
  OAI222_X1 U5979 ( .A1(n4849), .A2(n5721), .B1(n5716), .B2(n4924), .C1(n5715), 
        .C2(n4689), .ZN(U2891) );
  INV_X1 U5980 ( .A(DATAI_2_), .ZN(n6822) );
  OAI222_X1 U5981 ( .A1(n4850), .A2(n5721), .B1(n5716), .B2(n6822), .C1(n5715), 
        .C2(n4646), .ZN(U2889) );
  AOI21_X1 U5982 ( .B1(n4859), .B2(n4852), .A(n4853), .ZN(n4854) );
  AND2_X1 U5983 ( .A1(n4881), .A2(n4856), .ZN(n4857) );
  NOR2_X1 U5984 ( .A1(n4855), .A2(n4857), .ZN(n6414) );
  INV_X1 U5985 ( .A(n6414), .ZN(n6225) );
  OAI222_X1 U5986 ( .A1(n6232), .A2(n5670), .B1(n4858), .B2(n6266), .C1(n5672), 
        .C2(n6225), .ZN(U2855) );
  INV_X1 U5987 ( .A(EAX_REG_4__SCAN_IN), .ZN(n7003) );
  OAI222_X1 U5988 ( .A1(n6232), .A2(n5721), .B1(n5716), .B2(n4904), .C1(n7003), 
        .C2(n5715), .ZN(U2887) );
  XOR2_X1 U5989 ( .A(n4852), .B(n4859), .Z(n5622) );
  NOR2_X1 U5990 ( .A1(n6363), .A2(n5624), .ZN(n4862) );
  OAI22_X1 U5991 ( .A1(n5884), .A2(n4860), .B1(n6423), .B2(n6422), .ZN(n4861)
         );
  AOI211_X1 U5992 ( .C1(n5622), .C2(n6349), .A(n4862), .B(n4861), .ZN(n4867)
         );
  OR2_X1 U5993 ( .A1(n4864), .A2(n4863), .ZN(n6421) );
  NAND3_X1 U5994 ( .A1(n6421), .A2(n6358), .A3(n4865), .ZN(n4866) );
  NAND2_X1 U5995 ( .A1(n4867), .A2(n4866), .ZN(U2983) );
  XNOR2_X1 U5996 ( .A(n4851), .B(n4868), .ZN(n6215) );
  AOI22_X1 U5997 ( .A1(n5719), .A2(DATAI_5_), .B1(EAX_REG_5__SCAN_IN), .B2(
        n5718), .ZN(n4869) );
  OAI21_X1 U5998 ( .B1(n6215), .B2(n5721), .A(n4869), .ZN(U2886) );
  INV_X1 U5999 ( .A(n5622), .ZN(n4882) );
  INV_X1 U6000 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6292) );
  OAI222_X1 U6001 ( .A1(n5721), .A2(n4882), .B1(n5715), .B2(n6292), .C1(n4908), 
        .C2(n5716), .ZN(U2888) );
  NOR2_X1 U6002 ( .A1(n4870), .A2(n4788), .ZN(n4876) );
  NOR3_X1 U6003 ( .A1(n4876), .A2(n4875), .A3(FLUSH_REG_SCAN_IN), .ZN(n4873)
         );
  INV_X1 U6004 ( .A(n6747), .ZN(n4966) );
  NAND2_X1 U6005 ( .A1(n4874), .A2(n4966), .ZN(n4871) );
  NOR3_X1 U6006 ( .A1(n4876), .A2(n4875), .A3(n4874), .ZN(n4968) );
  AND2_X1 U6007 ( .A1(n5072), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6106) );
  INV_X1 U6008 ( .A(n3114), .ZN(n6521) );
  OAI22_X1 U6009 ( .A1(n4157), .A2(n6655), .B1(n6106), .B2(n6521), .ZN(n4877)
         );
  OAI21_X1 U6010 ( .B1(n4968), .B2(n4877), .A(n6448), .ZN(n4878) );
  OAI21_X1 U6011 ( .B1(n6448), .B2(n6651), .A(n4878), .ZN(U3465) );
  NAND2_X1 U6012 ( .A1(n4832), .A2(n4879), .ZN(n4880) );
  NAND2_X1 U6013 ( .A1(n4881), .A2(n4880), .ZN(n5623) );
  INV_X1 U6014 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4883) );
  OAI222_X1 U6015 ( .A1(n5672), .A2(n5623), .B1(n4883), .B2(n6266), .C1(n5670), 
        .C2(n4882), .ZN(U2856) );
  NOR2_X1 U6016 ( .A1(n4855), .A2(n4885), .ZN(n4886) );
  OR2_X1 U6017 ( .A1(n4884), .A2(n4886), .ZN(n6207) );
  OAI222_X1 U6018 ( .A1(n5672), .A2(n6207), .B1(n6209), .B2(n6266), .C1(n5670), 
        .C2(n6215), .ZN(U2854) );
  NAND2_X1 U6019 ( .A1(n5029), .A2(n6589), .ZN(n6519) );
  INV_X1 U6020 ( .A(n6519), .ZN(n4889) );
  NAND2_X1 U6021 ( .A1(n6518), .A2(n4889), .ZN(n5075) );
  NOR3_X1 U6022 ( .A1(n6452), .A2(n3601), .A3(n5212), .ZN(n4890) );
  OAI21_X1 U6023 ( .B1(n4890), .B2(n5888), .A(n6109), .ZN(n4892) );
  NAND2_X1 U6024 ( .A1(n4743), .A2(n3114), .ZN(n5214) );
  AND2_X1 U6025 ( .A1(n3104), .A2(n4786), .ZN(n5161) );
  INV_X1 U6026 ( .A(n5161), .ZN(n5258) );
  OR2_X1 U6027 ( .A1(n5214), .A2(n5258), .ZN(n4891) );
  NAND2_X1 U6028 ( .A1(n4892), .A2(n4894), .ZN(n4893) );
  NAND2_X1 U6029 ( .A1(n4929), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4903)
         );
  NAND2_X1 U6030 ( .A1(n6349), .A2(DATAI_29_), .ZN(n6699) );
  INV_X1 U6031 ( .A(n6699), .ZN(n5319) );
  INV_X1 U6032 ( .A(n4894), .ZN(n4895) );
  NAND2_X1 U6033 ( .A1(n4895), .A2(n6594), .ZN(n4897) );
  NAND2_X1 U6034 ( .A1(n5255), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4896) );
  OAI22_X1 U6035 ( .A1(n4932), .A2(n5325), .B1(n4931), .B2(n6628), .ZN(n4901)
         );
  AOI21_X1 U6036 ( .B1(n5319), .B2(n5286), .A(n4901), .ZN(n4902) );
  OAI211_X1 U6037 ( .C1(n5075), .C2(n6632), .A(n4903), .B(n4902), .ZN(U3145)
         );
  NAND2_X1 U6038 ( .A1(n4929), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4907)
         );
  NAND2_X1 U6039 ( .A1(n6349), .A2(DATAI_28_), .ZN(n6693) );
  INV_X1 U6040 ( .A(n6693), .ZN(n5356) );
  OR2_X1 U6041 ( .A1(n4930), .A2(n3445), .ZN(n6623) );
  OAI22_X1 U6042 ( .A1(n4932), .A2(n5361), .B1(n4931), .B2(n6623), .ZN(n4905)
         );
  AOI21_X1 U6043 ( .B1(n5356), .B2(n5286), .A(n4905), .ZN(n4906) );
  OAI211_X1 U6044 ( .C1(n5075), .C2(n6624), .A(n4907), .B(n4906), .ZN(U3144)
         );
  NAND2_X1 U6045 ( .A1(n6349), .A2(DATAI_19_), .ZN(n6619) );
  NAND2_X1 U6046 ( .A1(n4929), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4912)
         );
  NAND2_X1 U6047 ( .A1(n6349), .A2(DATAI_27_), .ZN(n6687) );
  INV_X1 U6048 ( .A(n6687), .ZN(n5340) );
  OAI22_X1 U6049 ( .A1(n4932), .A2(n5343), .B1(n4931), .B2(n6618), .ZN(n4910)
         );
  AOI21_X1 U6050 ( .B1(n5340), .B2(n5286), .A(n4910), .ZN(n4911) );
  OAI211_X1 U6051 ( .C1(n5075), .C2(n6619), .A(n4912), .B(n4911), .ZN(U3143)
         );
  NAND2_X1 U6052 ( .A1(n6349), .A2(DATAI_17_), .ZN(n6609) );
  NAND2_X1 U6053 ( .A1(n4929), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4916)
         );
  INV_X1 U6054 ( .A(n6675), .ZN(n5350) );
  OAI22_X1 U6055 ( .A1(n4932), .A2(n5353), .B1(n4931), .B2(n6608), .ZN(n4914)
         );
  AOI21_X1 U6056 ( .B1(n5350), .B2(n5286), .A(n4914), .ZN(n4915) );
  OAI211_X1 U6057 ( .C1(n5075), .C2(n6609), .A(n4916), .B(n4915), .ZN(U3141)
         );
  NAND2_X1 U6058 ( .A1(n4929), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4919)
         );
  NAND2_X1 U6059 ( .A1(n6349), .A2(DATAI_26_), .ZN(n6681) );
  OAI22_X1 U6060 ( .A1(n4932), .A2(n5338), .B1(n4931), .B2(n6613), .ZN(n4917)
         );
  AOI21_X1 U6061 ( .B1(n5335), .B2(n5286), .A(n4917), .ZN(n4918) );
  OAI211_X1 U6062 ( .C1(n5075), .C2(n6617), .A(n4919), .B(n4918), .ZN(U3142)
         );
  NAND2_X1 U6063 ( .A1(n4929), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4923)
         );
  OAI22_X1 U6064 ( .A1(n4932), .A2(n7081), .B1(n4931), .B2(n7072), .ZN(n4921)
         );
  AOI21_X1 U6065 ( .B1(n7077), .B2(n5286), .A(n4921), .ZN(n4922) );
  OAI211_X1 U6066 ( .C1(n5075), .C2(n7073), .A(n4923), .B(n4922), .ZN(U3146)
         );
  NAND2_X1 U6067 ( .A1(n6349), .A2(DATAI_16_), .ZN(n6591) );
  NAND2_X1 U6068 ( .A1(n4929), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4928)
         );
  NAND2_X1 U6069 ( .A1(n6349), .A2(DATAI_24_), .ZN(n6669) );
  INV_X1 U6070 ( .A(n6669), .ZN(n5345) );
  OAI22_X1 U6071 ( .A1(n4932), .A2(n5348), .B1(n4931), .B2(n6590), .ZN(n4926)
         );
  AOI21_X1 U6072 ( .B1(n5345), .B2(n5286), .A(n4926), .ZN(n4927) );
  OAI211_X1 U6073 ( .C1(n5075), .C2(n6591), .A(n4928), .B(n4927), .ZN(U3140)
         );
  NAND2_X1 U6074 ( .A1(n4929), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4935)
         );
  NAND2_X1 U6075 ( .A1(n6349), .A2(DATAI_31_), .ZN(n6716) );
  INV_X1 U6076 ( .A(n6716), .ZN(n5330) );
  INV_X1 U6077 ( .A(DATAI_7_), .ZN(n5069) );
  OAI22_X1 U6078 ( .A1(n4932), .A2(n5333), .B1(n4931), .B2(n6637), .ZN(n4933)
         );
  AOI21_X1 U6079 ( .B1(n5330), .B2(n5286), .A(n4933), .ZN(n4934) );
  OAI211_X1 U6080 ( .C1(n5075), .C2(n6638), .A(n4935), .B(n4934), .ZN(U3147)
         );
  NAND2_X1 U6081 ( .A1(n5029), .A2(n3601), .ZN(n6104) );
  INV_X1 U6082 ( .A(n4940), .ZN(n4936) );
  AOI21_X1 U6083 ( .B1(n4936), .B2(STATEBS16_REG_SCAN_IN), .A(n6655), .ZN(
        n4943) );
  INV_X1 U6084 ( .A(n4786), .ZN(n6099) );
  NAND2_X1 U6085 ( .A1(n6099), .A2(n3104), .ZN(n6657) );
  NOR2_X1 U6086 ( .A1(n6657), .A2(n4937), .ZN(n6496) );
  AND3_X1 U6087 ( .A1(n4975), .A2(n6781), .A3(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), 
        .ZN(n6491) );
  NAND2_X1 U6088 ( .A1(n6491), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n7071) );
  INV_X1 U6089 ( .A(n7071), .ZN(n4938) );
  AOI21_X1 U6090 ( .B1(n6496), .B2(n3114), .A(n4938), .ZN(n4942) );
  INV_X1 U6091 ( .A(n4942), .ZN(n4939) );
  NOR2_X1 U6092 ( .A1(n4940), .A2(n4157), .ZN(n5155) );
  OAI22_X1 U6093 ( .A1(n7074), .A2(n6638), .B1(n6637), .B2(n7071), .ZN(n4941)
         );
  AOI21_X1 U6094 ( .B1(n5330), .B2(n7076), .A(n4941), .ZN(n4946) );
  NAND2_X1 U6095 ( .A1(n4943), .A2(n4942), .ZN(n4944) );
  NAND2_X1 U6096 ( .A1(n7078), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4945) );
  OAI211_X1 U6097 ( .C1(n7082), .C2(n5333), .A(n4946), .B(n4945), .ZN(U3067)
         );
  OAI22_X1 U6098 ( .A1(n7074), .A2(n6617), .B1(n6613), .B2(n7071), .ZN(n4947)
         );
  AOI21_X1 U6099 ( .B1(n5335), .B2(n7076), .A(n4947), .ZN(n4949) );
  NAND2_X1 U6100 ( .A1(n7078), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4948) );
  OAI211_X1 U6101 ( .C1(n7082), .C2(n5338), .A(n4949), .B(n4948), .ZN(U3062)
         );
  OAI22_X1 U6102 ( .A1(n7074), .A2(n6619), .B1(n6618), .B2(n7071), .ZN(n4950)
         );
  AOI21_X1 U6103 ( .B1(n5340), .B2(n7076), .A(n4950), .ZN(n4952) );
  NAND2_X1 U6104 ( .A1(n7078), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4951) );
  OAI211_X1 U6105 ( .C1(n7082), .C2(n5343), .A(n4952), .B(n4951), .ZN(U3063)
         );
  OAI22_X1 U6106 ( .A1(n7074), .A2(n6591), .B1(n6590), .B2(n7071), .ZN(n4953)
         );
  AOI21_X1 U6107 ( .B1(n5345), .B2(n7076), .A(n4953), .ZN(n4955) );
  NAND2_X1 U6108 ( .A1(n7078), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4954) );
  OAI211_X1 U6109 ( .C1(n7082), .C2(n5348), .A(n4955), .B(n4954), .ZN(U3060)
         );
  OAI22_X1 U6110 ( .A1(n7074), .A2(n6609), .B1(n6608), .B2(n7071), .ZN(n4956)
         );
  AOI21_X1 U6111 ( .B1(n5350), .B2(n7076), .A(n4956), .ZN(n4958) );
  NAND2_X1 U6112 ( .A1(n7078), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4957) );
  OAI211_X1 U6113 ( .C1(n7082), .C2(n5353), .A(n4958), .B(n4957), .ZN(U3061)
         );
  OAI22_X1 U6114 ( .A1(n7074), .A2(n6624), .B1(n6623), .B2(n7071), .ZN(n4959)
         );
  AOI21_X1 U6115 ( .B1(n5356), .B2(n7076), .A(n4959), .ZN(n4961) );
  NAND2_X1 U6116 ( .A1(n7078), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4960) );
  OAI211_X1 U6117 ( .C1(n7082), .C2(n5361), .A(n4961), .B(n4960), .ZN(U3064)
         );
  OAI22_X1 U6118 ( .A1(n7074), .A2(n6632), .B1(n6628), .B2(n7071), .ZN(n4962)
         );
  AOI21_X1 U6119 ( .B1(n5319), .B2(n7076), .A(n4962), .ZN(n4964) );
  NAND2_X1 U6120 ( .A1(n7078), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4963) );
  OAI211_X1 U6121 ( .C1(n7082), .C2(n5325), .A(n4964), .B(n4963), .ZN(U3065)
         );
  INV_X1 U6122 ( .A(n4965), .ZN(n4974) );
  OAI21_X1 U6123 ( .B1(n4966), .B2(n6121), .A(n4967), .ZN(n4970) );
  OAI21_X1 U6124 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4811), .A(n4967), .ZN(
        n6718) );
  NOR2_X1 U6125 ( .A1(n6718), .A2(n4968), .ZN(n4969) );
  MUX2_X1 U6126 ( .A(n4970), .B(n4969), .S(STATE2_REG_0__SCAN_IN), .Z(n4972)
         );
  OAI211_X1 U6127 ( .C1(n4974), .C2(n4973), .A(n4972), .B(n4971), .ZN(U3148)
         );
  AND2_X1 U6128 ( .A1(n4976), .A2(n4975), .ZN(n6652) );
  INV_X1 U6129 ( .A(n5214), .ZN(n4978) );
  INV_X1 U6130 ( .A(n6657), .ZN(n4977) );
  AND2_X1 U6131 ( .A1(n6652), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4981)
         );
  AOI21_X1 U6132 ( .B1(n4978), .B2(n4977), .A(n4981), .ZN(n4986) );
  NOR2_X1 U6133 ( .A1(n4986), .A2(n6655), .ZN(n4979) );
  NOR2_X1 U6134 ( .A1(n4888), .A2(n3601), .ZN(n4980) );
  INV_X1 U6135 ( .A(n4981), .ZN(n5016) );
  NAND2_X1 U6136 ( .A1(n5252), .A2(n6711), .ZN(n4982) );
  OAI21_X1 U6137 ( .B1(n5016), .B2(n6637), .A(n4982), .ZN(n4983) );
  AOI21_X1 U6138 ( .B1(n5330), .B2(n6710), .A(n4983), .ZN(n4990) );
  INV_X1 U6139 ( .A(n4984), .ZN(n4985) );
  NOR2_X1 U6140 ( .A1(n4985), .A2(n6129), .ZN(n6105) );
  INV_X1 U6141 ( .A(n4986), .ZN(n4987) );
  OR3_X1 U6142 ( .A1(n6105), .A2(n6655), .A3(n4987), .ZN(n4988) );
  NAND2_X1 U6143 ( .A1(n5018), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4989)
         );
  OAI211_X1 U6144 ( .C1(n5021), .C2(n5333), .A(n4990), .B(n4989), .ZN(U3131)
         );
  INV_X1 U6145 ( .A(n7073), .ZN(n6702) );
  NAND2_X1 U6146 ( .A1(n5252), .A2(n6702), .ZN(n4991) );
  OAI21_X1 U6147 ( .B1(n5016), .B2(n7072), .A(n4991), .ZN(n4992) );
  AOI21_X1 U6148 ( .B1(n7077), .B2(n6710), .A(n4992), .ZN(n4994) );
  NAND2_X1 U6149 ( .A1(n5018), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4993)
         );
  OAI211_X1 U6150 ( .C1(n5021), .C2(n7081), .A(n4994), .B(n4993), .ZN(U3130)
         );
  INV_X1 U6151 ( .A(n6609), .ZN(n6672) );
  NAND2_X1 U6152 ( .A1(n5252), .A2(n6672), .ZN(n4995) );
  OAI21_X1 U6153 ( .B1(n5016), .B2(n6608), .A(n4995), .ZN(n4996) );
  AOI21_X1 U6154 ( .B1(n5350), .B2(n6710), .A(n4996), .ZN(n4998) );
  NAND2_X1 U6155 ( .A1(n5018), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4997)
         );
  OAI211_X1 U6156 ( .C1(n5021), .C2(n5353), .A(n4998), .B(n4997), .ZN(U3125)
         );
  INV_X1 U6157 ( .A(n6591), .ZN(n6666) );
  NAND2_X1 U6158 ( .A1(n5252), .A2(n6666), .ZN(n4999) );
  OAI21_X1 U6159 ( .B1(n5016), .B2(n6590), .A(n4999), .ZN(n5000) );
  AOI21_X1 U6160 ( .B1(n5345), .B2(n6710), .A(n5000), .ZN(n5002) );
  NAND2_X1 U6161 ( .A1(n5018), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n5001)
         );
  OAI211_X1 U6162 ( .C1(n5021), .C2(n5348), .A(n5002), .B(n5001), .ZN(U3124)
         );
  INV_X1 U6163 ( .A(n6632), .ZN(n6696) );
  NAND2_X1 U6164 ( .A1(n5252), .A2(n6696), .ZN(n5003) );
  OAI21_X1 U6165 ( .B1(n5016), .B2(n6628), .A(n5003), .ZN(n5004) );
  AOI21_X1 U6166 ( .B1(n5319), .B2(n6710), .A(n5004), .ZN(n5006) );
  NAND2_X1 U6167 ( .A1(n5018), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n5005)
         );
  OAI211_X1 U6168 ( .C1(n5021), .C2(n5325), .A(n5006), .B(n5005), .ZN(U3129)
         );
  NAND2_X1 U6169 ( .A1(n5252), .A2(n6684), .ZN(n5007) );
  OAI21_X1 U6170 ( .B1(n5016), .B2(n6618), .A(n5007), .ZN(n5008) );
  AOI21_X1 U6171 ( .B1(n5340), .B2(n6710), .A(n5008), .ZN(n5010) );
  NAND2_X1 U6172 ( .A1(n5018), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n5009)
         );
  OAI211_X1 U6173 ( .C1(n5021), .C2(n5343), .A(n5010), .B(n5009), .ZN(U3127)
         );
  INV_X1 U6174 ( .A(n6624), .ZN(n6690) );
  NAND2_X1 U6175 ( .A1(n5252), .A2(n6690), .ZN(n5011) );
  OAI21_X1 U6176 ( .B1(n5016), .B2(n6623), .A(n5011), .ZN(n5012) );
  AOI21_X1 U6177 ( .B1(n5356), .B2(n6710), .A(n5012), .ZN(n5014) );
  NAND2_X1 U6178 ( .A1(n5018), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n5013)
         );
  OAI211_X1 U6179 ( .C1(n5021), .C2(n5361), .A(n5014), .B(n5013), .ZN(U3128)
         );
  INV_X1 U6180 ( .A(n6617), .ZN(n6678) );
  NAND2_X1 U6181 ( .A1(n5252), .A2(n6678), .ZN(n5015) );
  OAI21_X1 U6182 ( .B1(n5016), .B2(n6613), .A(n5015), .ZN(n5017) );
  AOI21_X1 U6183 ( .B1(n5335), .B2(n6710), .A(n5017), .ZN(n5020) );
  NAND2_X1 U6184 ( .A1(n5018), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n5019)
         );
  OAI211_X1 U6185 ( .C1(n5021), .C2(n5338), .A(n5020), .B(n5019), .ZN(U3126)
         );
  OAI21_X1 U6186 ( .B1(n4884), .B2(n5023), .A(n5135), .ZN(n6396) );
  XOR2_X1 U6187 ( .A(n5024), .B(n5025), .Z(n6340) );
  INV_X1 U6188 ( .A(n6340), .ZN(n5065) );
  OAI222_X1 U6189 ( .A1(n6396), .A2(n5672), .B1(n5670), .B2(n5065), .C1(n5026), 
        .C2(n6266), .ZN(U2853) );
  OAI21_X1 U6190 ( .B1(n5032), .B2(n6655), .A(n6109), .ZN(n5035) );
  NOR2_X1 U6191 ( .A1(n4743), .A2(n6560), .ZN(n5077) );
  NOR2_X1 U6192 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5213) );
  NAND2_X1 U6193 ( .A1(n5213), .A2(n6781), .ZN(n5071) );
  OR2_X1 U6194 ( .A1(n5071), .A2(n6651), .ZN(n5058) );
  INV_X1 U6195 ( .A(n5058), .ZN(n5030) );
  AOI21_X1 U6196 ( .B1(n5077), .B2(n3114), .A(n5030), .ZN(n5034) );
  INV_X1 U6197 ( .A(n5034), .ZN(n5031) );
  INV_X1 U6198 ( .A(n5071), .ZN(n5037) );
  OAI22_X1 U6199 ( .A1(n5134), .A2(n6624), .B1(n6623), .B2(n5058), .ZN(n5033)
         );
  AOI21_X1 U6200 ( .B1(n5356), .B2(n5060), .A(n5033), .ZN(n5039) );
  NAND2_X1 U6201 ( .A1(n5035), .A2(n5034), .ZN(n5036) );
  NAND2_X1 U6202 ( .A1(n5061), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n5038) );
  OAI211_X1 U6203 ( .C1(n5064), .C2(n5361), .A(n5039), .B(n5038), .ZN(U3032)
         );
  OAI22_X1 U6204 ( .A1(n5134), .A2(n6619), .B1(n6618), .B2(n5058), .ZN(n5040)
         );
  AOI21_X1 U6205 ( .B1(n5340), .B2(n5060), .A(n5040), .ZN(n5042) );
  NAND2_X1 U6206 ( .A1(n5061), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n5041) );
  OAI211_X1 U6207 ( .C1(n5064), .C2(n5343), .A(n5042), .B(n5041), .ZN(U3031)
         );
  OAI22_X1 U6208 ( .A1(n5134), .A2(n7073), .B1(n7072), .B2(n5058), .ZN(n5043)
         );
  AOI21_X1 U6209 ( .B1(n7077), .B2(n5060), .A(n5043), .ZN(n5045) );
  NAND2_X1 U6210 ( .A1(n5061), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5044) );
  OAI211_X1 U6211 ( .C1(n5064), .C2(n7081), .A(n5045), .B(n5044), .ZN(U3034)
         );
  OAI22_X1 U6212 ( .A1(n5134), .A2(n6609), .B1(n6608), .B2(n5058), .ZN(n5046)
         );
  AOI21_X1 U6213 ( .B1(n5350), .B2(n5060), .A(n5046), .ZN(n5048) );
  NAND2_X1 U6214 ( .A1(n5061), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n5047) );
  OAI211_X1 U6215 ( .C1(n5064), .C2(n5353), .A(n5048), .B(n5047), .ZN(U3029)
         );
  OAI22_X1 U6216 ( .A1(n5134), .A2(n6638), .B1(n6637), .B2(n5058), .ZN(n5049)
         );
  AOI21_X1 U6217 ( .B1(n5330), .B2(n5060), .A(n5049), .ZN(n5051) );
  NAND2_X1 U6218 ( .A1(n5061), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5050) );
  OAI211_X1 U6219 ( .C1(n5064), .C2(n5333), .A(n5051), .B(n5050), .ZN(U3035)
         );
  OAI22_X1 U6220 ( .A1(n5134), .A2(n6617), .B1(n6613), .B2(n5058), .ZN(n5052)
         );
  AOI21_X1 U6221 ( .B1(n5335), .B2(n5060), .A(n5052), .ZN(n5054) );
  NAND2_X1 U6222 ( .A1(n5061), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n5053) );
  OAI211_X1 U6223 ( .C1(n5064), .C2(n5338), .A(n5054), .B(n5053), .ZN(U3030)
         );
  OAI22_X1 U6224 ( .A1(n5134), .A2(n6591), .B1(n6590), .B2(n5058), .ZN(n5055)
         );
  AOI21_X1 U6225 ( .B1(n5345), .B2(n5060), .A(n5055), .ZN(n5057) );
  NAND2_X1 U6226 ( .A1(n5061), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n5056) );
  OAI211_X1 U6227 ( .C1(n5064), .C2(n5348), .A(n5057), .B(n5056), .ZN(U3028)
         );
  OAI22_X1 U6228 ( .A1(n5134), .A2(n6632), .B1(n6628), .B2(n5058), .ZN(n5059)
         );
  AOI21_X1 U6229 ( .B1(n5319), .B2(n5060), .A(n5059), .ZN(n5063) );
  NAND2_X1 U6230 ( .A1(n5061), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n5062) );
  OAI211_X1 U6231 ( .C1(n5064), .C2(n5325), .A(n5063), .B(n5062), .ZN(U3033)
         );
  OAI222_X1 U6232 ( .A1(n5715), .A2(n5066), .B1(n4920), .B2(n5716), .C1(n5721), 
        .C2(n5065), .ZN(U2885) );
  XOR2_X1 U6233 ( .A(n5067), .B(n5150), .Z(n5210) );
  OAI222_X1 U6234 ( .A1(n5721), .A2(n6194), .B1(n5715), .B2(n4640), .C1(n5069), 
        .C2(n5716), .ZN(U2884) );
  AOI21_X1 U6235 ( .B1(n5310), .B2(n5075), .A(n6129), .ZN(n5070) );
  NOR3_X1 U6236 ( .A1(n5070), .A2(n5077), .A3(n6655), .ZN(n5074) );
  NOR2_X1 U6237 ( .A1(n5071), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5078)
         );
  NOR2_X1 U6238 ( .A1(n5078), .A2(n5072), .ZN(n5073) );
  INV_X1 U6239 ( .A(n6563), .ZN(n6649) );
  AOI21_X1 U6240 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6645), .A(n5100), .ZN(
        n6562) );
  OAI21_X1 U6241 ( .B1(n6649), .B2(n6603), .A(n6562), .ZN(n6493) );
  OR2_X1 U6242 ( .A1(n5076), .A2(n6603), .ZN(n5315) );
  NOR2_X1 U6243 ( .A1(n5315), .A2(n6645), .ZN(n6557) );
  AOI22_X1 U6244 ( .A1(n5077), .A2(n6594), .B1(n6557), .B2(n6649), .ZN(n5305)
         );
  INV_X1 U6245 ( .A(n5078), .ZN(n5304) );
  OAI22_X1 U6246 ( .A1(n5305), .A2(n5353), .B1(n6608), .B2(n5304), .ZN(n5080)
         );
  NOR2_X1 U6247 ( .A1(n5310), .A2(n6609), .ZN(n5079) );
  AOI211_X1 U6248 ( .C1(n5307), .C2(n5350), .A(n5080), .B(n5079), .ZN(n5081)
         );
  OAI21_X1 U6249 ( .B1(n5290), .B2(n5082), .A(n5081), .ZN(U3021) );
  OAI22_X1 U6250 ( .A1(n5305), .A2(n5333), .B1(n6637), .B2(n5304), .ZN(n5084)
         );
  NOR2_X1 U6251 ( .A1(n5310), .A2(n6638), .ZN(n5083) );
  AOI211_X1 U6252 ( .C1(n5307), .C2(n5330), .A(n5084), .B(n5083), .ZN(n5085)
         );
  OAI21_X1 U6253 ( .B1(n5290), .B2(n5086), .A(n5085), .ZN(U3027) );
  OAI22_X1 U6254 ( .A1(n5305), .A2(n5348), .B1(n6590), .B2(n5304), .ZN(n5088)
         );
  NOR2_X1 U6255 ( .A1(n5310), .A2(n6591), .ZN(n5087) );
  AOI211_X1 U6256 ( .C1(n5307), .C2(n5345), .A(n5088), .B(n5087), .ZN(n5089)
         );
  OAI21_X1 U6257 ( .B1(n5290), .B2(n5090), .A(n5089), .ZN(U3020) );
  OAI21_X1 U6258 ( .B1(n5093), .B2(n5092), .A(n5091), .ZN(n6404) );
  NAND2_X1 U6259 ( .A1(n6433), .A2(REIP_REG_5__SCAN_IN), .ZN(n6407) );
  OAI21_X1 U6260 ( .B1(n5884), .B2(n6960), .A(n6407), .ZN(n5095) );
  NOR2_X1 U6261 ( .A1(n6215), .A2(n5888), .ZN(n5094) );
  AOI211_X1 U6262 ( .C1(n6330), .C2(n6212), .A(n5095), .B(n5094), .ZN(n5096)
         );
  OAI21_X1 U6263 ( .B1(n6334), .B2(n6404), .A(n5096), .ZN(U2981) );
  OAI21_X1 U6264 ( .B1(n5097), .B2(n5131), .A(n6109), .ZN(n5098) );
  INV_X1 U6265 ( .A(n4743), .ZN(n6561) );
  INV_X1 U6266 ( .A(n3104), .ZN(n6101) );
  AND2_X1 U6267 ( .A1(n6101), .A2(n4786), .ZN(n5314) );
  NAND2_X1 U6268 ( .A1(n6561), .A2(n5314), .ZN(n6454) );
  AOI21_X1 U6269 ( .B1(n5098), .B2(n6454), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n5102) );
  NAND2_X1 U6270 ( .A1(n6456), .A2(n6781), .ZN(n6460) );
  NOR2_X1 U6271 ( .A1(n6460), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5105)
         );
  NOR2_X1 U6272 ( .A1(n6645), .A2(n6603), .ZN(n5099) );
  AND2_X1 U6273 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        STATE2_REG_2__SCAN_IN), .ZN(n5101) );
  NAND2_X1 U6274 ( .A1(n5127), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5108) );
  INV_X1 U6275 ( .A(n6454), .ZN(n5104) );
  NOR2_X1 U6276 ( .A1(n5315), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5103)
         );
  AOI22_X1 U6277 ( .A1(n5104), .A2(n6594), .B1(n6645), .B2(n5103), .ZN(n5129)
         );
  INV_X1 U6278 ( .A(n5105), .ZN(n5128) );
  OAI22_X1 U6279 ( .A1(n5129), .A2(n5325), .B1(n6628), .B2(n5128), .ZN(n5106)
         );
  AOI21_X1 U6280 ( .B1(n5131), .B2(n6696), .A(n5106), .ZN(n5107) );
  OAI211_X1 U6281 ( .C1(n5134), .C2(n6699), .A(n5108), .B(n5107), .ZN(U3041)
         );
  NAND2_X1 U6282 ( .A1(n5127), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5111) );
  OAI22_X1 U6283 ( .A1(n5129), .A2(n5348), .B1(n6590), .B2(n5128), .ZN(n5109)
         );
  AOI21_X1 U6284 ( .B1(n5131), .B2(n6666), .A(n5109), .ZN(n5110) );
  OAI211_X1 U6285 ( .C1(n5134), .C2(n6669), .A(n5111), .B(n5110), .ZN(U3036)
         );
  NAND2_X1 U6286 ( .A1(n5127), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5114) );
  OAI22_X1 U6287 ( .A1(n5129), .A2(n7081), .B1(n7072), .B2(n5128), .ZN(n5112)
         );
  AOI21_X1 U6288 ( .B1(n5131), .B2(n6702), .A(n5112), .ZN(n5113) );
  OAI211_X1 U6289 ( .C1(n5134), .C2(n6705), .A(n5114), .B(n5113), .ZN(U3042)
         );
  NAND2_X1 U6290 ( .A1(n5127), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5117) );
  OAI22_X1 U6291 ( .A1(n5129), .A2(n5333), .B1(n6637), .B2(n5128), .ZN(n5115)
         );
  AOI21_X1 U6292 ( .B1(n5131), .B2(n6711), .A(n5115), .ZN(n5116) );
  OAI211_X1 U6293 ( .C1(n5134), .C2(n6716), .A(n5117), .B(n5116), .ZN(U3043)
         );
  NAND2_X1 U6294 ( .A1(n5127), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5120) );
  OAI22_X1 U6295 ( .A1(n5129), .A2(n5361), .B1(n6623), .B2(n5128), .ZN(n5118)
         );
  AOI21_X1 U6296 ( .B1(n5131), .B2(n6690), .A(n5118), .ZN(n5119) );
  OAI211_X1 U6297 ( .C1(n5134), .C2(n6693), .A(n5120), .B(n5119), .ZN(U3040)
         );
  NAND2_X1 U6298 ( .A1(n5127), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5123) );
  OAI22_X1 U6299 ( .A1(n5129), .A2(n5343), .B1(n6618), .B2(n5128), .ZN(n5121)
         );
  AOI21_X1 U6300 ( .B1(n5131), .B2(n6684), .A(n5121), .ZN(n5122) );
  OAI211_X1 U6301 ( .C1(n5134), .C2(n6687), .A(n5123), .B(n5122), .ZN(U3039)
         );
  NAND2_X1 U6302 ( .A1(n5127), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5126) );
  OAI22_X1 U6303 ( .A1(n5129), .A2(n5338), .B1(n6613), .B2(n5128), .ZN(n5124)
         );
  AOI21_X1 U6304 ( .B1(n5131), .B2(n6678), .A(n5124), .ZN(n5125) );
  OAI211_X1 U6305 ( .C1(n5134), .C2(n6681), .A(n5126), .B(n5125), .ZN(U3038)
         );
  NAND2_X1 U6306 ( .A1(n5127), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5133) );
  OAI22_X1 U6307 ( .A1(n5129), .A2(n5353), .B1(n6608), .B2(n5128), .ZN(n5130)
         );
  AOI21_X1 U6308 ( .B1(n5131), .B2(n6672), .A(n5130), .ZN(n5132) );
  OAI211_X1 U6309 ( .C1(n5134), .C2(n6675), .A(n5133), .B(n5132), .ZN(U3037)
         );
  INV_X1 U6310 ( .A(n5135), .ZN(n5138) );
  OAI21_X1 U6311 ( .B1(n5138), .B2(n4323), .A(n5137), .ZN(n6188) );
  INV_X1 U6312 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5139) );
  OAI222_X1 U6313 ( .A1(n6188), .A2(n5672), .B1(n5670), .B2(n6194), .C1(n5139), 
        .C2(n6266), .ZN(U2852) );
  NAND2_X1 U6314 ( .A1(n5141), .A2(n5142), .ZN(n5143) );
  NAND2_X1 U6315 ( .A1(n5140), .A2(n5143), .ZN(n6328) );
  INV_X1 U6316 ( .A(n5145), .ZN(n5146) );
  AOI21_X1 U6317 ( .B1(n5147), .B2(n5144), .A(n5146), .ZN(n6084) );
  AOI22_X1 U6318 ( .A1(n6084), .A2(n6261), .B1(EBX_REG_11__SCAN_IN), .B2(n5659), .ZN(n5148) );
  OAI21_X1 U6319 ( .B1(n6328), .B2(n5670), .A(n5148), .ZN(U2848) );
  AOI22_X1 U6320 ( .A1(n5719), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n5718), .ZN(n5149) );
  OAI21_X1 U6321 ( .B1(n6328), .B2(n5721), .A(n5149), .ZN(U2880) );
  AND2_X1 U6322 ( .A1(n5067), .A2(n5150), .ZN(n5197) );
  NAND2_X1 U6323 ( .A1(n5197), .A2(n5196), .ZN(n5191) );
  INV_X1 U6324 ( .A(n5194), .ZN(n5151) );
  NOR2_X1 U6325 ( .A1(n5191), .A2(n5151), .ZN(n5192) );
  OAI21_X1 U6326 ( .B1(n5192), .B2(n5152), .A(n5141), .ZN(n5879) );
  AOI22_X1 U6327 ( .A1(n5719), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n5718), .ZN(n5153) );
  OAI21_X1 U6328 ( .B1(n5879), .B2(n5721), .A(n5153), .ZN(U2881) );
  INV_X1 U6329 ( .A(n5311), .ZN(n5154) );
  NOR3_X1 U6330 ( .A1(n5155), .A2(n5188), .A3(n6655), .ZN(n5156) );
  NAND2_X1 U6331 ( .A1(n5161), .A2(n6658), .ZN(n6522) );
  OAI21_X1 U6332 ( .B1(n5156), .B2(n6659), .A(n6522), .ZN(n5159) );
  NAND2_X1 U6333 ( .A1(n6526), .A2(n6651), .ZN(n5185) );
  NAND2_X1 U6334 ( .A1(n5185), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5157) );
  NAND4_X1 U6335 ( .A1(n5159), .A2(n5158), .A3(n5315), .A4(n5157), .ZN(n5184)
         );
  NAND2_X1 U6336 ( .A1(n5184), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5165) );
  NOR2_X1 U6337 ( .A1(n4743), .A2(n6655), .ZN(n5162) );
  INV_X1 U6338 ( .A(n6647), .ZN(n6490) );
  NOR2_X1 U6339 ( .A1(n6490), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5160)
         );
  AOI22_X1 U6340 ( .A1(n5162), .A2(n5161), .B1(n6645), .B2(n5160), .ZN(n5186)
         );
  OAI22_X1 U6341 ( .A1(n5186), .A2(n5333), .B1(n6637), .B2(n5185), .ZN(n5163)
         );
  AOI21_X1 U6342 ( .B1(n5188), .B2(n6711), .A(n5163), .ZN(n5164) );
  OAI211_X1 U6343 ( .C1(n7074), .C2(n6716), .A(n5165), .B(n5164), .ZN(U3075)
         );
  NAND2_X1 U6344 ( .A1(n5184), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5168) );
  OAI22_X1 U6345 ( .A1(n5186), .A2(n5343), .B1(n6618), .B2(n5185), .ZN(n5166)
         );
  AOI21_X1 U6346 ( .B1(n5188), .B2(n6684), .A(n5166), .ZN(n5167) );
  OAI211_X1 U6347 ( .C1(n7074), .C2(n6687), .A(n5168), .B(n5167), .ZN(U3071)
         );
  NAND2_X1 U6348 ( .A1(n5184), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5171) );
  OAI22_X1 U6349 ( .A1(n5186), .A2(n5353), .B1(n6608), .B2(n5185), .ZN(n5169)
         );
  AOI21_X1 U6350 ( .B1(n5188), .B2(n6672), .A(n5169), .ZN(n5170) );
  OAI211_X1 U6351 ( .C1(n7074), .C2(n6675), .A(n5171), .B(n5170), .ZN(U3069)
         );
  NAND2_X1 U6352 ( .A1(n5184), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5174) );
  OAI22_X1 U6353 ( .A1(n5186), .A2(n5338), .B1(n6613), .B2(n5185), .ZN(n5172)
         );
  AOI21_X1 U6354 ( .B1(n5188), .B2(n6678), .A(n5172), .ZN(n5173) );
  OAI211_X1 U6355 ( .C1(n7074), .C2(n6681), .A(n5174), .B(n5173), .ZN(U3070)
         );
  NAND2_X1 U6356 ( .A1(n5184), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5177) );
  OAI22_X1 U6357 ( .A1(n5186), .A2(n5361), .B1(n6623), .B2(n5185), .ZN(n5175)
         );
  AOI21_X1 U6358 ( .B1(n5188), .B2(n6690), .A(n5175), .ZN(n5176) );
  OAI211_X1 U6359 ( .C1(n7074), .C2(n6693), .A(n5177), .B(n5176), .ZN(U3072)
         );
  NAND2_X1 U6360 ( .A1(n5184), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5180) );
  OAI22_X1 U6361 ( .A1(n5186), .A2(n7081), .B1(n7072), .B2(n5185), .ZN(n5178)
         );
  AOI21_X1 U6362 ( .B1(n5188), .B2(n6702), .A(n5178), .ZN(n5179) );
  OAI211_X1 U6363 ( .C1(n7074), .C2(n6705), .A(n5180), .B(n5179), .ZN(U3074)
         );
  NAND2_X1 U6364 ( .A1(n5184), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5183) );
  OAI22_X1 U6365 ( .A1(n5186), .A2(n5325), .B1(n6628), .B2(n5185), .ZN(n5181)
         );
  AOI21_X1 U6366 ( .B1(n5188), .B2(n6696), .A(n5181), .ZN(n5182) );
  OAI211_X1 U6367 ( .C1(n7074), .C2(n6699), .A(n5183), .B(n5182), .ZN(U3073)
         );
  NAND2_X1 U6368 ( .A1(n5184), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n5190) );
  OAI22_X1 U6369 ( .A1(n5186), .A2(n5348), .B1(n6590), .B2(n5185), .ZN(n5187)
         );
  AOI21_X1 U6370 ( .B1(n5188), .B2(n6666), .A(n5187), .ZN(n5189) );
  OAI211_X1 U6371 ( .C1(n7074), .C2(n6669), .A(n5190), .B(n5189), .ZN(U3068)
         );
  INV_X1 U6372 ( .A(n5191), .ZN(n5198) );
  INV_X1 U6373 ( .A(n5192), .ZN(n5193) );
  OAI21_X1 U6374 ( .B1(n5198), .B2(n5194), .A(n5193), .ZN(n6161) );
  AOI22_X1 U6375 ( .A1(n5719), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n5718), .ZN(n5195) );
  OAI21_X1 U6376 ( .B1(n6161), .B2(n5721), .A(n5195), .ZN(U2882) );
  INV_X1 U6377 ( .A(n5196), .ZN(n5200) );
  INV_X1 U6378 ( .A(n5197), .ZN(n5199) );
  AOI21_X1 U6379 ( .B1(n5200), .B2(n5199), .A(n5198), .ZN(n6177) );
  INV_X1 U6380 ( .A(n6177), .ZN(n5204) );
  AOI22_X1 U6381 ( .A1(n5719), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n5718), .ZN(n5201) );
  OAI21_X1 U6382 ( .B1(n5204), .B2(n5721), .A(n5201), .ZN(U2883) );
  NAND2_X1 U6383 ( .A1(n5137), .A2(n5202), .ZN(n5203) );
  NAND2_X1 U6384 ( .A1(n6164), .A2(n5203), .ZN(n6172) );
  OAI222_X1 U6385 ( .A1(n5204), .A2(n5670), .B1(n7048), .B2(n6266), .C1(n6172), 
        .C2(n5672), .ZN(U2851) );
  OAI21_X1 U6386 ( .B1(n5207), .B2(n5206), .A(n3103), .ZN(n6384) );
  NAND2_X1 U6387 ( .A1(n6433), .A2(REIP_REG_7__SCAN_IN), .ZN(n6381) );
  NAND2_X1 U6388 ( .A1(n6354), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5208)
         );
  OAI211_X1 U6389 ( .C1(n6363), .C2(n6192), .A(n6381), .B(n5208), .ZN(n5209)
         );
  AOI21_X1 U6390 ( .B1(n5210), .B2(n6349), .A(n5209), .ZN(n5211) );
  OAI21_X1 U6391 ( .B1(n6384), .B2(n6334), .A(n5211), .ZN(U2979) );
  INV_X1 U6392 ( .A(n6567), .ZN(n5216) );
  NAND2_X1 U6393 ( .A1(n5213), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6559) );
  OR2_X1 U6394 ( .A1(n6559), .A2(n6651), .ZN(n5243) );
  OAI21_X1 U6395 ( .B1(n5214), .B2(n6560), .A(n5243), .ZN(n5222) );
  INV_X1 U6396 ( .A(n6559), .ZN(n5215) );
  OAI22_X1 U6397 ( .A1(n5244), .A2(n6591), .B1(n6590), .B2(n5243), .ZN(n5220)
         );
  AOI21_X1 U6398 ( .B1(n5345), .B2(n6584), .A(n5220), .ZN(n5224) );
  NAND2_X1 U6399 ( .A1(n6559), .A2(n6655), .ZN(n5221) );
  NAND2_X1 U6400 ( .A1(n5246), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n5223) );
  OAI211_X1 U6401 ( .C1(n5249), .C2(n5348), .A(n5224), .B(n5223), .ZN(U3092)
         );
  OAI22_X1 U6402 ( .A1(n5244), .A2(n7073), .B1(n7072), .B2(n5243), .ZN(n5225)
         );
  AOI21_X1 U6403 ( .B1(n7077), .B2(n6584), .A(n5225), .ZN(n5227) );
  NAND2_X1 U6404 ( .A1(n5246), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n5226) );
  OAI211_X1 U6405 ( .C1(n5249), .C2(n7081), .A(n5227), .B(n5226), .ZN(U3098)
         );
  OAI22_X1 U6406 ( .A1(n5244), .A2(n6632), .B1(n6628), .B2(n5243), .ZN(n5228)
         );
  AOI21_X1 U6407 ( .B1(n5319), .B2(n6584), .A(n5228), .ZN(n5230) );
  NAND2_X1 U6408 ( .A1(n5246), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n5229) );
  OAI211_X1 U6409 ( .C1(n5249), .C2(n5325), .A(n5230), .B(n5229), .ZN(U3097)
         );
  OAI22_X1 U6410 ( .A1(n5244), .A2(n6638), .B1(n6637), .B2(n5243), .ZN(n5231)
         );
  AOI21_X1 U6411 ( .B1(n5330), .B2(n6584), .A(n5231), .ZN(n5233) );
  NAND2_X1 U6412 ( .A1(n5246), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n5232) );
  OAI211_X1 U6413 ( .C1(n5249), .C2(n5333), .A(n5233), .B(n5232), .ZN(U3099)
         );
  OAI22_X1 U6414 ( .A1(n5244), .A2(n6619), .B1(n6618), .B2(n5243), .ZN(n5234)
         );
  AOI21_X1 U6415 ( .B1(n5340), .B2(n6584), .A(n5234), .ZN(n5236) );
  NAND2_X1 U6416 ( .A1(n5246), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n5235) );
  OAI211_X1 U6417 ( .C1(n5249), .C2(n5343), .A(n5236), .B(n5235), .ZN(U3095)
         );
  OAI22_X1 U6418 ( .A1(n5244), .A2(n6617), .B1(n6613), .B2(n5243), .ZN(n5237)
         );
  AOI21_X1 U6419 ( .B1(n5335), .B2(n6584), .A(n5237), .ZN(n5239) );
  NAND2_X1 U6420 ( .A1(n5246), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n5238) );
  OAI211_X1 U6421 ( .C1(n5249), .C2(n5338), .A(n5239), .B(n5238), .ZN(U3094)
         );
  OAI22_X1 U6422 ( .A1(n5244), .A2(n6609), .B1(n6608), .B2(n5243), .ZN(n5240)
         );
  AOI21_X1 U6423 ( .B1(n5350), .B2(n6584), .A(n5240), .ZN(n5242) );
  NAND2_X1 U6424 ( .A1(n5246), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n5241) );
  OAI211_X1 U6425 ( .C1(n5249), .C2(n5353), .A(n5242), .B(n5241), .ZN(U3093)
         );
  OAI22_X1 U6426 ( .A1(n5244), .A2(n6624), .B1(n6623), .B2(n5243), .ZN(n5245)
         );
  AOI21_X1 U6427 ( .B1(n5356), .B2(n6584), .A(n5245), .ZN(n5248) );
  NAND2_X1 U6428 ( .A1(n5246), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n5247) );
  OAI211_X1 U6429 ( .C1(n5249), .C2(n5361), .A(n5248), .B(n5247), .ZN(U3096)
         );
  XNOR2_X1 U6430 ( .A(n5140), .B(n3253), .ZN(n5872) );
  INV_X1 U6431 ( .A(n5872), .ZN(n5600) );
  AOI22_X1 U6432 ( .A1(n5719), .A2(DATAI_12_), .B1(EAX_REG_12__SCAN_IN), .B2(
        n5718), .ZN(n5251) );
  OAI21_X1 U6433 ( .B1(n5600), .B2(n5721), .A(n5251), .ZN(U2879) );
  NOR3_X1 U6434 ( .A1(n5252), .A2(n5286), .A3(n6655), .ZN(n5253) );
  OAI22_X1 U6435 ( .A1(n5253), .A2(n6659), .B1(n6658), .B2(n5258), .ZN(n5257)
         );
  AOI21_X1 U6436 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6781), .A(n5254), .ZN(
        n5321) );
  NAND2_X1 U6437 ( .A1(n5255), .A2(n6651), .ZN(n5283) );
  INV_X1 U6438 ( .A(n5315), .ZN(n6662) );
  AOI21_X1 U6439 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5283), .A(n6662), .ZN(
        n5256) );
  NAND3_X1 U6440 ( .A1(n5257), .A2(n5321), .A3(n5256), .ZN(n5282) );
  NAND2_X1 U6441 ( .A1(n5282), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5263)
         );
  NAND2_X1 U6442 ( .A1(n4743), .A2(n6594), .ZN(n6650) );
  OR2_X1 U6443 ( .A1(n6650), .A2(n5258), .ZN(n5260) );
  NAND3_X1 U6444 ( .A1(n6647), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6645), .ZN(n5259) );
  OAI22_X1 U6445 ( .A1(n5284), .A2(n5348), .B1(n6590), .B2(n5283), .ZN(n5261)
         );
  AOI21_X1 U6446 ( .B1(n5286), .B2(n6666), .A(n5261), .ZN(n5262) );
  OAI211_X1 U6447 ( .C1(n5289), .C2(n6669), .A(n5263), .B(n5262), .ZN(U3132)
         );
  NAND2_X1 U6448 ( .A1(n5282), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5266)
         );
  OAI22_X1 U6449 ( .A1(n5284), .A2(n5353), .B1(n6608), .B2(n5283), .ZN(n5264)
         );
  AOI21_X1 U6450 ( .B1(n5286), .B2(n6672), .A(n5264), .ZN(n5265) );
  OAI211_X1 U6451 ( .C1(n5289), .C2(n6675), .A(n5266), .B(n5265), .ZN(U3133)
         );
  NAND2_X1 U6452 ( .A1(n5282), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5269)
         );
  OAI22_X1 U6453 ( .A1(n5284), .A2(n5333), .B1(n6637), .B2(n5283), .ZN(n5267)
         );
  AOI21_X1 U6454 ( .B1(n5286), .B2(n6711), .A(n5267), .ZN(n5268) );
  OAI211_X1 U6455 ( .C1(n5289), .C2(n6716), .A(n5269), .B(n5268), .ZN(U3139)
         );
  NAND2_X1 U6456 ( .A1(n5282), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5272)
         );
  OAI22_X1 U6457 ( .A1(n5284), .A2(n7081), .B1(n7072), .B2(n5283), .ZN(n5270)
         );
  AOI21_X1 U6458 ( .B1(n5286), .B2(n6702), .A(n5270), .ZN(n5271) );
  OAI211_X1 U6459 ( .C1(n5289), .C2(n6705), .A(n5272), .B(n5271), .ZN(U3138)
         );
  NAND2_X1 U6460 ( .A1(n5282), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5275)
         );
  OAI22_X1 U6461 ( .A1(n5284), .A2(n5325), .B1(n6628), .B2(n5283), .ZN(n5273)
         );
  AOI21_X1 U6462 ( .B1(n5286), .B2(n6696), .A(n5273), .ZN(n5274) );
  OAI211_X1 U6463 ( .C1(n5289), .C2(n6699), .A(n5275), .B(n5274), .ZN(U3137)
         );
  NAND2_X1 U6464 ( .A1(n5282), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5278)
         );
  OAI22_X1 U6465 ( .A1(n5284), .A2(n5361), .B1(n6623), .B2(n5283), .ZN(n5276)
         );
  AOI21_X1 U6466 ( .B1(n5286), .B2(n6690), .A(n5276), .ZN(n5277) );
  OAI211_X1 U6467 ( .C1(n5289), .C2(n6693), .A(n5278), .B(n5277), .ZN(U3136)
         );
  NAND2_X1 U6468 ( .A1(n5282), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5281)
         );
  OAI22_X1 U6469 ( .A1(n5284), .A2(n5343), .B1(n6618), .B2(n5283), .ZN(n5279)
         );
  AOI21_X1 U6470 ( .B1(n5286), .B2(n6684), .A(n5279), .ZN(n5280) );
  OAI211_X1 U6471 ( .C1(n5289), .C2(n6687), .A(n5281), .B(n5280), .ZN(U3135)
         );
  NAND2_X1 U6472 ( .A1(n5282), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5288)
         );
  OAI22_X1 U6473 ( .A1(n5284), .A2(n5338), .B1(n6613), .B2(n5283), .ZN(n5285)
         );
  AOI21_X1 U6474 ( .B1(n5286), .B2(n6678), .A(n5285), .ZN(n5287) );
  OAI211_X1 U6475 ( .C1(n5289), .C2(n6681), .A(n5288), .B(n5287), .ZN(U3134)
         );
  INV_X1 U6476 ( .A(n5290), .ZN(n5303) );
  NAND2_X1 U6477 ( .A1(n5303), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5293) );
  OAI22_X1 U6478 ( .A1(n5305), .A2(n5325), .B1(n6628), .B2(n5304), .ZN(n5291)
         );
  AOI21_X1 U6479 ( .B1(n5307), .B2(n5319), .A(n5291), .ZN(n5292) );
  OAI211_X1 U6480 ( .C1(n5310), .C2(n6632), .A(n5293), .B(n5292), .ZN(U3025)
         );
  NAND2_X1 U6481 ( .A1(n5303), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5296) );
  OAI22_X1 U6482 ( .A1(n5305), .A2(n7081), .B1(n7072), .B2(n5304), .ZN(n5294)
         );
  AOI21_X1 U6483 ( .B1(n5307), .B2(n7077), .A(n5294), .ZN(n5295) );
  OAI211_X1 U6484 ( .C1(n5310), .C2(n7073), .A(n5296), .B(n5295), .ZN(U3026)
         );
  NAND2_X1 U6485 ( .A1(n5303), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5299) );
  OAI22_X1 U6486 ( .A1(n5305), .A2(n5361), .B1(n6623), .B2(n5304), .ZN(n5297)
         );
  AOI21_X1 U6487 ( .B1(n5307), .B2(n5356), .A(n5297), .ZN(n5298) );
  OAI211_X1 U6488 ( .C1(n5310), .C2(n6624), .A(n5299), .B(n5298), .ZN(U3024)
         );
  NAND2_X1 U6489 ( .A1(n5303), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5302) );
  OAI22_X1 U6490 ( .A1(n5305), .A2(n5343), .B1(n6618), .B2(n5304), .ZN(n5300)
         );
  AOI21_X1 U6491 ( .B1(n5307), .B2(n5340), .A(n5300), .ZN(n5301) );
  OAI211_X1 U6492 ( .C1(n5310), .C2(n6619), .A(n5302), .B(n5301), .ZN(U3023)
         );
  NAND2_X1 U6493 ( .A1(n5303), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5309) );
  OAI22_X1 U6494 ( .A1(n5305), .A2(n5338), .B1(n6613), .B2(n5304), .ZN(n5306)
         );
  AOI21_X1 U6495 ( .B1(n5307), .B2(n5335), .A(n5306), .ZN(n5308) );
  OAI211_X1 U6496 ( .C1(n5310), .C2(n6617), .A(n5309), .B(n5308), .ZN(U3022)
         );
  INV_X1 U6497 ( .A(n6644), .ZN(n5312) );
  OAI21_X1 U6498 ( .B1(n5357), .B2(n5312), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5313) );
  NAND2_X1 U6499 ( .A1(n5313), .A2(n6594), .ZN(n5322) );
  INV_X1 U6500 ( .A(n5322), .ZN(n5317) );
  NOR2_X1 U6501 ( .A1(n5315), .A2(n6781), .ZN(n5316) );
  AND2_X1 U6502 ( .A1(n6456), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6601)
         );
  NAND2_X1 U6503 ( .A1(n6601), .A2(n6651), .ZN(n5354) );
  OAI22_X1 U6504 ( .A1(n6644), .A2(n6632), .B1(n5354), .B2(n6628), .ZN(n5318)
         );
  AOI21_X1 U6505 ( .B1(n5357), .B2(n5319), .A(n5318), .ZN(n5324) );
  AOI21_X1 U6506 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5354), .A(n6647), .ZN(
        n5320) );
  NAND2_X1 U6507 ( .A1(n5358), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5323)
         );
  OAI211_X1 U6508 ( .C1(n5362), .C2(n5325), .A(n5324), .B(n5323), .ZN(U3105)
         );
  OAI22_X1 U6509 ( .A1(n6644), .A2(n7073), .B1(n5354), .B2(n7072), .ZN(n5326)
         );
  AOI21_X1 U6510 ( .B1(n5357), .B2(n7077), .A(n5326), .ZN(n5328) );
  NAND2_X1 U6511 ( .A1(n5358), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5327)
         );
  OAI211_X1 U6512 ( .C1(n5362), .C2(n7081), .A(n5328), .B(n5327), .ZN(U3106)
         );
  OAI22_X1 U6513 ( .A1(n6644), .A2(n6638), .B1(n5354), .B2(n6637), .ZN(n5329)
         );
  AOI21_X1 U6514 ( .B1(n5357), .B2(n5330), .A(n5329), .ZN(n5332) );
  NAND2_X1 U6515 ( .A1(n5358), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5331)
         );
  OAI211_X1 U6516 ( .C1(n5362), .C2(n5333), .A(n5332), .B(n5331), .ZN(U3107)
         );
  OAI22_X1 U6517 ( .A1(n6644), .A2(n6617), .B1(n5354), .B2(n6613), .ZN(n5334)
         );
  AOI21_X1 U6518 ( .B1(n5357), .B2(n5335), .A(n5334), .ZN(n5337) );
  NAND2_X1 U6519 ( .A1(n5358), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5336)
         );
  OAI211_X1 U6520 ( .C1(n5362), .C2(n5338), .A(n5337), .B(n5336), .ZN(U3102)
         );
  OAI22_X1 U6521 ( .A1(n6644), .A2(n6619), .B1(n5354), .B2(n6618), .ZN(n5339)
         );
  AOI21_X1 U6522 ( .B1(n5357), .B2(n5340), .A(n5339), .ZN(n5342) );
  NAND2_X1 U6523 ( .A1(n5358), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5341)
         );
  OAI211_X1 U6524 ( .C1(n5362), .C2(n5343), .A(n5342), .B(n5341), .ZN(U3103)
         );
  OAI22_X1 U6525 ( .A1(n6644), .A2(n6591), .B1(n5354), .B2(n6590), .ZN(n5344)
         );
  AOI21_X1 U6526 ( .B1(n5357), .B2(n5345), .A(n5344), .ZN(n5347) );
  NAND2_X1 U6527 ( .A1(n5358), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5346)
         );
  OAI211_X1 U6528 ( .C1(n5362), .C2(n5348), .A(n5347), .B(n5346), .ZN(U3100)
         );
  OAI22_X1 U6529 ( .A1(n6644), .A2(n6609), .B1(n5354), .B2(n6608), .ZN(n5349)
         );
  AOI21_X1 U6530 ( .B1(n5357), .B2(n5350), .A(n5349), .ZN(n5352) );
  NAND2_X1 U6531 ( .A1(n5358), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5351)
         );
  OAI211_X1 U6532 ( .C1(n5362), .C2(n5353), .A(n5352), .B(n5351), .ZN(U3101)
         );
  OAI22_X1 U6533 ( .A1(n6644), .A2(n6624), .B1(n5354), .B2(n6623), .ZN(n5355)
         );
  AOI21_X1 U6534 ( .B1(n5357), .B2(n5356), .A(n5355), .ZN(n5360) );
  NAND2_X1 U6535 ( .A1(n5358), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5359)
         );
  OAI211_X1 U6536 ( .C1(n5362), .C2(n5361), .A(n5360), .B(n5359), .ZN(U3104)
         );
  AOI21_X1 U6537 ( .B1(n5364), .B2(n5145), .A(n5363), .ZN(n6070) );
  INV_X1 U6538 ( .A(n6070), .ZN(n5366) );
  OAI222_X1 U6539 ( .A1(n5366), .A2(n5672), .B1(n5670), .B2(n5600), .C1(n5365), 
        .C2(n6266), .ZN(U2847) );
  AOI21_X1 U6540 ( .B1(n5367), .B2(n6119), .A(n6125), .ZN(n5373) );
  INV_X1 U6541 ( .A(n5368), .ZN(n5371) );
  OAI22_X1 U6542 ( .A1(n6121), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n5369), .ZN(n5370) );
  AOI21_X1 U6543 ( .B1(n6119), .B2(n5371), .A(n5370), .ZN(n5372) );
  OAI22_X1 U6544 ( .A1(n5373), .A2(n3269), .B1(n6125), .B2(n5372), .ZN(U3461)
         );
  AND2_X1 U6545 ( .A1(n5715), .A2(n5374), .ZN(n5375) );
  NAND2_X1 U6546 ( .A1(n5376), .A2(n5375), .ZN(n5378) );
  AOI22_X1 U6547 ( .A1(n5711), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n5718), .ZN(n5377) );
  NAND2_X1 U6548 ( .A1(n5378), .A2(n5377), .ZN(U2860) );
  NAND2_X1 U6549 ( .A1(n3402), .A2(n4316), .ZN(n5380) );
  OR2_X1 U6550 ( .A1(n5513), .A2(READREQUEST_REG_SCAN_IN), .ZN(n5379) );
  MUX2_X1 U6551 ( .A(n5380), .B(n5379), .S(n6741), .Z(U3474) );
  INV_X1 U6552 ( .A(n5726), .ZN(n5676) );
  INV_X1 U6553 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5643) );
  NAND3_X1 U6554 ( .A1(n4287), .A2(n5643), .A3(n5382), .ZN(n5383) );
  AND2_X1 U6555 ( .A1(n5384), .A2(n5383), .ZN(n5385) );
  NOR2_X1 U6556 ( .A1(n5399), .A2(n5386), .ZN(n5388) );
  OAI21_X1 U6557 ( .B1(n5388), .B2(REIP_REG_30__SCAN_IN), .A(n5387), .ZN(n5392) );
  INV_X1 U6558 ( .A(n5724), .ZN(n5390) );
  AOI22_X1 U6559 ( .A1(n6175), .A2(n5390), .B1(n6241), .B2(
        PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5391) );
  OAI211_X1 U6560 ( .C1(n5393), .C2(n6210), .A(n5392), .B(n5391), .ZN(n5394)
         );
  AOI21_X1 U6561 ( .B1(n5911), .B2(n3100), .A(n5394), .ZN(n5395) );
  OAI21_X1 U6562 ( .B1(n5676), .B2(n6193), .A(n5395), .ZN(U2797) );
  AOI22_X1 U6563 ( .A1(n6175), .A2(n5729), .B1(n6241), .B2(
        PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6564 ( .A1(n6249), .A2(EBX_REG_29__SCAN_IN), .ZN(n5396) );
  OAI211_X1 U6565 ( .C1(n5914), .C2(n6244), .A(n5397), .B(n5396), .ZN(n5398)
         );
  INV_X1 U6566 ( .A(n5398), .ZN(n5401) );
  MUX2_X1 U6567 ( .A(n5399), .B(n5411), .S(REIP_REG_29__SCAN_IN), .Z(n5400) );
  OAI211_X1 U6568 ( .C1(n5679), .C2(n6193), .A(n5401), .B(n5400), .ZN(U2798)
         );
  NAND2_X2 U6569 ( .A1(n5404), .A2(n4449), .ZN(n5743) );
  OAI22_X1 U6570 ( .A1(n6259), .A2(n5405), .B1(n5745), .B2(n6258), .ZN(n5410)
         );
  AOI21_X1 U6571 ( .B1(n5407), .B2(n5419), .A(n5406), .ZN(n5928) );
  INV_X1 U6572 ( .A(n5928), .ZN(n5408) );
  NOR2_X1 U6573 ( .A1(n5408), .A2(n6244), .ZN(n5409) );
  AOI211_X1 U6574 ( .C1(EBX_REG_28__SCAN_IN), .C2(n6249), .A(n5410), .B(n5409), 
        .ZN(n5414) );
  NAND2_X1 U6575 ( .A1(n5425), .A2(REIP_REG_27__SCAN_IN), .ZN(n5412) );
  MUX2_X1 U6576 ( .A(n5412), .B(n5411), .S(REIP_REG_28__SCAN_IN), .Z(n5413) );
  OAI211_X1 U6577 ( .C1(n5743), .C2(n6193), .A(n5414), .B(n5413), .ZN(U2799)
         );
  AOI21_X1 U6578 ( .B1(n5416), .B2(n5415), .A(n5402), .ZN(n5755) );
  INV_X1 U6579 ( .A(n5755), .ZN(n5684) );
  NAND2_X1 U6580 ( .A1(n5431), .A2(n5417), .ZN(n5418) );
  NAND2_X1 U6581 ( .A1(n5419), .A2(n5418), .ZN(n5939) );
  INV_X1 U6582 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5646) );
  OAI21_X1 U6583 ( .B1(n6210), .B2(n5646), .A(n5420), .ZN(n5421) );
  AOI21_X1 U6584 ( .B1(n5436), .B2(REIP_REG_27__SCAN_IN), .A(n5421), .ZN(n5422) );
  OAI21_X1 U6585 ( .B1(n5939), .B2(n6244), .A(n5422), .ZN(n5423) );
  AOI21_X1 U6586 ( .B1(n5425), .B2(n5424), .A(n5423), .ZN(n5426) );
  OAI21_X1 U6587 ( .B1(n5684), .B2(n6193), .A(n5426), .ZN(U2800) );
  INV_X1 U6588 ( .A(n5415), .ZN(n5428) );
  INV_X1 U6589 ( .A(n5765), .ZN(n5687) );
  OAI21_X1 U6590 ( .B1(n5430), .B2(n5432), .A(n5431), .ZN(n5647) );
  INV_X1 U6591 ( .A(n5647), .ZN(n5949) );
  AOI22_X1 U6592 ( .A1(n6175), .A2(n5762), .B1(n6241), .B2(
        PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5433) );
  OAI21_X1 U6593 ( .B1(n6210), .B2(n5648), .A(n5433), .ZN(n5434) );
  AOI21_X1 U6594 ( .B1(n5949), .B2(n3100), .A(n5434), .ZN(n5439) );
  NOR3_X1 U6595 ( .A1(n5456), .A2(n5454), .A3(n5435), .ZN(n5437) );
  OAI21_X1 U6596 ( .B1(n5437), .B2(REIP_REG_26__SCAN_IN), .A(n5436), .ZN(n5438) );
  OAI211_X1 U6597 ( .C1(n5687), .C2(n6193), .A(n5439), .B(n5438), .ZN(U2801)
         );
  OAI21_X1 U6598 ( .B1(n3137), .B2(n5441), .A(n5440), .ZN(n5780) );
  INV_X1 U6599 ( .A(n5442), .ZN(n5444) );
  INV_X1 U6600 ( .A(n4461), .ZN(n5443) );
  AOI21_X1 U6601 ( .B1(n5444), .B2(n5443), .A(n5430), .ZN(n5649) );
  XNOR2_X1 U6602 ( .A(REIP_REG_24__SCAN_IN), .B(REIP_REG_25__SCAN_IN), .ZN(
        n5445) );
  NOR2_X1 U6603 ( .A1(n5456), .A2(n5445), .ZN(n5449) );
  NAND2_X1 U6604 ( .A1(n5467), .A2(REIP_REG_25__SCAN_IN), .ZN(n5447) );
  AOI22_X1 U6605 ( .A1(n6175), .A2(n5768), .B1(n6241), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5446) );
  OAI211_X1 U6606 ( .C1(n6959), .C2(n6210), .A(n5447), .B(n5446), .ZN(n5448)
         );
  AOI211_X1 U6607 ( .C1(n5649), .C2(n6166), .A(n5449), .B(n5448), .ZN(n5450)
         );
  OAI21_X1 U6608 ( .B1(n5780), .B2(n6193), .A(n5450), .ZN(U2802) );
  INV_X1 U6609 ( .A(n5467), .ZN(n5455) );
  OAI22_X1 U6610 ( .A1(n6259), .A2(n3189), .B1(n5451), .B2(n6258), .ZN(n5452)
         );
  AOI21_X1 U6611 ( .B1(n6249), .B2(EBX_REG_24__SCAN_IN), .A(n5452), .ZN(n5453)
         );
  OAI21_X1 U6612 ( .B1(n5455), .B2(n5454), .A(n5453), .ZN(n5458) );
  NOR2_X1 U6613 ( .A1(n5456), .A2(REIP_REG_24__SCAN_IN), .ZN(n5457) );
  AOI211_X1 U6614 ( .C1(n3100), .C2(n5650), .A(n5458), .B(n5457), .ZN(n5459)
         );
  OAI21_X1 U6615 ( .B1(n5692), .B2(n6193), .A(n5459), .ZN(U2803) );
  AND2_X1 U6616 ( .A1(n4441), .A2(n5460), .ZN(n5461) );
  NAND2_X1 U6617 ( .A1(n4485), .A2(n5462), .ZN(n5463) );
  AND2_X1 U6618 ( .A1(n4376), .A2(n5463), .ZN(n5967) );
  INV_X1 U6619 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5465) );
  AOI22_X1 U6620 ( .A1(n6175), .A2(n5791), .B1(n6241), .B2(
        PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5464) );
  OAI21_X1 U6621 ( .B1(n6210), .B2(n5465), .A(n5464), .ZN(n5466) );
  AOI21_X1 U6622 ( .B1(n5967), .B2(n3100), .A(n5466), .ZN(n5470) );
  INV_X1 U6623 ( .A(n5478), .ZN(n5486) );
  NOR3_X1 U6624 ( .A1(n5486), .A2(n5472), .A3(n5795), .ZN(n5468) );
  OAI21_X1 U6625 ( .B1(n5468), .B2(REIP_REG_23__SCAN_IN), .A(n5467), .ZN(n5469) );
  OAI211_X1 U6626 ( .C1(n5789), .C2(n6193), .A(n5470), .B(n5469), .ZN(U2804)
         );
  XOR2_X1 U6627 ( .A(REIP_REG_22__SCAN_IN), .B(REIP_REG_21__SCAN_IN), .Z(n5477) );
  OAI22_X1 U6628 ( .A1(n6259), .A2(n6988), .B1(n5471), .B2(n6258), .ZN(n5474)
         );
  NOR2_X1 U6629 ( .A1(n5501), .A2(n5472), .ZN(n5473) );
  AOI211_X1 U6630 ( .C1(EBX_REG_22__SCAN_IN), .C2(n6249), .A(n5474), .B(n5473), 
        .ZN(n5475) );
  OAI21_X1 U6631 ( .B1(n5653), .B2(n6244), .A(n5475), .ZN(n5476) );
  AOI21_X1 U6632 ( .B1(n5478), .B2(n5477), .A(n5476), .ZN(n5479) );
  OAI21_X1 U6633 ( .B1(n5697), .B2(n6193), .A(n5479), .ZN(U2805) );
  XNOR2_X1 U6634 ( .A(n4439), .B(n5480), .ZN(n5799) );
  INV_X1 U6635 ( .A(n5799), .ZN(n5700) );
  AOI21_X1 U6636 ( .B1(n5483), .B2(n5482), .A(n5481), .ZN(n5975) );
  OAI22_X1 U6637 ( .A1(n6259), .A2(n6983), .B1(n5797), .B2(n6258), .ZN(n5484)
         );
  AOI21_X1 U6638 ( .B1(n6249), .B2(EBX_REG_21__SCAN_IN), .A(n5484), .ZN(n5485)
         );
  OAI21_X1 U6639 ( .B1(n5501), .B2(n5795), .A(n5485), .ZN(n5488) );
  NOR2_X1 U6640 ( .A1(n5486), .A2(REIP_REG_21__SCAN_IN), .ZN(n5487) );
  AOI211_X1 U6641 ( .C1(n5975), .C2(n3100), .A(n5488), .B(n5487), .ZN(n5489)
         );
  OAI21_X1 U6642 ( .B1(n5700), .B2(n6193), .A(n5489), .ZN(U2806) );
  OAI21_X1 U6643 ( .B1(n5490), .B2(n5491), .A(n4439), .ZN(n5807) );
  OAI22_X1 U6644 ( .A1(n6259), .A2(n3187), .B1(n5803), .B2(n6258), .ZN(n5500)
         );
  INV_X1 U6645 ( .A(EBX_REG_18__SCAN_IN), .ZN(n6953) );
  AOI21_X1 U6646 ( .B1(n4329), .B2(n6953), .A(n5492), .ZN(n5496) );
  INV_X1 U6647 ( .A(n5493), .ZN(n5494) );
  NOR2_X1 U6648 ( .A1(n5494), .A2(n5510), .ZN(n5495) );
  MUX2_X1 U6649 ( .A(n4364), .B(n5496), .S(n5495), .Z(n5497) );
  XOR2_X1 U6650 ( .A(n5498), .B(n5497), .Z(n5991) );
  NOR2_X1 U6651 ( .A1(n5991), .A2(n6244), .ZN(n5499) );
  AOI211_X1 U6652 ( .C1(EBX_REG_20__SCAN_IN), .C2(n6249), .A(n5500), .B(n5499), 
        .ZN(n5505) );
  INV_X1 U6653 ( .A(n5501), .ZN(n5502) );
  OAI21_X1 U6654 ( .B1(n5503), .B2(REIP_REG_20__SCAN_IN), .A(n5502), .ZN(n5504) );
  OAI211_X1 U6655 ( .C1(n5807), .C2(n6193), .A(n5505), .B(n5504), .ZN(U2807)
         );
  XNOR2_X1 U6656 ( .A(REIP_REG_18__SCAN_IN), .B(REIP_REG_19__SCAN_IN), .ZN(
        n5522) );
  AOI21_X1 U6658 ( .B1(n5508), .B2(n5507), .A(n5490), .ZN(n5812) );
  NAND2_X1 U6659 ( .A1(n5812), .A2(n6204), .ZN(n5521) );
  INV_X1 U6660 ( .A(n5510), .ZN(n5511) );
  XNOR2_X1 U6661 ( .A(n5509), .B(n5511), .ZN(n5997) );
  OR2_X1 U6662 ( .A1(n5527), .A2(n5512), .ZN(n5518) );
  NAND2_X1 U6663 ( .A1(n6241), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5514)
         );
  NAND2_X1 U6664 ( .A1(n6184), .A2(n5513), .ZN(n6190) );
  OAI211_X1 U6665 ( .C1(n6258), .C2(n5810), .A(n5514), .B(n6190), .ZN(n5515)
         );
  INV_X1 U6666 ( .A(n5515), .ZN(n5517) );
  NAND2_X1 U6667 ( .A1(n6249), .A2(EBX_REG_19__SCAN_IN), .ZN(n5516) );
  OAI211_X1 U6668 ( .C1(n6253), .C2(n5518), .A(n5517), .B(n5516), .ZN(n5519)
         );
  AOI21_X1 U6669 ( .B1(n5997), .B2(n3100), .A(n5519), .ZN(n5520) );
  OAI211_X1 U6670 ( .C1(n5530), .C2(n5522), .A(n5521), .B(n5520), .ZN(U2808)
         );
  INV_X1 U6672 ( .A(n5524), .ZN(n5536) );
  OAI21_X1 U6673 ( .B1(n5536), .B2(n3837), .A(n5507), .ZN(n5822) );
  OAI21_X1 U6674 ( .B1(n5493), .B2(n5526), .A(n5509), .ZN(n6006) );
  INV_X1 U6675 ( .A(n6006), .ZN(n5533) );
  NOR2_X1 U6676 ( .A1(n6253), .A2(n5527), .ZN(n5540) );
  AOI21_X1 U6677 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5540), .A(n6227), .ZN(n5529) );
  AOI22_X1 U6678 ( .A1(n6175), .A2(n5819), .B1(n6241), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5528) );
  OAI211_X1 U6679 ( .C1(n6210), .C2(n6953), .A(n5529), .B(n5528), .ZN(n5532)
         );
  NOR2_X1 U6680 ( .A1(n5530), .A2(REIP_REG_18__SCAN_IN), .ZN(n5531) );
  AOI211_X1 U6681 ( .C1(n5533), .C2(n6166), .A(n5532), .B(n5531), .ZN(n5534)
         );
  OAI21_X1 U6682 ( .B1(n5822), .B2(n6193), .A(n5534), .ZN(U2809) );
  AOI21_X1 U6683 ( .B1(n5537), .B2(n5535), .A(n5536), .ZN(n5830) );
  NOR2_X1 U6684 ( .A1(n3139), .A2(n5538), .ZN(n5539) );
  OR2_X1 U6685 ( .A1(n5493), .A2(n5539), .ZN(n6007) );
  OAI21_X1 U6686 ( .B1(REIP_REG_17__SCAN_IN), .B2(n5541), .A(n5540), .ZN(n5547) );
  NOR2_X1 U6687 ( .A1(n6210), .A2(n5657), .ZN(n5545) );
  INV_X1 U6688 ( .A(n5826), .ZN(n5543) );
  NAND2_X1 U6689 ( .A1(n6241), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5542)
         );
  OAI211_X1 U6690 ( .C1(n6258), .C2(n5543), .A(n5542), .B(n6190), .ZN(n5544)
         );
  NOR2_X1 U6691 ( .A1(n5545), .A2(n5544), .ZN(n5546) );
  OAI211_X1 U6692 ( .C1(n6244), .C2(n6007), .A(n5547), .B(n5546), .ZN(n5548)
         );
  AOI21_X1 U6693 ( .B1(n5830), .B2(n6204), .A(n5548), .ZN(n5549) );
  INV_X1 U6694 ( .A(n5549), .ZN(U2810) );
  OAI21_X1 U6695 ( .B1(n5550), .B2(n5551), .A(n5535), .ZN(n5835) );
  AND2_X1 U6696 ( .A1(n5569), .A2(n5552), .ZN(n5553) );
  NOR2_X1 U6697 ( .A1(n3139), .A2(n5553), .ZN(n6028) );
  NAND2_X1 U6698 ( .A1(n6184), .A2(n5554), .ZN(n5555) );
  NAND2_X1 U6699 ( .A1(n6186), .A2(n5555), .ZN(n5587) );
  INV_X1 U6700 ( .A(n5838), .ZN(n5557) );
  NAND2_X1 U6701 ( .A1(n6241), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5556)
         );
  OAI211_X1 U6702 ( .C1(n6258), .C2(n5557), .A(n5556), .B(n6190), .ZN(n5560)
         );
  XNOR2_X1 U6703 ( .A(REIP_REG_16__SCAN_IN), .B(REIP_REG_15__SCAN_IN), .ZN(
        n5558) );
  NOR2_X1 U6704 ( .A1(n5575), .A2(n5558), .ZN(n5559) );
  AOI211_X1 U6705 ( .C1(EBX_REG_16__SCAN_IN), .C2(n6249), .A(n5560), .B(n5559), 
        .ZN(n5561) );
  OAI21_X1 U6706 ( .B1(n5562), .B2(n5587), .A(n5561), .ZN(n5563) );
  AOI21_X1 U6707 ( .B1(n6028), .B2(n3100), .A(n5563), .ZN(n5564) );
  OAI21_X1 U6708 ( .B1(n5835), .B2(n6193), .A(n5564), .ZN(U2811) );
  AND2_X1 U6709 ( .A1(n5565), .A2(n5566), .ZN(n5567) );
  OR2_X1 U6710 ( .A1(n5567), .A2(n5550), .ZN(n5846) );
  INV_X1 U6711 ( .A(n5569), .ZN(n5570) );
  AOI21_X1 U6712 ( .B1(n5571), .B2(n5568), .A(n5570), .ZN(n6038) );
  INV_X1 U6713 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5572) );
  OAI22_X1 U6714 ( .A1(n6210), .A2(n5572), .B1(n5842), .B2(n6258), .ZN(n5577)
         );
  AOI21_X1 U6715 ( .B1(n6241), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6227), 
        .ZN(n5573) );
  OAI221_X1 U6716 ( .B1(REIP_REG_15__SCAN_IN), .B2(n5575), .C1(n5574), .C2(
        n5587), .A(n5573), .ZN(n5576) );
  AOI211_X1 U6717 ( .C1(n6038), .C2(n6166), .A(n5577), .B(n5576), .ZN(n5578)
         );
  OAI21_X1 U6718 ( .B1(n5846), .B2(n6193), .A(n5578), .ZN(U2812) );
  OAI21_X1 U6719 ( .B1(n5668), .B2(n5580), .A(n5568), .ZN(n6055) );
  OAI21_X1 U6720 ( .B1(n5581), .B2(n5582), .A(n5565), .ZN(n5855) );
  INV_X1 U6721 ( .A(n5855), .ZN(n5583) );
  NAND2_X1 U6722 ( .A1(n5583), .A2(n6204), .ZN(n5591) );
  AOI21_X1 U6723 ( .B1(n6241), .B2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6227), 
        .ZN(n5584) );
  OAI21_X1 U6724 ( .B1(n5851), .B2(n6258), .A(n5584), .ZN(n5589) );
  NOR2_X1 U6725 ( .A1(n6144), .A2(n5585), .ZN(n6152) );
  AOI21_X1 U6726 ( .B1(n6152), .B2(REIP_REG_13__SCAN_IN), .A(
        REIP_REG_14__SCAN_IN), .ZN(n5586) );
  NOR2_X1 U6727 ( .A1(n5587), .A2(n5586), .ZN(n5588) );
  AOI211_X1 U6728 ( .C1(EBX_REG_14__SCAN_IN), .C2(n6249), .A(n5589), .B(n5588), 
        .ZN(n5590) );
  OAI211_X1 U6729 ( .C1(n6055), .C2(n6244), .A(n5591), .B(n5590), .ZN(U2813)
         );
  NAND3_X1 U6730 ( .A1(n6237), .A2(n5596), .A3(n5593), .ZN(n5592) );
  OAI21_X1 U6731 ( .B1(n6258), .B2(n5870), .A(n5592), .ZN(n5598) );
  INV_X1 U6732 ( .A(n6184), .ZN(n6236) );
  INV_X1 U6733 ( .A(n5593), .ZN(n5594) );
  OAI21_X1 U6734 ( .B1(n6236), .B2(n5594), .A(n6186), .ZN(n6143) );
  AOI22_X1 U6735 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6249), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6241), .ZN(n5595) );
  OAI211_X1 U6736 ( .C1(n5596), .C2(n6143), .A(n5595), .B(n6190), .ZN(n5597)
         );
  AOI211_X1 U6737 ( .C1(n6070), .C2(n6166), .A(n5598), .B(n5597), .ZN(n5599)
         );
  OAI21_X1 U6738 ( .B1(n5600), .B2(n6193), .A(n5599), .ZN(U2815) );
  NOR2_X1 U6740 ( .A1(n6144), .A2(n5612), .ZN(n5613) );
  NAND2_X1 U6741 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5613), .ZN(n5611) );
  OAI33_X1 U6742 ( .A1(1'b0), .A2(n6143), .A3(n5601), .B1(REIP_REG_11__SCAN_IN), .B2(n5614), .B3(n5611), .ZN(n5603) );
  INV_X1 U6743 ( .A(n5603), .ZN(n5607) );
  AOI22_X1 U6744 ( .A1(n6084), .A2(n6166), .B1(n6249), .B2(EBX_REG_11__SCAN_IN), .ZN(n5604) );
  OAI211_X1 U6745 ( .C1(n6259), .C2(n7047), .A(n5604), .B(n6190), .ZN(n5605)
         );
  AOI21_X1 U6746 ( .B1(n6175), .B2(n6329), .A(n5605), .ZN(n5606) );
  OAI211_X1 U6747 ( .C1(n6193), .C2(n6328), .A(n5607), .B(n5606), .ZN(U2816)
         );
  INV_X1 U6748 ( .A(n5875), .ZN(n5617) );
  AOI21_X1 U6749 ( .B1(n6241), .B2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6227), 
        .ZN(n5610) );
  OAI21_X1 U6750 ( .B1(n6163), .B2(n5608), .A(n5144), .ZN(n5673) );
  INV_X1 U6751 ( .A(n5673), .ZN(n6366) );
  AOI22_X1 U6752 ( .A1(n6366), .A2(n6166), .B1(n6249), .B2(EBX_REG_10__SCAN_IN), .ZN(n5609) );
  OAI211_X1 U6753 ( .C1(REIP_REG_10__SCAN_IN), .C2(n5611), .A(n5610), .B(n5609), .ZN(n5616) );
  OAI21_X1 U6754 ( .B1(n6236), .B2(n5612), .A(n6186), .ZN(n6180) );
  NAND2_X1 U6755 ( .A1(n5613), .A2(n6158), .ZN(n6168) );
  AOI21_X1 U6756 ( .B1(n6180), .B2(n6168), .A(n5614), .ZN(n5615) );
  AOI211_X1 U6757 ( .C1(n6175), .C2(n5617), .A(n5616), .B(n5615), .ZN(n5618)
         );
  OAI21_X1 U6758 ( .B1(n6193), .B2(n5879), .A(n5618), .ZN(U2817) );
  INV_X1 U6759 ( .A(n6187), .ZN(n5619) );
  AOI21_X1 U6760 ( .B1(n6237), .B2(n5619), .A(n6236), .ZN(n6229) );
  NOR2_X1 U6761 ( .A1(n6235), .A2(n5636), .ZN(n5620) );
  AOI21_X1 U6762 ( .B1(n6184), .B2(n5620), .A(REIP_REG_3__SCAN_IN), .ZN(n5635)
         );
  OR2_X1 U6763 ( .A1(n5628), .A2(n3402), .ZN(n5621) );
  NAND2_X1 U6764 ( .A1(n5622), .A2(n6255), .ZN(n5634) );
  INV_X1 U6765 ( .A(n5623), .ZN(n6425) );
  NAND2_X1 U6766 ( .A1(n6166), .A2(n6425), .ZN(n5632) );
  INV_X1 U6767 ( .A(n5624), .ZN(n5625) );
  AOI22_X1 U6768 ( .A1(n6175), .A2(n5625), .B1(n6241), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5631) );
  NAND2_X1 U6769 ( .A1(n6249), .A2(EBX_REG_3__SCAN_IN), .ZN(n5630) );
  INV_X1 U6770 ( .A(n5626), .ZN(n5627) );
  NOR2_X1 U6771 ( .A1(n5628), .A2(n5627), .ZN(n6248) );
  NAND2_X1 U6772 ( .A1(n6248), .A2(n4743), .ZN(n5629) );
  OAI211_X1 U6773 ( .C1(n6229), .C2(n5635), .A(n5634), .B(n5633), .ZN(U2824)
         );
  NAND2_X1 U6774 ( .A1(n6237), .A2(n5636), .ZN(n6239) );
  AOI22_X1 U6775 ( .A1(n6241), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6236), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5637) );
  OAI211_X1 U6776 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6258), .A(n6239), 
        .B(n5637), .ZN(n5640) );
  INV_X1 U6777 ( .A(n6248), .ZN(n6223) );
  OAI22_X1 U6778 ( .A1(n6223), .A2(n6099), .B1(n6210), .B2(n5638), .ZN(n5639)
         );
  AOI211_X1 U6779 ( .C1(n3100), .C2(n4819), .A(n5640), .B(n5639), .ZN(n5641)
         );
  OAI21_X1 U6780 ( .B1(n6214), .B2(n5642), .A(n5641), .ZN(U2826) );
  INV_X1 U6781 ( .A(n5904), .ZN(n5644) );
  OAI22_X1 U6782 ( .A1(n5644), .A2(n5672), .B1(n6266), .B2(n5643), .ZN(U2828)
         );
  AOI22_X1 U6783 ( .A1(n5928), .A2(n6261), .B1(EBX_REG_28__SCAN_IN), .B2(n5659), .ZN(n5645) );
  OAI21_X1 U6784 ( .B1(n5743), .B2(n5670), .A(n5645), .ZN(U2831) );
  OAI222_X1 U6785 ( .A1(n5670), .A2(n5684), .B1(n5646), .B2(n6266), .C1(n5939), 
        .C2(n5672), .ZN(U2832) );
  OAI222_X1 U6786 ( .A1(n5670), .A2(n5687), .B1(n5648), .B2(n6266), .C1(n5647), 
        .C2(n5672), .ZN(U2833) );
  INV_X1 U6787 ( .A(n5649), .ZN(n5960) );
  OAI222_X1 U6788 ( .A1(n5780), .A2(n5670), .B1(n6959), .B2(n6266), .C1(n5960), 
        .C2(n5672), .ZN(U2834) );
  AOI22_X1 U6789 ( .A1(n5650), .A2(n6261), .B1(EBX_REG_24__SCAN_IN), .B2(n5659), .ZN(n5651) );
  OAI21_X1 U6790 ( .B1(n5692), .B2(n5670), .A(n5651), .ZN(U2835) );
  AOI22_X1 U6791 ( .A1(n5967), .A2(n6261), .B1(EBX_REG_23__SCAN_IN), .B2(n5659), .ZN(n5652) );
  OAI21_X1 U6792 ( .B1(n5789), .B2(n5670), .A(n5652), .ZN(U2836) );
  OAI222_X1 U6793 ( .A1(n5670), .A2(n5697), .B1(n5654), .B2(n6266), .C1(n5653), 
        .C2(n5672), .ZN(U2837) );
  AOI22_X1 U6794 ( .A1(n5975), .A2(n6261), .B1(EBX_REG_21__SCAN_IN), .B2(n5659), .ZN(n5655) );
  OAI21_X1 U6795 ( .B1(n5700), .B2(n5670), .A(n5655), .ZN(U2838) );
  OAI222_X1 U6796 ( .A1(n5991), .A2(n5672), .B1(n6881), .B2(n6266), .C1(n5807), 
        .C2(n5670), .ZN(U2839) );
  INV_X1 U6797 ( .A(n5812), .ZN(n5705) );
  AOI22_X1 U6798 ( .A1(n5997), .A2(n6261), .B1(EBX_REG_19__SCAN_IN), .B2(n5659), .ZN(n5656) );
  OAI21_X1 U6799 ( .B1(n5705), .B2(n5670), .A(n5656), .ZN(U2840) );
  OAI222_X1 U6800 ( .A1(n5822), .A2(n5670), .B1(n6953), .B2(n6266), .C1(n6006), 
        .C2(n5672), .ZN(U2841) );
  INV_X1 U6801 ( .A(n5830), .ZN(n5710) );
  OAI222_X1 U6802 ( .A1(n5710), .A2(n5670), .B1(n5657), .B2(n6266), .C1(n6007), 
        .C2(n5672), .ZN(U2842) );
  AOI22_X1 U6803 ( .A1(n6028), .A2(n6261), .B1(EBX_REG_16__SCAN_IN), .B2(n5659), .ZN(n5658) );
  OAI21_X1 U6804 ( .B1(n5835), .B2(n5670), .A(n5658), .ZN(U2843) );
  AOI22_X1 U6805 ( .A1(n6038), .A2(n6261), .B1(EBX_REG_15__SCAN_IN), .B2(n5659), .ZN(n5660) );
  OAI21_X1 U6806 ( .B1(n5846), .B2(n5670), .A(n5660), .ZN(U2844) );
  OAI222_X1 U6807 ( .A1(n5855), .A2(n5670), .B1(n5661), .B2(n6266), .C1(n6055), 
        .C2(n5672), .ZN(U2845) );
  NAND2_X1 U6808 ( .A1(n5663), .A2(n5664), .ZN(n5665) );
  NAND2_X1 U6809 ( .A1(n5662), .A2(n5665), .ZN(n6153) );
  INV_X1 U6810 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5669) );
  NOR2_X1 U6811 ( .A1(n5363), .A2(n5666), .ZN(n5667) );
  OR2_X1 U6812 ( .A1(n5668), .A2(n5667), .ZN(n6145) );
  OAI222_X1 U6813 ( .A1(n6153), .A2(n5670), .B1(n5669), .B2(n6266), .C1(n6145), 
        .C2(n5672), .ZN(U2846) );
  OAI222_X1 U6814 ( .A1(n5673), .A2(n5672), .B1(n5671), .B2(n6266), .C1(n5879), 
        .C2(n5670), .ZN(U2849) );
  AOI22_X1 U6815 ( .A1(n5711), .A2(DATAI_30_), .B1(n5718), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5675) );
  NAND2_X1 U6816 ( .A1(n5712), .A2(DATAI_14_), .ZN(n5674) );
  OAI211_X1 U6817 ( .C1(n5676), .C2(n5721), .A(n5675), .B(n5674), .ZN(U2861)
         );
  AOI22_X1 U6818 ( .A1(n5711), .A2(DATAI_29_), .B1(n5718), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U6819 ( .A1(n5712), .A2(DATAI_13_), .ZN(n5677) );
  OAI211_X1 U6820 ( .C1(n5679), .C2(n5721), .A(n5678), .B(n5677), .ZN(U2862)
         );
  AOI22_X1 U6821 ( .A1(n5711), .A2(DATAI_28_), .B1(n5718), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5681) );
  NAND2_X1 U6822 ( .A1(n5712), .A2(DATAI_12_), .ZN(n5680) );
  OAI211_X1 U6823 ( .C1(n5743), .C2(n5721), .A(n5681), .B(n5680), .ZN(U2863)
         );
  AOI22_X1 U6824 ( .A1(n5711), .A2(DATAI_27_), .B1(n5718), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U6825 ( .A1(n5712), .A2(DATAI_11_), .ZN(n5682) );
  OAI211_X1 U6826 ( .C1(n5684), .C2(n5721), .A(n5683), .B(n5682), .ZN(U2864)
         );
  AOI22_X1 U6827 ( .A1(n5711), .A2(DATAI_26_), .B1(n5718), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U6828 ( .A1(n5712), .A2(DATAI_10_), .ZN(n5685) );
  OAI211_X1 U6829 ( .C1(n5687), .C2(n5721), .A(n5686), .B(n5685), .ZN(U2865)
         );
  AOI22_X1 U6830 ( .A1(n5711), .A2(DATAI_25_), .B1(n5718), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U6831 ( .A1(n5712), .A2(DATAI_9_), .ZN(n5688) );
  OAI211_X1 U6832 ( .C1(n5780), .C2(n5721), .A(n5689), .B(n5688), .ZN(U2866)
         );
  AOI22_X1 U6833 ( .A1(n5711), .A2(DATAI_24_), .B1(n5718), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5691) );
  NAND2_X1 U6834 ( .A1(n5712), .A2(DATAI_8_), .ZN(n5690) );
  OAI211_X1 U6835 ( .C1(n5692), .C2(n5721), .A(n5691), .B(n5690), .ZN(U2867)
         );
  AOI22_X1 U6836 ( .A1(n5711), .A2(DATAI_23_), .B1(n5718), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5694) );
  NAND2_X1 U6837 ( .A1(n5712), .A2(DATAI_7_), .ZN(n5693) );
  OAI211_X1 U6838 ( .C1(n5789), .C2(n5721), .A(n5694), .B(n5693), .ZN(U2868)
         );
  AOI22_X1 U6839 ( .A1(n5711), .A2(DATAI_22_), .B1(n5718), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5696) );
  NAND2_X1 U6840 ( .A1(n5712), .A2(DATAI_6_), .ZN(n5695) );
  OAI211_X1 U6841 ( .C1(n5697), .C2(n5721), .A(n5696), .B(n5695), .ZN(U2869)
         );
  AOI22_X1 U6842 ( .A1(n5711), .A2(DATAI_21_), .B1(n5718), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5699) );
  NAND2_X1 U6843 ( .A1(n5712), .A2(DATAI_5_), .ZN(n5698) );
  OAI211_X1 U6844 ( .C1(n5700), .C2(n5721), .A(n5699), .B(n5698), .ZN(U2870)
         );
  AOI22_X1 U6845 ( .A1(n5711), .A2(DATAI_20_), .B1(n5718), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U6846 ( .A1(n5712), .A2(DATAI_4_), .ZN(n5701) );
  OAI211_X1 U6847 ( .C1(n5807), .C2(n5721), .A(n5702), .B(n5701), .ZN(U2871)
         );
  AOI22_X1 U6848 ( .A1(n5711), .A2(DATAI_19_), .B1(n5718), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5704) );
  NAND2_X1 U6849 ( .A1(n5712), .A2(DATAI_3_), .ZN(n5703) );
  OAI211_X1 U6850 ( .C1(n5705), .C2(n5721), .A(n5704), .B(n5703), .ZN(U2872)
         );
  AOI22_X1 U6851 ( .A1(n5711), .A2(DATAI_18_), .B1(n5718), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U6852 ( .A1(n5712), .A2(DATAI_2_), .ZN(n5706) );
  OAI211_X1 U6853 ( .C1(n5822), .C2(n5721), .A(n5707), .B(n5706), .ZN(U2873)
         );
  AOI22_X1 U6854 ( .A1(n5711), .A2(DATAI_17_), .B1(n5718), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5709) );
  NAND2_X1 U6855 ( .A1(n5712), .A2(DATAI_1_), .ZN(n5708) );
  OAI211_X1 U6856 ( .C1(n5710), .C2(n5721), .A(n5709), .B(n5708), .ZN(U2874)
         );
  AOI22_X1 U6857 ( .A1(n5711), .A2(DATAI_16_), .B1(n5718), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5714) );
  NAND2_X1 U6858 ( .A1(n5712), .A2(DATAI_0_), .ZN(n5713) );
  OAI211_X1 U6859 ( .C1(n5835), .C2(n5721), .A(n5714), .B(n5713), .ZN(U2875)
         );
  INV_X1 U6860 ( .A(DATAI_15_), .ZN(n6894) );
  INV_X1 U6861 ( .A(EAX_REG_15__SCAN_IN), .ZN(n7020) );
  OAI222_X1 U6862 ( .A1(n5846), .A2(n5721), .B1(n6894), .B2(n5716), .C1(n5715), 
        .C2(n7020), .ZN(U2876) );
  AOI22_X1 U6863 ( .A1(n5719), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n5718), .ZN(n5717) );
  OAI21_X1 U6864 ( .B1(n5855), .B2(n5721), .A(n5717), .ZN(U2877) );
  AOI22_X1 U6865 ( .A1(n5719), .A2(DATAI_13_), .B1(EAX_REG_13__SCAN_IN), .B2(
        n5718), .ZN(n5720) );
  OAI21_X1 U6866 ( .B1(n6153), .B2(n5721), .A(n5720), .ZN(U2878) );
  NAND2_X1 U6867 ( .A1(n6433), .A2(REIP_REG_30__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U6868 ( .A1(n6354), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5723)
         );
  OAI211_X1 U6869 ( .C1(n6363), .C2(n5724), .A(n5907), .B(n5723), .ZN(n5725)
         );
  AOI21_X1 U6870 ( .B1(n5726), .B2(n6349), .A(n5725), .ZN(n5727) );
  OAI21_X1 U6871 ( .B1(n5913), .B2(n6334), .A(n5727), .ZN(U2956) );
  XNOR2_X1 U6872 ( .A(n5728), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5923)
         );
  NAND2_X1 U6873 ( .A1(n6330), .A2(n5729), .ZN(n5730) );
  NAND2_X1 U6874 ( .A1(n6433), .A2(REIP_REG_29__SCAN_IN), .ZN(n5917) );
  OAI211_X1 U6875 ( .C1(n5884), .C2(n5731), .A(n5730), .B(n5917), .ZN(n5732)
         );
  OAI21_X1 U6876 ( .B1(n5923), .B2(n6334), .A(n5734), .ZN(U2957) );
  INV_X1 U6877 ( .A(n5735), .ZN(n5742) );
  INV_X1 U6878 ( .A(n5736), .ZN(n5737) );
  AND2_X1 U6879 ( .A1(n5737), .A2(n5757), .ZN(n5749) );
  INV_X1 U6880 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5937) );
  NAND2_X1 U6881 ( .A1(n5937), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5740) );
  NAND3_X1 U6882 ( .A1(n5735), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n6878), .ZN(n5739) );
  OAI211_X1 U6883 ( .C1(n5749), .C2(n5740), .A(n5739), .B(n5738), .ZN(n5741)
         );
  INV_X1 U6884 ( .A(n5743), .ZN(n5747) );
  NAND2_X1 U6885 ( .A1(n6433), .A2(REIP_REG_28__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U6886 ( .A1(n6354), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5744)
         );
  OAI211_X1 U6887 ( .C1(n6363), .C2(n5745), .A(n5924), .B(n5744), .ZN(n5746)
         );
  OAI21_X1 U6888 ( .B1(n5931), .B2(n6334), .A(n5748), .ZN(U2958) );
  NOR2_X1 U6889 ( .A1(n5735), .A2(n5749), .ZN(n5750) );
  XNOR2_X1 U6890 ( .A(n5750), .B(n5937), .ZN(n5943) );
  NAND2_X1 U6891 ( .A1(n6330), .A2(n5751), .ZN(n5752) );
  NAND2_X1 U6892 ( .A1(n6433), .A2(REIP_REG_27__SCAN_IN), .ZN(n5932) );
  OAI211_X1 U6893 ( .C1(n5884), .C2(n5753), .A(n5752), .B(n5932), .ZN(n5754)
         );
  AOI21_X1 U6894 ( .B1(n5755), .B2(n6349), .A(n5754), .ZN(n5756) );
  OAI21_X1 U6895 ( .B1(n5943), .B2(n6334), .A(n5756), .ZN(U2959) );
  INV_X1 U6896 ( .A(n5757), .ZN(n5759) );
  NAND2_X1 U6897 ( .A1(n5759), .A2(n5758), .ZN(n5761) );
  XOR2_X1 U6898 ( .A(n5761), .B(n5760), .Z(n5951) );
  NAND2_X1 U6899 ( .A1(n6330), .A2(n5762), .ZN(n5763) );
  NAND2_X1 U6900 ( .A1(n6433), .A2(REIP_REG_26__SCAN_IN), .ZN(n5946) );
  OAI211_X1 U6901 ( .C1(n5884), .C2(n6853), .A(n5763), .B(n5946), .ZN(n5764)
         );
  AOI21_X1 U6902 ( .B1(n5765), .B2(n6349), .A(n5764), .ZN(n5766) );
  OAI21_X1 U6903 ( .B1(n5951), .B2(n6334), .A(n5766), .ZN(U2960) );
  NAND2_X1 U6904 ( .A1(n6433), .A2(REIP_REG_25__SCAN_IN), .ZN(n5954) );
  OAI21_X1 U6905 ( .B1(n5884), .B2(n6906), .A(n5954), .ZN(n5767) );
  AOI21_X1 U6906 ( .B1(n6330), .B2(n5768), .A(n5767), .ZN(n5779) );
  NAND3_X1 U6907 ( .A1(n5771), .A2(n5770), .A3(n5986), .ZN(n5776) );
  INV_X1 U6908 ( .A(n5769), .ZN(n5773) );
  OAI21_X1 U6909 ( .B1(n5773), .B2(n5772), .A(n3107), .ZN(n5775) );
  XNOR2_X1 U6910 ( .A(n5848), .B(n6913), .ZN(n5774) );
  OAI211_X1 U6911 ( .C1(n5769), .C2(n5776), .A(n5775), .B(n5774), .ZN(n5777)
         );
  NAND2_X1 U6912 ( .A1(n5777), .A2(n5736), .ZN(n5952) );
  NAND2_X1 U6913 ( .A1(n5952), .A2(n6358), .ZN(n5778) );
  OAI211_X1 U6914 ( .C1(n5780), .C2(n5888), .A(n5779), .B(n5778), .ZN(U2961)
         );
  NAND2_X1 U6915 ( .A1(n3106), .A2(n5781), .ZN(n5782) );
  OR2_X1 U6916 ( .A1(n5783), .A2(n5782), .ZN(n5784) );
  XNOR2_X1 U6917 ( .A(n5787), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5969)
         );
  NAND2_X1 U6918 ( .A1(n6433), .A2(REIP_REG_23__SCAN_IN), .ZN(n5961) );
  OAI21_X1 U6919 ( .B1(n5884), .B2(n5788), .A(n5961), .ZN(n5790) );
  AOI21_X1 U6920 ( .B1(n5794), .B2(n5793), .A(n5792), .ZN(n5977) );
  NOR2_X1 U6921 ( .A1(n6423), .A2(n5795), .ZN(n5970) );
  AOI21_X1 U6922 ( .B1(n6354), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5970), 
        .ZN(n5796) );
  OAI21_X1 U6923 ( .B1(n5797), .B2(n6363), .A(n5796), .ZN(n5798) );
  AOI21_X1 U6924 ( .B1(n5799), .B2(n6349), .A(n5798), .ZN(n5800) );
  OAI21_X1 U6925 ( .B1(n5977), .B2(n6334), .A(n5800), .ZN(U2965) );
  XNOR2_X1 U6926 ( .A(n5802), .B(n5801), .ZN(n5978) );
  NAND2_X1 U6927 ( .A1(n5978), .A2(n6358), .ZN(n5806) );
  NOR2_X1 U6928 ( .A1(n6423), .A2(n4588), .ZN(n5988) );
  NOR2_X1 U6929 ( .A1(n6363), .A2(n5803), .ZN(n5804) );
  AOI211_X1 U6930 ( .C1(n6354), .C2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5988), 
        .B(n5804), .ZN(n5805) );
  OAI211_X1 U6931 ( .C1(n5888), .C2(n5807), .A(n5806), .B(n5805), .ZN(U2966)
         );
  XNOR2_X1 U6932 ( .A(n5769), .B(n5808), .ZN(n5999) );
  NAND2_X1 U6933 ( .A1(n6433), .A2(REIP_REG_19__SCAN_IN), .ZN(n5993) );
  NAND2_X1 U6934 ( .A1(n6354), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5809)
         );
  OAI211_X1 U6935 ( .C1(n6363), .C2(n5810), .A(n5993), .B(n5809), .ZN(n5811)
         );
  AOI21_X1 U6936 ( .B1(n5812), .B2(n6349), .A(n5811), .ZN(n5813) );
  OAI21_X1 U6937 ( .B1(n5999), .B2(n6334), .A(n5813), .ZN(U2967) );
  NAND3_X1 U6938 ( .A1(n5833), .A2(n4229), .A3(n6022), .ZN(n5823) );
  NAND3_X1 U6939 ( .A1(n5814), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5848), .ZN(n5824) );
  MUX2_X1 U6940 ( .A(n5823), .B(n5824), .S(INSTADDRPOINTER_REG_17__SCAN_IN), 
        .Z(n5815) );
  XNOR2_X1 U6941 ( .A(n5815), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6000)
         );
  NAND2_X1 U6942 ( .A1(n6000), .A2(n6358), .ZN(n5821) );
  NOR2_X1 U6943 ( .A1(n6423), .A2(n5816), .ZN(n6002) );
  NOR2_X1 U6944 ( .A1(n5884), .A2(n5817), .ZN(n5818) );
  AOI211_X1 U6945 ( .C1(n6330), .C2(n5819), .A(n6002), .B(n5818), .ZN(n5820)
         );
  OAI211_X1 U6946 ( .C1(n5888), .C2(n5822), .A(n5821), .B(n5820), .ZN(U2968)
         );
  NAND2_X1 U6947 ( .A1(n5824), .A2(n5823), .ZN(n5825) );
  XNOR2_X1 U6948 ( .A(n5825), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6016)
         );
  NAND2_X1 U6949 ( .A1(n6330), .A2(n5826), .ZN(n5827) );
  NAND2_X1 U6950 ( .A1(n6433), .A2(REIP_REG_17__SCAN_IN), .ZN(n6009) );
  OAI211_X1 U6951 ( .C1(n5884), .C2(n5828), .A(n5827), .B(n6009), .ZN(n5829)
         );
  AOI21_X1 U6952 ( .B1(n5830), .B2(n6349), .A(n5829), .ZN(n5831) );
  OAI21_X1 U6953 ( .B1(n6016), .B2(n6334), .A(n5831), .ZN(U2969) );
  XNOR2_X1 U6954 ( .A(n5848), .B(n6022), .ZN(n5832) );
  XNOR2_X1 U6955 ( .A(n5833), .B(n5832), .ZN(n6030) );
  NAND2_X1 U6956 ( .A1(n6433), .A2(REIP_REG_16__SCAN_IN), .ZN(n6024) );
  OAI21_X1 U6957 ( .B1(n5884), .B2(n5834), .A(n6024), .ZN(n5837) );
  NOR2_X1 U6958 ( .A1(n5835), .A2(n5888), .ZN(n5836) );
  AOI211_X1 U6959 ( .C1(n6330), .C2(n5838), .A(n5837), .B(n5836), .ZN(n5839)
         );
  OAI21_X1 U6960 ( .B1(n6334), .B2(n6030), .A(n5839), .ZN(U2970) );
  XNOR2_X1 U6961 ( .A(n5848), .B(n6035), .ZN(n5840) );
  XNOR2_X1 U6962 ( .A(n5841), .B(n5840), .ZN(n6031) );
  NAND2_X1 U6963 ( .A1(n6031), .A2(n6358), .ZN(n5845) );
  AND2_X1 U6964 ( .A1(n6433), .A2(REIP_REG_15__SCAN_IN), .ZN(n6032) );
  NOR2_X1 U6965 ( .A1(n6363), .A2(n5842), .ZN(n5843) );
  AOI211_X1 U6966 ( .C1(n6354), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6032), 
        .B(n5843), .ZN(n5844) );
  OAI211_X1 U6967 ( .C1(n5888), .C2(n5846), .A(n5845), .B(n5844), .ZN(U2971)
         );
  XNOR2_X1 U6968 ( .A(n5848), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5849)
         );
  XNOR2_X1 U6969 ( .A(n5847), .B(n5849), .ZN(n6041) );
  NAND2_X1 U6970 ( .A1(n6041), .A2(n6358), .ZN(n5854) );
  NOR2_X1 U6971 ( .A1(n6423), .A2(n5850), .ZN(n6052) );
  NOR2_X1 U6972 ( .A1(n6363), .A2(n5851), .ZN(n5852) );
  AOI211_X1 U6973 ( .C1(n6354), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6052), 
        .B(n5852), .ZN(n5853) );
  OAI211_X1 U6974 ( .C1(n5888), .C2(n5855), .A(n5854), .B(n5853), .ZN(U2972)
         );
  XNOR2_X1 U6975 ( .A(n5856), .B(n5857), .ZN(n6056) );
  NAND2_X1 U6976 ( .A1(n6056), .A2(n6358), .ZN(n5860) );
  AND2_X1 U6977 ( .A1(n6433), .A2(REIP_REG_13__SCAN_IN), .ZN(n6059) );
  NOR2_X1 U6978 ( .A1(n6363), .A2(n6157), .ZN(n5858) );
  AOI211_X1 U6979 ( .C1(n6354), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6059), 
        .B(n5858), .ZN(n5859) );
  OAI211_X1 U6980 ( .C1(n5888), .C2(n6153), .A(n5860), .B(n5859), .ZN(U2973)
         );
  NOR2_X1 U6981 ( .A1(n3107), .A2(n6364), .ZN(n5882) );
  AOI21_X1 U6982 ( .B1(n5861), .B2(n5880), .A(n5882), .ZN(n6073) );
  NAND2_X1 U6983 ( .A1(n6073), .A2(n5862), .ZN(n6075) );
  OAI21_X1 U6984 ( .B1(n6075), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n4229), 
        .ZN(n5863) );
  OAI21_X1 U6985 ( .B1(n6073), .B2(n5864), .A(n5863), .ZN(n5868) );
  INV_X1 U6986 ( .A(n5865), .ZN(n5866) );
  AOI21_X1 U6987 ( .B1(n4229), .B2(INSTADDRPOINTER_REG_12__SCAN_IN), .A(n5866), 
        .ZN(n5867) );
  XNOR2_X1 U6988 ( .A(n5868), .B(n5867), .ZN(n6072) );
  AND2_X1 U6989 ( .A1(n6433), .A2(REIP_REG_12__SCAN_IN), .ZN(n6069) );
  AOI21_X1 U6990 ( .B1(n6354), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6069), 
        .ZN(n5869) );
  OAI21_X1 U6991 ( .B1(n5870), .B2(n6363), .A(n5869), .ZN(n5871) );
  AOI21_X1 U6992 ( .B1(n5872), .B2(n6349), .A(n5871), .ZN(n5873) );
  OAI21_X1 U6993 ( .B1(n6072), .B2(n6334), .A(n5873), .ZN(U2974) );
  XNOR2_X1 U6994 ( .A(n3107), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5874)
         );
  XNOR2_X1 U6995 ( .A(n6073), .B(n5874), .ZN(n6369) );
  NAND2_X1 U6996 ( .A1(n6369), .A2(n6358), .ZN(n5878) );
  NOR2_X1 U6997 ( .A1(n6423), .A2(n5614), .ZN(n6365) );
  NOR2_X1 U6998 ( .A1(n6363), .A2(n5875), .ZN(n5876) );
  AOI211_X1 U6999 ( .C1(n6354), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6365), 
        .B(n5876), .ZN(n5877) );
  OAI211_X1 U7000 ( .C1(n5888), .C2(n5879), .A(n5878), .B(n5877), .ZN(U2976)
         );
  INV_X1 U7001 ( .A(n5880), .ZN(n5881) );
  NOR2_X1 U7002 ( .A1(n5882), .A2(n5881), .ZN(n5883) );
  XOR2_X1 U7003 ( .A(n5883), .B(n5861), .Z(n6377) );
  NAND2_X1 U7004 ( .A1(n6377), .A2(n6358), .ZN(n5887) );
  NAND2_X1 U7005 ( .A1(n6433), .A2(REIP_REG_9__SCAN_IN), .ZN(n6373) );
  OAI21_X1 U7006 ( .B1(n5884), .B2(n6159), .A(n6373), .ZN(n5885) );
  AOI21_X1 U7007 ( .B1(n6330), .B2(n6162), .A(n5885), .ZN(n5886) );
  OAI211_X1 U7008 ( .C1(n5888), .C2(n6161), .A(n5887), .B(n5886), .ZN(U2977)
         );
  OAI21_X1 U7009 ( .B1(n5891), .B2(n5890), .A(n5889), .ZN(n6097) );
  NOR2_X1 U7010 ( .A1(n6423), .A2(n6974), .ZN(n6094) );
  AOI21_X1 U7011 ( .B1(n6354), .B2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6094), 
        .ZN(n5892) );
  OAI21_X1 U7012 ( .B1(n6174), .B2(n6363), .A(n5892), .ZN(n5893) );
  AOI21_X1 U7013 ( .B1(n6177), .B2(n6349), .A(n5893), .ZN(n5894) );
  OAI21_X1 U7014 ( .B1(n6097), .B2(n6334), .A(n5894), .ZN(U2978) );
  INV_X1 U7015 ( .A(n5896), .ZN(n5897) );
  NAND2_X1 U7016 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5898) );
  NOR2_X1 U7017 ( .A1(n5953), .A2(n5898), .ZN(n5938) );
  NAND3_X1 U7018 ( .A1(n5938), .A2(n5916), .A3(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U7019 ( .A1(n7051), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5902) );
  NOR2_X1 U7020 ( .A1(n5944), .A2(n5898), .ZN(n5933) );
  NOR2_X1 U7021 ( .A1(n5944), .A2(n6394), .ZN(n5934) );
  AOI21_X1 U7022 ( .B1(n5916), .B2(n5933), .A(n5934), .ZN(n5915) );
  AOI21_X1 U7023 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .A(n6368), .ZN(n5899) );
  OAI21_X1 U7024 ( .B1(n5915), .B2(n5899), .A(INSTADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n5900) );
  OAI211_X1 U7025 ( .C1(n5909), .C2(n5902), .A(n5901), .B(n5900), .ZN(n5903)
         );
  AOI21_X1 U7026 ( .B1(n5904), .B2(n6435), .A(n5903), .ZN(n5905) );
  OAI21_X1 U7027 ( .B1(n5895), .B2(n6412), .A(n5905), .ZN(U2987) );
  INV_X1 U7028 ( .A(n5934), .ZN(n5906) );
  OAI211_X1 U7029 ( .C1(n5915), .C2(n3173), .A(INSTADDRPOINTER_REG_30__SCAN_IN), .B(n5906), .ZN(n5908) );
  OAI211_X1 U7030 ( .C1(n5909), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5908), .B(n5907), .ZN(n5910) );
  AOI21_X1 U7031 ( .B1(n5911), .B2(n6435), .A(n5910), .ZN(n5912) );
  INV_X1 U7032 ( .A(n5914), .ZN(n5921) );
  INV_X1 U7033 ( .A(n5915), .ZN(n5919) );
  NAND3_X1 U7034 ( .A1(n5938), .A2(n5916), .A3(n3173), .ZN(n5918) );
  OAI211_X1 U7035 ( .C1(n5919), .C2(n3173), .A(n5918), .B(n5917), .ZN(n5920)
         );
  AOI21_X1 U7036 ( .B1(n5921), .B2(n6435), .A(n5920), .ZN(n5922) );
  OAI21_X1 U7037 ( .B1(n5923), .B2(n6412), .A(n5922), .ZN(U2989) );
  XNOR2_X1 U7038 ( .A(n6878), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5927)
         );
  INV_X1 U7039 ( .A(n5924), .ZN(n5926) );
  NOR3_X1 U7040 ( .A1(n5934), .A2(n5933), .A3(n6878), .ZN(n5925) );
  AOI211_X1 U7041 ( .C1(n5938), .C2(n5927), .A(n5926), .B(n5925), .ZN(n5930)
         );
  NAND2_X1 U7042 ( .A1(n5928), .A2(n6435), .ZN(n5929) );
  OAI211_X1 U7043 ( .C1(n5931), .C2(n6412), .A(n5930), .B(n5929), .ZN(U2990)
         );
  INV_X1 U7044 ( .A(n5932), .ZN(n5936) );
  NOR3_X1 U7045 ( .A1(n5934), .A2(n5933), .A3(n5937), .ZN(n5935) );
  AOI211_X1 U7046 ( .C1(n5938), .C2(n5937), .A(n5936), .B(n5935), .ZN(n5942)
         );
  INV_X1 U7047 ( .A(n5939), .ZN(n5940) );
  NAND2_X1 U7048 ( .A1(n5940), .A2(n6435), .ZN(n5941) );
  OAI211_X1 U7049 ( .C1(n5943), .C2(n6412), .A(n5942), .B(n5941), .ZN(U2991)
         );
  XNOR2_X1 U7050 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5947) );
  NAND2_X1 U7051 ( .A1(n5944), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5945) );
  OAI211_X1 U7052 ( .C1(n5953), .C2(n5947), .A(n5946), .B(n5945), .ZN(n5948)
         );
  AOI21_X1 U7053 ( .B1(n5949), .B2(n6435), .A(n5948), .ZN(n5950) );
  OAI21_X1 U7054 ( .B1(n5951), .B2(n6412), .A(n5950), .ZN(U2992) );
  NAND2_X1 U7055 ( .A1(n5952), .A2(n6440), .ZN(n5959) );
  INV_X1 U7056 ( .A(n5953), .ZN(n5957) );
  OAI21_X1 U7057 ( .B1(n5955), .B2(n6913), .A(n5954), .ZN(n5956) );
  AOI21_X1 U7058 ( .B1(n5957), .B2(n6913), .A(n5956), .ZN(n5958) );
  OAI211_X1 U7059 ( .C1(n6397), .C2(n5960), .A(n5959), .B(n5958), .ZN(U2993)
         );
  INV_X1 U7060 ( .A(n5961), .ZN(n5962) );
  AOI21_X1 U7061 ( .B1(n5963), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n5962), 
        .ZN(n5964) );
  OAI21_X1 U7062 ( .B1(n5965), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n5964), 
        .ZN(n5966) );
  AOI21_X1 U7063 ( .B1(n5967), .B2(n6435), .A(n5966), .ZN(n5968) );
  OAI21_X1 U7064 ( .B1(n5969), .B2(n6412), .A(n5968), .ZN(U2995) );
  AOI21_X1 U7065 ( .B1(n5971), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5970), 
        .ZN(n5972) );
  OAI21_X1 U7066 ( .B1(n5973), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5972), 
        .ZN(n5974) );
  AOI21_X1 U7067 ( .B1(n5975), .B2(n6435), .A(n5974), .ZN(n5976) );
  OAI21_X1 U7068 ( .B1(n5977), .B2(n6412), .A(n5976), .ZN(U2997) );
  NAND2_X1 U7069 ( .A1(n5978), .A2(n6440), .ZN(n5990) );
  OR2_X1 U7070 ( .A1(n6392), .A2(n5979), .ZN(n5982) );
  OAI21_X1 U7071 ( .B1(n6010), .B2(n5980), .A(n6017), .ZN(n5981) );
  AND2_X1 U7072 ( .A1(n5982), .A2(n5981), .ZN(n6011) );
  OAI21_X1 U7073 ( .B1(n5983), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n6011), 
        .ZN(n6003) );
  INV_X1 U7074 ( .A(n6003), .ZN(n5984) );
  OAI21_X1 U7075 ( .B1(n6368), .B2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n5984), 
        .ZN(n5992) );
  NOR3_X1 U7076 ( .A1(n5995), .A2(n5986), .A3(n5985), .ZN(n5987) );
  AOI211_X1 U7077 ( .C1(INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n5992), .A(n5988), .B(n5987), .ZN(n5989) );
  OAI211_X1 U7078 ( .C1(n6397), .C2(n5991), .A(n5990), .B(n5989), .ZN(U2998)
         );
  NAND2_X1 U7079 ( .A1(n5992), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5994) );
  OAI211_X1 U7080 ( .C1(n5995), .C2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5994), .B(n5993), .ZN(n5996) );
  AOI21_X1 U7081 ( .B1(n5997), .B2(n6435), .A(n5996), .ZN(n5998) );
  OAI21_X1 U7082 ( .B1(n5999), .B2(n6412), .A(n5998), .ZN(U2999) );
  NAND2_X1 U7083 ( .A1(n6000), .A2(n6440), .ZN(n6005) );
  NOR3_X1 U7084 ( .A1(n6008), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n6010), 
        .ZN(n6001) );
  AOI211_X1 U7085 ( .C1(INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n6003), .A(n6002), .B(n6001), .ZN(n6004) );
  OAI211_X1 U7086 ( .C1(n6397), .C2(n6006), .A(n6005), .B(n6004), .ZN(U3000)
         );
  INV_X1 U7087 ( .A(n6007), .ZN(n6014) );
  NOR2_X1 U7088 ( .A1(n6008), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6013)
         );
  OAI21_X1 U7089 ( .B1(n6011), .B2(n6010), .A(n6009), .ZN(n6012) );
  AOI211_X1 U7090 ( .C1(n6014), .C2(n6435), .A(n6013), .B(n6012), .ZN(n6015)
         );
  OAI21_X1 U7091 ( .B1(n6016), .B2(n6412), .A(n6015), .ZN(U3001) );
  NAND3_X1 U7092 ( .A1(n6079), .A2(n6023), .A3(n6035), .ZN(n6034) );
  INV_X1 U7093 ( .A(n6023), .ZN(n6021) );
  NAND2_X1 U7094 ( .A1(n6017), .A2(n6045), .ZN(n6020) );
  OR2_X1 U7095 ( .A1(n6392), .A2(n6018), .ZN(n6019) );
  NAND2_X1 U7096 ( .A1(n6020), .A2(n6019), .ZN(n6042) );
  AOI21_X1 U7097 ( .B1(n6021), .B2(n6394), .A(n6042), .ZN(n6036) );
  AOI21_X1 U7098 ( .B1(n6034), .B2(n6036), .A(n6022), .ZN(n6027) );
  NAND4_X1 U7099 ( .A1(n6079), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n6023), .A4(n6022), .ZN(n6025) );
  NAND2_X1 U7100 ( .A1(n6025), .A2(n6024), .ZN(n6026) );
  AOI211_X1 U7101 ( .C1(n6028), .C2(n6435), .A(n6027), .B(n6026), .ZN(n6029)
         );
  OAI21_X1 U7102 ( .B1(n6030), .B2(n6412), .A(n6029), .ZN(U3002) );
  INV_X1 U7103 ( .A(n6031), .ZN(n6040) );
  INV_X1 U7104 ( .A(n6032), .ZN(n6033) );
  OAI211_X1 U7105 ( .C1(n6036), .C2(n6035), .A(n6034), .B(n6033), .ZN(n6037)
         );
  AOI21_X1 U7106 ( .B1(n6038), .B2(n6435), .A(n6037), .ZN(n6039) );
  OAI21_X1 U7107 ( .B1(n6040), .B2(n6412), .A(n6039), .ZN(U3003) );
  NAND2_X1 U7108 ( .A1(n6041), .A2(n6440), .ZN(n6054) );
  NAND2_X1 U7109 ( .A1(n6394), .A2(n6064), .ZN(n6043) );
  INV_X1 U7110 ( .A(n6042), .ZN(n6082) );
  OAI211_X1 U7111 ( .C1(INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n6044), .A(n6043), .B(n6082), .ZN(n6060) );
  INV_X1 U7112 ( .A(n6045), .ZN(n6048) );
  OAI21_X1 U7113 ( .B1(n6048), .B2(n6047), .A(n6046), .ZN(n6050) );
  AOI21_X1 U7114 ( .B1(n6079), .B2(INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6049) );
  AOI211_X1 U7115 ( .C1(INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n6050), .A(n6064), .B(n6049), .ZN(n6051) );
  AOI211_X1 U7116 ( .C1(INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n6060), .A(n6052), .B(n6051), .ZN(n6053) );
  OAI211_X1 U7117 ( .C1(n6397), .C2(n6055), .A(n6054), .B(n6053), .ZN(U3004)
         );
  NAND2_X1 U7118 ( .A1(n6056), .A2(n6440), .ZN(n6062) );
  INV_X1 U7119 ( .A(n6079), .ZN(n6057) );
  NOR3_X1 U7120 ( .A1(n6057), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n6064), 
        .ZN(n6058) );
  AOI211_X1 U7121 ( .C1(INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n6060), .A(n6059), .B(n6058), .ZN(n6061) );
  OAI211_X1 U7122 ( .C1(n6397), .C2(n6145), .A(n6062), .B(n6061), .ZN(U3005)
         );
  INV_X1 U7123 ( .A(n6063), .ZN(n6065) );
  OAI21_X1 U7124 ( .B1(n6065), .B2(n6436), .A(n6064), .ZN(n6067) );
  AOI21_X1 U7125 ( .B1(n6079), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6066) );
  AOI21_X1 U7126 ( .B1(n6082), .B2(n6067), .A(n6066), .ZN(n6068) );
  AOI211_X1 U7127 ( .C1(n6070), .C2(n6435), .A(n6069), .B(n6068), .ZN(n6071)
         );
  OAI21_X1 U7128 ( .B1(n6072), .B2(n6412), .A(n6071), .ZN(U3006) );
  INV_X1 U7129 ( .A(n6073), .ZN(n6074) );
  AOI22_X1 U7130 ( .A1(n4229), .A2(n6075), .B1(n6074), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6078) );
  XNOR2_X1 U7131 ( .A(n3106), .B(n6081), .ZN(n6077) );
  XNOR2_X1 U7132 ( .A(n6078), .B(n6077), .ZN(n6335) );
  NAND2_X1 U7133 ( .A1(n6079), .A2(n6081), .ZN(n6080) );
  NAND2_X1 U7134 ( .A1(n6433), .A2(REIP_REG_11__SCAN_IN), .ZN(n6326) );
  OAI211_X1 U7135 ( .C1(n6082), .C2(n6081), .A(n6080), .B(n6326), .ZN(n6083)
         );
  AOI21_X1 U7136 ( .B1(n6084), .B2(n6435), .A(n6083), .ZN(n6085) );
  OAI21_X1 U7137 ( .B1(n6335), .B2(n6412), .A(n6085), .ZN(U3007) );
  INV_X1 U7138 ( .A(n6172), .ZN(n6095) );
  OAI221_X1 U7139 ( .B1(n6437), .B2(n6436), .C1(n6443), .C2(n6436), .A(n6086), 
        .ZN(n6431) );
  INV_X1 U7140 ( .A(n6431), .ZN(n6403) );
  NAND2_X1 U7141 ( .A1(n6087), .A2(n6403), .ZN(n6402) );
  NOR2_X1 U7142 ( .A1(n6401), .A2(n6402), .ZN(n6386) );
  OAI21_X1 U7143 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6386), .ZN(n6092) );
  INV_X1 U7144 ( .A(n6088), .ZN(n6089) );
  OAI22_X1 U7145 ( .A1(n6436), .A2(n6391), .B1(n6392), .B2(n6089), .ZN(n6090)
         );
  AOI21_X1 U7146 ( .B1(n6436), .B2(n6091), .A(n6090), .ZN(n6390) );
  OAI22_X1 U7147 ( .A1(n6367), .A2(n6092), .B1(n6390), .B2(n6858), .ZN(n6093)
         );
  AOI211_X1 U7148 ( .C1(n6435), .C2(n6095), .A(n6094), .B(n6093), .ZN(n6096)
         );
  OAI21_X1 U7149 ( .B1(n6412), .B2(n6097), .A(n6096), .ZN(U3010) );
  NAND2_X1 U7150 ( .A1(n4888), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6595) );
  OAI211_X1 U7151 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n4888), .A(n6595), .B(
        n6594), .ZN(n6098) );
  OAI21_X1 U7152 ( .B1(n6106), .B2(n6099), .A(n6098), .ZN(n6100) );
  MUX2_X1 U7153 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n6100), .S(n6448), 
        .Z(U3464) );
  XNOR2_X1 U7154 ( .A(n6452), .B(n6595), .ZN(n6102) );
  OAI22_X1 U7155 ( .A1(n6102), .A2(n6655), .B1(n6101), .B2(n6106), .ZN(n6103)
         );
  MUX2_X1 U7156 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n6103), .S(n6448), 
        .Z(U3463) );
  INV_X1 U7157 ( .A(n5028), .ZN(n6108) );
  NOR2_X1 U7158 ( .A1(n6104), .A2(n6595), .ZN(n6529) );
  NOR3_X1 U7159 ( .A1(n6105), .A2(n6593), .A3(n6529), .ZN(n6107) );
  OAI222_X1 U7160 ( .A1(n6109), .A2(n6108), .B1(n6655), .B2(n6107), .C1(n6106), 
        .C2(n6561), .ZN(n6110) );
  MUX2_X1 U7161 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n6110), .S(n6448), 
        .Z(U3462) );
  INV_X1 U7162 ( .A(n6111), .ZN(n6116) );
  NAND3_X1 U7163 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6112), .A3(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7164 ( .A1(n6113), .A2(n6119), .ZN(n6114) );
  OAI211_X1 U7165 ( .C1(n6116), .C2(n4788), .A(n6115), .B(n6114), .ZN(n6117)
         );
  MUX2_X1 U7166 ( .A(n6117), .B(n6756), .S(n6125), .Z(U3460) );
  INV_X1 U7167 ( .A(n6118), .ZN(n6124) );
  INV_X1 U7168 ( .A(n6119), .ZN(n6123) );
  INV_X1 U7169 ( .A(n6120), .ZN(n6122) );
  OAI22_X1 U7170 ( .A1(n6124), .A2(n6123), .B1(n6122), .B2(n6121), .ZN(n6126)
         );
  MUX2_X1 U7171 ( .A(n6126), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6125), 
        .Z(U3456) );
  AND2_X1 U7172 ( .A1(n6295), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  NOR2_X1 U7173 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n6128) );
  OAI21_X1 U7174 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6128), .A(n4598), .ZN(n6127)
         );
  OAI21_X1 U7175 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n4598), .A(n6127), .ZN(
        U2791) );
  OAI21_X1 U7176 ( .B1(BS16_N), .B2(n6128), .A(n6730), .ZN(n6729) );
  OAI21_X1 U7177 ( .B1(n6730), .B2(n6129), .A(n6729), .ZN(U2792) );
  AND2_X1 U7178 ( .A1(n6130), .A2(n6717), .ZN(n6740) );
  OAI21_X1 U7179 ( .B1(n6740), .B2(n6872), .A(n6334), .ZN(U2793) );
  INV_X1 U7180 ( .A(DATAWIDTH_REG_18__SCAN_IN), .ZN(n7006) );
  INV_X1 U7181 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6938) );
  INV_X1 U7182 ( .A(DATAWIDTH_REG_30__SCAN_IN), .ZN(n6990) );
  INV_X1 U7183 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6841) );
  NAND4_X1 U7184 ( .A1(n7006), .A2(n6938), .A3(n6990), .A4(n6841), .ZN(n6131)
         );
  AOI211_X1 U7185 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_8__SCAN_IN), .B(n6131), 
        .ZN(n6140) );
  NOR4_X1 U7186 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n6139) );
  NOR4_X1 U7187 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(DATAWIDTH_REG_27__SCAN_IN), .ZN(n6138)
         );
  NOR4_X1 U7188 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(DATAWIDTH_REG_25__SCAN_IN), .ZN(n6132)
         );
  INV_X1 U7189 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6954) );
  NAND2_X1 U7190 ( .A1(n6132), .A2(n6954), .ZN(n6766) );
  NOR4_X1 U7191 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6135) );
  NOR4_X1 U7192 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_21__SCAN_IN), .A4(
        DATAWIDTH_REG_29__SCAN_IN), .ZN(n6134) );
  NOR4_X1 U7193 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_31__SCAN_IN), .A4(
        DATAWIDTH_REG_2__SCAN_IN), .ZN(n6133) );
  NAND3_X1 U7194 ( .A1(n6135), .A2(n6134), .A3(n6133), .ZN(n6136) );
  NOR2_X1 U7195 ( .A1(n6766), .A2(n6136), .ZN(n6137) );
  NAND4_X1 U7196 ( .A1(n6140), .A2(n6139), .A3(n6138), .A4(n6137), .ZN(n6736)
         );
  NOR2_X1 U7197 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6736), .ZN(n6737) );
  INV_X1 U7198 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6951) );
  OR4_X1 U7199 ( .A1(n6736), .A2(DATAWIDTH_REG_1__SCAN_IN), .A3(
        REIP_REG_0__SCAN_IN), .A4(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6141) );
  OAI221_X1 U7200 ( .B1(n6737), .B2(n6951), .C1(n6737), .C2(n6736), .A(n6141), 
        .ZN(U2794) );
  INV_X1 U7201 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6821) );
  AOI22_X1 U7202 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(n6736), .B1(n6737), 
        .B2(n6821), .ZN(n6142) );
  NAND2_X1 U7203 ( .A1(n6142), .A2(n6141), .ZN(U2795) );
  OAI21_X1 U7204 ( .B1(REIP_REG_12__SCAN_IN), .B2(n6144), .A(n6143), .ZN(n6150) );
  INV_X1 U7205 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6148) );
  INV_X1 U7206 ( .A(n6145), .ZN(n6146) );
  AOI22_X1 U7207 ( .A1(n6146), .A2(n6166), .B1(n6249), .B2(EBX_REG_13__SCAN_IN), .ZN(n6147) );
  OAI211_X1 U7208 ( .C1(n6259), .C2(n6148), .A(n6147), .B(n6190), .ZN(n6149)
         );
  AOI221_X1 U7209 ( .B1(n6152), .B2(n6151), .C1(n6150), .C2(
        REIP_REG_13__SCAN_IN), .A(n6149), .ZN(n6156) );
  INV_X1 U7210 ( .A(n6153), .ZN(n6154) );
  NAND2_X1 U7211 ( .A1(n6154), .A2(n6204), .ZN(n6155) );
  OAI211_X1 U7212 ( .C1(n6258), .C2(n6157), .A(n6156), .B(n6155), .ZN(U2814)
         );
  OAI22_X1 U7213 ( .A1(n6159), .A2(n6259), .B1(n6158), .B2(n6180), .ZN(n6160)
         );
  AOI211_X1 U7214 ( .C1(n6249), .C2(EBX_REG_9__SCAN_IN), .A(n6227), .B(n6160), 
        .ZN(n6170) );
  INV_X1 U7215 ( .A(n6161), .ZN(n6263) );
  AOI22_X1 U7216 ( .A1(n6263), .A2(n6204), .B1(n6175), .B2(n6162), .ZN(n6169)
         );
  AOI21_X1 U7217 ( .B1(n6165), .B2(n6164), .A(n6163), .ZN(n6375) );
  NAND2_X1 U7218 ( .A1(n6375), .A2(n3100), .ZN(n6167) );
  NAND4_X1 U7219 ( .A1(n6170), .A2(n6169), .A3(n6168), .A4(n6167), .ZN(U2818)
         );
  AND2_X1 U7220 ( .A1(n6237), .A2(n6171), .ZN(n6189) );
  AOI21_X1 U7221 ( .B1(REIP_REG_7__SCAN_IN), .B2(n6189), .A(
        REIP_REG_8__SCAN_IN), .ZN(n6181) );
  OAI22_X1 U7222 ( .A1(n6244), .A2(n6172), .B1(n6210), .B2(n7048), .ZN(n6173)
         );
  AOI211_X1 U7223 ( .C1(n6241), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6227), 
        .B(n6173), .ZN(n6179) );
  INV_X1 U7224 ( .A(n6174), .ZN(n6176) );
  AOI22_X1 U7225 ( .A1(n6177), .A2(n6204), .B1(n6176), .B2(n6175), .ZN(n6178)
         );
  OAI211_X1 U7226 ( .C1(n6181), .C2(n6180), .A(n6179), .B(n6178), .ZN(U2819)
         );
  INV_X1 U7227 ( .A(n6182), .ZN(n6183) );
  NAND2_X1 U7228 ( .A1(n6184), .A2(n6183), .ZN(n6185) );
  NAND2_X1 U7229 ( .A1(n6186), .A2(n6185), .ZN(n6219) );
  NAND2_X1 U7230 ( .A1(n6237), .A2(n6187), .ZN(n6224) );
  NOR2_X1 U7231 ( .A1(n7024), .A2(n6224), .ZN(n6206) );
  NAND3_X1 U7232 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6206), .A3(n6395), .ZN(n6202) );
  INV_X1 U7233 ( .A(n6188), .ZN(n6383) );
  AOI22_X1 U7234 ( .A1(n6189), .A2(n6198), .B1(n6166), .B2(n6383), .ZN(n6191)
         );
  OAI211_X1 U7235 ( .C1(n6259), .C2(n6847), .A(n6191), .B(n6190), .ZN(n6196)
         );
  OAI22_X1 U7236 ( .A1(n6194), .A2(n6193), .B1(n6192), .B2(n6258), .ZN(n6195)
         );
  AOI211_X1 U7237 ( .C1(EBX_REG_7__SCAN_IN), .C2(n6249), .A(n6196), .B(n6195), 
        .ZN(n6197) );
  OAI221_X1 U7238 ( .B1(n6198), .B2(n6219), .C1(n6198), .C2(n6202), .A(n6197), 
        .ZN(U2820) );
  OAI22_X1 U7239 ( .A1(n6199), .A2(n6259), .B1(n6244), .B2(n6396), .ZN(n6200)
         );
  AOI211_X1 U7240 ( .C1(n6249), .C2(EBX_REG_6__SCAN_IN), .A(n6227), .B(n6200), 
        .ZN(n6201) );
  OAI211_X1 U7241 ( .C1(n6395), .C2(n6219), .A(n6202), .B(n6201), .ZN(n6203)
         );
  AOI21_X1 U7242 ( .B1(n6204), .B2(n6340), .A(n6203), .ZN(n6205) );
  OAI21_X1 U7243 ( .B1(n6343), .B2(n6258), .A(n6205), .ZN(U2821) );
  NOR2_X1 U7244 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6206), .ZN(n6220) );
  INV_X1 U7245 ( .A(n6207), .ZN(n6405) );
  AOI21_X1 U7246 ( .B1(n6241), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n6227), 
        .ZN(n6208) );
  OAI21_X1 U7247 ( .B1(n6210), .B2(n6209), .A(n6208), .ZN(n6211) );
  AOI21_X1 U7248 ( .B1(n3100), .B2(n6405), .A(n6211), .ZN(n6218) );
  INV_X1 U7249 ( .A(n6212), .ZN(n6213) );
  OAI22_X1 U7250 ( .A1(n6215), .A2(n6214), .B1(n6213), .B2(n6258), .ZN(n6216)
         );
  INV_X1 U7251 ( .A(n6216), .ZN(n6217) );
  OAI211_X1 U7252 ( .C1(n6220), .C2(n6219), .A(n6218), .B(n6217), .ZN(U2822)
         );
  INV_X1 U7253 ( .A(n6221), .ZN(n6222) );
  OAI22_X1 U7254 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6224), .B1(n6223), .B2(n6222), .ZN(n6231) );
  NOR2_X1 U7255 ( .A1(n6244), .A2(n6225), .ZN(n6226) );
  AOI211_X1 U7256 ( .C1(n6241), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6227), 
        .B(n6226), .ZN(n6228) );
  OAI21_X1 U7257 ( .B1(n6229), .B2(n7024), .A(n6228), .ZN(n6230) );
  AOI211_X1 U7258 ( .C1(EBX_REG_4__SCAN_IN), .C2(n6249), .A(n6231), .B(n6230), 
        .ZN(n6234) );
  INV_X1 U7259 ( .A(n6232), .ZN(n6348) );
  NAND2_X1 U7260 ( .A1(n6348), .A2(n6255), .ZN(n6233) );
  OAI211_X1 U7261 ( .C1(n6258), .C2(n6353), .A(n6234), .B(n6233), .ZN(U2823)
         );
  NOR2_X1 U7262 ( .A1(n6236), .A2(n6235), .ZN(n6240) );
  AOI21_X1 U7263 ( .B1(n6237), .B2(REIP_REG_1__SCAN_IN), .A(
        REIP_REG_2__SCAN_IN), .ZN(n6238) );
  AOI21_X1 U7264 ( .B1(n6240), .B2(n6239), .A(n6238), .ZN(n6246) );
  AOI22_X1 U7265 ( .A1(EBX_REG_2__SCAN_IN), .A2(n6249), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n6241), .ZN(n6243) );
  NAND2_X1 U7266 ( .A1(n6248), .A2(n3104), .ZN(n6242) );
  OAI211_X1 U7267 ( .C1(n6244), .C2(n6432), .A(n6243), .B(n6242), .ZN(n6245)
         );
  AOI211_X1 U7268 ( .C1(n6359), .C2(n6255), .A(n6246), .B(n6245), .ZN(n6247)
         );
  OAI21_X1 U7269 ( .B1(n6362), .B2(n6258), .A(n6247), .ZN(U2825) );
  INV_X1 U7270 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n6260) );
  AOI22_X1 U7271 ( .A1(n6249), .A2(EBX_REG_0__SCAN_IN), .B1(n6248), .B2(n3114), 
        .ZN(n6252) );
  NAND2_X1 U7272 ( .A1(n6166), .A2(n6250), .ZN(n6251) );
  OAI211_X1 U7273 ( .C1(n6253), .C2(n6891), .A(n6252), .B(n6251), .ZN(n6254)
         );
  AOI21_X1 U7274 ( .B1(n6256), .B2(n6255), .A(n6254), .ZN(n6257) );
  OAI221_X1 U7275 ( .B1(n6260), .B2(n6259), .C1(n6260), .C2(n6258), .A(n6257), 
        .ZN(U2827) );
  INV_X1 U7276 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6265) );
  AOI22_X1 U7277 ( .A1(n6263), .A2(n6262), .B1(n6261), .B2(n6375), .ZN(n6264)
         );
  OAI21_X1 U7278 ( .B1(n6266), .B2(n6265), .A(n6264), .ZN(U2850) );
  INV_X1 U7279 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n6837) );
  AOI22_X1 U7280 ( .A1(n6272), .A2(EAX_REG_24__SCAN_IN), .B1(n6744), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n6267) );
  OAI21_X1 U7281 ( .B1(n6837), .B2(n6285), .A(n6267), .ZN(U2899) );
  INV_X1 U7282 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n7023) );
  AOI22_X1 U7283 ( .A1(n6272), .A2(EAX_REG_23__SCAN_IN), .B1(n6744), .B2(
        UWORD_REG_7__SCAN_IN), .ZN(n6268) );
  OAI21_X1 U7284 ( .B1(n7023), .B2(n6285), .A(n6268), .ZN(U2900) );
  INV_X1 U7285 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n6809) );
  AOI22_X1 U7286 ( .A1(n6272), .A2(EAX_REG_22__SCAN_IN), .B1(n6744), .B2(
        UWORD_REG_6__SCAN_IN), .ZN(n6269) );
  OAI21_X1 U7287 ( .B1(n6809), .B2(n6285), .A(n6269), .ZN(U2901) );
  AOI22_X1 U7288 ( .A1(n6295), .A2(DATAO_REG_19__SCAN_IN), .B1(n6272), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n6270) );
  OAI21_X1 U7289 ( .B1(n6280), .B2(n4659), .A(n6270), .ZN(U2904) );
  INV_X1 U7290 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n6856) );
  AOI22_X1 U7291 ( .A1(n6272), .A2(EAX_REG_18__SCAN_IN), .B1(n6744), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n6271) );
  OAI21_X1 U7292 ( .B1(n6856), .B2(n6285), .A(n6271), .ZN(U2905) );
  INV_X1 U7293 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n7011) );
  AOI22_X1 U7294 ( .A1(n6295), .A2(DATAO_REG_16__SCAN_IN), .B1(n6272), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6273) );
  OAI21_X1 U7295 ( .B1(n6280), .B2(n7011), .A(n6273), .ZN(U2907) );
  AOI22_X1 U7296 ( .A1(n6744), .A2(LWORD_REG_15__SCAN_IN), .B1(n6295), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6274) );
  OAI21_X1 U7297 ( .B1(n7020), .B2(n6297), .A(n6274), .ZN(U2908) );
  INV_X1 U7298 ( .A(LWORD_REG_14__SCAN_IN), .ZN(n7009) );
  AOI22_X1 U7299 ( .A1(EAX_REG_14__SCAN_IN), .A2(n6288), .B1(n6295), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6275) );
  OAI21_X1 U7300 ( .B1(n6280), .B2(n7009), .A(n6275), .ZN(U2909) );
  INV_X1 U7301 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n6838) );
  AOI22_X1 U7302 ( .A1(EAX_REG_13__SCAN_IN), .A2(n6288), .B1(n6744), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n6276) );
  OAI21_X1 U7303 ( .B1(n6838), .B2(n6285), .A(n6276), .ZN(U2910) );
  INV_X1 U7304 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6278) );
  AOI22_X1 U7305 ( .A1(n6744), .A2(LWORD_REG_12__SCAN_IN), .B1(n6295), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6277) );
  OAI21_X1 U7306 ( .B1(n6278), .B2(n6297), .A(n6277), .ZN(U2911) );
  INV_X1 U7307 ( .A(LWORD_REG_11__SCAN_IN), .ZN(n7016) );
  AOI22_X1 U7308 ( .A1(EAX_REG_11__SCAN_IN), .A2(n6288), .B1(n6295), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6279) );
  OAI21_X1 U7309 ( .B1(n6280), .B2(n7016), .A(n6279), .ZN(U2912) );
  AOI222_X1 U7310 ( .A1(n6295), .A2(DATAO_REG_10__SCAN_IN), .B1(n6288), .B2(
        EAX_REG_10__SCAN_IN), .C1(n6744), .C2(LWORD_REG_10__SCAN_IN), .ZN(
        n6281) );
  INV_X1 U7311 ( .A(n6281), .ZN(U2913) );
  INV_X1 U7312 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6283) );
  AOI22_X1 U7313 ( .A1(n6744), .A2(LWORD_REG_9__SCAN_IN), .B1(n6295), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6282) );
  OAI21_X1 U7314 ( .B1(n6283), .B2(n6297), .A(n6282), .ZN(U2914) );
  INV_X1 U7315 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n6909) );
  AOI22_X1 U7316 ( .A1(EAX_REG_8__SCAN_IN), .A2(n6288), .B1(n6744), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n6284) );
  OAI21_X1 U7317 ( .B1(n6909), .B2(n6285), .A(n6284), .ZN(U2915) );
  AOI22_X1 U7318 ( .A1(n6744), .A2(LWORD_REG_7__SCAN_IN), .B1(n6295), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6286) );
  OAI21_X1 U7319 ( .B1(n4640), .B2(n6297), .A(n6286), .ZN(U2916) );
  AOI222_X1 U7320 ( .A1(n6295), .A2(DATAO_REG_6__SCAN_IN), .B1(n6288), .B2(
        EAX_REG_6__SCAN_IN), .C1(n6744), .C2(LWORD_REG_6__SCAN_IN), .ZN(n6287)
         );
  INV_X1 U7321 ( .A(n6287), .ZN(U2917) );
  AOI222_X1 U7322 ( .A1(n6295), .A2(DATAO_REG_5__SCAN_IN), .B1(n6288), .B2(
        EAX_REG_5__SCAN_IN), .C1(n6744), .C2(LWORD_REG_5__SCAN_IN), .ZN(n6289)
         );
  INV_X1 U7323 ( .A(n6289), .ZN(U2918) );
  AOI22_X1 U7324 ( .A1(n6744), .A2(LWORD_REG_4__SCAN_IN), .B1(n6295), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6290) );
  OAI21_X1 U7325 ( .B1(n7003), .B2(n6297), .A(n6290), .ZN(U2919) );
  AOI22_X1 U7326 ( .A1(n6744), .A2(LWORD_REG_3__SCAN_IN), .B1(n6295), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6291) );
  OAI21_X1 U7327 ( .B1(n6292), .B2(n6297), .A(n6291), .ZN(U2920) );
  AOI22_X1 U7328 ( .A1(n6744), .A2(LWORD_REG_2__SCAN_IN), .B1(n6295), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6293) );
  OAI21_X1 U7329 ( .B1(n4646), .B2(n6297), .A(n6293), .ZN(U2921) );
  AOI22_X1 U7330 ( .A1(n6744), .A2(LWORD_REG_1__SCAN_IN), .B1(n6295), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6294) );
  OAI21_X1 U7331 ( .B1(n6855), .B2(n6297), .A(n6294), .ZN(U2922) );
  AOI22_X1 U7332 ( .A1(n6744), .A2(LWORD_REG_0__SCAN_IN), .B1(n6295), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6296) );
  OAI21_X1 U7333 ( .B1(n4689), .B2(n6297), .A(n6296), .ZN(U2923) );
  AOI22_X1 U7334 ( .A1(n6304), .A2(DATAI_0_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n6323), .ZN(n6298) );
  OAI21_X1 U7335 ( .B1(n7011), .B2(n6325), .A(n6298), .ZN(U2924) );
  AOI22_X1 U7336 ( .A1(EAX_REG_24__SCAN_IN), .A2(n6323), .B1(n6319), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n6299) );
  NAND2_X1 U7337 ( .A1(n6304), .A2(DATAI_8_), .ZN(n6311) );
  NAND2_X1 U7338 ( .A1(n6299), .A2(n6311), .ZN(U2932) );
  AOI22_X1 U7339 ( .A1(EAX_REG_26__SCAN_IN), .A2(n6323), .B1(n6319), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U7340 ( .A1(n6304), .A2(DATAI_10_), .ZN(n6313) );
  NAND2_X1 U7341 ( .A1(n6300), .A2(n6313), .ZN(U2934) );
  INV_X1 U7342 ( .A(DATAI_11_), .ZN(n6301) );
  NOR2_X1 U7343 ( .A1(n6308), .A2(n6301), .ZN(n6315) );
  AOI21_X1 U7344 ( .B1(n6319), .B2(UWORD_REG_11__SCAN_IN), .A(n6315), .ZN(
        n6302) );
  OAI21_X1 U7345 ( .B1(n4003), .B2(n6310), .A(n6302), .ZN(U2935) );
  AOI22_X1 U7346 ( .A1(EAX_REG_28__SCAN_IN), .A2(n6323), .B1(n6319), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U7347 ( .A1(n6304), .A2(DATAI_12_), .ZN(n6317) );
  NAND2_X1 U7348 ( .A1(n6303), .A2(n6317), .ZN(U2936) );
  NAND2_X1 U7349 ( .A1(n6304), .A2(DATAI_13_), .ZN(n6320) );
  INV_X1 U7350 ( .A(n6320), .ZN(n6305) );
  AOI21_X1 U7351 ( .B1(n6319), .B2(UWORD_REG_13__SCAN_IN), .A(n6305), .ZN(
        n6306) );
  OAI21_X1 U7352 ( .B1(n4048), .B2(n6310), .A(n6306), .ZN(U2937) );
  INV_X1 U7353 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6903) );
  INV_X1 U7354 ( .A(DATAI_14_), .ZN(n6307) );
  NOR2_X1 U7355 ( .A1(n6308), .A2(n6307), .ZN(n6322) );
  AOI21_X1 U7356 ( .B1(n6319), .B2(UWORD_REG_14__SCAN_IN), .A(n6322), .ZN(
        n6309) );
  OAI21_X1 U7357 ( .B1(n6903), .B2(n6310), .A(n6309), .ZN(U2938) );
  AOI22_X1 U7358 ( .A1(EAX_REG_8__SCAN_IN), .A2(n6323), .B1(n6319), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n6312) );
  NAND2_X1 U7359 ( .A1(n6312), .A2(n6311), .ZN(U2947) );
  AOI22_X1 U7360 ( .A1(EAX_REG_10__SCAN_IN), .A2(n6323), .B1(
        LWORD_REG_10__SCAN_IN), .B2(n6319), .ZN(n6314) );
  NAND2_X1 U7361 ( .A1(n6314), .A2(n6313), .ZN(U2949) );
  AOI21_X1 U7362 ( .B1(n6323), .B2(EAX_REG_11__SCAN_IN), .A(n6315), .ZN(n6316)
         );
  OAI21_X1 U7363 ( .B1(n7016), .B2(n6325), .A(n6316), .ZN(U2950) );
  AOI22_X1 U7364 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6323), .B1(n6319), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n6318) );
  NAND2_X1 U7365 ( .A1(n6318), .A2(n6317), .ZN(U2951) );
  AOI22_X1 U7366 ( .A1(EAX_REG_13__SCAN_IN), .A2(n6323), .B1(n6319), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n6321) );
  NAND2_X1 U7367 ( .A1(n6321), .A2(n6320), .ZN(U2952) );
  AOI21_X1 U7368 ( .B1(n6323), .B2(EAX_REG_14__SCAN_IN), .A(n6322), .ZN(n6324)
         );
  OAI21_X1 U7369 ( .B1(n7009), .B2(n6325), .A(n6324), .ZN(U2953) );
  INV_X1 U7370 ( .A(n6326), .ZN(n6327) );
  AOI21_X1 U7371 ( .B1(n6354), .B2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6327), 
        .ZN(n6333) );
  INV_X1 U7372 ( .A(n6328), .ZN(n6331) );
  AOI22_X1 U7373 ( .A1(n6331), .A2(n6349), .B1(n6330), .B2(n6329), .ZN(n6332)
         );
  OAI211_X1 U7374 ( .C1(n6335), .C2(n6334), .A(n6333), .B(n6332), .ZN(U2975)
         );
  AOI22_X1 U7375 ( .A1(n6354), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .B1(n6433), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n6342) );
  OAI21_X1 U7376 ( .B1(n6338), .B2(n6337), .A(n6336), .ZN(n6339) );
  INV_X1 U7377 ( .A(n6339), .ZN(n6399) );
  AOI22_X1 U7378 ( .A1(n6399), .A2(n6358), .B1(n6349), .B2(n6340), .ZN(n6341)
         );
  OAI211_X1 U7379 ( .C1(n6363), .C2(n6343), .A(n6342), .B(n6341), .ZN(U2980)
         );
  AOI22_X1 U7380 ( .A1(n6354), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n6433), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n6352) );
  OR2_X1 U7381 ( .A1(n6345), .A2(n6344), .ZN(n6346) );
  NAND2_X1 U7382 ( .A1(n6347), .A2(n6346), .ZN(n6413) );
  INV_X1 U7383 ( .A(n6413), .ZN(n6350) );
  AOI22_X1 U7384 ( .A1(n6350), .A2(n6358), .B1(n6349), .B2(n6348), .ZN(n6351)
         );
  OAI211_X1 U7385 ( .C1(n6363), .C2(n6353), .A(n6352), .B(n6351), .ZN(U2982)
         );
  AOI22_X1 U7386 ( .A1(n6354), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n6433), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6361) );
  XNOR2_X1 U7387 ( .A(n6355), .B(n6442), .ZN(n6357) );
  XNOR2_X1 U7388 ( .A(n6357), .B(n6356), .ZN(n6441) );
  AOI22_X1 U7389 ( .A1(n6359), .A2(n6349), .B1(n6358), .B2(n6441), .ZN(n6360)
         );
  OAI211_X1 U7390 ( .C1(n6363), .C2(n6362), .A(n6361), .B(n6360), .ZN(U2984)
         );
  NAND2_X1 U7391 ( .A1(n6367), .A2(n6386), .ZN(n6380) );
  AOI22_X1 U7392 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n5862), .B1(
        INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6364), .ZN(n6372) );
  AOI21_X1 U7393 ( .B1(n6366), .B2(n6435), .A(n6365), .ZN(n6371) );
  OAI21_X1 U7394 ( .B1(n6368), .B2(n6367), .A(n6390), .ZN(n6376) );
  AOI22_X1 U7395 ( .A1(n6369), .A2(n6440), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6376), .ZN(n6370) );
  OAI211_X1 U7396 ( .C1(n6380), .C2(n6372), .A(n6371), .B(n6370), .ZN(U3008)
         );
  INV_X1 U7397 ( .A(n6373), .ZN(n6374) );
  AOI21_X1 U7398 ( .B1(n6375), .B2(n6435), .A(n6374), .ZN(n6379) );
  AOI22_X1 U7399 ( .A1(n6377), .A2(n6440), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6376), .ZN(n6378) );
  OAI211_X1 U7400 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6380), .A(n6379), 
        .B(n6378), .ZN(U3009) );
  INV_X1 U7401 ( .A(n6381), .ZN(n6382) );
  AOI21_X1 U7402 ( .B1(n6383), .B2(n6435), .A(n6382), .ZN(n6388) );
  INV_X1 U7403 ( .A(n6384), .ZN(n6385) );
  AOI22_X1 U7404 ( .A1(n6386), .A2(n6389), .B1(n6385), .B2(n6440), .ZN(n6387)
         );
  OAI211_X1 U7405 ( .C1(n6390), .C2(n6389), .A(n6388), .B(n6387), .ZN(U3011)
         );
  OAI22_X1 U7406 ( .A1(n6392), .A2(n6437), .B1(n6436), .B2(n6391), .ZN(n6439)
         );
  AOI21_X1 U7407 ( .B1(n6394), .B2(n6393), .A(n6439), .ZN(n6410) );
  OAI22_X1 U7408 ( .A1(n6397), .A2(n6396), .B1(n6395), .B2(n6423), .ZN(n6398)
         );
  AOI21_X1 U7409 ( .B1(n6399), .B2(n6440), .A(n6398), .ZN(n6400) );
  OAI221_X1 U7410 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n6402), .C1(n6401), .C2(n6410), .A(n6400), .ZN(U3012) );
  NOR2_X1 U7411 ( .A1(n6430), .A2(n6420), .ZN(n6411) );
  AOI21_X1 U7412 ( .B1(n6411), .B2(n6403), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6409) );
  INV_X1 U7413 ( .A(n6404), .ZN(n6406) );
  AOI22_X1 U7414 ( .A1(n6406), .A2(n6440), .B1(n6435), .B2(n6405), .ZN(n6408)
         );
  OAI211_X1 U7415 ( .C1(n6410), .C2(n6409), .A(n6408), .B(n6407), .ZN(U3013)
         );
  AOI21_X1 U7416 ( .B1(n6436), .B2(n6438), .A(n6439), .ZN(n6429) );
  AOI211_X1 U7417 ( .C1(n6430), .C2(n6420), .A(n6411), .B(n6431), .ZN(n6418)
         );
  NOR2_X1 U7418 ( .A1(n6413), .A2(n6412), .ZN(n6417) );
  NAND2_X1 U7419 ( .A1(n6435), .A2(n6414), .ZN(n6415) );
  OAI21_X1 U7420 ( .B1(n7024), .B2(n6423), .A(n6415), .ZN(n6416) );
  NOR3_X1 U7421 ( .A1(n6418), .A2(n6417), .A3(n6416), .ZN(n6419) );
  OAI21_X1 U7422 ( .B1(n6429), .B2(n6420), .A(n6419), .ZN(U3014) );
  NAND3_X1 U7423 ( .A1(n6421), .A2(n6440), .A3(n4865), .ZN(n6427) );
  NOR2_X1 U7424 ( .A1(n6423), .A2(n6422), .ZN(n6424) );
  AOI21_X1 U7425 ( .B1(n6435), .B2(n6425), .A(n6424), .ZN(n6426) );
  AND2_X1 U7426 ( .A1(n6427), .A2(n6426), .ZN(n6428) );
  OAI221_X1 U7427 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n6431), .C1(n6430), .C2(n6429), .A(n6428), .ZN(U3015) );
  INV_X1 U7428 ( .A(n6432), .ZN(n6434) );
  AOI22_X1 U7429 ( .A1(n6435), .A2(n6434), .B1(n6433), .B2(REIP_REG_2__SCAN_IN), .ZN(n6447) );
  OAI221_X1 U7430 ( .B1(n6438), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .C1(n6438), .C2(n6437), .A(n6436), .ZN(n6446) );
  AOI22_X1 U7431 ( .A1(n6441), .A2(n6440), .B1(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6439), .ZN(n6445) );
  NAND3_X1 U7432 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6443), .A3(n6442), 
        .ZN(n6444) );
  NAND4_X1 U7433 ( .A1(n6447), .A2(n6446), .A3(n6445), .A4(n6444), .ZN(U3016)
         );
  NOR2_X1 U7434 ( .A1(n7040), .A2(n6448), .ZN(U3019) );
  OAI22_X1 U7435 ( .A1(n6517), .A2(n6591), .B1(n6590), .B2(n6483), .ZN(n6450)
         );
  INV_X1 U7436 ( .A(n6450), .ZN(n6464) );
  INV_X1 U7437 ( .A(n6595), .ZN(n6451) );
  NAND2_X1 U7438 ( .A1(n6452), .A2(n6451), .ZN(n6453) );
  OAI21_X1 U7439 ( .B1(n6593), .B2(n6453), .A(n6594), .ZN(n6462) );
  OR2_X1 U7440 ( .A1(n6454), .A2(n6521), .ZN(n6455) );
  INV_X1 U7441 ( .A(n6461), .ZN(n6459) );
  INV_X1 U7442 ( .A(n6456), .ZN(n6458) );
  INV_X1 U7443 ( .A(n6523), .ZN(n6457) );
  AOI21_X1 U7444 ( .B1(n6458), .B2(n6655), .A(n6457), .ZN(n6599) );
  OAI211_X1 U7445 ( .C1(n6462), .C2(n6459), .A(n6599), .B(n6781), .ZN(n6486)
         );
  OAI22_X1 U7446 ( .A1(n6462), .A2(n6461), .B1(n6603), .B2(n6460), .ZN(n6485)
         );
  AOI22_X1 U7447 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6486), .B1(n6654), 
        .B2(n6485), .ZN(n6463) );
  OAI211_X1 U7448 ( .C1(n6669), .C2(n6489), .A(n6464), .B(n6463), .ZN(U3044)
         );
  OAI22_X1 U7449 ( .A1(n6517), .A2(n6609), .B1(n6608), .B2(n6483), .ZN(n6465)
         );
  INV_X1 U7450 ( .A(n6465), .ZN(n6467) );
  AOI22_X1 U7451 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6486), .B1(n6671), 
        .B2(n6485), .ZN(n6466) );
  OAI211_X1 U7452 ( .C1(n6489), .C2(n6675), .A(n6467), .B(n6466), .ZN(U3045)
         );
  OAI22_X1 U7453 ( .A1(n6489), .A2(n6681), .B1(n6613), .B2(n6483), .ZN(n6468)
         );
  INV_X1 U7454 ( .A(n6468), .ZN(n6470) );
  AOI22_X1 U7455 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6486), .B1(n6677), 
        .B2(n6485), .ZN(n6469) );
  OAI211_X1 U7456 ( .C1(n6617), .C2(n6517), .A(n6470), .B(n6469), .ZN(U3046)
         );
  OAI22_X1 U7457 ( .A1(n6517), .A2(n6619), .B1(n6618), .B2(n6483), .ZN(n6471)
         );
  INV_X1 U7458 ( .A(n6471), .ZN(n6473) );
  AOI22_X1 U7459 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6486), .B1(n6683), 
        .B2(n6485), .ZN(n6472) );
  OAI211_X1 U7460 ( .C1(n6489), .C2(n6687), .A(n6473), .B(n6472), .ZN(U3047)
         );
  OAI22_X1 U7461 ( .A1(n6517), .A2(n6624), .B1(n6623), .B2(n6483), .ZN(n6474)
         );
  INV_X1 U7462 ( .A(n6474), .ZN(n6476) );
  AOI22_X1 U7463 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6486), .B1(n6689), 
        .B2(n6485), .ZN(n6475) );
  OAI211_X1 U7464 ( .C1(n6489), .C2(n6693), .A(n6476), .B(n6475), .ZN(U3048)
         );
  OAI22_X1 U7465 ( .A1(n6489), .A2(n6699), .B1(n6628), .B2(n6483), .ZN(n6477)
         );
  INV_X1 U7466 ( .A(n6477), .ZN(n6479) );
  AOI22_X1 U7467 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6486), .B1(n6695), 
        .B2(n6485), .ZN(n6478) );
  OAI211_X1 U7468 ( .C1(n6632), .C2(n6517), .A(n6479), .B(n6478), .ZN(U3049)
         );
  OAI22_X1 U7469 ( .A1(n6517), .A2(n7073), .B1(n7072), .B2(n6483), .ZN(n6480)
         );
  INV_X1 U7470 ( .A(n6480), .ZN(n6482) );
  AOI22_X1 U7471 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6486), .B1(n6701), 
        .B2(n6485), .ZN(n6481) );
  OAI211_X1 U7472 ( .C1(n6489), .C2(n6705), .A(n6482), .B(n6481), .ZN(U3050)
         );
  OAI22_X1 U7473 ( .A1(n6517), .A2(n6638), .B1(n6637), .B2(n6483), .ZN(n6484)
         );
  INV_X1 U7474 ( .A(n6484), .ZN(n6488) );
  AOI22_X1 U7475 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6486), .B1(n6708), 
        .B2(n6485), .ZN(n6487) );
  OAI211_X1 U7476 ( .C1(n6489), .C2(n6716), .A(n6488), .B(n6487), .ZN(U3051)
         );
  OAI33_X1 U7477 ( .A1(n4743), .A2(n6657), .A3(n6655), .B1(n6563), .B2(n6490), 
        .B3(n6645), .ZN(n6513) );
  INV_X1 U7478 ( .A(n6590), .ZN(n6653) );
  NAND2_X1 U7479 ( .A1(n6491), .A2(n6651), .ZN(n6494) );
  INV_X1 U7480 ( .A(n6494), .ZN(n6512) );
  AOI22_X1 U7481 ( .A1(n6513), .A2(n6654), .B1(n6653), .B2(n6512), .ZN(n6499)
         );
  NOR2_X1 U7482 ( .A1(n7076), .A2(n6655), .ZN(n6492) );
  AOI21_X1 U7483 ( .B1(n6492), .B2(n6517), .A(n6659), .ZN(n6497) );
  AOI211_X1 U7484 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6494), .A(n6662), .B(
        n6493), .ZN(n6495) );
  AOI22_X1 U7485 ( .A1(n6514), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n6666), 
        .B2(n7076), .ZN(n6498) );
  OAI211_X1 U7486 ( .C1(n6669), .C2(n6517), .A(n6499), .B(n6498), .ZN(U3052)
         );
  INV_X1 U7487 ( .A(n6608), .ZN(n6670) );
  AOI22_X1 U7488 ( .A1(n6513), .A2(n6671), .B1(n6670), .B2(n6512), .ZN(n6501)
         );
  AOI22_X1 U7489 ( .A1(n6514), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n6672), 
        .B2(n7076), .ZN(n6500) );
  OAI211_X1 U7490 ( .C1(n6675), .C2(n6517), .A(n6501), .B(n6500), .ZN(U3053)
         );
  INV_X1 U7491 ( .A(n6613), .ZN(n6676) );
  AOI22_X1 U7492 ( .A1(n6513), .A2(n6677), .B1(n6676), .B2(n6512), .ZN(n6503)
         );
  AOI22_X1 U7493 ( .A1(n6514), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n6678), 
        .B2(n7076), .ZN(n6502) );
  OAI211_X1 U7494 ( .C1(n6681), .C2(n6517), .A(n6503), .B(n6502), .ZN(U3054)
         );
  INV_X1 U7495 ( .A(n6618), .ZN(n6682) );
  AOI22_X1 U7496 ( .A1(n3143), .A2(n6683), .B1(n6682), .B2(n6512), .ZN(n6505)
         );
  AOI22_X1 U7497 ( .A1(n6514), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n6684), 
        .B2(n7076), .ZN(n6504) );
  OAI211_X1 U7498 ( .C1(n6687), .C2(n6517), .A(n6505), .B(n6504), .ZN(U3055)
         );
  INV_X1 U7499 ( .A(n6623), .ZN(n6688) );
  AOI22_X1 U7500 ( .A1(n6513), .A2(n6689), .B1(n6688), .B2(n6512), .ZN(n6507)
         );
  AOI22_X1 U7501 ( .A1(n6514), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n6690), 
        .B2(n7076), .ZN(n6506) );
  OAI211_X1 U7502 ( .C1(n6693), .C2(n6517), .A(n6507), .B(n6506), .ZN(U3056)
         );
  INV_X1 U7503 ( .A(n6628), .ZN(n6694) );
  AOI22_X1 U7504 ( .A1(n3143), .A2(n6695), .B1(n6694), .B2(n6512), .ZN(n6509)
         );
  AOI22_X1 U7505 ( .A1(n6514), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n6696), 
        .B2(n7076), .ZN(n6508) );
  OAI211_X1 U7506 ( .C1(n6699), .C2(n6517), .A(n6509), .B(n6508), .ZN(U3057)
         );
  INV_X1 U7507 ( .A(n7072), .ZN(n6700) );
  AOI22_X1 U7508 ( .A1(n3143), .A2(n6701), .B1(n6700), .B2(n6512), .ZN(n6511)
         );
  AOI22_X1 U7509 ( .A1(n6514), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n6702), 
        .B2(n7076), .ZN(n6510) );
  OAI211_X1 U7510 ( .C1(n6705), .C2(n6517), .A(n6511), .B(n6510), .ZN(U3058)
         );
  INV_X1 U7511 ( .A(n6637), .ZN(n6707) );
  AOI22_X1 U7512 ( .A1(n3143), .A2(n6708), .B1(n6707), .B2(n6512), .ZN(n6516)
         );
  AOI22_X1 U7513 ( .A1(n6514), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n6711), 
        .B2(n7076), .ZN(n6515) );
  OAI211_X1 U7514 ( .C1(n6716), .C2(n6517), .A(n6516), .B(n6515), .ZN(U3059)
         );
  OAI22_X1 U7515 ( .A1(n6551), .A2(n6669), .B1(n6550), .B2(n6590), .ZN(n6520)
         );
  INV_X1 U7516 ( .A(n6520), .ZN(n6531) );
  OAI21_X1 U7517 ( .B1(n6522), .B2(n6521), .A(n6550), .ZN(n6525) );
  OR3_X1 U7518 ( .A1(n6529), .A2(n6655), .A3(n6525), .ZN(n6524) );
  OAI211_X1 U7519 ( .C1(n6526), .C2(n6594), .A(n6524), .B(n6523), .ZN(n6554)
         );
  NAND2_X1 U7520 ( .A1(n6525), .A2(n6594), .ZN(n6528) );
  INV_X1 U7521 ( .A(n6526), .ZN(n6527) );
  OAI22_X1 U7522 ( .A1(n6529), .A2(n6528), .B1(n6527), .B2(n6603), .ZN(n6553)
         );
  AOI22_X1 U7523 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6554), .B1(n6654), 
        .B2(n6553), .ZN(n6530) );
  OAI211_X1 U7524 ( .C1(n6591), .C2(n6588), .A(n6531), .B(n6530), .ZN(U3076)
         );
  OAI22_X1 U7525 ( .A1(n6551), .A2(n6675), .B1(n6550), .B2(n6608), .ZN(n6532)
         );
  INV_X1 U7526 ( .A(n6532), .ZN(n6534) );
  AOI22_X1 U7527 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6554), .B1(n6671), 
        .B2(n6553), .ZN(n6533) );
  OAI211_X1 U7528 ( .C1(n6609), .C2(n6588), .A(n6534), .B(n6533), .ZN(U3077)
         );
  OAI22_X1 U7529 ( .A1(n6551), .A2(n6681), .B1(n6550), .B2(n6613), .ZN(n6535)
         );
  INV_X1 U7530 ( .A(n6535), .ZN(n6537) );
  AOI22_X1 U7531 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6554), .B1(n6677), 
        .B2(n6553), .ZN(n6536) );
  OAI211_X1 U7532 ( .C1(n6617), .C2(n6588), .A(n6537), .B(n6536), .ZN(U3078)
         );
  OAI22_X1 U7533 ( .A1(n6551), .A2(n6687), .B1(n6550), .B2(n6618), .ZN(n6538)
         );
  INV_X1 U7534 ( .A(n6538), .ZN(n6540) );
  AOI22_X1 U7535 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6554), .B1(n6683), 
        .B2(n6553), .ZN(n6539) );
  OAI211_X1 U7536 ( .C1(n6619), .C2(n6588), .A(n6540), .B(n6539), .ZN(U3079)
         );
  OAI22_X1 U7537 ( .A1(n6551), .A2(n6693), .B1(n6550), .B2(n6623), .ZN(n6541)
         );
  INV_X1 U7538 ( .A(n6541), .ZN(n6543) );
  AOI22_X1 U7539 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6554), .B1(n6689), 
        .B2(n6553), .ZN(n6542) );
  OAI211_X1 U7540 ( .C1(n6624), .C2(n6588), .A(n6543), .B(n6542), .ZN(U3080)
         );
  OAI22_X1 U7541 ( .A1(n6551), .A2(n6699), .B1(n6550), .B2(n6628), .ZN(n6544)
         );
  INV_X1 U7542 ( .A(n6544), .ZN(n6546) );
  AOI22_X1 U7543 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6554), .B1(n6695), 
        .B2(n6553), .ZN(n6545) );
  OAI211_X1 U7544 ( .C1(n6632), .C2(n6588), .A(n6546), .B(n6545), .ZN(U3081)
         );
  OAI22_X1 U7545 ( .A1(n6551), .A2(n6705), .B1(n6550), .B2(n7072), .ZN(n6547)
         );
  INV_X1 U7546 ( .A(n6547), .ZN(n6549) );
  AOI22_X1 U7547 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6554), .B1(n6701), 
        .B2(n6553), .ZN(n6548) );
  OAI211_X1 U7548 ( .C1(n7073), .C2(n6588), .A(n6549), .B(n6548), .ZN(U3082)
         );
  OAI22_X1 U7549 ( .A1(n6551), .A2(n6716), .B1(n6550), .B2(n6637), .ZN(n6552)
         );
  INV_X1 U7550 ( .A(n6552), .ZN(n6556) );
  AOI22_X1 U7551 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6554), .B1(n6708), 
        .B2(n6553), .ZN(n6555) );
  OAI211_X1 U7552 ( .C1(n6638), .C2(n6588), .A(n6556), .B(n6555), .ZN(U3083)
         );
  INV_X1 U7553 ( .A(n6557), .ZN(n6558) );
  OAI22_X1 U7554 ( .A1(n6650), .A2(n6560), .B1(n6649), .B2(n6558), .ZN(n6583)
         );
  OR2_X1 U7555 ( .A1(n6559), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6564)
         );
  INV_X1 U7556 ( .A(n6564), .ZN(n6582) );
  AOI22_X1 U7557 ( .A1(n6583), .A2(n6654), .B1(n6653), .B2(n6582), .ZN(n6569)
         );
  OAI22_X1 U7558 ( .A1(n6588), .A2(n6659), .B1(n6561), .B2(n6560), .ZN(n6566)
         );
  OAI21_X1 U7559 ( .B1(n6563), .B2(n6603), .A(n6562), .ZN(n6661) );
  AOI211_X1 U7560 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6564), .A(n6647), .B(
        n6661), .ZN(n6565) );
  AOI22_X1 U7561 ( .A1(n6585), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6666), 
        .B2(n6584), .ZN(n6568) );
  OAI211_X1 U7562 ( .C1(n6669), .C2(n6588), .A(n6569), .B(n6568), .ZN(U3084)
         );
  AOI22_X1 U7563 ( .A1(n6583), .A2(n6671), .B1(n6670), .B2(n6582), .ZN(n6571)
         );
  AOI22_X1 U7564 ( .A1(n6585), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6672), 
        .B2(n6584), .ZN(n6570) );
  OAI211_X1 U7565 ( .C1(n6675), .C2(n6588), .A(n6571), .B(n6570), .ZN(U3085)
         );
  AOI22_X1 U7566 ( .A1(n6583), .A2(n6677), .B1(n6676), .B2(n6582), .ZN(n6573)
         );
  AOI22_X1 U7567 ( .A1(n6585), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6678), 
        .B2(n6584), .ZN(n6572) );
  OAI211_X1 U7568 ( .C1(n6681), .C2(n6588), .A(n6573), .B(n6572), .ZN(U3086)
         );
  AOI22_X1 U7569 ( .A1(n6583), .A2(n6683), .B1(n6682), .B2(n6582), .ZN(n6575)
         );
  AOI22_X1 U7570 ( .A1(n6585), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6684), 
        .B2(n6584), .ZN(n6574) );
  OAI211_X1 U7571 ( .C1(n6687), .C2(n6588), .A(n6575), .B(n6574), .ZN(U3087)
         );
  AOI22_X1 U7572 ( .A1(n6583), .A2(n6689), .B1(n6688), .B2(n6582), .ZN(n6577)
         );
  AOI22_X1 U7573 ( .A1(n6585), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6690), 
        .B2(n6584), .ZN(n6576) );
  OAI211_X1 U7574 ( .C1(n6693), .C2(n6588), .A(n6577), .B(n6576), .ZN(U3088)
         );
  AOI22_X1 U7575 ( .A1(n6583), .A2(n6695), .B1(n6694), .B2(n6582), .ZN(n6579)
         );
  AOI22_X1 U7576 ( .A1(n6585), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6696), 
        .B2(n6584), .ZN(n6578) );
  OAI211_X1 U7577 ( .C1(n6699), .C2(n6588), .A(n6579), .B(n6578), .ZN(U3089)
         );
  AOI22_X1 U7578 ( .A1(n6583), .A2(n6701), .B1(n6700), .B2(n6582), .ZN(n6581)
         );
  AOI22_X1 U7579 ( .A1(n6585), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6702), 
        .B2(n6584), .ZN(n6580) );
  OAI211_X1 U7580 ( .C1(n6705), .C2(n6588), .A(n6581), .B(n6580), .ZN(U3090)
         );
  AOI22_X1 U7581 ( .A1(n6583), .A2(n6708), .B1(n6707), .B2(n6582), .ZN(n6587)
         );
  AOI22_X1 U7582 ( .A1(n6585), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6711), 
        .B2(n6584), .ZN(n6586) );
  OAI211_X1 U7583 ( .C1(n6716), .C2(n6588), .A(n6587), .B(n6586), .ZN(U3091)
         );
  AND2_X1 U7584 ( .A1(n6601), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6597)
         );
  INV_X1 U7585 ( .A(n6597), .ZN(n6636) );
  OAI22_X1 U7586 ( .A1(n6715), .A2(n6591), .B1(n6590), .B2(n6636), .ZN(n6592)
         );
  INV_X1 U7587 ( .A(n6592), .ZN(n6607) );
  INV_X1 U7588 ( .A(n6593), .ZN(n6596) );
  OAI21_X1 U7589 ( .B1(n6596), .B2(n6595), .A(n6594), .ZN(n6605) );
  AOI21_X1 U7590 ( .B1(n6598), .B2(n3114), .A(n6597), .ZN(n6604) );
  INV_X1 U7591 ( .A(n6604), .ZN(n6600) );
  OAI211_X1 U7592 ( .C1(n6605), .C2(n6600), .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n6599), .ZN(n6641) );
  INV_X1 U7593 ( .A(n6601), .ZN(n6602) );
  OAI22_X1 U7594 ( .A1(n6605), .A2(n6604), .B1(n6603), .B2(n6602), .ZN(n6640)
         );
  AOI22_X1 U7595 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6641), .B1(n6654), 
        .B2(n6640), .ZN(n6606) );
  OAI211_X1 U7596 ( .C1(n6669), .C2(n6644), .A(n6607), .B(n6606), .ZN(U3108)
         );
  OAI22_X1 U7597 ( .A1(n6715), .A2(n6609), .B1(n6608), .B2(n6636), .ZN(n6610)
         );
  INV_X1 U7598 ( .A(n6610), .ZN(n6612) );
  AOI22_X1 U7599 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6641), .B1(n6671), 
        .B2(n6640), .ZN(n6611) );
  OAI211_X1 U7600 ( .C1(n6675), .C2(n6644), .A(n6612), .B(n6611), .ZN(U3109)
         );
  OAI22_X1 U7601 ( .A1(n6644), .A2(n6681), .B1(n6613), .B2(n6636), .ZN(n6614)
         );
  INV_X1 U7602 ( .A(n6614), .ZN(n6616) );
  AOI22_X1 U7603 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6641), .B1(n6677), 
        .B2(n6640), .ZN(n6615) );
  OAI211_X1 U7604 ( .C1(n6617), .C2(n6715), .A(n6616), .B(n6615), .ZN(U3110)
         );
  OAI22_X1 U7605 ( .A1(n6715), .A2(n6619), .B1(n6618), .B2(n6636), .ZN(n6620)
         );
  INV_X1 U7606 ( .A(n6620), .ZN(n6622) );
  AOI22_X1 U7607 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6641), .B1(n6683), 
        .B2(n6640), .ZN(n6621) );
  OAI211_X1 U7608 ( .C1(n6687), .C2(n6644), .A(n6622), .B(n6621), .ZN(U3111)
         );
  OAI22_X1 U7609 ( .A1(n6715), .A2(n6624), .B1(n6623), .B2(n6636), .ZN(n6625)
         );
  INV_X1 U7610 ( .A(n6625), .ZN(n6627) );
  AOI22_X1 U7611 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6641), .B1(n6689), 
        .B2(n6640), .ZN(n6626) );
  OAI211_X1 U7612 ( .C1(n6693), .C2(n6644), .A(n6627), .B(n6626), .ZN(U3112)
         );
  OAI22_X1 U7613 ( .A1(n6644), .A2(n6699), .B1(n6628), .B2(n6636), .ZN(n6629)
         );
  INV_X1 U7614 ( .A(n6629), .ZN(n6631) );
  AOI22_X1 U7615 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6641), .B1(n6695), 
        .B2(n6640), .ZN(n6630) );
  OAI211_X1 U7616 ( .C1(n6632), .C2(n6715), .A(n6631), .B(n6630), .ZN(U3113)
         );
  OAI22_X1 U7617 ( .A1(n6644), .A2(n6705), .B1(n7072), .B2(n6636), .ZN(n6633)
         );
  INV_X1 U7618 ( .A(n6633), .ZN(n6635) );
  AOI22_X1 U7619 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6641), .B1(n6701), 
        .B2(n6640), .ZN(n6634) );
  OAI211_X1 U7620 ( .C1(n7073), .C2(n6715), .A(n6635), .B(n6634), .ZN(U3114)
         );
  OAI22_X1 U7621 ( .A1(n6715), .A2(n6638), .B1(n6637), .B2(n6636), .ZN(n6639)
         );
  INV_X1 U7622 ( .A(n6639), .ZN(n6643) );
  AOI22_X1 U7623 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6641), .B1(n6708), 
        .B2(n6640), .ZN(n6642) );
  OAI211_X1 U7624 ( .C1(n6716), .C2(n6644), .A(n6643), .B(n6642), .ZN(U3115)
         );
  INV_X1 U7625 ( .A(n6645), .ZN(n6646) );
  NAND2_X1 U7626 ( .A1(n6647), .A2(n6646), .ZN(n6648) );
  OAI22_X1 U7627 ( .A1(n6650), .A2(n6657), .B1(n6649), .B2(n6648), .ZN(n6709)
         );
  NAND2_X1 U7628 ( .A1(n6652), .A2(n6651), .ZN(n6663) );
  AOI22_X1 U7629 ( .A1(n6709), .A2(n6654), .B1(n6653), .B2(n6706), .ZN(n6668)
         );
  INV_X1 U7630 ( .A(n6715), .ZN(n6656) );
  NOR3_X1 U7631 ( .A1(n6656), .A2(n6710), .A3(n6655), .ZN(n6660) );
  OAI22_X1 U7632 ( .A1(n6660), .A2(n6659), .B1(n6658), .B2(n6657), .ZN(n6665)
         );
  AOI211_X1 U7633 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6663), .A(n6662), .B(
        n6661), .ZN(n6664) );
  NAND2_X1 U7634 ( .A1(n6665), .A2(n6664), .ZN(n6712) );
  AOI22_X1 U7635 ( .A1(n6712), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n6666), 
        .B2(n6710), .ZN(n6667) );
  OAI211_X1 U7636 ( .C1(n6669), .C2(n6715), .A(n6668), .B(n6667), .ZN(U3116)
         );
  AOI22_X1 U7637 ( .A1(n6709), .A2(n6671), .B1(n6670), .B2(n6706), .ZN(n6674)
         );
  AOI22_X1 U7638 ( .A1(n6712), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n6672), 
        .B2(n6710), .ZN(n6673) );
  OAI211_X1 U7639 ( .C1(n6675), .C2(n6715), .A(n6674), .B(n6673), .ZN(U3117)
         );
  AOI22_X1 U7640 ( .A1(n6709), .A2(n6677), .B1(n6676), .B2(n6706), .ZN(n6680)
         );
  AOI22_X1 U7641 ( .A1(n6712), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n6678), 
        .B2(n6710), .ZN(n6679) );
  OAI211_X1 U7642 ( .C1(n6681), .C2(n6715), .A(n6680), .B(n6679), .ZN(U3118)
         );
  AOI22_X1 U7643 ( .A1(n6709), .A2(n6683), .B1(n6682), .B2(n6706), .ZN(n6686)
         );
  AOI22_X1 U7644 ( .A1(n6712), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n6684), 
        .B2(n6710), .ZN(n6685) );
  OAI211_X1 U7645 ( .C1(n6687), .C2(n6715), .A(n6686), .B(n6685), .ZN(U3119)
         );
  AOI22_X1 U7646 ( .A1(n6709), .A2(n6689), .B1(n6688), .B2(n6706), .ZN(n6692)
         );
  AOI22_X1 U7647 ( .A1(n6712), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n6690), 
        .B2(n6710), .ZN(n6691) );
  OAI211_X1 U7648 ( .C1(n6693), .C2(n6715), .A(n6692), .B(n6691), .ZN(U3120)
         );
  AOI22_X1 U7649 ( .A1(n6709), .A2(n6695), .B1(n6694), .B2(n6706), .ZN(n6698)
         );
  AOI22_X1 U7650 ( .A1(n6712), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n6696), 
        .B2(n6710), .ZN(n6697) );
  OAI211_X1 U7651 ( .C1(n6699), .C2(n6715), .A(n6698), .B(n6697), .ZN(U3121)
         );
  AOI22_X1 U7652 ( .A1(n6709), .A2(n6701), .B1(n6700), .B2(n6706), .ZN(n6704)
         );
  AOI22_X1 U7653 ( .A1(n6712), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n6702), 
        .B2(n6710), .ZN(n6703) );
  OAI211_X1 U7654 ( .C1(n6705), .C2(n6715), .A(n6704), .B(n6703), .ZN(U3122)
         );
  AOI22_X1 U7655 ( .A1(n6709), .A2(n6708), .B1(n6707), .B2(n6706), .ZN(n6714)
         );
  AOI22_X1 U7656 ( .A1(n6712), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n6711), 
        .B2(n6710), .ZN(n6713) );
  OAI211_X1 U7657 ( .C1(n6716), .C2(n6715), .A(n6714), .B(n6713), .ZN(U3123)
         );
  AOI21_X1 U7658 ( .B1(n3267), .B2(n4811), .A(n6717), .ZN(n6721) );
  OAI211_X1 U7659 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(STATE2_REG_1__SCAN_IN), .B(n6718), .ZN(n6719) );
  OAI211_X1 U7660 ( .C1(n6722), .C2(n6721), .A(n6720), .B(n6719), .ZN(U3149)
         );
  OAI221_X1 U7661 ( .B1(STATE2_REG_2__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(STATE2_REG_2__SCAN_IN), .C2(n4811), .A(n6723), .ZN(n6725) );
  OAI21_X1 U7662 ( .B1(n6747), .B2(n6725), .A(n6724), .ZN(U3150) );
  AND2_X1 U7663 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6726), .ZN(U3151) );
  NOR2_X1 U7664 ( .A1(n6730), .A2(n6990), .ZN(U3152) );
  AND2_X1 U7665 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6726), .ZN(U3153) );
  AND2_X1 U7666 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6726), .ZN(U3154) );
  INV_X1 U7667 ( .A(DATAWIDTH_REG_27__SCAN_IN), .ZN(n6888) );
  NOR2_X1 U7668 ( .A1(n6730), .A2(n6888), .ZN(U3155) );
  AND2_X1 U7669 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6726), .ZN(U3156) );
  INV_X1 U7670 ( .A(DATAWIDTH_REG_25__SCAN_IN), .ZN(n7050) );
  NOR2_X1 U7671 ( .A1(n6730), .A2(n7050), .ZN(U3157) );
  INV_X1 U7672 ( .A(DATAWIDTH_REG_24__SCAN_IN), .ZN(n7002) );
  NOR2_X1 U7673 ( .A1(n6730), .A2(n7002), .ZN(U3158) );
  AND2_X1 U7674 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6726), .ZN(U3159) );
  NOR2_X1 U7675 ( .A1(n6730), .A2(n6938), .ZN(U3160) );
  AND2_X1 U7676 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6726), .ZN(U3161) );
  INV_X1 U7677 ( .A(DATAWIDTH_REG_20__SCAN_IN), .ZN(n6827) );
  NOR2_X1 U7678 ( .A1(n6730), .A2(n6827), .ZN(U3162) );
  AND2_X1 U7679 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6726), .ZN(U3163) );
  NOR2_X1 U7680 ( .A1(n6730), .A2(n7006), .ZN(U3164) );
  AND2_X1 U7681 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6726), .ZN(U3165) );
  INV_X1 U7682 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6876) );
  NOR2_X1 U7683 ( .A1(n6730), .A2(n6876), .ZN(U3166) );
  AND2_X1 U7684 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6726), .ZN(U3167) );
  AND2_X1 U7685 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6726), .ZN(U3168) );
  INV_X1 U7686 ( .A(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6859) );
  NOR2_X1 U7687 ( .A1(n6730), .A2(n6859), .ZN(U3169) );
  AND2_X1 U7688 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6726), .ZN(U3170) );
  AND2_X1 U7689 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6726), .ZN(U3171) );
  NOR2_X1 U7690 ( .A1(n6730), .A2(n6954), .ZN(U3172) );
  NOR2_X1 U7691 ( .A1(n6730), .A2(n6841), .ZN(U3173) );
  AND2_X1 U7692 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6726), .ZN(U3174) );
  INV_X1 U7693 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6921) );
  NOR2_X1 U7694 ( .A1(n6730), .A2(n6921), .ZN(U3175) );
  AND2_X1 U7695 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6726), .ZN(U3176) );
  INV_X1 U7696 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6843) );
  NOR2_X1 U7697 ( .A1(n6730), .A2(n6843), .ZN(U3177) );
  AND2_X1 U7698 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6726), .ZN(U3178) );
  AND2_X1 U7699 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6726), .ZN(U3179) );
  AND2_X1 U7700 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6726), .ZN(U3180) );
  OAI22_X1 U7701 ( .A1(n4598), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n6752), .ZN(n6727) );
  INV_X1 U7702 ( .A(n6727), .ZN(U3445) );
  MUX2_X1 U7703 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n4598), .Z(U3446) );
  INV_X1 U7704 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n6957) );
  AOI22_X1 U7705 ( .A1(n6752), .A2(n6951), .B1(n6957), .B2(n4598), .ZN(U3447)
         );
  INV_X1 U7706 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6735) );
  INV_X1 U7707 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6950) );
  AOI22_X1 U7708 ( .A1(n6752), .A2(n6735), .B1(n6950), .B2(n4598), .ZN(U3448)
         );
  OAI21_X1 U7709 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6730), .A(n6729), .ZN(
        n6728) );
  INV_X1 U7710 ( .A(n6728), .ZN(U3451) );
  OAI21_X1 U7711 ( .B1(n6730), .B2(n6821), .A(n6729), .ZN(U3452) );
  NAND2_X1 U7712 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n6734) );
  INV_X1 U7713 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6731) );
  OAI211_X1 U7714 ( .C1(n6731), .C2(n6891), .A(n6821), .B(n6737), .ZN(n6733)
         );
  NAND2_X1 U7715 ( .A1(BYTEENABLE_REG_2__SCAN_IN), .A2(n6736), .ZN(n6732) );
  OAI211_X1 U7716 ( .C1(n6734), .C2(n6736), .A(n6733), .B(n6732), .ZN(U3468)
         );
  AOI22_X1 U7717 ( .A1(n6737), .A2(n6891), .B1(n6736), .B2(n6735), .ZN(U3469)
         );
  INV_X1 U7718 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6973) );
  AOI22_X1 U7719 ( .A1(n6752), .A2(READREQUEST_REG_SCAN_IN), .B1(n6973), .B2(
        n4598), .ZN(U3470) );
  INV_X1 U7720 ( .A(MORE_REG_SCAN_IN), .ZN(n6875) );
  INV_X1 U7721 ( .A(n6740), .ZN(n6738) );
  AOI22_X1 U7722 ( .A1(n6740), .A2(n6739), .B1(n6875), .B2(n6738), .ZN(U3471)
         );
  INV_X1 U7723 ( .A(n6741), .ZN(n6742) );
  AOI211_X1 U7724 ( .C1(n6744), .C2(n4811), .A(n6743), .B(n6742), .ZN(n6751)
         );
  OAI211_X1 U7725 ( .C1(n6746), .C2(STATEBS16_REG_SCAN_IN), .A(n6745), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6748) );
  AOI21_X1 U7726 ( .B1(n6748), .B2(STATE2_REG_0__SCAN_IN), .A(n6747), .ZN(
        n6750) );
  NAND2_X1 U7727 ( .A1(n6751), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6749) );
  OAI21_X1 U7728 ( .B1(n6751), .B2(n6750), .A(n6749), .ZN(U3472) );
  OAI22_X1 U7729 ( .A1(n4598), .A2(MEMORYFETCH_REG_SCAN_IN), .B1(
        M_IO_N_REG_SCAN_IN), .B2(n6752), .ZN(n6753) );
  INV_X1 U7730 ( .A(n6753), .ZN(U3473) );
  NAND4_X1 U7731 ( .A1(DATAO_REG_18__SCAN_IN), .A2(EAX_REG_1__SCAN_IN), .A3(
        ADDRESS_REG_18__SCAN_IN), .A4(n6862), .ZN(n6754) );
  NOR3_X1 U7732 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(
        DATAO_REG_25__SCAN_IN), .A3(n6754), .ZN(n6765) );
  INV_X1 U7733 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n6840) );
  NOR4_X1 U7734 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAO_REG_24__SCAN_IN), 
        .A3(n6838), .A4(n6840), .ZN(n6755) );
  NAND3_X1 U7735 ( .A1(NA_N), .A2(DATAWIDTH_REG_5__SCAN_IN), .A3(n6755), .ZN(
        n6763) );
  INV_X1 U7736 ( .A(DATAI_26_), .ZN(n6825) );
  NOR4_X1 U7737 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(DATAI_2_), .A3(
        DATAWIDTH_REG_1__SCAN_IN), .A4(n6825), .ZN(n6761) );
  INV_X1 U7738 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n6831) );
  NOR4_X1 U7739 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(
        INSTQUEUE_REG_10__3__SCAN_IN), .A3(DATAO_REG_5__SCAN_IN), .A4(n6831), 
        .ZN(n6760) );
  NOR4_X1 U7740 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(
        INSTQUEUE_REG_2__6__SCAN_IN), .A3(n5090), .A4(n6811), .ZN(n6759) );
  INV_X1 U7741 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n6757) );
  NOR4_X1 U7742 ( .A1(n6809), .A2(n6757), .A3(n6756), .A4(DATAI_31_), .ZN(
        n6758) );
  NAND4_X1 U7743 ( .A1(n6761), .A2(n6760), .A3(n6759), .A4(n6758), .ZN(n6762)
         );
  NOR4_X1 U7744 ( .A1(INSTQUEUE_REG_8__6__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .A3(n6763), .A4(n6762), .ZN(n6764) );
  NAND4_X1 U7745 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6765), .A3(n6764), 
        .A4(n6858), .ZN(n6805) );
  INV_X1 U7746 ( .A(DATAI_18_), .ZN(n6912) );
  NOR4_X1 U7747 ( .A1(n6906), .A2(n4646), .A3(n6912), .A4(n6910), .ZN(n6769)
         );
  NOR4_X1 U7748 ( .A1(EAX_REG_30__SCAN_IN), .A2(DATAO_REG_8__SCAN_IN), .A3(
        n6907), .A4(n6913), .ZN(n6768) );
  NOR4_X1 U7749 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(
        INSTQUEUE_REG_5__2__SCAN_IN), .A3(DATAI_24_), .A4(n6766), .ZN(n6767)
         );
  AND4_X1 U7750 ( .A1(n6769), .A2(n6768), .A3(UWORD_REG_3__SCAN_IN), .A4(n6767), .ZN(n6776) );
  NAND4_X1 U7751 ( .A1(INSTADDRPOINTER_REG_31__SCAN_IN), .A2(DATAI_16_), .A3(
        n6770), .A4(n7008), .ZN(n6774) );
  NAND4_X1 U7752 ( .A1(EAX_REG_4__SCAN_IN), .A2(UWORD_REG_0__SCAN_IN), .A3(
        LWORD_REG_14__SCAN_IN), .A4(n4725), .ZN(n6773) );
  INV_X1 U7753 ( .A(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n7041) );
  INV_X1 U7754 ( .A(EAX_REG_21__SCAN_IN), .ZN(n7033) );
  NAND4_X1 U7755 ( .A1(INSTQUEUE_REG_6__3__SCAN_IN), .A2(
        INSTQUEUE_REG_14__3__SCAN_IN), .A3(n7041), .A4(n7033), .ZN(n6772) );
  NAND4_X1 U7756 ( .A1(EBX_REG_8__SCAN_IN), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .A3(DATAO_REG_10__SCAN_IN), .A4(n3782), .ZN(n6771) );
  NOR4_X1 U7757 ( .A1(n6774), .A2(n6773), .A3(n6772), .A4(n6771), .ZN(n6775)
         );
  NAND2_X1 U7758 ( .A1(n6776), .A2(n6775), .ZN(n6804) );
  NAND4_X1 U7759 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6878), .A3(n6881), 
        .A4(n6892), .ZN(n6780) );
  NAND4_X1 U7760 ( .A1(MORE_REG_SCAN_IN), .A2(ADDRESS_REG_11__SCAN_IN), .A3(
        DATAWIDTH_REG_16__SCAN_IN), .A4(n6872), .ZN(n6779) );
  NAND4_X1 U7761 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .A3(DATAI_15_), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n6778) );
  INV_X1 U7762 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n6895) );
  NAND4_X1 U7763 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), 
        .A3(n4048), .A4(n6895), .ZN(n6777) );
  OR4_X1 U7764 ( .A1(n6780), .A2(n6779), .A3(n6778), .A4(n6777), .ZN(n6803) );
  NAND4_X1 U7765 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(EAX_REG_27__SCAN_IN), 
        .A3(BYTEENABLE_REG_1__SCAN_IN), .A4(n6953), .ZN(n6787) );
  INV_X1 U7766 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n6782) );
  NAND4_X1 U7767 ( .A1(n6782), .A2(n6781), .A3(INSTQUEUE_REG_3__4__SCAN_IN), 
        .A4(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n6786) );
  INV_X1 U7768 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n6784) );
  AND2_X1 U7769 ( .A1(REIP_REG_4__SCAN_IN), .A2(REIP_REG_5__SCAN_IN), .ZN(
        n6783) );
  NAND4_X1 U7770 ( .A1(n6784), .A2(n7040), .A3(DATAWIDTH_REG_30__SCAN_IN), 
        .A4(n6783), .ZN(n6785) );
  NOR3_X1 U7771 ( .A1(n6787), .A2(n6786), .A3(n6785), .ZN(n6793) );
  NAND4_X1 U7772 ( .A1(EBX_REG_25__SCAN_IN), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .A3(BE_N_REG_0__SCAN_IN), .A4(BE_N_REG_1__SCAN_IN), .ZN(n6790) );
  INV_X1 U7773 ( .A(DATAI_29_), .ZN(n6788) );
  NAND4_X1 U7774 ( .A1(n6788), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .A3(
        INSTQUEUE_REG_3__7__SCAN_IN), .A4(ADDRESS_REG_23__SCAN_IN), .ZN(n6789)
         );
  NOR2_X1 U7775 ( .A1(n6790), .A2(n6789), .ZN(n6792) );
  INV_X1 U7776 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n6989) );
  INV_X1 U7777 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n6982) );
  INV_X1 U7778 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n6986) );
  AND4_X1 U7779 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n6982), .A3(n6986), 
        .A4(n6988), .ZN(n6791) );
  NAND4_X1 U7780 ( .A1(n6793), .A2(n6792), .A3(n6989), .A4(n6791), .ZN(n6796)
         );
  NOR4_X1 U7781 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(HOLD), .A3(
        LWORD_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6794) );
  NAND3_X1 U7782 ( .A1(BE_N_REG_3__SCAN_IN), .A2(n6794), .A3(n5817), .ZN(n6795) );
  NOR2_X1 U7783 ( .A1(n6796), .A2(n6795), .ZN(n6801) );
  NOR4_X1 U7784 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(
        INSTQUEUE_REG_11__3__SCAN_IN), .A3(DATAO_REG_23__SCAN_IN), .A4(n7006), 
        .ZN(n6800) );
  INV_X1 U7785 ( .A(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n7018) );
  NOR4_X1 U7786 ( .A1(DATAI_19_), .A2(D_C_N_REG_SCAN_IN), .A3(n7020), .A4(
        n7018), .ZN(n6799) );
  INV_X1 U7787 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n6967) );
  NAND4_X1 U7788 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(
        INSTQUEUE_REG_13__3__SCAN_IN), .A3(REIP_REG_8__SCAN_IN), .A4(n6967), 
        .ZN(n6797) );
  NOR3_X1 U7789 ( .A1(M_IO_N_REG_SCAN_IN), .A2(W_R_N_REG_SCAN_IN), .A3(n6797), 
        .ZN(n6798) );
  NAND4_X1 U7790 ( .A1(n6801), .A2(n6800), .A3(n6799), .A4(n6798), .ZN(n6802)
         );
  NOR4_X1 U7791 ( .A1(n6805), .A2(n6804), .A3(n6803), .A4(n6802), .ZN(n6806)
         );
  NOR2_X1 U7792 ( .A1(n6806), .A2(LWORD_REG_11__SCAN_IN), .ZN(n7070) );
  INV_X1 U7793 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6808) );
  AOI22_X1 U7794 ( .A1(n6809), .A2(keyinput27), .B1(n6808), .B2(keyinput54), 
        .ZN(n6807) );
  OAI221_X1 U7795 ( .B1(n6809), .B2(keyinput27), .C1(n6808), .C2(keyinput54), 
        .A(n6807), .ZN(n6819) );
  AOI22_X1 U7796 ( .A1(n5090), .A2(keyinput75), .B1(keyinput107), .B2(n6811), 
        .ZN(n6810) );
  OAI221_X1 U7797 ( .B1(n5090), .B2(keyinput75), .C1(n6811), .C2(keyinput107), 
        .A(n6810), .ZN(n6818) );
  INV_X1 U7798 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n6812) );
  XOR2_X1 U7799 ( .A(n6812), .B(keyinput10), .Z(n6816) );
  XNOR2_X1 U7800 ( .A(keyinput21), .B(DATAI_31_), .ZN(n6815) );
  XNOR2_X1 U7801 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .B(keyinput90), .ZN(n6814)
         );
  XNOR2_X1 U7802 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .B(keyinput106), .ZN(n6813) );
  NAND4_X1 U7803 ( .A1(n6816), .A2(n6815), .A3(n6814), .A4(n6813), .ZN(n6817)
         );
  NOR3_X1 U7804 ( .A1(n6819), .A2(n6818), .A3(n6817), .ZN(n6870) );
  AOI22_X1 U7805 ( .A1(n6822), .A2(keyinput65), .B1(keyinput17), .B2(n6821), 
        .ZN(n6820) );
  OAI221_X1 U7806 ( .B1(n6822), .B2(keyinput65), .C1(n6821), .C2(keyinput17), 
        .A(n6820), .ZN(n6835) );
  INV_X1 U7807 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n6824) );
  AOI22_X1 U7808 ( .A1(n6825), .A2(keyinput121), .B1(n6824), .B2(keyinput2), 
        .ZN(n6823) );
  OAI221_X1 U7809 ( .B1(n6825), .B2(keyinput121), .C1(n6824), .C2(keyinput2), 
        .A(n6823), .ZN(n6834) );
  INV_X1 U7810 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n6828) );
  AOI22_X1 U7811 ( .A1(n6828), .A2(keyinput33), .B1(keyinput48), .B2(n6827), 
        .ZN(n6826) );
  OAI221_X1 U7812 ( .B1(n6828), .B2(keyinput33), .C1(n6827), .C2(keyinput48), 
        .A(n6826), .ZN(n6833) );
  INV_X1 U7813 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6830) );
  AOI22_X1 U7814 ( .A1(n6831), .A2(keyinput60), .B1(keyinput49), .B2(n6830), 
        .ZN(n6829) );
  OAI221_X1 U7815 ( .B1(n6831), .B2(keyinput60), .C1(n6830), .C2(keyinput49), 
        .A(n6829), .ZN(n6832) );
  NOR4_X1 U7816 ( .A1(n6835), .A2(n6834), .A3(n6833), .A4(n6832), .ZN(n6869)
         );
  AOI22_X1 U7817 ( .A1(n6838), .A2(keyinput67), .B1(keyinput31), .B2(n6837), 
        .ZN(n6836) );
  OAI221_X1 U7818 ( .B1(n6838), .B2(keyinput67), .C1(n6837), .C2(keyinput31), 
        .A(n6836), .ZN(n6851) );
  AOI22_X1 U7819 ( .A1(n6841), .A2(keyinput63), .B1(keyinput43), .B2(n6840), 
        .ZN(n6839) );
  OAI221_X1 U7820 ( .B1(n6841), .B2(keyinput63), .C1(n6840), .C2(keyinput43), 
        .A(n6839), .ZN(n6850) );
  AOI22_X1 U7821 ( .A1(n6844), .A2(keyinput110), .B1(keyinput76), .B2(n6843), 
        .ZN(n6842) );
  OAI221_X1 U7822 ( .B1(n6844), .B2(keyinput110), .C1(n6843), .C2(keyinput76), 
        .A(n6842), .ZN(n6849) );
  INV_X1 U7823 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n6846) );
  AOI22_X1 U7824 ( .A1(n6847), .A2(keyinput38), .B1(n6846), .B2(keyinput97), 
        .ZN(n6845) );
  OAI221_X1 U7825 ( .B1(n6847), .B2(keyinput38), .C1(n6846), .C2(keyinput97), 
        .A(n6845), .ZN(n6848) );
  NOR4_X1 U7826 ( .A1(n6851), .A2(n6850), .A3(n6849), .A4(n6848), .ZN(n6868)
         );
  AOI22_X1 U7827 ( .A1(n6853), .A2(keyinput62), .B1(keyinput100), .B2(n4726), 
        .ZN(n6852) );
  OAI221_X1 U7828 ( .B1(n6853), .B2(keyinput62), .C1(n4726), .C2(keyinput100), 
        .A(n6852), .ZN(n6866) );
  AOI22_X1 U7829 ( .A1(n6856), .A2(keyinput119), .B1(n6855), .B2(keyinput6), 
        .ZN(n6854) );
  OAI221_X1 U7830 ( .B1(n6856), .B2(keyinput119), .C1(n6855), .C2(keyinput6), 
        .A(n6854), .ZN(n6865) );
  AOI22_X1 U7831 ( .A1(n6859), .A2(keyinput77), .B1(n6858), .B2(keyinput72), 
        .ZN(n6857) );
  OAI221_X1 U7832 ( .B1(n6859), .B2(keyinput77), .C1(n6858), .C2(keyinput72), 
        .A(n6857), .ZN(n6864) );
  AOI22_X1 U7833 ( .A1(n6862), .A2(keyinput18), .B1(keyinput115), .B2(n6861), 
        .ZN(n6860) );
  OAI221_X1 U7834 ( .B1(n6862), .B2(keyinput18), .C1(n6861), .C2(keyinput115), 
        .A(n6860), .ZN(n6863) );
  NOR4_X1 U7835 ( .A1(n6866), .A2(n6865), .A3(n6864), .A4(n6863), .ZN(n6867)
         );
  NAND4_X1 U7836 ( .A1(n6870), .A2(n6869), .A3(n6868), .A4(n6867), .ZN(n7068)
         );
  AOI22_X1 U7837 ( .A1(n6873), .A2(keyinput61), .B1(n6872), .B2(keyinput117), 
        .ZN(n6871) );
  OAI221_X1 U7838 ( .B1(n6873), .B2(keyinput61), .C1(n6872), .C2(keyinput117), 
        .A(n6871), .ZN(n6886) );
  AOI22_X1 U7839 ( .A1(n6876), .A2(keyinput15), .B1(n6875), .B2(keyinput126), 
        .ZN(n6874) );
  OAI221_X1 U7840 ( .B1(n6876), .B2(keyinput15), .C1(n6875), .C2(keyinput126), 
        .A(n6874), .ZN(n6885) );
  AOI22_X1 U7841 ( .A1(n6879), .A2(keyinput3), .B1(n6878), .B2(keyinput96), 
        .ZN(n6877) );
  OAI221_X1 U7842 ( .B1(n6879), .B2(keyinput3), .C1(n6878), .C2(keyinput96), 
        .A(n6877), .ZN(n6884) );
  AOI22_X1 U7843 ( .A1(n6882), .A2(keyinput4), .B1(n6881), .B2(keyinput109), 
        .ZN(n6880) );
  OAI221_X1 U7844 ( .B1(n6882), .B2(keyinput4), .C1(n6881), .C2(keyinput109), 
        .A(n6880), .ZN(n6883) );
  NOR4_X1 U7845 ( .A1(n6886), .A2(n6885), .A3(n6884), .A4(n6883), .ZN(n6934)
         );
  AOI22_X1 U7846 ( .A1(n6889), .A2(keyinput127), .B1(keyinput79), .B2(n6888), 
        .ZN(n6887) );
  OAI221_X1 U7847 ( .B1(n6889), .B2(keyinput127), .C1(n6888), .C2(keyinput79), 
        .A(n6887), .ZN(n6901) );
  AOI22_X1 U7848 ( .A1(n6892), .A2(keyinput108), .B1(keyinput99), .B2(n6891), 
        .ZN(n6890) );
  OAI221_X1 U7849 ( .B1(n6892), .B2(keyinput108), .C1(n6891), .C2(keyinput99), 
        .A(n6890), .ZN(n6900) );
  AOI22_X1 U7850 ( .A1(n4048), .A2(keyinput105), .B1(keyinput113), .B2(n6894), 
        .ZN(n6893) );
  OAI221_X1 U7851 ( .B1(n4048), .B2(keyinput105), .C1(n6894), .C2(keyinput113), 
        .A(n6893), .ZN(n6899) );
  XOR2_X1 U7852 ( .A(n6895), .B(keyinput125), .Z(n6897) );
  XNOR2_X1 U7853 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .B(keyinput56), .ZN(n6896)
         );
  NAND2_X1 U7854 ( .A1(n6897), .A2(n6896), .ZN(n6898) );
  NOR4_X1 U7855 ( .A1(n6901), .A2(n6900), .A3(n6899), .A4(n6898), .ZN(n6933)
         );
  INV_X1 U7856 ( .A(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n6904) );
  AOI22_X1 U7857 ( .A1(n6904), .A2(keyinput112), .B1(keyinput82), .B2(n6903), 
        .ZN(n6902) );
  OAI221_X1 U7858 ( .B1(n6904), .B2(keyinput112), .C1(n6903), .C2(keyinput82), 
        .A(n6902), .ZN(n6917) );
  AOI22_X1 U7859 ( .A1(n6907), .A2(keyinput98), .B1(keyinput80), .B2(n6906), 
        .ZN(n6905) );
  OAI221_X1 U7860 ( .B1(n6907), .B2(keyinput98), .C1(n6906), .C2(keyinput80), 
        .A(n6905), .ZN(n6916) );
  AOI22_X1 U7861 ( .A1(n6910), .A2(keyinput24), .B1(keyinput123), .B2(n6909), 
        .ZN(n6908) );
  OAI221_X1 U7862 ( .B1(n6910), .B2(keyinput24), .C1(n6909), .C2(keyinput123), 
        .A(n6908), .ZN(n6915) );
  AOI22_X1 U7863 ( .A1(n6913), .A2(keyinput55), .B1(keyinput58), .B2(n6912), 
        .ZN(n6911) );
  OAI221_X1 U7864 ( .B1(n6913), .B2(keyinput55), .C1(n6912), .C2(keyinput58), 
        .A(n6911), .ZN(n6914) );
  NOR4_X1 U7865 ( .A1(n6917), .A2(n6916), .A3(n6915), .A4(n6914), .ZN(n6932)
         );
  INV_X1 U7866 ( .A(DATAI_24_), .ZN(n6919) );
  AOI22_X1 U7867 ( .A1(n6919), .A2(keyinput12), .B1(keyinput102), .B2(n4659), 
        .ZN(n6918) );
  OAI221_X1 U7868 ( .B1(n6919), .B2(keyinput12), .C1(n4659), .C2(keyinput102), 
        .A(n6918), .ZN(n6930) );
  INV_X1 U7869 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n6922) );
  AOI22_X1 U7870 ( .A1(n6922), .A2(keyinput92), .B1(keyinput13), .B2(n6921), 
        .ZN(n6920) );
  OAI221_X1 U7871 ( .B1(n6922), .B2(keyinput92), .C1(n6921), .C2(keyinput13), 
        .A(n6920), .ZN(n6929) );
  INV_X1 U7872 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n6924) );
  AOI22_X1 U7873 ( .A1(n4646), .A2(keyinput71), .B1(n6924), .B2(keyinput41), 
        .ZN(n6923) );
  OAI221_X1 U7874 ( .B1(n4646), .B2(keyinput71), .C1(n6924), .C2(keyinput41), 
        .A(n6923), .ZN(n6928) );
  XNOR2_X1 U7875 ( .A(INSTQUEUE_REG_3__7__SCAN_IN), .B(keyinput28), .ZN(n6926)
         );
  XNOR2_X1 U7876 ( .A(keyinput53), .B(DATAI_29_), .ZN(n6925) );
  NAND2_X1 U7877 ( .A1(n6926), .A2(n6925), .ZN(n6927) );
  NOR4_X1 U7878 ( .A1(n6930), .A2(n6929), .A3(n6928), .A4(n6927), .ZN(n6931)
         );
  NAND4_X1 U7879 ( .A1(n6934), .A2(n6933), .A3(n6932), .A4(n6931), .ZN(n7067)
         );
  AOI22_X1 U7880 ( .A1(n5817), .A2(keyinput25), .B1(keyinput40), .B2(n6936), 
        .ZN(n6935) );
  OAI221_X1 U7881 ( .B1(n5817), .B2(keyinput25), .C1(n6936), .C2(keyinput40), 
        .A(n6935), .ZN(n6948) );
  AOI22_X1 U7882 ( .A1(n6782), .A2(keyinput51), .B1(keyinput22), .B2(n6938), 
        .ZN(n6937) );
  OAI221_X1 U7883 ( .B1(n6782), .B2(keyinput51), .C1(n6938), .C2(keyinput22), 
        .A(n6937), .ZN(n6947) );
  INV_X1 U7884 ( .A(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n6941) );
  AOI22_X1 U7885 ( .A1(n6941), .A2(keyinput8), .B1(keyinput44), .B2(n6940), 
        .ZN(n6939) );
  OAI221_X1 U7886 ( .B1(n6941), .B2(keyinput8), .C1(n6940), .C2(keyinput44), 
        .A(n6939), .ZN(n6946) );
  INV_X1 U7887 ( .A(LWORD_REG_10__SCAN_IN), .ZN(n6942) );
  XOR2_X1 U7888 ( .A(keyinput50), .B(n6942), .Z(n6944) );
  XNOR2_X1 U7889 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .B(keyinput94), .ZN(n6943)
         );
  NAND2_X1 U7890 ( .A1(n6944), .A2(n6943), .ZN(n6945) );
  NOR4_X1 U7891 ( .A1(n6948), .A2(n6947), .A3(n6946), .A4(n6945), .ZN(n7000)
         );
  AOI22_X1 U7892 ( .A1(n6951), .A2(keyinput118), .B1(keyinput95), .B2(n6950), 
        .ZN(n6949) );
  OAI221_X1 U7893 ( .B1(n6951), .B2(keyinput118), .C1(n6950), .C2(keyinput95), 
        .A(n6949), .ZN(n6964) );
  AOI22_X1 U7894 ( .A1(n6954), .A2(keyinput69), .B1(n6953), .B2(keyinput87), 
        .ZN(n6952) );
  OAI221_X1 U7895 ( .B1(n6954), .B2(keyinput69), .C1(n6953), .C2(keyinput87), 
        .A(n6952), .ZN(n6963) );
  INV_X1 U7896 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n6956) );
  AOI22_X1 U7897 ( .A1(n6957), .A2(keyinput32), .B1(keyinput0), .B2(n6956), 
        .ZN(n6955) );
  OAI221_X1 U7898 ( .B1(n6957), .B2(keyinput32), .C1(n6956), .C2(keyinput0), 
        .A(n6955), .ZN(n6962) );
  AOI22_X1 U7899 ( .A1(n6960), .A2(keyinput101), .B1(n6959), .B2(keyinput1), 
        .ZN(n6958) );
  OAI221_X1 U7900 ( .B1(n6960), .B2(keyinput101), .C1(n6959), .C2(keyinput1), 
        .A(n6958), .ZN(n6961) );
  NOR4_X1 U7901 ( .A1(n6964), .A2(n6963), .A3(n6962), .A4(n6961), .ZN(n6999)
         );
  INV_X1 U7902 ( .A(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n6966) );
  AOI22_X1 U7903 ( .A1(n6967), .A2(keyinput66), .B1(keyinput26), .B2(n6966), 
        .ZN(n6965) );
  OAI221_X1 U7904 ( .B1(n6967), .B2(keyinput66), .C1(n6966), .C2(keyinput26), 
        .A(n6965), .ZN(n6980) );
  INV_X1 U7905 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n6970) );
  INV_X1 U7906 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n6969) );
  AOI22_X1 U7907 ( .A1(n6970), .A2(keyinput104), .B1(keyinput114), .B2(n6969), 
        .ZN(n6968) );
  OAI221_X1 U7908 ( .B1(n6970), .B2(keyinput104), .C1(n6969), .C2(keyinput114), 
        .A(n6968), .ZN(n6979) );
  INV_X1 U7909 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n6972) );
  AOI22_X1 U7910 ( .A1(n6973), .A2(keyinput91), .B1(n6972), .B2(keyinput68), 
        .ZN(n6971) );
  OAI221_X1 U7911 ( .B1(n6973), .B2(keyinput91), .C1(n6972), .C2(keyinput68), 
        .A(n6971), .ZN(n6978) );
  XOR2_X1 U7912 ( .A(n6974), .B(keyinput37), .Z(n6976) );
  XNOR2_X1 U7913 ( .A(n6756), .B(keyinput19), .ZN(n6975) );
  NAND2_X1 U7914 ( .A1(n6976), .A2(n6975), .ZN(n6977) );
  NOR4_X1 U7915 ( .A1(n6980), .A2(n6979), .A3(n6978), .A4(n6977), .ZN(n6998)
         );
  AOI22_X1 U7916 ( .A1(n6983), .A2(keyinput29), .B1(n6982), .B2(keyinput52), 
        .ZN(n6981) );
  OAI221_X1 U7917 ( .B1(n6983), .B2(keyinput29), .C1(n6982), .C2(keyinput52), 
        .A(n6981), .ZN(n6996) );
  INV_X1 U7918 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6985) );
  AOI22_X1 U7919 ( .A1(n6986), .A2(keyinput88), .B1(keyinput9), .B2(n6985), 
        .ZN(n6984) );
  OAI221_X1 U7920 ( .B1(n6986), .B2(keyinput88), .C1(n6985), .C2(keyinput9), 
        .A(n6984), .ZN(n6995) );
  AOI22_X1 U7921 ( .A1(n6989), .A2(keyinput57), .B1(n6988), .B2(keyinput120), 
        .ZN(n6987) );
  OAI221_X1 U7922 ( .B1(n6989), .B2(keyinput57), .C1(n6988), .C2(keyinput120), 
        .A(n6987), .ZN(n6994) );
  XOR2_X1 U7923 ( .A(n6990), .B(keyinput122), .Z(n6992) );
  XNOR2_X1 U7924 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .B(keyinput116), .ZN(n6991) );
  NAND2_X1 U7925 ( .A1(n6992), .A2(n6991), .ZN(n6993) );
  NOR4_X1 U7926 ( .A1(n6996), .A2(n6995), .A3(n6994), .A4(n6993), .ZN(n6997)
         );
  NAND4_X1 U7927 ( .A1(n7000), .A2(n6999), .A3(n6998), .A4(n6997), .ZN(n7066)
         );
  AOI22_X1 U7928 ( .A1(n7003), .A2(keyinput70), .B1(keyinput93), .B2(n7002), 
        .ZN(n7001) );
  OAI221_X1 U7929 ( .B1(n7003), .B2(keyinput70), .C1(n7002), .C2(keyinput93), 
        .A(n7001), .ZN(n7015) );
  INV_X1 U7930 ( .A(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n7005) );
  AOI22_X1 U7931 ( .A1(n7006), .A2(keyinput78), .B1(n7005), .B2(keyinput59), 
        .ZN(n7004) );
  OAI221_X1 U7932 ( .B1(n7006), .B2(keyinput78), .C1(n7005), .C2(keyinput59), 
        .A(n7004), .ZN(n7014) );
  AOI22_X1 U7933 ( .A1(n7009), .A2(keyinput30), .B1(n7008), .B2(keyinput84), 
        .ZN(n7007) );
  OAI221_X1 U7934 ( .B1(n7009), .B2(keyinput30), .C1(n7008), .C2(keyinput84), 
        .A(n7007), .ZN(n7013) );
  AOI22_X1 U7935 ( .A1(n4725), .A2(keyinput36), .B1(keyinput45), .B2(n7011), 
        .ZN(n7010) );
  OAI221_X1 U7936 ( .B1(n4725), .B2(keyinput36), .C1(n7011), .C2(keyinput45), 
        .A(n7010), .ZN(n7012) );
  NOR4_X1 U7937 ( .A1(n7015), .A2(n7014), .A3(n7013), .A4(n7012), .ZN(n7064)
         );
  AOI22_X1 U7938 ( .A1(keyinput124), .A2(n7018), .B1(keyinput14), .B2(n7016), 
        .ZN(n7017) );
  OAI21_X1 U7939 ( .B1(n7018), .B2(keyinput124), .A(n7017), .ZN(n7031) );
  INV_X1 U7940 ( .A(D_C_N_REG_SCAN_IN), .ZN(n7021) );
  AOI22_X1 U7941 ( .A1(n7021), .A2(keyinput74), .B1(n7020), .B2(keyinput89), 
        .ZN(n7019) );
  OAI221_X1 U7942 ( .B1(n7021), .B2(keyinput74), .C1(n7020), .C2(keyinput89), 
        .A(n7019), .ZN(n7030) );
  AOI22_X1 U7943 ( .A1(n7024), .A2(keyinput23), .B1(keyinput47), .B2(n7023), 
        .ZN(n7022) );
  OAI221_X1 U7944 ( .B1(n7024), .B2(keyinput23), .C1(n7023), .C2(keyinput47), 
        .A(n7022), .ZN(n7029) );
  INV_X1 U7945 ( .A(DATAI_19_), .ZN(n7027) );
  INV_X1 U7946 ( .A(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n7026) );
  AOI22_X1 U7947 ( .A1(n7027), .A2(keyinput34), .B1(n7026), .B2(keyinput20), 
        .ZN(n7025) );
  OAI221_X1 U7948 ( .B1(n7027), .B2(keyinput34), .C1(n7026), .C2(keyinput20), 
        .A(n7025), .ZN(n7028) );
  NOR4_X1 U7949 ( .A1(n7031), .A2(n7030), .A3(n7029), .A4(n7028), .ZN(n7063)
         );
  INV_X1 U7950 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n7034) );
  AOI22_X1 U7951 ( .A1(n7034), .A2(keyinput83), .B1(keyinput11), .B2(n7033), 
        .ZN(n7032) );
  OAI221_X1 U7952 ( .B1(n7034), .B2(keyinput83), .C1(n7033), .C2(keyinput11), 
        .A(n7032), .ZN(n7045) );
  INV_X1 U7953 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n7036) );
  AOI22_X1 U7954 ( .A1(n3782), .A2(keyinput5), .B1(n7036), .B2(keyinput42), 
        .ZN(n7035) );
  OAI221_X1 U7955 ( .B1(n3782), .B2(keyinput5), .C1(n7036), .C2(keyinput42), 
        .A(n7035), .ZN(n7044) );
  INV_X1 U7956 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n7038) );
  AOI22_X1 U7957 ( .A1(n4003), .A2(keyinput39), .B1(n7038), .B2(keyinput7), 
        .ZN(n7037) );
  OAI221_X1 U7958 ( .B1(n4003), .B2(keyinput39), .C1(n7038), .C2(keyinput7), 
        .A(n7037), .ZN(n7043) );
  AOI22_X1 U7959 ( .A1(n7041), .A2(keyinput16), .B1(n7040), .B2(keyinput85), 
        .ZN(n7039) );
  OAI221_X1 U7960 ( .B1(n7041), .B2(keyinput16), .C1(n7040), .C2(keyinput85), 
        .A(n7039), .ZN(n7042) );
  NOR4_X1 U7961 ( .A1(n7045), .A2(n7044), .A3(n7043), .A4(n7042), .ZN(n7062)
         );
  AOI22_X1 U7962 ( .A1(n7048), .A2(keyinput73), .B1(keyinput86), .B2(n7047), 
        .ZN(n7046) );
  OAI221_X1 U7963 ( .B1(n7048), .B2(keyinput73), .C1(n7047), .C2(keyinput86), 
        .A(n7046), .ZN(n7060) );
  AOI22_X1 U7964 ( .A1(n7051), .A2(keyinput81), .B1(keyinput46), .B2(n7050), 
        .ZN(n7049) );
  OAI221_X1 U7965 ( .B1(n7051), .B2(keyinput81), .C1(n7050), .C2(keyinput46), 
        .A(n7049), .ZN(n7059) );
  INV_X1 U7966 ( .A(DATAI_16_), .ZN(n7054) );
  INV_X1 U7967 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n7053) );
  AOI22_X1 U7968 ( .A1(n7054), .A2(keyinput35), .B1(keyinput103), .B2(n7053), 
        .ZN(n7052) );
  OAI221_X1 U7969 ( .B1(n7054), .B2(keyinput35), .C1(n7053), .C2(keyinput103), 
        .A(n7052), .ZN(n7058) );
  XNOR2_X1 U7970 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(keyinput64), .ZN(
        n7056) );
  XNOR2_X1 U7971 ( .A(keyinput111), .B(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n7055) );
  NAND2_X1 U7972 ( .A1(n7056), .A2(n7055), .ZN(n7057) );
  NOR4_X1 U7973 ( .A1(n7060), .A2(n7059), .A3(n7058), .A4(n7057), .ZN(n7061)
         );
  NAND4_X1 U7974 ( .A1(n7064), .A2(n7063), .A3(n7062), .A4(n7061), .ZN(n7065)
         );
  NOR4_X1 U7975 ( .A1(n7068), .A2(n7067), .A3(n7066), .A4(n7065), .ZN(n7069)
         );
  OAI21_X1 U7976 ( .B1(keyinput14), .B2(n7070), .A(n7069), .ZN(n7084) );
  OAI22_X1 U7977 ( .A1(n7074), .A2(n7073), .B1(n7072), .B2(n7071), .ZN(n7075)
         );
  AOI21_X1 U7978 ( .B1(n7077), .B2(n7076), .A(n7075), .ZN(n7080) );
  NAND2_X1 U7979 ( .A1(n7078), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n7079) );
  OAI211_X1 U7980 ( .C1(n7082), .C2(n7081), .A(n7080), .B(n7079), .ZN(n7083)
         );
  XNOR2_X1 U7981 ( .A(n7084), .B(n7083), .ZN(U3066) );
  AND4_X1 U4377 ( .A1(n3304), .A2(n3303), .A3(n3302), .A4(n3301), .ZN(n3305)
         );
  CLKBUF_X1 U3572 ( .A(n6076), .Z(n3105) );
  CLKBUF_X1 U3597 ( .A(n3423), .Z(n3788) );
  NAND2_X2 U3700 ( .A1(n3277), .A2(n4677), .ZN(n3362) );
  CLKBUF_X1 U3705 ( .A(n3636), .Z(n3114) );
  CLKBUF_X1 U4018 ( .A(n3412), .Z(n4925) );
  CLKBUF_X1 U4101 ( .A(n5523), .Z(n5524) );
  CLKBUF_X1 U4180 ( .A(n5068), .Z(n5150) );
  AND2_X2 U4239 ( .A1(n5430), .A2(n3228), .ZN(n5406) );
  CLKBUF_X1 U6657 ( .A(n5027), .Z(n5028) );
  CLKBUF_X1 U6671 ( .A(n5506), .Z(n5507) );
endmodule

