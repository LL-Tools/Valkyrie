

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4303, n4304, n4305, n4306, n4307, n4308, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380;

  INV_X4 U4809 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NAND2_X1 U4810 ( .A1(n5470), .A2(n5469), .ZN(n9578) );
  OR2_X1 U4811 ( .A1(n7318), .A2(n10101), .ZN(n10102) );
  INV_X1 U4812 ( .A(n4310), .ZN(n9192) );
  INV_X2 U4813 ( .A(n8584), .ZN(n8591) );
  INV_X1 U4814 ( .A(n5746), .ZN(n5976) );
  BUF_X1 U4815 ( .A(n9100), .Z(n6472) );
  CLKBUF_X2 U4816 ( .A(n8172), .Z(n4312) );
  XNOR2_X2 U4817 ( .A(n5726), .B(n5710), .ZN(n9100) );
  OR2_X1 U4818 ( .A1(n6096), .A2(n6095), .ZN(n4441) );
  NAND2_X1 U4819 ( .A1(n4500), .A2(n4370), .ZN(n8888) );
  INV_X1 U4820 ( .A(n5772), .ZN(n5949) );
  NAND2_X1 U4821 ( .A1(n8440), .A2(n8603), .ZN(n8584) );
  NAND2_X1 U4822 ( .A1(n8208), .A2(n5769), .ZN(n8491) );
  NAND2_X1 U4823 ( .A1(n8450), .A2(n8451), .ZN(n10255) );
  NOR2_X1 U4824 ( .A1(n9578), .A2(n9577), .ZN(n9581) );
  NAND2_X1 U4825 ( .A1(n4955), .A2(n5364), .ZN(n5272) );
  INV_X1 U4826 ( .A(n8623), .ZN(n8482) );
  NAND2_X1 U4828 ( .A1(n6883), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6922) );
  OAI21_X1 U4829 ( .B1(n8773), .B2(n6057), .A(n6058), .ZN(n8765) );
  CLKBUF_X3 U4830 ( .A(n5761), .Z(n8565) );
  INV_X1 U4831 ( .A(n8624), .ZN(n7265) );
  AND3_X1 U4832 ( .A1(n6130), .A2(n6129), .A3(n6128), .ZN(n6135) );
  NAND2_X1 U4833 ( .A1(n9243), .A2(n7761), .ZN(n9252) );
  NAND2_X1 U4834 ( .A1(n9215), .A2(n7795), .ZN(n9146) );
  NAND2_X1 U4835 ( .A1(n5547), .A2(n5546), .ZN(n9203) );
  XNOR2_X1 U4836 ( .A(n8765), .B(n8764), .ZN(n4519) );
  INV_X1 U4837 ( .A(n8436), .ZN(n8311) );
  XNOR2_X1 U4838 ( .A(n5748), .B(n5763), .ZN(n6372) );
  NAND4_X2 U4839 ( .A1(n5018), .A2(n5017), .A3(n5016), .A4(n5015), .ZN(n8050)
         );
  INV_X1 U4840 ( .A(n5614), .ZN(n10147) );
  OR2_X1 U4841 ( .A1(n6237), .A2(n6236), .ZN(n8169) );
  AOI211_X1 U4842 ( .C1(n10223), .C2(n9715), .A(n9714), .B(n9713), .ZN(n9785)
         );
  AND2_X1 U4843 ( .A1(n6605), .A2(n6604), .ZN(n8345) );
  INV_X2 U4844 ( .A(n9663), .ZN(n10130) );
  NAND2_X1 U4845 ( .A1(n6412), .A2(n8727), .ZN(n6416) );
  NOR2_X2 U4846 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n6094) );
  NAND2_X2 U4847 ( .A1(n9401), .A2(n10180), .ZN(n10124) );
  OAI21_X2 U4848 ( .B1(n7458), .B2(n5622), .A(n7973), .ZN(n7510) );
  XNOR2_X2 U4849 ( .A(n4751), .B(n6445), .ZN(n6883) );
  AND3_X2 U4850 ( .A1(n6091), .A2(n5707), .A3(n5706), .ZN(n6085) );
  NAND2_X1 U4851 ( .A1(n7092), .A2(n7091), .ZN(n8388) );
  AND2_X2 U4852 ( .A1(n4984), .A2(SI_1_), .ZN(n5030) );
  NOR2_X2 U4853 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n6121) );
  XNOR2_X2 U4854 ( .A(n5614), .B(n8050), .ZN(n10145) );
  NOR2_X1 U4855 ( .A1(n5705), .A2(n5854), .ZN(n5708) );
  NOR3_X1 U4856 ( .A1(n8876), .A2(n8890), .A3(n8403), .ZN(n8404) );
  AOI21_X2 U4857 ( .B1(n9223), .B2(n9225), .A(n9224), .ZN(n9227) );
  NAND2_X2 U4858 ( .A1(n7717), .A2(n7716), .ZN(n9223) );
  OR2_X2 U4859 ( .A1(n9401), .A2(n10180), .ZN(n7949) );
  XNOR2_X2 U4860 ( .A(n5010), .B(n5009), .ZN(n6639) );
  OAI21_X2 U4861 ( .B1(n7377), .B2(n5869), .A(n5868), .ZN(n7556) );
  OAI22_X2 U4862 ( .A1(n7344), .A2(n5851), .B1(n7539), .B2(n7451), .ZN(n7377)
         );
  NOR2_X2 U4863 ( .A1(n8228), .A2(n8227), .ZN(n8231) );
  XNOR2_X2 U4864 ( .A(n5383), .B(n5382), .ZN(n8151) );
  AOI21_X2 U4865 ( .B1(n6338), .B2(P1_REG1_REG_4__SCAN_IN), .A(n9431), .ZN(
        n9444) );
  AND2_X2 U4866 ( .A1(n9433), .A2(n9434), .ZN(n9431) );
  AOI21_X1 U4867 ( .B1(n4519), .B2(n10257), .A(n4516), .ZN(n9016) );
  NAND2_X1 U4868 ( .A1(n8779), .A2(n8786), .ZN(n4879) );
  OAI21_X1 U4869 ( .B1(n8812), .B2(n4901), .A(n4385), .ZN(n6191) );
  NAND2_X1 U4870 ( .A1(n8080), .A2(n8079), .ZN(n8142) );
  XNOR2_X1 U4871 ( .A(n6216), .B(n6215), .ZN(n7910) );
  NAND2_X1 U4872 ( .A1(n9546), .A2(n5638), .ZN(n8021) );
  INV_X1 U4873 ( .A(n9203), .ZN(n4303) );
  NAND2_X1 U4874 ( .A1(n5453), .A2(n5452), .ZN(n9731) );
  NAND2_X1 U4875 ( .A1(n7495), .A2(n6405), .ZN(n6406) );
  NAND2_X1 U4876 ( .A1(n5415), .A2(n5414), .ZN(n5430) );
  NAND2_X1 U4877 ( .A1(n7342), .A2(n8477), .ZN(n7379) );
  NAND2_X1 U4878 ( .A1(n10224), .A2(n9211), .ZN(n7969) );
  NAND2_X1 U4879 ( .A1(n5155), .A2(n5154), .ZN(n10224) );
  INV_X1 U4880 ( .A(n7539), .ZN(n7263) );
  INV_X1 U4881 ( .A(n7354), .ZN(n7206) );
  INV_X1 U4882 ( .A(n5754), .ZN(n10278) );
  NAND2_X1 U4883 ( .A1(n5760), .A2(n5759), .ZN(n10260) );
  CLKBUF_X2 U4884 ( .A(n5046), .Z(n5647) );
  CLKBUF_X1 U4885 ( .A(n5746), .Z(n8363) );
  BUF_X2 U4886 ( .A(n4337), .Z(n8366) );
  NAND2_X2 U4887 ( .A1(n8189), .A2(n10002), .ZN(n5014) );
  INV_X2 U4888 ( .A(n6641), .ZN(n5517) );
  INV_X2 U4889 ( .A(n5073), .ZN(n5659) );
  INV_X2 U4890 ( .A(n5073), .ZN(n4304) );
  INV_X1 U4891 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5837) );
  OR2_X1 U4892 ( .A1(n9788), .A2(n9773), .ZN(n4418) );
  OR2_X1 U4893 ( .A1(n8612), .A2(n4423), .ZN(n8615) );
  AOI21_X1 U4894 ( .B1(n8601), .B2(n8600), .A(n8599), .ZN(n8612) );
  AOI211_X1 U4895 ( .C1(n8167), .C2(n8166), .A(n8165), .B(n8164), .ZN(n8181)
         );
  MUX2_X1 U4896 ( .A(n9786), .B(n9785), .S(n10232), .Z(n9787) );
  AOI21_X1 U4897 ( .B1(n6199), .B2(n6511), .A(n6510), .ZN(n6512) );
  MUX2_X1 U4898 ( .A(n6249), .B(n9867), .S(n10230), .Z(n6247) );
  MUX2_X1 U4899 ( .A(n6249), .B(n6248), .S(n10245), .Z(n6250) );
  NOR2_X1 U4900 ( .A1(n9719), .A2(n4428), .ZN(n4427) );
  NOR2_X1 U4901 ( .A1(n9792), .A2(n4426), .ZN(n4425) );
  AOI21_X1 U4902 ( .B1(n6199), .B2(n6198), .A(n6197), .ZN(n6200) );
  OR2_X1 U4903 ( .A1(n8581), .A2(n8577), .ZN(n8589) );
  CLKBUF_X1 U4904 ( .A(n9621), .Z(n4422) );
  AND2_X1 U4905 ( .A1(n9710), .A2(n9709), .ZN(n9781) );
  NAND2_X1 U4906 ( .A1(n9621), .A2(n4664), .ZN(n4663) );
  NAND2_X1 U4907 ( .A1(n5409), .A2(n5408), .ZN(n9621) );
  NAND2_X1 U4908 ( .A1(n4746), .A2(n6416), .ZN(n8730) );
  OAI21_X1 U4909 ( .B1(n8169), .B2(n9373), .A(n8102), .ZN(n8107) );
  OAI21_X1 U4910 ( .B1(n4879), .B2(n4472), .A(n4469), .ZN(n6256) );
  NAND2_X1 U4911 ( .A1(n9532), .A2(n4818), .ZN(n4817) );
  AND2_X1 U4912 ( .A1(n8365), .A2(n8364), .ZN(n9012) );
  NAND2_X1 U4913 ( .A1(n4545), .A2(n9552), .ZN(n9532) );
  NAND2_X1 U4914 ( .A1(n9567), .A2(n9550), .ZN(n4545) );
  OAI21_X1 U4915 ( .B1(n4318), .B2(n4921), .A(n4376), .ZN(n4920) );
  OR2_X2 U4916 ( .A1(n9715), .A2(n9116), .ZN(n8080) );
  NAND2_X1 U4917 ( .A1(n9564), .A2(n5637), .ZN(n9567) );
  NAND2_X2 U4918 ( .A1(n5524), .A2(n5523), .ZN(n9715) );
  NAND2_X1 U4919 ( .A1(n9375), .A2(n4303), .ZN(n8042) );
  NOR2_X1 U4920 ( .A1(n9789), .A2(n9812), .ZN(n4426) );
  NAND2_X1 U4921 ( .A1(n9607), .A2(n5636), .ZN(n9564) );
  NOR2_X1 U4922 ( .A1(n9789), .A2(n9743), .ZN(n4428) );
  AOI21_X1 U4923 ( .B1(n4870), .B2(n4876), .A(n4395), .ZN(n4869) );
  NAND2_X1 U4924 ( .A1(n8426), .A2(n8554), .ZN(n8786) );
  AOI21_X1 U4925 ( .B1(n4665), .B2(n4662), .A(n4661), .ZN(n4660) );
  NAND2_X1 U4926 ( .A1(n6207), .A2(SI_29_), .ZN(n6223) );
  NAND2_X1 U4927 ( .A1(n4645), .A2(n4412), .ZN(n10080) );
  OAI21_X1 U4928 ( .B1(n10000), .B2(n5039), .A(n5670), .ZN(n5688) );
  NAND2_X1 U4929 ( .A1(n7759), .A2(n7758), .ZN(n9243) );
  AOI21_X1 U4930 ( .B1(n4593), .B2(n4931), .A(n4592), .ZN(n4591) );
  NAND2_X1 U4931 ( .A1(n6048), .A2(n6047), .ZN(n9024) );
  AND2_X1 U4932 ( .A1(n4873), .A2(n4871), .ZN(n4870) );
  NAND2_X1 U4933 ( .A1(n4770), .A2(n5505), .ZN(n9546) );
  XNOR2_X1 U4934 ( .A(n5522), .B(n5521), .ZN(n9098) );
  NAND2_X1 U4935 ( .A1(n4884), .A2(n4331), .ZN(n8874) );
  NAND2_X1 U4936 ( .A1(n5285), .A2(n5284), .ZN(n7626) );
  OAI211_X1 U4937 ( .C1(n5669), .C2(n5668), .A(n5667), .B(n5666), .ZN(n10000)
         );
  NOR2_X1 U4938 ( .A1(n9598), .A2(n7803), .ZN(n4661) );
  AND2_X1 U4939 ( .A1(n4811), .A2(n4557), .ZN(n4556) );
  NAND2_X1 U4940 ( .A1(n5489), .A2(n5488), .ZN(n9558) );
  CLKBUF_X1 U4941 ( .A(n8916), .Z(n4308) );
  XNOR2_X1 U4942 ( .A(n5515), .B(n5532), .ZN(n7678) );
  OAI21_X1 U4943 ( .B1(n6007), .B2(n4835), .A(n4465), .ZN(n4463) );
  AOI21_X1 U4944 ( .B1(n8855), .B2(n4908), .A(n4906), .ZN(n4905) );
  AOI21_X1 U4945 ( .B1(n8828), .B2(n8829), .A(n8814), .ZN(n4465) );
  NAND2_X1 U4946 ( .A1(n6017), .A2(n6016), .ZN(n9042) );
  INV_X1 U4947 ( .A(n4908), .ZN(n4907) );
  NAND2_X1 U4948 ( .A1(n6009), .A2(n6008), .ZN(n9048) );
  NAND2_X1 U4949 ( .A1(n5436), .A2(n5435), .ZN(n9806) );
  AND2_X1 U4950 ( .A1(n4325), .A2(n4810), .ZN(n4809) );
  OR2_X1 U4951 ( .A1(n8980), .A2(n8893), .ZN(n8532) );
  AND2_X1 U4952 ( .A1(n8077), .A2(n8083), .ZN(n9657) );
  XNOR2_X1 U4953 ( .A(n5462), .B(n5461), .ZN(n7576) );
  NAND2_X1 U4954 ( .A1(n6406), .A2(n6904), .ZN(n6407) );
  INV_X1 U4955 ( .A(n8881), .ZN(n8980) );
  OR2_X1 U4956 ( .A1(n9754), .A2(n5632), .ZN(n8076) );
  OAI21_X1 U4957 ( .B1(n7580), .B2(n5892), .A(n5893), .ZN(n7639) );
  OR2_X1 U4958 ( .A1(n8976), .A2(n8873), .ZN(n8536) );
  NAND2_X1 U4959 ( .A1(n5988), .A2(n5987), .ZN(n9054) );
  AND2_X1 U4960 ( .A1(n5963), .A2(n5962), .ZN(n8881) );
  INV_X1 U4961 ( .A(n4777), .ZN(n5481) );
  NAND2_X1 U4962 ( .A1(n5978), .A2(n5977), .ZN(n8976) );
  NAND2_X1 U4963 ( .A1(n7028), .A2(n7027), .ZN(n7026) );
  OR2_X1 U4964 ( .A1(n10023), .A2(n10022), .ZN(n4640) );
  NAND2_X1 U4965 ( .A1(n5998), .A2(n5997), .ZN(n9060) );
  OR2_X1 U4966 ( .A1(n7143), .A2(n5039), .ZN(n5372) );
  OAI22_X1 U4967 ( .A1(n5430), .A2(n4778), .B1(n4783), .B2(n4780), .ZN(n4777)
         );
  AOI21_X1 U4968 ( .B1(n7615), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7610), .ZN(
        n10023) );
  OAI21_X1 U4969 ( .B1(n7498), .B2(n7497), .A(n7496), .ZN(n7500) );
  NAND2_X1 U4970 ( .A1(n8285), .A2(n6536), .ZN(n7017) );
  AND2_X1 U4971 ( .A1(n8528), .A2(n8518), .ZN(n8915) );
  NAND2_X1 U4972 ( .A1(n5942), .A2(n5941), .ZN(n9073) );
  AND2_X1 U4973 ( .A1(n7371), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7498) );
  NAND2_X1 U4974 ( .A1(n5338), .A2(n5337), .ZN(n9828) );
  NAND2_X1 U4975 ( .A1(n9307), .A2(n7727), .ZN(n8064) );
  NAND2_X1 U4976 ( .A1(n4382), .A2(n7387), .ZN(n7658) );
  NAND2_X1 U4977 ( .A1(n5315), .A2(n5314), .ZN(n9764) );
  NAND2_X1 U4978 ( .A1(n5933), .A2(n5932), .ZN(n8986) );
  NAND2_X1 U4979 ( .A1(n5911), .A2(n5910), .ZN(n9092) );
  NAND2_X1 U4980 ( .A1(n5899), .A2(n5898), .ZN(n8436) );
  NAND2_X1 U4981 ( .A1(n5811), .A2(n5810), .ZN(n7245) );
  NAND2_X1 U4982 ( .A1(n5293), .A2(n5292), .ZN(n9835) );
  NAND2_X1 U4983 ( .A1(n5884), .A2(n5883), .ZN(n7840) );
  NAND2_X1 U4984 ( .A1(n5309), .A2(n5308), .ZN(n5331) );
  AND2_X1 U4985 ( .A1(n5245), .A2(n5262), .ZN(n6819) );
  AND2_X1 U4986 ( .A1(n5265), .A2(n5226), .ZN(n6790) );
  NOR2_X1 U4987 ( .A1(n10323), .A2(n6509), .ZN(n6510) );
  NAND2_X1 U4988 ( .A1(n5861), .A2(n5860), .ZN(n8481) );
  NAND2_X1 U4989 ( .A1(n5872), .A2(n5871), .ZN(n8997) );
  NAND2_X1 U4990 ( .A1(n5208), .A2(n5207), .ZN(n9169) );
  AND2_X1 U4991 ( .A1(n8470), .A2(n8500), .ZN(n8393) );
  OR2_X1 U4992 ( .A1(n5221), .A2(n5220), .ZN(n4791) );
  INV_X1 U4993 ( .A(n6537), .ZN(n10299) );
  AND2_X1 U4994 ( .A1(n5096), .A2(n5118), .ZN(n6658) );
  AND4_X1 U4995 ( .A1(n5820), .A2(n5819), .A3(n5818), .A4(n5817), .ZN(n7297)
         );
  NAND2_X1 U4996 ( .A1(n6194), .A2(n8613), .ZN(n6518) );
  CLKBUF_X1 U4997 ( .A(n6159), .Z(n8739) );
  NAND4_X2 U4998 ( .A1(n5778), .A2(n5777), .A3(n5776), .A4(n5775), .ZN(n8626)
         );
  CLKBUF_X3 U4999 ( .A(n7710), .Z(n7861) );
  AND3_X1 U5000 ( .A1(n5768), .A2(n5767), .A3(n4499), .ZN(n10285) );
  NAND4_X1 U5001 ( .A1(n5051), .A2(n5050), .A3(n5049), .A4(n5048), .ZN(n9399)
         );
  INV_X1 U5002 ( .A(n6159), .ZN(n6194) );
  BUF_X1 U5003 ( .A(n6833), .Z(n9402) );
  NAND4_X2 U5004 ( .A1(n5745), .A2(n5744), .A3(n5743), .A4(n5742), .ZN(n8627)
         );
  AND2_X2 U5005 ( .A1(n6831), .A2(n6832), .ZN(n7710) );
  NAND4_X1 U5006 ( .A1(n4999), .A2(n4998), .A3(n4997), .A4(n4996), .ZN(n7000)
         );
  BUF_X2 U5007 ( .A(n5046), .Z(n5682) );
  CLKBUF_X3 U5008 ( .A(n5047), .Z(n6240) );
  BUF_X2 U5009 ( .A(n5773), .Z(n5914) );
  INV_X1 U5010 ( .A(n5102), .ZN(n5552) );
  INV_X4 U5011 ( .A(n5039), .ZN(n6217) );
  XNOR2_X1 U5012 ( .A(n5576), .B(P1_IR_REG_21__SCAN_IN), .ZN(n8172) );
  CLKBUF_X2 U5013 ( .A(n5727), .Z(n5773) );
  AND2_X1 U5014 ( .A1(n5957), .A2(n5956), .ZN(n5960) );
  AND2_X1 U5015 ( .A1(n5718), .A2(n5716), .ZN(n5727) );
  NAND2_X1 U5016 ( .A1(n5762), .A2(n5517), .ZN(n5746) );
  NAND2_X1 U5017 ( .A1(n5014), .A2(n6640), .ZN(n5039) );
  XNOR2_X1 U5018 ( .A(n6098), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8440) );
  AND2_X1 U5019 ( .A1(n4772), .A2(n5187), .ZN(n4462) );
  MUX2_X1 U5020 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9107), .S(n5762), .Z(n9004) );
  AOI21_X1 U5021 ( .B1(n5181), .B2(n4773), .A(n5180), .ZN(n4772) );
  NAND2_X1 U5022 ( .A1(n7895), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4966) );
  NOR2_X1 U5023 ( .A1(n5164), .A2(n4776), .ZN(n4775) );
  XNOR2_X1 U5024 ( .A(n6099), .B(n6100), .ZN(n8613) );
  NAND2_X1 U5025 ( .A1(n5188), .A2(n5186), .ZN(n5201) );
  NAND2_X1 U5026 ( .A1(n4441), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6099) );
  OR2_X1 U5027 ( .A1(n4977), .A2(n5290), .ZN(n4979) );
  NAND2_X1 U5028 ( .A1(n5369), .A2(n5368), .ZN(n5575) );
  NAND2_X1 U5029 ( .A1(n5569), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4981) );
  OAI21_X1 U5030 ( .B1(n4799), .B2(SI_3_), .A(n5076), .ZN(n5035) );
  NOR2_X1 U5031 ( .A1(n4989), .A2(n9949), .ZN(n5027) );
  XNOR2_X1 U5032 ( .A(n5178), .B(SI_9_), .ZN(n5181) );
  NAND2_X1 U5033 ( .A1(n5074), .A2(SI_5_), .ZN(n5119) );
  XNOR2_X1 U5034 ( .A(n5143), .B(SI_8_), .ZN(n5164) );
  XNOR2_X1 U5035 ( .A(n5779), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6434) );
  OAI21_X1 U5036 ( .B1(n5464), .B2(P1_DATAO_REG_0__SCAN_IN), .A(n4988), .ZN(
        n4989) );
  INV_X1 U5037 ( .A(n5272), .ZN(n4305) );
  NAND4_X1 U5038 ( .A1(n5708), .A2(n5709), .A3(n5856), .A4(n4710), .ZN(n6118)
         );
  AND3_X1 U5039 ( .A1(n4962), .A2(n4961), .A3(n5587), .ZN(n4963) );
  NAND2_X1 U5040 ( .A1(n5012), .A2(n5011), .ZN(n5363) );
  OR2_X1 U5041 ( .A1(n5765), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5789) );
  CLKBUF_X2 U5042 ( .A(n4974), .Z(n5012) );
  NAND3_X1 U5043 ( .A1(n9922), .A2(n5701), .A3(n5790), .ZN(n5855) );
  INV_X1 U5044 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6157) );
  NOR2_X1 U5045 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4951) );
  NOR2_X2 U5046 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n6091) );
  NOR2_X1 U5047 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n6083) );
  NOR2_X1 U5048 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5360) );
  INV_X1 U5049 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5790) );
  NOR2_X1 U5050 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5955) );
  INV_X4 U5051 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U5052 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9922) );
  CLKBUF_X1 U5053 ( .A(n7089), .Z(n4306) );
  CLKBUF_X1 U5054 ( .A(n7900), .Z(n4307) );
  INV_X2 U5055 ( .A(n5065), .ZN(n6239) );
  NAND2_X1 U5056 ( .A1(n9098), .A2(n6217), .ZN(n5524) );
  NAND2_X1 U5057 ( .A1(n7678), .A2(n6217), .ZN(n4770) );
  OR2_X2 U5058 ( .A1(n8646), .A2(n4383), .ZN(n4751) );
  NAND2_X2 U5059 ( .A1(n4420), .A2(n8544), .ZN(n8812) );
  OAI21_X2 U5060 ( .B1(n7626), .B2(n5301), .A(n5302), .ZN(n9689) );
  AOI21_X2 U5061 ( .B1(n7017), .B2(n7018), .A(n6539), .ZN(n7028) );
  AND2_X2 U5062 ( .A1(n4487), .A2(n4485), .ZN(n5073) );
  INV_X2 U5063 ( .A(n5659), .ZN(n6641) );
  INV_X1 U5064 ( .A(n5073), .ZN(n5500) );
  OR2_X2 U5065 ( .A1(n6924), .A2(n4729), .ZN(n4728) );
  NAND2_X2 U5066 ( .A1(n6590), .A2(n6589), .ZN(n8317) );
  BUF_X4 U5067 ( .A(n9113), .Z(n4310) );
  NAND2_X1 U5068 ( .A1(n6838), .A2(n6837), .ZN(n9113) );
  XNOR2_X1 U5069 ( .A(n6372), .B(n10271), .ZN(n6770) );
  NAND2_X4 U5070 ( .A1(n6498), .A2(n9100), .ZN(n5762) );
  XNOR2_X2 U5071 ( .A(n5725), .B(n5724), .ZN(n6498) );
  BUF_X8 U5072 ( .A(n8367), .Z(n4311) );
  NAND3_X2 U5073 ( .A1(n5734), .A2(n5733), .A3(n5732), .ZN(n6168) );
  INV_X1 U5074 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5706) );
  NAND2_X1 U5075 ( .A1(n8043), .A2(n8042), .ZN(n8094) );
  OR2_X1 U5076 ( .A1(n9036), .A2(n8783), .ZN(n8555) );
  AND2_X1 U5077 ( .A1(n6189), .A2(n8819), .ZN(n8430) );
  NAND2_X1 U5078 ( .A1(n4916), .A2(n4914), .ZN(n6609) );
  AOI21_X1 U5079 ( .B1(n4920), .B2(n4918), .A(n4915), .ZN(n4914) );
  NOR2_X1 U5080 ( .A1(n6599), .A2(n8767), .ZN(n4915) );
  INV_X1 U5081 ( .A(n8366), .ZN(n6262) );
  AND2_X1 U5082 ( .A1(n6613), .A2(n8591), .ZN(n10262) );
  INV_X2 U5083 ( .A(n8565), .ZN(n8563) );
  OR2_X1 U5084 ( .A1(n5541), .A2(n5540), .ZN(n5544) );
  NAND2_X1 U5085 ( .A1(n9301), .A2(n4314), .ZN(n4859) );
  INV_X1 U5086 ( .A(n9657), .ZN(n4558) );
  OAI21_X1 U5087 ( .B1(n4393), .B2(n4785), .A(n5461), .ZN(n4784) );
  NAND2_X1 U5088 ( .A1(n5222), .A2(SI_12_), .ZN(n5264) );
  AND2_X1 U5089 ( .A1(n5223), .A2(n4351), .ZN(n4790) );
  INV_X1 U5090 ( .A(n5224), .ZN(n5223) );
  OR2_X1 U5091 ( .A1(n8997), .A2(n8484), .ZN(n8483) );
  NAND2_X1 U5092 ( .A1(n6768), .A2(n6396), .ZN(n6397) );
  AOI21_X1 U5093 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n6660), .A(n8641), .ZN(
        n6375) );
  OR2_X1 U5094 ( .A1(n7918), .A2(n8569), .ZN(n8586) );
  AND2_X1 U5095 ( .A1(n5990), .A2(n5989), .ZN(n5992) );
  INV_X1 U5096 ( .A(n5999), .ZN(n5990) );
  AND2_X1 U5097 ( .A1(n6083), .A2(n9923), .ZN(n4752) );
  AOI21_X1 U5098 ( .B1(n4832), .B2(n4833), .A(n4971), .ZN(n4834) );
  NAND2_X1 U5099 ( .A1(n4969), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4833) );
  NAND2_X1 U5100 ( .A1(n9999), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4832) );
  AND2_X1 U5101 ( .A1(n9587), .A2(n9588), .ZN(n5636) );
  NOR2_X1 U5102 ( .A1(n5209), .A2(n7188), .ZN(n5195) );
  AND2_X1 U5103 ( .A1(n8042), .A2(n8027), .ZN(n5641) );
  INV_X1 U5104 ( .A(n4680), .ZN(n4679) );
  NAND2_X1 U5105 ( .A1(n4791), .A2(n4790), .ZN(n5265) );
  NAND2_X1 U5106 ( .A1(n4923), .A2(n4338), .ZN(n4922) );
  NAND2_X1 U5107 ( .A1(n4601), .A2(n4600), .ZN(n4599) );
  NAND2_X1 U5108 ( .A1(n4340), .A2(n4604), .ZN(n4600) );
  OR2_X1 U5109 ( .A1(n4602), .A2(n4340), .ZN(n4601) );
  NAND2_X1 U5110 ( .A1(n8483), .A2(n8505), .ZN(n6559) );
  INV_X1 U5111 ( .A(n5731), .ZN(n5772) );
  NAND2_X1 U5112 ( .A1(n8184), .A2(n5717), .ZN(n5731) );
  XNOR2_X1 U5113 ( .A(n6375), .B(n4750), .ZN(n6888) );
  INV_X1 U5114 ( .A(n7491), .ZN(n4733) );
  NAND2_X1 U5115 ( .A1(n4605), .A2(n8662), .ZN(n4609) );
  INV_X1 U5116 ( .A(n6380), .ZN(n4605) );
  AOI21_X1 U5117 ( .B1(n4321), .B2(n4461), .A(n4373), .ZN(n4457) );
  NAND2_X1 U5118 ( .A1(n5769), .A2(n10285), .ZN(n5771) );
  NAND2_X1 U5119 ( .A1(n5762), .A2(n6641), .ZN(n5761) );
  INV_X1 U5120 ( .A(n4902), .ZN(n4901) );
  OR2_X1 U5121 ( .A1(n6182), .A2(n6181), .ZN(n6183) );
  OR2_X1 U5122 ( .A1(n6307), .A2(n8603), .ZN(n10304) );
  INV_X2 U5123 ( .A(n6641), .ZN(n6640) );
  INV_X1 U5124 ( .A(n6240), .ZN(n5686) );
  NAND2_X1 U5125 ( .A1(n4655), .A2(n4654), .ZN(n4657) );
  AOI21_X1 U5126 ( .B1(n9443), .B2(n4658), .A(n9456), .ZN(n4654) );
  OR2_X1 U5127 ( .A1(n5098), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5148) );
  NAND2_X1 U5128 ( .A1(n8043), .A2(n8097), .ZN(n8138) );
  OR2_X1 U5129 ( .A1(n5506), .A2(n7874), .ZN(n5550) );
  OR2_X1 U5130 ( .A1(n4554), .A2(n4553), .ZN(n4552) );
  OR2_X1 U5131 ( .A1(n8050), .A2(n10147), .ZN(n5019) );
  INV_X1 U5132 ( .A(n5641), .ZN(n8139) );
  INV_X1 U5133 ( .A(n5672), .ZN(n9507) );
  INV_X1 U5134 ( .A(n4666), .ZN(n4665) );
  OAI21_X1 U5135 ( .B1(n4316), .B2(n9624), .A(n5445), .ZN(n4666) );
  NAND2_X1 U5136 ( .A1(n4437), .A2(n6217), .ZN(n5275) );
  INV_X1 U5137 ( .A(n6822), .ZN(n4437) );
  INV_X2 U5138 ( .A(n6218), .ZN(n5384) );
  OR2_X1 U5139 ( .A1(n5586), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n5567) );
  NAND2_X1 U5140 ( .A1(n4484), .A2(n4344), .ZN(n5381) );
  INV_X1 U5141 ( .A(n5201), .ZN(n5187) );
  NAND2_X1 U5142 ( .A1(n4771), .A2(n5146), .ZN(n5182) );
  NAND2_X1 U5143 ( .A1(n5142), .A2(n4775), .ZN(n4771) );
  NAND2_X1 U5144 ( .A1(n6073), .A2(n6072), .ZN(n8576) );
  NAND2_X1 U5145 ( .A1(n6080), .A2(n6079), .ZN(n8766) );
  OAI21_X1 U5146 ( .B1(n6113), .B2(n8871), .A(n6112), .ZN(n6313) );
  NOR2_X1 U5147 ( .A1(n6111), .A2(n6110), .ZN(n6112) );
  NOR2_X1 U5148 ( .A1(n8234), .A2(n8908), .ZN(n6110) );
  NOR2_X1 U5149 ( .A1(n4353), .A2(n4849), .ZN(n4848) );
  INV_X1 U5150 ( .A(n9206), .ZN(n4849) );
  NAND2_X1 U5151 ( .A1(n9450), .A2(n9451), .ZN(n9449) );
  NAND2_X1 U5152 ( .A1(n4544), .A2(n7963), .ZN(n7970) );
  OR3_X1 U5153 ( .A1(n8502), .A2(n6174), .A3(n8501), .ZN(n8508) );
  OAI211_X1 U5154 ( .C1(n7981), .C2(n4523), .A(n4522), .B(n4521), .ZN(n7982)
         );
  NAND2_X1 U5155 ( .A1(n4526), .A2(n4524), .ZN(n4521) );
  INV_X1 U5156 ( .A(n4524), .ZN(n4523) );
  NOR2_X1 U5157 ( .A1(n5630), .A2(n8039), .ZN(n4534) );
  AND2_X1 U5158 ( .A1(n7998), .A2(n8083), .ZN(n4529) );
  AOI21_X1 U5159 ( .B1(n8525), .B2(n8584), .A(n4721), .ZN(n4720) );
  INV_X1 U5160 ( .A(n8542), .ZN(n4718) );
  NAND2_X1 U5161 ( .A1(n4381), .A2(n4566), .ZN(n8425) );
  NOR2_X1 U5162 ( .A1(n4708), .A2(n4707), .ZN(n4706) );
  NAND2_X1 U5163 ( .A1(n8555), .A2(n8591), .ZN(n4707) );
  INV_X1 U5164 ( .A(n8553), .ZN(n4709) );
  AOI21_X1 U5165 ( .B1(n4716), .B2(n4714), .A(n4424), .ZN(n8552) );
  NAND2_X1 U5166 ( .A1(n8548), .A2(n8790), .ZN(n4424) );
  NOR2_X1 U5167 ( .A1(n4715), .A2(n4372), .ZN(n4714) );
  INV_X1 U5168 ( .A(n7685), .ZN(n4866) );
  INV_X1 U5169 ( .A(n5446), .ZN(n4785) );
  INV_X1 U5170 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5704) );
  INV_X1 U5171 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U5172 ( .A1(n5639), .A2(n4676), .ZN(n4675) );
  INV_X1 U5173 ( .A(n5514), .ZN(n4676) );
  AOI21_X1 U5174 ( .B1(n5639), .B2(n4674), .A(n4379), .ZN(n4673) );
  INV_X1 U5175 ( .A(n5513), .ZN(n4674) );
  NAND2_X1 U5176 ( .A1(n4677), .A2(n5498), .ZN(n4669) );
  NOR2_X1 U5177 ( .A1(n4675), .A2(n4672), .ZN(n4671) );
  INV_X1 U5178 ( .A(n4677), .ZN(n4672) );
  INV_X1 U5179 ( .A(n5463), .ZN(n4780) );
  NOR2_X1 U5180 ( .A1(n4785), .A2(n4780), .ZN(n4779) );
  INV_X1 U5181 ( .A(n4937), .ZN(n4781) );
  NAND2_X1 U5182 ( .A1(n4483), .A2(n5380), .ZN(n4482) );
  INV_X1 U5183 ( .A(n5395), .ZN(n4483) );
  NOR2_X1 U5184 ( .A1(n4482), .A2(n4479), .ZN(n4478) );
  INV_X1 U5185 ( .A(n5349), .ZN(n4479) );
  OAI21_X1 U5186 ( .B1(n6564), .B2(n4927), .A(n8191), .ZN(n4926) );
  OR2_X1 U5187 ( .A1(n8949), .A2(n8379), .ZN(n8594) );
  OR2_X1 U5188 ( .A1(n6397), .A2(n6647), .ZN(n4739) );
  NOR2_X1 U5189 ( .A1(n6459), .A2(n7472), .ZN(n4432) );
  NAND2_X1 U5190 ( .A1(n8714), .A2(n4410), .ZN(n6412) );
  NAND2_X1 U5191 ( .A1(n4748), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4747) );
  NOR2_X1 U5192 ( .A1(n6071), .A2(n4476), .ZN(n4475) );
  INV_X1 U5193 ( .A(n6058), .ZN(n4476) );
  INV_X1 U5194 ( .A(n6046), .ZN(n4471) );
  OR2_X1 U5195 ( .A1(n4474), .A2(n6071), .ZN(n4473) );
  NAND2_X1 U5196 ( .A1(n6057), .A2(n6058), .ZN(n4474) );
  AND2_X1 U5197 ( .A1(n5943), .A2(n4577), .ZN(n4576) );
  INV_X1 U5198 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n4577) );
  INV_X1 U5199 ( .A(n5945), .ZN(n5944) );
  AND2_X1 U5200 ( .A1(n5900), .A2(n4574), .ZN(n4573) );
  INV_X1 U5201 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n4574) );
  INV_X1 U5202 ( .A(n5902), .ZN(n5901) );
  NOR2_X1 U5203 ( .A1(n5862), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n4571) );
  INV_X1 U5204 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n4565) );
  NOR2_X1 U5205 ( .A1(n8383), .A2(n4893), .ZN(n4892) );
  INV_X1 U5206 ( .A(n8426), .ZN(n4893) );
  OR2_X1 U5207 ( .A1(n9018), .A2(n8234), .ZN(n8561) );
  OR2_X1 U5208 ( .A1(n9024), .A2(n8782), .ZN(n8558) );
  OR2_X1 U5209 ( .A1(n7451), .A2(n7263), .ZN(n8477) );
  OR2_X1 U5210 ( .A1(n7339), .A2(n7297), .ZN(n8470) );
  NOR2_X1 U5211 ( .A1(n7090), .A2(n4510), .ZN(n4509) );
  INV_X1 U5212 ( .A(n6170), .ZN(n4510) );
  INV_X1 U5213 ( .A(n6082), .ZN(n6084) );
  INV_X1 U5214 ( .A(n4856), .ZN(n4855) );
  OAI21_X1 U5215 ( .B1(n4858), .B2(n4857), .A(n7746), .ZN(n4856) );
  NAND2_X1 U5216 ( .A1(n4354), .A2(n4860), .ZN(n4857) );
  INV_X1 U5217 ( .A(n4550), .ZN(n4549) );
  OAI21_X1 U5218 ( .B1(n8138), .B2(n8042), .A(n10140), .ZN(n4550) );
  INV_X1 U5219 ( .A(n8083), .ZN(n4559) );
  NOR2_X1 U5220 ( .A1(n4813), .A2(n4812), .ZN(n4811) );
  NOR2_X1 U5221 ( .A1(n4819), .A2(n8130), .ZN(n4554) );
  NOR2_X1 U5222 ( .A1(n5230), .A2(n4494), .ZN(n4493) );
  NAND2_X1 U5223 ( .A1(n7227), .A2(n10116), .ZN(n7938) );
  NAND2_X1 U5224 ( .A1(n10138), .A2(n10137), .ZN(n4825) );
  XNOR2_X1 U5225 ( .A(n6833), .B(n5002), .ZN(n5612) );
  OR2_X1 U5226 ( .A1(n9546), .A2(n5638), .ZN(n8079) );
  AND2_X1 U5227 ( .A1(n4963), .A2(n4822), .ZN(n4821) );
  AND2_X1 U5228 ( .A1(n4978), .A2(n4980), .ZN(n4822) );
  XNOR2_X1 U5229 ( .A(n5394), .B(SI_19_), .ZN(n5395) );
  XNOR2_X1 U5230 ( .A(n5347), .B(SI_17_), .ZN(n5349) );
  NOR2_X1 U5231 ( .A1(n5328), .A2(n5327), .ZN(n5330) );
  OAI21_X1 U5232 ( .B1(n5222), .B2(SI_12_), .A(n5264), .ZN(n5224) );
  NAND2_X1 U5233 ( .A1(n5183), .A2(SI_10_), .ZN(n5188) );
  INV_X1 U5234 ( .A(n5141), .ZN(n4776) );
  AOI21_X1 U5235 ( .B1(n4911), .B2(n4913), .A(n4361), .ZN(n4909) );
  INV_X1 U5236 ( .A(n4588), .ZN(n4587) );
  OAI21_X1 U5237 ( .B1(n4319), .B2(n4589), .A(n6553), .ZN(n4588) );
  AND2_X1 U5238 ( .A1(n7593), .A2(n6552), .ZN(n6553) );
  INV_X1 U5239 ( .A(n6551), .ZN(n4589) );
  NOR2_X1 U5240 ( .A1(n6596), .A2(n4924), .ZN(n4923) );
  NOR2_X1 U5241 ( .A1(n4338), .A2(n8318), .ZN(n4924) );
  OR2_X1 U5242 ( .A1(n8414), .A2(n8413), .ZN(n8598) );
  NAND2_X1 U5243 ( .A1(n6104), .A2(n6103), .ZN(n8373) );
  INV_X1 U5244 ( .A(n7916), .ZN(n6104) );
  INV_X1 U5245 ( .A(n5949), .ZN(n8368) );
  NAND2_X1 U5246 ( .A1(n4760), .A2(n4763), .ZN(n6796) );
  OR2_X1 U5247 ( .A1(n4762), .A2(n4761), .ZN(n4758) );
  AND2_X1 U5248 ( .A1(n4754), .A2(n8637), .ZN(n6742) );
  NAND2_X1 U5249 ( .A1(n6727), .A2(n4755), .ZN(n4754) );
  NOR2_X1 U5250 ( .A1(n4324), .A2(n4756), .ZN(n4755) );
  NAND2_X1 U5251 ( .A1(n6888), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6915) );
  NAND2_X1 U5252 ( .A1(n4350), .A2(n7050), .ZN(n6376) );
  INV_X1 U5253 ( .A(n4632), .ZN(n4629) );
  NAND2_X1 U5254 ( .A1(n4635), .A2(n6683), .ZN(n4626) );
  NAND2_X1 U5255 ( .A1(n4745), .A2(n8662), .ZN(n4744) );
  AND2_X1 U5256 ( .A1(n8674), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4608) );
  NAND2_X1 U5257 ( .A1(n4749), .A2(n6487), .ZN(n4748) );
  INV_X1 U5258 ( .A(n6412), .ZN(n4749) );
  NAND3_X1 U5259 ( .A1(n4638), .A2(n4411), .A3(n4636), .ZN(n6385) );
  NOR2_X1 U5260 ( .A1(n8743), .A2(n6493), .ZN(n6500) );
  NAND2_X1 U5261 ( .A1(n6385), .A2(n8727), .ZN(n6389) );
  OR2_X1 U5262 ( .A1(n8722), .A2(n8983), .ZN(n8720) );
  INV_X1 U5263 ( .A(n8735), .ZN(n4622) );
  OAI21_X1 U5264 ( .B1(n4408), .B2(n4621), .A(n4620), .ZN(n4619) );
  NOR2_X1 U5265 ( .A1(n6386), .A2(n4622), .ZN(n4621) );
  NAND2_X1 U5266 ( .A1(n4408), .A2(n8735), .ZN(n4620) );
  INV_X1 U5267 ( .A(n8775), .ZN(n8234) );
  NOR2_X1 U5268 ( .A1(n8569), .A2(n8910), .ZN(n6111) );
  NAND2_X1 U5269 ( .A1(n6062), .A2(n6061), .ZN(n6074) );
  INV_X1 U5270 ( .A(n6063), .ZN(n6062) );
  NAND2_X1 U5271 ( .A1(n5992), .A2(n5991), .ZN(n6010) );
  INV_X1 U5272 ( .A(n8833), .ZN(n8858) );
  NAND2_X1 U5273 ( .A1(n5944), .A2(n5943), .ZN(n5964) );
  OR2_X1 U5274 ( .A1(n5934), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U5275 ( .A1(n5880), .A2(n5879), .ZN(n7580) );
  NAND2_X1 U5276 ( .A1(n4571), .A2(n4570), .ZN(n5886) );
  INV_X1 U5277 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n4570) );
  OR2_X1 U5278 ( .A1(n5803), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5825) );
  AOI21_X1 U5279 ( .B1(n4892), .B2(n4708), .A(n4890), .ZN(n4889) );
  INV_X1 U5280 ( .A(n8558), .ZN(n4890) );
  INV_X1 U5281 ( .A(n4892), .ZN(n4891) );
  AND2_X1 U5282 ( .A1(n8561), .A2(n8562), .ZN(n8764) );
  NAND2_X1 U5283 ( .A1(n8766), .A2(n10261), .ZN(n4518) );
  NAND2_X1 U5284 ( .A1(n8775), .A2(n10261), .ZN(n4445) );
  NAND2_X1 U5285 ( .A1(n8423), .A2(n9030), .ZN(n8426) );
  AND2_X1 U5286 ( .A1(n8558), .A2(n8557), .ZN(n8774) );
  NOR2_X1 U5287 ( .A1(n8430), .A2(n8429), .ZN(n4902) );
  CLKBUF_X1 U5288 ( .A(n8802), .Z(n8803) );
  OR2_X1 U5289 ( .A1(n8430), .A2(n8384), .ZN(n8804) );
  NAND2_X1 U5290 ( .A1(n8812), .A2(n8550), .ZN(n4903) );
  AND2_X1 U5291 ( .A1(n8543), .A2(n8536), .ZN(n4908) );
  NAND2_X1 U5292 ( .A1(n8544), .A2(n8545), .ZN(n8828) );
  NAND2_X1 U5293 ( .A1(n8860), .A2(n8859), .ZN(n8862) );
  OAI21_X1 U5294 ( .B1(n7583), .B2(n6179), .A(n8511), .ZN(n7646) );
  INV_X1 U5295 ( .A(n8910), .ZN(n10261) );
  OR2_X1 U5296 ( .A1(n8565), .A2(n6667), .ZN(n4499) );
  NOR2_X1 U5297 ( .A1(n4899), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4897) );
  NAND2_X1 U5298 ( .A1(n5710), .A2(n6119), .ZN(n4899) );
  INV_X1 U5299 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7188) );
  OR2_X1 U5300 ( .A1(n5169), .A2(n5158), .ZN(n5209) );
  AND2_X1 U5301 ( .A1(n9149), .A2(n7806), .ZN(n7807) );
  NAND2_X1 U5302 ( .A1(n4853), .A2(n4852), .ZN(n4851) );
  NOR2_X1 U5303 ( .A1(n9204), .A2(n9371), .ZN(n4852) );
  INV_X1 U5304 ( .A(n9205), .ZN(n4853) );
  NAND2_X1 U5305 ( .A1(n9216), .A2(n9217), .ZN(n9215) );
  INV_X1 U5306 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5230) );
  INV_X1 U5307 ( .A(n9194), .ZN(n9115) );
  NAND2_X1 U5308 ( .A1(n4840), .A2(n4838), .ZN(n4837) );
  INV_X1 U5309 ( .A(n7119), .ZN(n4838) );
  NAND3_X1 U5310 ( .A1(n6968), .A2(n6967), .A3(n4840), .ZN(n4836) );
  AND2_X1 U5311 ( .A1(n9322), .A2(n4939), .ZN(n7716) );
  OR2_X1 U5312 ( .A1(n9160), .A2(n7715), .ZN(n4939) );
  AND2_X1 U5313 ( .A1(n7869), .A2(n7866), .ZN(n7867) );
  AND3_X1 U5314 ( .A1(n5323), .A2(n5322), .A3(n5321), .ZN(n7750) );
  AND4_X1 U5315 ( .A1(n5200), .A2(n5199), .A3(n5198), .A4(n5197), .ZN(n7711)
         );
  AND4_X1 U5316 ( .A1(n5163), .A2(n5162), .A3(n5161), .A4(n5160), .ZN(n9211)
         );
  INV_X1 U5317 ( .A(n5021), .ZN(n5065) );
  NAND2_X1 U5318 ( .A1(n9448), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n4658) );
  OR2_X1 U5319 ( .A1(n9444), .A2(n9443), .ZN(n4659) );
  NOR2_X1 U5320 ( .A1(n7611), .A2(n7612), .ZN(n7610) );
  NOR2_X1 U5321 ( .A1(n10048), .A2(n4453), .ZN(n10059) );
  AND2_X1 U5322 ( .A1(n6351), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4453) );
  NAND2_X1 U5323 ( .A1(n10059), .A2(n10060), .ZN(n10058) );
  AOI21_X1 U5324 ( .B1(n10064), .B2(n4648), .A(n4414), .ZN(n4647) );
  INV_X1 U5325 ( .A(n6325), .ZN(n4648) );
  NAND2_X1 U5326 ( .A1(n4646), .A2(n10064), .ZN(n4645) );
  INV_X1 U5327 ( .A(n10043), .ZN(n4646) );
  XNOR2_X1 U5328 ( .A(n4454), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n6353) );
  NAND2_X1 U5329 ( .A1(n10074), .A2(n6352), .ZN(n4454) );
  OR2_X1 U5330 ( .A1(n10016), .A2(n10012), .ZN(n10030) );
  NAND2_X1 U5331 ( .A1(n4549), .A2(n8138), .ZN(n4548) );
  AND2_X1 U5332 ( .A1(n8148), .A2(n6931), .ZN(n9313) );
  AND2_X1 U5333 ( .A1(n5550), .A2(n5507), .ZN(n7873) );
  NAND2_X1 U5334 ( .A1(n9652), .A2(n8083), .ZN(n9640) );
  NAND2_X1 U5335 ( .A1(n9653), .A2(n9657), .ZN(n9652) );
  NAND2_X1 U5336 ( .A1(n4555), .A2(n4554), .ZN(n7627) );
  NAND2_X1 U5337 ( .A1(n7521), .A2(n5624), .ZN(n7653) );
  NAND2_X1 U5338 ( .A1(n7510), .A2(n7509), .ZN(n7521) );
  NAND2_X1 U5339 ( .A1(n7937), .A2(n4815), .ZN(n4814) );
  AND3_X1 U5340 ( .A1(n4802), .A2(n4803), .A3(n10201), .ZN(n10119) );
  NAND2_X1 U5341 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5067) );
  NAND2_X1 U5342 ( .A1(n4520), .A2(n7948), .ZN(n7070) );
  NAND2_X1 U5343 ( .A1(n10125), .A2(n8052), .ZN(n4520) );
  NAND2_X1 U5344 ( .A1(n7401), .A2(n7481), .ZN(n6837) );
  AND2_X1 U5345 ( .A1(n8044), .A2(n9563), .ZN(n9587) );
  NAND2_X1 U5346 ( .A1(n5418), .A2(n5417), .ZN(n7786) );
  NOR2_X1 U5347 ( .A1(n4684), .A2(n4377), .ZN(n4683) );
  INV_X1 U5348 ( .A(n5379), .ZN(n4684) );
  OR2_X1 U5349 ( .A1(n9672), .A2(n5378), .ZN(n4685) );
  NOR2_X1 U5350 ( .A1(n5014), .A2(n4650), .ZN(n4686) );
  NAND2_X1 U5351 ( .A1(n6641), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4800) );
  OR2_X1 U5352 ( .A1(n6837), .A2(n8106), .ZN(n10213) );
  NAND2_X1 U5353 ( .A1(n5572), .A2(n5571), .ZN(n9995) );
  NAND2_X1 U5354 ( .A1(n5516), .A2(n5531), .ZN(n5522) );
  NAND2_X1 U5355 ( .A1(n5515), .A2(n5532), .ZN(n5516) );
  INV_X1 U5356 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5563) );
  INV_X1 U5357 ( .A(n5447), .ZN(n4786) );
  AND2_X1 U5358 ( .A1(n5463), .A2(n5451), .ZN(n5461) );
  INV_X1 U5359 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5560) );
  NAND2_X1 U5360 ( .A1(n5583), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5576) );
  OAI21_X1 U5361 ( .B1(n5575), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5581) );
  NOR2_X1 U5362 ( .A1(n5363), .A2(n5362), .ZN(n5365) );
  NAND2_X1 U5363 ( .A1(n5244), .A2(n5243), .ZN(n5262) );
  NAND2_X1 U5364 ( .A1(n5270), .A2(n5269), .ZN(n5287) );
  NOR2_X1 U5365 ( .A1(n5268), .A2(n5267), .ZN(n5269) );
  INV_X1 U5366 ( .A(n5146), .ZN(n4773) );
  NOR2_X1 U5367 ( .A1(n5125), .A2(n5124), .ZN(n5126) );
  NAND2_X1 U5368 ( .A1(n5290), .A2(n5011), .ZN(n4652) );
  AOI21_X1 U5369 ( .B1(n8822), .B2(n5914), .A(n6014), .ZN(n8243) );
  NOR2_X1 U5370 ( .A1(n4597), .A2(n8345), .ZN(n4595) );
  AND2_X1 U5371 ( .A1(n4599), .A2(n4387), .ZN(n4597) );
  NAND2_X1 U5372 ( .A1(n4599), .A2(n4603), .ZN(n4598) );
  OR2_X1 U5373 ( .A1(n4340), .A2(n8280), .ZN(n4603) );
  NAND2_X1 U5374 ( .A1(n7880), .A2(n6563), .ZN(n8307) );
  NAND2_X1 U5375 ( .A1(n6056), .A2(n6055), .ZN(n8767) );
  NAND2_X1 U5376 ( .A1(n6024), .A2(n6023), .ZN(n8819) );
  AND3_X1 U5377 ( .A1(n5757), .A2(n5756), .A3(n5755), .ZN(n5760) );
  NAND2_X1 U5378 ( .A1(n4337), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U5379 ( .A1(n5772), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5745) );
  NOR2_X1 U5380 ( .A1(n4738), .A2(n4731), .ZN(n7493) );
  NAND2_X1 U5381 ( .A1(n4730), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4731) );
  INV_X1 U5382 ( .A(n8751), .ZN(n8663) );
  AND2_X1 U5383 ( .A1(n4332), .A2(n4609), .ZN(n8676) );
  NAND2_X1 U5384 ( .A1(n4766), .A2(n6478), .ZN(n4765) );
  INV_X1 U5385 ( .A(n6382), .ZN(n4766) );
  NAND2_X1 U5386 ( .A1(n6382), .A2(n8693), .ZN(n6383) );
  OAI21_X1 U5387 ( .B1(n8654), .B2(n6505), .A(n8328), .ZN(n4439) );
  AOI21_X1 U5388 ( .B1(n6270), .B2(n6269), .A(n6268), .ZN(n6275) );
  NAND2_X1 U5389 ( .A1(n6273), .A2(n4935), .ZN(n6274) );
  OR2_X1 U5390 ( .A1(n10000), .A2(n8565), .ZN(n6255) );
  AND2_X1 U5391 ( .A1(n10269), .A2(n6308), .ZN(n8945) );
  OR2_X1 U5392 ( .A1(n5762), .A2(n4433), .ZN(n5738) );
  NAND2_X1 U5393 ( .A1(n6306), .A2(n6662), .ZN(n10253) );
  INV_X1 U5394 ( .A(n8880), .ZN(n8929) );
  AND2_X1 U5395 ( .A1(n8576), .A2(n10300), .ZN(n6114) );
  NAND2_X1 U5396 ( .A1(n6028), .A2(n6027), .ZN(n9036) );
  NOR2_X1 U5397 ( .A1(n4851), .A2(n4846), .ZN(n4845) );
  AND2_X1 U5398 ( .A1(n9205), .A2(n9349), .ZN(n4850) );
  INV_X1 U5399 ( .A(n7867), .ZN(n4846) );
  OR2_X1 U5400 ( .A1(n9126), .A2(n4851), .ZN(n4847) );
  NAND2_X2 U5401 ( .A1(n5372), .A2(n5371), .ZN(n9754) );
  NAND2_X1 U5402 ( .A1(n5557), .A2(n5556), .ZN(n9375) );
  OR2_X1 U5403 ( .A1(n9200), .A2(n5552), .ZN(n5557) );
  NAND2_X1 U5404 ( .A1(n5444), .A2(n5443), .ZN(n9381) );
  OR2_X1 U5405 ( .A1(n9613), .A2(n5552), .ZN(n5444) );
  XNOR2_X1 U5406 ( .A(n9414), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9420) );
  NAND2_X1 U5407 ( .A1(n9435), .A2(n4367), .ZN(n9450) );
  AND2_X1 U5408 ( .A1(n5099), .A2(n5148), .ZN(n9462) );
  NOR2_X1 U5409 ( .A1(n7404), .A2(n4451), .ZN(n7618) );
  NOR2_X1 U5410 ( .A1(n6346), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4451) );
  NAND2_X1 U5411 ( .A1(n7618), .A2(n7617), .ZN(n7616) );
  NOR2_X1 U5412 ( .A1(n10020), .A2(n10019), .ZN(n10018) );
  NAND2_X1 U5413 ( .A1(n5600), .A2(n9996), .ZN(n9660) );
  NAND2_X1 U5414 ( .A1(n5688), .A2(n9771), .ZN(n5698) );
  AND2_X1 U5415 ( .A1(n7844), .A2(n10248), .ZN(n4827) );
  NOR2_X1 U5416 ( .A1(n10248), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n4826) );
  OR2_X1 U5417 ( .A1(n6245), .A2(n6826), .ZN(n10245) );
  NAND2_X1 U5418 ( .A1(n4421), .A2(n5690), .ZN(n6296) );
  AND2_X1 U5419 ( .A1(n5676), .A2(n5675), .ZN(n5678) );
  AND2_X1 U5420 ( .A1(n5654), .A2(n9198), .ZN(n7845) );
  NOR2_X1 U5421 ( .A1(n10232), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n4828) );
  NAND2_X1 U5422 ( .A1(n8186), .A2(n6217), .ZN(n5547) );
  OR2_X1 U5423 ( .A1(n6687), .A2(n5039), .ZN(n5208) );
  NAND2_X1 U5424 ( .A1(n8444), .A2(n8443), .ZN(n4699) );
  NAND2_X1 U5425 ( .A1(n6521), .A2(n8445), .ZN(n4698) );
  NAND2_X1 U5426 ( .A1(n4696), .A2(n8591), .ZN(n4695) );
  INV_X1 U5427 ( .A(n8446), .ZN(n4696) );
  AND2_X1 U5428 ( .A1(n8065), .A2(n4375), .ZN(n4528) );
  NAND2_X1 U5429 ( .A1(n7965), .A2(n7971), .ZN(n7966) );
  NAND2_X1 U5430 ( .A1(n7970), .A2(n7964), .ZN(n7965) );
  NAND2_X1 U5431 ( .A1(n4348), .A2(n4525), .ZN(n4524) );
  INV_X1 U5432 ( .A(n8069), .ZN(n4525) );
  OAI211_X1 U5433 ( .C1(n7976), .C2(n8061), .A(n7975), .B(n8168), .ZN(n7981)
         );
  OAI21_X1 U5434 ( .B1(n4693), .B2(n4692), .A(n4690), .ZN(n8514) );
  OAI211_X1 U5435 ( .C1(n8508), .C2(n8506), .A(n8490), .B(n4328), .ZN(n4693)
         );
  AOI21_X1 U5436 ( .B1(n4691), .B2(n7583), .A(n8439), .ZN(n4690) );
  NOR2_X1 U5437 ( .A1(n8890), .A2(n4703), .ZN(n4702) );
  NOR2_X1 U5438 ( .A1(n8518), .A2(n8591), .ZN(n4703) );
  NAND2_X1 U5439 ( .A1(n7984), .A2(n4368), .ZN(n4530) );
  AOI21_X1 U5440 ( .B1(n8524), .B2(n8591), .A(n4713), .ZN(n4712) );
  NAND2_X1 U5441 ( .A1(n4378), .A2(n4719), .ZN(n4713) );
  NOR2_X1 U5442 ( .A1(n4717), .A2(n8547), .ZN(n4715) );
  INV_X1 U5443 ( .A(n8079), .ZN(n8023) );
  INV_X1 U5444 ( .A(n8427), .ZN(n4564) );
  NAND2_X1 U5445 ( .A1(n10278), .A2(n8627), .ZN(n8451) );
  AND2_X1 U5446 ( .A1(n9024), .A2(n8782), .ZN(n8383) );
  INV_X1 U5447 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n9923) );
  NAND2_X1 U5448 ( .A1(n4314), .A2(n7725), .ZN(n4860) );
  INV_X1 U5449 ( .A(n4859), .ZN(n4858) );
  INV_X1 U5450 ( .A(n4865), .ZN(n4864) );
  OAI211_X1 U5451 ( .C1(n4867), .C2(n4866), .A(n7697), .B(n7696), .ZN(n4865)
         );
  OR2_X1 U5452 ( .A1(n9275), .A2(n9207), .ZN(n7696) );
  NAND2_X1 U5453 ( .A1(n4864), .A2(n4866), .ZN(n4862) );
  INV_X1 U5454 ( .A(n8002), .ZN(n4813) );
  INV_X1 U5455 ( .A(n8000), .ZN(n4812) );
  NAND2_X1 U5456 ( .A1(n7937), .A2(n8114), .ZN(n8054) );
  INV_X1 U5457 ( .A(n9375), .ZN(n5558) );
  OAI21_X1 U5458 ( .B1(n4682), .B2(n4681), .A(n5407), .ZN(n4680) );
  INV_X1 U5459 ( .A(n5378), .ZN(n4681) );
  INV_X1 U5460 ( .A(n4683), .ZN(n4682) );
  AND2_X1 U5461 ( .A1(n5077), .A2(n5076), .ZN(n5078) );
  AND2_X1 U5462 ( .A1(n4347), .A2(n4918), .ZN(n4917) );
  INV_X1 U5463 ( .A(n8335), .ZN(n4918) );
  AND2_X1 U5464 ( .A1(n4912), .A2(n8325), .ZN(n4911) );
  OR2_X1 U5465 ( .A1(n8266), .A2(n4913), .ZN(n4912) );
  INV_X1 U5466 ( .A(n6578), .ZN(n4913) );
  NOR2_X1 U5467 ( .A1(n4346), .A2(n8280), .ZN(n4602) );
  XNOR2_X1 U5468 ( .A(n6526), .B(n10285), .ZN(n6533) );
  NOR2_X1 U5469 ( .A1(n6920), .A2(n7289), .ZN(n4729) );
  OAI21_X1 U5470 ( .B1(n4335), .B2(n6914), .A(n4633), .ZN(n4632) );
  NOR2_X1 U5471 ( .A1(n6914), .A2(n10321), .ZN(n4628) );
  NOR2_X1 U5472 ( .A1(n6914), .A2(n4631), .ZN(n4630) );
  NAND2_X1 U5473 ( .A1(n6683), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4631) );
  NAND2_X1 U5474 ( .A1(n4612), .A2(n4611), .ZN(n4610) );
  NAND2_X1 U5475 ( .A1(n7172), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4611) );
  NAND2_X1 U5476 ( .A1(n7500), .A2(n6379), .ZN(n6380) );
  OR2_X1 U5477 ( .A1(n8576), .A2(n8582), .ZN(n6253) );
  INV_X1 U5478 ( .A(n8562), .ZN(n4888) );
  NAND2_X1 U5479 ( .A1(n6026), .A2(n4460), .ZN(n4459) );
  INV_X1 U5480 ( .A(n6025), .ZN(n4460) );
  INV_X1 U5481 ( .A(n6026), .ZN(n4461) );
  INV_X1 U5482 ( .A(n6030), .ZN(n6029) );
  INV_X1 U5483 ( .A(n8627), .ZN(n5752) );
  NAND2_X1 U5484 ( .A1(n4902), .A2(n4904), .ZN(n4900) );
  INV_X1 U5485 ( .A(n8854), .ZN(n4468) );
  NAND2_X1 U5486 ( .A1(n4467), .A2(n4323), .ZN(n4466) );
  INV_X1 U5487 ( .A(n6007), .ZN(n4467) );
  NOR2_X1 U5488 ( .A1(n4323), .A2(n5986), .ZN(n4835) );
  INV_X1 U5489 ( .A(n8541), .ZN(n4906) );
  INV_X1 U5490 ( .A(n4503), .ZN(n4502) );
  OAI22_X1 U5491 ( .A1(n5919), .A2(n4504), .B1(n8933), .B2(n6567), .ZN(n4503)
         );
  NAND2_X1 U5492 ( .A1(n7637), .A2(n4505), .ZN(n4504) );
  INV_X1 U5493 ( .A(n7636), .ZN(n4505) );
  NAND2_X1 U5494 ( .A1(n7637), .A2(n4507), .ZN(n4506) );
  INV_X1 U5495 ( .A(n5919), .ZN(n4507) );
  NAND2_X1 U5496 ( .A1(n6696), .A2(n6695), .ZN(n8442) );
  NOR2_X1 U5497 ( .A1(n5908), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n5957) );
  AND2_X1 U5498 ( .A1(n5858), .A2(n5857), .ZN(n4442) );
  INV_X1 U5499 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4486) );
  NOR2_X1 U5500 ( .A1(n9334), .A2(n4878), .ZN(n4877) );
  INV_X1 U5501 ( .A(n7767), .ZN(n4878) );
  AND2_X1 U5502 ( .A1(n4407), .A2(n7231), .ZN(n4867) );
  INV_X1 U5503 ( .A(n9180), .ZN(n4871) );
  INV_X1 U5504 ( .A(n9189), .ZN(n7801) );
  NAND2_X1 U5505 ( .A1(n8096), .A2(n8095), .ZN(n8099) );
  INV_X1 U5506 ( .A(n8094), .ZN(n8095) );
  AND2_X1 U5507 ( .A1(n4640), .A2(n4639), .ZN(n6323) );
  NAND2_X1 U5508 ( .A1(n10026), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n4639) );
  OR2_X1 U5509 ( .A1(n5490), .A2(n7831), .ZN(n5506) );
  NOR2_X1 U5510 ( .A1(n9154), .A2(n9315), .ZN(n4498) );
  INV_X1 U5511 ( .A(n5438), .ZN(n5437) );
  INV_X1 U5512 ( .A(n5317), .ZN(n5316) );
  NOR2_X1 U5513 ( .A1(n5339), .A2(n4496), .ZN(n4495) );
  NAND2_X1 U5514 ( .A1(n5316), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5340) );
  OR2_X1 U5515 ( .A1(n5295), .A2(n5294), .ZN(n5317) );
  NOR2_X1 U5516 ( .A1(n9169), .A2(n7553), .ZN(n4804) );
  INV_X1 U5517 ( .A(n5067), .ZN(n4491) );
  NAND2_X1 U5518 ( .A1(n4670), .A2(n4667), .ZN(n5672) );
  INV_X1 U5519 ( .A(n4668), .ZN(n4667) );
  OAI21_X1 U5520 ( .B1(n4675), .B2(n4669), .A(n4673), .ZN(n4668) );
  NAND2_X1 U5521 ( .A1(n9378), .A2(n9558), .ZN(n4677) );
  AND2_X1 U5522 ( .A1(n4665), .A2(n4356), .ZN(n4664) );
  AND2_X1 U5523 ( .A1(n4316), .A2(n4356), .ZN(n4662) );
  AND3_X1 U5524 ( .A1(n4809), .A2(n4808), .A3(n7670), .ZN(n9646) );
  NAND2_X1 U5525 ( .A1(n6639), .A2(n6640), .ZN(n4688) );
  NAND2_X1 U5526 ( .A1(n5499), .A2(n5539), .ZN(n5515) );
  AND2_X1 U5527 ( .A1(n5531), .A2(n5504), .ZN(n5532) );
  NAND2_X1 U5528 ( .A1(n4781), .A2(n4779), .ZN(n4778) );
  INV_X1 U5529 ( .A(n4784), .ZN(n4783) );
  AND2_X1 U5530 ( .A1(n5482), .A2(n5468), .ZN(n5480) );
  INV_X1 U5531 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U5532 ( .A1(n4477), .A2(n4480), .ZN(n5411) );
  INV_X1 U5533 ( .A(n4481), .ZN(n4480) );
  OAI22_X1 U5534 ( .A1(n4344), .A2(n4482), .B1(n5394), .B2(SI_19_), .ZN(n4481)
         );
  AOI21_X1 U5535 ( .B1(n4790), .B2(n5220), .A(n4380), .ZN(n4789) );
  AND2_X1 U5536 ( .A1(n5120), .A2(n5119), .ZN(n5121) );
  NAND2_X1 U5537 ( .A1(n6253), .A2(n6251), .ZN(n8412) );
  NAND2_X1 U5538 ( .A1(n7026), .A2(n4363), .ZN(n7202) );
  AOI21_X1 U5539 ( .B1(n4930), .B2(n8218), .A(n4362), .ZN(n4593) );
  INV_X1 U5540 ( .A(n8240), .ZN(n4592) );
  NAND2_X1 U5541 ( .A1(n7295), .A2(n6551), .ZN(n7589) );
  XNOR2_X1 U5542 ( .A(n6526), .B(n6522), .ZN(n6523) );
  XNOR2_X1 U5543 ( .A(n10278), .B(n6526), .ZN(n6527) );
  NAND2_X1 U5544 ( .A1(n6576), .A2(n8266), .ZN(n8268) );
  INV_X1 U5545 ( .A(n8248), .ZN(n4921) );
  INV_X1 U5546 ( .A(n4926), .ZN(n4925) );
  AND2_X1 U5547 ( .A1(n8373), .A2(n8372), .ZN(n8413) );
  NAND2_X1 U5548 ( .A1(n5772), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5755) );
  OR2_X1 U5549 ( .A1(n6617), .A2(n6366), .ZN(n6420) );
  INV_X1 U5550 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6754) );
  NAND2_X1 U5551 ( .A1(n6398), .A2(n6718), .ZN(n6722) );
  OAI21_X1 U5552 ( .B1(n6374), .B2(n4324), .A(n4313), .ZN(n8637) );
  OR2_X1 U5553 ( .A1(n4324), .A2(n6723), .ZN(n4753) );
  AOI21_X1 U5554 ( .B1(n6740), .B2(n6739), .A(n6439), .ZN(n8631) );
  OR2_X1 U5555 ( .A1(n5821), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U5556 ( .A1(n4402), .A2(n7164), .ZN(n7166) );
  XNOR2_X1 U5557 ( .A(n4610), .B(n7367), .ZN(n7371) );
  AND2_X1 U5558 ( .A1(n4610), .A2(n4769), .ZN(n7497) );
  NAND2_X1 U5559 ( .A1(n5896), .A2(n5895), .ZN(n5908) );
  INV_X1 U5560 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5895) );
  INV_X1 U5561 ( .A(n5894), .ZN(n5896) );
  OR2_X1 U5562 ( .A1(n8656), .A2(n8655), .ZN(n8659) );
  INV_X1 U5563 ( .A(n4747), .ZN(n4746) );
  OAI21_X1 U5564 ( .B1(n8743), .B2(n8742), .A(n8741), .ZN(n8747) );
  NAND2_X1 U5565 ( .A1(n8586), .A2(n8360), .ZN(n6271) );
  OR2_X1 U5566 ( .A1(n6074), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n7916) );
  INV_X1 U5567 ( .A(n4475), .ZN(n4472) );
  AND2_X1 U5568 ( .A1(n4389), .A2(n4470), .ZN(n4469) );
  NAND2_X1 U5569 ( .A1(n4475), .A2(n4471), .ZN(n4470) );
  OR2_X1 U5570 ( .A1(n6049), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U5571 ( .A1(n6029), .A2(n4563), .ZN(n6049) );
  NOR2_X1 U5572 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n4563) );
  OR2_X1 U5573 ( .A1(n6018), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6030) );
  OR2_X1 U5574 ( .A1(n6010), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U5575 ( .A1(n5944), .A2(n4333), .ZN(n5999) );
  INV_X1 U5576 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n4575) );
  INV_X1 U5577 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n4572) );
  NAND2_X1 U5578 ( .A1(n5901), .A2(n4573), .ZN(n5924) );
  NAND2_X1 U5579 ( .A1(n5901), .A2(n5900), .ZN(n5912) );
  NAND2_X1 U5580 ( .A1(n4569), .A2(n5885), .ZN(n5902) );
  INV_X1 U5581 ( .A(n5886), .ZN(n4569) );
  INV_X1 U5582 ( .A(n6559), .ZN(n8399) );
  INV_X1 U5583 ( .A(n4571), .ZN(n5873) );
  NAND2_X1 U5584 ( .A1(n6173), .A2(n8500), .ZN(n4883) );
  NAND2_X1 U5585 ( .A1(n5844), .A2(n5843), .ZN(n5862) );
  INV_X1 U5586 ( .A(n5845), .ZN(n5844) );
  NAND2_X1 U5587 ( .A1(n4561), .A2(n4560), .ZN(n5845) );
  INV_X1 U5588 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n4560) );
  INV_X1 U5589 ( .A(n5827), .ZN(n4561) );
  AND2_X1 U5590 ( .A1(n7254), .A2(n8469), .ZN(n8392) );
  NAND2_X1 U5591 ( .A1(n4562), .A2(n5815), .ZN(n5827) );
  INV_X1 U5592 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5815) );
  INV_X1 U5593 ( .A(n5825), .ZN(n4562) );
  CLKBUF_X1 U5594 ( .A(n7134), .Z(n7251) );
  NAND2_X1 U5595 ( .A1(n4511), .A2(n6170), .ZN(n7094) );
  AND2_X1 U5596 ( .A1(n5794), .A2(n5793), .ZN(n6537) );
  INV_X1 U5597 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5782) );
  NAND2_X1 U5598 ( .A1(n8213), .A2(n4565), .ZN(n5783) );
  NAND2_X1 U5599 ( .A1(n10249), .A2(n8450), .ZN(n6982) );
  OR2_X1 U5600 ( .A1(n10304), .A2(n8440), .ZN(n6305) );
  AND2_X1 U5601 ( .A1(n6283), .A2(n8584), .ZN(n6304) );
  AND2_X1 U5602 ( .A1(n8758), .A2(n8757), .ZN(n9010) );
  INV_X1 U5603 ( .A(n8774), .ZN(n4447) );
  NAND2_X1 U5604 ( .A1(n8550), .A2(n8428), .ZN(n8813) );
  AOI21_X1 U5605 ( .B1(n8854), .B2(n5986), .A(n4323), .ZN(n8841) );
  AND2_X1 U5606 ( .A1(n5952), .A2(n5951), .ZN(n8911) );
  NAND2_X1 U5607 ( .A1(n4500), .A2(n4502), .ZN(n8923) );
  OR2_X1 U5608 ( .A1(n6521), .A2(n4700), .ZN(n9003) );
  INV_X1 U5609 ( .A(n8442), .ZN(n4700) );
  INV_X1 U5610 ( .A(n10302), .ZN(n10300) );
  AND2_X1 U5611 ( .A1(n6617), .A2(n6158), .ZN(n6662) );
  AND2_X1 U5612 ( .A1(n5709), .A2(n6119), .ZN(n4434) );
  XNOR2_X1 U5613 ( .A(n6087), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8603) );
  XNOR2_X1 U5614 ( .A(n5975), .B(P2_IR_REG_19__SCAN_IN), .ZN(n6159) );
  OR2_X1 U5615 ( .A1(n5834), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5836) );
  OR2_X1 U5616 ( .A1(n5795), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5797) );
  NAND2_X1 U5617 ( .A1(n6393), .A2(n5763), .ZN(n5765) );
  XNOR2_X1 U5618 ( .A(n5735), .B(n4623), .ZN(n6717) );
  INV_X1 U5619 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4623) );
  INV_X1 U5620 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5132) );
  AND2_X1 U5621 ( .A1(n7737), .A2(n7736), .ZN(n9136) );
  AOI21_X1 U5622 ( .B1(n4875), .B2(n4877), .A(n4874), .ZN(n4873) );
  INV_X1 U5623 ( .A(n9335), .ZN(n4874) );
  INV_X1 U5624 ( .A(n9253), .ZN(n4875) );
  INV_X1 U5625 ( .A(n4877), .ZN(n4876) );
  AND2_X1 U5626 ( .A1(n9119), .A2(n9118), .ZN(n9204) );
  OR2_X1 U5627 ( .A1(n5399), .A2(n9296), .ZN(n5420) );
  NAND2_X1 U5628 ( .A1(n5195), .A2(n4493), .ZN(n5253) );
  OR2_X1 U5629 ( .A1(n9238), .A2(n7757), .ZN(n4934) );
  NAND2_X1 U5630 ( .A1(n4836), .A2(n4366), .ZN(n7224) );
  INV_X1 U5631 ( .A(n7123), .ZN(n4839) );
  NOR2_X1 U5632 ( .A1(n7805), .A2(n7804), .ZN(n9262) );
  AND2_X1 U5633 ( .A1(n7818), .A2(n7817), .ZN(n9261) );
  AND2_X1 U5634 ( .A1(n6969), .A2(n6970), .ZN(n6967) );
  NAND2_X1 U5635 ( .A1(n4863), .A2(n7685), .ZN(n9274) );
  NAND2_X1 U5636 ( .A1(n9346), .A2(n4867), .ZN(n4863) );
  NAND2_X1 U5637 ( .A1(n5419), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5438) );
  INV_X1 U5638 ( .A(n5420), .ZN(n5419) );
  NAND2_X1 U5639 ( .A1(n7792), .A2(n7794), .ZN(n7795) );
  INV_X1 U5640 ( .A(n9391), .ZN(n7977) );
  NAND2_X1 U5641 ( .A1(n5316), .A2(n4495), .ZN(n5373) );
  NAND2_X1 U5642 ( .A1(n7765), .A2(n7766), .ZN(n7767) );
  NAND2_X1 U5643 ( .A1(n9252), .A2(n9253), .ZN(n9251) );
  INV_X1 U5644 ( .A(n9313), .ZN(n9351) );
  OR2_X1 U5645 ( .A1(n7819), .A2(n7818), .ZN(n7858) );
  OR2_X1 U5646 ( .A1(n6870), .A2(n6931), .ZN(n9353) );
  INV_X1 U5647 ( .A(n9353), .ZN(n9314) );
  AND2_X1 U5648 ( .A1(n8040), .A2(n4542), .ZN(n4541) );
  NAND2_X1 U5649 ( .A1(n9503), .A2(n8168), .ZN(n4542) );
  NAND2_X1 U5650 ( .A1(n8036), .A2(n8035), .ZN(n4543) );
  NOR2_X1 U5651 ( .A1(n8038), .A2(n4355), .ZN(n4792) );
  AOI21_X1 U5652 ( .B1(n9526), .B2(n5529), .A(n5528), .ZN(n9116) );
  AND4_X1 U5653 ( .A1(n5215), .A2(n5214), .A3(n5213), .A4(n5212), .ZN(n7460)
         );
  AND4_X1 U5654 ( .A1(n5072), .A2(n5071), .A3(n5070), .A4(n5069), .ZN(n9352)
         );
  INV_X1 U5655 ( .A(n4834), .ZN(n4830) );
  AND2_X1 U5656 ( .A1(n6328), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6637) );
  AND2_X1 U5657 ( .A1(n4657), .A2(n4656), .ZN(n9471) );
  NAND2_X1 U5658 ( .A1(n9462), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n4656) );
  NOR2_X1 U5659 ( .A1(n9469), .A2(n4644), .ZN(n9485) );
  AND2_X1 U5660 ( .A1(n9476), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n4644) );
  NOR2_X1 U5661 ( .A1(n9485), .A2(n9484), .ZN(n9483) );
  NOR2_X1 U5662 ( .A1(n9483), .A2(n4643), .ZN(n7009) );
  AND2_X1 U5663 ( .A1(n9490), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n4643) );
  NAND2_X1 U5664 ( .A1(n7009), .A2(n7010), .ZN(n7008) );
  OR2_X1 U5665 ( .A1(n5205), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5227) );
  AOI21_X1 U5666 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n7196), .A(n7191), .ZN(
        n7308) );
  NOR2_X1 U5667 ( .A1(n7306), .A2(n4642), .ZN(n7408) );
  AND2_X1 U5668 ( .A1(n7311), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4642) );
  NAND2_X1 U5669 ( .A1(n7408), .A2(n7409), .ZN(n7407) );
  NAND2_X1 U5670 ( .A1(n7407), .A2(n4641), .ZN(n7611) );
  OR2_X1 U5671 ( .A1(n6346), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n4641) );
  XNOR2_X1 U5672 ( .A(n6323), .B(n4450), .ZN(n10033) );
  NOR2_X1 U5673 ( .A1(n10033), .A2(n10032), .ZN(n10031) );
  NOR2_X1 U5674 ( .A1(n10018), .A2(n4405), .ZN(n6349) );
  OR2_X1 U5675 ( .A1(n10057), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4452) );
  NAND2_X1 U5676 ( .A1(n4339), .A2(n10076), .ZN(n10074) );
  NOR2_X1 U5677 ( .A1(n4807), .A2(n9503), .ZN(n4805) );
  AND2_X1 U5678 ( .A1(n9537), .A2(n8047), .ZN(n4818) );
  NAND2_X1 U5679 ( .A1(n8143), .A2(n5635), .ZN(n9607) );
  AND2_X1 U5680 ( .A1(n9646), .A2(n9813), .ZN(n9628) );
  NAND2_X1 U5681 ( .A1(n9628), .A2(n9612), .ZN(n9611) );
  OR2_X1 U5682 ( .A1(n5387), .A2(n9184), .ZN(n5399) );
  AND2_X1 U5683 ( .A1(n7670), .A2(n5608), .ZN(n9673) );
  AND2_X1 U5684 ( .A1(n4555), .A2(n8068), .ZN(n4948) );
  AND2_X1 U5685 ( .A1(n4493), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n4492) );
  OR2_X1 U5686 ( .A1(n5277), .A2(n5276), .ZN(n5295) );
  NAND2_X1 U5687 ( .A1(n7387), .A2(n4320), .ZN(n7528) );
  NAND2_X1 U5688 ( .A1(n5195), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5231) );
  NAND2_X1 U5689 ( .A1(n7390), .A2(n7971), .ZN(n7458) );
  CLKBUF_X1 U5690 ( .A(n7383), .Z(n7386) );
  CLKBUF_X1 U5691 ( .A(n7276), .Z(n7277) );
  OR2_X1 U5692 ( .A1(n5133), .A2(n5132), .ZN(n5169) );
  NOR2_X1 U5693 ( .A1(n10116), .A2(n7320), .ZN(n4801) );
  NAND2_X1 U5694 ( .A1(n7937), .A2(n7936), .ZN(n10108) );
  NAND2_X1 U5695 ( .A1(n4802), .A2(n4803), .ZN(n10117) );
  OR2_X1 U5696 ( .A1(n6837), .A2(n8171), .ZN(n9693) );
  NAND2_X1 U5697 ( .A1(n4491), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5104) );
  NAND2_X1 U5698 ( .A1(n4825), .A2(n4823), .ZN(n10125) );
  NOR2_X1 U5699 ( .A1(n5616), .A2(n4824), .ZN(n4823) );
  INV_X1 U5700 ( .A(n5615), .ZN(n4824) );
  NAND2_X1 U5701 ( .A1(n4825), .A2(n5615), .ZN(n7947) );
  NOR2_X1 U5702 ( .A1(n10146), .A2(n10147), .ZN(n10151) );
  INV_X1 U5703 ( .A(n9693), .ZN(n10148) );
  INV_X1 U5704 ( .A(n5612), .ZN(n8119) );
  NAND2_X1 U5705 ( .A1(n4817), .A2(n4816), .ZN(n5643) );
  AND2_X1 U5706 ( .A1(n5640), .A2(n8021), .ZN(n4816) );
  AND2_X1 U5707 ( .A1(n8079), .A2(n8021), .ZN(n9537) );
  AND2_X1 U5708 ( .A1(n8047), .A2(n8020), .ZN(n9552) );
  XNOR2_X1 U5709 ( .A(n9578), .B(n8015), .ZN(n9571) );
  NAND2_X1 U5710 ( .A1(n9689), .A2(n9690), .ZN(n5325) );
  AOI22_X1 U5711 ( .A1(n5384), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6236), .B2(
        n9462), .ZN(n5100) );
  AND2_X1 U5712 ( .A1(n10095), .A2(n9779), .ZN(n10195) );
  INV_X1 U5713 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4964) );
  INV_X1 U5714 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4978) );
  XNOR2_X1 U5715 ( .A(n5562), .B(P1_IR_REG_25__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U5716 ( .A1(n5567), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U5717 ( .A1(n4787), .A2(n5429), .ZN(n5448) );
  INV_X1 U5718 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5368) );
  INV_X1 U5719 ( .A(n5367), .ZN(n5369) );
  CLKBUF_X1 U5720 ( .A(n5272), .Z(n5289) );
  NAND2_X1 U5721 ( .A1(n4791), .A2(n4351), .ZN(n5225) );
  NAND2_X1 U5722 ( .A1(n5142), .A2(n5141), .ZN(n5165) );
  NAND2_X1 U5723 ( .A1(n4455), .A2(n5028), .ZN(n4992) );
  OR2_X1 U5724 ( .A1(n5073), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4988) );
  NAND2_X1 U5725 ( .A1(n7026), .A2(n6542), .ZN(n7204) );
  NAND2_X1 U5726 ( .A1(n8305), .A2(n6566), .ZN(n8192) );
  AND4_X1 U5727 ( .A1(n5878), .A2(n5877), .A3(n5876), .A4(n5875), .ZN(n8484)
         );
  NAND2_X1 U5728 ( .A1(n6582), .A2(n6581), .ZN(n8219) );
  AND2_X1 U5729 ( .A1(n8373), .A2(n6108), .ZN(n8569) );
  OR2_X1 U5730 ( .A1(n6521), .A2(n6520), .ZN(n6785) );
  AOI21_X1 U5731 ( .B1(n4587), .B2(n4589), .A(n4586), .ZN(n4585) );
  INV_X1 U5732 ( .A(n6560), .ZN(n4586) );
  AND2_X1 U5733 ( .A1(n6036), .A2(n6035), .ZN(n8783) );
  NAND2_X1 U5734 ( .A1(n4919), .A2(n4318), .ZN(n8247) );
  NAND2_X1 U5735 ( .A1(n8317), .A2(n4923), .ZN(n4919) );
  NAND2_X1 U5736 ( .A1(n4929), .A2(n4319), .ZN(n7295) );
  AOI21_X1 U5737 ( .B1(n8836), .B2(n6103), .A(n5996), .ZN(n8301) );
  NAND2_X1 U5738 ( .A1(n8219), .A2(n6585), .ZN(n8297) );
  NAND2_X1 U5739 ( .A1(n8268), .A2(n6578), .ZN(n8326) );
  AOI21_X1 U5740 ( .B1(n8317), .B2(n4347), .A(n4920), .ZN(n8334) );
  INV_X1 U5741 ( .A(n8341), .ZN(n8355) );
  NAND2_X1 U5742 ( .A1(n8614), .A2(n8613), .ZN(n4423) );
  INV_X1 U5743 ( .A(n8413), .ZN(n8758) );
  NAND2_X1 U5744 ( .A1(n6069), .A2(n6068), .ZN(n8775) );
  INV_X1 U5745 ( .A(n8783), .ZN(n8805) );
  INV_X1 U5746 ( .A(n8301), .ZN(n8846) );
  INV_X1 U5747 ( .A(n8892), .ZN(n8924) );
  NAND4_X1 U5748 ( .A1(n5891), .A2(n5890), .A3(n5889), .A4(n5888), .ZN(n8621)
         );
  OR2_X1 U5749 ( .A1(n6707), .A2(n10311), .ZN(n6708) );
  NAND2_X1 U5750 ( .A1(n6430), .A2(n6429), .ZN(n6794) );
  NAND2_X1 U5751 ( .A1(n4431), .A2(n4430), .ZN(n6792) );
  INV_X1 U5752 ( .A(n6795), .ZN(n4430) );
  INV_X1 U5753 ( .A(n6794), .ZN(n4431) );
  AOI21_X1 U5754 ( .B1(n6741), .B2(n8637), .A(n8638), .ZN(n8641) );
  AOI21_X1 U5755 ( .B1(n6915), .B2(n4335), .A(n6914), .ZN(n6913) );
  AOI21_X1 U5756 ( .B1(n6922), .B2(n4315), .A(n6921), .ZN(n6924) );
  INV_X1 U5757 ( .A(n4738), .ZN(n4735) );
  INV_X1 U5758 ( .A(n4730), .ZN(n7492) );
  AND2_X1 U5759 ( .A1(n4330), .A2(n4744), .ZN(n8684) );
  NAND2_X1 U5760 ( .A1(n4609), .A2(n6381), .ZN(n8651) );
  AND2_X1 U5761 ( .A1(n8682), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4743) );
  AND2_X1 U5762 ( .A1(n4607), .A2(n4606), .ZN(n8678) );
  AND2_X1 U5763 ( .A1(n8701), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4637) );
  NAND2_X1 U5764 ( .A1(n8702), .A2(n8701), .ZN(n4638) );
  AND2_X1 U5765 ( .A1(n8639), .A2(n4616), .ZN(n4614) );
  NAND2_X1 U5766 ( .A1(n8639), .A2(n4617), .ZN(n4615) );
  NAND2_X1 U5767 ( .A1(n4619), .A2(n4413), .ZN(n4617) );
  INV_X1 U5768 ( .A(n9092), .ZN(n8933) );
  NAND2_X1 U5769 ( .A1(n6986), .A2(n5771), .ZN(n7062) );
  INV_X1 U5770 ( .A(n10285), .ZN(n8208) );
  INV_X1 U5771 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8213) );
  NAND2_X1 U5772 ( .A1(n8359), .A2(n8358), .ZN(n8949) );
  NOR2_X1 U5773 ( .A1(n10323), .A2(n8953), .ZN(n4515) );
  NAND2_X1 U5774 ( .A1(n6060), .A2(n6059), .ZN(n9018) );
  NAND2_X1 U5775 ( .A1(n4886), .A2(n4889), .ZN(n8763) );
  OR2_X1 U5776 ( .A1(n6192), .A2(n4891), .ZN(n4886) );
  NAND2_X1 U5777 ( .A1(n4518), .A2(n4517), .ZN(n4516) );
  NAND2_X1 U5778 ( .A1(n8767), .A2(n10262), .ZN(n4517) );
  AOI21_X1 U5779 ( .B1(n4446), .B2(n10257), .A(n4443), .ZN(n9022) );
  NAND2_X1 U5780 ( .A1(n4445), .A2(n4444), .ZN(n4443) );
  XNOR2_X1 U5781 ( .A(n8773), .B(n4447), .ZN(n4446) );
  NAND2_X1 U5782 ( .A1(n4568), .A2(n10262), .ZN(n4444) );
  NAND2_X1 U5783 ( .A1(n4894), .A2(n8426), .ZN(n8772) );
  NAND2_X1 U5784 ( .A1(n6192), .A2(n8554), .ZN(n4894) );
  INV_X1 U5785 ( .A(n6192), .ZN(n8787) );
  NAND2_X1 U5786 ( .A1(n4458), .A2(n6026), .ZN(n8793) );
  NAND2_X1 U5787 ( .A1(n8803), .A2(n6025), .ZN(n4458) );
  NAND2_X1 U5788 ( .A1(n4903), .A2(n4902), .ZN(n8791) );
  NAND2_X1 U5789 ( .A1(n4903), .A2(n8428), .ZN(n8801) );
  NAND2_X1 U5790 ( .A1(n8862), .A2(n4908), .ZN(n8826) );
  NAND2_X1 U5791 ( .A1(n8862), .A2(n8536), .ZN(n8840) );
  NAND2_X1 U5792 ( .A1(n5923), .A2(n5922), .ZN(n9085) );
  NAND2_X1 U5793 ( .A1(n6185), .A2(n8432), .ZN(n8921) );
  NAND2_X1 U5794 ( .A1(n7639), .A2(n7636), .ZN(n4501) );
  NAND2_X1 U5795 ( .A1(n5842), .A2(n5841), .ZN(n7451) );
  INV_X1 U5796 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5714) );
  OAI21_X1 U5797 ( .B1(n6118), .B2(n4899), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5725) );
  NAND2_X1 U5798 ( .A1(n6120), .A2(n4581), .ZN(n9103) );
  AOI21_X1 U5799 ( .B1(n6118), .B2(n4583), .A(n4582), .ZN(n4581) );
  NOR2_X1 U5800 ( .A1(n6119), .A2(n5711), .ZN(n4583) );
  AND2_X1 U5801 ( .A1(n6119), .A2(n5711), .ZN(n4582) );
  INV_X1 U5802 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n9854) );
  INV_X1 U5803 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6682) );
  INV_X1 U5804 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4983) );
  CLKBUF_X1 U5805 ( .A(n6717), .Z(n4433) );
  NAND2_X1 U5806 ( .A1(n9346), .A2(n7231), .ZN(n7686) );
  AND2_X1 U5807 ( .A1(n9127), .A2(n9126), .ZN(n9197) );
  NAND2_X1 U5808 ( .A1(n4872), .A2(n4873), .ZN(n9182) );
  OR2_X1 U5809 ( .A1(n9252), .A2(n4876), .ZN(n4872) );
  INV_X1 U5810 ( .A(n7155), .ZN(n10168) );
  INV_X1 U5811 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4538) );
  INV_X1 U5812 ( .A(n10010), .ZN(n4537) );
  NOR2_X1 U5813 ( .A1(n9227), .A2(n7726), .ZN(n9300) );
  NAND2_X1 U5814 ( .A1(n9251), .A2(n7767), .ZN(n9338) );
  AND2_X1 U5815 ( .A1(n6830), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9364) );
  INV_X1 U5816 ( .A(n9364), .ZN(n9342) );
  AND2_X1 U5817 ( .A1(n6874), .A2(n6871), .ZN(n9349) );
  INV_X1 U5818 ( .A(n9366), .ZN(n9356) );
  INV_X1 U5819 ( .A(n9369), .ZN(n9332) );
  NAND2_X1 U5820 ( .A1(n5512), .A2(n5511), .ZN(n9377) );
  NAND2_X1 U5821 ( .A1(n5477), .A2(n5476), .ZN(n9379) );
  OR2_X1 U5822 ( .A1(n9576), .A2(n5552), .ZN(n5477) );
  NAND4_X2 U5823 ( .A1(n5026), .A2(n5025), .A3(n5024), .A4(n5023), .ZN(n9401)
         );
  OR2_X1 U5824 ( .A1(n5065), .A2(n5022), .ZN(n5024) );
  AND2_X1 U5825 ( .A1(n6356), .A2(n6355), .ZN(n10014) );
  NAND2_X1 U5826 ( .A1(n9449), .A2(n4369), .ZN(n9464) );
  NAND2_X1 U5827 ( .A1(n9464), .A2(n9465), .ZN(n9463) );
  AND2_X1 U5828 ( .A1(n4659), .A2(n4658), .ZN(n9457) );
  NAND2_X1 U5829 ( .A1(n7312), .A2(n4398), .ZN(n7405) );
  NOR2_X1 U5830 ( .A1(n7405), .A2(n7406), .ZN(n7404) );
  AND2_X1 U5831 ( .A1(n7616), .A2(n6347), .ZN(n10020) );
  INV_X1 U5832 ( .A(n4640), .ZN(n10021) );
  XNOR2_X1 U5833 ( .A(n6349), .B(n4450), .ZN(n10036) );
  NOR2_X1 U5834 ( .A1(n10036), .A2(n10035), .ZN(n10034) );
  NOR2_X1 U5835 ( .A1(n10050), .A2(n10049), .ZN(n10048) );
  NAND2_X1 U5836 ( .A1(n10063), .A2(n10064), .ZN(n10062) );
  NAND2_X1 U5837 ( .A1(n10043), .A2(n6325), .ZN(n10063) );
  NAND2_X1 U5838 ( .A1(n4645), .A2(n4647), .ZN(n10078) );
  INV_X1 U5839 ( .A(n6353), .ZN(n6362) );
  AOI21_X1 U5840 ( .B1(n9507), .B2(n9506), .A(n9505), .ZN(n9509) );
  INV_X1 U5841 ( .A(n8138), .ZN(n9508) );
  NAND2_X1 U5842 ( .A1(n5680), .A2(n4326), .ZN(n4546) );
  XNOR2_X1 U5843 ( .A(n5550), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9526) );
  INV_X1 U5844 ( .A(n9731), .ZN(n9598) );
  NAND2_X1 U5845 ( .A1(n9640), .A2(n8000), .ZN(n9623) );
  NAND2_X1 U5846 ( .A1(n7627), .A2(n7989), .ZN(n9700) );
  INV_X1 U5847 ( .A(n9776), .ZN(n9143) );
  NAND2_X1 U5848 ( .A1(n4814), .A2(n5621), .ZN(n7392) );
  INV_X1 U5849 ( .A(n9660), .ZN(n10143) );
  INV_X1 U5850 ( .A(n9708), .ZN(n10154) );
  AND2_X1 U5851 ( .A1(n7909), .A2(n9709), .ZN(n6249) );
  INV_X1 U5852 ( .A(n9503), .ZN(n9784) );
  OAI21_X1 U5853 ( .B1(n4422), .B2(n4316), .A(n4665), .ZN(n9586) );
  NAND2_X1 U5854 ( .A1(n4422), .A2(n9624), .ZN(n9602) );
  NAND2_X1 U5855 ( .A1(n4685), .A2(n4683), .ZN(n9637) );
  NAND2_X1 U5856 ( .A1(n4685), .A2(n5379), .ZN(n9658) );
  NAND2_X2 U5857 ( .A1(n5386), .A2(n5385), .ZN(n9822) );
  AND2_X2 U5858 ( .A1(n6246), .A2(n6826), .ZN(n10232) );
  OAI211_X1 U5859 ( .C1(n6223), .C2(n6234), .A(n6233), .B(n6232), .ZN(n8361)
         );
  MUX2_X1 U5860 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5568), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n5570) );
  INV_X1 U5861 ( .A(n5584), .ZN(n10009) );
  XNOR2_X1 U5862 ( .A(n5564), .B(n5563), .ZN(n7625) );
  NAND2_X1 U5863 ( .A1(n4782), .A2(n5446), .ZN(n5462) );
  NAND2_X1 U5864 ( .A1(n4787), .A2(n4393), .ZN(n4782) );
  NAND2_X1 U5865 ( .A1(n4484), .A2(n4336), .ZN(n5356) );
  NAND2_X1 U5866 ( .A1(n5287), .A2(n5271), .ZN(n6822) );
  NAND2_X1 U5867 ( .A1(n4774), .A2(n4772), .ZN(n5202) );
  INV_X1 U5868 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5147) );
  XNOR2_X1 U5869 ( .A(n4449), .B(n5040), .ZN(n9414) );
  NAND2_X1 U5870 ( .A1(n5363), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4449) );
  OAI21_X1 U5871 ( .B1(n5012), .B2(n4653), .A(n4652), .ZN(n4651) );
  NAND2_X1 U5872 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4653) );
  NAND2_X1 U5873 ( .A1(n4976), .A2(n4975), .ZN(n6680) );
  NAND2_X1 U5874 ( .A1(n4598), .A2(n6606), .ZN(n4596) );
  NAND2_X1 U5875 ( .A1(n4765), .A2(n6383), .ZN(n8688) );
  NOR2_X1 U5876 ( .A1(n6392), .A2(n4439), .ZN(n4438) );
  NAND2_X1 U5877 ( .A1(n6313), .A2(n10269), .ZN(n6314) );
  INV_X1 U5878 ( .A(n6312), .ZN(n6315) );
  OAI21_X1 U5879 ( .B1(n6277), .B2(n6292), .A(n6291), .ZN(n6293) );
  OAI21_X1 U5880 ( .B1(n9016), .B2(n10320), .A(n4512), .ZN(P2_U3486) );
  INV_X1 U5881 ( .A(n4513), .ZN(n4512) );
  OAI21_X1 U5882 ( .B1(n9021), .B2(n8992), .A(n4514), .ZN(n4513) );
  NOR2_X1 U5883 ( .A1(n4394), .A2(n4515), .ZN(n4514) );
  NOR2_X1 U5884 ( .A1(n10308), .A2(n6196), .ZN(n6197) );
  NAND2_X1 U5885 ( .A1(n4352), .A2(n4846), .ZN(n4844) );
  NAND2_X1 U5886 ( .A1(n5655), .A2(n9663), .ZN(n5656) );
  AND2_X1 U5887 ( .A1(n5698), .A2(n5697), .ZN(n5699) );
  NOR2_X1 U5888 ( .A1(n7850), .A2(n7849), .ZN(n7851) );
  AND2_X1 U5889 ( .A1(n9203), .A2(n9771), .ZN(n7849) );
  AOI21_X1 U5890 ( .B1(n7845), .B2(n4827), .A(n4826), .ZN(n7850) );
  OAI21_X1 U5891 ( .B1(n9510), .B2(n9812), .A(n6298), .ZN(n6299) );
  NOR2_X1 U5892 ( .A1(n7847), .A2(n7846), .ZN(n7848) );
  AND2_X1 U5893 ( .A1(n9203), .A2(n9836), .ZN(n7846) );
  AOI21_X1 U5894 ( .B1(n7845), .B2(n4829), .A(n4828), .ZN(n7847) );
  INV_X1 U5895 ( .A(n4971), .ZN(n7911) );
  INV_X1 U5896 ( .A(n6750), .ZN(n4756) );
  AND2_X1 U5897 ( .A1(n4753), .A2(n4756), .ZN(n4313) );
  NAND2_X1 U5898 ( .A1(n7732), .A2(n7731), .ZN(n4314) );
  NAND2_X1 U5899 ( .A1(n4751), .A2(n4750), .ZN(n4315) );
  NAND2_X1 U5900 ( .A1(n9601), .A2(n4949), .ZN(n4316) );
  NAND2_X1 U5901 ( .A1(n9525), .A2(n4806), .ZN(n4317) );
  INV_X1 U5902 ( .A(n4931), .ZN(n4930) );
  NAND2_X1 U5903 ( .A1(n6586), .A2(n6585), .ZN(n4931) );
  INV_X1 U5904 ( .A(n8068), .ZN(n4819) );
  AND2_X1 U5905 ( .A1(n4922), .A2(n6595), .ZN(n4318) );
  AND2_X1 U5906 ( .A1(n6548), .A2(n6547), .ZN(n4319) );
  NAND2_X1 U5907 ( .A1(n6380), .A2(n6904), .ZN(n6381) );
  AND2_X1 U5908 ( .A1(n9234), .A2(n4804), .ZN(n4320) );
  NAND2_X1 U5909 ( .A1(n4568), .A2(n4567), .ZN(n8554) );
  INV_X1 U5910 ( .A(n8554), .ZN(n4708) );
  OAI21_X1 U5911 ( .B1(n6582), .B2(n4931), .A(n4593), .ZN(n8239) );
  AND2_X1 U5912 ( .A1(n4459), .A2(n8794), .ZN(n4321) );
  AND3_X1 U5913 ( .A1(n4765), .A2(n6383), .A3(P2_REG1_REG_15__SCAN_IN), .ZN(
        n4322) );
  NOR2_X1 U5914 ( .A1(n5985), .A2(n8855), .ZN(n4323) );
  NOR2_X1 U5915 ( .A1(n6434), .A2(n10316), .ZN(n4324) );
  INV_X1 U5916 ( .A(n6683), .ZN(n7050) );
  AND2_X1 U5917 ( .A1(n9679), .A2(n5608), .ZN(n4325) );
  NAND2_X1 U5918 ( .A1(n8511), .A2(n8510), .ZN(n7583) );
  INV_X1 U5919 ( .A(n9558), .ZN(n9722) );
  NOR2_X1 U5920 ( .A1(n9611), .A2(n9731), .ZN(n5609) );
  AND2_X1 U5921 ( .A1(n4549), .A2(n4374), .ZN(n4326) );
  AND2_X1 U5922 ( .A1(n4764), .A2(n6373), .ZN(n4327) );
  AND2_X1 U5923 ( .A1(n4689), .A2(n4357), .ZN(n4328) );
  AND2_X1 U5924 ( .A1(n5627), .A2(n7989), .ZN(n4329) );
  AND2_X1 U5925 ( .A1(n6407), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4330) );
  AND2_X1 U5926 ( .A1(n6188), .A2(n8520), .ZN(n4331) );
  AND2_X1 U5927 ( .A1(n6381), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4332) );
  NAND2_X1 U5928 ( .A1(n7387), .A2(n4804), .ZN(n7463) );
  AND2_X1 U5929 ( .A1(n4576), .A2(n4575), .ZN(n4333) );
  OR2_X1 U5930 ( .A1(n7106), .A2(n10131), .ZN(n4334) );
  OR2_X1 U5931 ( .A1(n6375), .A2(n6445), .ZN(n4335) );
  OR2_X1 U5932 ( .A1(n5348), .A2(SI_17_), .ZN(n4336) );
  NOR2_X2 U5933 ( .A1(n5718), .A2(n5717), .ZN(n4337) );
  INV_X1 U5934 ( .A(n4568), .ZN(n8423) );
  NAND2_X1 U5935 ( .A1(n6045), .A2(n6044), .ZN(n4568) );
  AND2_X1 U5936 ( .A1(n6591), .A2(n8243), .ZN(n4338) );
  AND2_X1 U5937 ( .A1(n10058), .A2(n4452), .ZN(n4339) );
  CLKBUF_X3 U5938 ( .A(n5102), .Z(n5529) );
  AND2_X1 U5939 ( .A1(n8276), .A2(n8819), .ZN(n4340) );
  OAI21_X1 U5940 ( .B1(n9227), .B2(n4860), .A(n4859), .ZN(n9133) );
  AND2_X1 U5941 ( .A1(n6172), .A2(n8500), .ZN(n4341) );
  AND2_X1 U5942 ( .A1(n9525), .A2(n9529), .ZN(n4342) );
  OR2_X1 U5943 ( .A1(n8626), .A2(n8289), .ZN(n4343) );
  AND2_X1 U5944 ( .A1(n4336), .A2(n5354), .ZN(n4344) );
  NAND2_X1 U5945 ( .A1(n7262), .A2(n7261), .ZN(n4929) );
  OR2_X1 U5946 ( .A1(n8393), .A2(n7248), .ZN(n4345) );
  OR2_X1 U5947 ( .A1(n8276), .A2(n8819), .ZN(n4346) );
  AND2_X1 U5948 ( .A1(n8248), .A2(n4923), .ZN(n4347) );
  AND2_X1 U5949 ( .A1(n8064), .A2(n7988), .ZN(n4348) );
  AND2_X1 U5950 ( .A1(n4343), .A2(n5771), .ZN(n4349) );
  AND2_X1 U5951 ( .A1(n4629), .A2(n4627), .ZN(n4350) );
  OR2_X1 U5952 ( .A1(n5219), .A2(SI_11_), .ZN(n4351) );
  AND2_X1 U5953 ( .A1(n9126), .A2(n4850), .ZN(n4352) );
  NAND2_X1 U5954 ( .A1(n4501), .A2(n7637), .ZN(n8934) );
  AND3_X1 U5955 ( .A1(n9205), .A2(n9349), .A3(n9204), .ZN(n4353) );
  OR2_X1 U5956 ( .A1(n7743), .A2(n9136), .ZN(n4354) );
  NAND2_X1 U5957 ( .A1(n7070), .A2(n8111), .ZN(n7937) );
  AND2_X1 U5958 ( .A1(n9784), .A2(n8039), .ZN(n4355) );
  OR2_X1 U5959 ( .A1(n9731), .A2(n9380), .ZN(n4356) );
  INV_X1 U5960 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5798) );
  INV_X1 U5961 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4980) );
  AND3_X1 U5962 ( .A1(n8488), .A2(n8487), .A3(n8489), .ZN(n4357) );
  AND2_X1 U5963 ( .A1(n5727), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n4358) );
  AND2_X1 U5964 ( .A1(n6275), .A2(n6274), .ZN(n7914) );
  NAND2_X1 U5965 ( .A1(n4638), .A2(n4636), .ZN(n4359) );
  NOR2_X1 U5966 ( .A1(n8901), .A2(n5953), .ZN(n4360) );
  NAND2_X1 U5967 ( .A1(n4884), .A2(n8520), .ZN(n8875) );
  AND2_X1 U5968 ( .A1(n6580), .A2(n8893), .ZN(n4361) );
  AND2_X1 U5969 ( .A1(n6587), .A2(n8858), .ZN(n4362) );
  AND2_X1 U5970 ( .A1(n5859), .A2(n6096), .ZN(n6459) );
  INV_X1 U5971 ( .A(n7728), .ZN(n9307) );
  AND2_X1 U5972 ( .A1(n5251), .A2(n5250), .ZN(n7728) );
  OR2_X1 U5973 ( .A1(n9048), .A2(n8243), .ZN(n8428) );
  NAND2_X1 U5974 ( .A1(n4442), .A2(n5856), .ZN(n6096) );
  AND2_X1 U5975 ( .A1(n6543), .A2(n6542), .ZN(n4363) );
  AND2_X1 U5976 ( .A1(n4748), .A2(n6416), .ZN(n4364) );
  NAND2_X1 U5977 ( .A1(n9828), .A2(n9386), .ZN(n4365) );
  AND2_X1 U5978 ( .A1(n4837), .A2(n4839), .ZN(n4366) );
  INV_X1 U5979 ( .A(n5688), .ZN(n9510) );
  INV_X1 U5980 ( .A(n7553), .ZN(n9333) );
  NAND2_X1 U5981 ( .A1(n5194), .A2(n5193), .ZN(n7553) );
  OR2_X1 U5982 ( .A1(n9429), .A2(n6339), .ZN(n4367) );
  AND2_X1 U5983 ( .A1(n7983), .A2(n4534), .ZN(n4368) );
  NAND2_X1 U5984 ( .A1(n4348), .A2(n7980), .ZN(n4526) );
  OR2_X1 U5985 ( .A1(n6644), .A2(n7073), .ZN(n4369) );
  AND2_X1 U5986 ( .A1(n4502), .A2(n4360), .ZN(n4370) );
  INV_X1 U5987 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5011) );
  AND2_X1 U5988 ( .A1(n8219), .A2(n4930), .ZN(n4371) );
  NAND2_X1 U5989 ( .A1(n5398), .A2(n5397), .ZN(n9816) );
  INV_X1 U5990 ( .A(n9816), .ZN(n4808) );
  OR2_X1 U5991 ( .A1(n8813), .A2(n8546), .ZN(n4372) );
  NOR2_X1 U5992 ( .A1(n9036), .A2(n8805), .ZN(n4373) );
  INV_X1 U5993 ( .A(n8550), .ZN(n4904) );
  INV_X1 U5994 ( .A(n4807), .ZN(n4806) );
  NAND2_X1 U5995 ( .A1(n9529), .A2(n4303), .ZN(n4807) );
  NAND2_X1 U5996 ( .A1(n8042), .A2(n8138), .ZN(n4374) );
  INV_X1 U5997 ( .A(n10260), .ZN(n5769) );
  INV_X1 U5998 ( .A(n9822), .ZN(n4810) );
  AND2_X1 U5999 ( .A1(n7972), .A2(n8039), .ZN(n4375) );
  NAND2_X1 U6000 ( .A1(n6597), .A2(n8423), .ZN(n4376) );
  AND2_X1 U6001 ( .A1(n9822), .A2(n9384), .ZN(n4377) );
  INV_X1 U6002 ( .A(n9234), .ZN(n7515) );
  AND2_X1 U6003 ( .A1(n5229), .A2(n5228), .ZN(n9234) );
  OR2_X1 U6004 ( .A1(n9054), .A2(n8301), .ZN(n8544) );
  AND2_X1 U6005 ( .A1(n8542), .A2(n4720), .ZN(n4378) );
  NOR2_X1 U6006 ( .A1(n9715), .A2(n9376), .ZN(n4379) );
  NAND2_X1 U6007 ( .A1(n5264), .A2(n5263), .ZN(n4380) );
  NAND2_X1 U6008 ( .A1(n6190), .A2(n8555), .ZN(n4381) );
  AND2_X1 U6009 ( .A1(n4320), .A2(n7728), .ZN(n4382) );
  AND2_X1 U6010 ( .A1(n6660), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4383) );
  INV_X1 U6011 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5290) );
  INV_X1 U6012 ( .A(n4969), .ZN(n9999) );
  AND2_X1 U6013 ( .A1(n8076), .A2(n7925), .ZN(n4384) );
  INV_X1 U6014 ( .A(n7989), .ZN(n4553) );
  AND2_X1 U6015 ( .A1(n8553), .A2(n4900), .ZN(n4385) );
  INV_X1 U6016 ( .A(n6566), .ZN(n4927) );
  AND2_X1 U6017 ( .A1(n4524), .A2(n4528), .ZN(n4386) );
  NAND2_X1 U6018 ( .A1(n4346), .A2(n8280), .ZN(n4387) );
  INV_X1 U6019 ( .A(n8526), .ZN(n4896) );
  AND2_X1 U6020 ( .A1(n8590), .A2(n8594), .ZN(n4388) );
  AND2_X1 U6021 ( .A1(n4473), .A2(n6070), .ZN(n4389) );
  AND2_X1 U6022 ( .A1(n4862), .A2(n7702), .ZN(n4390) );
  INV_X1 U6023 ( .A(n4634), .ZN(n4633) );
  NOR2_X1 U6024 ( .A1(n6920), .A2(n7335), .ZN(n4634) );
  AND2_X1 U6025 ( .A1(n4847), .A2(n4848), .ZN(n4391) );
  OR2_X1 U6026 ( .A1(n9060), .A2(n8858), .ZN(n8543) );
  AND2_X1 U6027 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_REG3_REG_6__SCAN_IN), 
        .ZN(n4392) );
  XNOR2_X1 U6028 ( .A(n5822), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6445) );
  INV_X1 U6029 ( .A(n6445), .ZN(n4750) );
  AND2_X1 U6030 ( .A1(n7387), .A2(n7421), .ZN(n7388) );
  NAND2_X1 U6031 ( .A1(n5766), .A2(n5789), .ZN(n6647) );
  AND2_X1 U6032 ( .A1(n5429), .A2(n4786), .ZN(n4393) );
  AND2_X1 U6033 ( .A1(n9018), .A2(n8994), .ZN(n4394) );
  NAND2_X1 U6034 ( .A1(n6038), .A2(n6037), .ZN(n9030) );
  INV_X1 U6035 ( .A(n9030), .ZN(n4567) );
  NAND2_X1 U6036 ( .A1(n7670), .A2(n4325), .ZN(n9664) );
  AND2_X1 U6037 ( .A1(n7780), .A2(n7779), .ZN(n4395) );
  NAND2_X1 U6038 ( .A1(n4928), .A2(n6564), .ZN(n8305) );
  NAND2_X1 U6039 ( .A1(n4929), .A2(n6547), .ZN(n7293) );
  AND2_X1 U6040 ( .A1(n6407), .A2(n4744), .ZN(n4396) );
  INV_X1 U6041 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n4494) );
  NOR2_X1 U6042 ( .A1(n9300), .A2(n9301), .ZN(n4397) );
  OR2_X1 U6043 ( .A1(n6700), .A2(n7462), .ZN(n4398) );
  NAND2_X1 U6044 ( .A1(n4735), .A2(n4730), .ZN(n4399) );
  NAND2_X1 U6045 ( .A1(n4742), .A2(n4741), .ZN(n4400) );
  AND2_X1 U6046 ( .A1(n4836), .A2(n4837), .ZN(n4401) );
  INV_X1 U6047 ( .A(n9378), .ZN(n7684) );
  NAND2_X1 U6048 ( .A1(n5497), .A2(n5496), .ZN(n9378) );
  AND2_X1 U6049 ( .A1(n6376), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4402) );
  AND2_X1 U6050 ( .A1(n4495), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n4403) );
  NAND2_X1 U6051 ( .A1(n6255), .A2(n8566), .ZN(n7918) );
  AND2_X1 U6052 ( .A1(n4573), .A2(n4572), .ZN(n4404) );
  NOR2_X1 U6053 ( .A1(n10192), .A2(n10131), .ZN(n4802) );
  INV_X1 U6054 ( .A(n10039), .ZN(n4450) );
  AND2_X1 U6055 ( .A1(n10026), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4405) );
  NAND2_X1 U6056 ( .A1(n6742), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6741) );
  OR2_X1 U6057 ( .A1(n6821), .A2(n6408), .ZN(n4406) );
  OR2_X1 U6058 ( .A1(n7236), .A2(n7235), .ZN(n4407) );
  XOR2_X1 U6059 ( .A(n8739), .B(n8977), .Z(n4408) );
  OR2_X1 U6060 ( .A1(n6821), .A2(n8993), .ZN(n4409) );
  OR2_X1 U6061 ( .A1(n6994), .A2(n6411), .ZN(n4410) );
  OR2_X1 U6062 ( .A1(n6994), .A2(n6384), .ZN(n4411) );
  AND2_X1 U6063 ( .A1(n4647), .A2(n4649), .ZN(n4412) );
  INV_X1 U6064 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n4496) );
  INV_X1 U6065 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n4497) );
  OR2_X1 U6066 ( .A1(n4408), .A2(n4622), .ZN(n4413) );
  NOR2_X1 U6067 ( .A1(n10057), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n4414) );
  NAND2_X1 U6068 ( .A1(n4408), .A2(n6386), .ZN(n4618) );
  NAND2_X1 U6069 ( .A1(n7164), .A2(n6376), .ZN(n4415) );
  AND2_X1 U6070 ( .A1(n4498), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n4416) );
  NAND2_X1 U6071 ( .A1(n4619), .A2(n4618), .ZN(n4616) );
  XNOR2_X1 U6072 ( .A(n5870), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7367) );
  INV_X1 U6073 ( .A(n7367), .ZN(n4769) );
  AND2_X1 U6074 ( .A1(n4763), .A2(n6724), .ZN(n4417) );
  INV_X1 U6075 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n4737) );
  INV_X1 U6076 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4490) );
  INV_X1 U6077 ( .A(n4650), .ZN(n6940) );
  OR2_X1 U6078 ( .A1(n5013), .A2(n4651), .ZN(n4650) );
  INV_X1 U6079 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n4761) );
  NAND2_X1 U6080 ( .A1(n4738), .A2(n4736), .ZN(n4734) );
  INV_X1 U6081 ( .A(n6169), .ZN(n8387) );
  NAND2_X1 U6082 ( .A1(n7034), .A2(n6521), .ZN(n7035) );
  AND2_X2 U6083 ( .A1(n8446), .A2(n8447), .ZN(n7034) );
  NAND2_X1 U6084 ( .A1(n8943), .A2(n8431), .ZN(n6185) );
  NAND2_X1 U6085 ( .A1(n6192), .A2(n4889), .ZN(n4885) );
  INV_X2 U6086 ( .A(n7044), .ZN(n6522) );
  NAND3_X2 U6087 ( .A1(n5736), .A2(n5737), .A3(n5738), .ZN(n7044) );
  NAND3_X1 U6088 ( .A1(n4305), .A2(n4821), .A3(n4831), .ZN(n4967) );
  NAND2_X1 U6089 ( .A1(n7156), .A2(n5613), .ZN(n10138) );
  INV_X1 U6090 ( .A(n8041), .ZN(n8179) );
  NAND2_X1 U6091 ( .A1(n4535), .A2(n4531), .ZN(n4429) );
  OAI21_X1 U6092 ( .B1(n8018), .B2(n8017), .A(n8016), .ZN(n8019) );
  OAI21_X1 U6093 ( .B1(n7946), .B2(n7945), .A(n8168), .ZN(n4544) );
  NAND2_X1 U6094 ( .A1(n4419), .A2(n4418), .ZN(P1_U3549) );
  MUX2_X1 U6095 ( .A(n9716), .B(n9785), .S(n10248), .Z(n4419) );
  NAND2_X1 U6096 ( .A1(n4558), .A2(n8083), .ZN(n4557) );
  NAND2_X1 U6097 ( .A1(n5381), .A2(n5380), .ZN(n5396) );
  OAI21_X2 U6098 ( .B1(n8860), .B2(n4907), .A(n4905), .ZN(n4420) );
  AND2_X2 U6099 ( .A1(n6191), .A2(n8555), .ZN(n6192) );
  NAND3_X1 U6100 ( .A1(n5677), .A2(n5679), .A3(n5678), .ZN(n4421) );
  NAND2_X1 U6101 ( .A1(n5064), .A2(n5063), .ZN(n7068) );
  OAI21_X4 U6102 ( .B1(n9572), .B2(n5479), .A(n5478), .ZN(n9549) );
  OAI21_X1 U6103 ( .B1(n4304), .B2(n4983), .A(n4982), .ZN(n4984) );
  NAND2_X1 U6104 ( .A1(n4688), .A2(n4800), .ZN(n4687) );
  NAND2_X1 U6105 ( .A1(n5005), .A2(n4455), .ZN(n5010) );
  NAND2_X1 U6106 ( .A1(n4732), .A2(n4734), .ZN(n7495) );
  INV_X1 U6107 ( .A(n6393), .ZN(n4580) );
  NAND3_X1 U6108 ( .A1(n8589), .A2(n4436), .A3(n4388), .ZN(n8597) );
  NAND4_X1 U6109 ( .A1(n4705), .A2(n8556), .A3(n4564), .A4(n8774), .ZN(n8560)
         );
  NAND2_X1 U6110 ( .A1(n4701), .A2(n8523), .ZN(n8531) );
  NAND2_X1 U6111 ( .A1(n4435), .A2(n8515), .ZN(n8527) );
  INV_X1 U6112 ( .A(n4692), .ZN(n4691) );
  NAND2_X1 U6113 ( .A1(n7223), .A2(n7224), .ZN(n9347) );
  NAND2_X2 U6114 ( .A1(n9172), .A2(n9173), .ZN(n6968) );
  NAND2_X2 U6115 ( .A1(n7824), .A2(n7823), .ZN(n7868) );
  NAND2_X1 U6116 ( .A1(n6374), .A2(n6723), .ZN(n6727) );
  INV_X1 U6117 ( .A(n7168), .ZN(n4612) );
  NOR2_X4 U6118 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6393) );
  CLKBUF_X2 U6119 ( .A(n6372), .Z(n4448) );
  NAND2_X1 U6120 ( .A1(n7051), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7182) );
  NAND2_X2 U6121 ( .A1(n6798), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6797) );
  AND2_X2 U6122 ( .A1(n4739), .A2(n6719), .ZN(n6798) );
  NAND2_X1 U6123 ( .A1(n8738), .A2(n8737), .ZN(n4726) );
  NAND2_X4 U6124 ( .A1(n5014), .A2(n6641), .ZN(n6218) );
  OAI21_X1 U6125 ( .B1(n9790), .B2(n9838), .A(n4425), .ZN(P1_U3516) );
  OAI21_X1 U6126 ( .B1(n9790), .B2(n9773), .A(n4427), .ZN(P1_U3548) );
  NAND2_X1 U6127 ( .A1(n4429), .A2(n4532), .ZN(n4533) );
  NAND3_X1 U6128 ( .A1(n5028), .A2(n5029), .A3(n5027), .ZN(n5033) );
  NAND2_X1 U6129 ( .A1(n4986), .A2(n4985), .ZN(n5028) );
  NAND2_X1 U6130 ( .A1(n7925), .A2(n7924), .ZN(n8109) );
  NAND2_X1 U6131 ( .A1(n6457), .A2(n6456), .ZN(n7176) );
  NAND2_X1 U6132 ( .A1(n6448), .A2(n6884), .ZN(n6910) );
  INV_X1 U6133 ( .A(n4723), .ZN(n4722) );
  OAI21_X1 U6134 ( .B1(n8179), .B2(n8178), .A(n8177), .ZN(n8180) );
  AOI21_X1 U6135 ( .B1(n8724), .B2(n8723), .A(n6488), .ZN(n6489) );
  NOR2_X1 U6136 ( .A1(n7935), .A2(n7934), .ZN(n8001) );
  NAND2_X1 U6137 ( .A1(n4540), .A2(n4539), .ZN(n8041) );
  NAND2_X2 U6138 ( .A1(n4740), .A2(n4744), .ZN(n4742) );
  NOR2_X1 U6139 ( .A1(n7179), .A2(n4432), .ZN(n6404) );
  NOR2_X1 U6140 ( .A1(n8433), .A2(n8526), .ZN(n4895) );
  AOI21_X1 U6141 ( .B1(n4889), .B2(n4891), .A(n4888), .ZN(n4887) );
  NAND3_X1 U6142 ( .A1(n7134), .A2(n4341), .A3(n6175), .ZN(n4881) );
  NAND2_X1 U6143 ( .A1(n7089), .A2(n8464), .ZN(n7134) );
  OAI21_X2 U6144 ( .B1(n7379), .B2(n8476), .A(n8504), .ZN(n7561) );
  NAND2_X1 U6145 ( .A1(n8874), .A2(n8532), .ZN(n8860) );
  NAND2_X1 U6146 ( .A1(n6254), .A2(n6253), .ZN(n8378) );
  NAND2_X1 U6147 ( .A1(n6982), .A2(n8387), .ZN(n6981) );
  NAND4_X1 U6148 ( .A1(n4434), .A2(n5856), .A3(n5708), .A4(n4710), .ZN(n6120)
         );
  AND2_X1 U6149 ( .A1(n5728), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5729) );
  NAND2_X1 U6150 ( .A1(n8514), .A2(n8944), .ZN(n4435) );
  NOR2_X2 U6151 ( .A1(n6082), .A2(n5855), .ZN(n5709) );
  NAND2_X1 U6152 ( .A1(n8588), .A2(n8587), .ZN(n4436) );
  NAND2_X1 U6153 ( .A1(n4704), .A2(n4702), .ZN(n4701) );
  NAND2_X1 U6154 ( .A1(n4712), .A2(n8534), .ZN(n4716) );
  OAI21_X1 U6155 ( .B1(n4543), .B2(n4793), .A(n4792), .ZN(n4539) );
  OAI21_X1 U6156 ( .B1(n4543), .B2(n9503), .A(n4541), .ZN(n4540) );
  NAND2_X1 U6157 ( .A1(n8019), .A2(n4798), .ZN(n4797) );
  NOR2_X1 U6158 ( .A1(n5179), .A2(SI_9_), .ZN(n5180) );
  NAND2_X1 U6159 ( .A1(n7653), .A2(n4329), .ZN(n4551) );
  NAND2_X1 U6160 ( .A1(n6868), .A2(n6867), .ZN(n6955) );
  NAND2_X1 U6161 ( .A1(n6857), .A2(n6856), .ZN(n6866) );
  NAND3_X1 U6162 ( .A1(n6506), .A2(n6504), .A3(n4438), .ZN(P2_U3200) );
  NAND2_X1 U6163 ( .A1(n4440), .A2(n6525), .ZN(n6807) );
  NAND2_X1 U6164 ( .A1(n6784), .A2(n6785), .ZN(n4440) );
  NAND2_X1 U6165 ( .A1(n4578), .A2(n6569), .ZN(n8255) );
  NAND2_X1 U6166 ( .A1(n4910), .A2(n4909), .ZN(n8217) );
  AOI21_X2 U6167 ( .B1(n8317), .B2(n8318), .A(n4338), .ZN(n8277) );
  XNOR2_X2 U6168 ( .A(n8378), .B(n6271), .ZN(n7919) );
  NAND2_X1 U6169 ( .A1(n8886), .A2(n8519), .ZN(n4884) );
  NAND2_X1 U6170 ( .A1(n6397), .A2(n6647), .ZN(n6719) );
  NOR2_X1 U6171 ( .A1(n4728), .A2(n6683), .ZN(n4727) );
  NOR2_X2 U6172 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4974) );
  INV_X1 U6173 ( .A(n5030), .ZN(n4455) );
  NAND2_X1 U6174 ( .A1(n8802), .A2(n4321), .ZN(n4456) );
  NAND2_X1 U6175 ( .A1(n4456), .A2(n4457), .ZN(n8779) );
  NAND2_X1 U6176 ( .A1(n4774), .A2(n4462), .ZN(n5204) );
  NAND3_X1 U6177 ( .A1(n4464), .A2(n4463), .A3(n8813), .ZN(n8817) );
  NAND3_X1 U6178 ( .A1(n4468), .A2(n4466), .A3(n4465), .ZN(n4464) );
  NAND2_X1 U6179 ( .A1(n4879), .A2(n6046), .ZN(n8773) );
  XNOR2_X1 U6180 ( .A(n6256), .B(n6081), .ZN(n6113) );
  NAND2_X1 U6181 ( .A1(n5350), .A2(n5349), .ZN(n4484) );
  NAND2_X1 U6182 ( .A1(n5350), .A2(n4478), .ZN(n4477) );
  INV_X1 U6183 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4489) );
  INV_X1 U6184 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4488) );
  NAND3_X1 U6185 ( .A1(n4486), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4485) );
  NAND3_X1 U6186 ( .A1(n4490), .A2(n4489), .A3(n4488), .ZN(n4487) );
  NAND2_X1 U6187 ( .A1(n4491), .A2(n4392), .ZN(n5133) );
  NAND2_X1 U6188 ( .A1(n5195), .A2(n4492), .ZN(n5277) );
  NAND2_X1 U6189 ( .A1(n5316), .A2(n4403), .ZN(n5387) );
  NAND2_X1 U6190 ( .A1(n5437), .A2(n4498), .ZN(n5471) );
  NAND2_X1 U6191 ( .A1(n5437), .A2(n4416), .ZN(n5490) );
  NAND2_X1 U6192 ( .A1(n5437), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5454) );
  OR2_X2 U6193 ( .A1(n7639), .A2(n4506), .ZN(n4500) );
  NAND2_X1 U6194 ( .A1(n4511), .A2(n4509), .ZN(n4508) );
  NAND2_X1 U6195 ( .A1(n4349), .A2(n6986), .ZN(n4511) );
  NAND2_X1 U6196 ( .A1(n4508), .A2(n7091), .ZN(n7137) );
  NAND2_X1 U6197 ( .A1(n6120), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5726) );
  NAND2_X1 U6198 ( .A1(n7967), .A2(n4528), .ZN(n4527) );
  NAND2_X1 U6199 ( .A1(n7967), .A2(n4386), .ZN(n4522) );
  NAND3_X1 U6200 ( .A1(n4527), .A2(n7981), .A3(n7980), .ZN(n7987) );
  INV_X1 U6201 ( .A(n8005), .ZN(n4532) );
  NAND3_X1 U6202 ( .A1(n4530), .A2(n7999), .A3(n4529), .ZN(n4531) );
  NAND2_X1 U6203 ( .A1(n4533), .A2(n8004), .ZN(n8007) );
  AND2_X1 U6204 ( .A1(n8001), .A2(n4536), .ZN(n4535) );
  AND2_X1 U6205 ( .A1(n8000), .A2(n9622), .ZN(n4536) );
  INV_X1 U6206 ( .A(n6901), .ZN(n7151) );
  MUX2_X1 U6207 ( .A(n4538), .B(n4537), .S(n5014), .Z(n6901) );
  XNOR2_X2 U6208 ( .A(n4981), .B(n4980), .ZN(n10002) );
  XNOR2_X2 U6209 ( .A(n4979), .B(n4978), .ZN(n8189) );
  OR2_X1 U6210 ( .A1(n5680), .A2(n4548), .ZN(n4547) );
  NAND3_X1 U6211 ( .A1(n4547), .A2(n4546), .A3(n5687), .ZN(n9516) );
  NAND3_X2 U6212 ( .A1(n4551), .A2(n4552), .A3(n9701), .ZN(n9699) );
  NAND2_X1 U6213 ( .A1(n7653), .A2(n5627), .ZN(n4555) );
  OAI21_X2 U6214 ( .B1(n9653), .B2(n4559), .A(n4556), .ZN(n8143) );
  MUX2_X1 U6215 ( .A(n6643), .B(n5751), .S(n5073), .Z(n5007) );
  MUX2_X1 U6216 ( .A(n7574), .B(n7579), .S(n6641), .Z(n5449) );
  NAND3_X1 U6217 ( .A1(n5621), .A2(n8120), .A3(n4814), .ZN(n7390) );
  NAND2_X1 U6218 ( .A1(n6029), .A2(n9846), .ZN(n6039) );
  NAND2_X1 U6219 ( .A1(n6040), .A2(n6049), .ZN(n8785) );
  NAND3_X1 U6220 ( .A1(n8213), .A2(n5782), .A3(n4565), .ZN(n5803) );
  NOR2_X1 U6221 ( .A1(n8786), .A2(n8549), .ZN(n4566) );
  NAND2_X1 U6222 ( .A1(n5901), .A2(n4404), .ZN(n5934) );
  NAND2_X1 U6223 ( .A1(n5944), .A2(n4576), .ZN(n5979) );
  NAND2_X1 U6224 ( .A1(n8255), .A2(n6570), .ZN(n6575) );
  NAND2_X1 U6225 ( .A1(n4579), .A2(n4925), .ZN(n4578) );
  NAND2_X1 U6226 ( .A1(n8307), .A2(n6566), .ZN(n4579) );
  NAND2_X1 U6227 ( .A1(n4580), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5748) );
  INV_X2 U6228 ( .A(n6526), .ZN(n6600) );
  NAND2_X1 U6229 ( .A1(n4929), .A2(n4587), .ZN(n4584) );
  NAND2_X1 U6230 ( .A1(n4584), .A2(n4585), .ZN(n7882) );
  NAND2_X1 U6231 ( .A1(n4590), .A2(n4591), .ZN(n6590) );
  NAND2_X1 U6232 ( .A1(n6582), .A2(n4593), .ZN(n4590) );
  NAND2_X1 U6233 ( .A1(n8277), .A2(n4595), .ZN(n4594) );
  OAI211_X1 U6234 ( .C1(n8277), .C2(n4596), .A(n4594), .B(n8284), .ZN(P2_U3169) );
  XNOR2_X1 U6235 ( .A(n8277), .B(n8276), .ZN(n8278) );
  INV_X1 U6236 ( .A(n8280), .ZN(n4604) );
  NAND3_X1 U6237 ( .A1(n4609), .A2(n6381), .A3(n4608), .ZN(n4607) );
  NAND2_X1 U6238 ( .A1(n8675), .A2(n8674), .ZN(n4606) );
  NAND3_X1 U6239 ( .A1(n4607), .A2(n4409), .A3(n4606), .ZN(n6382) );
  NAND2_X1 U6240 ( .A1(n6387), .A2(n6386), .ZN(n8736) );
  NAND2_X1 U6241 ( .A1(n6387), .A2(n4614), .ZN(n4613) );
  OAI211_X1 U6242 ( .C1(n6387), .C2(n4615), .A(n8755), .B(n4613), .ZN(n4723)
         );
  NAND2_X1 U6243 ( .A1(n6888), .A2(n4628), .ZN(n4627) );
  OAI211_X1 U6244 ( .C1(n4335), .C2(n4626), .A(n4625), .B(n4624), .ZN(n6377)
         );
  NAND2_X1 U6245 ( .A1(n4634), .A2(n6683), .ZN(n4624) );
  NAND2_X1 U6246 ( .A1(n6888), .A2(n4630), .ZN(n4625) );
  INV_X1 U6247 ( .A(n6914), .ZN(n4635) );
  NAND3_X1 U6248 ( .A1(n4765), .A2(n4637), .A3(n6383), .ZN(n4636) );
  INV_X1 U6249 ( .A(n10077), .ZN(n4649) );
  MUX2_X1 U6250 ( .A(n10235), .B(P1_REG1_REG_2__SCAN_IN), .S(n4650), .Z(n6939)
         );
  NAND2_X1 U6251 ( .A1(n9444), .A2(n4658), .ZN(n4655) );
  INV_X1 U6252 ( .A(n4659), .ZN(n9442) );
  INV_X1 U6253 ( .A(n4657), .ZN(n9455) );
  NAND2_X2 U6254 ( .A1(n4663), .A2(n4660), .ZN(n9572) );
  OAI21_X1 U6255 ( .B1(n9549), .B2(n5498), .A(n4677), .ZN(n9538) );
  NAND2_X1 U6256 ( .A1(n9549), .A2(n4671), .ZN(n4670) );
  OAI21_X2 U6257 ( .B1(n9538), .B2(n5514), .A(n5513), .ZN(n9520) );
  NAND2_X1 U6258 ( .A1(n9672), .A2(n4683), .ZN(n4678) );
  NAND2_X1 U6259 ( .A1(n4678), .A2(n4679), .ZN(n5409) );
  INV_X2 U6260 ( .A(n5014), .ZN(n6236) );
  AOI21_X2 U6261 ( .B1(n4687), .B2(n5014), .A(n4686), .ZN(n5614) );
  NAND2_X1 U6262 ( .A1(n8473), .A2(n4694), .ZN(n4689) );
  NAND2_X1 U6263 ( .A1(n8512), .A2(n8513), .ZN(n4692) );
  INV_X1 U6264 ( .A(n8506), .ZN(n4694) );
  NAND3_X1 U6265 ( .A1(n4697), .A2(n8449), .A3(n4695), .ZN(n8456) );
  NAND3_X1 U6266 ( .A1(n4699), .A2(n8446), .A3(n4698), .ZN(n4697) );
  NAND3_X1 U6267 ( .A1(n8517), .A2(n8591), .A3(n8518), .ZN(n4704) );
  OAI21_X1 U6268 ( .B1(n8552), .B2(n4709), .A(n4706), .ZN(n4705) );
  AND2_X2 U6269 ( .A1(n6085), .A2(n4752), .ZN(n4710) );
  INV_X1 U6270 ( .A(n4711), .ZN(n4717) );
  OAI21_X1 U6271 ( .B1(n8540), .B2(n4718), .A(n8544), .ZN(n4711) );
  INV_X1 U6272 ( .A(n8547), .ZN(n4719) );
  INV_X1 U6273 ( .A(n8535), .ZN(n4721) );
  AOI21_X2 U6274 ( .B1(n10113), .B2(n5112), .A(n4938), .ZN(n7317) );
  NAND2_X1 U6275 ( .A1(n5325), .A2(n5324), .ZN(n7666) );
  NOR2_X1 U6276 ( .A1(n6324), .A2(n10031), .ZN(n10045) );
  NAND2_X1 U6277 ( .A1(n6363), .A2(n8175), .ZN(n6364) );
  NAND2_X1 U6278 ( .A1(n4724), .A2(n4722), .ZN(P2_U3201) );
  NAND2_X1 U6279 ( .A1(n4725), .A2(n8740), .ZN(n4724) );
  XNOR2_X1 U6280 ( .A(n4726), .B(n8745), .ZN(n4725) );
  NOR2_X2 U6281 ( .A1(n6403), .A2(n4727), .ZN(n7051) );
  AND2_X2 U6282 ( .A1(n4728), .A2(n6683), .ZN(n6403) );
  CLKBUF_X1 U6283 ( .A(n4736), .Z(n4730) );
  AOI21_X2 U6284 ( .B1(n4736), .B2(n4737), .A(n4733), .ZN(n4732) );
  OR2_X2 U6285 ( .A1(n6404), .A2(n7367), .ZN(n4736) );
  AND2_X2 U6286 ( .A1(n6404), .A2(n7367), .ZN(n4738) );
  NAND2_X1 U6287 ( .A1(n8683), .A2(n8682), .ZN(n4741) );
  AND2_X2 U6288 ( .A1(n6407), .A2(n4743), .ZN(n4740) );
  NAND3_X1 U6289 ( .A1(n4742), .A2(n4406), .A3(n4741), .ZN(n6409) );
  INV_X1 U6290 ( .A(n6406), .ZN(n4745) );
  NAND2_X1 U6291 ( .A1(n4747), .A2(n6416), .ZN(n6414) );
  INV_X1 U6292 ( .A(n5765), .ZN(n5856) );
  INV_X1 U6293 ( .A(n6765), .ZN(n4757) );
  OAI22_X1 U6294 ( .A1(n4758), .A2(n4757), .B1(n4761), .B2(n6647), .ZN(n4760)
         );
  NAND2_X1 U6295 ( .A1(n4759), .A2(n6647), .ZN(n6724) );
  NAND2_X1 U6296 ( .A1(n6765), .A2(n6373), .ZN(n4759) );
  NAND2_X1 U6297 ( .A1(n4327), .A2(n6765), .ZN(n4763) );
  INV_X1 U6298 ( .A(n6373), .ZN(n4762) );
  INV_X1 U6299 ( .A(n6647), .ZN(n4764) );
  NAND2_X1 U6300 ( .A1(n6376), .A2(n4768), .ZN(n4767) );
  OAI21_X1 U6301 ( .B1(n7164), .B2(n7165), .A(n4767), .ZN(n7168) );
  NOR2_X1 U6302 ( .A1(n7165), .A2(n7469), .ZN(n4768) );
  NAND3_X1 U6303 ( .A1(n5142), .A2(n4775), .A3(n5181), .ZN(n4774) );
  NAND2_X2 U6304 ( .A1(n5127), .A2(n5126), .ZN(n5142) );
  OR2_X1 U6305 ( .A1(n5430), .A2(n4937), .ZN(n4787) );
  NAND2_X1 U6306 ( .A1(n4788), .A2(n4789), .ZN(n5270) );
  NAND2_X1 U6307 ( .A1(n5221), .A2(n4790), .ZN(n4788) );
  NAND2_X1 U6308 ( .A1(n9503), .A2(n9373), .ZN(n4793) );
  NAND2_X1 U6309 ( .A1(n4794), .A2(n8028), .ZN(n8034) );
  NAND2_X1 U6310 ( .A1(n4795), .A2(n8039), .ZN(n4794) );
  NAND2_X1 U6311 ( .A1(n4796), .A2(n8026), .ZN(n4795) );
  NAND3_X1 U6312 ( .A1(n8024), .A2(n8080), .A3(n4797), .ZN(n4796) );
  INV_X1 U6313 ( .A(n8089), .ZN(n4798) );
  NAND2_X1 U6314 ( .A1(n4799), .A2(SI_3_), .ZN(n5076) );
  MUX2_X1 U6315 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n5073), .Z(n4799) );
  NAND3_X1 U6316 ( .A1(n4802), .A2(n4803), .A3(n4801), .ZN(n7318) );
  INV_X1 U6317 ( .A(n7106), .ZN(n4803) );
  NAND3_X1 U6318 ( .A1(n9525), .A2(n9510), .A3(n4806), .ZN(n9497) );
  NAND3_X1 U6319 ( .A1(n9525), .A2(n9510), .A3(n4805), .ZN(n9498) );
  NAND2_X1 U6320 ( .A1(n4809), .A2(n7670), .ZN(n9665) );
  NAND3_X1 U6321 ( .A1(n4305), .A2(n4963), .A3(n4831), .ZN(n5569) );
  NOR2_X1 U6322 ( .A1(n8123), .A2(n8115), .ZN(n4815) );
  NAND2_X1 U6323 ( .A1(n4817), .A2(n8021), .ZN(n9521) );
  NOR2_X1 U6324 ( .A1(n4820), .A2(n5272), .ZN(n4977) );
  NAND3_X1 U6325 ( .A1(n4831), .A2(n4963), .A3(n4980), .ZN(n4820) );
  AND2_X1 U6326 ( .A1(n7844), .A2(n10232), .ZN(n4829) );
  NAND3_X1 U6327 ( .A1(n4970), .A2(n4972), .A3(n4830), .ZN(n6833) );
  INV_X1 U6328 ( .A(n4959), .ZN(n4831) );
  NOR2_X2 U6329 ( .A1(n5272), .A2(n4959), .ZN(n5559) );
  NOR2_X1 U6330 ( .A1(n4971), .A2(n4969), .ZN(n5021) );
  NOR2_X2 U6331 ( .A1(n4971), .A2(n9999), .ZN(n5046) );
  NAND2_X1 U6332 ( .A1(n8817), .A2(n6015), .ZN(n8802) );
  NAND2_X1 U6333 ( .A1(n6968), .A2(n6967), .ZN(n7122) );
  INV_X1 U6334 ( .A(n7120), .ZN(n4840) );
  INV_X1 U6335 ( .A(n7868), .ZN(n4843) );
  NAND2_X1 U6336 ( .A1(n7868), .A2(n7867), .ZN(n9127) );
  NAND4_X1 U6337 ( .A1(n4842), .A2(n4844), .A3(n4391), .A4(n4841), .ZN(
        P1_U3220) );
  NAND2_X1 U6338 ( .A1(n7868), .A2(n4845), .ZN(n4841) );
  NAND2_X1 U6339 ( .A1(n4843), .A2(n4352), .ZN(n4842) );
  NAND2_X1 U6340 ( .A1(n4854), .A2(n4855), .ZN(n7759) );
  NAND3_X1 U6341 ( .A1(n9227), .A2(n4354), .A3(n4859), .ZN(n4854) );
  NAND2_X1 U6342 ( .A1(n9346), .A2(n4864), .ZN(n4861) );
  NAND2_X1 U6343 ( .A1(n4861), .A2(n4390), .ZN(n9159) );
  NAND2_X1 U6344 ( .A1(n9252), .A2(n4870), .ZN(n4868) );
  NAND2_X1 U6345 ( .A1(n4868), .A2(n4869), .ZN(n9292) );
  OAI21_X2 U6346 ( .B1(n7245), .B2(n4345), .A(n5833), .ZN(n7344) );
  NAND2_X1 U6347 ( .A1(n5770), .A2(n6169), .ZN(n6986) );
  AND2_X2 U6348 ( .A1(n4881), .A2(n4880), .ZN(n7342) );
  NAND3_X1 U6349 ( .A1(n6173), .A2(n8500), .A3(n6175), .ZN(n4880) );
  NAND2_X1 U6350 ( .A1(n4882), .A2(n4883), .ZN(n7343) );
  NAND2_X1 U6351 ( .A1(n4341), .A2(n7251), .ZN(n4882) );
  NAND2_X1 U6352 ( .A1(n4885), .A2(n4887), .ZN(n6193) );
  NAND2_X1 U6353 ( .A1(n6185), .A2(n4895), .ZN(n6186) );
  NAND2_X1 U6354 ( .A1(n4898), .A2(n4897), .ZN(n5713) );
  INV_X1 U6355 ( .A(n6118), .ZN(n4898) );
  NOR2_X2 U6356 ( .A1(n5713), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n7900) );
  NAND2_X1 U6357 ( .A1(n6576), .A2(n4911), .ZN(n4910) );
  NAND2_X1 U6358 ( .A1(n8317), .A2(n4917), .ZN(n4916) );
  INV_X1 U6359 ( .A(n8307), .ZN(n4928) );
  NAND2_X1 U6360 ( .A1(n6203), .A2(n6202), .ZN(n6210) );
  OR3_X1 U6361 ( .A1(n6203), .A2(n6208), .A3(n5665), .ZN(n5666) );
  XNOR2_X1 U6362 ( .A(n6203), .B(n6202), .ZN(n8186) );
  INV_X1 U6363 ( .A(n7845), .ZN(n5655) );
  NOR2_X1 U6364 ( .A1(n8841), .A2(n8839), .ZN(n8842) );
  NAND2_X1 U6365 ( .A1(n5747), .A2(n6639), .ZN(n5750) );
  OAI211_X1 U6366 ( .C1(n5746), .C2(n5751), .A(n5750), .B(n5749), .ZN(n5754)
         );
  INV_X1 U6367 ( .A(n5717), .ZN(n5716) );
  XNOR2_X1 U6368 ( .A(n9507), .B(n8139), .ZN(n7852) );
  INV_X1 U6369 ( .A(n5037), .ZN(n5034) );
  NAND2_X1 U6370 ( .A1(n5265), .A2(n5264), .ZN(n5244) );
  INV_X1 U6371 ( .A(n7840), .ZN(n6176) );
  AOI21_X1 U6372 ( .B1(n6359), .B2(n8151), .A(n6358), .ZN(n6365) );
  AND2_X1 U6373 ( .A1(n7334), .A2(n8151), .ZN(n8106) );
  NAND2_X1 U6374 ( .A1(n7035), .A2(n8446), .ZN(n10250) );
  AND2_X2 U6375 ( .A1(n4971), .A2(n9999), .ZN(n5047) );
  INV_X1 U6376 ( .A(n9525), .ZN(n9542) );
  CLKBUF_X1 U6377 ( .A(n7561), .Z(n7644) );
  NAND2_X1 U6378 ( .A1(n5204), .A2(n5188), .ZN(n5221) );
  AOI21_X2 U6379 ( .B1(n8888), .B2(n5973), .A(n4936), .ZN(n8854) );
  AND2_X1 U6380 ( .A1(n6629), .A2(n6628), .ZN(n7019) );
  INV_X1 U6381 ( .A(n8345), .ZN(n6606) );
  AND2_X1 U6382 ( .A1(n6280), .A2(n6279), .ZN(n4932) );
  OR2_X1 U6383 ( .A1(n10310), .A2(n10302), .ZN(n9078) );
  INV_X1 U6384 ( .A(n9078), .ZN(n6278) );
  INV_X1 U6385 ( .A(n9088), .ZN(n6198) );
  INV_X1 U6386 ( .A(n8992), .ZN(n6511) );
  INV_X1 U6387 ( .A(n8172), .ZN(n7401) );
  NAND2_X2 U6388 ( .A1(n5601), .A2(n9660), .ZN(n9663) );
  OR2_X1 U6389 ( .A1(n6844), .A2(n6843), .ZN(n4933) );
  AND2_X1 U6390 ( .A1(n6272), .A2(n10257), .ZN(n4935) );
  NOR2_X1 U6391 ( .A1(n5972), .A2(n8869), .ZN(n4936) );
  AND2_X1 U6392 ( .A1(n5427), .A2(n5426), .ZN(n4937) );
  NOR2_X1 U6393 ( .A1(n5111), .A2(n10114), .ZN(n4938) );
  INV_X1 U6394 ( .A(n8430), .ZN(n6190) );
  OR2_X1 U6395 ( .A1(n8169), .A2(n9743), .ZN(n4940) );
  OR2_X1 U6396 ( .A1(n8169), .A2(n9812), .ZN(n4941) );
  XNOR2_X1 U6397 ( .A(n6252), .B(n6081), .ZN(n6508) );
  AND3_X1 U6398 ( .A1(n6085), .A2(n6084), .A3(n6083), .ZN(n4942) );
  AND2_X1 U6399 ( .A1(n7457), .A2(n7393), .ZN(n4943) );
  INV_X1 U6400 ( .A(n7505), .ZN(n6378) );
  OR2_X1 U6401 ( .A1(n9082), .A2(n9081), .ZN(P2_U3438) );
  OR2_X1 U6402 ( .A1(n8988), .A2(n8987), .ZN(P2_U3475) );
  OR2_X1 U6403 ( .A1(n8920), .A2(n8919), .ZN(P2_U3217) );
  INV_X1 U6404 ( .A(n8396), .ZN(n6175) );
  AND2_X1 U6405 ( .A1(n6635), .A2(n6634), .ZN(n4947) );
  NAND2_X1 U6406 ( .A1(n9806), .A2(n9381), .ZN(n4949) );
  OR2_X1 U6407 ( .A1(n8576), .A2(n8766), .ZN(n4950) );
  INV_X1 U6408 ( .A(n8412), .ZN(n6081) );
  NAND2_X1 U6409 ( .A1(n7962), .A2(n8039), .ZN(n7963) );
  OR2_X1 U6410 ( .A1(n9571), .A2(n8014), .ZN(n8017) );
  INV_X1 U6411 ( .A(n5639), .ZN(n5640) );
  INV_X1 U6412 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U6413 ( .A1(n8445), .A2(n8613), .ZN(n6516) );
  NAND2_X1 U6414 ( .A1(n4312), .A2(n7334), .ZN(n6836) );
  INV_X1 U6415 ( .A(n8130), .ZN(n5629) );
  OR2_X1 U6416 ( .A1(n5533), .A2(n5532), .ZN(n5537) );
  INV_X1 U6417 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5710) );
  INV_X1 U6418 ( .A(n8766), .ZN(n8582) );
  INV_X1 U6419 ( .A(n8500), .ZN(n6174) );
  INV_X1 U6420 ( .A(n5855), .ZN(n5857) );
  OAI21_X1 U6421 ( .B1(n4312), .B2(n8175), .A(n6836), .ZN(n6838) );
  AND2_X1 U6422 ( .A1(n8140), .A2(n8097), .ZN(n8098) );
  AND2_X1 U6423 ( .A1(n9508), .A2(n5674), .ZN(n5671) );
  INV_X1 U6424 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4960) );
  INV_X1 U6425 ( .A(n5326), .ZN(n5328) );
  NAND2_X1 U6426 ( .A1(n6378), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6379) );
  INV_X1 U6427 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5843) );
  NAND2_X1 U6428 ( .A1(n5974), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5975) );
  INV_X1 U6429 ( .A(n6999), .ZN(n6856) );
  AND2_X1 U6430 ( .A1(n9242), .A2(n4934), .ZN(n7758) );
  INV_X1 U6431 ( .A(n9390), .ZN(n7727) );
  OR2_X1 U6432 ( .A1(n6826), .A2(n6825), .ZN(n6869) );
  INV_X1 U6433 ( .A(n9995), .ZN(n5692) );
  INV_X1 U6434 ( .A(n5542), .ZN(n5543) );
  INV_X1 U6435 ( .A(n5244), .ZN(n5241) );
  NAND2_X1 U6436 ( .A1(n5113), .A2(SI_7_), .ZN(n5141) );
  NOR2_X1 U6437 ( .A1(n5082), .A2(n5081), .ZN(n5083) );
  INV_X1 U6438 ( .A(n6633), .ZN(n6634) );
  NAND2_X1 U6439 ( .A1(n8417), .A2(n8445), .ZN(n8418) );
  INV_X1 U6440 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5724) );
  INV_X1 U6441 ( .A(n8767), .ZN(n8782) );
  AND2_X1 U6442 ( .A1(n5970), .A2(n5969), .ZN(n8893) );
  INV_X1 U6443 ( .A(n8937), .ZN(n8194) );
  OR2_X1 U6444 ( .A1(n6656), .A2(n6142), .ZN(n6286) );
  NAND2_X1 U6445 ( .A1(n6790), .A2(n8563), .ZN(n5884) );
  INV_X1 U6446 ( .A(n10262), .ZN(n8908) );
  OR2_X1 U6447 ( .A1(n6947), .A2(n6195), .ZN(n10265) );
  INV_X1 U6448 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5763) );
  NAND2_X1 U6449 ( .A1(n9292), .A2(n9293), .ZN(n9291) );
  OR2_X1 U6450 ( .A1(n6878), .A2(n8157), .ZN(n9366) );
  NAND2_X1 U6451 ( .A1(n5344), .A2(n4365), .ZN(n5346) );
  OR2_X1 U6452 ( .A1(n9693), .A2(n8151), .ZN(n5693) );
  INV_X1 U6453 ( .A(n9380), .ZN(n7803) );
  OR2_X1 U6454 ( .A1(n7081), .A2(n5604), .ZN(n10095) );
  AND2_X1 U6455 ( .A1(n5539), .A2(n5487), .ZN(n5534) );
  XNOR2_X1 U6456 ( .A(n5219), .B(SI_11_), .ZN(n5220) );
  INV_X1 U6457 ( .A(n8819), .ZN(n8321) );
  INV_X1 U6458 ( .A(n8339), .ZN(n8348) );
  INV_X1 U6459 ( .A(n8350), .ZN(n8336) );
  XNOR2_X1 U6460 ( .A(n6527), .B(n8210), .ZN(n6808) );
  NAND2_X1 U6461 ( .A1(n6611), .A2(n10253), .ZN(n8341) );
  AND3_X1 U6462 ( .A1(n5938), .A2(n5937), .A3(n5936), .ZN(n8892) );
  AND2_X1 U6463 ( .A1(n6417), .A2(n8744), .ZN(n8740) );
  AND2_X1 U6464 ( .A1(n10323), .A2(n10300), .ZN(n8994) );
  AND4_X1 U6465 ( .A1(n6618), .A2(n6286), .A3(n6662), .A4(n6285), .ZN(n6303)
         );
  INV_X1 U6466 ( .A(n6508), .ZN(n6199) );
  OR2_X1 U6467 ( .A1(n6622), .A2(n6612), .ZN(n6166) );
  NAND2_X1 U6468 ( .A1(n6879), .A2(n9660), .ZN(n9369) );
  INV_X1 U6469 ( .A(n10047), .ZN(n10075) );
  INV_X1 U6470 ( .A(n10069), .ZN(n10083) );
  INV_X1 U6471 ( .A(n10030), .ZN(n10081) );
  INV_X1 U6472 ( .A(n10201), .ZN(n10116) );
  INV_X1 U6473 ( .A(n10185), .ZN(n10131) );
  INV_X1 U6474 ( .A(n9697), .ZN(n10142) );
  AND2_X1 U6475 ( .A1(n10248), .A2(n10223), .ZN(n9771) );
  INV_X1 U6476 ( .A(n10213), .ZN(n10223) );
  INV_X1 U6477 ( .A(n9812), .ZN(n9836) );
  INV_X1 U6478 ( .A(n10195), .ZN(n10221) );
  NAND2_X1 U6479 ( .A1(n5574), .A2(n9998), .ZN(n6826) );
  INV_X1 U6480 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5000) );
  INV_X1 U6481 ( .A(n8243), .ZN(n8832) );
  INV_X1 U6482 ( .A(n8748), .ZN(n8654) );
  INV_X1 U6483 ( .A(n8753), .ZN(n8657) );
  OR2_X1 U6484 ( .A1(n6758), .A2(n8744), .ZN(n8756) );
  INV_X1 U6485 ( .A(n8945), .ZN(n8932) );
  INV_X1 U6486 ( .A(n10269), .ZN(n10272) );
  INV_X1 U6487 ( .A(n10323), .ZN(n10320) );
  OR2_X1 U6488 ( .A1(n10310), .A2(n10295), .ZN(n9088) );
  NAND2_X1 U6489 ( .A1(n6662), .A2(n6661), .ZN(n6672) );
  INV_X1 U6490 ( .A(n6459), .ZN(n7172) );
  INV_X1 U6491 ( .A(n9349), .ZN(n9371) );
  INV_X1 U6492 ( .A(n7460), .ZN(n9393) );
  INV_X1 U6493 ( .A(n10014), .ZN(n10089) );
  AND2_X1 U6494 ( .A1(n5657), .A2(n5656), .ZN(n5658) );
  NAND2_X1 U6495 ( .A1(n9663), .A2(n5605), .ZN(n9708) );
  INV_X1 U6496 ( .A(n10153), .ZN(n9667) );
  INV_X2 U6497 ( .A(n10245), .ZN(n10248) );
  INV_X1 U6498 ( .A(n7786), .ZN(n9813) );
  INV_X1 U6499 ( .A(n10232), .ZN(n10230) );
  INV_X1 U6500 ( .A(n10163), .ZN(n10160) );
  AND2_X1 U6501 ( .A1(n9996), .A2(n9995), .ZN(n10163) );
  INV_X1 U6502 ( .A(n7894), .ZN(n10005) );
  INV_X1 U6503 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10328) );
  INV_X1 U6504 ( .A(n8628), .ZN(P2_U3893) );
  NAND2_X1 U6505 ( .A1(n6315), .A2(n6314), .ZN(P2_U3205) );
  INV_X1 U6506 ( .A(n9400), .ZN(P1_U3973) );
  NAND2_X1 U6507 ( .A1(n6365), .A2(n6364), .ZN(P1_U3262) );
  OAI21_X1 U6508 ( .B1(n7852), .B2(n9708), .A(n5658), .ZN(P1_U3265) );
  NOR2_X2 U6509 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5361) );
  NAND3_X1 U6510 ( .A1(n4974), .A2(n4951), .A3(n5361), .ZN(n5098) );
  INV_X1 U6511 ( .A(n5098), .ZN(n4955) );
  NOR2_X1 U6512 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4954) );
  NOR2_X1 U6513 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4953) );
  NOR2_X1 U6514 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4952) );
  NOR2_X2 U6515 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5190) );
  AND4_X2 U6516 ( .A1(n4954), .A2(n4953), .A3(n4952), .A4(n5190), .ZN(n5364)
         );
  NOR2_X1 U6517 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n4958) );
  NOR2_X1 U6518 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4957) );
  NOR2_X1 U6519 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n4956) );
  NAND4_X1 U6520 ( .A1(n5360), .A2(n4958), .A3(n4957), .A4(n4956), .ZN(n4959)
         );
  NAND2_X1 U6521 ( .A1(n5563), .A2(n4960), .ZN(n5566) );
  INV_X1 U6522 ( .A(n5566), .ZN(n4962) );
  NOR2_X1 U6523 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n4961) );
  INV_X1 U6524 ( .A(n4967), .ZN(n4965) );
  NAND2_X1 U6525 ( .A1(n4965), .A2(n4964), .ZN(n7895) );
  XNOR2_X2 U6526 ( .A(n4966), .B(P1_IR_REG_30__SCAN_IN), .ZN(n4971) );
  NAND2_X1 U6527 ( .A1(n4967), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4968) );
  XNOR2_X2 U6528 ( .A(n4968), .B(P1_IR_REG_29__SCAN_IN), .ZN(n4969) );
  AND2_X2 U6529 ( .A1(n4971), .A2(n4969), .ZN(n5102) );
  NAND2_X1 U6530 ( .A1(n5102), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n4970) );
  NAND2_X1 U6531 ( .A1(n5047), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4972) );
  NAND2_X1 U6532 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4973) );
  MUX2_X1 U6533 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4973), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n4976) );
  INV_X1 U6534 ( .A(n5012), .ZN(n4975) );
  INV_X1 U6535 ( .A(n6680), .ZN(n9409) );
  NAND2_X1 U6536 ( .A1(n4304), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4982) );
  INV_X1 U6537 ( .A(n4984), .ZN(n4986) );
  INV_X1 U6538 ( .A(SI_1_), .ZN(n4985) );
  INV_X1 U6539 ( .A(n4992), .ZN(n4990) );
  INV_X1 U6540 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n4987) );
  NAND2_X1 U6541 ( .A1(n4990), .A2(n5027), .ZN(n5005) );
  INV_X1 U6542 ( .A(n5027), .ZN(n4991) );
  NAND2_X1 U6543 ( .A1(n4992), .A2(n4991), .ZN(n4993) );
  NAND2_X1 U6544 ( .A1(n5005), .A2(n4993), .ZN(n6679) );
  NAND2_X1 U6545 ( .A1(n6641), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4994) );
  OAI211_X1 U6546 ( .C1(n6679), .C2(n6641), .A(n5014), .B(n4994), .ZN(n4995)
         );
  OAI21_X1 U6547 ( .B1(n9409), .B2(n5014), .A(n4995), .ZN(n5002) );
  NAND2_X1 U6548 ( .A1(n5102), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n4999) );
  NAND2_X1 U6549 ( .A1(n5046), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4998) );
  NAND2_X1 U6550 ( .A1(n5047), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n4997) );
  NAND2_X1 U6551 ( .A1(n5021), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n4996) );
  NOR2_X1 U6552 ( .A1(n6641), .A2(n9949), .ZN(n5001) );
  XNOR2_X1 U6553 ( .A(n5001), .B(n5000), .ZN(n10010) );
  NAND2_X1 U6554 ( .A1(n7000), .A2(n7151), .ZN(n7147) );
  NAND2_X1 U6555 ( .A1(n5612), .A2(n7147), .ZN(n5004) );
  INV_X1 U6556 ( .A(n5002), .ZN(n7155) );
  OR2_X1 U6557 ( .A1(n9402), .A2(n7155), .ZN(n5003) );
  NAND2_X1 U6558 ( .A1(n5004), .A2(n5003), .ZN(n10144) );
  INV_X1 U6559 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5751) );
  INV_X1 U6560 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6643) );
  INV_X1 U6561 ( .A(SI_2_), .ZN(n5006) );
  NAND2_X1 U6562 ( .A1(n5007), .A2(n5006), .ZN(n5029) );
  INV_X1 U6563 ( .A(n5007), .ZN(n5008) );
  NAND2_X1 U6564 ( .A1(n5008), .A2(SI_2_), .ZN(n5031) );
  NAND2_X1 U6565 ( .A1(n5029), .A2(n5031), .ZN(n5009) );
  INV_X1 U6566 ( .A(n5363), .ZN(n5013) );
  NAND2_X1 U6567 ( .A1(n5102), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5018) );
  NAND2_X1 U6568 ( .A1(n5046), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5017) );
  NAND2_X1 U6569 ( .A1(n5047), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5016) );
  NAND2_X1 U6570 ( .A1(n5021), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5015) );
  NAND2_X1 U6571 ( .A1(n10144), .A2(n10145), .ZN(n5020) );
  NAND2_X1 U6572 ( .A1(n5020), .A2(n5019), .ZN(n7105) );
  NAND2_X1 U6573 ( .A1(n5046), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5026) );
  NAND2_X1 U6574 ( .A1(n5047), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5025) );
  INV_X1 U6575 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5022) );
  INV_X1 U6576 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7108) );
  NAND2_X1 U6577 ( .A1(n5529), .A2(n7108), .ZN(n5023) );
  NAND2_X1 U6578 ( .A1(n5030), .A2(n5029), .ZN(n5032) );
  NAND3_X1 U6579 ( .A1(n5033), .A2(n5032), .A3(n5031), .ZN(n5037) );
  NAND2_X1 U6580 ( .A1(n5034), .A2(n5035), .ZN(n5038) );
  INV_X1 U6581 ( .A(n5035), .ZN(n5036) );
  NAND2_X1 U6582 ( .A1(n5037), .A2(n5036), .ZN(n5079) );
  NAND2_X1 U6583 ( .A1(n5038), .A2(n5079), .ZN(n6667) );
  OR2_X1 U6584 ( .A1(n6667), .A2(n5039), .ZN(n5043) );
  INV_X1 U6585 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6668) );
  OR2_X1 U6586 ( .A1(n6218), .A2(n6668), .ZN(n5042) );
  INV_X1 U6587 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5040) );
  OR2_X1 U6588 ( .A1(n5014), .A2(n9414), .ZN(n5041) );
  AND3_X2 U6589 ( .A1(n5043), .A2(n5042), .A3(n5041), .ZN(n10180) );
  NAND2_X2 U6590 ( .A1(n7949), .A2(n10124), .ZN(n8110) );
  NAND2_X1 U6591 ( .A1(n7105), .A2(n8110), .ZN(n5045) );
  INV_X1 U6592 ( .A(n10180), .ZN(n9175) );
  OR2_X1 U6593 ( .A1(n9401), .A2(n9175), .ZN(n5044) );
  NAND2_X1 U6594 ( .A1(n5045), .A2(n5044), .ZN(n10132) );
  OAI21_X1 U6595 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n5067), .ZN(n6972) );
  OR2_X1 U6596 ( .A1(n5552), .A2(n6972), .ZN(n5051) );
  NAND2_X1 U6597 ( .A1(n6239), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5050) );
  NAND2_X1 U6598 ( .A1(n5046), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5049) );
  NAND2_X1 U6599 ( .A1(n6240), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5048) );
  AND2_X1 U6600 ( .A1(n5079), .A2(n5076), .ZN(n5055) );
  MUX2_X1 U6601 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n4304), .Z(n5052) );
  NAND2_X1 U6602 ( .A1(n5052), .A2(SI_4_), .ZN(n5077) );
  INV_X1 U6603 ( .A(n5052), .ZN(n5054) );
  INV_X1 U6604 ( .A(SI_4_), .ZN(n5053) );
  NAND2_X1 U6605 ( .A1(n5054), .A2(n5053), .ZN(n5080) );
  NAND2_X1 U6606 ( .A1(n5077), .A2(n5080), .ZN(n5056) );
  NAND2_X1 U6607 ( .A1(n5055), .A2(n5056), .ZN(n5059) );
  INV_X1 U6608 ( .A(n5055), .ZN(n5058) );
  INV_X1 U6609 ( .A(n5056), .ZN(n5057) );
  NAND2_X1 U6610 ( .A1(n5058), .A2(n5057), .ZN(n5075) );
  AND2_X1 U6611 ( .A1(n5059), .A2(n5075), .ZN(n6651) );
  NAND2_X1 U6612 ( .A1(n6651), .A2(n6217), .ZN(n5062) );
  OR2_X1 U6613 ( .A1(n5363), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n5060) );
  NAND2_X1 U6614 ( .A1(n5060), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5087) );
  XNOR2_X1 U6615 ( .A(n5087), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6338) );
  AOI22_X1 U6616 ( .A1(n5384), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n6236), .B2(
        n6338), .ZN(n5061) );
  AND2_X2 U6617 ( .A1(n5062), .A2(n5061), .ZN(n10185) );
  XNOR2_X1 U6618 ( .A(n9399), .B(n10185), .ZN(n10133) );
  NAND2_X1 U6619 ( .A1(n10132), .A2(n10133), .ZN(n5064) );
  INV_X1 U6620 ( .A(n9399), .ZN(n7071) );
  NAND2_X1 U6621 ( .A1(n7071), .A2(n10185), .ZN(n5063) );
  INV_X2 U6622 ( .A(n5065), .ZN(n5683) );
  NAND2_X1 U6623 ( .A1(n5683), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5072) );
  NAND2_X1 U6624 ( .A1(n5647), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5071) );
  NAND2_X1 U6625 ( .A1(n6240), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5070) );
  INV_X1 U6626 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5066) );
  NAND2_X1 U6627 ( .A1(n5067), .A2(n5066), .ZN(n5068) );
  NAND2_X1 U6628 ( .A1(n5104), .A2(n5068), .ZN(n7127) );
  OR2_X1 U6629 ( .A1(n5552), .A2(n7127), .ZN(n5069) );
  INV_X1 U6630 ( .A(n5073), .ZN(n5464) );
  MUX2_X1 U6631 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5500), .Z(n5074) );
  OAI21_X1 U6632 ( .B1(n5074), .B2(SI_5_), .A(n5119), .ZN(n5082) );
  NAND3_X1 U6633 ( .A1(n5075), .A2(n5077), .A3(n5082), .ZN(n5085) );
  NAND2_X1 U6634 ( .A1(n5079), .A2(n5078), .ZN(n5084) );
  INV_X1 U6635 ( .A(n5080), .ZN(n5081) );
  NAND2_X1 U6636 ( .A1(n5084), .A2(n5083), .ZN(n5122) );
  NAND2_X1 U6637 ( .A1(n5085), .A2(n5122), .ZN(n6649) );
  OR2_X1 U6638 ( .A1(n6649), .A2(n5039), .ZN(n5091) );
  INV_X1 U6639 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5086) );
  NAND2_X1 U6640 ( .A1(n5087), .A2(n5086), .ZN(n5088) );
  NAND2_X1 U6641 ( .A1(n5088), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5089) );
  XNOR2_X1 U6642 ( .A(n5089), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9448) );
  AOI22_X1 U6643 ( .A1(n5384), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6236), .B2(
        n9448), .ZN(n5090) );
  NAND2_X1 U6644 ( .A1(n5091), .A2(n5090), .ZN(n10192) );
  NAND2_X1 U6645 ( .A1(n9352), .A2(n10192), .ZN(n7936) );
  INV_X1 U6646 ( .A(n9352), .ZN(n9398) );
  INV_X1 U6647 ( .A(n10192), .ZN(n7118) );
  NAND2_X1 U6648 ( .A1(n9398), .A2(n7118), .ZN(n8111) );
  NAND2_X1 U6649 ( .A1(n7936), .A2(n8111), .ZN(n7069) );
  NAND2_X1 U6650 ( .A1(n7068), .A2(n7069), .ZN(n10113) );
  OR2_X1 U6651 ( .A1(n9398), .A2(n10192), .ZN(n10112) );
  NAND2_X1 U6652 ( .A1(n5122), .A2(n5119), .ZN(n5095) );
  MUX2_X1 U6653 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5500), .Z(n5092) );
  NAND2_X1 U6654 ( .A1(n5092), .A2(SI_6_), .ZN(n5120) );
  INV_X1 U6655 ( .A(n5092), .ZN(n5093) );
  INV_X1 U6656 ( .A(SI_6_), .ZN(n9903) );
  NAND2_X1 U6657 ( .A1(n5093), .A2(n9903), .ZN(n5123) );
  AND2_X1 U6658 ( .A1(n5120), .A2(n5123), .ZN(n5094) );
  OR2_X1 U6659 ( .A1(n5095), .A2(n5094), .ZN(n5096) );
  NAND2_X1 U6660 ( .A1(n5095), .A2(n5094), .ZN(n5118) );
  NAND2_X1 U6661 ( .A1(n6658), .A2(n6217), .ZN(n5101) );
  NAND2_X1 U6662 ( .A1(n5098), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5097) );
  MUX2_X1 U6663 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5097), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5099) );
  AND2_X2 U6664 ( .A1(n5101), .A2(n5100), .ZN(n10201) );
  NAND2_X1 U6665 ( .A1(n5682), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5109) );
  NAND2_X1 U6666 ( .A1(n6240), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5108) );
  INV_X1 U6667 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U6668 ( .A1(n5104), .A2(n5103), .ZN(n5105) );
  AND2_X1 U6669 ( .A1(n5133), .A2(n5105), .ZN(n10111) );
  NAND2_X1 U6670 ( .A1(n5529), .A2(n10111), .ZN(n5107) );
  NAND2_X1 U6671 ( .A1(n6239), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5106) );
  NAND4_X1 U6672 ( .A1(n5109), .A2(n5108), .A3(n5107), .A4(n5106), .ZN(n9397)
         );
  INV_X1 U6673 ( .A(n9397), .ZN(n7227) );
  NAND2_X1 U6674 ( .A1(n10201), .A2(n7227), .ZN(n5110) );
  AND2_X1 U6675 ( .A1(n10112), .A2(n5110), .ZN(n5112) );
  INV_X1 U6676 ( .A(n5110), .ZN(n5111) );
  NAND2_X1 U6677 ( .A1(n10201), .A2(n9397), .ZN(n7953) );
  NAND2_X1 U6678 ( .A1(n7953), .A2(n7938), .ZN(n10114) );
  MUX2_X1 U6679 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5464), .Z(n5113) );
  INV_X1 U6680 ( .A(n5113), .ZN(n5115) );
  INV_X1 U6681 ( .A(SI_7_), .ZN(n5114) );
  NAND2_X1 U6682 ( .A1(n5115), .A2(n5114), .ZN(n5116) );
  NAND2_X1 U6683 ( .A1(n5141), .A2(n5116), .ZN(n5124) );
  AND2_X1 U6684 ( .A1(n5124), .A2(n5120), .ZN(n5117) );
  NAND2_X1 U6685 ( .A1(n5118), .A2(n5117), .ZN(n5128) );
  NAND2_X1 U6686 ( .A1(n5122), .A2(n5121), .ZN(n5127) );
  INV_X1 U6687 ( .A(n5123), .ZN(n5125) );
  NAND2_X1 U6688 ( .A1(n5128), .A2(n5142), .ZN(n6670) );
  OR2_X1 U6689 ( .A1(n6670), .A2(n5039), .ZN(n5131) );
  NAND2_X1 U6690 ( .A1(n5148), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5129) );
  XNOR2_X1 U6691 ( .A(n5129), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9476) );
  AOI22_X1 U6692 ( .A1(n5384), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6236), .B2(
        n9476), .ZN(n5130) );
  AND2_X2 U6693 ( .A1(n5131), .A2(n5130), .ZN(n10207) );
  NAND2_X1 U6694 ( .A1(n5683), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5138) );
  NAND2_X1 U6695 ( .A1(n5647), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5137) );
  NAND2_X1 U6696 ( .A1(n5133), .A2(n5132), .ZN(n5134) );
  AND2_X1 U6697 ( .A1(n5169), .A2(n5134), .ZN(n7319) );
  NAND2_X1 U6698 ( .A1(n5529), .A2(n7319), .ZN(n5136) );
  NAND2_X1 U6699 ( .A1(n6240), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5135) );
  NAND4_X1 U6700 ( .A1(n5138), .A2(n5137), .A3(n5136), .A4(n5135), .ZN(n9396)
         );
  NAND2_X1 U6701 ( .A1(n10207), .A2(n9396), .ZN(n5620) );
  INV_X1 U6702 ( .A(n9396), .ZN(n9354) );
  INV_X1 U6703 ( .A(n10207), .ZN(n7320) );
  NAND2_X1 U6704 ( .A1(n9354), .A2(n7320), .ZN(n7940) );
  NAND2_X1 U6705 ( .A1(n5620), .A2(n7940), .ZN(n7957) );
  NAND2_X1 U6706 ( .A1(n7317), .A2(n7957), .ZN(n5140) );
  NAND2_X1 U6707 ( .A1(n10207), .A2(n9354), .ZN(n5139) );
  NAND2_X1 U6708 ( .A1(n5140), .A2(n5139), .ZN(n7276) );
  MUX2_X1 U6709 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n5464), .Z(n5143) );
  INV_X1 U6710 ( .A(n5143), .ZN(n5145) );
  INV_X1 U6711 ( .A(SI_8_), .ZN(n5144) );
  NAND2_X1 U6712 ( .A1(n5145), .A2(n5144), .ZN(n5146) );
  MUX2_X1 U6713 ( .A(n6682), .B(n5147), .S(n5500), .Z(n5178) );
  XNOR2_X1 U6714 ( .A(n5182), .B(n5181), .ZN(n6681) );
  NAND2_X1 U6715 ( .A1(n6681), .A2(n6217), .ZN(n5155) );
  INV_X1 U6716 ( .A(n5148), .ZN(n5150) );
  INV_X1 U6717 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5149) );
  NAND2_X1 U6718 ( .A1(n5150), .A2(n5149), .ZN(n5189) );
  NAND2_X1 U6719 ( .A1(n5189), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5166) );
  INV_X1 U6720 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5151) );
  NAND2_X1 U6721 ( .A1(n5166), .A2(n5151), .ZN(n5152) );
  NAND2_X1 U6722 ( .A1(n5152), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5153) );
  XNOR2_X1 U6723 ( .A(n5153), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6343) );
  AOI22_X1 U6724 ( .A1(n5384), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6236), .B2(
        n6343), .ZN(n5154) );
  NAND2_X1 U6725 ( .A1(n5647), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5163) );
  NAND2_X1 U6726 ( .A1(n6240), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5162) );
  NAND2_X1 U6727 ( .A1(n5683), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5161) );
  INV_X1 U6728 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5157) );
  INV_X1 U6729 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5156) );
  OAI21_X1 U6730 ( .B1(n5169), .B2(n5157), .A(n5156), .ZN(n5159) );
  NAND2_X1 U6731 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n5158) );
  NAND2_X1 U6732 ( .A1(n5159), .A2(n5209), .ZN(n9285) );
  OR2_X1 U6733 ( .A1(n5552), .A2(n9285), .ZN(n5160) );
  OR2_X1 U6734 ( .A1(n10224), .A2(n9211), .ZN(n7964) );
  NAND2_X1 U6735 ( .A1(n7964), .A2(n7969), .ZN(n7278) );
  XNOR2_X1 U6736 ( .A(n5165), .B(n5164), .ZN(n6664) );
  NAND2_X1 U6737 ( .A1(n6664), .A2(n6217), .ZN(n5168) );
  XNOR2_X1 U6738 ( .A(n5166), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9490) );
  AOI22_X1 U6739 ( .A1(n5384), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6236), .B2(
        n9490), .ZN(n5167) );
  NAND2_X1 U6740 ( .A1(n5168), .A2(n5167), .ZN(n10101) );
  XNOR2_X1 U6741 ( .A(n5169), .B(P1_REG3_REG_8__SCAN_IN), .ZN(n10099) );
  NAND2_X1 U6742 ( .A1(n5529), .A2(n10099), .ZN(n5173) );
  NAND2_X1 U6743 ( .A1(n5682), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5172) );
  NAND2_X1 U6744 ( .A1(n6240), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5171) );
  NAND2_X1 U6745 ( .A1(n6239), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5170) );
  NAND4_X1 U6746 ( .A1(n5173), .A2(n5172), .A3(n5171), .A4(n5170), .ZN(n9395)
         );
  NAND2_X1 U6747 ( .A1(n10101), .A2(n9395), .ZN(n10090) );
  AND2_X1 U6748 ( .A1(n7278), .A2(n10090), .ZN(n5174) );
  NAND2_X1 U6749 ( .A1(n7276), .A2(n5174), .ZN(n5177) );
  NOR2_X1 U6750 ( .A1(n10101), .A2(n9395), .ZN(n10092) );
  INV_X1 U6751 ( .A(n9211), .ZN(n9394) );
  NOR2_X1 U6752 ( .A1(n10224), .A2(n9394), .ZN(n5175) );
  AOI21_X1 U6753 ( .B1(n7278), .B2(n10092), .A(n5175), .ZN(n5176) );
  NAND2_X1 U6754 ( .A1(n5177), .A2(n5176), .ZN(n7383) );
  INV_X1 U6755 ( .A(n5178), .ZN(n5179) );
  MUX2_X1 U6756 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n4304), .Z(n5183) );
  INV_X1 U6757 ( .A(n5183), .ZN(n5185) );
  INV_X1 U6758 ( .A(SI_10_), .ZN(n5184) );
  NAND2_X1 U6759 ( .A1(n5185), .A2(n5184), .ZN(n5186) );
  MUX2_X1 U6760 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n5517), .Z(n5219) );
  XNOR2_X1 U6761 ( .A(n5221), .B(n5220), .ZN(n6699) );
  NAND2_X1 U6762 ( .A1(n6699), .A2(n6217), .ZN(n5194) );
  INV_X1 U6763 ( .A(n5189), .ZN(n5191) );
  NAND2_X1 U6764 ( .A1(n5191), .A2(n5190), .ZN(n5205) );
  NAND2_X1 U6765 ( .A1(n5227), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5192) );
  XNOR2_X1 U6766 ( .A(n5192), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7311) );
  AOI22_X1 U6767 ( .A1(n5384), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6236), .B2(
        n7311), .ZN(n5193) );
  NAND2_X1 U6768 ( .A1(n5683), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5200) );
  NAND2_X1 U6769 ( .A1(n5647), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5199) );
  NAND2_X1 U6770 ( .A1(n6240), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5198) );
  INV_X1 U6771 ( .A(n5195), .ZN(n5211) );
  NAND2_X1 U6772 ( .A1(n5211), .A2(n4494), .ZN(n5196) );
  NAND2_X1 U6773 ( .A1(n5231), .A2(n5196), .ZN(n9326) );
  OR2_X1 U6774 ( .A1(n5552), .A2(n9326), .ZN(n5197) );
  OR2_X1 U6775 ( .A1(n7553), .A2(n7711), .ZN(n7973) );
  NAND2_X1 U6776 ( .A1(n7553), .A2(n7711), .ZN(n7972) );
  NAND2_X1 U6777 ( .A1(n7973), .A2(n7972), .ZN(n7457) );
  NAND2_X1 U6778 ( .A1(n5202), .A2(n5201), .ZN(n5203) );
  NAND2_X1 U6779 ( .A1(n5204), .A2(n5203), .ZN(n6687) );
  NAND2_X1 U6780 ( .A1(n5205), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5206) );
  XNOR2_X1 U6781 ( .A(n5206), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7196) );
  AOI22_X1 U6782 ( .A1(n5384), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6236), .B2(
        n7196), .ZN(n5207) );
  NAND2_X1 U6783 ( .A1(n6239), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5215) );
  NAND2_X1 U6784 ( .A1(n5682), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5214) );
  NAND2_X1 U6785 ( .A1(n6240), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5213) );
  NAND2_X1 U6786 ( .A1(n5209), .A2(n7188), .ZN(n5210) );
  NAND2_X1 U6787 ( .A1(n5211), .A2(n5210), .ZN(n9167) );
  OR2_X1 U6788 ( .A1(n5552), .A2(n9167), .ZN(n5212) );
  OR2_X1 U6789 ( .A1(n9169), .A2(n7460), .ZN(n8062) );
  NAND2_X1 U6790 ( .A1(n9169), .A2(n7460), .ZN(n7971) );
  NAND2_X1 U6791 ( .A1(n8062), .A2(n7971), .ZN(n7393) );
  NAND2_X1 U6792 ( .A1(n7383), .A2(n4943), .ZN(n5218) );
  NOR2_X1 U6793 ( .A1(n9169), .A2(n9393), .ZN(n7454) );
  INV_X1 U6794 ( .A(n7711), .ZN(n9392) );
  NOR2_X1 U6795 ( .A1(n7553), .A2(n9392), .ZN(n5216) );
  AOI21_X1 U6796 ( .B1(n7457), .B2(n7454), .A(n5216), .ZN(n5217) );
  NAND2_X1 U6797 ( .A1(n5218), .A2(n5217), .ZN(n7513) );
  MUX2_X1 U6798 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6640), .Z(n5222) );
  NAND2_X1 U6799 ( .A1(n5225), .A2(n5224), .ZN(n5226) );
  NAND2_X1 U6800 ( .A1(n6790), .A2(n6217), .ZN(n5229) );
  OAI21_X1 U6801 ( .B1(n5227), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5247) );
  XNOR2_X1 U6802 ( .A(n5247), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6346) );
  AOI22_X1 U6803 ( .A1(n5384), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6236), .B2(
        n6346), .ZN(n5228) );
  NAND2_X1 U6804 ( .A1(n5647), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5236) );
  NAND2_X1 U6805 ( .A1(n6240), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5235) );
  NAND2_X1 U6806 ( .A1(n5231), .A2(n5230), .ZN(n5232) );
  AND2_X1 U6807 ( .A1(n5253), .A2(n5232), .ZN(n9231) );
  NAND2_X1 U6808 ( .A1(n5529), .A2(n9231), .ZN(n5234) );
  NAND2_X1 U6809 ( .A1(n6239), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5233) );
  NAND4_X1 U6810 ( .A1(n5236), .A2(n5235), .A3(n5234), .A4(n5233), .ZN(n9391)
         );
  NAND2_X1 U6811 ( .A1(n9234), .A2(n9391), .ZN(n7974) );
  NAND2_X1 U6812 ( .A1(n7515), .A2(n7977), .ZN(n8065) );
  NAND2_X1 U6813 ( .A1(n7974), .A2(n8065), .ZN(n8124) );
  NAND2_X1 U6814 ( .A1(n7513), .A2(n8124), .ZN(n7512) );
  NAND2_X1 U6815 ( .A1(n9234), .A2(n7977), .ZN(n5237) );
  NAND2_X1 U6816 ( .A1(n7512), .A2(n5237), .ZN(n7531) );
  MUX2_X1 U6817 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n5517), .Z(n5238) );
  NAND2_X1 U6818 ( .A1(n5238), .A2(SI_13_), .ZN(n5263) );
  INV_X1 U6819 ( .A(n5238), .ZN(n5240) );
  INV_X1 U6820 ( .A(SI_13_), .ZN(n5239) );
  NAND2_X1 U6821 ( .A1(n5240), .A2(n5239), .ZN(n5266) );
  NAND2_X1 U6822 ( .A1(n5263), .A2(n5266), .ZN(n5242) );
  NAND2_X1 U6823 ( .A1(n5241), .A2(n5242), .ZN(n5245) );
  INV_X1 U6824 ( .A(n5242), .ZN(n5243) );
  NAND2_X1 U6825 ( .A1(n6819), .A2(n6217), .ZN(n5251) );
  INV_X1 U6826 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5246) );
  NAND2_X1 U6827 ( .A1(n5247), .A2(n5246), .ZN(n5248) );
  NAND2_X1 U6828 ( .A1(n5248), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5249) );
  XNOR2_X1 U6829 ( .A(n5249), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7615) );
  AOI22_X1 U6830 ( .A1(n6236), .A2(n7615), .B1(n5384), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n5250) );
  NAND2_X1 U6831 ( .A1(n5682), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5258) );
  NAND2_X1 U6832 ( .A1(n6239), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5257) );
  INV_X1 U6833 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U6834 ( .A1(n5253), .A2(n5252), .ZN(n5254) );
  AND2_X1 U6835 ( .A1(n5277), .A2(n5254), .ZN(n9302) );
  NAND2_X1 U6836 ( .A1(n5529), .A2(n9302), .ZN(n5256) );
  NAND2_X1 U6837 ( .A1(n6240), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5255) );
  NAND4_X1 U6838 ( .A1(n5258), .A2(n5257), .A3(n5256), .A4(n5255), .ZN(n9390)
         );
  NAND2_X1 U6839 ( .A1(n7728), .A2(n9390), .ZN(n8069) );
  NAND2_X1 U6840 ( .A1(n8069), .A2(n8064), .ZN(n7530) );
  NAND2_X1 U6841 ( .A1(n7531), .A2(n7530), .ZN(n7529) );
  NAND2_X1 U6842 ( .A1(n7728), .A2(n7727), .ZN(n5259) );
  NAND2_X1 U6843 ( .A1(n7529), .A2(n5259), .ZN(n7652) );
  MUX2_X1 U6844 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6640), .Z(n5260) );
  NAND2_X1 U6845 ( .A1(n5260), .A2(SI_14_), .ZN(n5286) );
  OAI21_X1 U6846 ( .B1(n5260), .B2(SI_14_), .A(n5286), .ZN(n5268) );
  AND2_X1 U6847 ( .A1(n5268), .A2(n5263), .ZN(n5261) );
  NAND2_X1 U6848 ( .A1(n5262), .A2(n5261), .ZN(n5271) );
  INV_X1 U6849 ( .A(n5266), .ZN(n5267) );
  NAND2_X1 U6850 ( .A1(n5289), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5273) );
  XNOR2_X1 U6851 ( .A(n5273), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10026) );
  AOI22_X1 U6852 ( .A1(n5384), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6236), .B2(
        n10026), .ZN(n5274) );
  NAND2_X2 U6853 ( .A1(n5275), .A2(n5274), .ZN(n9776) );
  NAND2_X1 U6854 ( .A1(n5647), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5282) );
  NAND2_X1 U6855 ( .A1(n5683), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5281) );
  INV_X1 U6856 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5276) );
  NAND2_X1 U6857 ( .A1(n5277), .A2(n5276), .ZN(n5278) );
  AND2_X1 U6858 ( .A1(n5295), .A2(n5278), .ZN(n9140) );
  NAND2_X1 U6859 ( .A1(n5529), .A2(n9140), .ZN(n5280) );
  NAND2_X1 U6860 ( .A1(n6240), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5279) );
  NAND4_X1 U6861 ( .A1(n5282), .A2(n5281), .A3(n5280), .A4(n5279), .ZN(n9389)
         );
  NAND2_X1 U6862 ( .A1(n9776), .A2(n9389), .ZN(n5283) );
  NAND2_X1 U6863 ( .A1(n7652), .A2(n5283), .ZN(n5285) );
  INV_X1 U6864 ( .A(n9389), .ZN(n5625) );
  NAND2_X1 U6865 ( .A1(n9143), .A2(n5625), .ZN(n5284) );
  NAND2_X1 U6866 ( .A1(n5287), .A2(n5286), .ZN(n5306) );
  MUX2_X1 U6867 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6640), .Z(n5307) );
  XNOR2_X1 U6868 ( .A(n5307), .B(SI_15_), .ZN(n5288) );
  XNOR2_X1 U6869 ( .A(n5306), .B(n5288), .ZN(n6977) );
  NAND2_X1 U6870 ( .A1(n6977), .A2(n6217), .ZN(n5293) );
  NOR2_X1 U6871 ( .A1(n5289), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5312) );
  OR2_X1 U6872 ( .A1(n5312), .A2(n5290), .ZN(n5291) );
  XNOR2_X1 U6873 ( .A(n5291), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10039) );
  AOI22_X1 U6874 ( .A1(n5384), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6236), .B2(
        n10039), .ZN(n5292) );
  NAND2_X1 U6875 ( .A1(n5682), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5300) );
  INV_X1 U6876 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5294) );
  NAND2_X1 U6877 ( .A1(n5295), .A2(n5294), .ZN(n5296) );
  AND2_X1 U6878 ( .A1(n5317), .A2(n5296), .ZN(n9363) );
  NAND2_X1 U6879 ( .A1(n5529), .A2(n9363), .ZN(n5299) );
  NAND2_X1 U6880 ( .A1(n6240), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5298) );
  NAND2_X1 U6881 ( .A1(n6239), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5297) );
  NAND4_X1 U6882 ( .A1(n5300), .A2(n5299), .A3(n5298), .A4(n5297), .ZN(n9388)
         );
  NOR2_X1 U6883 ( .A1(n9835), .A2(n9388), .ZN(n5301) );
  NAND2_X1 U6884 ( .A1(n9835), .A2(n9388), .ZN(n5302) );
  INV_X1 U6885 ( .A(n5307), .ZN(n5304) );
  INV_X1 U6886 ( .A(SI_15_), .ZN(n5303) );
  NAND2_X1 U6887 ( .A1(n5304), .A2(n5303), .ZN(n5305) );
  NAND2_X1 U6888 ( .A1(n5306), .A2(n5305), .ZN(n5309) );
  NAND2_X1 U6889 ( .A1(n5307), .A2(SI_15_), .ZN(n5308) );
  MUX2_X1 U6890 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n6640), .Z(n5326) );
  XNOR2_X1 U6891 ( .A(n5326), .B(SI_16_), .ZN(n5310) );
  XNOR2_X1 U6892 ( .A(n5331), .B(n5310), .ZN(n6992) );
  NAND2_X1 U6893 ( .A1(n6992), .A2(n6217), .ZN(n5315) );
  INV_X1 U6894 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5311) );
  NAND2_X1 U6895 ( .A1(n5312), .A2(n5311), .ZN(n5313) );
  NAND2_X1 U6896 ( .A1(n5313), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5334) );
  XNOR2_X1 U6897 ( .A(n5334), .B(P1_IR_REG_16__SCAN_IN), .ZN(n6351) );
  AOI22_X1 U6898 ( .A1(n5384), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6236), .B2(
        n6351), .ZN(n5314) );
  NAND2_X1 U6899 ( .A1(n5317), .A2(n4496), .ZN(n5318) );
  NAND2_X1 U6900 ( .A1(n5340), .A2(n5318), .ZN(n9246) );
  OR2_X1 U6901 ( .A1(n9246), .A2(n5552), .ZN(n5323) );
  NAND2_X1 U6902 ( .A1(n5683), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5320) );
  NAND2_X1 U6903 ( .A1(n5682), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5319) );
  AND2_X1 U6904 ( .A1(n5320), .A2(n5319), .ZN(n5322) );
  NAND2_X1 U6905 ( .A1(n6240), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5321) );
  OR2_X1 U6906 ( .A1(n9764), .A2(n7750), .ZN(n7990) );
  NAND2_X1 U6907 ( .A1(n9764), .A2(n7750), .ZN(n8075) );
  NAND2_X1 U6908 ( .A1(n7990), .A2(n8075), .ZN(n9690) );
  INV_X1 U6909 ( .A(n7750), .ZN(n9387) );
  NAND2_X1 U6910 ( .A1(n9764), .A2(n9387), .ZN(n5324) );
  INV_X1 U6911 ( .A(n7666), .ZN(n5344) );
  INV_X1 U6912 ( .A(SI_16_), .ZN(n5327) );
  NAND2_X1 U6913 ( .A1(n5328), .A2(n5327), .ZN(n5329) );
  OAI21_X2 U6914 ( .B1(n5331), .B2(n5330), .A(n5329), .ZN(n5350) );
  INV_X1 U6915 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7146) );
  INV_X1 U6916 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5332) );
  MUX2_X1 U6917 ( .A(n7146), .B(n5332), .S(n6640), .Z(n5347) );
  XNOR2_X1 U6918 ( .A(n5350), .B(n5349), .ZN(n7087) );
  NAND2_X1 U6919 ( .A1(n7087), .A2(n6217), .ZN(n5338) );
  INV_X1 U6920 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U6921 ( .A1(n5334), .A2(n5333), .ZN(n5335) );
  NAND2_X1 U6922 ( .A1(n5335), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5336) );
  XNOR2_X1 U6923 ( .A(n5336), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10057) );
  AOI22_X1 U6924 ( .A1(n5384), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6236), .B2(
        n10057), .ZN(n5337) );
  INV_X1 U6925 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6926 ( .A1(n5340), .A2(n5339), .ZN(n5341) );
  NAND2_X1 U6927 ( .A1(n5373), .A2(n5341), .ZN(n7673) );
  AOI22_X1 U6928 ( .A1(n5683), .A2(P1_REG0_REG_17__SCAN_IN), .B1(n5682), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U6929 ( .A1(n6240), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5342) );
  OAI211_X1 U6930 ( .C1(n7673), .C2(n5552), .A(n5343), .B(n5342), .ZN(n9386)
         );
  OR2_X1 U6931 ( .A1(n9828), .A2(n9386), .ZN(n5345) );
  NAND2_X1 U6932 ( .A1(n5346), .A2(n5345), .ZN(n9672) );
  INV_X1 U6933 ( .A(n5347), .ZN(n5348) );
  MUX2_X1 U6934 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5517), .Z(n5351) );
  NAND2_X1 U6935 ( .A1(n5351), .A2(SI_18_), .ZN(n5380) );
  INV_X1 U6936 ( .A(n5351), .ZN(n5352) );
  INV_X1 U6937 ( .A(SI_18_), .ZN(n9928) );
  NAND2_X1 U6938 ( .A1(n5352), .A2(n9928), .ZN(n5353) );
  NAND2_X1 U6939 ( .A1(n5380), .A2(n5353), .ZN(n5355) );
  INV_X1 U6940 ( .A(n5355), .ZN(n5354) );
  NAND2_X1 U6941 ( .A1(n5356), .A2(n5355), .ZN(n5357) );
  NAND2_X1 U6942 ( .A1(n5381), .A2(n5357), .ZN(n7143) );
  NOR2_X1 U6943 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5359) );
  INV_X1 U6944 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5358) );
  NAND4_X1 U6945 ( .A1(n5361), .A2(n5360), .A3(n5359), .A4(n5358), .ZN(n5362)
         );
  NAND2_X1 U6946 ( .A1(n5365), .A2(n5364), .ZN(n5367) );
  NAND2_X1 U6947 ( .A1(n5367), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5366) );
  MUX2_X1 U6948 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5366), .S(
        P1_IR_REG_18__SCAN_IN), .Z(n5370) );
  AND2_X1 U6949 ( .A1(n5370), .A2(n5575), .ZN(n10082) );
  AOI22_X1 U6950 ( .A1(n5384), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6236), .B2(
        n10082), .ZN(n5371) );
  INV_X1 U6951 ( .A(n5683), .ZN(n5494) );
  INV_X1 U6952 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U6953 ( .A1(n5373), .A2(n4497), .ZN(n5374) );
  NAND2_X1 U6954 ( .A1(n5387), .A2(n5374), .ZN(n9676) );
  OR2_X1 U6955 ( .A1(n9676), .A2(n5552), .ZN(n5376) );
  AOI22_X1 U6956 ( .A1(n6240), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n5647), .B2(
        P1_REG1_REG_18__SCAN_IN), .ZN(n5375) );
  OAI211_X1 U6957 ( .C1(n5494), .C2(n5377), .A(n5376), .B(n5375), .ZN(n9385)
         );
  NOR2_X1 U6958 ( .A1(n9754), .A2(n9385), .ZN(n5378) );
  NAND2_X1 U6959 ( .A1(n9754), .A2(n9385), .ZN(n5379) );
  MUX2_X1 U6960 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n5517), .Z(n5394) );
  XNOR2_X1 U6961 ( .A(n5396), .B(n5395), .ZN(n7243) );
  NAND2_X1 U6962 ( .A1(n7243), .A2(n6217), .ZN(n5386) );
  NAND2_X1 U6963 ( .A1(n5575), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5383) );
  INV_X1 U6964 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5382) );
  INV_X2 U6965 ( .A(n8151), .ZN(n8175) );
  AOI22_X1 U6966 ( .A1(n5384), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6236), .B2(
        n8175), .ZN(n5385) );
  INV_X1 U6967 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9184) );
  NAND2_X1 U6968 ( .A1(n5387), .A2(n9184), .ZN(n5388) );
  NAND2_X1 U6969 ( .A1(n5399), .A2(n5388), .ZN(n9661) );
  OR2_X1 U6970 ( .A1(n9661), .A2(n5552), .ZN(n5393) );
  INV_X1 U6971 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9662) );
  NAND2_X1 U6972 ( .A1(n5682), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U6973 ( .A1(n6239), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5389) );
  OAI211_X1 U6974 ( .C1(n5686), .C2(n9662), .A(n5390), .B(n5389), .ZN(n5391)
         );
  INV_X1 U6975 ( .A(n5391), .ZN(n5392) );
  NAND2_X1 U6976 ( .A1(n5393), .A2(n5392), .ZN(n9384) );
  INV_X1 U6977 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7332) );
  MUX2_X1 U6978 ( .A(n9854), .B(n7332), .S(n5659), .Z(n5413) );
  XNOR2_X1 U6979 ( .A(n5413), .B(SI_20_), .ZN(n5410) );
  XNOR2_X1 U6980 ( .A(n5411), .B(n5410), .ZN(n7303) );
  NAND2_X1 U6981 ( .A1(n7303), .A2(n6217), .ZN(n5398) );
  OR2_X1 U6982 ( .A1(n6218), .A2(n7332), .ZN(n5397) );
  INV_X1 U6983 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9296) );
  NAND2_X1 U6984 ( .A1(n5399), .A2(n9296), .ZN(n5400) );
  NAND2_X1 U6985 ( .A1(n5420), .A2(n5400), .ZN(n9295) );
  INV_X1 U6986 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U6987 ( .A1(n5647), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5402) );
  NAND2_X1 U6988 ( .A1(n5683), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5401) );
  OAI211_X1 U6989 ( .C1(n5686), .C2(n5403), .A(n5402), .B(n5401), .ZN(n5404)
         );
  INV_X1 U6990 ( .A(n5404), .ZN(n5405) );
  OAI21_X1 U6991 ( .B1(n9295), .B2(n5552), .A(n5405), .ZN(n9383) );
  OR2_X1 U6992 ( .A1(n9816), .A2(n9383), .ZN(n5406) );
  OR2_X1 U6993 ( .A1(n9822), .A2(n9384), .ZN(n9636) );
  AND2_X1 U6994 ( .A1(n5406), .A2(n9636), .ZN(n5407) );
  NAND2_X1 U6995 ( .A1(n9816), .A2(n9383), .ZN(n5408) );
  NAND2_X1 U6996 ( .A1(n5411), .A2(n5410), .ZN(n5415) );
  INV_X1 U6997 ( .A(SI_20_), .ZN(n5412) );
  NAND2_X1 U6998 ( .A1(n5413), .A2(n5412), .ZN(n5414) );
  INV_X1 U6999 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7398) );
  INV_X1 U7000 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7403) );
  MUX2_X1 U7001 ( .A(n7398), .B(n7403), .S(n5659), .Z(n5427) );
  XNOR2_X1 U7002 ( .A(n5427), .B(SI_21_), .ZN(n5416) );
  XNOR2_X1 U7003 ( .A(n5430), .B(n5416), .ZN(n7397) );
  NAND2_X1 U7004 ( .A1(n7397), .A2(n6217), .ZN(n5418) );
  OR2_X1 U7005 ( .A1(n6218), .A2(n7403), .ZN(n5417) );
  INV_X1 U7006 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9219) );
  NAND2_X1 U7007 ( .A1(n5420), .A2(n9219), .ZN(n5421) );
  AND2_X1 U7008 ( .A1(n5438), .A2(n5421), .ZN(n9630) );
  INV_X1 U7009 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U7010 ( .A1(n5683), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5423) );
  NAND2_X1 U7011 ( .A1(n5647), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5422) );
  OAI211_X1 U7012 ( .C1(n5424), .C2(n5686), .A(n5423), .B(n5422), .ZN(n5425)
         );
  AOI21_X1 U7013 ( .B1(n9630), .B2(n5529), .A(n5425), .ZN(n7790) );
  OR2_X1 U7014 ( .A1(n7786), .A2(n7790), .ZN(n8002) );
  NAND2_X1 U7015 ( .A1(n7786), .A2(n7790), .ZN(n8003) );
  NAND2_X1 U7016 ( .A1(n8002), .A2(n8003), .ZN(n9624) );
  INV_X1 U7017 ( .A(n7790), .ZN(n9382) );
  NAND2_X1 U7018 ( .A1(n7786), .A2(n9382), .ZN(n9601) );
  INV_X1 U7019 ( .A(SI_21_), .ZN(n5426) );
  INV_X1 U7020 ( .A(n5427), .ZN(n5428) );
  NAND2_X1 U7021 ( .A1(n5428), .A2(SI_21_), .ZN(n5429) );
  INV_X1 U7022 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7485) );
  INV_X1 U7023 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7482) );
  MUX2_X1 U7024 ( .A(n7485), .B(n7482), .S(n5659), .Z(n5432) );
  INV_X1 U7025 ( .A(SI_22_), .ZN(n5431) );
  NAND2_X1 U7026 ( .A1(n5432), .A2(n5431), .ZN(n5446) );
  INV_X1 U7027 ( .A(n5432), .ZN(n5433) );
  NAND2_X1 U7028 ( .A1(n5433), .A2(SI_22_), .ZN(n5434) );
  NAND2_X1 U7029 ( .A1(n5446), .A2(n5434), .ZN(n5447) );
  XNOR2_X1 U7030 ( .A(n5448), .B(n5447), .ZN(n7480) );
  NAND2_X1 U7031 ( .A1(n7480), .A2(n6217), .ZN(n5436) );
  OR2_X1 U7032 ( .A1(n6218), .A2(n7482), .ZN(n5435) );
  INV_X1 U7033 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9315) );
  NAND2_X1 U7034 ( .A1(n5438), .A2(n9315), .ZN(n5439) );
  NAND2_X1 U7035 ( .A1(n5454), .A2(n5439), .ZN(n9613) );
  INV_X1 U7036 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9914) );
  NAND2_X1 U7037 ( .A1(n6240), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U7038 ( .A1(n5647), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5440) );
  OAI211_X1 U7039 ( .C1(n5494), .C2(n9914), .A(n5441), .B(n5440), .ZN(n5442)
         );
  INV_X1 U7040 ( .A(n5442), .ZN(n5443) );
  OR2_X1 U7041 ( .A1(n9806), .A2(n9381), .ZN(n5445) );
  INV_X1 U7042 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7579) );
  INV_X1 U7043 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7574) );
  INV_X1 U7044 ( .A(SI_23_), .ZN(n9878) );
  NAND2_X1 U7045 ( .A1(n5449), .A2(n9878), .ZN(n5463) );
  INV_X1 U7046 ( .A(n5449), .ZN(n5450) );
  NAND2_X1 U7047 ( .A1(n5450), .A2(SI_23_), .ZN(n5451) );
  NAND2_X1 U7048 ( .A1(n7576), .A2(n6217), .ZN(n5453) );
  OR2_X1 U7049 ( .A1(n6218), .A2(n7574), .ZN(n5452) );
  INV_X1 U7050 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9154) );
  NAND2_X1 U7051 ( .A1(n5454), .A2(n9154), .ZN(n5455) );
  AND2_X1 U7052 ( .A1(n5471), .A2(n5455), .ZN(n9595) );
  NAND2_X1 U7053 ( .A1(n9595), .A2(n5529), .ZN(n5460) );
  INV_X1 U7054 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9940) );
  NAND2_X1 U7055 ( .A1(n5647), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U7056 ( .A1(n6240), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5456) );
  OAI211_X1 U7057 ( .C1(n5494), .C2(n9940), .A(n5457), .B(n5456), .ZN(n5458)
         );
  INV_X1 U7058 ( .A(n5458), .ZN(n5459) );
  NAND2_X1 U7059 ( .A1(n5460), .A2(n5459), .ZN(n9380) );
  INV_X1 U7060 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7622) );
  INV_X1 U7061 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7623) );
  MUX2_X1 U7062 ( .A(n7622), .B(n7623), .S(n5659), .Z(n5466) );
  INV_X1 U7063 ( .A(SI_24_), .ZN(n5465) );
  NAND2_X1 U7064 ( .A1(n5466), .A2(n5465), .ZN(n5482) );
  INV_X1 U7065 ( .A(n5466), .ZN(n5467) );
  NAND2_X1 U7066 ( .A1(n5467), .A2(SI_24_), .ZN(n5468) );
  XNOR2_X1 U7067 ( .A(n5481), .B(n5480), .ZN(n7621) );
  NAND2_X1 U7068 ( .A1(n7621), .A2(n6217), .ZN(n5470) );
  OR2_X1 U7069 ( .A1(n6218), .A2(n7623), .ZN(n5469) );
  INV_X1 U7070 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9269) );
  NAND2_X1 U7071 ( .A1(n5471), .A2(n9269), .ZN(n5472) );
  NAND2_X1 U7072 ( .A1(n5490), .A2(n5472), .ZN(n9576) );
  INV_X1 U7073 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9575) );
  NAND2_X1 U7074 ( .A1(n6239), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U7075 ( .A1(n5682), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5473) );
  OAI211_X1 U7076 ( .C1(n9575), .C2(n5686), .A(n5474), .B(n5473), .ZN(n5475)
         );
  INV_X1 U7077 ( .A(n5475), .ZN(n5476) );
  AND2_X1 U7078 ( .A1(n9578), .A2(n9379), .ZN(n5479) );
  OR2_X1 U7079 ( .A1(n9578), .A2(n9379), .ZN(n5478) );
  NAND2_X1 U7080 ( .A1(n5481), .A2(n5480), .ZN(n5483) );
  NAND2_X1 U7081 ( .A1(n5483), .A2(n5482), .ZN(n5536) );
  INV_X1 U7082 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7664) );
  INV_X1 U7083 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10006) );
  MUX2_X1 U7084 ( .A(n7664), .B(n10006), .S(n5659), .Z(n5485) );
  INV_X1 U7085 ( .A(SI_25_), .ZN(n5484) );
  NAND2_X1 U7086 ( .A1(n5485), .A2(n5484), .ZN(n5539) );
  INV_X1 U7087 ( .A(n5485), .ZN(n5486) );
  NAND2_X1 U7088 ( .A1(n5486), .A2(SI_25_), .ZN(n5487) );
  XNOR2_X1 U7089 ( .A(n5536), .B(n5534), .ZN(n7663) );
  NAND2_X1 U7090 ( .A1(n7663), .A2(n6217), .ZN(n5489) );
  OR2_X1 U7091 ( .A1(n6218), .A2(n10006), .ZN(n5488) );
  INV_X1 U7092 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n7831) );
  NAND2_X1 U7093 ( .A1(n5490), .A2(n7831), .ZN(n5491) );
  AND2_X1 U7094 ( .A1(n5506), .A2(n5491), .ZN(n7830) );
  NAND2_X1 U7095 ( .A1(n7830), .A2(n5529), .ZN(n5497) );
  INV_X1 U7096 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9915) );
  NAND2_X1 U7097 ( .A1(n6240), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U7098 ( .A1(n5682), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5492) );
  OAI211_X1 U7099 ( .C1(n5494), .C2(n9915), .A(n5493), .B(n5492), .ZN(n5495)
         );
  INV_X1 U7100 ( .A(n5495), .ZN(n5496) );
  NOR2_X1 U7101 ( .A1(n9558), .A2(n9378), .ZN(n5498) );
  NAND2_X1 U7102 ( .A1(n5536), .A2(n5534), .ZN(n5499) );
  INV_X1 U7103 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9102) );
  INV_X1 U7104 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7679) );
  MUX2_X1 U7105 ( .A(n9102), .B(n7679), .S(n5659), .Z(n5502) );
  INV_X1 U7106 ( .A(SI_26_), .ZN(n5501) );
  NAND2_X1 U7107 ( .A1(n5502), .A2(n5501), .ZN(n5531) );
  INV_X1 U7108 ( .A(n5502), .ZN(n5503) );
  NAND2_X1 U7109 ( .A1(n5503), .A2(SI_26_), .ZN(n5504) );
  OR2_X1 U7110 ( .A1(n6218), .A2(n7679), .ZN(n5505) );
  INV_X1 U7111 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n7874) );
  NAND2_X1 U7112 ( .A1(n5506), .A2(n7874), .ZN(n5507) );
  NAND2_X1 U7113 ( .A1(n7873), .A2(n5102), .ZN(n5512) );
  INV_X1 U7114 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9540) );
  NAND2_X1 U7115 ( .A1(n5647), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5509) );
  NAND2_X1 U7116 ( .A1(n5683), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5508) );
  OAI211_X1 U7117 ( .C1(n9540), .C2(n5686), .A(n5509), .B(n5508), .ZN(n5510)
         );
  INV_X1 U7118 ( .A(n5510), .ZN(n5511) );
  AND2_X1 U7119 ( .A1(n9546), .A2(n9377), .ZN(n5514) );
  OR2_X1 U7120 ( .A1(n9546), .A2(n9377), .ZN(n5513) );
  INV_X1 U7121 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9099) );
  INV_X1 U7122 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10004) );
  MUX2_X1 U7123 ( .A(n9099), .B(n10004), .S(n5659), .Z(n5519) );
  INV_X1 U7124 ( .A(SI_27_), .ZN(n5518) );
  NAND2_X1 U7125 ( .A1(n5519), .A2(n5518), .ZN(n5530) );
  INV_X1 U7126 ( .A(n5519), .ZN(n5520) );
  NAND2_X1 U7127 ( .A1(n5520), .A2(SI_27_), .ZN(n5542) );
  AND2_X1 U7128 ( .A1(n5530), .A2(n5542), .ZN(n5521) );
  OR2_X1 U7129 ( .A1(n6218), .A2(n10004), .ZN(n5523) );
  INV_X1 U7130 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U7131 ( .A1(n5682), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U7132 ( .A1(n6239), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5525) );
  OAI211_X1 U7133 ( .C1(n5527), .C2(n5686), .A(n5526), .B(n5525), .ZN(n5528)
         );
  NAND2_X1 U7134 ( .A1(n9715), .A2(n9116), .ZN(n8025) );
  NAND2_X1 U7135 ( .A1(n8080), .A2(n8025), .ZN(n5639) );
  INV_X1 U7136 ( .A(n9116), .ZN(n9376) );
  AND2_X1 U7137 ( .A1(n5531), .A2(n5530), .ZN(n5538) );
  INV_X1 U7138 ( .A(n5538), .ZN(n5533) );
  AND2_X1 U7139 ( .A1(n5534), .A2(n5537), .ZN(n5535) );
  NAND2_X1 U7140 ( .A1(n5536), .A2(n5535), .ZN(n5545) );
  INV_X1 U7141 ( .A(n5537), .ZN(n5541) );
  AND2_X1 U7142 ( .A1(n5539), .A2(n5538), .ZN(n5540) );
  AOI21_X2 U7143 ( .B1(n5545), .B2(n5544), .A(n5543), .ZN(n6203) );
  INV_X1 U7144 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8188) );
  INV_X1 U7145 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9842) );
  MUX2_X1 U7146 ( .A(n8188), .B(n9842), .S(n5659), .Z(n5661) );
  XNOR2_X1 U7147 ( .A(n5661), .B(SI_28_), .ZN(n6202) );
  OR2_X1 U7148 ( .A1(n6218), .A2(n9842), .ZN(n5546) );
  NAND2_X1 U7149 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5548) );
  NOR2_X1 U7150 ( .A1(n5550), .A2(n5548), .ZN(n5651) );
  INV_X1 U7151 ( .A(n5651), .ZN(n9512) );
  INV_X1 U7152 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5549) );
  INV_X1 U7153 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9199) );
  OAI21_X1 U7154 ( .B1(n5550), .B2(n5549), .A(n9199), .ZN(n5551) );
  NAND2_X1 U7155 ( .A1(n9512), .A2(n5551), .ZN(n9200) );
  INV_X1 U7156 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U7157 ( .A1(n5683), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5554) );
  NAND2_X1 U7158 ( .A1(n5682), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5553) );
  OAI211_X1 U7159 ( .C1(n5606), .C2(n5686), .A(n5554), .B(n5553), .ZN(n5555)
         );
  INV_X1 U7160 ( .A(n5555), .ZN(n5556) );
  NAND2_X1 U7161 ( .A1(n9203), .A2(n5558), .ZN(n8027) );
  NAND2_X1 U7162 ( .A1(n5559), .A2(n5560), .ZN(n5586) );
  NAND2_X1 U7163 ( .A1(n5564), .A2(n5563), .ZN(n5561) );
  NAND2_X1 U7164 ( .A1(n5561), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5562) );
  NAND2_X1 U7165 ( .A1(n10009), .A2(P1_B_REG_SCAN_IN), .ZN(n5565) );
  MUX2_X1 U7166 ( .A(P1_B_REG_SCAN_IN), .B(n5565), .S(n7625), .Z(n5572) );
  OAI21_X1 U7167 ( .B1(n5567), .B2(n5566), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5568) );
  NAND2_X1 U7168 ( .A1(n5570), .A2(n5569), .ZN(n7680) );
  INV_X1 U7169 ( .A(n7680), .ZN(n5571) );
  INV_X1 U7170 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U7171 ( .A1(n5692), .A2(n5573), .ZN(n5574) );
  NAND2_X1 U7172 ( .A1(n7680), .A2(n7625), .ZN(n9998) );
  INV_X1 U7173 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U7174 ( .A1(n5581), .A2(n5580), .ZN(n5583) );
  INV_X1 U7175 ( .A(n5559), .ZN(n5577) );
  NAND2_X1 U7176 ( .A1(n5577), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5578) );
  MUX2_X1 U7177 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5578), .S(
        P1_IR_REG_22__SCAN_IN), .Z(n5579) );
  NAND2_X1 U7178 ( .A1(n5579), .A2(n5586), .ZN(n7481) );
  INV_X1 U7179 ( .A(n7481), .ZN(n8159) );
  NAND2_X1 U7180 ( .A1(n4312), .A2(n8159), .ZN(n6870) );
  OR2_X1 U7181 ( .A1(n5581), .A2(n5580), .ZN(n5582) );
  NAND2_X1 U7182 ( .A1(n5583), .A2(n5582), .ZN(n7334) );
  NOR2_X1 U7183 ( .A1(n7680), .A2(n7625), .ZN(n5585) );
  NAND2_X2 U7184 ( .A1(n5585), .A2(n5584), .ZN(n6832) );
  NAND2_X1 U7185 ( .A1(n5586), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5588) );
  XNOR2_X1 U7186 ( .A(n5588), .B(n5587), .ZN(n6328) );
  OAI211_X1 U7187 ( .C1(n6870), .C2(n8106), .A(n6832), .B(n6328), .ZN(n6827)
         );
  NOR2_X1 U7188 ( .A1(n6827), .A2(P1_U3086), .ZN(n5696) );
  NOR4_X1 U7189 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n5592) );
  NOR4_X1 U7190 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5591) );
  NOR4_X1 U7191 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n5590) );
  NOR4_X1 U7192 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n5589) );
  AND4_X1 U7193 ( .A1(n5592), .A2(n5591), .A3(n5590), .A4(n5589), .ZN(n5597)
         );
  NOR2_X1 U7194 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .ZN(
        n9930) );
  NOR4_X1 U7195 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5595) );
  NOR4_X1 U7196 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n5594) );
  NOR4_X1 U7197 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n5593) );
  AND4_X1 U7198 ( .A1(n9930), .A2(n5595), .A3(n5594), .A4(n5593), .ZN(n5596)
         );
  NAND2_X1 U7199 ( .A1(n5597), .A2(n5596), .ZN(n5691) );
  INV_X1 U7200 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n5598) );
  OR2_X1 U7201 ( .A1(n5691), .A2(n5598), .ZN(n5599) );
  NAND2_X1 U7202 ( .A1(n5692), .A2(n5599), .ZN(n6824) );
  NAND2_X1 U7203 ( .A1(n10009), .A2(n7680), .ZN(n9997) );
  NAND4_X1 U7204 ( .A1(n6826), .A2(n5696), .A3(n6824), .A4(n9997), .ZN(n5601)
         );
  INV_X1 U7205 ( .A(n7334), .ZN(n8171) );
  INV_X1 U7206 ( .A(n5693), .ZN(n5600) );
  NAND2_X1 U7207 ( .A1(n6832), .A2(n6637), .ZN(n8158) );
  INV_X1 U7208 ( .A(n8158), .ZN(n9996) );
  INV_X1 U7209 ( .A(n8106), .ZN(n8157) );
  OR2_X1 U7210 ( .A1(n6870), .A2(n8157), .ZN(n5602) );
  NAND2_X1 U7211 ( .A1(n5602), .A2(n6837), .ZN(n7081) );
  NAND2_X1 U7212 ( .A1(n8159), .A2(n8151), .ZN(n5603) );
  AND2_X1 U7213 ( .A1(n8157), .A2(n5603), .ZN(n5604) );
  AND2_X1 U7214 ( .A1(n7334), .A2(n8175), .ZN(n8105) );
  NAND2_X1 U7215 ( .A1(n4312), .A2(n8105), .ZN(n7148) );
  NAND2_X1 U7216 ( .A1(n10095), .A2(n7148), .ZN(n5605) );
  NOR2_X1 U7217 ( .A1(n6837), .A2(n7334), .ZN(n6876) );
  NAND2_X1 U7218 ( .A1(n9663), .A2(n6876), .ZN(n9697) );
  OAI22_X1 U7219 ( .A1(n9200), .A2(n9660), .B1(n5606), .B2(n9663), .ZN(n5611)
         );
  NOR2_X1 U7220 ( .A1(n9835), .A2(n9764), .ZN(n7669) );
  INV_X1 U7221 ( .A(n7669), .ZN(n5607) );
  NOR2_X1 U7222 ( .A1(n9828), .A2(n5607), .ZN(n5608) );
  NAND2_X1 U7223 ( .A1(n10168), .A2(n6901), .ZN(n10146) );
  NAND2_X1 U7224 ( .A1(n10151), .A2(n10180), .ZN(n7106) );
  NOR2_X2 U7225 ( .A1(n10102), .A2(n10224), .ZN(n7387) );
  INV_X1 U7226 ( .A(n9169), .ZN(n7421) );
  NOR2_X4 U7227 ( .A1(n7658), .A2(n9776), .ZN(n7670) );
  INV_X1 U7228 ( .A(n9754), .ZN(n9679) );
  INV_X1 U7229 ( .A(n9806), .ZN(n9612) );
  INV_X1 U7230 ( .A(n5609), .ZN(n9577) );
  NAND2_X1 U7231 ( .A1(n9722), .A2(n9581), .ZN(n9557) );
  NOR2_X2 U7232 ( .A1(n9557), .A2(n9546), .ZN(n9525) );
  OAI211_X1 U7233 ( .C1(n4303), .C2(n4342), .A(n4317), .B(n10148), .ZN(n7844)
         );
  NOR2_X2 U7234 ( .A1(n10130), .A2(n8175), .ZN(n10153) );
  NOR2_X1 U7235 ( .A1(n7844), .A2(n9667), .ZN(n5610) );
  AOI211_X1 U7236 ( .C1(n10142), .C2(n9203), .A(n5611), .B(n5610), .ZN(n5657)
         );
  NOR2_X1 U7237 ( .A1(n7000), .A2(n6901), .ZN(n7157) );
  NAND2_X1 U7238 ( .A1(n8119), .A2(n7157), .ZN(n7156) );
  OR2_X1 U7239 ( .A1(n9402), .A2(n10168), .ZN(n5613) );
  INV_X1 U7240 ( .A(n10145), .ZN(n10137) );
  OR2_X1 U7241 ( .A1(n8050), .A2(n5614), .ZN(n5615) );
  INV_X1 U7242 ( .A(n7949), .ZN(n5616) );
  NAND2_X1 U7243 ( .A1(n9399), .A2(n10185), .ZN(n7951) );
  AND2_X1 U7244 ( .A1(n10124), .A2(n7951), .ZN(n8052) );
  NAND2_X1 U7245 ( .A1(n7071), .A2(n10131), .ZN(n7948) );
  AND2_X1 U7246 ( .A1(n7938), .A2(n7936), .ZN(n8114) );
  INV_X1 U7247 ( .A(n9395), .ZN(n5618) );
  NAND2_X1 U7248 ( .A1(n10101), .A2(n5618), .ZN(n7941) );
  NAND2_X1 U7249 ( .A1(n7969), .A2(n7941), .ZN(n7959) );
  INV_X1 U7250 ( .A(n7940), .ZN(n5617) );
  OR2_X1 U7251 ( .A1(n7959), .A2(n5617), .ZN(n8123) );
  OR2_X1 U7252 ( .A1(n10101), .A2(n5618), .ZN(n7271) );
  NAND2_X1 U7253 ( .A1(n7964), .A2(n7271), .ZN(n7945) );
  NAND2_X1 U7254 ( .A1(n7945), .A2(n7969), .ZN(n5619) );
  NAND2_X1 U7255 ( .A1(n8123), .A2(n5619), .ZN(n8059) );
  AND2_X1 U7256 ( .A1(n7271), .A2(n5620), .ZN(n7956) );
  NAND3_X1 U7257 ( .A1(n7964), .A2(n7956), .A3(n7953), .ZN(n8122) );
  NAND2_X1 U7258 ( .A1(n8059), .A2(n8122), .ZN(n5621) );
  INV_X1 U7259 ( .A(n7972), .ZN(n5622) );
  INV_X1 U7260 ( .A(n8124), .ZN(n7509) );
  INV_X1 U7261 ( .A(n7974), .ZN(n5623) );
  NOR2_X1 U7262 ( .A1(n7530), .A2(n5623), .ZN(n5624) );
  NAND2_X1 U7263 ( .A1(n9143), .A2(n9389), .ZN(n8068) );
  NAND2_X1 U7264 ( .A1(n9776), .A2(n5625), .ZN(n7988) );
  NAND2_X1 U7265 ( .A1(n8068), .A2(n7988), .ZN(n7985) );
  INV_X1 U7266 ( .A(n8064), .ZN(n5626) );
  NOR2_X1 U7267 ( .A1(n7985), .A2(n5626), .ZN(n5627) );
  INV_X1 U7268 ( .A(n9388), .ZN(n5628) );
  OR2_X1 U7269 ( .A1(n9835), .A2(n5628), .ZN(n7991) );
  NAND2_X1 U7270 ( .A1(n9835), .A2(n5628), .ZN(n7989) );
  NAND2_X1 U7271 ( .A1(n7991), .A2(n7989), .ZN(n8130) );
  INV_X1 U7272 ( .A(n9690), .ZN(n9701) );
  INV_X1 U7273 ( .A(n9386), .ZN(n9339) );
  OR2_X1 U7274 ( .A1(n9828), .A2(n9339), .ZN(n9680) );
  NAND2_X1 U7275 ( .A1(n9828), .A2(n9339), .ZN(n7924) );
  NAND2_X1 U7276 ( .A1(n9680), .A2(n7924), .ZN(n7993) );
  INV_X1 U7277 ( .A(n8075), .ZN(n5630) );
  NOR2_X1 U7278 ( .A1(n7993), .A2(n5630), .ZN(n5631) );
  NAND2_X1 U7279 ( .A1(n9699), .A2(n5631), .ZN(n9681) );
  INV_X1 U7280 ( .A(n9385), .ZN(n5632) );
  NAND2_X1 U7281 ( .A1(n9754), .A2(n5632), .ZN(n7925) );
  AND2_X1 U7282 ( .A1(n4384), .A2(n9680), .ZN(n5633) );
  NAND2_X1 U7283 ( .A1(n9681), .A2(n5633), .ZN(n9682) );
  NAND2_X1 U7284 ( .A1(n9682), .A2(n7925), .ZN(n9653) );
  INV_X1 U7285 ( .A(n9384), .ZN(n9340) );
  OR2_X1 U7286 ( .A1(n9822), .A2(n9340), .ZN(n8077) );
  NAND2_X1 U7287 ( .A1(n9822), .A2(n9340), .ZN(n8083) );
  INV_X1 U7288 ( .A(n9383), .ZN(n8108) );
  OR2_X1 U7289 ( .A1(n9816), .A2(n8108), .ZN(n8000) );
  INV_X1 U7290 ( .A(n9381), .ZN(n5634) );
  OR2_X2 U7291 ( .A1(n9806), .A2(n5634), .ZN(n9588) );
  NAND2_X1 U7292 ( .A1(n9806), .A2(n5634), .ZN(n8008) );
  NAND2_X1 U7293 ( .A1(n9588), .A2(n8008), .ZN(n9604) );
  NAND2_X1 U7294 ( .A1(n9816), .A2(n8108), .ZN(n9622) );
  NAND2_X1 U7295 ( .A1(n8003), .A2(n9622), .ZN(n7922) );
  AND2_X1 U7296 ( .A1(n7922), .A2(n8002), .ZN(n9605) );
  NOR2_X1 U7297 ( .A1(n9604), .A2(n9605), .ZN(n5635) );
  OR2_X1 U7298 ( .A1(n9731), .A2(n7803), .ZN(n8044) );
  NAND2_X1 U7299 ( .A1(n9731), .A2(n7803), .ZN(n9563) );
  INV_X1 U7300 ( .A(n9563), .ZN(n8045) );
  INV_X1 U7301 ( .A(n9379), .ZN(n8015) );
  NOR2_X1 U7302 ( .A1(n8045), .A2(n9571), .ZN(n5637) );
  OR2_X1 U7303 ( .A1(n9578), .A2(n8015), .ZN(n9550) );
  OR2_X1 U7304 ( .A1(n9558), .A2(n7684), .ZN(n8047) );
  NAND2_X1 U7305 ( .A1(n9558), .A2(n7684), .ZN(n8020) );
  INV_X1 U7306 ( .A(n9377), .ZN(n5638) );
  INV_X1 U7307 ( .A(n8047), .ZN(n8022) );
  NAND2_X1 U7308 ( .A1(n5643), .A2(n8080), .ZN(n5642) );
  NAND2_X1 U7309 ( .A1(n5642), .A2(n5641), .ZN(n5680) );
  NAND3_X1 U7310 ( .A1(n8139), .A2(n8080), .A3(n5643), .ZN(n5646) );
  NAND2_X1 U7311 ( .A1(n4312), .A2(n8171), .ZN(n5645) );
  NAND2_X1 U7312 ( .A1(n8159), .A2(n8175), .ZN(n5644) );
  NAND2_X1 U7313 ( .A1(n5645), .A2(n5644), .ZN(n10140) );
  NAND3_X1 U7314 ( .A1(n5680), .A2(n5646), .A3(n10140), .ZN(n5654) );
  INV_X1 U7315 ( .A(n6870), .ZN(n8148) );
  INV_X1 U7316 ( .A(n8189), .ZN(n6931) );
  OR2_X1 U7317 ( .A1(n9116), .A2(n9351), .ZN(n5653) );
  INV_X1 U7318 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9511) );
  NAND2_X1 U7319 ( .A1(n5647), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5649) );
  NAND2_X1 U7320 ( .A1(n6239), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5648) );
  OAI211_X1 U7321 ( .C1(n9511), .C2(n5686), .A(n5649), .B(n5648), .ZN(n5650)
         );
  AOI21_X1 U7322 ( .B1(n5651), .B2(n5102), .A(n5650), .ZN(n7222) );
  OR2_X1 U7323 ( .A1(n7222), .A2(n9353), .ZN(n5652) );
  AND2_X1 U7324 ( .A1(n5653), .A2(n5652), .ZN(n9198) );
  MUX2_X1 U7325 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n5659), .Z(n6205) );
  XNOR2_X1 U7326 ( .A(n6205), .B(SI_29_), .ZN(n5665) );
  INV_X1 U7327 ( .A(n5665), .ZN(n5660) );
  AOI21_X1 U7328 ( .B1(n5660), .B2(SI_28_), .A(n5661), .ZN(n5669) );
  INV_X1 U7329 ( .A(SI_28_), .ZN(n5662) );
  INV_X1 U7330 ( .A(n5661), .ZN(n5664) );
  AOI21_X1 U7331 ( .B1(n5665), .B2(n5662), .A(n5664), .ZN(n5668) );
  NAND2_X1 U7332 ( .A1(n5664), .A2(SI_28_), .ZN(n5663) );
  NAND3_X1 U7333 ( .A1(n6203), .A2(n5665), .A3(n5663), .ZN(n5667) );
  NOR2_X1 U7334 ( .A1(n5664), .A2(SI_28_), .ZN(n6208) );
  INV_X1 U7335 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10001) );
  OR2_X1 U7336 ( .A1(n6218), .A2(n10001), .ZN(n5670) );
  OR2_X1 U7337 ( .A1(n5688), .A2(n7222), .ZN(n8043) );
  NAND2_X1 U7338 ( .A1(n5688), .A2(n7222), .ZN(n8097) );
  NAND2_X1 U7339 ( .A1(n9203), .A2(n9375), .ZN(n5674) );
  NAND2_X1 U7340 ( .A1(n5672), .A2(n5671), .ZN(n5679) );
  OR2_X1 U7341 ( .A1(n9203), .A2(n9375), .ZN(n9506) );
  INV_X1 U7342 ( .A(n9506), .ZN(n5673) );
  AND2_X1 U7343 ( .A1(n7481), .A2(n8175), .ZN(n8039) );
  NAND2_X1 U7344 ( .A1(n8039), .A2(n7334), .ZN(n9779) );
  AOI21_X1 U7345 ( .B1(n9508), .B2(n5673), .A(n10195), .ZN(n5676) );
  INV_X1 U7346 ( .A(n5674), .ZN(n9505) );
  NAND2_X1 U7347 ( .A1(n8138), .A2(n9505), .ZN(n5675) );
  NAND3_X1 U7348 ( .A1(n9507), .A2(n8138), .A3(n9506), .ZN(n5677) );
  INV_X1 U7349 ( .A(n10002), .ZN(n10012) );
  AND2_X1 U7350 ( .A1(n10012), .A2(P1_B_REG_SCAN_IN), .ZN(n5681) );
  NOR2_X1 U7351 ( .A1(n9353), .A2(n5681), .ZN(n6244) );
  INV_X1 U7352 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9501) );
  NAND2_X1 U7353 ( .A1(n5682), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U7354 ( .A1(n5683), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5684) );
  OAI211_X1 U7355 ( .C1(n5686), .C2(n9501), .A(n5685), .B(n5684), .ZN(n9374)
         );
  AOI22_X1 U7356 ( .A1(n9375), .A2(n9313), .B1(n6244), .B2(n9374), .ZN(n5687)
         );
  AOI21_X1 U7357 ( .B1(n4317), .B2(n5688), .A(n9693), .ZN(n5689) );
  AND2_X1 U7358 ( .A1(n9497), .A2(n5689), .ZN(n9515) );
  NOR2_X1 U7359 ( .A1(n9516), .A2(n9515), .ZN(n5690) );
  OAI21_X1 U7360 ( .B1(n9995), .B2(P1_D_REG_1__SCAN_IN), .A(n9997), .ZN(n5695)
         );
  NAND2_X1 U7361 ( .A1(n5692), .A2(n5691), .ZN(n5694) );
  NAND4_X1 U7362 ( .A1(n5696), .A2(n5695), .A3(n5694), .A4(n5693), .ZN(n6245)
         );
  NAND2_X1 U7363 ( .A1(n6296), .A2(n10248), .ZN(n5700) );
  NAND2_X1 U7364 ( .A1(n10245), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U7365 ( .A1(n5700), .A2(n5699), .ZN(P1_U3551) );
  NAND2_X1 U7366 ( .A1(n5955), .A2(n6094), .ZN(n6082) );
  INV_X2 U7367 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5701) );
  NAND3_X1 U7368 ( .A1(n6121), .A2(n5702), .A3(n6157), .ZN(n5705) );
  NAND4_X1 U7369 ( .A1(n5837), .A2(n5798), .A3(n5704), .A4(n5703), .ZN(n5854)
         );
  NOR2_X1 U7370 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5707) );
  INV_X1 U7371 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5711) );
  OR2_X2 U7372 ( .A1(n7900), .A2(n5711), .ZN(n5712) );
  XNOR2_X2 U7373 ( .A(n5712), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5718) );
  INV_X1 U7374 ( .A(n5718), .ZN(n8184) );
  NAND2_X1 U7375 ( .A1(n5713), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5715) );
  XNOR2_X2 U7376 ( .A(n5715), .B(n5714), .ZN(n5717) );
  NAND2_X1 U7377 ( .A1(n5772), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5722) );
  AND2_X2 U7378 ( .A1(n5718), .A2(n5717), .ZN(n5728) );
  INV_X1 U7379 ( .A(n5728), .ZN(n5758) );
  INV_X1 U7380 ( .A(n5758), .ZN(n5741) );
  NAND2_X1 U7381 ( .A1(n5741), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U7382 ( .A1(n5773), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5720) );
  NAND2_X1 U7383 ( .A1(n4337), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5719) );
  NAND4_X2 U7384 ( .A1(n5722), .A2(n5721), .A3(n5720), .A4(n5719), .ZN(n6695)
         );
  NAND2_X1 U7385 ( .A1(n6641), .A2(SI_0_), .ZN(n5723) );
  XNOR2_X1 U7386 ( .A(n5723), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9107) );
  NAND2_X1 U7387 ( .A1(n6695), .A2(n9004), .ZN(n7036) );
  NOR2_X1 U7388 ( .A1(n4358), .A2(n5729), .ZN(n5734) );
  INV_X1 U7389 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5730) );
  OR2_X1 U7390 ( .A1(n5731), .A2(n5730), .ZN(n5733) );
  NAND2_X1 U7391 ( .A1(n4337), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5732) );
  INV_X2 U7392 ( .A(n6168), .ZN(n10256) );
  NAND2_X1 U7393 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5735) );
  OR2_X1 U7394 ( .A1(n5746), .A2(n4983), .ZN(n5737) );
  OR2_X1 U7395 ( .A1(n5761), .A2(n6679), .ZN(n5736) );
  OAI21_X1 U7396 ( .B1(n7036), .B2(n10256), .A(n6522), .ZN(n5740) );
  NAND2_X1 U7397 ( .A1(n7036), .A2(n10256), .ZN(n5739) );
  NAND2_X1 U7398 ( .A1(n5740), .A2(n5739), .ZN(n5753) );
  NAND2_X1 U7399 ( .A1(n5773), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5743) );
  NAND2_X1 U7400 ( .A1(n5741), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5742) );
  INV_X1 U7401 ( .A(n5761), .ZN(n5747) );
  OR2_X1 U7402 ( .A1(n5762), .A2(n4448), .ZN(n5749) );
  NAND2_X2 U7403 ( .A1(n5752), .A2(n5754), .ZN(n8450) );
  NAND2_X1 U7404 ( .A1(n5753), .A2(n10255), .ZN(n6983) );
  OR2_X1 U7405 ( .A1(n8627), .A2(n5754), .ZN(n6984) );
  NAND2_X1 U7406 ( .A1(n6983), .A2(n6984), .ZN(n5770) );
  NAND2_X1 U7407 ( .A1(n4337), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5757) );
  NAND2_X1 U7408 ( .A1(n5773), .A2(n8213), .ZN(n5756) );
  NAND2_X1 U7409 ( .A1(n5741), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5759) );
  INV_X1 U7410 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6646) );
  OR2_X1 U7411 ( .A1(n5746), .A2(n6646), .ZN(n5768) );
  NAND2_X1 U7412 ( .A1(n5765), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5764) );
  MUX2_X1 U7413 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5764), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5766) );
  OR2_X1 U7414 ( .A1(n5762), .A2(n6647), .ZN(n5767) );
  NAND2_X1 U7415 ( .A1(n10260), .A2(n10285), .ZN(n8459) );
  NAND2_X1 U7416 ( .A1(n8491), .A2(n8459), .ZN(n6169) );
  NAND2_X1 U7417 ( .A1(n4311), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5778) );
  NAND2_X1 U7418 ( .A1(n5772), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5777) );
  NAND2_X1 U7419 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5774) );
  NAND2_X1 U7420 ( .A1(n5783), .A2(n5774), .ZN(n8292) );
  NAND2_X1 U7421 ( .A1(n5914), .A2(n8292), .ZN(n5776) );
  NAND2_X1 U7422 ( .A1(n8366), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5775) );
  NAND2_X1 U7423 ( .A1(n6651), .A2(n8563), .ZN(n5781) );
  INV_X2 U7424 ( .A(n5762), .ZN(n6368) );
  NAND2_X1 U7425 ( .A1(n5789), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5779) );
  AOI22_X1 U7426 ( .A1(n5976), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n6368), .B2(
        n6434), .ZN(n5780) );
  NAND2_X1 U7427 ( .A1(n5781), .A2(n5780), .ZN(n8289) );
  NAND2_X1 U7428 ( .A1(n8626), .A2(n8289), .ZN(n6170) );
  INV_X4 U7429 ( .A(n5949), .ZN(n6259) );
  NAND2_X1 U7430 ( .A1(n6259), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U7431 ( .A1(n8366), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5787) );
  NAND2_X1 U7432 ( .A1(n5783), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5784) );
  NAND2_X1 U7433 ( .A1(n5803), .A2(n5784), .ZN(n7093) );
  NAND2_X1 U7434 ( .A1(n5914), .A2(n7093), .ZN(n5786) );
  NAND2_X1 U7435 ( .A1(n4311), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5785) );
  AND4_X2 U7436 ( .A1(n5788), .A2(n5787), .A3(n5786), .A4(n5785), .ZN(n7139)
         );
  INV_X2 U7437 ( .A(n7139), .ZN(n8625) );
  OR2_X1 U7438 ( .A1(n6649), .A2(n8565), .ZN(n5794) );
  INV_X1 U7439 ( .A(n5789), .ZN(n5791) );
  NAND2_X1 U7440 ( .A1(n5791), .A2(n5790), .ZN(n5795) );
  NAND2_X1 U7441 ( .A1(n5795), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5792) );
  XNOR2_X1 U7442 ( .A(n5792), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6750) );
  AOI22_X1 U7443 ( .A1(n5976), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6368), .B2(
        n6750), .ZN(n5793) );
  AND2_X1 U7444 ( .A1(n8625), .A2(n10299), .ZN(n7090) );
  NAND2_X1 U7445 ( .A1(n7139), .A2(n6537), .ZN(n7091) );
  NAND2_X1 U7446 ( .A1(n6658), .A2(n8563), .ZN(n5802) );
  NAND2_X1 U7447 ( .A1(n5797), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5796) );
  MUX2_X1 U7448 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5796), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5800) );
  INV_X1 U7449 ( .A(n5797), .ZN(n5799) );
  NAND2_X1 U7450 ( .A1(n5799), .A2(n5798), .ZN(n5821) );
  NAND2_X1 U7451 ( .A1(n5800), .A2(n5821), .ZN(n6660) );
  INV_X1 U7452 ( .A(n6660), .ZN(n8636) );
  AOI22_X1 U7453 ( .A1(n5976), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6368), .B2(
        n8636), .ZN(n5801) );
  NAND2_X1 U7454 ( .A1(n5802), .A2(n5801), .ZN(n7217) );
  NAND2_X1 U7455 ( .A1(n6259), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U7456 ( .A1(n4311), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5807) );
  NAND2_X1 U7457 ( .A1(n5803), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U7458 ( .A1(n5825), .A2(n5804), .ZN(n7216) );
  NAND2_X1 U7459 ( .A1(n5914), .A2(n7216), .ZN(n5806) );
  NAND2_X1 U7460 ( .A1(n8366), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5805) );
  NAND4_X1 U7461 ( .A1(n5808), .A2(n5807), .A3(n5806), .A4(n5805), .ZN(n7354)
         );
  NAND2_X1 U7462 ( .A1(n7217), .A2(n7354), .ZN(n5809) );
  NAND2_X1 U7463 ( .A1(n7137), .A2(n5809), .ZN(n5811) );
  INV_X1 U7464 ( .A(n7217), .ZN(n7029) );
  NAND2_X1 U7465 ( .A1(n7029), .A2(n7206), .ZN(n5810) );
  NAND2_X1 U7466 ( .A1(n6664), .A2(n8563), .ZN(n5814) );
  NAND2_X1 U7467 ( .A1(n5834), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5812) );
  XNOR2_X1 U7468 ( .A(n5812), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6920) );
  AOI22_X1 U7469 ( .A1(n5976), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6368), .B2(
        n6920), .ZN(n5813) );
  NAND2_X1 U7470 ( .A1(n5814), .A2(n5813), .ZN(n7339) );
  NAND2_X1 U7471 ( .A1(n6259), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5820) );
  INV_X1 U7472 ( .A(n4311), .ZN(n6053) );
  INV_X2 U7473 ( .A(n5758), .ZN(n8367) );
  NAND2_X1 U7474 ( .A1(n4311), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5819) );
  NAND2_X1 U7475 ( .A1(n5827), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5816) );
  NAND2_X1 U7476 ( .A1(n5845), .A2(n5816), .ZN(n7290) );
  NAND2_X1 U7477 ( .A1(n5914), .A2(n7290), .ZN(n5818) );
  NAND2_X1 U7478 ( .A1(n8366), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5817) );
  NAND2_X1 U7479 ( .A1(n7339), .A2(n7297), .ZN(n8500) );
  OR2_X1 U7480 ( .A1(n6670), .A2(n8565), .ZN(n5824) );
  NAND2_X1 U7481 ( .A1(n5821), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5822) );
  AOI22_X1 U7482 ( .A1(n5976), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6368), .B2(
        n6445), .ZN(n5823) );
  NAND2_X1 U7483 ( .A1(n5824), .A2(n5823), .ZN(n7350) );
  NAND2_X1 U7484 ( .A1(n6259), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5831) );
  NAND2_X1 U7485 ( .A1(n8366), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U7486 ( .A1(n5825), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5826) );
  NAND2_X1 U7487 ( .A1(n5827), .A2(n5826), .ZN(n7360) );
  NAND2_X1 U7488 ( .A1(n5914), .A2(n7360), .ZN(n5829) );
  NAND2_X1 U7489 ( .A1(n5741), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5828) );
  NAND4_X1 U7490 ( .A1(n5831), .A2(n5830), .A3(n5829), .A4(n5828), .ZN(n8624)
         );
  NOR2_X1 U7491 ( .A1(n7350), .A2(n8624), .ZN(n7248) );
  INV_X1 U7492 ( .A(n8393), .ZN(n5832) );
  AND2_X1 U7493 ( .A1(n7350), .A2(n8624), .ZN(n7246) );
  INV_X1 U7494 ( .A(n7297), .ZN(n7355) );
  AOI22_X1 U7495 ( .A1(n5832), .A2(n7246), .B1(n7355), .B2(n7339), .ZN(n5833)
         );
  NAND2_X1 U7496 ( .A1(n6681), .A2(n8563), .ZN(n5842) );
  NAND2_X1 U7497 ( .A1(n5836), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5835) );
  MUX2_X1 U7498 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5835), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n5839) );
  INV_X1 U7499 ( .A(n5836), .ZN(n5838) );
  NAND2_X1 U7500 ( .A1(n5838), .A2(n5837), .ZN(n5852) );
  NAND2_X1 U7501 ( .A1(n5839), .A2(n5852), .ZN(n6683) );
  OAI22_X1 U7502 ( .A1(n6683), .A2(n5762), .B1(n8363), .B2(n6682), .ZN(n5840)
         );
  INV_X1 U7503 ( .A(n5840), .ZN(n5841) );
  NAND2_X1 U7504 ( .A1(n8368), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U7505 ( .A1(n4311), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U7506 ( .A1(n5845), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5846) );
  NAND2_X1 U7507 ( .A1(n5862), .A2(n5846), .ZN(n7450) );
  NAND2_X1 U7508 ( .A1(n5914), .A2(n7450), .ZN(n5848) );
  NAND2_X1 U7509 ( .A1(n8366), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5847) );
  NAND4_X1 U7510 ( .A1(n5850), .A2(n5849), .A3(n5848), .A4(n5847), .ZN(n7539)
         );
  AND2_X1 U7511 ( .A1(n7451), .A2(n7539), .ZN(n5851) );
  OR2_X1 U7512 ( .A1(n6687), .A2(n8565), .ZN(n5861) );
  NAND2_X1 U7513 ( .A1(n5852), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5853) );
  MUX2_X1 U7514 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5853), .S(
        P2_IR_REG_10__SCAN_IN), .Z(n5859) );
  NOR2_X1 U7515 ( .A1(n5854), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5858) );
  AOI22_X1 U7516 ( .A1(n6459), .A2(n6368), .B1(n5976), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U7517 ( .A1(n6259), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U7518 ( .A1(n8366), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U7519 ( .A1(n5862), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5863) );
  NAND2_X1 U7520 ( .A1(n5873), .A2(n5863), .ZN(n7544) );
  NAND2_X1 U7521 ( .A1(n5914), .A2(n7544), .ZN(n5865) );
  NAND2_X1 U7522 ( .A1(n4311), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5864) );
  NAND4_X1 U7523 ( .A1(n5867), .A2(n5866), .A3(n5865), .A4(n5864), .ZN(n8623)
         );
  NOR2_X1 U7524 ( .A1(n8481), .A2(n8623), .ZN(n5869) );
  NAND2_X1 U7525 ( .A1(n8481), .A2(n8623), .ZN(n5868) );
  NAND2_X1 U7526 ( .A1(n6699), .A2(n8563), .ZN(n5872) );
  NAND2_X1 U7527 ( .A1(n6096), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5870) );
  AOI22_X1 U7528 ( .A1(n5976), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6368), .B2(
        n7367), .ZN(n5871) );
  NAND2_X1 U7529 ( .A1(n4311), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U7530 ( .A1(n8368), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U7531 ( .A1(n5873), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U7532 ( .A1(n5886), .A2(n5874), .ZN(n7597) );
  NAND2_X1 U7533 ( .A1(n5914), .A2(n7597), .ZN(n5876) );
  NAND2_X1 U7534 ( .A1(n8366), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U7535 ( .A1(n8997), .A2(n8484), .ZN(n8505) );
  NAND2_X1 U7536 ( .A1(n7556), .A2(n6559), .ZN(n5880) );
  INV_X1 U7537 ( .A(n8484), .ZN(n8622) );
  NAND2_X1 U7538 ( .A1(n8997), .A2(n8622), .ZN(n5879) );
  INV_X1 U7539 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5881) );
  NAND2_X1 U7540 ( .A1(n6086), .A2(n5881), .ZN(n5894) );
  NAND2_X1 U7541 ( .A1(n5894), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5882) );
  XNOR2_X1 U7542 ( .A(n5882), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7505) );
  AOI22_X1 U7543 ( .A1(n5976), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6368), .B2(
        n7505), .ZN(n5883) );
  NAND2_X1 U7544 ( .A1(n4311), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5891) );
  NAND2_X1 U7545 ( .A1(n6259), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5890) );
  INV_X1 U7546 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5885) );
  NAND2_X1 U7547 ( .A1(n5886), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5887) );
  NAND2_X1 U7548 ( .A1(n5902), .A2(n5887), .ZN(n7886) );
  NAND2_X1 U7549 ( .A1(n6103), .A2(n7886), .ZN(n5889) );
  NAND2_X1 U7550 ( .A1(n8366), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5888) );
  AND2_X1 U7551 ( .A1(n7840), .A2(n8621), .ZN(n5892) );
  INV_X1 U7552 ( .A(n8621), .ZN(n8310) );
  NAND2_X1 U7553 ( .A1(n6176), .A2(n8310), .ZN(n5893) );
  NAND2_X1 U7554 ( .A1(n6819), .A2(n8563), .ZN(n5899) );
  NAND2_X1 U7555 ( .A1(n5908), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5897) );
  XNOR2_X1 U7556 ( .A(n5897), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8662) );
  AOI22_X1 U7557 ( .A1(n5976), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6368), .B2(
        n8662), .ZN(n5898) );
  NAND2_X1 U7558 ( .A1(n4311), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U7559 ( .A1(n6259), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5906) );
  INV_X1 U7560 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U7561 ( .A1(n5902), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U7562 ( .A1(n5912), .A2(n5903), .ZN(n8314) );
  NAND2_X1 U7563 ( .A1(n5914), .A2(n8314), .ZN(n5905) );
  NAND2_X1 U7564 ( .A1(n8366), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5904) );
  NAND4_X1 U7565 ( .A1(n5907), .A2(n5906), .A3(n5905), .A4(n5904), .ZN(n8937)
         );
  NAND2_X1 U7566 ( .A1(n8436), .A2(n8937), .ZN(n7636) );
  NAND2_X1 U7567 ( .A1(n8311), .A2(n8194), .ZN(n7637) );
  OR2_X1 U7568 ( .A1(n6822), .A2(n8565), .ZN(n5911) );
  INV_X1 U7569 ( .A(n5957), .ZN(n5909) );
  NAND2_X1 U7570 ( .A1(n5909), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5929) );
  XNOR2_X1 U7571 ( .A(n5929), .B(P2_IR_REG_14__SCAN_IN), .ZN(n6821) );
  AOI22_X1 U7572 ( .A1(n5976), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6368), .B2(
        n6821), .ZN(n5910) );
  NAND2_X1 U7573 ( .A1(n5912), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U7574 ( .A1(n5924), .A2(n5913), .ZN(n8941) );
  NAND2_X1 U7575 ( .A1(n8941), .A2(n6103), .ZN(n5918) );
  NAND2_X1 U7576 ( .A1(n4311), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U7577 ( .A1(n6259), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5916) );
  NAND2_X1 U7578 ( .A1(n8366), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5915) );
  NAND4_X1 U7579 ( .A1(n5918), .A2(n5917), .A3(n5916), .A4(n5915), .ZN(n8925)
         );
  NOR2_X1 U7580 ( .A1(n9092), .A2(n8925), .ZN(n5919) );
  INV_X1 U7581 ( .A(n8925), .ZN(n6567) );
  NAND2_X1 U7582 ( .A1(n6977), .A2(n8563), .ZN(n5923) );
  INV_X1 U7583 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U7584 ( .A1(n5929), .A2(n6088), .ZN(n5920) );
  NAND2_X1 U7585 ( .A1(n5920), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5921) );
  XNOR2_X1 U7586 ( .A(n5921), .B(P2_IR_REG_15__SCAN_IN), .ZN(n6478) );
  AOI22_X1 U7587 ( .A1(n5976), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6478), .B2(
        n6368), .ZN(n5922) );
  INV_X1 U7588 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8989) );
  NAND2_X1 U7589 ( .A1(n5924), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5925) );
  NAND2_X1 U7590 ( .A1(n5934), .A2(n5925), .ZN(n8928) );
  NAND2_X1 U7591 ( .A1(n8928), .A2(n6103), .ZN(n5927) );
  AOI22_X1 U7592 ( .A1(n6259), .A2(P2_REG0_REG_15__SCAN_IN), .B1(n4311), .B2(
        P2_REG2_REG_15__SCAN_IN), .ZN(n5926) );
  OAI211_X1 U7593 ( .C1(n6262), .C2(n8989), .A(n5927), .B(n5926), .ZN(n8936)
         );
  AND2_X1 U7594 ( .A1(n9085), .A2(n8936), .ZN(n8901) );
  NAND2_X1 U7595 ( .A1(n6992), .A2(n8563), .ZN(n5933) );
  OAI21_X1 U7596 ( .B1(P2_IR_REG_15__SCAN_IN), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7597 ( .A1(n5929), .A2(n5928), .ZN(n5930) );
  OR2_X1 U7598 ( .A1(n5930), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5939) );
  NAND2_X1 U7599 ( .A1(n5930), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5931) );
  AND2_X1 U7600 ( .A1(n5939), .A2(n5931), .ZN(n6994) );
  AOI22_X1 U7601 ( .A1(n5976), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6994), .B2(
        n6368), .ZN(n5932) );
  NAND2_X1 U7602 ( .A1(n5934), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5935) );
  NAND2_X1 U7603 ( .A1(n5945), .A2(n5935), .ZN(n8917) );
  NAND2_X1 U7604 ( .A1(n8917), .A2(n6103), .ZN(n5938) );
  AOI22_X1 U7605 ( .A1(n8366), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n6259), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n5937) );
  NAND2_X1 U7606 ( .A1(n4311), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5936) );
  AND2_X1 U7607 ( .A1(n8986), .A2(n8924), .ZN(n5953) );
  NAND2_X1 U7608 ( .A1(n7087), .A2(n8563), .ZN(n5942) );
  NAND2_X1 U7609 ( .A1(n5939), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5940) );
  XNOR2_X1 U7610 ( .A(n5940), .B(P2_IR_REG_17__SCAN_IN), .ZN(n6487) );
  AOI22_X1 U7611 ( .A1(n6487), .A2(n6368), .B1(n5976), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n5941) );
  INV_X1 U7612 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5943) );
  NAND2_X1 U7613 ( .A1(n5945), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U7614 ( .A1(n5964), .A2(n5946), .ZN(n8898) );
  NAND2_X1 U7615 ( .A1(n8898), .A2(n6103), .ZN(n5952) );
  INV_X1 U7616 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9943) );
  NAND2_X1 U7617 ( .A1(n4311), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U7618 ( .A1(n8366), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5947) );
  OAI211_X1 U7619 ( .C1(n5949), .C2(n9943), .A(n5948), .B(n5947), .ZN(n5950)
         );
  INV_X1 U7620 ( .A(n5950), .ZN(n5951) );
  XNOR2_X1 U7621 ( .A(n9073), .B(n8911), .ZN(n8890) );
  OR2_X1 U7622 ( .A1(n8986), .A2(n8892), .ZN(n8528) );
  NAND2_X1 U7623 ( .A1(n8986), .A2(n8892), .ZN(n8518) );
  INV_X1 U7624 ( .A(n8915), .ZN(n6187) );
  OR2_X1 U7625 ( .A1(n9085), .A2(n8936), .ZN(n8903) );
  AND2_X1 U7626 ( .A1(n6187), .A2(n8903), .ZN(n8902) );
  OR2_X1 U7627 ( .A1(n5953), .A2(n8902), .ZN(n8887) );
  AND2_X1 U7628 ( .A1(n8890), .A2(n8887), .ZN(n8868) );
  OR2_X1 U7629 ( .A1(n7143), .A2(n8565), .ZN(n5963) );
  NOR2_X1 U7630 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5954) );
  AND2_X1 U7631 ( .A1(n5955), .A2(n5954), .ZN(n5956) );
  INV_X1 U7632 ( .A(n5960), .ZN(n5958) );
  NAND2_X1 U7633 ( .A1(n5958), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5959) );
  MUX2_X1 U7634 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5959), .S(
        P2_IR_REG_18__SCAN_IN), .Z(n5961) );
  INV_X1 U7635 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U7636 ( .A1(n5960), .A2(n6090), .ZN(n5974) );
  NAND2_X1 U7637 ( .A1(n5961), .A2(n5974), .ZN(n8742) );
  INV_X1 U7638 ( .A(n8742), .ZN(n6501) );
  AOI22_X1 U7639 ( .A1(n6368), .A2(n6501), .B1(n5976), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7640 ( .A1(n5964), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U7641 ( .A1(n5979), .A2(n5965), .ZN(n8878) );
  NAND2_X1 U7642 ( .A1(n8878), .A2(n6103), .ZN(n5970) );
  INV_X1 U7643 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8981) );
  NAND2_X1 U7644 ( .A1(n8368), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5967) );
  NAND2_X1 U7645 ( .A1(n4311), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5966) );
  OAI211_X1 U7646 ( .C1(n6262), .C2(n8981), .A(n5967), .B(n5966), .ZN(n5968)
         );
  INV_X1 U7647 ( .A(n5968), .ZN(n5969) );
  NAND2_X1 U7648 ( .A1(n8881), .A2(n8893), .ZN(n5971) );
  AND2_X1 U7649 ( .A1(n8868), .A2(n5971), .ZN(n5973) );
  INV_X1 U7650 ( .A(n5971), .ZN(n5972) );
  INV_X1 U7651 ( .A(n8911), .ZN(n8327) );
  NAND2_X1 U7652 ( .A1(n9073), .A2(n8327), .ZN(n8869) );
  INV_X1 U7653 ( .A(n8893), .ZN(n6817) );
  NAND2_X1 U7654 ( .A1(n8980), .A2(n6817), .ZN(n8853) );
  NAND2_X1 U7655 ( .A1(n7243), .A2(n8563), .ZN(n5978) );
  AOI22_X1 U7656 ( .A1(n8739), .A2(n6368), .B1(n5976), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n5977) );
  NAND2_X1 U7657 ( .A1(n5979), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5980) );
  NAND2_X1 U7658 ( .A1(n5999), .A2(n5980), .ZN(n8863) );
  INV_X1 U7659 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8977) );
  NAND2_X1 U7660 ( .A1(n4311), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U7661 ( .A1(n6259), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5981) );
  OAI211_X1 U7662 ( .C1(n8977), .C2(n6262), .A(n5982), .B(n5981), .ZN(n5983)
         );
  AOI21_X1 U7663 ( .B1(n8863), .B2(n5914), .A(n5983), .ZN(n8873) );
  INV_X1 U7664 ( .A(n8873), .ZN(n8847) );
  NAND2_X1 U7665 ( .A1(n8976), .A2(n8847), .ZN(n5984) );
  AND2_X1 U7666 ( .A1(n8853), .A2(n5984), .ZN(n5986) );
  INV_X1 U7667 ( .A(n5984), .ZN(n5985) );
  NAND2_X1 U7668 ( .A1(n8976), .A2(n8873), .ZN(n8535) );
  NAND2_X1 U7669 ( .A1(n8536), .A2(n8535), .ZN(n8855) );
  NAND2_X1 U7670 ( .A1(n7397), .A2(n8563), .ZN(n5988) );
  OR2_X1 U7671 ( .A1(n8363), .A2(n7398), .ZN(n5987) );
  INV_X1 U7672 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5989) );
  INV_X1 U7673 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5991) );
  INV_X1 U7674 ( .A(n5992), .ZN(n6001) );
  NAND2_X1 U7675 ( .A1(n6001), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5993) );
  NAND2_X1 U7676 ( .A1(n6010), .A2(n5993), .ZN(n8836) );
  INV_X1 U7677 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8969) );
  NAND2_X1 U7678 ( .A1(n4311), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U7679 ( .A1(n6259), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5994) );
  OAI211_X1 U7680 ( .C1(n8969), .C2(n6262), .A(n5995), .B(n5994), .ZN(n5996)
         );
  NAND2_X1 U7681 ( .A1(n9054), .A2(n8301), .ZN(n8545) );
  NAND2_X1 U7682 ( .A1(n7303), .A2(n8563), .ZN(n5998) );
  OR2_X1 U7683 ( .A1(n8363), .A2(n9854), .ZN(n5997) );
  NAND2_X1 U7684 ( .A1(n5999), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U7685 ( .A1(n6001), .A2(n6000), .ZN(n8850) );
  NAND2_X1 U7686 ( .A1(n8850), .A2(n6103), .ZN(n6006) );
  INV_X1 U7687 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8972) );
  NAND2_X1 U7688 ( .A1(n4311), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U7689 ( .A1(n8368), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6002) );
  OAI211_X1 U7690 ( .C1(n8972), .C2(n6262), .A(n6003), .B(n6002), .ZN(n6004)
         );
  INV_X1 U7691 ( .A(n6004), .ZN(n6005) );
  NAND2_X1 U7692 ( .A1(n6006), .A2(n6005), .ZN(n8833) );
  NAND2_X1 U7693 ( .A1(n9060), .A2(n8858), .ZN(n8825) );
  NAND2_X1 U7694 ( .A1(n8543), .A2(n8825), .ZN(n8844) );
  NAND2_X1 U7695 ( .A1(n8828), .A2(n8844), .ZN(n6007) );
  NOR2_X1 U7696 ( .A1(n9060), .A2(n8833), .ZN(n8829) );
  NOR2_X1 U7697 ( .A1(n9054), .A2(n8846), .ZN(n8814) );
  NAND2_X1 U7698 ( .A1(n7480), .A2(n8563), .ZN(n6009) );
  OR2_X1 U7699 ( .A1(n8363), .A2(n7485), .ZN(n6008) );
  NAND2_X1 U7700 ( .A1(n6010), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7701 ( .A1(n6018), .A2(n6011), .ZN(n8822) );
  INV_X1 U7702 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8966) );
  NAND2_X1 U7703 ( .A1(n4311), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6013) );
  NAND2_X1 U7704 ( .A1(n6259), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6012) );
  OAI211_X1 U7705 ( .C1(n8966), .C2(n6262), .A(n6013), .B(n6012), .ZN(n6014)
         );
  NAND2_X1 U7706 ( .A1(n9048), .A2(n8243), .ZN(n8550) );
  OR2_X1 U7707 ( .A1(n9048), .A2(n8832), .ZN(n6015) );
  NAND2_X1 U7708 ( .A1(n7576), .A2(n8563), .ZN(n6017) );
  OR2_X1 U7709 ( .A1(n8363), .A2(n7579), .ZN(n6016) );
  NAND2_X1 U7710 ( .A1(n6018), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U7711 ( .A1(n6030), .A2(n6019), .ZN(n8808) );
  NAND2_X1 U7712 ( .A1(n8808), .A2(n6103), .ZN(n6024) );
  INV_X1 U7713 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9952) );
  NAND2_X1 U7714 ( .A1(n6259), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6021) );
  NAND2_X1 U7715 ( .A1(n4311), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6020) );
  OAI211_X1 U7716 ( .C1(n6262), .C2(n9952), .A(n6021), .B(n6020), .ZN(n6022)
         );
  INV_X1 U7717 ( .A(n6022), .ZN(n6023) );
  NAND2_X1 U7718 ( .A1(n9042), .A2(n8819), .ZN(n6025) );
  OR2_X1 U7719 ( .A1(n9042), .A2(n8819), .ZN(n6026) );
  NAND2_X1 U7720 ( .A1(n7621), .A2(n8563), .ZN(n6028) );
  OR2_X1 U7721 ( .A1(n8363), .A2(n7622), .ZN(n6027) );
  INV_X1 U7722 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9846) );
  NAND2_X1 U7723 ( .A1(n6030), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7724 ( .A1(n6039), .A2(n6031), .ZN(n8798) );
  NAND2_X1 U7725 ( .A1(n8798), .A2(n6103), .ZN(n6036) );
  INV_X1 U7726 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8961) );
  NAND2_X1 U7727 ( .A1(n8368), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6033) );
  NAND2_X1 U7728 ( .A1(n5741), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6032) );
  OAI211_X1 U7729 ( .C1(n6262), .C2(n8961), .A(n6033), .B(n6032), .ZN(n6034)
         );
  INV_X1 U7730 ( .A(n6034), .ZN(n6035) );
  NAND2_X1 U7731 ( .A1(n9036), .A2(n8783), .ZN(n8422) );
  NAND2_X1 U7732 ( .A1(n8555), .A2(n8422), .ZN(n8794) );
  NAND2_X1 U7733 ( .A1(n7663), .A2(n8563), .ZN(n6038) );
  OR2_X1 U7734 ( .A1(n8363), .A2(n7664), .ZN(n6037) );
  NAND2_X1 U7735 ( .A1(n6039), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7736 ( .A1(n8785), .A2(n6103), .ZN(n6045) );
  INV_X1 U7737 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8958) );
  NAND2_X1 U7738 ( .A1(n4311), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6042) );
  NAND2_X1 U7739 ( .A1(n8368), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6041) );
  OAI211_X1 U7740 ( .C1(n8958), .C2(n6262), .A(n6042), .B(n6041), .ZN(n6043)
         );
  INV_X1 U7741 ( .A(n6043), .ZN(n6044) );
  OR2_X1 U7742 ( .A1(n9030), .A2(n4568), .ZN(n6046) );
  NAND2_X1 U7743 ( .A1(n7678), .A2(n8563), .ZN(n6048) );
  OR2_X1 U7744 ( .A1(n8363), .A2(n9102), .ZN(n6047) );
  NAND2_X1 U7745 ( .A1(n6049), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U7746 ( .A1(n6063), .A2(n6050), .ZN(n8776) );
  NAND2_X1 U7747 ( .A1(n8776), .A2(n5914), .ZN(n6056) );
  INV_X1 U7748 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9904) );
  NAND2_X1 U7749 ( .A1(n8366), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U7750 ( .A1(n6259), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6051) );
  OAI211_X1 U7751 ( .C1(n6053), .C2(n9904), .A(n6052), .B(n6051), .ZN(n6054)
         );
  INV_X1 U7752 ( .A(n6054), .ZN(n6055) );
  NOR2_X1 U7753 ( .A1(n9024), .A2(n8767), .ZN(n6057) );
  NAND2_X1 U7754 ( .A1(n9024), .A2(n8767), .ZN(n6058) );
  NAND2_X1 U7755 ( .A1(n9098), .A2(n8563), .ZN(n6060) );
  OR2_X1 U7756 ( .A1(n8363), .A2(n9099), .ZN(n6059) );
  INV_X1 U7757 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7758 ( .A1(n6063), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7759 ( .A1(n6074), .A2(n6064), .ZN(n8769) );
  NAND2_X1 U7760 ( .A1(n8769), .A2(n6103), .ZN(n6069) );
  INV_X1 U7761 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8953) );
  NAND2_X1 U7762 ( .A1(n6259), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6066) );
  NAND2_X1 U7763 ( .A1(n4311), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6065) );
  OAI211_X1 U7764 ( .C1(n8953), .C2(n6262), .A(n6066), .B(n6065), .ZN(n6067)
         );
  INV_X1 U7765 ( .A(n6067), .ZN(n6068) );
  AND2_X1 U7766 ( .A1(n9018), .A2(n8775), .ZN(n6071) );
  OR2_X1 U7767 ( .A1(n9018), .A2(n8775), .ZN(n6070) );
  NAND2_X1 U7768 ( .A1(n8186), .A2(n8563), .ZN(n6073) );
  OR2_X1 U7769 ( .A1(n8363), .A2(n8188), .ZN(n6072) );
  NAND2_X1 U7770 ( .A1(n6074), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7771 ( .A1(n7916), .A2(n6075), .ZN(n8232) );
  NAND2_X1 U7772 ( .A1(n8232), .A2(n6103), .ZN(n6080) );
  INV_X1 U7773 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U7774 ( .A1(n5728), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U7775 ( .A1(n6259), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6076) );
  OAI211_X1 U7776 ( .C1(n6509), .C2(n6262), .A(n6077), .B(n6076), .ZN(n6078)
         );
  INV_X1 U7777 ( .A(n6078), .ZN(n6079) );
  NAND2_X1 U7778 ( .A1(n8576), .A2(n8582), .ZN(n6251) );
  INV_X1 U7779 ( .A(n6096), .ZN(n6086) );
  NAND2_X1 U7780 ( .A1(n6086), .A2(n4942), .ZN(n6115) );
  NAND2_X1 U7781 ( .A1(n6115), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7782 ( .A1(n8739), .A2(n8603), .ZN(n6102) );
  INV_X1 U7783 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6089) );
  AND3_X1 U7784 ( .A1(n6090), .A2(n6089), .A3(n6088), .ZN(n6093) );
  NOR2_X1 U7785 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n6092) );
  NAND4_X1 U7786 ( .A1(n6094), .A2(n6093), .A3(n6092), .A4(n6091), .ZN(n6095)
         );
  INV_X1 U7787 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6100) );
  NAND2_X1 U7788 ( .A1(n6099), .A2(n6100), .ZN(n6097) );
  NAND2_X1 U7789 ( .A1(n6097), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6098) );
  INV_X1 U7790 ( .A(n8613), .ZN(n8610) );
  NAND2_X1 U7791 ( .A1(n8440), .A2(n8610), .ZN(n6101) );
  NAND2_X2 U7792 ( .A1(n6102), .A2(n6101), .ZN(n10257) );
  INV_X1 U7793 ( .A(n10257), .ZN(n8871) );
  INV_X1 U7794 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n7915) );
  NAND2_X1 U7795 ( .A1(n8368), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U7796 ( .A1(n8366), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6105) );
  OAI211_X1 U7797 ( .C1(n7915), .C2(n6053), .A(n6106), .B(n6105), .ZN(n6107)
         );
  INV_X1 U7798 ( .A(n6107), .ZN(n6108) );
  INV_X1 U7799 ( .A(n6498), .ZN(n6494) );
  INV_X1 U7800 ( .A(n6472), .ZN(n8744) );
  NAND2_X1 U7801 ( .A1(n6494), .A2(n8744), .ZN(n6109) );
  NAND2_X1 U7802 ( .A1(n5762), .A2(n6109), .ZN(n6614) );
  NAND2_X1 U7803 ( .A1(n6614), .A2(n8591), .ZN(n8910) );
  INV_X1 U7804 ( .A(n6614), .ZN(n6613) );
  INV_X2 U7805 ( .A(n8440), .ZN(n8445) );
  INV_X1 U7806 ( .A(n8603), .ZN(n7483) );
  NAND2_X1 U7807 ( .A1(n8445), .A2(n7483), .ZN(n10302) );
  NOR2_X1 U7808 ( .A1(n6313), .A2(n6114), .ZN(n6507) );
  OAI21_X2 U7809 ( .B1(n6115), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6156) );
  NAND2_X1 U7810 ( .A1(n6156), .A2(n6157), .ZN(n6127) );
  NAND2_X1 U7811 ( .A1(n6127), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6137) );
  INV_X1 U7812 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U7813 ( .A1(n6137), .A2(n6136), .ZN(n6138) );
  NAND2_X1 U7814 ( .A1(n6138), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6117) );
  INV_X1 U7815 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6116) );
  XNOR2_X1 U7816 ( .A(n6117), .B(n6116), .ZN(n7665) );
  INV_X1 U7817 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U7818 ( .A1(n7665), .A2(n9103), .ZN(n6133) );
  INV_X1 U7819 ( .A(n9103), .ZN(n6130) );
  INV_X1 U7820 ( .A(n6127), .ZN(n6125) );
  INV_X1 U7821 ( .A(P2_B_REG_SCAN_IN), .ZN(n6122) );
  AOI22_X1 U7822 ( .A1(n6121), .A2(P2_B_REG_SCAN_IN), .B1(
        P2_IR_REG_24__SCAN_IN), .B2(n6122), .ZN(n6123) );
  INV_X1 U7823 ( .A(n6123), .ZN(n6124) );
  NAND2_X1 U7824 ( .A1(n6125), .A2(n6124), .ZN(n6129) );
  XNOR2_X1 U7825 ( .A(P2_IR_REG_24__SCAN_IN), .B(P2_B_REG_SCAN_IN), .ZN(n6126)
         );
  NAND3_X1 U7826 ( .A1(n6127), .A2(P2_IR_REG_25__SCAN_IN), .A3(n6126), .ZN(
        n6128) );
  INV_X1 U7827 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7828 ( .A1(n6135), .A2(n6131), .ZN(n6132) );
  NAND2_X1 U7829 ( .A1(n6133), .A2(n6132), .ZN(n6656) );
  INV_X1 U7830 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U7831 ( .A1(n6135), .A2(n6134), .ZN(n6141) );
  OR2_X1 U7832 ( .A1(n6137), .A2(n6136), .ZN(n6139) );
  NAND2_X1 U7833 ( .A1(n6139), .A2(n6138), .ZN(n6153) );
  NAND2_X1 U7834 ( .A1(n6153), .A2(n9103), .ZN(n6140) );
  AND2_X2 U7835 ( .A1(n6141), .A2(n6140), .ZN(n6514) );
  INV_X1 U7836 ( .A(n6514), .ZN(n6142) );
  NOR2_X1 U7837 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .ZN(
        n6146) );
  NOR4_X1 U7838 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n6145) );
  NOR4_X1 U7839 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6144) );
  NOR4_X1 U7840 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6143) );
  NAND4_X1 U7841 ( .A1(n6146), .A2(n6145), .A3(n6144), .A4(n6143), .ZN(n6152)
         );
  NOR4_X1 U7842 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6150) );
  NOR4_X1 U7843 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6149) );
  NOR4_X1 U7844 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6148) );
  NOR4_X1 U7845 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6147) );
  NAND4_X1 U7846 ( .A1(n6150), .A2(n6149), .A3(n6148), .A4(n6147), .ZN(n6151)
         );
  OAI21_X1 U7847 ( .B1(n6152), .B2(n6151), .A(n6135), .ZN(n6285) );
  INV_X1 U7848 ( .A(n6285), .ZN(n6164) );
  OR2_X1 U7849 ( .A1(n6286), .A2(n6164), .ZN(n6616) );
  INV_X1 U7850 ( .A(n7665), .ZN(n6155) );
  NOR2_X1 U7851 ( .A1(n6153), .A2(n9103), .ZN(n6154) );
  NAND2_X1 U7852 ( .A1(n6155), .A2(n6154), .ZN(n6617) );
  XNOR2_X1 U7853 ( .A(n6156), .B(n6157), .ZN(n7577) );
  AND2_X1 U7854 ( .A1(n7577), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6158) );
  INV_X1 U7855 ( .A(n6662), .ZN(n6657) );
  NOR2_X1 U7856 ( .A1(n6616), .A2(n6657), .ZN(n6610) );
  OR2_X1 U7857 ( .A1(n6518), .A2(n8584), .ZN(n6625) );
  NAND2_X1 U7858 ( .A1(n8610), .A2(n8603), .ZN(n6160) );
  NOR2_X1 U7859 ( .A1(n6160), .A2(n8440), .ZN(n6161) );
  NAND2_X1 U7860 ( .A1(n8739), .A2(n6161), .ZN(n6619) );
  NAND2_X1 U7861 ( .A1(n6625), .A2(n6619), .ZN(n6162) );
  NAND2_X1 U7862 ( .A1(n6610), .A2(n6162), .ZN(n6167) );
  NAND2_X1 U7863 ( .A1(n8739), .A2(n8613), .ZN(n6307) );
  NAND2_X1 U7864 ( .A1(n6307), .A2(n10300), .ZN(n10251) );
  AND2_X1 U7865 ( .A1(n8584), .A2(n10302), .ZN(n6163) );
  NAND2_X1 U7866 ( .A1(n6619), .A2(n6163), .ZN(n6602) );
  AND2_X1 U7867 ( .A1(n10251), .A2(n6602), .ZN(n6622) );
  NOR2_X1 U7868 ( .A1(n6514), .A2(n6164), .ZN(n6165) );
  AND2_X1 U7869 ( .A1(n6165), .A2(n6656), .ZN(n6626) );
  NAND2_X1 U7870 ( .A1(n6626), .A2(n6662), .ZN(n6612) );
  AND2_X2 U7871 ( .A1(n6167), .A2(n6166), .ZN(n10310) );
  INV_X2 U7872 ( .A(n10310), .ZN(n10308) );
  OR2_X1 U7873 ( .A1(n6507), .A2(n10310), .ZN(n6201) );
  NAND2_X1 U7874 ( .A1(n6168), .A2(n6522), .ZN(n8447) );
  NAND2_X2 U7875 ( .A1(n10256), .A2(n7044), .ZN(n8446) );
  INV_X1 U7876 ( .A(n9004), .ZN(n6696) );
  NOR2_X1 U7877 ( .A1(n6695), .A2(n6696), .ZN(n6521) );
  INV_X1 U7878 ( .A(n10255), .ZN(n8385) );
  NAND2_X1 U7879 ( .A1(n10250), .A2(n8385), .ZN(n10249) );
  NAND2_X1 U7880 ( .A1(n6981), .A2(n8491), .ZN(n7061) );
  NAND2_X1 U7881 ( .A1(n4343), .A2(n6170), .ZN(n8457) );
  NAND2_X1 U7882 ( .A1(n7061), .A2(n8457), .ZN(n6171) );
  INV_X1 U7883 ( .A(n8289), .ZN(n10290) );
  OR2_X1 U7884 ( .A1(n8626), .A2(n10290), .ZN(n8461) );
  NAND2_X1 U7885 ( .A1(n6171), .A2(n8461), .ZN(n7089) );
  NAND2_X1 U7886 ( .A1(n6537), .A2(n8625), .ZN(n8464) );
  NAND2_X1 U7887 ( .A1(n7217), .A2(n7206), .ZN(n8466) );
  NAND2_X1 U7888 ( .A1(n7139), .A2(n10299), .ZN(n7135) );
  NAND2_X1 U7889 ( .A1(n8466), .A2(n7135), .ZN(n8460) );
  AND2_X1 U7890 ( .A1(n7350), .A2(n7265), .ZN(n8501) );
  NOR2_X1 U7891 ( .A1(n8460), .A2(n8501), .ZN(n6172) );
  NAND2_X1 U7892 ( .A1(n7029), .A2(n7354), .ZN(n8465) );
  OR2_X1 U7893 ( .A1(n7350), .A2(n7265), .ZN(n8469) );
  OAI211_X1 U7894 ( .C1(n8501), .C2(n8465), .A(n8470), .B(n8469), .ZN(n6173)
         );
  NAND2_X1 U7895 ( .A1(n7451), .A2(n7263), .ZN(n8503) );
  NAND2_X1 U7896 ( .A1(n8477), .A2(n8503), .ZN(n8396) );
  NOR2_X1 U7897 ( .A1(n8481), .A2(n8482), .ZN(n8476) );
  NAND2_X1 U7898 ( .A1(n8481), .A2(n8482), .ZN(n8504) );
  NAND2_X1 U7899 ( .A1(n6176), .A2(n8621), .ZN(n8511) );
  AND2_X1 U7900 ( .A1(n8399), .A2(n8511), .ZN(n7643) );
  NOR2_X1 U7901 ( .A1(n8436), .A2(n8194), .ZN(n6181) );
  INV_X1 U7902 ( .A(n6181), .ZN(n6177) );
  AND2_X1 U7903 ( .A1(n7643), .A2(n6177), .ZN(n6178) );
  NAND2_X1 U7904 ( .A1(n7561), .A2(n6178), .ZN(n6184) );
  NAND2_X1 U7905 ( .A1(n7840), .A2(n8310), .ZN(n8510) );
  INV_X1 U7906 ( .A(n8505), .ZN(n6179) );
  NAND2_X1 U7907 ( .A1(n8436), .A2(n8194), .ZN(n6180) );
  AND2_X1 U7908 ( .A1(n7646), .A2(n6180), .ZN(n6182) );
  NAND2_X1 U7909 ( .A1(n6184), .A2(n6183), .ZN(n8943) );
  NAND2_X1 U7910 ( .A1(n8933), .A2(n8925), .ZN(n8431) );
  NAND2_X1 U7911 ( .A1(n9092), .A2(n6567), .ZN(n8432) );
  INV_X1 U7912 ( .A(n8936), .ZN(n8909) );
  AND2_X1 U7913 ( .A1(n9085), .A2(n8909), .ZN(n8526) );
  OR2_X1 U7914 ( .A1(n9085), .A2(n8909), .ZN(n8516) );
  NAND2_X1 U7915 ( .A1(n6186), .A2(n8516), .ZN(n8916) );
  OAI21_X2 U7916 ( .B1(n8916), .B2(n6187), .A(n8518), .ZN(n8886) );
  INV_X1 U7917 ( .A(n8890), .ZN(n8519) );
  NAND2_X1 U7918 ( .A1(n9073), .A2(n8911), .ZN(n8520) );
  NAND2_X1 U7919 ( .A1(n8980), .A2(n8893), .ZN(n8521) );
  NAND2_X1 U7920 ( .A1(n8532), .A2(n8521), .ZN(n8876) );
  INV_X1 U7921 ( .A(n8876), .ZN(n6188) );
  INV_X1 U7922 ( .A(n8855), .ZN(n8859) );
  AND2_X1 U7923 ( .A1(n8545), .A2(n8825), .ZN(n8541) );
  INV_X1 U7924 ( .A(n9042), .ZN(n6189) );
  NAND2_X1 U7925 ( .A1(n9042), .A2(n8321), .ZN(n8790) );
  AND2_X1 U7926 ( .A1(n8422), .A2(n8790), .ZN(n8553) );
  NAND2_X1 U7927 ( .A1(n9018), .A2(n8234), .ZN(n8562) );
  NAND2_X1 U7928 ( .A1(n6193), .A2(n8561), .ZN(n6252) );
  NAND2_X1 U7929 ( .A1(n6625), .A2(n10302), .ZN(n6947) );
  NAND2_X1 U7930 ( .A1(n6194), .A2(n8603), .ZN(n6282) );
  AND2_X1 U7931 ( .A1(n6518), .A2(n6282), .ZN(n6195) );
  NAND2_X1 U7932 ( .A1(n10265), .A2(n10304), .ZN(n10293) );
  INV_X1 U7933 ( .A(n10293), .ZN(n10295) );
  INV_X1 U7934 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6196) );
  NAND2_X1 U7935 ( .A1(n6201), .A2(n6200), .ZN(P2_U3455) );
  INV_X1 U7936 ( .A(n6208), .ZN(n6204) );
  NAND2_X1 U7937 ( .A1(n6210), .A2(n6204), .ZN(n6206) );
  INV_X1 U7938 ( .A(n6205), .ZN(n6209) );
  NAND2_X1 U7939 ( .A1(n6206), .A2(n6209), .ZN(n6207) );
  NOR2_X1 U7940 ( .A1(n6209), .A2(n6208), .ZN(n6211) );
  NAND2_X1 U7941 ( .A1(n6211), .A2(n6210), .ZN(n6226) );
  NAND2_X1 U7942 ( .A1(n6223), .A2(n6226), .ZN(n6216) );
  INV_X1 U7943 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7912) );
  INV_X1 U7944 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8357) );
  MUX2_X1 U7945 ( .A(n7912), .B(n8357), .S(n6641), .Z(n6213) );
  INV_X1 U7946 ( .A(SI_30_), .ZN(n6212) );
  NAND2_X1 U7947 ( .A1(n6213), .A2(n6212), .ZN(n6227) );
  INV_X1 U7948 ( .A(n6213), .ZN(n6214) );
  NAND2_X1 U7949 ( .A1(n6214), .A2(SI_30_), .ZN(n6224) );
  NAND2_X1 U7950 ( .A1(n6227), .A2(n6224), .ZN(n6215) );
  NAND2_X1 U7951 ( .A1(n7910), .A2(n6217), .ZN(n6220) );
  OR2_X1 U7952 ( .A1(n6218), .A2(n7912), .ZN(n6219) );
  NAND2_X2 U7953 ( .A1(n6220), .A2(n6219), .ZN(n9503) );
  INV_X1 U7954 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6235) );
  MUX2_X1 U7955 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6641), .Z(n6222) );
  INV_X1 U7956 ( .A(SI_31_), .ZN(n6221) );
  XNOR2_X1 U7957 ( .A(n6222), .B(n6221), .ZN(n6225) );
  NAND2_X1 U7958 ( .A1(n6225), .A2(n6227), .ZN(n6234) );
  INV_X1 U7959 ( .A(n6225), .ZN(n6229) );
  NAND4_X1 U7960 ( .A1(n6223), .A2(n6224), .A3(n6226), .A4(n6229), .ZN(n6233)
         );
  NAND3_X1 U7961 ( .A1(n6226), .A2(n6225), .A3(n6224), .ZN(n6231) );
  INV_X1 U7962 ( .A(n6227), .ZN(n6228) );
  XNOR2_X1 U7963 ( .A(n6229), .B(n6228), .ZN(n6230) );
  NAND2_X1 U7964 ( .A1(n6231), .A2(n6230), .ZN(n6232) );
  MUX2_X1 U7965 ( .A(n6235), .B(n8361), .S(n5659), .Z(n6237) );
  XNOR2_X1 U7966 ( .A(n9498), .B(n8169), .ZN(n6238) );
  NAND2_X1 U7967 ( .A1(n6238), .A2(n10148), .ZN(n7909) );
  NAND2_X1 U7968 ( .A1(n6239), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U7969 ( .A1(n5682), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6242) );
  NAND2_X1 U7970 ( .A1(n6240), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6241) );
  NAND3_X1 U7971 ( .A1(n6243), .A2(n6242), .A3(n6241), .ZN(n9373) );
  NAND2_X1 U7972 ( .A1(n9373), .A2(n6244), .ZN(n9709) );
  INV_X1 U7973 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9867) );
  INV_X1 U7974 ( .A(n6245), .ZN(n6246) );
  NAND2_X1 U7975 ( .A1(n10232), .A2(n10223), .ZN(n9812) );
  NAND2_X1 U7976 ( .A1(n6247), .A2(n4941), .ZN(P1_U3521) );
  INV_X1 U7977 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6248) );
  INV_X1 U7978 ( .A(n9771), .ZN(n9743) );
  NAND2_X1 U7979 ( .A1(n6250), .A2(n4940), .ZN(P1_U3553) );
  NAND2_X1 U7980 ( .A1(n6252), .A2(n6251), .ZN(n6254) );
  INV_X1 U7981 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9097) );
  OR2_X1 U7982 ( .A1(n8363), .A2(n9097), .ZN(n8566) );
  NAND2_X1 U7983 ( .A1(n7918), .A2(n8569), .ZN(n8360) );
  NAND2_X1 U7984 ( .A1(n7919), .A2(n10293), .ZN(n6276) );
  INV_X1 U7985 ( .A(n6256), .ZN(n6257) );
  NAND2_X1 U7986 ( .A1(n6257), .A2(n4950), .ZN(n6270) );
  INV_X1 U7987 ( .A(n8576), .ZN(n8587) );
  OAI211_X1 U7988 ( .C1(n8587), .C2(n8582), .A(n6271), .B(n10257), .ZN(n6258)
         );
  INV_X1 U7989 ( .A(n6258), .ZN(n6269) );
  NAND3_X1 U7990 ( .A1(n8576), .A2(n8766), .A3(n10257), .ZN(n6267) );
  INV_X1 U7991 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8952) );
  NAND2_X1 U7992 ( .A1(n4311), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6261) );
  NAND2_X1 U7993 ( .A1(n6259), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6260) );
  OAI211_X1 U7994 ( .C1(n8952), .C2(n6262), .A(n6261), .B(n6260), .ZN(n6263)
         );
  INV_X1 U7995 ( .A(n6263), .ZN(n6264) );
  NAND2_X1 U7996 ( .A1(n8373), .A2(n6264), .ZN(n8619) );
  AND2_X1 U7997 ( .A1(n5762), .A2(P2_B_REG_SCAN_IN), .ZN(n6265) );
  NOR2_X1 U7998 ( .A1(n8910), .A2(n6265), .ZN(n8757) );
  AOI22_X1 U7999 ( .A1(n10262), .A2(n8766), .B1(n8619), .B2(n8757), .ZN(n6266)
         );
  OAI21_X1 U8000 ( .B1(n6271), .B2(n6267), .A(n6266), .ZN(n6268) );
  INV_X1 U8001 ( .A(n6270), .ZN(n6273) );
  INV_X1 U8002 ( .A(n6271), .ZN(n6272) );
  NAND2_X1 U8003 ( .A1(n6276), .A2(n7914), .ZN(n6290) );
  NAND2_X1 U8004 ( .A1(n6290), .A2(n10308), .ZN(n6281) );
  INV_X1 U8005 ( .A(n7918), .ZN(n6277) );
  NAND2_X1 U8006 ( .A1(n7918), .A2(n6278), .ZN(n6280) );
  NAND2_X1 U8007 ( .A1(n10310), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U8008 ( .A1(n6281), .A2(n4932), .ZN(P2_U3456) );
  NAND2_X1 U8009 ( .A1(n6305), .A2(n6514), .ZN(n6284) );
  OR2_X1 U8010 ( .A1(n6282), .A2(n8613), .ZN(n6283) );
  NAND2_X1 U8011 ( .A1(n6284), .A2(n6304), .ZN(n6289) );
  NAND2_X1 U8012 ( .A1(n6518), .A2(n8591), .ZN(n6618) );
  INV_X1 U8013 ( .A(n6304), .ZN(n6287) );
  NAND2_X1 U8014 ( .A1(n6287), .A2(n6656), .ZN(n6288) );
  AND3_X2 U8015 ( .A1(n6289), .A2(n6303), .A3(n6288), .ZN(n10323) );
  NAND2_X1 U8016 ( .A1(n6290), .A2(n10323), .ZN(n6295) );
  INV_X1 U8017 ( .A(n8994), .ZN(n6292) );
  NAND2_X1 U8018 ( .A1(n10320), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6291) );
  INV_X1 U8019 ( .A(n6293), .ZN(n6294) );
  NAND2_X1 U8020 ( .A1(n6295), .A2(n6294), .ZN(P2_U3488) );
  NAND2_X1 U8021 ( .A1(n6296), .A2(n10232), .ZN(n6301) );
  INV_X1 U8022 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6297) );
  OR2_X1 U8023 ( .A1(n10232), .A2(n6297), .ZN(n6298) );
  INV_X1 U8024 ( .A(n6299), .ZN(n6300) );
  NAND2_X1 U8025 ( .A1(n6301), .A2(n6300), .ZN(P1_U3519) );
  NAND2_X1 U8026 ( .A1(n6304), .A2(n6656), .ZN(n6302) );
  OAI211_X1 U8027 ( .C1(n6304), .C2(n6514), .A(n6303), .B(n6302), .ZN(n6309)
         );
  INV_X1 U8028 ( .A(n6305), .ZN(n6306) );
  NAND2_X2 U8029 ( .A1(n6309), .A2(n10253), .ZN(n10269) );
  OR2_X1 U8030 ( .A1(n6307), .A2(n8445), .ZN(n7353) );
  NAND2_X1 U8031 ( .A1(n10265), .A2(n7353), .ZN(n6308) );
  INV_X2 U8032 ( .A(n10253), .ZN(n8942) );
  AOI22_X1 U8033 ( .A1(n8232), .A2(n8942), .B1(n10272), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n6311) );
  OR2_X1 U8034 ( .A1(n6309), .A2(n10251), .ZN(n8880) );
  NAND2_X1 U8035 ( .A1(n8576), .A2(n8929), .ZN(n6310) );
  OAI211_X1 U8036 ( .C1(n6508), .C2(n8932), .A(n6311), .B(n6310), .ZN(n6312)
         );
  INV_X1 U8037 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9760) );
  XNOR2_X1 U8038 ( .A(n10057), .B(n9760), .ZN(n10064) );
  OR2_X1 U8039 ( .A1(n6351), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6325) );
  INV_X1 U8040 ( .A(n6351), .ZN(n10046) );
  XNOR2_X1 U8041 ( .A(n10046), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n10044) );
  INV_X1 U8042 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10235) );
  INV_X1 U8043 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10233) );
  MUX2_X1 U8044 ( .A(n10233), .B(P1_REG1_REG_1__SCAN_IN), .S(n6680), .Z(n9405)
         );
  AND2_X1 U8045 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9404) );
  NAND2_X1 U8046 ( .A1(n9405), .A2(n9404), .ZN(n9403) );
  NAND2_X1 U8047 ( .A1(n9409), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6316) );
  NAND2_X1 U8048 ( .A1(n9403), .A2(n6316), .ZN(n6938) );
  NAND2_X1 U8049 ( .A1(n6939), .A2(n6938), .ZN(n6937) );
  NAND2_X1 U8050 ( .A1(n6940), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6317) );
  NAND2_X1 U8051 ( .A1(n6937), .A2(n6317), .ZN(n9422) );
  XNOR2_X1 U8052 ( .A(n9414), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9423) );
  NAND2_X1 U8053 ( .A1(n9422), .A2(n9423), .ZN(n9421) );
  INV_X1 U8054 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6318) );
  OR2_X1 U8055 ( .A1(n9414), .A2(n6318), .ZN(n6319) );
  NAND2_X1 U8056 ( .A1(n9421), .A2(n6319), .ZN(n9433) );
  INV_X1 U8057 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6320) );
  XNOR2_X1 U8058 ( .A(n6338), .B(n6320), .ZN(n9434) );
  INV_X1 U8059 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6321) );
  MUX2_X1 U8060 ( .A(n6321), .B(P1_REG1_REG_5__SCAN_IN), .S(n9448), .Z(n9443)
         );
  XNOR2_X1 U8061 ( .A(n9462), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n9456) );
  INV_X1 U8062 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6322) );
  MUX2_X1 U8063 ( .A(n6322), .B(P1_REG1_REG_7__SCAN_IN), .S(n9476), .Z(n9470)
         );
  NOR2_X1 U8064 ( .A1(n9471), .A2(n9470), .ZN(n9469) );
  XNOR2_X1 U8065 ( .A(n9490), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n9484) );
  INV_X1 U8066 ( .A(n6343), .ZN(n7012) );
  XNOR2_X1 U8067 ( .A(n7012), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n7010) );
  OAI21_X1 U8068 ( .B1(n6343), .B2(P1_REG1_REG_9__SCAN_IN), .A(n7008), .ZN(
        n7192) );
  XNOR2_X1 U8069 ( .A(n7196), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n7193) );
  NOR2_X1 U8070 ( .A1(n7192), .A2(n7193), .ZN(n7191) );
  XNOR2_X1 U8071 ( .A(n7311), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n7307) );
  NOR2_X1 U8072 ( .A1(n7308), .A2(n7307), .ZN(n7306) );
  INV_X1 U8073 ( .A(n6346), .ZN(n7411) );
  XNOR2_X1 U8074 ( .A(n7411), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n7409) );
  XNOR2_X1 U8075 ( .A(n7615), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n7612) );
  XNOR2_X1 U8076 ( .A(n10026), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n10022) );
  NOR2_X1 U8077 ( .A1(n6323), .A2(n4450), .ZN(n6324) );
  INV_X1 U8078 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10032) );
  NAND2_X1 U8079 ( .A1(n10044), .A2(n10045), .ZN(n10043) );
  NAND2_X1 U8080 ( .A1(n10082), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6326) );
  OAI21_X1 U8081 ( .B1(n10082), .B2(P1_REG1_REG_18__SCAN_IN), .A(n6326), .ZN(
        n10077) );
  NAND2_X1 U8082 ( .A1(n10080), .A2(n6326), .ZN(n6327) );
  XNOR2_X1 U8083 ( .A(n6327), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n6360) );
  OR2_X1 U8084 ( .A1(n6328), .A2(P1_U3086), .ZN(n8162) );
  NAND2_X1 U8085 ( .A1(n8158), .A2(n8162), .ZN(n6355) );
  INV_X1 U8086 ( .A(n6328), .ZN(n6329) );
  OR2_X1 U8087 ( .A1(n6870), .A2(n6329), .ZN(n6330) );
  AND2_X1 U8088 ( .A1(n6330), .A2(n5014), .ZN(n6354) );
  NAND2_X1 U8089 ( .A1(n6355), .A2(n6354), .ZN(n10016) );
  OR2_X1 U8090 ( .A1(n8189), .A2(n10002), .ZN(n6331) );
  OR2_X1 U8091 ( .A1(n10016), .A2(n6331), .ZN(n10047) );
  INV_X1 U8092 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9874) );
  MUX2_X1 U8093 ( .A(P1_REG2_REG_18__SCAN_IN), .B(n9874), .S(n10082), .Z(
        n10076) );
  NOR2_X1 U8094 ( .A1(n10057), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6332) );
  AOI21_X1 U8095 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n10057), .A(n6332), .ZN(
        n10060) );
  INV_X1 U8096 ( .A(n7311), .ZN(n6700) );
  INV_X1 U8097 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7462) );
  INV_X1 U8098 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6345) );
  INV_X1 U8099 ( .A(n7196), .ZN(n6684) );
  INV_X1 U8100 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6344) );
  INV_X1 U8101 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6342) );
  INV_X1 U8102 ( .A(n9490), .ZN(n6677) );
  INV_X1 U8103 ( .A(n9476), .ZN(n6669) );
  INV_X1 U8104 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6341) );
  INV_X1 U8105 ( .A(n9462), .ZN(n6675) );
  INV_X1 U8106 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6340) );
  INV_X1 U8107 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7073) );
  INV_X1 U8108 ( .A(n9448), .ZN(n6644) );
  INV_X1 U8109 ( .A(n6338), .ZN(n9429) );
  INV_X1 U8110 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6339) );
  INV_X1 U8111 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6333) );
  MUX2_X1 U8112 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6333), .S(n6940), .Z(n6936)
         );
  INV_X1 U8113 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7150) );
  MUX2_X1 U8114 ( .A(n7150), .B(P1_REG2_REG_1__SCAN_IN), .S(n6680), .Z(n9408)
         );
  AND2_X1 U8115 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9407) );
  NAND2_X1 U8116 ( .A1(n9408), .A2(n9407), .ZN(n9406) );
  NAND2_X1 U8117 ( .A1(n9409), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6334) );
  NAND2_X1 U8118 ( .A1(n9406), .A2(n6334), .ZN(n6935) );
  NAND2_X1 U8119 ( .A1(n6936), .A2(n6935), .ZN(n6934) );
  NAND2_X1 U8120 ( .A1(n6940), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U8121 ( .A1(n6934), .A2(n6335), .ZN(n9419) );
  NAND2_X1 U8122 ( .A1(n9419), .A2(n9420), .ZN(n9418) );
  INV_X1 U8123 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6336) );
  OR2_X1 U8124 ( .A1(n9414), .A2(n6336), .ZN(n6337) );
  NAND2_X1 U8125 ( .A1(n9418), .A2(n6337), .ZN(n9436) );
  XNOR2_X1 U8126 ( .A(n6338), .B(n6339), .ZN(n9437) );
  NAND2_X1 U8127 ( .A1(n9436), .A2(n9437), .ZN(n9435) );
  MUX2_X1 U8128 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7073), .S(n9448), .Z(n9451)
         );
  XOR2_X1 U8129 ( .A(n9462), .B(P1_REG2_REG_6__SCAN_IN), .Z(n9465) );
  OAI21_X1 U8130 ( .B1(n6675), .B2(n6340), .A(n9463), .ZN(n9479) );
  MUX2_X1 U8131 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n6341), .S(n9476), .Z(n9478)
         );
  NAND2_X1 U8132 ( .A1(n9479), .A2(n9478), .ZN(n9477) );
  OAI21_X1 U8133 ( .B1(n6669), .B2(n6341), .A(n9477), .ZN(n9493) );
  XOR2_X1 U8134 ( .A(n9490), .B(P1_REG2_REG_8__SCAN_IN), .Z(n9492) );
  NAND2_X1 U8135 ( .A1(n9493), .A2(n9492), .ZN(n9491) );
  OAI21_X1 U8136 ( .B1(n6342), .B2(n6677), .A(n9491), .ZN(n7006) );
  XNOR2_X1 U8137 ( .A(n6343), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n7007) );
  NOR2_X1 U8138 ( .A1(n7006), .A2(n7007), .ZN(n7005) );
  AOI21_X1 U8139 ( .B1(n7012), .B2(n6344), .A(n7005), .ZN(n7199) );
  XOR2_X1 U8140 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n7196), .Z(n7198) );
  NAND2_X1 U8141 ( .A1(n7199), .A2(n7198), .ZN(n7197) );
  OAI21_X1 U8142 ( .B1(n6345), .B2(n6684), .A(n7197), .ZN(n7314) );
  MUX2_X1 U8143 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n7462), .S(n7311), .Z(n7313)
         );
  NAND2_X1 U8144 ( .A1(n7314), .A2(n7313), .ZN(n7312) );
  XNOR2_X1 U8145 ( .A(n6346), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n7406) );
  XOR2_X1 U8146 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n7615), .Z(n7617) );
  NAND2_X1 U8147 ( .A1(n7615), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6347) );
  NAND2_X1 U8148 ( .A1(n10026), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6348) );
  OAI21_X1 U8149 ( .B1(n10026), .B2(P1_REG2_REG_14__SCAN_IN), .A(n6348), .ZN(
        n10019) );
  NOR2_X1 U8150 ( .A1(n6349), .A2(n4450), .ZN(n6350) );
  INV_X1 U8151 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10035) );
  NOR2_X1 U8152 ( .A1(n6350), .A2(n10034), .ZN(n10050) );
  INV_X1 U8153 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9859) );
  AOI22_X1 U8154 ( .A1(n6351), .A2(n9859), .B1(P1_REG2_REG_16__SCAN_IN), .B2(
        n10046), .ZN(n10049) );
  NAND2_X1 U8155 ( .A1(n10082), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6352) );
  OAI22_X1 U8156 ( .A1(n6360), .A2(n10030), .B1(n10047), .B2(n6353), .ZN(n6359) );
  INV_X1 U8157 ( .A(n6354), .ZN(n6356) );
  NAND2_X1 U8158 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n6357) );
  OAI21_X1 U8159 ( .B1(n10089), .B2(n4489), .A(n6357), .ZN(n6358) );
  NAND2_X1 U8160 ( .A1(n10081), .A2(n6360), .ZN(n6361) );
  OR2_X1 U8161 ( .A1(n10016), .A2(n6931), .ZN(n10069) );
  OAI211_X1 U8162 ( .C1(n10047), .C2(n6362), .A(n6361), .B(n10069), .ZN(n6363)
         );
  INV_X1 U8163 ( .A(n7577), .ZN(n6366) );
  OR2_X1 U8164 ( .A1(n8584), .A2(n6366), .ZN(n6367) );
  NAND2_X1 U8165 ( .A1(n6420), .A2(n6367), .ZN(n6390) );
  OR2_X1 U8166 ( .A1(n6390), .A2(n6368), .ZN(n6369) );
  NAND2_X1 U8167 ( .A1(n6369), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  OR2_X2 U8168 ( .A1(n6420), .A2(P2_U3151), .ZN(n8628) );
  INV_X1 U8169 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n6384) );
  INV_X1 U8170 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8993) );
  INV_X1 U8171 ( .A(n6920), .ZN(n6665) );
  AND2_X1 U8172 ( .A1(n6754), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6370) );
  NAND2_X1 U8173 ( .A1(n6393), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6371) );
  OAI21_X1 U8174 ( .B1(n6717), .B2(n6370), .A(n6371), .ZN(n6707) );
  INV_X1 U8175 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10311) );
  NAND2_X1 U8176 ( .A1(n6708), .A2(n6371), .ZN(n6766) );
  INV_X1 U8177 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10313) );
  XNOR2_X1 U8178 ( .A(n4448), .B(n10313), .ZN(n6767) );
  NAND2_X1 U8179 ( .A1(n6766), .A2(n6767), .ZN(n6765) );
  NAND2_X1 U8180 ( .A1(n4448), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U8181 ( .A1(n6796), .A2(n6724), .ZN(n6374) );
  XNOR2_X1 U8182 ( .A(n6434), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n6723) );
  INV_X1 U8183 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10316) );
  XNOR2_X1 U8184 ( .A(n6660), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n8638) );
  XNOR2_X1 U8185 ( .A(n6920), .B(n7335), .ZN(n6914) );
  INV_X1 U8186 ( .A(n6377), .ZN(n7164) );
  INV_X1 U8187 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7476) );
  XNOR2_X1 U8188 ( .A(n6459), .B(n7476), .ZN(n7165) );
  XNOR2_X1 U8189 ( .A(n7505), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n7496) );
  INV_X1 U8190 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9908) );
  INV_X1 U8191 ( .A(n8662), .ZN(n6904) );
  INV_X1 U8192 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8652) );
  INV_X1 U8193 ( .A(n6381), .ZN(n8675) );
  XNOR2_X1 U8194 ( .A(n6821), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n8674) );
  INV_X1 U8195 ( .A(n6478), .ZN(n8693) );
  INV_X1 U8196 ( .A(n6383), .ZN(n8702) );
  XNOR2_X1 U8197 ( .A(n6994), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8701) );
  INV_X1 U8198 ( .A(n6487), .ZN(n8727) );
  OAI21_X1 U8199 ( .B1(n6385), .B2(n8727), .A(n6389), .ZN(n8722) );
  INV_X1 U8200 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8983) );
  NAND2_X1 U8201 ( .A1(n8720), .A2(n6389), .ZN(n6387) );
  NAND2_X1 U8202 ( .A1(n8742), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8735) );
  OAI21_X1 U8203 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n8742), .A(n8735), .ZN(
        n6388) );
  INV_X1 U8204 ( .A(n6388), .ZN(n6386) );
  NAND3_X1 U8205 ( .A1(n8720), .A2(n6389), .A3(n6388), .ZN(n6391) );
  OR2_X1 U8206 ( .A1(n6390), .A2(P2_U3151), .ZN(n6496) );
  NOR2_X1 U8207 ( .A1(n6496), .A2(n6498), .ZN(n6417) );
  INV_X1 U8208 ( .A(n6417), .ZN(n6758) );
  AOI21_X1 U8209 ( .B1(n8736), .B2(n6391), .A(n8756), .ZN(n6392) );
  INV_X1 U8210 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n6411) );
  INV_X1 U8211 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6408) );
  AND2_X1 U8212 ( .A1(n6754), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6394) );
  NAND2_X1 U8213 ( .A1(n6393), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6395) );
  OAI21_X1 U8214 ( .B1(n6717), .B2(n6394), .A(n6395), .ZN(n6710) );
  INV_X1 U8215 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7043) );
  OR2_X1 U8216 ( .A1(n6710), .A2(n7043), .ZN(n6711) );
  NAND2_X1 U8217 ( .A1(n6711), .A2(n6395), .ZN(n6769) );
  INV_X1 U8218 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10271) );
  NAND2_X1 U8219 ( .A1(n6769), .A2(n6770), .ZN(n6768) );
  NAND2_X1 U8220 ( .A1(n4448), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6396) );
  NAND2_X1 U8221 ( .A1(n6797), .A2(n6719), .ZN(n6398) );
  XNOR2_X1 U8222 ( .A(n6434), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n6718) );
  INV_X1 U8223 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7064) );
  OR2_X1 U8224 ( .A1(n6434), .A2(n7064), .ZN(n6399) );
  NAND2_X1 U8225 ( .A1(n6722), .A2(n6399), .ZN(n6400) );
  NAND2_X1 U8226 ( .A1(n6400), .A2(n4756), .ZN(n8642) );
  INV_X1 U8227 ( .A(n6400), .ZN(n6401) );
  NAND2_X1 U8228 ( .A1(n6401), .A2(n6750), .ZN(n6402) );
  AND2_X2 U8229 ( .A1(n8642), .A2(n6402), .ZN(n6744) );
  NAND2_X2 U8230 ( .A1(n6744), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8644) );
  XNOR2_X1 U8231 ( .A(n6660), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n8643) );
  AOI21_X1 U8232 ( .B1(n8644), .B2(n8642), .A(n8643), .ZN(n8646) );
  INV_X1 U8233 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7289) );
  XNOR2_X1 U8234 ( .A(n6920), .B(n7289), .ZN(n6921) );
  INV_X1 U8235 ( .A(n6403), .ZN(n7180) );
  INV_X1 U8236 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7472) );
  XNOR2_X1 U8237 ( .A(n6459), .B(n7472), .ZN(n7181) );
  AOI21_X2 U8238 ( .B1(n7182), .B2(n7180), .A(n7181), .ZN(n7179) );
  XNOR2_X1 U8239 ( .A(n7505), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n7491) );
  INV_X1 U8240 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7585) );
  NAND2_X1 U8241 ( .A1(n6378), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6405) );
  INV_X1 U8242 ( .A(n6407), .ZN(n8683) );
  XNOR2_X1 U8243 ( .A(n6821), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n8682) );
  NAND2_X1 U8244 ( .A1(n6409), .A2(n8693), .ZN(n6410) );
  OAI21_X1 U8245 ( .B1(n6409), .B2(n8693), .A(n6410), .ZN(n8694) );
  INV_X1 U8246 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8927) );
  NOR2_X2 U8247 ( .A1(n8694), .A2(n8927), .ZN(n8711) );
  INV_X1 U8248 ( .A(n6410), .ZN(n8710) );
  XNOR2_X1 U8249 ( .A(n6994), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n8709) );
  OAI21_X2 U8250 ( .B1(n8711), .B2(n8710), .A(n8709), .ZN(n8714) );
  INV_X1 U8251 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8897) );
  NAND2_X1 U8252 ( .A1(n8742), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8737) );
  OAI21_X1 U8253 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8742), .A(n8737), .ZN(
        n6415) );
  INV_X1 U8254 ( .A(n6415), .ZN(n6413) );
  NAND2_X1 U8255 ( .A1(n6414), .A2(n6413), .ZN(n8738) );
  NAND3_X1 U8256 ( .A1(n8730), .A2(n6416), .A3(n6415), .ZN(n6418) );
  INV_X1 U8257 ( .A(n8740), .ZN(n8712) );
  AOI21_X1 U8258 ( .B1(n8738), .B2(n6418), .A(n8712), .ZN(n6419) );
  INV_X1 U8259 ( .A(n6419), .ZN(n6506) );
  INV_X1 U8260 ( .A(n6420), .ZN(n6421) );
  NOR2_X1 U8261 ( .A1(P2_U3150), .A2(n6421), .ZN(n8748) );
  INV_X1 U8262 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n6505) );
  MUX2_X1 U8263 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n9100), .Z(n6425) );
  INV_X1 U8264 ( .A(n4433), .ZN(n6422) );
  XNOR2_X1 U8265 ( .A(n6425), .B(n6422), .ZN(n6703) );
  INV_X1 U8266 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6424) );
  INV_X1 U8267 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6423) );
  MUX2_X1 U8268 ( .A(n6424), .B(n6423), .S(n9100), .Z(n6753) );
  NAND2_X1 U8269 ( .A1(n6753), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6757) );
  NAND2_X1 U8270 ( .A1(n6703), .A2(n6757), .ZN(n6427) );
  NAND2_X1 U8271 ( .A1(n6425), .A2(n4433), .ZN(n6426) );
  NAND2_X1 U8272 ( .A1(n6427), .A2(n6426), .ZN(n6764) );
  MUX2_X1 U8273 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n9100), .Z(n6428) );
  INV_X1 U8274 ( .A(n4448), .ZN(n6777) );
  XNOR2_X1 U8275 ( .A(n6428), .B(n6777), .ZN(n6763) );
  NAND2_X1 U8276 ( .A1(n6764), .A2(n6763), .ZN(n6430) );
  NAND2_X1 U8277 ( .A1(n6428), .A2(n4448), .ZN(n6429) );
  MUX2_X1 U8278 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n9100), .Z(n6431) );
  XNOR2_X1 U8279 ( .A(n6431), .B(n6647), .ZN(n6795) );
  MUX2_X1 U8280 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n6472), .Z(n6435) );
  XNOR2_X1 U8281 ( .A(n6435), .B(n6434), .ZN(n6734) );
  INV_X1 U8282 ( .A(n6431), .ZN(n6432) );
  NAND2_X1 U8283 ( .A1(n6432), .A2(n4764), .ZN(n6732) );
  AND2_X1 U8284 ( .A1(n6734), .A2(n6732), .ZN(n6433) );
  NAND2_X1 U8285 ( .A1(n6792), .A2(n6433), .ZN(n6733) );
  INV_X1 U8286 ( .A(n6434), .ZN(n6738) );
  NAND2_X1 U8287 ( .A1(n6435), .A2(n6738), .ZN(n6436) );
  NAND2_X1 U8288 ( .A1(n6733), .A2(n6436), .ZN(n6740) );
  MUX2_X1 U8289 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n6472), .Z(n6437) );
  XNOR2_X1 U8290 ( .A(n6437), .B(n6750), .ZN(n6739) );
  INV_X1 U8291 ( .A(n6437), .ZN(n6438) );
  NOR2_X1 U8292 ( .A1(n6438), .A2(n6750), .ZN(n6439) );
  INV_X1 U8293 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7215) );
  INV_X1 U8294 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6440) );
  MUX2_X1 U8295 ( .A(n7215), .B(n6440), .S(n6472), .Z(n6441) );
  NAND2_X1 U8296 ( .A1(n6441), .A2(n8636), .ZN(n6886) );
  INV_X1 U8297 ( .A(n6441), .ZN(n6442) );
  NAND2_X1 U8298 ( .A1(n6442), .A2(n6660), .ZN(n6443) );
  AND2_X1 U8299 ( .A1(n6886), .A2(n6443), .ZN(n8630) );
  NAND2_X1 U8300 ( .A1(n8631), .A2(n8630), .ZN(n8629) );
  NAND2_X1 U8301 ( .A1(n8629), .A2(n6886), .ZN(n6448) );
  INV_X1 U8302 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7362) );
  INV_X1 U8303 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10321) );
  MUX2_X1 U8304 ( .A(n7362), .B(n10321), .S(n6472), .Z(n6444) );
  NAND2_X1 U8305 ( .A1(n6444), .A2(n6445), .ZN(n6906) );
  INV_X1 U8306 ( .A(n6444), .ZN(n6446) );
  NAND2_X1 U8307 ( .A1(n6446), .A2(n4750), .ZN(n6447) );
  AND2_X1 U8308 ( .A1(n6906), .A2(n6447), .ZN(n6884) );
  NAND2_X1 U8309 ( .A1(n6910), .A2(n6906), .ZN(n6452) );
  MUX2_X1 U8310 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n6472), .Z(n6449) );
  NAND2_X1 U8311 ( .A1(n6665), .A2(n6449), .ZN(n6451) );
  INV_X1 U8312 ( .A(n6449), .ZN(n6450) );
  NAND2_X1 U8313 ( .A1(n6450), .A2(n6920), .ZN(n7053) );
  AND2_X1 U8314 ( .A1(n6451), .A2(n7053), .ZN(n6908) );
  NAND2_X1 U8315 ( .A1(n6452), .A2(n6908), .ZN(n7054) );
  NAND2_X1 U8316 ( .A1(n7054), .A2(n7053), .ZN(n6457) );
  INV_X1 U8317 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7448) );
  INV_X1 U8318 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7469) );
  MUX2_X1 U8319 ( .A(n7448), .B(n7469), .S(n6472), .Z(n6453) );
  NAND2_X1 U8320 ( .A1(n7050), .A2(n6453), .ZN(n7175) );
  INV_X1 U8321 ( .A(n6453), .ZN(n6454) );
  NAND2_X1 U8322 ( .A1(n6683), .A2(n6454), .ZN(n6455) );
  NAND2_X1 U8323 ( .A1(n7175), .A2(n6455), .ZN(n7052) );
  INV_X1 U8324 ( .A(n7052), .ZN(n6456) );
  NAND2_X1 U8325 ( .A1(n7176), .A2(n7175), .ZN(n6461) );
  MUX2_X1 U8326 ( .A(n7472), .B(n7476), .S(n6472), .Z(n6458) );
  OR2_X1 U8327 ( .A1(n6459), .A2(n6458), .ZN(n6460) );
  NAND2_X1 U8328 ( .A1(n6459), .A2(n6458), .ZN(n6462) );
  AND2_X1 U8329 ( .A1(n6460), .A2(n6462), .ZN(n7173) );
  NAND2_X1 U8330 ( .A1(n6461), .A2(n7173), .ZN(n7178) );
  NAND2_X1 U8331 ( .A1(n7178), .A2(n6462), .ZN(n7366) );
  MUX2_X1 U8332 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n9100), .Z(n6463) );
  XNOR2_X1 U8333 ( .A(n6463), .B(n7367), .ZN(n7365) );
  NAND2_X1 U8334 ( .A1(n7366), .A2(n7365), .ZN(n7364) );
  INV_X1 U8335 ( .A(n6463), .ZN(n6464) );
  NAND2_X1 U8336 ( .A1(n6464), .A2(n7367), .ZN(n6465) );
  NAND2_X1 U8337 ( .A1(n7364), .A2(n6465), .ZN(n7490) );
  MUX2_X1 U8338 ( .A(n7585), .B(n9908), .S(n9100), .Z(n6466) );
  AND2_X1 U8339 ( .A1(n6466), .A2(n7505), .ZN(n7486) );
  OR2_X1 U8340 ( .A1(n7490), .A2(n7486), .ZN(n6468) );
  INV_X1 U8341 ( .A(n6466), .ZN(n6467) );
  NAND2_X1 U8342 ( .A1(n6467), .A2(n6378), .ZN(n7487) );
  NAND2_X1 U8343 ( .A1(n6468), .A2(n7487), .ZN(n8656) );
  MUX2_X1 U8344 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n6472), .Z(n6469) );
  XNOR2_X1 U8345 ( .A(n6469), .B(n6904), .ZN(n8655) );
  INV_X1 U8346 ( .A(n6469), .ZN(n6470) );
  NAND2_X1 U8347 ( .A1(n6470), .A2(n8662), .ZN(n6471) );
  NAND2_X1 U8348 ( .A1(n8659), .A2(n6471), .ZN(n8670) );
  MUX2_X1 U8349 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n6472), .Z(n6473) );
  XNOR2_X1 U8350 ( .A(n6473), .B(n6821), .ZN(n8669) );
  NAND2_X1 U8351 ( .A1(n8670), .A2(n8669), .ZN(n8668) );
  INV_X1 U8352 ( .A(n6473), .ZN(n6474) );
  NAND2_X1 U8353 ( .A1(n6474), .A2(n6821), .ZN(n6475) );
  NAND2_X1 U8354 ( .A1(n8668), .A2(n6475), .ZN(n8690) );
  MUX2_X1 U8355 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n9100), .Z(n6476) );
  XNOR2_X1 U8356 ( .A(n6478), .B(n6476), .ZN(n8689) );
  NAND2_X1 U8357 ( .A1(n8690), .A2(n8689), .ZN(n6480) );
  INV_X1 U8358 ( .A(n6476), .ZN(n6477) );
  NAND2_X1 U8359 ( .A1(n6478), .A2(n6477), .ZN(n6479) );
  NAND2_X1 U8360 ( .A1(n6480), .A2(n6479), .ZN(n8705) );
  MUX2_X1 U8361 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n9100), .Z(n6481) );
  XNOR2_X1 U8362 ( .A(n6994), .B(n6481), .ZN(n8704) );
  NAND2_X1 U8363 ( .A1(n8705), .A2(n8704), .ZN(n6484) );
  INV_X1 U8364 ( .A(n6481), .ZN(n6482) );
  NAND2_X1 U8365 ( .A1(n6994), .A2(n6482), .ZN(n6483) );
  NAND2_X1 U8366 ( .A1(n6484), .A2(n6483), .ZN(n8724) );
  MUX2_X1 U8367 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n9100), .Z(n6485) );
  XNOR2_X1 U8368 ( .A(n6487), .B(n6485), .ZN(n8723) );
  INV_X1 U8369 ( .A(n6485), .ZN(n6486) );
  AND2_X1 U8370 ( .A1(n6487), .A2(n6486), .ZN(n6488) );
  MUX2_X1 U8371 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n6472), .Z(n6490) );
  AND2_X1 U8372 ( .A1(n6489), .A2(n6490), .ZN(n8743) );
  INV_X1 U8373 ( .A(n6489), .ZN(n6492) );
  INV_X1 U8374 ( .A(n6490), .ZN(n6491) );
  NAND2_X1 U8375 ( .A1(n6492), .A2(n6491), .ZN(n8741) );
  INV_X1 U8376 ( .A(n8741), .ZN(n6493) );
  INV_X1 U8377 ( .A(n6500), .ZN(n6495) );
  NOR2_X1 U8378 ( .A1(n8628), .A2(n6494), .ZN(n8753) );
  NAND2_X1 U8379 ( .A1(n6495), .A2(n8753), .ZN(n6503) );
  INV_X1 U8380 ( .A(n6496), .ZN(n6497) );
  NAND2_X1 U8381 ( .A1(n6497), .A2(n8744), .ZN(n6499) );
  MUX2_X1 U8382 ( .A(n8628), .B(n6499), .S(n6498), .Z(n8751) );
  AOI21_X1 U8383 ( .B1(n6500), .B2(P2_U3893), .A(n8663), .ZN(n6502) );
  MUX2_X1 U8384 ( .A(n6503), .B(n6502), .S(n6501), .Z(n6504) );
  NAND2_X1 U8385 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8328) );
  OR2_X1 U8386 ( .A1(n6507), .A2(n10320), .ZN(n6513) );
  NAND2_X1 U8387 ( .A1(n10323), .A2(n10293), .ZN(n8992) );
  NAND2_X1 U8388 ( .A1(n6513), .A2(n6512), .ZN(P2_U3487) );
  AOI21_X1 U8389 ( .B1(n6514), .B2(n8445), .A(n8613), .ZN(n6515) );
  INV_X1 U8390 ( .A(n6515), .ZN(n6517) );
  NAND2_X1 U8391 ( .A1(n6517), .A2(n6516), .ZN(n6519) );
  NAND2_X2 U8392 ( .A1(n6519), .A2(n6518), .ZN(n6526) );
  NOR2_X1 U8393 ( .A1(n6526), .A2(n9004), .ZN(n6520) );
  XNOR2_X1 U8394 ( .A(n6523), .B(n10256), .ZN(n6784) );
  INV_X1 U8395 ( .A(n6523), .ZN(n6524) );
  NAND2_X1 U8396 ( .A1(n6524), .A2(n10256), .ZN(n6525) );
  INV_X1 U8397 ( .A(n8627), .ZN(n8210) );
  NAND2_X1 U8398 ( .A1(n6807), .A2(n6808), .ZN(n6530) );
  INV_X1 U8399 ( .A(n6527), .ZN(n6528) );
  NAND2_X1 U8400 ( .A1(n6528), .A2(n8210), .ZN(n6529) );
  NAND2_X1 U8401 ( .A1(n6530), .A2(n6529), .ZN(n8205) );
  INV_X1 U8402 ( .A(n8205), .ZN(n6532) );
  XNOR2_X1 U8403 ( .A(n6533), .B(n10260), .ZN(n8204) );
  INV_X1 U8404 ( .A(n8204), .ZN(n6531) );
  NAND2_X1 U8405 ( .A1(n6532), .A2(n6531), .ZN(n8206) );
  NAND2_X1 U8406 ( .A1(n6533), .A2(n10260), .ZN(n6534) );
  AND2_X1 U8407 ( .A1(n8206), .A2(n6534), .ZN(n8287) );
  INV_X4 U8408 ( .A(n6600), .ZN(n8229) );
  XNOR2_X1 U8409 ( .A(n8229), .B(n8289), .ZN(n6535) );
  XNOR2_X1 U8410 ( .A(n6535), .B(n8626), .ZN(n8286) );
  NAND2_X1 U8411 ( .A1(n8287), .A2(n8286), .ZN(n8285) );
  INV_X1 U8412 ( .A(n8626), .ZN(n7020) );
  NAND2_X1 U8413 ( .A1(n6535), .A2(n7020), .ZN(n6536) );
  XNOR2_X1 U8414 ( .A(n6537), .B(n8229), .ZN(n6538) );
  XNOR2_X1 U8415 ( .A(n6538), .B(n7139), .ZN(n7018) );
  NOR2_X1 U8416 ( .A1(n6538), .A2(n8625), .ZN(n6539) );
  XNOR2_X1 U8417 ( .A(n7217), .B(n8229), .ZN(n6540) );
  XNOR2_X1 U8418 ( .A(n6540), .B(n7354), .ZN(n7027) );
  INV_X1 U8419 ( .A(n6540), .ZN(n6541) );
  NAND2_X1 U8420 ( .A1(n6541), .A2(n7354), .ZN(n6542) );
  XNOR2_X1 U8421 ( .A(n7350), .B(n8229), .ZN(n6544) );
  XNOR2_X1 U8422 ( .A(n6544), .B(n7265), .ZN(n7205) );
  INV_X1 U8423 ( .A(n7205), .ZN(n6543) );
  NAND2_X1 U8424 ( .A1(n6544), .A2(n7265), .ZN(n6545) );
  NAND2_X1 U8425 ( .A1(n7202), .A2(n6545), .ZN(n7262) );
  XNOR2_X1 U8426 ( .A(n7339), .B(n8229), .ZN(n6546) );
  XNOR2_X1 U8427 ( .A(n6546), .B(n7355), .ZN(n7261) );
  NAND2_X1 U8428 ( .A1(n6546), .A2(n7297), .ZN(n6547) );
  XNOR2_X1 U8429 ( .A(n7451), .B(n8229), .ZN(n6549) );
  XNOR2_X1 U8430 ( .A(n6549), .B(n7263), .ZN(n7294) );
  INV_X1 U8431 ( .A(n7294), .ZN(n6548) );
  INV_X1 U8432 ( .A(n6549), .ZN(n6550) );
  NAND2_X1 U8433 ( .A1(n6550), .A2(n7539), .ZN(n6551) );
  XNOR2_X1 U8434 ( .A(n6559), .B(n6600), .ZN(n7593) );
  XNOR2_X1 U8435 ( .A(n8481), .B(n6600), .ZN(n7590) );
  OR2_X1 U8436 ( .A1(n7590), .A2(n8623), .ZN(n6552) );
  NAND2_X1 U8437 ( .A1(n8229), .A2(n8623), .ZN(n6554) );
  OAI22_X1 U8438 ( .A1(n8481), .A2(n6554), .B1(n8484), .B2(n8229), .ZN(n6558)
         );
  NOR2_X1 U8439 ( .A1(n8482), .A2(n8229), .ZN(n6555) );
  AOI22_X1 U8440 ( .A1(n8481), .A2(n6555), .B1(n8229), .B2(n8622), .ZN(n6556)
         );
  NAND2_X1 U8441 ( .A1(n6559), .A2(n6556), .ZN(n6557) );
  OAI21_X1 U8442 ( .B1(n6559), .B2(n6558), .A(n6557), .ZN(n6560) );
  XNOR2_X1 U8443 ( .A(n7840), .B(n8229), .ZN(n6561) );
  XNOR2_X1 U8444 ( .A(n6561), .B(n8621), .ZN(n7881) );
  NAND2_X1 U8445 ( .A1(n7882), .A2(n7881), .ZN(n7880) );
  INV_X1 U8446 ( .A(n6561), .ZN(n6562) );
  NAND2_X1 U8447 ( .A1(n6562), .A2(n8621), .ZN(n6563) );
  XNOR2_X1 U8448 ( .A(n8436), .B(n8229), .ZN(n6565) );
  XNOR2_X1 U8449 ( .A(n6565), .B(n8194), .ZN(n8308) );
  INV_X1 U8450 ( .A(n8308), .ZN(n6564) );
  NAND2_X1 U8451 ( .A1(n6565), .A2(n8194), .ZN(n6566) );
  XNOR2_X1 U8452 ( .A(n9092), .B(n8229), .ZN(n6568) );
  XNOR2_X1 U8453 ( .A(n6568), .B(n8925), .ZN(n8191) );
  NAND2_X1 U8454 ( .A1(n6568), .A2(n6567), .ZN(n6569) );
  XNOR2_X1 U8455 ( .A(n8986), .B(n6600), .ZN(n8254) );
  XNOR2_X1 U8456 ( .A(n9085), .B(n6600), .ZN(n8256) );
  AND2_X1 U8457 ( .A1(n8256), .A2(n8936), .ZN(n8257) );
  AOI21_X1 U8458 ( .B1(n8254), .B2(n8924), .A(n8257), .ZN(n6570) );
  INV_X1 U8459 ( .A(n8254), .ZN(n8267) );
  OAI21_X1 U8460 ( .B1(n8256), .B2(n8936), .A(n8924), .ZN(n6573) );
  AND2_X1 U8461 ( .A1(n8892), .A2(n8909), .ZN(n6572) );
  INV_X1 U8462 ( .A(n8256), .ZN(n6571) );
  AOI22_X1 U8463 ( .A1(n8267), .A2(n6573), .B1(n6572), .B2(n6571), .ZN(n6574)
         );
  NAND2_X1 U8464 ( .A1(n6575), .A2(n6574), .ZN(n6576) );
  XNOR2_X1 U8465 ( .A(n9073), .B(n8229), .ZN(n6577) );
  XNOR2_X1 U8466 ( .A(n6577), .B(n8327), .ZN(n8266) );
  NAND2_X1 U8467 ( .A1(n6577), .A2(n8911), .ZN(n6578) );
  XNOR2_X1 U8468 ( .A(n8881), .B(n8229), .ZN(n6579) );
  XNOR2_X1 U8469 ( .A(n6579), .B(n8893), .ZN(n8325) );
  INV_X1 U8470 ( .A(n6579), .ZN(n6580) );
  INV_X1 U8471 ( .A(n8217), .ZN(n6582) );
  XNOR2_X1 U8472 ( .A(n8976), .B(n8229), .ZN(n6583) );
  XNOR2_X1 U8473 ( .A(n6583), .B(n8873), .ZN(n8218) );
  INV_X1 U8474 ( .A(n8218), .ZN(n6581) );
  INV_X1 U8475 ( .A(n6583), .ZN(n6584) );
  NAND2_X1 U8476 ( .A1(n6584), .A2(n8847), .ZN(n6585) );
  XNOR2_X1 U8477 ( .A(n9060), .B(n8229), .ZN(n6587) );
  XNOR2_X1 U8478 ( .A(n6587), .B(n8858), .ZN(n8298) );
  INV_X1 U8479 ( .A(n8298), .ZN(n6586) );
  XNOR2_X1 U8480 ( .A(n9054), .B(n8229), .ZN(n6588) );
  XNOR2_X1 U8481 ( .A(n6588), .B(n8846), .ZN(n8240) );
  NAND2_X1 U8482 ( .A1(n6588), .A2(n8301), .ZN(n6589) );
  XNOR2_X1 U8483 ( .A(n9048), .B(n8229), .ZN(n6591) );
  XNOR2_X1 U8484 ( .A(n6591), .B(n8832), .ZN(n8318) );
  XNOR2_X1 U8485 ( .A(n9036), .B(n8229), .ZN(n8279) );
  XNOR2_X1 U8486 ( .A(n9042), .B(n6600), .ZN(n8276) );
  INV_X1 U8487 ( .A(n8276), .ZN(n6592) );
  OAI22_X1 U8488 ( .A1(n8279), .A2(n8783), .B1(n8321), .B2(n6592), .ZN(n6596)
         );
  OAI21_X1 U8489 ( .B1(n8276), .B2(n8819), .A(n8805), .ZN(n6594) );
  NOR2_X1 U8490 ( .A1(n8805), .A2(n8819), .ZN(n6593) );
  AOI22_X1 U8491 ( .A1(n6594), .A2(n8279), .B1(n6593), .B2(n6592), .ZN(n6595)
         );
  XNOR2_X1 U8492 ( .A(n9030), .B(n8229), .ZN(n6597) );
  XNOR2_X1 U8493 ( .A(n6597), .B(n4568), .ZN(n8248) );
  XNOR2_X1 U8494 ( .A(n9024), .B(n8229), .ZN(n6598) );
  XNOR2_X1 U8495 ( .A(n6598), .B(n8782), .ZN(n8335) );
  INV_X1 U8496 ( .A(n6598), .ZN(n6599) );
  XNOR2_X1 U8497 ( .A(n9018), .B(n6600), .ZN(n6601) );
  NAND2_X1 U8498 ( .A1(n6601), .A2(n8775), .ZN(n8226) );
  OAI21_X1 U8499 ( .B1(n6601), .B2(n8775), .A(n8226), .ZN(n6608) );
  NAND2_X1 U8500 ( .A1(n6609), .A2(n6608), .ZN(n6607) );
  INV_X1 U8501 ( .A(n6602), .ZN(n6603) );
  NAND2_X1 U8502 ( .A1(n6610), .A2(n6603), .ZN(n6605) );
  OR2_X1 U8503 ( .A1(n6612), .A2(n6619), .ZN(n6604) );
  NAND2_X1 U8504 ( .A1(n6607), .A2(n6606), .ZN(n6636) );
  NOR2_X1 U8505 ( .A1(n6609), .A2(n6608), .ZN(n8228) );
  NAND2_X1 U8506 ( .A1(n6610), .A2(n10300), .ZN(n6611) );
  NAND2_X1 U8507 ( .A1(n9018), .A2(n8341), .ZN(n6635) );
  NOR2_X1 U8508 ( .A1(n6612), .A2(n6625), .ZN(n6615) );
  NAND2_X1 U8509 ( .A1(n6615), .A2(n6613), .ZN(n8339) );
  NAND2_X1 U8510 ( .A1(n6615), .A2(n6614), .ZN(n8350) );
  NAND2_X1 U8511 ( .A1(n8766), .A2(n8336), .ZN(n6632) );
  INV_X1 U8512 ( .A(n6616), .ZN(n6623) );
  AND3_X1 U8513 ( .A1(n6618), .A2(n6617), .A3(n7577), .ZN(n6621) );
  OR2_X1 U8514 ( .A1(n6626), .A2(n6619), .ZN(n6620) );
  OAI211_X1 U8515 ( .C1(n6623), .C2(n6622), .A(n6621), .B(n6620), .ZN(n6624)
         );
  NAND2_X1 U8516 ( .A1(n6624), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6629) );
  NOR2_X1 U8517 ( .A1(n6657), .A2(n6625), .ZN(n8606) );
  INV_X1 U8518 ( .A(n6626), .ZN(n6627) );
  NAND2_X1 U8519 ( .A1(n8606), .A2(n6627), .ZN(n6628) );
  AOI22_X1 U8520 ( .A1(n8769), .A2(n8352), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n6631) );
  OAI211_X1 U8521 ( .C1(n8782), .C2(n8339), .A(n6632), .B(n6631), .ZN(n6633)
         );
  OAI21_X1 U8522 ( .B1(n6636), .B2(n8228), .A(n4947), .ZN(P2_U3154) );
  INV_X1 U8523 ( .A(n6637), .ZN(n6638) );
  OR2_X2 U8524 ( .A1(n6832), .A2(n6638), .ZN(n9400) );
  AND2_X1 U8525 ( .A1(n6641), .A2(P2_U3151), .ZN(n7575) );
  INV_X2 U8526 ( .A(n7575), .ZN(n9106) );
  INV_X1 U8527 ( .A(n6639), .ZN(n6642) );
  NAND2_X1 U8528 ( .A1(n5659), .A2(P2_U3151), .ZN(n9101) );
  INV_X1 U8529 ( .A(n9101), .ZN(n7902) );
  INV_X1 U8530 ( .A(n7902), .ZN(n8187) );
  OAI222_X1 U8531 ( .A1(n4448), .A2(P2_U3151), .B1(n9106), .B2(n6642), .C1(
        n8187), .C2(n5751), .ZN(P2_U3293) );
  NAND2_X1 U8532 ( .A1(n6641), .A2(P1_U3086), .ZN(n7913) );
  AND2_X1 U8533 ( .A1(n5659), .A2(P1_U3086), .ZN(n7572) );
  INV_X2 U8534 ( .A(n7572), .ZN(n10008) );
  OAI222_X1 U8535 ( .A1(n7913), .A2(n6643), .B1(n10008), .B2(n6642), .C1(
        P1_U3086), .C2(n4650), .ZN(P1_U3353) );
  INV_X1 U8536 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6645) );
  OAI222_X1 U8537 ( .A1(n7913), .A2(n6645), .B1(n10008), .B2(n6649), .C1(n6644), .C2(P1_U3086), .ZN(P1_U3350) );
  OAI222_X1 U8538 ( .A1(n9106), .A2(n6667), .B1(n6647), .B2(P2_U3151), .C1(
        n6646), .C2(n8187), .ZN(P2_U3292) );
  OAI222_X1 U8539 ( .A1(n9106), .A2(n6679), .B1(n4433), .B2(P2_U3151), .C1(
        n4983), .C2(n8187), .ZN(P2_U3294) );
  INV_X1 U8540 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6648) );
  OAI222_X1 U8541 ( .A1(n9106), .A2(n6649), .B1(n4756), .B2(P2_U3151), .C1(
        n6648), .C2(n8187), .ZN(P2_U3290) );
  INV_X1 U8542 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6650) );
  OAI222_X1 U8543 ( .A1(n9106), .A2(n6670), .B1(n4750), .B2(P2_U3151), .C1(
        n6650), .C2(n8187), .ZN(P2_U3288) );
  INV_X1 U8544 ( .A(n6651), .ZN(n6653) );
  INV_X1 U8545 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6652) );
  OAI222_X1 U8546 ( .A1(n9106), .A2(n6653), .B1(n6738), .B2(P2_U3151), .C1(
        n6652), .C2(n8187), .ZN(P2_U3291) );
  INV_X1 U8547 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6654) );
  OAI222_X1 U8548 ( .A1(n7913), .A2(n6654), .B1(n10008), .B2(n6653), .C1(n9429), .C2(P1_U3086), .ZN(P1_U3351) );
  NAND2_X1 U8549 ( .A1(n6657), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6655) );
  OAI21_X1 U8550 ( .B1(n6657), .B2(n6656), .A(n6655), .ZN(P2_U3377) );
  INV_X1 U8551 ( .A(n6658), .ZN(n6674) );
  INV_X1 U8552 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6659) );
  OAI222_X1 U8553 ( .A1(n9106), .A2(n6674), .B1(n6660), .B2(P2_U3151), .C1(
        n6659), .C2(n8187), .ZN(P2_U3289) );
  INV_X1 U8554 ( .A(n6135), .ZN(n6661) );
  AND4_X1 U8555 ( .A1(n6153), .A2(P2_STATE_REG_SCAN_IN), .A3(n9103), .A4(n7577), .ZN(n6663) );
  AOI21_X1 U8556 ( .B1(n6672), .B2(n6134), .A(n6663), .ZN(P2_U3376) );
  INV_X1 U8557 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6666) );
  INV_X1 U8558 ( .A(n6664), .ZN(n6676) );
  OAI222_X1 U8559 ( .A1(n8187), .A2(n6666), .B1(n9106), .B2(n6676), .C1(
        P2_U3151), .C2(n6665), .ZN(P2_U3287) );
  AND2_X1 U8560 ( .A1(n6672), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8561 ( .A1(n6672), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8562 ( .A1(n6672), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8563 ( .A1(n6672), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8564 ( .A1(n6672), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8565 ( .A1(n6672), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8566 ( .A1(n6672), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8567 ( .A1(n6672), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8568 ( .A1(n6672), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8569 ( .A1(n6672), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8570 ( .A1(n6672), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8571 ( .A1(n6672), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8572 ( .A1(n6672), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8573 ( .A1(n6672), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8574 ( .A1(n6672), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8575 ( .A1(n6672), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8576 ( .A1(n6672), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8577 ( .A1(n6672), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8578 ( .A1(n6672), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8579 ( .A1(n6672), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8580 ( .A1(n6672), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8581 ( .A1(n6672), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8582 ( .A1(n6672), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8583 ( .A1(n6672), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8584 ( .A1(n6672), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8585 ( .A1(n6672), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8586 ( .A1(n6672), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8587 ( .A1(n6672), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  INV_X1 U8588 ( .A(n7913), .ZN(n7894) );
  OAI222_X1 U8589 ( .A1(n10005), .A2(n6668), .B1(n10008), .B2(n6667), .C1(
        n9414), .C2(P1_U3086), .ZN(P1_U3352) );
  INV_X1 U8590 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6671) );
  OAI222_X1 U8591 ( .A1(n10005), .A2(n6671), .B1(n10008), .B2(n6670), .C1(
        n6669), .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U8592 ( .A(n6672), .ZN(n6673) );
  INV_X1 U8593 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n9882) );
  NOR2_X1 U8594 ( .A1(n6673), .A2(n9882), .ZN(P2_U3254) );
  INV_X1 U8595 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n9944) );
  NOR2_X1 U8596 ( .A1(n6673), .A2(n9944), .ZN(P2_U3251) );
  INV_X1 U8597 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9894) );
  OAI222_X1 U8598 ( .A1(P1_U3086), .A2(n6675), .B1(n10005), .B2(n9894), .C1(
        n6674), .C2(n10008), .ZN(P1_U3349) );
  INV_X1 U8599 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6694) );
  OAI222_X1 U8600 ( .A1(P1_U3086), .A2(n6677), .B1(n10008), .B2(n6676), .C1(
        n10005), .C2(n6694), .ZN(P1_U3347) );
  INV_X1 U8601 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6678) );
  OAI222_X1 U8602 ( .A1(P1_U3086), .A2(n6680), .B1(n10008), .B2(n6679), .C1(
        n6678), .C2(n10005), .ZN(P1_U3354) );
  NOR2_X1 U8603 ( .A1(n10014), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8604 ( .A(n6681), .ZN(n6686) );
  OAI222_X1 U8605 ( .A1(n9106), .A2(n6686), .B1(n6683), .B2(P2_U3151), .C1(
        n6682), .C2(n8187), .ZN(P2_U3286) );
  INV_X1 U8606 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6685) );
  OAI222_X1 U8607 ( .A1(n7913), .A2(n6685), .B1(n10008), .B2(n6687), .C1(n6684), .C2(P1_U3086), .ZN(P1_U3345) );
  OAI222_X1 U8608 ( .A1(P1_U3086), .A2(n7012), .B1(n7913), .B2(n5147), .C1(
        n6686), .C2(n10008), .ZN(P1_U3346) );
  INV_X1 U8609 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6688) );
  OAI222_X1 U8610 ( .A1(n8187), .A2(n6688), .B1(n7172), .B2(P2_U3151), .C1(
        n9106), .C2(n6687), .ZN(P2_U3285) );
  NAND2_X1 U8611 ( .A1(n8050), .A2(P1_U3973), .ZN(n6689) );
  OAI21_X1 U8612 ( .B1(P1_U3973), .B2(n5751), .A(n6689), .ZN(P1_U3556) );
  NAND2_X1 U8613 ( .A1(n7000), .A2(P1_U3973), .ZN(n6690) );
  OAI21_X1 U8614 ( .B1(P1_U3973), .B2(n4987), .A(n6690), .ZN(P1_U3554) );
  NAND2_X1 U8615 ( .A1(P2_U3893), .A2(n7539), .ZN(n6691) );
  OAI21_X1 U8616 ( .B1(P2_U3893), .B2(n5147), .A(n6691), .ZN(P2_U3500) );
  NAND2_X1 U8617 ( .A1(P2_U3893), .A2(n7354), .ZN(n6692) );
  OAI21_X1 U8618 ( .B1(P2_U3893), .B2(n9894), .A(n6692), .ZN(P2_U3497) );
  NAND2_X1 U8619 ( .A1(n7355), .A2(P2_U3893), .ZN(n6693) );
  OAI21_X1 U8620 ( .B1(P2_U3893), .B2(n6694), .A(n6693), .ZN(P2_U3499) );
  INV_X1 U8621 ( .A(n9003), .ZN(n8386) );
  NAND2_X1 U8622 ( .A1(n7019), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6811) );
  NAND2_X1 U8623 ( .A1(n6811), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6698) );
  AOI22_X1 U8624 ( .A1(n8336), .A2(n6168), .B1(n8341), .B2(n9004), .ZN(n6697)
         );
  OAI211_X1 U8625 ( .C1(n8345), .C2(n8386), .A(n6698), .B(n6697), .ZN(P2_U3172) );
  INV_X1 U8626 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9948) );
  INV_X1 U8627 ( .A(n6699), .ZN(n6701) );
  OAI222_X1 U8628 ( .A1(n8187), .A2(n9948), .B1(n9106), .B2(n6701), .C1(
        P2_U3151), .C2(n4769), .ZN(P2_U3284) );
  INV_X1 U8629 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6702) );
  OAI222_X1 U8630 ( .A1(n7913), .A2(n6702), .B1(n10008), .B2(n6701), .C1(
        P1_U3086), .C2(n6700), .ZN(P1_U3344) );
  XOR2_X1 U8631 ( .A(n6703), .B(n6757), .Z(n6706) );
  INV_X1 U8632 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6704) );
  OAI22_X1 U8633 ( .A1(n8654), .A2(n10328), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6704), .ZN(n6705) );
  AOI21_X1 U8634 ( .B1(n8753), .B2(n6706), .A(n6705), .ZN(n6716) );
  INV_X1 U8635 ( .A(n8756), .ZN(n8639) );
  INV_X1 U8636 ( .A(n6707), .ZN(n6709) );
  OAI21_X1 U8637 ( .B1(n6709), .B2(P2_REG1_REG_1__SCAN_IN), .A(n6708), .ZN(
        n6714) );
  INV_X1 U8638 ( .A(n6710), .ZN(n6712) );
  OAI21_X1 U8639 ( .B1(n6712), .B2(P2_REG2_REG_1__SCAN_IN), .A(n6711), .ZN(
        n6713) );
  AOI22_X1 U8640 ( .A1(n8639), .A2(n6714), .B1(n8740), .B2(n6713), .ZN(n6715)
         );
  OAI211_X1 U8641 ( .C1(n4433), .C2(n8751), .A(n6716), .B(n6715), .ZN(P2_U3183) );
  INV_X1 U8642 ( .A(n6718), .ZN(n6720) );
  NAND3_X1 U8643 ( .A1(n6797), .A2(n6720), .A3(n6719), .ZN(n6721) );
  AOI21_X1 U8644 ( .B1(n6722), .B2(n6721), .A(n8712), .ZN(n6731) );
  INV_X1 U8645 ( .A(n6723), .ZN(n6725) );
  NAND3_X1 U8646 ( .A1(n6796), .A2(n6725), .A3(n6724), .ZN(n6726) );
  AOI21_X1 U8647 ( .B1(n6727), .B2(n6726), .A(n8756), .ZN(n6730) );
  INV_X1 U8648 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6728) );
  NAND2_X1 U8649 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n8290) );
  OAI21_X1 U8650 ( .B1(n8654), .B2(n6728), .A(n8290), .ZN(n6729) );
  NOR3_X1 U8651 ( .A1(n6731), .A2(n6730), .A3(n6729), .ZN(n6737) );
  AND2_X1 U8652 ( .A1(n6792), .A2(n6732), .ZN(n6735) );
  OAI211_X1 U8653 ( .C1(n6735), .C2(n6734), .A(n8753), .B(n6733), .ZN(n6736)
         );
  OAI211_X1 U8654 ( .C1(n8751), .C2(n6738), .A(n6737), .B(n6736), .ZN(P2_U3186) );
  XNOR2_X1 U8655 ( .A(n6740), .B(n6739), .ZN(n6752) );
  OAI21_X1 U8656 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n6742), .A(n6741), .ZN(
        n6743) );
  INV_X1 U8657 ( .A(n6743), .ZN(n6748) );
  AND2_X1 U8658 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7022) );
  AOI21_X1 U8659 ( .B1(n8748), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n7022), .ZN(
        n6747) );
  OAI21_X1 U8660 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n6744), .A(n8644), .ZN(
        n6745) );
  NAND2_X1 U8661 ( .A1(n8740), .A2(n6745), .ZN(n6746) );
  OAI211_X1 U8662 ( .C1(n6748), .C2(n8756), .A(n6747), .B(n6746), .ZN(n6749)
         );
  AOI21_X1 U8663 ( .B1(n6750), .B2(n8663), .A(n6749), .ZN(n6751) );
  OAI21_X1 U8664 ( .B1(n8657), .B2(n6752), .A(n6751), .ZN(P2_U3187) );
  INV_X1 U8665 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6762) );
  INV_X1 U8666 ( .A(n6753), .ZN(n6755) );
  NAND2_X1 U8667 ( .A1(n6755), .A2(n6754), .ZN(n6756) );
  AOI22_X1 U8668 ( .A1(n6758), .A2(n8657), .B1(n6757), .B2(n6756), .ZN(n6759)
         );
  AOI21_X1 U8669 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n6759), .ZN(
        n6761) );
  NAND2_X1 U8670 ( .A1(n8663), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6760) );
  OAI211_X1 U8671 ( .C1(n8654), .C2(n6762), .A(n6761), .B(n6760), .ZN(P2_U3182) );
  XNOR2_X1 U8672 ( .A(n6764), .B(n6763), .ZN(n6775) );
  OAI21_X1 U8673 ( .B1(n6767), .B2(n6766), .A(n6765), .ZN(n6772) );
  OAI21_X1 U8674 ( .B1(n6770), .B2(n6769), .A(n6768), .ZN(n6771) );
  AOI22_X1 U8675 ( .A1(n8639), .A2(n6772), .B1(n8740), .B2(n6771), .ZN(n6774)
         );
  AOI22_X1 U8676 ( .A1(n8748), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3151), .ZN(n6773) );
  OAI211_X1 U8677 ( .C1(n8657), .C2(n6775), .A(n6774), .B(n6773), .ZN(n6776)
         );
  AOI21_X1 U8678 ( .B1(n6777), .B2(n8663), .A(n6776), .ZN(n6778) );
  INV_X1 U8679 ( .A(n6778), .ZN(P2_U3184) );
  INV_X1 U8680 ( .A(n10140), .ZN(n9642) );
  NAND2_X1 U8681 ( .A1(n7000), .A2(n6901), .ZN(n8051) );
  INV_X1 U8682 ( .A(n8051), .ZN(n6779) );
  NOR2_X1 U8683 ( .A1(n7157), .A2(n6779), .ZN(n8113) );
  AOI21_X1 U8684 ( .B1(n10195), .B2(n9642), .A(n8113), .ZN(n6782) );
  INV_X1 U8685 ( .A(n9402), .ZN(n6875) );
  NOR2_X1 U8686 ( .A1(n6875), .A2(n9353), .ZN(n7078) );
  INV_X1 U8687 ( .A(n6837), .ZN(n6780) );
  NAND2_X1 U8688 ( .A1(n7151), .A2(n6780), .ZN(n7086) );
  INV_X1 U8689 ( .A(n7086), .ZN(n6781) );
  NOR3_X1 U8690 ( .A1(n6782), .A2(n7078), .A3(n6781), .ZN(n10165) );
  NAND2_X1 U8691 ( .A1(n10245), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6783) );
  OAI21_X1 U8692 ( .B1(n10165), .B2(n10245), .A(n6783), .ZN(P1_U3522) );
  XOR2_X1 U8693 ( .A(n6784), .B(n6785), .Z(n6789) );
  AOI22_X1 U8694 ( .A1(n8336), .A2(n8627), .B1(n8348), .B2(n6695), .ZN(n6786)
         );
  OAI21_X1 U8695 ( .B1(n6522), .B2(n8355), .A(n6786), .ZN(n6787) );
  AOI21_X1 U8696 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n6811), .A(n6787), .ZN(
        n6788) );
  OAI21_X1 U8697 ( .B1(n8345), .B2(n6789), .A(n6788), .ZN(P2_U3162) );
  INV_X1 U8698 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6791) );
  INV_X1 U8699 ( .A(n6790), .ZN(n6814) );
  OAI222_X1 U8700 ( .A1(n7913), .A2(n6791), .B1(n10008), .B2(n6814), .C1(n7411), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8701 ( .A(n6792), .ZN(n6793) );
  AOI21_X1 U8702 ( .B1(n6795), .B2(n6794), .A(n6793), .ZN(n6805) );
  INV_X1 U8703 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6802) );
  OAI21_X1 U8704 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n4417), .A(n6796), .ZN(
        n6800) );
  OAI21_X1 U8705 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n6798), .A(n6797), .ZN(
        n6799) );
  AOI22_X1 U8706 ( .A1(n8639), .A2(n6800), .B1(n8740), .B2(n6799), .ZN(n6801)
         );
  NAND2_X1 U8707 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8209) );
  OAI211_X1 U8708 ( .C1(n8654), .C2(n6802), .A(n6801), .B(n8209), .ZN(n6803)
         );
  AOI21_X1 U8709 ( .B1(n4764), .B2(n8663), .A(n6803), .ZN(n6804) );
  OAI21_X1 U8710 ( .B1(n6805), .B2(n8657), .A(n6804), .ZN(P2_U3185) );
  NAND2_X1 U8711 ( .A1(n8327), .A2(P2_U3893), .ZN(n6806) );
  OAI21_X1 U8712 ( .B1(P2_U3893), .B2(n5332), .A(n6806), .ZN(P2_U3508) );
  XOR2_X1 U8713 ( .A(n6807), .B(n6808), .Z(n6813) );
  AOI22_X1 U8714 ( .A1(n8348), .A2(n6168), .B1(n8336), .B2(n10260), .ZN(n6809)
         );
  OAI21_X1 U8715 ( .B1(n10278), .B2(n8355), .A(n6809), .ZN(n6810) );
  AOI21_X1 U8716 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n6811), .A(n6810), .ZN(
        n6812) );
  OAI21_X1 U8717 ( .B1(n6813), .B2(n8345), .A(n6812), .ZN(P2_U3177) );
  INV_X1 U8718 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6815) );
  OAI222_X1 U8719 ( .A1(n8187), .A2(n6815), .B1(n6378), .B2(P2_U3151), .C1(
        n9106), .C2(n6814), .ZN(P2_U3283) );
  AOI22_X1 U8720 ( .A1(n10026), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n7894), .ZN(n6816) );
  OAI21_X1 U8721 ( .B1(n6822), .B2(n10008), .A(n6816), .ZN(P1_U3341) );
  INV_X1 U8722 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7132) );
  NAND2_X1 U8723 ( .A1(n6817), .A2(P2_U3893), .ZN(n6818) );
  OAI21_X1 U8724 ( .B1(P2_U3893), .B2(n7132), .A(n6818), .ZN(P2_U3509) );
  INV_X1 U8725 ( .A(n6819), .ZN(n6903) );
  AOI22_X1 U8726 ( .A1(n7615), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n7894), .ZN(n6820) );
  OAI21_X1 U8727 ( .B1(n6903), .B2(n10008), .A(n6820), .ZN(P1_U3342) );
  INV_X1 U8728 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6823) );
  INV_X1 U8729 ( .A(n6821), .ZN(n8673) );
  OAI222_X1 U8730 ( .A1(n9101), .A2(n6823), .B1(n8673), .B2(P2_U3151), .C1(
        n9106), .C2(n6822), .ZN(P2_U3281) );
  NAND2_X1 U8731 ( .A1(n6824), .A2(n9997), .ZN(n6825) );
  OAI21_X1 U8732 ( .B1(n6876), .B2(n10213), .A(n6869), .ZN(n6829) );
  INV_X1 U8733 ( .A(n6827), .ZN(n6828) );
  NAND2_X1 U8734 ( .A1(n6829), .A2(n6828), .ZN(n6830) );
  NOR2_X1 U8735 ( .A1(n9364), .A2(P1_U3086), .ZN(n6896) );
  INV_X1 U8736 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6882) );
  AND2_X1 U8737 ( .A1(n4312), .A2(n7334), .ZN(n6831) );
  AND2_X4 U8738 ( .A1(n6836), .A2(n6832), .ZN(n9189) );
  NAND2_X1 U8739 ( .A1(n9189), .A2(n7155), .ZN(n6835) );
  NAND2_X1 U8740 ( .A1(n6833), .A2(n7710), .ZN(n6834) );
  NAND2_X1 U8741 ( .A1(n6835), .A2(n6834), .ZN(n6839) );
  XNOR2_X1 U8742 ( .A(n6839), .B(n4310), .ZN(n6844) );
  NAND2_X1 U8743 ( .A1(n8106), .A2(n7481), .ZN(n6840) );
  AND2_X1 U8744 ( .A1(n7148), .A2(n6840), .ZN(n6841) );
  AND2_X2 U8745 ( .A1(n6841), .A2(n6832), .ZN(n9194) );
  AND2_X1 U8746 ( .A1(n7710), .A2(n7155), .ZN(n6842) );
  AOI21_X1 U8747 ( .B1(n9402), .B2(n9194), .A(n6842), .ZN(n6843) );
  NAND2_X1 U8748 ( .A1(n6844), .A2(n6843), .ZN(n6865) );
  NAND2_X1 U8749 ( .A1(n6865), .A2(n4933), .ZN(n6998) );
  INV_X1 U8750 ( .A(n6998), .ZN(n6857) );
  NAND2_X1 U8751 ( .A1(n7000), .A2(n7710), .ZN(n6846) );
  NAND2_X1 U8752 ( .A1(n9189), .A2(n7151), .ZN(n6845) );
  NAND2_X1 U8753 ( .A1(n6846), .A2(n6845), .ZN(n6852) );
  INV_X1 U8754 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6847) );
  NOR2_X1 U8755 ( .A1(n6832), .A2(n6847), .ZN(n6848) );
  OR2_X1 U8756 ( .A1(n6852), .A2(n6848), .ZN(n6897) );
  NAND2_X1 U8757 ( .A1(n7000), .A2(n9194), .ZN(n6851) );
  INV_X1 U8758 ( .A(n6832), .ZN(n6849) );
  AOI22_X1 U8759 ( .A1(n7710), .A2(n7151), .B1(n6849), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n6850) );
  NAND2_X1 U8760 ( .A1(n6851), .A2(n6850), .ZN(n6898) );
  NAND2_X1 U8761 ( .A1(n6897), .A2(n6898), .ZN(n6855) );
  INV_X1 U8762 ( .A(n6852), .ZN(n6853) );
  NAND2_X1 U8763 ( .A1(n6853), .A2(n4310), .ZN(n6854) );
  NAND2_X1 U8764 ( .A1(n6855), .A2(n6854), .ZN(n6999) );
  INV_X1 U8765 ( .A(n6866), .ZN(n6997) );
  INV_X1 U8766 ( .A(n6865), .ZN(n6864) );
  NAND2_X1 U8767 ( .A1(n8050), .A2(n7710), .ZN(n6859) );
  NAND2_X1 U8768 ( .A1(n10147), .A2(n9189), .ZN(n6858) );
  NAND2_X1 U8769 ( .A1(n6859), .A2(n6858), .ZN(n6860) );
  XNOR2_X1 U8770 ( .A(n6860), .B(n4310), .ZN(n6862) );
  AOI22_X1 U8771 ( .A1(n8050), .A2(n9194), .B1(n10147), .B2(n7710), .ZN(n6861)
         );
  OR2_X1 U8772 ( .A1(n6862), .A2(n6861), .ZN(n6863) );
  NAND2_X1 U8773 ( .A1(n6862), .A2(n6861), .ZN(n6954) );
  AND2_X1 U8774 ( .A1(n6863), .A2(n6954), .ZN(n6867) );
  NOR3_X1 U8775 ( .A1(n6997), .A2(n6864), .A3(n6867), .ZN(n6873) );
  NAND2_X1 U8776 ( .A1(n6866), .A2(n6865), .ZN(n6868) );
  INV_X1 U8777 ( .A(n6955), .ZN(n6872) );
  NOR2_X1 U8778 ( .A1(n6869), .A2(n8158), .ZN(n6874) );
  AND2_X1 U8779 ( .A1(n10213), .A2(n6870), .ZN(n6871) );
  OAI21_X1 U8780 ( .B1(n6873), .B2(n6872), .A(n9349), .ZN(n6881) );
  INV_X1 U8781 ( .A(n6874), .ZN(n6878) );
  INV_X1 U8782 ( .A(n9401), .ZN(n6971) );
  OAI22_X1 U8783 ( .A1(n6875), .A2(n9351), .B1(n6971), .B2(n9353), .ZN(n10139)
         );
  INV_X1 U8784 ( .A(n6876), .ZN(n6877) );
  OR2_X1 U8785 ( .A1(n6878), .A2(n6877), .ZN(n6879) );
  AOI22_X1 U8786 ( .A1(n9356), .A2(n10139), .B1(n9369), .B2(n10147), .ZN(n6880) );
  OAI211_X1 U8787 ( .C1(n6896), .C2(n6882), .A(n6881), .B(n6880), .ZN(P1_U3237) );
  OAI21_X1 U8788 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n6883), .A(n6922), .ZN(
        n6894) );
  INV_X1 U8789 ( .A(n6884), .ZN(n6885) );
  NAND3_X1 U8790 ( .A1(n8629), .A2(n6886), .A3(n6885), .ZN(n6887) );
  AOI21_X1 U8791 ( .B1(n6910), .B2(n6887), .A(n8657), .ZN(n6893) );
  OAI21_X1 U8792 ( .B1(P2_REG1_REG_7__SCAN_IN), .B2(n6888), .A(n6915), .ZN(
        n6889) );
  NAND2_X1 U8793 ( .A1(n6889), .A2(n8639), .ZN(n6891) );
  AND2_X1 U8794 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7208) );
  AOI21_X1 U8795 ( .B1(n8748), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7208), .ZN(
        n6890) );
  OAI211_X1 U8796 ( .C1(n8751), .C2(n4750), .A(n6891), .B(n6890), .ZN(n6892)
         );
  AOI211_X1 U8797 ( .C1(n8740), .C2(n6894), .A(n6893), .B(n6892), .ZN(n6895)
         );
  INV_X1 U8798 ( .A(n6895), .ZN(P2_U3189) );
  INV_X1 U8799 ( .A(n6896), .ZN(n7002) );
  NAND2_X1 U8800 ( .A1(n7002), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6900) );
  XOR2_X1 U8801 ( .A(n6898), .B(n6897), .Z(n6929) );
  AOI22_X1 U8802 ( .A1(n6929), .A2(n9349), .B1(n9356), .B2(n7078), .ZN(n6899)
         );
  OAI211_X1 U8803 ( .C1(n9332), .C2(n6901), .A(n6900), .B(n6899), .ZN(P1_U3232) );
  INV_X1 U8804 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7244) );
  NAND2_X1 U8805 ( .A1(n8847), .A2(P2_U3893), .ZN(n6902) );
  OAI21_X1 U8806 ( .B1(P2_U3893), .B2(n7244), .A(n6902), .ZN(P2_U3510) );
  INV_X1 U8807 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6905) );
  OAI222_X1 U8808 ( .A1(n9101), .A2(n6905), .B1(n6904), .B2(P2_U3151), .C1(
        n9106), .C2(n6903), .ZN(P2_U3282) );
  INV_X1 U8809 ( .A(n6906), .ZN(n6907) );
  NOR2_X1 U8810 ( .A1(n6908), .A2(n6907), .ZN(n6911) );
  INV_X1 U8811 ( .A(n7054), .ZN(n6909) );
  AOI21_X1 U8812 ( .B1(n6911), .B2(n6910), .A(n6909), .ZN(n6927) );
  INV_X1 U8813 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n6912) );
  NAND2_X1 U8814 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7264) );
  OAI21_X1 U8815 ( .B1(n8654), .B2(n6912), .A(n7264), .ZN(n6919) );
  INV_X1 U8816 ( .A(n6913), .ZN(n6917) );
  NAND3_X1 U8817 ( .A1(n6915), .A2(n6914), .A3(n4335), .ZN(n6916) );
  AOI21_X1 U8818 ( .B1(n6917), .B2(n6916), .A(n8756), .ZN(n6918) );
  AOI211_X1 U8819 ( .C1(n8663), .C2(n6920), .A(n6919), .B(n6918), .ZN(n6926)
         );
  AND3_X1 U8820 ( .A1(n6922), .A2(n6921), .A3(n4315), .ZN(n6923) );
  OAI21_X1 U8821 ( .B1(n6924), .B2(n6923), .A(n8740), .ZN(n6925) );
  OAI211_X1 U8822 ( .C1(n6927), .C2(n8657), .A(n6926), .B(n6925), .ZN(P2_U3190) );
  NOR2_X1 U8823 ( .A1(n10002), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6928) );
  NOR2_X1 U8824 ( .A1(n6928), .A2(n8189), .ZN(n10011) );
  INV_X1 U8825 ( .A(n6929), .ZN(n6930) );
  MUX2_X1 U8826 ( .A(n9407), .B(n6930), .S(n10002), .Z(n6932) );
  NAND2_X1 U8827 ( .A1(n6932), .A2(n6931), .ZN(n6933) );
  OAI211_X1 U8828 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n10011), .A(n6933), .B(
        P1_U3973), .ZN(n9441) );
  INV_X1 U8829 ( .A(n9441), .ZN(n6946) );
  OAI211_X1 U8830 ( .C1(n6936), .C2(n6935), .A(n10075), .B(n6934), .ZN(n6944)
         );
  OAI211_X1 U8831 ( .C1(n6939), .C2(n6938), .A(n10081), .B(n6937), .ZN(n6943)
         );
  AOI22_X1 U8832 ( .A1(n10014), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6942) );
  NAND2_X1 U8833 ( .A1(n10083), .A2(n6940), .ZN(n6941) );
  NAND4_X1 U8834 ( .A1(n6944), .A2(n6943), .A3(n6942), .A4(n6941), .ZN(n6945)
         );
  OR2_X1 U8835 ( .A1(n6946), .A2(n6945), .ZN(P1_U3245) );
  INV_X1 U8836 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6950) );
  INV_X1 U8837 ( .A(n6947), .ZN(n6948) );
  NAND2_X1 U8838 ( .A1(n9003), .A2(n6948), .ZN(n6949) );
  OR2_X1 U8839 ( .A1(n10256), .A2(n8910), .ZN(n9006) );
  OAI211_X1 U8840 ( .C1(n10253), .C2(n6950), .A(n6949), .B(n9006), .ZN(n6951)
         );
  MUX2_X1 U8841 ( .A(n6951), .B(P2_REG2_REG_0__SCAN_IN), .S(n10272), .Z(n6952)
         );
  AOI21_X1 U8842 ( .B1(n8929), .B2(n9004), .A(n6952), .ZN(n6953) );
  INV_X1 U8843 ( .A(n6953), .ZN(P2_U3233) );
  NAND2_X1 U8844 ( .A1(n6955), .A2(n6954), .ZN(n9172) );
  NAND2_X1 U8845 ( .A1(n9401), .A2(n7710), .ZN(n6957) );
  NAND2_X1 U8846 ( .A1(n9175), .A2(n9189), .ZN(n6956) );
  NAND2_X1 U8847 ( .A1(n6957), .A2(n6956), .ZN(n6958) );
  XNOR2_X1 U8848 ( .A(n6958), .B(n9192), .ZN(n6964) );
  AOI22_X1 U8849 ( .A1(n9401), .A2(n9194), .B1(n7710), .B2(n9175), .ZN(n6965)
         );
  XNOR2_X1 U8850 ( .A(n6964), .B(n6965), .ZN(n9173) );
  NAND2_X1 U8851 ( .A1(n9399), .A2(n7710), .ZN(n6960) );
  OR2_X1 U8852 ( .A1(n10185), .A2(n7801), .ZN(n6959) );
  NAND2_X1 U8853 ( .A1(n6960), .A2(n6959), .ZN(n6961) );
  XNOR2_X1 U8854 ( .A(n6961), .B(n4310), .ZN(n7114) );
  NAND2_X1 U8855 ( .A1(n9399), .A2(n9194), .ZN(n6963) );
  OR2_X1 U8856 ( .A1(n10185), .A2(n7791), .ZN(n6962) );
  NAND2_X1 U8857 ( .A1(n6963), .A2(n6962), .ZN(n7115) );
  XNOR2_X1 U8858 ( .A(n7114), .B(n7115), .ZN(n6969) );
  INV_X1 U8859 ( .A(n6964), .ZN(n6966) );
  NAND2_X1 U8860 ( .A1(n6966), .A2(n6965), .ZN(n6970) );
  NAND2_X1 U8861 ( .A1(n7122), .A2(n9349), .ZN(n6976) );
  AOI21_X1 U8862 ( .B1(n6968), .B2(n6970), .A(n6969), .ZN(n6975) );
  OAI22_X1 U8863 ( .A1(n6971), .A2(n9351), .B1(n9352), .B2(n9353), .ZN(n10127)
         );
  AND2_X1 U8864 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9427) );
  AOI21_X1 U8865 ( .B1(n9356), .B2(n10127), .A(n9427), .ZN(n6974) );
  INV_X1 U8866 ( .A(n6972), .ZN(n10129) );
  AOI22_X1 U8867 ( .A1(n9369), .A2(n10131), .B1(n9364), .B2(n10129), .ZN(n6973) );
  OAI211_X1 U8868 ( .C1(n6976), .C2(n6975), .A(n6974), .B(n6973), .ZN(P1_U3230) );
  INV_X1 U8869 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6978) );
  INV_X1 U8870 ( .A(n6977), .ZN(n6979) );
  OAI222_X1 U8871 ( .A1(n7913), .A2(n6978), .B1(n10008), .B2(n6979), .C1(
        P1_U3086), .C2(n4450), .ZN(P1_U3340) );
  INV_X1 U8872 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6980) );
  OAI222_X1 U8873 ( .A1(n8187), .A2(n6980), .B1(n9106), .B2(n6979), .C1(
        P2_U3151), .C2(n8693), .ZN(P2_U3280) );
  OAI21_X1 U8874 ( .B1(n6982), .B2(n8387), .A(n6981), .ZN(n10287) );
  INV_X1 U8875 ( .A(n10287), .ZN(n6991) );
  INV_X1 U8876 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6988) );
  NAND3_X1 U8877 ( .A1(n6983), .A2(n8387), .A3(n6984), .ZN(n6985) );
  NAND2_X1 U8878 ( .A1(n6986), .A2(n6985), .ZN(n6987) );
  AOI222_X1 U8879 ( .A1(n10257), .A2(n6987), .B1(n8626), .B2(n10261), .C1(
        n8627), .C2(n10262), .ZN(n10284) );
  MUX2_X1 U8880 ( .A(n6988), .B(n10284), .S(n10269), .Z(n6990) );
  AOI22_X1 U8881 ( .A1(n8929), .A2(n8208), .B1(n8942), .B2(n8213), .ZN(n6989)
         );
  OAI211_X1 U8882 ( .C1(n6991), .C2(n8932), .A(n6990), .B(n6989), .ZN(P2_U3230) );
  INV_X1 U8883 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6993) );
  INV_X1 U8884 ( .A(n6992), .ZN(n6995) );
  OAI222_X1 U8885 ( .A1(n10005), .A2(n6993), .B1(n10008), .B2(n6995), .C1(
        P1_U3086), .C2(n10046), .ZN(P1_U3339) );
  INV_X1 U8886 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6996) );
  INV_X1 U8887 ( .A(n6994), .ZN(n8708) );
  OAI222_X1 U8888 ( .A1(n9101), .A2(n6996), .B1(n9106), .B2(n6995), .C1(
        P2_U3151), .C2(n8708), .ZN(P2_U3279) );
  AOI21_X1 U8889 ( .B1(n6999), .B2(n6998), .A(n6997), .ZN(n7004) );
  AOI22_X1 U8890 ( .A1(n9314), .A2(n8050), .B1(n7000), .B2(n9313), .ZN(n7160)
         );
  OAI22_X1 U8891 ( .A1(n9332), .A2(n10168), .B1(n7160), .B2(n9366), .ZN(n7001)
         );
  AOI21_X1 U8892 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n7002), .A(n7001), .ZN(
        n7003) );
  OAI21_X1 U8893 ( .B1(n7004), .B2(n9371), .A(n7003), .ZN(P1_U3222) );
  AOI21_X1 U8894 ( .B1(n7007), .B2(n7006), .A(n7005), .ZN(n7016) );
  OAI21_X1 U8895 ( .B1(n7010), .B2(n7009), .A(n7008), .ZN(n7014) );
  AND2_X1 U8896 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9283) );
  AOI21_X1 U8897 ( .B1(n10014), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9283), .ZN(
        n7011) );
  OAI21_X1 U8898 ( .B1(n10069), .B2(n7012), .A(n7011), .ZN(n7013) );
  AOI21_X1 U8899 ( .B1(n7014), .B2(n10081), .A(n7013), .ZN(n7015) );
  OAI21_X1 U8900 ( .B1(n7016), .B2(n10047), .A(n7015), .ZN(P1_U3252) );
  XOR2_X1 U8901 ( .A(n7018), .B(n7017), .Z(n7025) );
  AOI22_X1 U8902 ( .A1(n8336), .A2(n7354), .B1(n8341), .B2(n10299), .ZN(n7024)
         );
  INV_X2 U8903 ( .A(n7019), .ZN(n8352) );
  NOR2_X1 U8904 ( .A1(n8339), .A2(n7020), .ZN(n7021) );
  AOI211_X1 U8905 ( .C1(n7093), .C2(n8352), .A(n7022), .B(n7021), .ZN(n7023)
         );
  OAI211_X1 U8906 ( .C1(n7025), .C2(n8345), .A(n7024), .B(n7023), .ZN(P2_U3167) );
  OAI211_X1 U8907 ( .C1(n7028), .C2(n7027), .A(n7026), .B(n6606), .ZN(n7033)
         );
  NAND2_X1 U8908 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8633) );
  OAI21_X1 U8909 ( .B1(n8339), .B2(n7139), .A(n8633), .ZN(n7031) );
  OAI22_X1 U8910 ( .A1(n8355), .A2(n7029), .B1(n7265), .B2(n8350), .ZN(n7030)
         );
  AOI211_X1 U8911 ( .C1(n7216), .C2(n8352), .A(n7031), .B(n7030), .ZN(n7032)
         );
  NAND2_X1 U8912 ( .A1(n7033), .A2(n7032), .ZN(P2_U3179) );
  INV_X1 U8913 ( .A(n7353), .ZN(n10268) );
  OAI21_X1 U8914 ( .B1(n7034), .B2(n6521), .A(n7035), .ZN(n10277) );
  INV_X1 U8915 ( .A(n7036), .ZN(n7037) );
  NOR2_X1 U8916 ( .A1(n7034), .A2(n7037), .ZN(n10254) );
  AOI21_X1 U8917 ( .B1(n7037), .B2(n7034), .A(n10254), .ZN(n7041) );
  AOI22_X1 U8918 ( .A1(n10261), .A2(n8627), .B1(n6695), .B2(n10262), .ZN(n7040) );
  INV_X1 U8919 ( .A(n10265), .ZN(n7038) );
  NAND2_X1 U8920 ( .A1(n10277), .A2(n7038), .ZN(n7039) );
  OAI211_X1 U8921 ( .C1(n7041), .C2(n8871), .A(n7040), .B(n7039), .ZN(n10275)
         );
  AOI21_X1 U8922 ( .B1(n10268), .B2(n10277), .A(n10275), .ZN(n7042) );
  MUX2_X1 U8923 ( .A(n7043), .B(n7042), .S(n10269), .Z(n7046) );
  NAND2_X1 U8924 ( .A1(n8929), .A2(n7044), .ZN(n7045) );
  OAI211_X1 U8925 ( .C1(n10253), .C2(n6704), .A(n7046), .B(n7045), .ZN(
        P2_U3232) );
  INV_X1 U8926 ( .A(n7166), .ZN(n7047) );
  AOI21_X1 U8927 ( .B1(n7469), .B2(n4415), .A(n7047), .ZN(n7060) );
  INV_X1 U8928 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7048) );
  NAND2_X1 U8929 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7298) );
  OAI21_X1 U8930 ( .B1(n8654), .B2(n7048), .A(n7298), .ZN(n7049) );
  AOI21_X1 U8931 ( .B1(n7050), .B2(n8663), .A(n7049), .ZN(n7059) );
  OAI21_X1 U8932 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n7051), .A(n7182), .ZN(
        n7057) );
  NAND3_X1 U8933 ( .A1(n7054), .A2(n7053), .A3(n7052), .ZN(n7055) );
  AOI21_X1 U8934 ( .B1(n7176), .B2(n7055), .A(n8657), .ZN(n7056) );
  AOI21_X1 U8935 ( .B1(n7057), .B2(n8740), .A(n7056), .ZN(n7058) );
  OAI211_X1 U8936 ( .C1(n7060), .C2(n8756), .A(n7059), .B(n7058), .ZN(P2_U3191) );
  XNOR2_X1 U8937 ( .A(n7061), .B(n8457), .ZN(n10292) );
  INV_X1 U8938 ( .A(n10292), .ZN(n7067) );
  XOR2_X1 U8939 ( .A(n7062), .B(n8457), .Z(n7063) );
  AOI222_X1 U8940 ( .A1(n10257), .A2(n7063), .B1(n10260), .B2(n10262), .C1(
        n8625), .C2(n10261), .ZN(n10289) );
  MUX2_X1 U8941 ( .A(n7064), .B(n10289), .S(n10269), .Z(n7066) );
  AOI22_X1 U8942 ( .A1(n8929), .A2(n8289), .B1(n8942), .B2(n8292), .ZN(n7065)
         );
  OAI211_X1 U8943 ( .C1(n7067), .C2(n8932), .A(n7066), .B(n7065), .ZN(P2_U3229) );
  XOR2_X1 U8944 ( .A(n7069), .B(n7068), .Z(n10196) );
  XOR2_X1 U8945 ( .A(n7070), .B(n7069), .Z(n7072) );
  OAI22_X1 U8946 ( .A1(n7071), .A2(n9351), .B1(n7227), .B2(n9353), .ZN(n7126)
         );
  AOI21_X1 U8947 ( .B1(n7072), .B2(n10140), .A(n7126), .ZN(n10194) );
  MUX2_X1 U8948 ( .A(n10194), .B(n7073), .S(n10130), .Z(n7077) );
  INV_X1 U8949 ( .A(n10117), .ZN(n7074) );
  AOI211_X1 U8950 ( .C1(n10192), .C2(n4334), .A(n9693), .B(n7074), .ZN(n10191)
         );
  OAI22_X1 U8951 ( .A1(n9697), .A2(n7118), .B1(n9660), .B2(n7127), .ZN(n7075)
         );
  AOI21_X1 U8952 ( .B1(n10191), .B2(n10153), .A(n7075), .ZN(n7076) );
  OAI211_X1 U8953 ( .C1(n10196), .C2(n9708), .A(n7077), .B(n7076), .ZN(
        P1_U3288) );
  NOR2_X1 U8954 ( .A1(n7086), .A2(n7334), .ZN(n7079) );
  AOI211_X1 U8955 ( .C1(n10143), .C2(P1_REG3_REG_0__SCAN_IN), .A(n7079), .B(
        n7078), .ZN(n7080) );
  OAI21_X1 U8956 ( .B1(n8113), .B2(n7081), .A(n7080), .ZN(n7084) );
  INV_X1 U8957 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7082) );
  NOR2_X1 U8958 ( .A1(n9663), .A2(n7082), .ZN(n7083) );
  AOI21_X1 U8959 ( .B1(n7084), .B2(n9663), .A(n7083), .ZN(n7085) );
  OAI21_X1 U8960 ( .B1(n9667), .B2(n7086), .A(n7085), .ZN(P1_U3293) );
  INV_X1 U8961 ( .A(n7087), .ZN(n7145) );
  AOI22_X1 U8962 ( .A1(n10057), .A2(P1_STATE_REG_SCAN_IN), .B1(n7894), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n7088) );
  OAI21_X1 U8963 ( .B1(n7145), .B2(n10008), .A(n7088), .ZN(P1_U3338) );
  INV_X1 U8964 ( .A(n7090), .ZN(n7092) );
  XOR2_X1 U8965 ( .A(n4306), .B(n8388), .Z(n10296) );
  AOI22_X1 U8966 ( .A1(n8929), .A2(n10299), .B1(n8942), .B2(n7093), .ZN(n7100)
         );
  XNOR2_X1 U8967 ( .A(n7094), .B(n8388), .ZN(n7095) );
  NAND2_X1 U8968 ( .A1(n7095), .A2(n10257), .ZN(n7097) );
  AOI22_X1 U8969 ( .A1(n10262), .A2(n8626), .B1(n7354), .B2(n10261), .ZN(n7096) );
  NAND2_X1 U8970 ( .A1(n7097), .A2(n7096), .ZN(n10298) );
  MUX2_X1 U8971 ( .A(n10298), .B(P2_REG2_REG_5__SCAN_IN), .S(n10272), .Z(n7098) );
  INV_X1 U8972 ( .A(n7098), .ZN(n7099) );
  OAI211_X1 U8973 ( .C1(n10296), .C2(n8932), .A(n7100), .B(n7099), .ZN(
        P2_U3228) );
  XNOR2_X1 U8974 ( .A(n7947), .B(n8110), .ZN(n7104) );
  NAND2_X1 U8975 ( .A1(n8050), .A2(n9313), .ZN(n7102) );
  NAND2_X1 U8976 ( .A1(n9399), .A2(n9314), .ZN(n7101) );
  NAND2_X1 U8977 ( .A1(n7102), .A2(n7101), .ZN(n9176) );
  INV_X1 U8978 ( .A(n9176), .ZN(n7103) );
  OAI21_X1 U8979 ( .B1(n7104), .B2(n9642), .A(n7103), .ZN(n10181) );
  INV_X1 U8980 ( .A(n10181), .ZN(n7113) );
  XNOR2_X1 U8981 ( .A(n8110), .B(n7105), .ZN(n10183) );
  OAI211_X1 U8982 ( .C1(n10151), .C2(n10180), .A(n10148), .B(n7106), .ZN(
        n10179) );
  INV_X1 U8983 ( .A(n10179), .ZN(n7107) );
  NAND2_X1 U8984 ( .A1(n10153), .A2(n7107), .ZN(n7110) );
  AOI22_X1 U8985 ( .A1(n10130), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10143), .B2(
        n7108), .ZN(n7109) );
  OAI211_X1 U8986 ( .C1(n9697), .C2(n10180), .A(n7110), .B(n7109), .ZN(n7111)
         );
  AOI21_X1 U8987 ( .B1(n10183), .B2(n10154), .A(n7111), .ZN(n7112) );
  OAI21_X1 U8988 ( .B1(n7113), .B2(n10130), .A(n7112), .ZN(P1_U3290) );
  INV_X1 U8989 ( .A(n7114), .ZN(n7116) );
  NAND2_X1 U8990 ( .A1(n7116), .A2(n7115), .ZN(n7119) );
  OAI22_X1 U8991 ( .A1(n9352), .A2(n7791), .B1(n7118), .B2(n7801), .ZN(n7117)
         );
  XNOR2_X1 U8992 ( .A(n7117), .B(n4310), .ZN(n7120) );
  OAI22_X1 U8993 ( .A1(n9352), .A2(n9115), .B1(n7118), .B2(n7791), .ZN(n7123)
         );
  INV_X1 U8994 ( .A(n7224), .ZN(n7125) );
  AND2_X1 U8995 ( .A1(n7120), .A2(n7119), .ZN(n7121) );
  NAND2_X1 U8996 ( .A1(n7122), .A2(n7121), .ZN(n7223) );
  NAND2_X1 U8997 ( .A1(n4401), .A2(n7223), .ZN(n7124) );
  AOI22_X1 U8998 ( .A1(n7125), .A2(n7223), .B1(n7124), .B2(n7123), .ZN(n7131)
         );
  AOI22_X1 U8999 ( .A1(n9356), .A2(n7126), .B1(P1_REG3_REG_5__SCAN_IN), .B2(
        P1_U3086), .ZN(n7130) );
  INV_X1 U9000 ( .A(n7127), .ZN(n7128) );
  AOI22_X1 U9001 ( .A1(n9369), .A2(n10192), .B1(n9364), .B2(n7128), .ZN(n7129)
         );
  OAI211_X1 U9002 ( .C1(n7131), .C2(n9371), .A(n7130), .B(n7129), .ZN(P1_U3227) );
  INV_X1 U9003 ( .A(n10082), .ZN(n7133) );
  OAI222_X1 U9004 ( .A1(P1_U3086), .A2(n7133), .B1(n10005), .B2(n7132), .C1(
        n7143), .C2(n10008), .ZN(P1_U3337) );
  NAND2_X1 U9005 ( .A1(n7251), .A2(n7135), .ZN(n7136) );
  XNOR2_X1 U9006 ( .A(n7217), .B(n7354), .ZN(n8391) );
  XNOR2_X1 U9007 ( .A(n7136), .B(n8391), .ZN(n7212) );
  XNOR2_X1 U9008 ( .A(n7137), .B(n8391), .ZN(n7138) );
  OAI222_X1 U9009 ( .A1(n8910), .A2(n7265), .B1(n8908), .B2(n7139), .C1(n7138), 
        .C2(n8871), .ZN(n7213) );
  AOI21_X1 U9010 ( .B1(n10293), .B2(n7212), .A(n7213), .ZN(n7142) );
  AOI22_X1 U9011 ( .A1(n6278), .A2(n7217), .B1(n10310), .B2(
        P2_REG0_REG_6__SCAN_IN), .ZN(n7140) );
  OAI21_X1 U9012 ( .B1(n7142), .B2(n10310), .A(n7140), .ZN(P2_U3408) );
  AOI22_X1 U9013 ( .A1(n8994), .A2(n7217), .B1(n10320), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n7141) );
  OAI21_X1 U9014 ( .B1(n7142), .B2(n10320), .A(n7141), .ZN(P2_U3465) );
  INV_X1 U9015 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7144) );
  OAI222_X1 U9016 ( .A1(n9101), .A2(n7144), .B1(n8742), .B2(P2_U3151), .C1(
        n9106), .C2(n7143), .ZN(P2_U3277) );
  OAI222_X1 U9017 ( .A1(n9101), .A2(n7146), .B1(n8727), .B2(P2_U3151), .C1(
        n9106), .C2(n7145), .ZN(P2_U3278) );
  XNOR2_X1 U9018 ( .A(n7147), .B(n8119), .ZN(n10166) );
  NOR2_X1 U9019 ( .A1(n10130), .A2(n7148), .ZN(n10105) );
  INV_X1 U9020 ( .A(n10105), .ZN(n7163) );
  INV_X1 U9021 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7149) );
  OAI22_X1 U9022 ( .A1(n9663), .A2(n7150), .B1(n7149), .B2(n9660), .ZN(n7154)
         );
  AOI21_X1 U9023 ( .B1(n7155), .B2(n7151), .A(n9693), .ZN(n7152) );
  NAND2_X1 U9024 ( .A1(n7152), .A2(n10146), .ZN(n10167) );
  NOR2_X1 U9025 ( .A1(n9667), .A2(n10167), .ZN(n7153) );
  AOI211_X1 U9026 ( .C1(n10142), .C2(n7155), .A(n7154), .B(n7153), .ZN(n7162)
         );
  OAI21_X1 U9027 ( .B1(n8119), .B2(n7157), .A(n7156), .ZN(n7158) );
  NAND2_X1 U9028 ( .A1(n7158), .A2(n10140), .ZN(n7159) );
  OAI211_X1 U9029 ( .C1(n10166), .C2(n10095), .A(n7160), .B(n7159), .ZN(n10169) );
  NAND2_X1 U9030 ( .A1(n10169), .A2(n9663), .ZN(n7161) );
  OAI211_X1 U9031 ( .C1(n10166), .C2(n7163), .A(n7162), .B(n7161), .ZN(
        P1_U3292) );
  AND3_X1 U9032 ( .A1(n7166), .A2(n7165), .A3(n7164), .ZN(n7167) );
  OAI21_X1 U9033 ( .B1(n7168), .B2(n7167), .A(n8639), .ZN(n7171) );
  NAND2_X1 U9034 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7540) );
  INV_X1 U9035 ( .A(n7540), .ZN(n7169) );
  AOI21_X1 U9036 ( .B1(n8748), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7169), .ZN(
        n7170) );
  OAI211_X1 U9037 ( .C1(n8751), .C2(n7172), .A(n7171), .B(n7170), .ZN(n7187)
         );
  INV_X1 U9038 ( .A(n7173), .ZN(n7174) );
  NAND3_X1 U9039 ( .A1(n7176), .A2(n7175), .A3(n7174), .ZN(n7177) );
  AOI21_X1 U9040 ( .B1(n7178), .B2(n7177), .A(n8657), .ZN(n7186) );
  INV_X1 U9041 ( .A(n7179), .ZN(n7184) );
  NAND3_X1 U9042 ( .A1(n7182), .A2(n7181), .A3(n7180), .ZN(n7183) );
  AOI21_X1 U9043 ( .B1(n7184), .B2(n7183), .A(n8712), .ZN(n7185) );
  OR3_X1 U9044 ( .A1(n7187), .A2(n7186), .A3(n7185), .ZN(P2_U3192) );
  INV_X1 U9045 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7190) );
  NOR2_X1 U9046 ( .A1(n7188), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9164) );
  INV_X1 U9047 ( .A(n9164), .ZN(n7189) );
  OAI21_X1 U9048 ( .B1(n10089), .B2(n7190), .A(n7189), .ZN(n7195) );
  AOI211_X1 U9049 ( .C1(n7193), .C2(n7192), .A(n10030), .B(n7191), .ZN(n7194)
         );
  AOI211_X1 U9050 ( .C1(n10083), .C2(n7196), .A(n7195), .B(n7194), .ZN(n7201)
         );
  OAI211_X1 U9051 ( .C1(n7199), .C2(n7198), .A(n7197), .B(n10075), .ZN(n7200)
         );
  NAND2_X1 U9052 ( .A1(n7201), .A2(n7200), .ZN(P1_U3253) );
  INV_X1 U9053 ( .A(n7202), .ZN(n7203) );
  AOI21_X1 U9054 ( .B1(n7205), .B2(n7204), .A(n7203), .ZN(n7211) );
  AOI22_X1 U9055 ( .A1(n8336), .A2(n7355), .B1(n8341), .B2(n7350), .ZN(n7210)
         );
  NOR2_X1 U9056 ( .A1(n8339), .A2(n7206), .ZN(n7207) );
  AOI211_X1 U9057 ( .C1(n7360), .C2(n8352), .A(n7208), .B(n7207), .ZN(n7209)
         );
  OAI211_X1 U9058 ( .C1(n7211), .C2(n8345), .A(n7210), .B(n7209), .ZN(P2_U3153) );
  INV_X1 U9059 ( .A(n7212), .ZN(n7220) );
  INV_X1 U9060 ( .A(n7213), .ZN(n7214) );
  MUX2_X1 U9061 ( .A(n7215), .B(n7214), .S(n10269), .Z(n7219) );
  AOI22_X1 U9062 ( .A1(n8929), .A2(n7217), .B1(n8942), .B2(n7216), .ZN(n7218)
         );
  OAI211_X1 U9063 ( .C1(n7220), .C2(n8932), .A(n7219), .B(n7218), .ZN(P2_U3227) );
  NAND2_X1 U9064 ( .A1(n9400), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7221) );
  OAI21_X1 U9065 ( .B1(n7222), .B2(n9400), .A(n7221), .ZN(P1_U3583) );
  NAND2_X1 U9066 ( .A1(n9397), .A2(n7861), .ZN(n7225) );
  OAI21_X1 U9067 ( .B1(n10201), .B2(n7801), .A(n7225), .ZN(n7226) );
  XNOR2_X1 U9068 ( .A(n7226), .B(n4310), .ZN(n7228) );
  OAI22_X1 U9069 ( .A1(n10201), .A2(n7791), .B1(n7227), .B2(n9115), .ZN(n7229)
         );
  XNOR2_X1 U9070 ( .A(n7228), .B(n7229), .ZN(n9348) );
  NAND2_X2 U9071 ( .A1(n9347), .A2(n9348), .ZN(n9346) );
  INV_X1 U9072 ( .A(n7229), .ZN(n7230) );
  NAND2_X1 U9073 ( .A1(n7228), .A2(n7230), .ZN(n7231) );
  NAND2_X1 U9074 ( .A1(n9396), .A2(n7710), .ZN(n7232) );
  OAI21_X1 U9075 ( .B1(n10207), .B2(n7801), .A(n7232), .ZN(n7233) );
  XNOR2_X1 U9076 ( .A(n7233), .B(n9192), .ZN(n7236) );
  NAND2_X1 U9077 ( .A1(n9396), .A2(n9194), .ZN(n7234) );
  OAI21_X1 U9078 ( .B1(n10207), .B2(n7791), .A(n7234), .ZN(n7235) );
  NAND2_X1 U9079 ( .A1(n7236), .A2(n7235), .ZN(n7685) );
  NAND2_X1 U9080 ( .A1(n4407), .A2(n7685), .ZN(n7237) );
  XNOR2_X1 U9081 ( .A(n7686), .B(n7237), .ZN(n7242) );
  NAND2_X1 U9082 ( .A1(n9397), .A2(n9313), .ZN(n7239) );
  NAND2_X1 U9083 ( .A1(n9395), .A2(n9314), .ZN(n7238) );
  NAND2_X1 U9084 ( .A1(n7239), .A2(n7238), .ZN(n7325) );
  AOI22_X1 U9085 ( .A1(n9356), .A2(n7325), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n7241) );
  AOI22_X1 U9086 ( .A1(n9369), .A2(n7320), .B1(n9364), .B2(n7319), .ZN(n7240)
         );
  OAI211_X1 U9087 ( .C1(n7242), .C2(n9371), .A(n7241), .B(n7240), .ZN(P1_U3213) );
  INV_X1 U9088 ( .A(n7243), .ZN(n7878) );
  OAI222_X1 U9089 ( .A1(P1_U3086), .A2(n8151), .B1(n10008), .B2(n7878), .C1(
        n10005), .C2(n7244), .ZN(P1_U3336) );
  INV_X1 U9090 ( .A(n7246), .ZN(n7247) );
  OAI21_X1 U9091 ( .B1(n7245), .B2(n7248), .A(n7247), .ZN(n7249) );
  XNOR2_X1 U9092 ( .A(n7249), .B(n8393), .ZN(n7250) );
  AOI222_X1 U9093 ( .A1(n10257), .A2(n7250), .B1(n7539), .B2(n10261), .C1(
        n8624), .C2(n10262), .ZN(n7341) );
  INV_X1 U9094 ( .A(n7251), .ZN(n7253) );
  NAND2_X1 U9095 ( .A1(n8460), .A2(n8465), .ZN(n8498) );
  INV_X1 U9096 ( .A(n8498), .ZN(n7252) );
  AOI21_X1 U9097 ( .B1(n7253), .B2(n8465), .A(n7252), .ZN(n7352) );
  INV_X1 U9098 ( .A(n8501), .ZN(n7254) );
  NAND2_X1 U9099 ( .A1(n7352), .A2(n8392), .ZN(n7351) );
  NAND2_X1 U9100 ( .A1(n7351), .A2(n8469), .ZN(n7255) );
  XNOR2_X1 U9101 ( .A(n7255), .B(n8393), .ZN(n7336) );
  INV_X1 U9102 ( .A(n7336), .ZN(n7259) );
  INV_X1 U9103 ( .A(n7339), .ZN(n7257) );
  INV_X1 U9104 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7256) );
  OAI22_X1 U9105 ( .A1(n7257), .A2(n9078), .B1(n10308), .B2(n7256), .ZN(n7258)
         );
  AOI21_X1 U9106 ( .B1(n7259), .B2(n6198), .A(n7258), .ZN(n7260) );
  OAI21_X1 U9107 ( .B1(n7341), .B2(n10310), .A(n7260), .ZN(P2_U3414) );
  XOR2_X1 U9108 ( .A(n7262), .B(n7261), .Z(n7270) );
  NOR2_X1 U9109 ( .A1(n8350), .A2(n7263), .ZN(n7267) );
  OAI21_X1 U9110 ( .B1(n8339), .B2(n7265), .A(n7264), .ZN(n7266) );
  AOI211_X1 U9111 ( .C1(n7290), .C2(n8352), .A(n7267), .B(n7266), .ZN(n7269)
         );
  NAND2_X1 U9112 ( .A1(n8341), .A2(n7339), .ZN(n7268) );
  OAI211_X1 U9113 ( .C1(n7270), .C2(n8345), .A(n7269), .B(n7268), .ZN(P2_U3161) );
  NAND2_X1 U9114 ( .A1(n8054), .A2(n7953), .ZN(n7322) );
  OR2_X1 U9115 ( .A1(n7322), .A2(n7957), .ZN(n7324) );
  NAND2_X1 U9116 ( .A1(n7324), .A2(n7940), .ZN(n10093) );
  INV_X1 U9117 ( .A(n7941), .ZN(n7272) );
  OAI21_X1 U9118 ( .B1(n10093), .B2(n7272), .A(n7271), .ZN(n7273) );
  XNOR2_X1 U9119 ( .A(n7273), .B(n7278), .ZN(n7274) );
  NAND2_X1 U9120 ( .A1(n7274), .A2(n10140), .ZN(n7275) );
  NAND2_X1 U9121 ( .A1(n9395), .A2(n9313), .ZN(n9281) );
  NAND2_X1 U9122 ( .A1(n7275), .A2(n9281), .ZN(n10228) );
  INV_X1 U9123 ( .A(n10228), .ZN(n7288) );
  OAI21_X1 U9124 ( .B1(n7277), .B2(n10092), .A(n10090), .ZN(n7280) );
  INV_X1 U9125 ( .A(n7278), .ZN(n7279) );
  XNOR2_X1 U9126 ( .A(n7280), .B(n7279), .ZN(n10222) );
  INV_X1 U9127 ( .A(n10224), .ZN(n7281) );
  XNOR2_X1 U9128 ( .A(n10102), .B(n7281), .ZN(n7283) );
  NAND2_X1 U9129 ( .A1(n9393), .A2(n9314), .ZN(n9282) );
  INV_X1 U9130 ( .A(n9282), .ZN(n7282) );
  AOI21_X1 U9131 ( .B1(n7283), .B2(n10148), .A(n7282), .ZN(n10226) );
  OAI22_X1 U9132 ( .A1(n9663), .A2(n6344), .B1(n9285), .B2(n9660), .ZN(n7284)
         );
  AOI21_X1 U9133 ( .B1(n10142), .B2(n10224), .A(n7284), .ZN(n7285) );
  OAI21_X1 U9134 ( .B1(n10226), .B2(n9667), .A(n7285), .ZN(n7286) );
  AOI21_X1 U9135 ( .B1(n10222), .B2(n10154), .A(n7286), .ZN(n7287) );
  OAI21_X1 U9136 ( .B1(n7288), .B2(n10130), .A(n7287), .ZN(P1_U3284) );
  MUX2_X1 U9137 ( .A(n7289), .B(n7341), .S(n10269), .Z(n7292) );
  AOI22_X1 U9138 ( .A1(n8929), .A2(n7339), .B1(n8942), .B2(n7290), .ZN(n7291)
         );
  OAI211_X1 U9139 ( .C1(n7336), .C2(n8932), .A(n7292), .B(n7291), .ZN(P2_U3225) );
  INV_X1 U9140 ( .A(n7451), .ZN(n7471) );
  AOI21_X1 U9141 ( .B1(n7293), .B2(n7294), .A(n8345), .ZN(n7296) );
  NAND2_X1 U9142 ( .A1(n7296), .A2(n7295), .ZN(n7302) );
  NOR2_X1 U9143 ( .A1(n8339), .A2(n7297), .ZN(n7300) );
  OAI21_X1 U9144 ( .B1(n8350), .B2(n8482), .A(n7298), .ZN(n7299) );
  AOI211_X1 U9145 ( .C1(n7450), .C2(n8352), .A(n7300), .B(n7299), .ZN(n7301)
         );
  OAI211_X1 U9146 ( .C1(n7471), .C2(n8355), .A(n7302), .B(n7301), .ZN(P2_U3171) );
  INV_X1 U9147 ( .A(n7303), .ZN(n7333) );
  OAI222_X1 U9148 ( .A1(n9106), .A2(n7333), .B1(P2_U3151), .B2(n8613), .C1(
        n9854), .C2(n9101), .ZN(P2_U3275) );
  INV_X1 U9149 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7305) );
  AND2_X1 U9150 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9328) );
  INV_X1 U9151 ( .A(n9328), .ZN(n7304) );
  OAI21_X1 U9152 ( .B1(n10089), .B2(n7305), .A(n7304), .ZN(n7310) );
  AOI211_X1 U9153 ( .C1(n7308), .C2(n7307), .A(n10030), .B(n7306), .ZN(n7309)
         );
  AOI211_X1 U9154 ( .C1(n10083), .C2(n7311), .A(n7310), .B(n7309), .ZN(n7316)
         );
  OAI211_X1 U9155 ( .C1(n7314), .C2(n7313), .A(n7312), .B(n10075), .ZN(n7315)
         );
  NAND2_X1 U9156 ( .A1(n7316), .A2(n7315), .ZN(P1_U3254) );
  XNOR2_X1 U9157 ( .A(n7317), .B(n7957), .ZN(n10205) );
  OAI211_X1 U9158 ( .C1(n10119), .C2(n10207), .A(n10148), .B(n7318), .ZN(
        n10206) );
  AOI22_X1 U9159 ( .A1(n10142), .A2(n7320), .B1(n7319), .B2(n10143), .ZN(n7321) );
  OAI21_X1 U9160 ( .B1(n10206), .B2(n9667), .A(n7321), .ZN(n7330) );
  INV_X1 U9161 ( .A(n10095), .ZN(n7657) );
  NAND2_X1 U9162 ( .A1(n10205), .A2(n7657), .ZN(n7328) );
  NAND2_X1 U9163 ( .A1(n7322), .A2(n7957), .ZN(n7323) );
  NAND2_X1 U9164 ( .A1(n7324), .A2(n7323), .ZN(n7326) );
  AOI21_X1 U9165 ( .B1(n7326), .B2(n10140), .A(n7325), .ZN(n7327) );
  NAND2_X1 U9166 ( .A1(n7328), .A2(n7327), .ZN(n10210) );
  MUX2_X1 U9167 ( .A(n10210), .B(P1_REG2_REG_7__SCAN_IN), .S(n10130), .Z(n7329) );
  AOI211_X1 U9168 ( .C1(n10105), .C2(n10205), .A(n7330), .B(n7329), .ZN(n7331)
         );
  INV_X1 U9169 ( .A(n7331), .ZN(P1_U3286) );
  OAI222_X1 U9170 ( .A1(P1_U3086), .A2(n7334), .B1(n10008), .B2(n7333), .C1(
        n7332), .C2(n10005), .ZN(P1_U3335) );
  INV_X1 U9171 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7335) );
  NOR2_X1 U9172 ( .A1(n10323), .A2(n7335), .ZN(n7338) );
  NOR2_X1 U9173 ( .A1(n7336), .A2(n8992), .ZN(n7337) );
  AOI211_X1 U9174 ( .C1(n8994), .C2(n7339), .A(n7338), .B(n7337), .ZN(n7340)
         );
  OAI21_X1 U9175 ( .B1(n7341), .B2(n10320), .A(n7340), .ZN(P2_U3467) );
  INV_X1 U9176 ( .A(n10304), .ZN(n10282) );
  OAI21_X1 U9177 ( .B1(n7343), .B2(n6175), .A(n7342), .ZN(n7348) );
  INV_X1 U9178 ( .A(n7348), .ZN(n7447) );
  XOR2_X1 U9179 ( .A(n8396), .B(n7344), .Z(n7345) );
  NAND2_X1 U9180 ( .A1(n7345), .A2(n10257), .ZN(n7347) );
  AOI22_X1 U9181 ( .A1(n7355), .A2(n10262), .B1(n10261), .B2(n8623), .ZN(n7346) );
  OAI211_X1 U9182 ( .C1(n7348), .C2(n10265), .A(n7347), .B(n7346), .ZN(n7446)
         );
  AOI21_X1 U9183 ( .B1(n10282), .B2(n7447), .A(n7446), .ZN(n7468) );
  AOI22_X1 U9184 ( .A1(n6278), .A2(n7451), .B1(P2_REG0_REG_9__SCAN_IN), .B2(
        n10310), .ZN(n7349) );
  OAI21_X1 U9185 ( .B1(n7468), .B2(n10310), .A(n7349), .ZN(P2_U3417) );
  INV_X1 U9186 ( .A(n7350), .ZN(n10303) );
  OAI21_X1 U9187 ( .B1(n7352), .B2(n8392), .A(n7351), .ZN(n10305) );
  NOR2_X1 U9188 ( .A1(n10305), .A2(n7353), .ZN(n7359) );
  AOI22_X1 U9189 ( .A1(n7355), .A2(n10261), .B1(n10262), .B2(n7354), .ZN(n7358) );
  INV_X1 U9190 ( .A(n8392), .ZN(n8497) );
  XNOR2_X1 U9191 ( .A(n7245), .B(n8497), .ZN(n7356) );
  NAND2_X1 U9192 ( .A1(n7356), .A2(n10257), .ZN(n7357) );
  OAI211_X1 U9193 ( .C1(n10305), .C2(n10265), .A(n7358), .B(n7357), .ZN(n10307) );
  AOI211_X1 U9194 ( .C1(n8942), .C2(n7360), .A(n7359), .B(n10307), .ZN(n7361)
         );
  MUX2_X1 U9195 ( .A(n7362), .B(n7361), .S(n10269), .Z(n7363) );
  OAI21_X1 U9196 ( .B1(n10303), .B2(n8880), .A(n7363), .ZN(P2_U3226) );
  AOI21_X1 U9197 ( .B1(n4737), .B2(n4399), .A(n7493), .ZN(n7375) );
  OAI21_X1 U9198 ( .B1(n7366), .B2(n7365), .A(n7364), .ZN(n7370) );
  INV_X1 U9199 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n9848) );
  NAND2_X1 U9200 ( .A1(n8663), .A2(n7367), .ZN(n7368) );
  NAND2_X1 U9201 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7594) );
  OAI211_X1 U9202 ( .C1(n9848), .C2(n8654), .A(n7368), .B(n7594), .ZN(n7369)
         );
  AOI21_X1 U9203 ( .B1(n7370), .B2(n8753), .A(n7369), .ZN(n7374) );
  NOR2_X1 U9204 ( .A1(n7371), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7372) );
  OAI21_X1 U9205 ( .B1(n7372), .B2(n7498), .A(n8639), .ZN(n7373) );
  OAI211_X1 U9206 ( .C1(n7375), .C2(n8712), .A(n7374), .B(n7373), .ZN(P2_U3193) );
  INV_X1 U9207 ( .A(n8504), .ZN(n7376) );
  OR2_X1 U9208 ( .A1(n8476), .A2(n7376), .ZN(n8397) );
  XNOR2_X1 U9209 ( .A(n7377), .B(n8397), .ZN(n7378) );
  AOI222_X1 U9210 ( .A1(n10257), .A2(n7378), .B1(n8622), .B2(n10261), .C1(
        n7539), .C2(n10262), .ZN(n7475) );
  AOI22_X1 U9211 ( .A1(n6278), .A2(n8481), .B1(n10310), .B2(
        P2_REG0_REG_10__SCAN_IN), .ZN(n7382) );
  XOR2_X1 U9212 ( .A(n7379), .B(n8397), .Z(n7479) );
  INV_X1 U9213 ( .A(n7479), .ZN(n7380) );
  NAND2_X1 U9214 ( .A1(n7380), .A2(n6198), .ZN(n7381) );
  OAI211_X1 U9215 ( .C1(n7475), .C2(n10310), .A(n7382), .B(n7381), .ZN(
        P2_U3420) );
  INV_X1 U9216 ( .A(n7386), .ZN(n7384) );
  INV_X1 U9217 ( .A(n7393), .ZN(n8120) );
  NOR2_X1 U9218 ( .A1(n7384), .A2(n8120), .ZN(n7455) );
  INV_X1 U9219 ( .A(n7455), .ZN(n7385) );
  OAI21_X1 U9220 ( .B1(n7386), .B2(n7393), .A(n7385), .ZN(n7416) );
  INV_X1 U9221 ( .A(n7387), .ZN(n7389) );
  AOI211_X1 U9222 ( .C1(n9169), .C2(n7389), .A(n9693), .B(n7388), .ZN(n7417)
         );
  INV_X1 U9223 ( .A(n7390), .ZN(n7391) );
  AOI21_X1 U9224 ( .B1(n7393), .B2(n7392), .A(n7391), .ZN(n7395) );
  OAI22_X1 U9225 ( .A1(n7711), .A2(n9353), .B1(n9211), .B2(n9351), .ZN(n9165)
         );
  INV_X1 U9226 ( .A(n9165), .ZN(n7394) );
  OAI21_X1 U9227 ( .B1(n7395), .B2(n9642), .A(n7394), .ZN(n7423) );
  AOI211_X1 U9228 ( .C1(n7416), .C2(n10221), .A(n7417), .B(n7423), .ZN(n7400)
         );
  AOI22_X1 U9229 ( .A1(n9169), .A2(n9836), .B1(P1_REG0_REG_10__SCAN_IN), .B2(
        n10230), .ZN(n7396) );
  OAI21_X1 U9230 ( .B1(n7400), .B2(n10230), .A(n7396), .ZN(P1_U3483) );
  INV_X1 U9231 ( .A(n7397), .ZN(n7402) );
  OAI222_X1 U9232 ( .A1(n9106), .A2(n7402), .B1(P2_U3151), .B2(n8445), .C1(
        n7398), .C2(n9101), .ZN(P2_U3274) );
  AOI22_X1 U9233 ( .A1(n9169), .A2(n9771), .B1(P1_REG1_REG_10__SCAN_IN), .B2(
        n10245), .ZN(n7399) );
  OAI21_X1 U9234 ( .B1(n7400), .B2(n10245), .A(n7399), .ZN(P1_U3532) );
  OAI222_X1 U9235 ( .A1(n10005), .A2(n7403), .B1(n10008), .B2(n7402), .C1(
        n7401), .C2(P1_U3086), .ZN(P1_U3334) );
  AOI21_X1 U9236 ( .B1(n7406), .B2(n7405), .A(n7404), .ZN(n7415) );
  OAI21_X1 U9237 ( .B1(n7409), .B2(n7408), .A(n7407), .ZN(n7413) );
  NAND2_X1 U9238 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9228) );
  NAND2_X1 U9239 ( .A1(n10014), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n7410) );
  OAI211_X1 U9240 ( .C1(n10069), .C2(n7411), .A(n9228), .B(n7410), .ZN(n7412)
         );
  AOI21_X1 U9241 ( .B1(n7413), .B2(n10081), .A(n7412), .ZN(n7414) );
  OAI21_X1 U9242 ( .B1(n7415), .B2(n10047), .A(n7414), .ZN(P1_U3255) );
  INV_X1 U9243 ( .A(n7416), .ZN(n7425) );
  NAND2_X1 U9244 ( .A1(n7417), .A2(n10153), .ZN(n7420) );
  INV_X1 U9245 ( .A(n9167), .ZN(n7418) );
  AOI22_X1 U9246 ( .A1(n10130), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7418), .B2(
        n10143), .ZN(n7419) );
  OAI211_X1 U9247 ( .C1(n7421), .C2(n9697), .A(n7420), .B(n7419), .ZN(n7422)
         );
  AOI21_X1 U9248 ( .B1(n9663), .B2(n7423), .A(n7422), .ZN(n7424) );
  OAI21_X1 U9249 ( .B1(n7425), .B2(n9708), .A(n7424), .ZN(P1_U3283) );
  INV_X1 U9250 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10330) );
  INV_X1 U9251 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10073) );
  INV_X1 U9252 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7426) );
  AOI22_X1 U9253 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .B1(n10073), .B2(n7426), .ZN(n10335) );
  NOR2_X1 U9254 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(P2_ADDR_REG_16__SCAN_IN), 
        .ZN(n7427) );
  AOI21_X1 U9255 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n7427), .ZN(n10338) );
  NOR2_X1 U9256 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7428) );
  AOI21_X1 U9257 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7428), .ZN(n10341) );
  NOR2_X1 U9258 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7429) );
  AOI21_X1 U9259 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7429), .ZN(n10344) );
  NOR2_X1 U9260 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7430) );
  AOI21_X1 U9261 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7430), .ZN(n10347) );
  NOR2_X1 U9262 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7431) );
  AOI21_X1 U9263 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7431), .ZN(n10350) );
  NOR2_X1 U9264 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7432) );
  AOI21_X1 U9265 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7432), .ZN(n10353) );
  NOR2_X1 U9266 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7433) );
  AOI21_X1 U9267 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7433), .ZN(n10356) );
  NOR2_X1 U9268 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7434) );
  AOI21_X1 U9269 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7434), .ZN(n10365) );
  NOR2_X1 U9270 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7435) );
  AOI21_X1 U9271 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7435), .ZN(n10371) );
  NOR2_X1 U9272 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7436) );
  AOI21_X1 U9273 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7436), .ZN(n10368) );
  NOR2_X1 U9274 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7437) );
  AOI21_X1 U9275 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7437), .ZN(n10359) );
  NOR2_X1 U9276 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(P2_ADDR_REG_5__SCAN_IN), 
        .ZN(n7438) );
  AOI21_X1 U9277 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n7438), .ZN(n10362) );
  AND2_X1 U9278 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7439) );
  NOR2_X1 U9279 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7439), .ZN(n10325) );
  INV_X1 U9280 ( .A(n10325), .ZN(n10326) );
  NAND3_X1 U9281 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10327) );
  NAND2_X1 U9282 ( .A1(n10328), .A2(n10327), .ZN(n10324) );
  NAND2_X1 U9283 ( .A1(n10326), .A2(n10324), .ZN(n10374) );
  NAND2_X1 U9284 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7440) );
  OAI21_X1 U9285 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7440), .ZN(n10373) );
  NOR2_X1 U9286 ( .A1(n10374), .A2(n10373), .ZN(n10372) );
  AOI21_X1 U9287 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10372), .ZN(n10377) );
  NAND2_X1 U9288 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7441) );
  OAI21_X1 U9289 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7441), .ZN(n10376) );
  NOR2_X1 U9290 ( .A1(n10377), .A2(n10376), .ZN(n10375) );
  AOI21_X1 U9291 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10375), .ZN(n10380) );
  NOR2_X1 U9292 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7442) );
  AOI21_X1 U9293 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7442), .ZN(n10379) );
  NAND2_X1 U9294 ( .A1(n10380), .A2(n10379), .ZN(n10378) );
  OAI21_X1 U9295 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10378), .ZN(n10361) );
  NAND2_X1 U9296 ( .A1(n10362), .A2(n10361), .ZN(n10360) );
  OAI21_X1 U9297 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10360), .ZN(n10358) );
  NAND2_X1 U9298 ( .A1(n10359), .A2(n10358), .ZN(n10357) );
  OAI21_X1 U9299 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10357), .ZN(n10367) );
  NAND2_X1 U9300 ( .A1(n10368), .A2(n10367), .ZN(n10366) );
  OAI21_X1 U9301 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10366), .ZN(n10370) );
  NAND2_X1 U9302 ( .A1(n10371), .A2(n10370), .ZN(n10369) );
  OAI21_X1 U9303 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10369), .ZN(n10364) );
  NAND2_X1 U9304 ( .A1(n10365), .A2(n10364), .ZN(n10363) );
  OAI21_X1 U9305 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10363), .ZN(n10355) );
  NAND2_X1 U9306 ( .A1(n10356), .A2(n10355), .ZN(n10354) );
  OAI21_X1 U9307 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10354), .ZN(n10352) );
  NAND2_X1 U9308 ( .A1(n10353), .A2(n10352), .ZN(n10351) );
  OAI21_X1 U9309 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10351), .ZN(n10349) );
  NAND2_X1 U9310 ( .A1(n10350), .A2(n10349), .ZN(n10348) );
  OAI21_X1 U9311 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10348), .ZN(n10346) );
  NAND2_X1 U9312 ( .A1(n10347), .A2(n10346), .ZN(n10345) );
  OAI21_X1 U9313 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10345), .ZN(n10343) );
  NAND2_X1 U9314 ( .A1(n10344), .A2(n10343), .ZN(n10342) );
  OAI21_X1 U9315 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10342), .ZN(n10340) );
  NAND2_X1 U9316 ( .A1(n10341), .A2(n10340), .ZN(n10339) );
  OAI21_X1 U9317 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10339), .ZN(n10337) );
  NAND2_X1 U9318 ( .A1(n10338), .A2(n10337), .ZN(n10336) );
  OAI21_X1 U9319 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10336), .ZN(n10334) );
  NAND2_X1 U9320 ( .A1(n10335), .A2(n10334), .ZN(n10333) );
  OAI21_X1 U9321 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10333), .ZN(n10331) );
  NOR2_X1 U9322 ( .A1(n10330), .A2(n10331), .ZN(n7443) );
  NAND2_X1 U9323 ( .A1(n10330), .A2(n10331), .ZN(n10329) );
  OAI21_X1 U9324 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7443), .A(n10329), .ZN(
        n7445) );
  XNOR2_X1 U9325 ( .A(n4490), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7444) );
  XNOR2_X1 U9326 ( .A(n7445), .B(n7444), .ZN(ADD_1068_U4) );
  AOI21_X1 U9327 ( .B1(n10268), .B2(n7447), .A(n7446), .ZN(n7449) );
  MUX2_X1 U9328 ( .A(n7449), .B(n7448), .S(n10272), .Z(n7453) );
  AOI22_X1 U9329 ( .A1(n8929), .A2(n7451), .B1(n8942), .B2(n7450), .ZN(n7452)
         );
  NAND2_X1 U9330 ( .A1(n7453), .A2(n7452), .ZN(P2_U3224) );
  NOR2_X1 U9331 ( .A1(n7455), .A2(n7454), .ZN(n7456) );
  INV_X1 U9332 ( .A(n7457), .ZN(n8126) );
  XNOR2_X1 U9333 ( .A(n7456), .B(n8126), .ZN(n7551) );
  XNOR2_X1 U9334 ( .A(n7458), .B(n7457), .ZN(n7459) );
  NOR2_X1 U9335 ( .A1(n7459), .A2(n9642), .ZN(n7461) );
  OAI22_X1 U9336 ( .A1(n7977), .A2(n9353), .B1(n7460), .B2(n9351), .ZN(n9329)
         );
  AOI211_X1 U9337 ( .C1(n7551), .C2(n7657), .A(n7461), .B(n9329), .ZN(n7548)
         );
  MUX2_X1 U9338 ( .A(n7462), .B(n7548), .S(n9663), .Z(n7467) );
  OAI211_X1 U9339 ( .C1(n7388), .C2(n9333), .A(n10148), .B(n7463), .ZN(n7547)
         );
  NOR2_X1 U9340 ( .A1(n7547), .A2(n9667), .ZN(n7465) );
  OAI22_X1 U9341 ( .A1(n9333), .A2(n9697), .B1(n9326), .B2(n9660), .ZN(n7464)
         );
  AOI211_X1 U9342 ( .C1(n7551), .C2(n10105), .A(n7465), .B(n7464), .ZN(n7466)
         );
  NAND2_X1 U9343 ( .A1(n7467), .A2(n7466), .ZN(P1_U3282) );
  MUX2_X1 U9344 ( .A(n7469), .B(n7468), .S(n10323), .Z(n7470) );
  OAI21_X1 U9345 ( .B1(n7471), .B2(n6292), .A(n7470), .ZN(P2_U3468) );
  MUX2_X1 U9346 ( .A(n7472), .B(n7475), .S(n10269), .Z(n7474) );
  AOI22_X1 U9347 ( .A1(n8481), .A2(n8929), .B1(n8942), .B2(n7544), .ZN(n7473)
         );
  OAI211_X1 U9348 ( .C1(n7479), .C2(n8932), .A(n7474), .B(n7473), .ZN(P2_U3223) );
  MUX2_X1 U9349 ( .A(n7476), .B(n7475), .S(n10323), .Z(n7478) );
  NAND2_X1 U9350 ( .A1(n8481), .A2(n8994), .ZN(n7477) );
  OAI211_X1 U9351 ( .C1(n7479), .C2(n8992), .A(n7478), .B(n7477), .ZN(P2_U3469) );
  INV_X1 U9352 ( .A(n7480), .ZN(n7484) );
  OAI222_X1 U9353 ( .A1(n10005), .A2(n7482), .B1(n10008), .B2(n7484), .C1(
        P1_U3086), .C2(n7481), .ZN(P1_U3333) );
  OAI222_X1 U9354 ( .A1(n8187), .A2(n7485), .B1(n9106), .B2(n7484), .C1(n7483), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  INV_X1 U9355 ( .A(n7486), .ZN(n7488) );
  NAND2_X1 U9356 ( .A1(n7488), .A2(n7487), .ZN(n7489) );
  XNOR2_X1 U9357 ( .A(n7490), .B(n7489), .ZN(n7508) );
  OR3_X1 U9358 ( .A1(n7493), .A2(n7492), .A3(n7491), .ZN(n7494) );
  AOI21_X1 U9359 ( .B1(n7495), .B2(n7494), .A(n8712), .ZN(n7502) );
  OR3_X1 U9360 ( .A1(n7498), .A2(n7497), .A3(n7496), .ZN(n7499) );
  AOI21_X1 U9361 ( .B1(n7500), .B2(n7499), .A(n8756), .ZN(n7501) );
  NOR2_X1 U9362 ( .A1(n7502), .A2(n7501), .ZN(n7507) );
  INV_X1 U9363 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7503) );
  NAND2_X1 U9364 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7883) );
  OAI21_X1 U9365 ( .B1(n8654), .B2(n7503), .A(n7883), .ZN(n7504) );
  AOI21_X1 U9366 ( .B1(n7505), .B2(n8663), .A(n7504), .ZN(n7506) );
  OAI211_X1 U9367 ( .C1(n8657), .C2(n7508), .A(n7507), .B(n7506), .ZN(P2_U3194) );
  XNOR2_X1 U9368 ( .A(n7510), .B(n7509), .ZN(n7511) );
  AOI22_X1 U9369 ( .A1(n9392), .A2(n9313), .B1(n9314), .B2(n9390), .ZN(n9229)
         );
  OAI21_X1 U9370 ( .B1(n7511), .B2(n9642), .A(n9229), .ZN(n7566) );
  INV_X1 U9371 ( .A(n7566), .ZN(n7520) );
  OAI21_X1 U9372 ( .B1(n7513), .B2(n8124), .A(n7512), .ZN(n7568) );
  INV_X1 U9373 ( .A(n7463), .ZN(n7514) );
  OAI211_X1 U9374 ( .C1(n7514), .C2(n9234), .A(n10148), .B(n7528), .ZN(n7565)
         );
  AOI22_X1 U9375 ( .A1(n10130), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9231), .B2(
        n10143), .ZN(n7517) );
  NAND2_X1 U9376 ( .A1(n7515), .A2(n10142), .ZN(n7516) );
  OAI211_X1 U9377 ( .C1(n7565), .C2(n9667), .A(n7517), .B(n7516), .ZN(n7518)
         );
  AOI21_X1 U9378 ( .B1(n7568), .B2(n10154), .A(n7518), .ZN(n7519) );
  OAI21_X1 U9379 ( .B1(n7520), .B2(n10130), .A(n7519), .ZN(P1_U3281) );
  INV_X1 U9380 ( .A(n7653), .ZN(n7523) );
  INV_X1 U9381 ( .A(n7530), .ZN(n8127) );
  AOI21_X1 U9382 ( .B1(n7521), .B2(n7974), .A(n8127), .ZN(n7522) );
  OAI21_X1 U9383 ( .B1(n7523), .B2(n7522), .A(n10140), .ZN(n7526) );
  NAND2_X1 U9384 ( .A1(n9389), .A2(n9314), .ZN(n7525) );
  NAND2_X1 U9385 ( .A1(n9391), .A2(n9313), .ZN(n7524) );
  AND2_X1 U9386 ( .A1(n7525), .A2(n7524), .ZN(n9305) );
  NAND2_X1 U9387 ( .A1(n7526), .A2(n9305), .ZN(n7606) );
  INV_X1 U9388 ( .A(n7658), .ZN(n7527) );
  AOI211_X1 U9389 ( .C1(n9307), .C2(n7528), .A(n9693), .B(n7527), .ZN(n7602)
         );
  NOR2_X1 U9390 ( .A1(n7606), .A2(n7602), .ZN(n7538) );
  AOI22_X1 U9391 ( .A1(n9307), .A2(n9836), .B1(P1_REG0_REG_13__SCAN_IN), .B2(
        n10230), .ZN(n7534) );
  OAI21_X1 U9392 ( .B1(n7531), .B2(n7530), .A(n7529), .ZN(n7601) );
  NAND2_X1 U9393 ( .A1(n10232), .A2(n10221), .ZN(n9838) );
  INV_X1 U9394 ( .A(n9838), .ZN(n7532) );
  NAND2_X1 U9395 ( .A1(n7601), .A2(n7532), .ZN(n7533) );
  OAI211_X1 U9396 ( .C1(n7538), .C2(n10230), .A(n7534), .B(n7533), .ZN(
        P1_U3492) );
  AOI22_X1 U9397 ( .A1(n9307), .A2(n9771), .B1(P1_REG1_REG_13__SCAN_IN), .B2(
        n10245), .ZN(n7537) );
  NAND2_X1 U9398 ( .A1(n10248), .A2(n10221), .ZN(n9773) );
  INV_X1 U9399 ( .A(n9773), .ZN(n7535) );
  NAND2_X1 U9400 ( .A1(n7601), .A2(n7535), .ZN(n7536) );
  OAI211_X1 U9401 ( .C1(n7538), .C2(n10245), .A(n7537), .B(n7536), .ZN(
        P1_U3535) );
  XNOR2_X1 U9402 ( .A(n7589), .B(n8623), .ZN(n7591) );
  XOR2_X1 U9403 ( .A(n7590), .B(n7591), .Z(n7546) );
  NAND2_X1 U9404 ( .A1(n8348), .A2(n7539), .ZN(n7541) );
  OAI211_X1 U9405 ( .C1(n8484), .C2(n8350), .A(n7541), .B(n7540), .ZN(n7543)
         );
  INV_X1 U9406 ( .A(n8481), .ZN(n8480) );
  NOR2_X1 U9407 ( .A1(n8480), .A2(n8355), .ZN(n7542) );
  AOI211_X1 U9408 ( .C1(n7544), .C2(n8352), .A(n7543), .B(n7542), .ZN(n7545)
         );
  OAI21_X1 U9409 ( .B1(n7546), .B2(n8345), .A(n7545), .ZN(P2_U3157) );
  INV_X1 U9410 ( .A(n9779), .ZN(n10219) );
  INV_X1 U9411 ( .A(n7547), .ZN(n7550) );
  INV_X1 U9412 ( .A(n7548), .ZN(n7549) );
  AOI211_X1 U9413 ( .C1(n10219), .C2(n7551), .A(n7550), .B(n7549), .ZN(n7555)
         );
  AOI22_X1 U9414 ( .A1(n7553), .A2(n9836), .B1(P1_REG0_REG_11__SCAN_IN), .B2(
        n10230), .ZN(n7552) );
  OAI21_X1 U9415 ( .B1(n7555), .B2(n10230), .A(n7552), .ZN(P1_U3486) );
  AOI22_X1 U9416 ( .A1(n7553), .A2(n9771), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n10245), .ZN(n7554) );
  OAI21_X1 U9417 ( .B1(n7555), .B2(n10245), .A(n7554), .ZN(P1_U3533) );
  XNOR2_X1 U9418 ( .A(n7556), .B(n8399), .ZN(n7557) );
  NAND2_X1 U9419 ( .A1(n7557), .A2(n10257), .ZN(n7559) );
  AOI22_X1 U9420 ( .A1(n10262), .A2(n8623), .B1(n8621), .B2(n10261), .ZN(n7558) );
  NAND2_X1 U9421 ( .A1(n7559), .A2(n7558), .ZN(n9002) );
  AOI21_X1 U9422 ( .B1(n8942), .B2(n7597), .A(n9002), .ZN(n7560) );
  MUX2_X1 U9423 ( .A(n4737), .B(n7560), .S(n10269), .Z(n7564) );
  NAND2_X1 U9424 ( .A1(n7644), .A2(n8399), .ZN(n7582) );
  OR2_X1 U9425 ( .A1(n7644), .A2(n8399), .ZN(n7562) );
  NAND2_X1 U9426 ( .A1(n7582), .A2(n7562), .ZN(n8998) );
  AOI22_X1 U9427 ( .A1(n8998), .A2(n8945), .B1(n8929), .B2(n8997), .ZN(n7563)
         );
  NAND2_X1 U9428 ( .A1(n7564), .A2(n7563), .ZN(P2_U3222) );
  OAI21_X1 U9429 ( .B1(n9234), .B2(n10213), .A(n7565), .ZN(n7567) );
  AOI211_X1 U9430 ( .C1(n10221), .C2(n7568), .A(n7567), .B(n7566), .ZN(n7571)
         );
  NAND2_X1 U9431 ( .A1(n10230), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7569) );
  OAI21_X1 U9432 ( .B1(n7571), .B2(n10230), .A(n7569), .ZN(P1_U3489) );
  NAND2_X1 U9433 ( .A1(n10245), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7570) );
  OAI21_X1 U9434 ( .B1(n7571), .B2(n10245), .A(n7570), .ZN(P1_U3534) );
  NAND2_X1 U9435 ( .A1(n7576), .A2(n7572), .ZN(n7573) );
  OAI211_X1 U9436 ( .C1(n7574), .C2(n7913), .A(n7573), .B(n8162), .ZN(P1_U3332) );
  NAND2_X1 U9437 ( .A1(n7576), .A2(n7575), .ZN(n7578) );
  OR2_X1 U9438 ( .A1(n7577), .A2(P2_U3151), .ZN(n8609) );
  OAI211_X1 U9439 ( .C1(n7579), .C2(n9101), .A(n7578), .B(n8609), .ZN(P2_U3272) );
  XNOR2_X1 U9440 ( .A(n7580), .B(n7583), .ZN(n7581) );
  OAI222_X1 U9441 ( .A1(n8910), .A2(n8194), .B1(n8908), .B2(n8484), .C1(n7581), 
        .C2(n8871), .ZN(n7835) );
  AOI21_X1 U9442 ( .B1(n8942), .B2(n7886), .A(n7835), .ZN(n7588) );
  NAND2_X1 U9443 ( .A1(n7582), .A2(n8505), .ZN(n7584) );
  INV_X1 U9444 ( .A(n7583), .ZN(n8509) );
  XNOR2_X1 U9445 ( .A(n7584), .B(n8509), .ZN(n7841) );
  OAI22_X1 U9446 ( .A1(n6176), .A2(n8880), .B1(n7585), .B2(n10269), .ZN(n7586)
         );
  AOI21_X1 U9447 ( .B1(n7841), .B2(n8945), .A(n7586), .ZN(n7587) );
  OAI21_X1 U9448 ( .B1(n7588), .B2(n10272), .A(n7587), .ZN(P2_U3221) );
  OAI22_X1 U9449 ( .A1(n7591), .A2(n7590), .B1(n8623), .B2(n7589), .ZN(n7592)
         );
  XOR2_X1 U9450 ( .A(n7593), .B(n7592), .Z(n7600) );
  NAND2_X1 U9451 ( .A1(n8348), .A2(n8623), .ZN(n7595) );
  OAI211_X1 U9452 ( .C1(n8310), .C2(n8350), .A(n7595), .B(n7594), .ZN(n7596)
         );
  AOI21_X1 U9453 ( .B1(n7597), .B2(n8352), .A(n7596), .ZN(n7599) );
  NAND2_X1 U9454 ( .A1(n8997), .A2(n8341), .ZN(n7598) );
  OAI211_X1 U9455 ( .C1(n7600), .C2(n8345), .A(n7599), .B(n7598), .ZN(P2_U3176) );
  INV_X1 U9456 ( .A(n7601), .ZN(n7608) );
  NAND2_X1 U9457 ( .A1(n7602), .A2(n10153), .ZN(n7604) );
  AOI22_X1 U9458 ( .A1(n10130), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9302), .B2(
        n10143), .ZN(n7603) );
  OAI211_X1 U9459 ( .C1(n7728), .C2(n9697), .A(n7604), .B(n7603), .ZN(n7605)
         );
  AOI21_X1 U9460 ( .B1(n9663), .B2(n7606), .A(n7605), .ZN(n7607) );
  OAI21_X1 U9461 ( .B1(n7608), .B2(n9708), .A(n7607), .ZN(P1_U3280) );
  NAND2_X1 U9462 ( .A1(n10014), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n7609) );
  NAND2_X1 U9463 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9303) );
  NAND2_X1 U9464 ( .A1(n7609), .A2(n9303), .ZN(n7614) );
  AOI211_X1 U9465 ( .C1(n7612), .C2(n7611), .A(n10030), .B(n7610), .ZN(n7613)
         );
  AOI211_X1 U9466 ( .C1(n10083), .C2(n7615), .A(n7614), .B(n7613), .ZN(n7620)
         );
  OAI211_X1 U9467 ( .C1(n7618), .C2(n7617), .A(n7616), .B(n10075), .ZN(n7619)
         );
  NAND2_X1 U9468 ( .A1(n7620), .A2(n7619), .ZN(P1_U3256) );
  INV_X1 U9469 ( .A(n7621), .ZN(n7624) );
  OAI222_X1 U9470 ( .A1(n9106), .A2(n7624), .B1(P2_U3151), .B2(n6153), .C1(
        n7622), .C2(n9101), .ZN(P2_U3271) );
  OAI222_X1 U9471 ( .A1(n7625), .A2(P1_U3086), .B1(n10008), .B2(n7624), .C1(
        n7623), .C2(n10005), .ZN(P1_U3331) );
  XOR2_X1 U9472 ( .A(n7626), .B(n8130), .Z(n9839) );
  INV_X1 U9473 ( .A(n9363), .ZN(n7630) );
  OAI21_X1 U9474 ( .B1(n4948), .B2(n5629), .A(n7627), .ZN(n7629) );
  AOI22_X1 U9475 ( .A1(n9387), .A2(n9314), .B1(n9313), .B2(n9389), .ZN(n9367)
         );
  INV_X1 U9476 ( .A(n9367), .ZN(n7628) );
  AOI21_X1 U9477 ( .B1(n7629), .B2(n10140), .A(n7628), .ZN(n9769) );
  OAI21_X1 U9478 ( .B1(n7630), .B2(n9660), .A(n9769), .ZN(n7634) );
  INV_X1 U9479 ( .A(n9835), .ZN(n7631) );
  NAND2_X1 U9480 ( .A1(n7670), .A2(n7631), .ZN(n9694) );
  OAI211_X1 U9481 ( .C1(n7670), .C2(n7631), .A(n9694), .B(n10148), .ZN(n9768)
         );
  AOI22_X1 U9482 ( .A1(n9835), .A2(n10142), .B1(P1_REG2_REG_15__SCAN_IN), .B2(
        n10130), .ZN(n7632) );
  OAI21_X1 U9483 ( .B1(n9768), .B2(n9667), .A(n7632), .ZN(n7633) );
  AOI21_X1 U9484 ( .B1(n7634), .B2(n9663), .A(n7633), .ZN(n7635) );
  OAI21_X1 U9485 ( .B1(n9839), .B2(n9708), .A(n7635), .ZN(P1_U3278) );
  NAND2_X1 U9486 ( .A1(n7637), .A2(n7636), .ZN(n8513) );
  INV_X1 U9487 ( .A(n8513), .ZN(n7638) );
  XNOR2_X1 U9488 ( .A(n7639), .B(n7638), .ZN(n7640) );
  NAND2_X1 U9489 ( .A1(n7640), .A2(n10257), .ZN(n7642) );
  AOI22_X1 U9490 ( .A1(n10261), .A2(n8925), .B1(n8621), .B2(n10262), .ZN(n7641) );
  NAND2_X1 U9491 ( .A1(n7642), .A2(n7641), .ZN(n7890) );
  MUX2_X1 U9492 ( .A(n7890), .B(P2_REG0_REG_13__SCAN_IN), .S(n10310), .Z(n7649) );
  NAND2_X1 U9493 ( .A1(n7644), .A2(n7643), .ZN(n7645) );
  AND2_X1 U9494 ( .A1(n7646), .A2(n7645), .ZN(n7647) );
  XNOR2_X1 U9495 ( .A(n7647), .B(n8513), .ZN(n7893) );
  OAI22_X1 U9496 ( .A1(n7893), .A2(n9088), .B1(n8311), .B2(n9078), .ZN(n7648)
         );
  OR2_X1 U9497 ( .A1(n7649), .A2(n7648), .ZN(P2_U3429) );
  MUX2_X1 U9498 ( .A(n7890), .B(P2_REG1_REG_13__SCAN_IN), .S(n10320), .Z(n7651) );
  OAI22_X1 U9499 ( .A1(n7893), .A2(n8992), .B1(n8311), .B2(n6292), .ZN(n7650)
         );
  OR2_X1 U9500 ( .A1(n7651), .A2(n7650), .ZN(P2_U3472) );
  XNOR2_X1 U9501 ( .A(n7652), .B(n7985), .ZN(n9774) );
  NAND2_X1 U9502 ( .A1(n7653), .A2(n8064), .ZN(n7654) );
  XNOR2_X1 U9503 ( .A(n7654), .B(n7985), .ZN(n7655) );
  AOI22_X1 U9504 ( .A1(n9314), .A2(n9388), .B1(n9390), .B2(n9313), .ZN(n9138)
         );
  OAI21_X1 U9505 ( .B1(n7655), .B2(n9642), .A(n9138), .ZN(n7656) );
  AOI21_X1 U9506 ( .B1(n9774), .B2(n7657), .A(n7656), .ZN(n9778) );
  AOI211_X1 U9507 ( .C1(n9776), .C2(n7658), .A(n9693), .B(n7670), .ZN(n9775)
         );
  NAND2_X1 U9508 ( .A1(n9775), .A2(n10153), .ZN(n7660) );
  AOI22_X1 U9509 ( .A1(n10130), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9140), .B2(
        n10143), .ZN(n7659) );
  OAI211_X1 U9510 ( .C1(n9143), .C2(n9697), .A(n7660), .B(n7659), .ZN(n7661)
         );
  AOI21_X1 U9511 ( .B1(n10105), .B2(n9774), .A(n7661), .ZN(n7662) );
  OAI21_X1 U9512 ( .B1(n9778), .B2(n10130), .A(n7662), .ZN(P1_U3279) );
  INV_X1 U9513 ( .A(n7663), .ZN(n10007) );
  OAI222_X1 U9514 ( .A1(n9106), .A2(n10007), .B1(P2_U3151), .B2(n7665), .C1(
        n7664), .C2(n9101), .ZN(P2_U3270) );
  XNOR2_X1 U9515 ( .A(n7666), .B(n7993), .ZN(n9831) );
  NAND2_X1 U9516 ( .A1(n9699), .A2(n8075), .ZN(n7667) );
  XNOR2_X1 U9517 ( .A(n7667), .B(n7993), .ZN(n7668) );
  AOI22_X1 U9518 ( .A1(n9385), .A2(n9314), .B1(n9313), .B2(n9387), .ZN(n9255)
         );
  OAI21_X1 U9519 ( .B1(n7668), .B2(n9642), .A(n9255), .ZN(n9759) );
  INV_X1 U9520 ( .A(n9828), .ZN(n9260) );
  NAND2_X1 U9521 ( .A1(n7670), .A2(n7669), .ZN(n9691) );
  NAND2_X1 U9522 ( .A1(n9691), .A2(n9828), .ZN(n7671) );
  NAND2_X1 U9523 ( .A1(n7671), .A2(n10148), .ZN(n7672) );
  NOR2_X1 U9524 ( .A1(n9673), .A2(n7672), .ZN(n9758) );
  NAND2_X1 U9525 ( .A1(n9758), .A2(n10153), .ZN(n7675) );
  INV_X1 U9526 ( .A(n7673), .ZN(n9257) );
  AOI22_X1 U9527 ( .A1(n10130), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9257), .B2(
        n10143), .ZN(n7674) );
  OAI211_X1 U9528 ( .C1(n9260), .C2(n9697), .A(n7675), .B(n7674), .ZN(n7676)
         );
  AOI21_X1 U9529 ( .B1(n9759), .B2(n9663), .A(n7676), .ZN(n7677) );
  OAI21_X1 U9530 ( .B1(n9831), .B2(n9708), .A(n7677), .ZN(P1_U3276) );
  INV_X1 U9531 ( .A(n7678), .ZN(n9105) );
  OAI222_X1 U9532 ( .A1(n7680), .A2(P1_U3086), .B1(n10008), .B2(n9105), .C1(
        n7679), .C2(n10005), .ZN(P1_U3329) );
  NAND2_X1 U9533 ( .A1(n9558), .A2(n9189), .ZN(n7682) );
  NAND2_X1 U9534 ( .A1(n9378), .A2(n7861), .ZN(n7681) );
  NAND2_X1 U9535 ( .A1(n7682), .A2(n7681), .ZN(n7683) );
  XNOR2_X1 U9536 ( .A(n7683), .B(n4310), .ZN(n7857) );
  OAI22_X1 U9537 ( .A1(n9722), .A2(n7791), .B1(n7684), .B2(n9115), .ZN(n7855)
         );
  XNOR2_X1 U9538 ( .A(n7857), .B(n7855), .ZN(n7826) );
  NAND2_X1 U9539 ( .A1(n10224), .A2(n9189), .ZN(n7688) );
  NAND2_X1 U9540 ( .A1(n9394), .A2(n7861), .ZN(n7687) );
  NAND2_X1 U9541 ( .A1(n7688), .A2(n7687), .ZN(n7689) );
  XNOR2_X1 U9542 ( .A(n7689), .B(n4310), .ZN(n9277) );
  NOR2_X1 U9543 ( .A1(n9211), .A2(n9115), .ZN(n7690) );
  AOI21_X1 U9544 ( .B1(n10224), .B2(n7861), .A(n7690), .ZN(n7698) );
  NAND2_X1 U9545 ( .A1(n9277), .A2(n7698), .ZN(n7697) );
  NAND2_X1 U9546 ( .A1(n10101), .A2(n9189), .ZN(n7692) );
  NAND2_X1 U9547 ( .A1(n9395), .A2(n7861), .ZN(n7691) );
  NAND2_X1 U9548 ( .A1(n7692), .A2(n7691), .ZN(n7693) );
  XNOR2_X1 U9549 ( .A(n7693), .B(n9192), .ZN(n9275) );
  NAND2_X1 U9550 ( .A1(n10101), .A2(n7861), .ZN(n7695) );
  NAND2_X1 U9551 ( .A1(n9395), .A2(n9194), .ZN(n7694) );
  NAND2_X1 U9552 ( .A1(n7695), .A2(n7694), .ZN(n9207) );
  INV_X1 U9553 ( .A(n7698), .ZN(n9276) );
  AOI21_X1 U9554 ( .B1(n9275), .B2(n9207), .A(n9276), .ZN(n7700) );
  NAND3_X1 U9555 ( .A1(n9275), .A2(n9276), .A3(n9207), .ZN(n7699) );
  OAI21_X1 U9556 ( .B1(n7700), .B2(n9277), .A(n7699), .ZN(n7701) );
  INV_X1 U9557 ( .A(n7701), .ZN(n7702) );
  NAND2_X1 U9558 ( .A1(n9169), .A2(n9189), .ZN(n7704) );
  NAND2_X1 U9559 ( .A1(n9393), .A2(n7861), .ZN(n7703) );
  NAND2_X1 U9560 ( .A1(n7704), .A2(n7703), .ZN(n7705) );
  XNOR2_X1 U9561 ( .A(n7705), .B(n9192), .ZN(n7714) );
  NAND2_X1 U9562 ( .A1(n9169), .A2(n7861), .ZN(n7707) );
  NAND2_X1 U9563 ( .A1(n9393), .A2(n9194), .ZN(n7706) );
  NAND2_X1 U9564 ( .A1(n7707), .A2(n7706), .ZN(n9163) );
  OR2_X1 U9565 ( .A1(n7714), .A2(n9163), .ZN(n7708) );
  NAND2_X1 U9566 ( .A1(n9159), .A2(n7708), .ZN(n7717) );
  OAI22_X1 U9567 ( .A1(n9333), .A2(n7801), .B1(n7711), .B2(n7791), .ZN(n7709)
         );
  XOR2_X1 U9568 ( .A(n4310), .B(n7709), .Z(n7713) );
  INV_X1 U9569 ( .A(n7710), .ZN(n7791) );
  OAI22_X1 U9570 ( .A1(n9333), .A2(n7791), .B1(n7711), .B2(n9115), .ZN(n7712)
         );
  NOR2_X1 U9571 ( .A1(n7713), .A2(n7712), .ZN(n7718) );
  AOI21_X1 U9572 ( .B1(n7713), .B2(n7712), .A(n7718), .ZN(n9322) );
  INV_X1 U9573 ( .A(n7714), .ZN(n9160) );
  INV_X1 U9574 ( .A(n9163), .ZN(n7715) );
  INV_X1 U9575 ( .A(n7718), .ZN(n9225) );
  OAI22_X1 U9576 ( .A1(n9234), .A2(n7801), .B1(n7977), .B2(n7791), .ZN(n7719)
         );
  XNOR2_X1 U9577 ( .A(n7719), .B(n4310), .ZN(n7721) );
  OAI22_X1 U9578 ( .A1(n9234), .A2(n7791), .B1(n7977), .B2(n9115), .ZN(n7722)
         );
  INV_X1 U9579 ( .A(n7722), .ZN(n7720) );
  NAND2_X1 U9580 ( .A1(n7721), .A2(n7720), .ZN(n7725) );
  INV_X1 U9581 ( .A(n7721), .ZN(n7723) );
  NAND2_X1 U9582 ( .A1(n7723), .A2(n7722), .ZN(n7724) );
  NAND2_X1 U9583 ( .A1(n7725), .A2(n7724), .ZN(n9224) );
  INV_X1 U9584 ( .A(n7725), .ZN(n7726) );
  OAI22_X1 U9585 ( .A1(n7728), .A2(n7791), .B1(n7727), .B2(n9115), .ZN(n7730)
         );
  OAI22_X1 U9586 ( .A1(n7728), .A2(n7801), .B1(n7727), .B2(n7791), .ZN(n7729)
         );
  XNOR2_X1 U9587 ( .A(n7729), .B(n4310), .ZN(n7732) );
  XOR2_X1 U9588 ( .A(n7730), .B(n7732), .Z(n9301) );
  INV_X1 U9589 ( .A(n7730), .ZN(n7731) );
  NAND2_X1 U9590 ( .A1(n9776), .A2(n9189), .ZN(n7734) );
  NAND2_X1 U9591 ( .A1(n9389), .A2(n7861), .ZN(n7733) );
  NAND2_X1 U9592 ( .A1(n7734), .A2(n7733), .ZN(n7735) );
  XNOR2_X1 U9593 ( .A(n7735), .B(n4310), .ZN(n7743) );
  NAND2_X1 U9594 ( .A1(n9776), .A2(n7861), .ZN(n7737) );
  NAND2_X1 U9595 ( .A1(n9389), .A2(n9194), .ZN(n7736) );
  NAND2_X1 U9596 ( .A1(n9835), .A2(n9189), .ZN(n7739) );
  NAND2_X1 U9597 ( .A1(n9388), .A2(n7861), .ZN(n7738) );
  NAND2_X1 U9598 ( .A1(n7739), .A2(n7738), .ZN(n7740) );
  XNOR2_X1 U9599 ( .A(n7740), .B(n9192), .ZN(n7756) );
  NAND2_X1 U9600 ( .A1(n9835), .A2(n7710), .ZN(n7742) );
  NAND2_X1 U9601 ( .A1(n9388), .A2(n9194), .ZN(n7741) );
  NAND2_X1 U9602 ( .A1(n7742), .A2(n7741), .ZN(n9362) );
  INV_X1 U9603 ( .A(n7743), .ZN(n9134) );
  INV_X1 U9604 ( .A(n9136), .ZN(n7744) );
  OAI22_X1 U9605 ( .A1(n7756), .A2(n9362), .B1(n9134), .B2(n7744), .ZN(n7745)
         );
  INV_X1 U9606 ( .A(n7745), .ZN(n7746) );
  NAND2_X1 U9607 ( .A1(n9764), .A2(n9189), .ZN(n7748) );
  NAND2_X1 U9608 ( .A1(n9387), .A2(n7861), .ZN(n7747) );
  NAND2_X1 U9609 ( .A1(n7748), .A2(n7747), .ZN(n7749) );
  XNOR2_X1 U9610 ( .A(n7749), .B(n4310), .ZN(n7753) );
  INV_X1 U9611 ( .A(n7753), .ZN(n7755) );
  NOR2_X1 U9612 ( .A1(n7750), .A2(n9115), .ZN(n7751) );
  AOI21_X1 U9613 ( .B1(n9764), .B2(n7861), .A(n7751), .ZN(n7752) );
  INV_X1 U9614 ( .A(n7752), .ZN(n7754) );
  AND2_X1 U9615 ( .A1(n7753), .A2(n7752), .ZN(n7760) );
  AOI21_X1 U9616 ( .B1(n7755), .B2(n7754), .A(n7760), .ZN(n9242) );
  INV_X1 U9617 ( .A(n7756), .ZN(n9238) );
  INV_X1 U9618 ( .A(n9362), .ZN(n7757) );
  INV_X1 U9619 ( .A(n7760), .ZN(n7761) );
  AOI22_X1 U9620 ( .A1(n9828), .A2(n7861), .B1(n9194), .B2(n9386), .ZN(n7766)
         );
  NAND2_X1 U9621 ( .A1(n9828), .A2(n9189), .ZN(n7763) );
  NAND2_X1 U9622 ( .A1(n9386), .A2(n7710), .ZN(n7762) );
  NAND2_X1 U9623 ( .A1(n7763), .A2(n7762), .ZN(n7764) );
  XNOR2_X1 U9624 ( .A(n7764), .B(n4310), .ZN(n7765) );
  XOR2_X1 U9625 ( .A(n7766), .B(n7765), .Z(n9253) );
  NAND2_X1 U9626 ( .A1(n9754), .A2(n9189), .ZN(n7769) );
  NAND2_X1 U9627 ( .A1(n9385), .A2(n7861), .ZN(n7768) );
  NAND2_X1 U9628 ( .A1(n7769), .A2(n7768), .ZN(n7770) );
  XNOR2_X1 U9629 ( .A(n7770), .B(n9192), .ZN(n7774) );
  NAND2_X1 U9630 ( .A1(n9754), .A2(n7861), .ZN(n7772) );
  NAND2_X1 U9631 ( .A1(n9385), .A2(n9194), .ZN(n7771) );
  NAND2_X1 U9632 ( .A1(n7772), .A2(n7771), .ZN(n7773) );
  NOR2_X1 U9633 ( .A1(n7774), .A2(n7773), .ZN(n9334) );
  NAND2_X1 U9634 ( .A1(n7774), .A2(n7773), .ZN(n9335) );
  NAND2_X1 U9635 ( .A1(n9822), .A2(n9189), .ZN(n7776) );
  NAND2_X1 U9636 ( .A1(n9384), .A2(n7861), .ZN(n7775) );
  NAND2_X1 U9637 ( .A1(n7776), .A2(n7775), .ZN(n7777) );
  XNOR2_X1 U9638 ( .A(n7777), .B(n4310), .ZN(n7780) );
  AND2_X1 U9639 ( .A1(n9384), .A2(n9194), .ZN(n7778) );
  AOI21_X1 U9640 ( .B1(n9822), .B2(n7861), .A(n7778), .ZN(n7779) );
  NOR2_X1 U9641 ( .A1(n7780), .A2(n7779), .ZN(n9180) );
  AOI22_X1 U9642 ( .A1(n9816), .A2(n9189), .B1(n7861), .B2(n9383), .ZN(n7781)
         );
  XNOR2_X1 U9643 ( .A(n7781), .B(n4310), .ZN(n7783) );
  OAI22_X1 U9644 ( .A1(n4808), .A2(n7791), .B1(n8108), .B2(n9115), .ZN(n7782)
         );
  NOR2_X1 U9645 ( .A1(n7783), .A2(n7782), .ZN(n7784) );
  AOI21_X1 U9646 ( .B1(n7783), .B2(n7782), .A(n7784), .ZN(n9293) );
  INV_X1 U9647 ( .A(n7784), .ZN(n7785) );
  NAND2_X1 U9648 ( .A1(n9291), .A2(n7785), .ZN(n9216) );
  NAND2_X1 U9649 ( .A1(n7786), .A2(n9189), .ZN(n7788) );
  OR2_X1 U9650 ( .A1(n7790), .A2(n7791), .ZN(n7787) );
  NAND2_X1 U9651 ( .A1(n7788), .A2(n7787), .ZN(n7789) );
  XNOR2_X1 U9652 ( .A(n7789), .B(n4310), .ZN(n7792) );
  OAI22_X1 U9653 ( .A1(n9813), .A2(n7791), .B1(n7790), .B2(n9115), .ZN(n7793)
         );
  XNOR2_X1 U9654 ( .A(n7792), .B(n7793), .ZN(n9217) );
  INV_X1 U9655 ( .A(n7793), .ZN(n7794) );
  NAND2_X1 U9656 ( .A1(n9806), .A2(n9189), .ZN(n7797) );
  NAND2_X1 U9657 ( .A1(n9381), .A2(n7861), .ZN(n7796) );
  NAND2_X1 U9658 ( .A1(n7797), .A2(n7796), .ZN(n7798) );
  XNOR2_X1 U9659 ( .A(n7798), .B(n9192), .ZN(n9144) );
  NAND2_X1 U9660 ( .A1(n9806), .A2(n7861), .ZN(n7800) );
  NAND2_X1 U9661 ( .A1(n9381), .A2(n9194), .ZN(n7799) );
  NAND2_X1 U9662 ( .A1(n7800), .A2(n7799), .ZN(n9312) );
  NOR2_X1 U9663 ( .A1(n9144), .A2(n9312), .ZN(n7808) );
  OAI22_X1 U9664 ( .A1(n9598), .A2(n7801), .B1(n7803), .B2(n7791), .ZN(n7802)
         );
  XOR2_X1 U9665 ( .A(n4310), .B(n7802), .Z(n7805) );
  OAI22_X1 U9666 ( .A1(n9598), .A2(n7791), .B1(n7803), .B2(n9115), .ZN(n7804)
         );
  AOI21_X1 U9667 ( .B1(n7805), .B2(n7804), .A(n9262), .ZN(n9149) );
  NAND2_X1 U9668 ( .A1(n9144), .A2(n9312), .ZN(n7806) );
  OAI21_X2 U9669 ( .B1(n9146), .B2(n7808), .A(n7807), .ZN(n9150) );
  INV_X1 U9670 ( .A(n9262), .ZN(n7820) );
  NAND2_X1 U9671 ( .A1(n9150), .A2(n7820), .ZN(n7854) );
  NAND2_X1 U9672 ( .A1(n9578), .A2(n9189), .ZN(n7810) );
  NAND2_X1 U9673 ( .A1(n9379), .A2(n7861), .ZN(n7809) );
  NAND2_X1 U9674 ( .A1(n7810), .A2(n7809), .ZN(n7811) );
  XNOR2_X1 U9675 ( .A(n7811), .B(n4310), .ZN(n7813) );
  AND2_X1 U9676 ( .A1(n9379), .A2(n9194), .ZN(n7812) );
  AOI21_X1 U9677 ( .B1(n9578), .B2(n7861), .A(n7812), .ZN(n7814) );
  NAND2_X1 U9678 ( .A1(n7813), .A2(n7814), .ZN(n7818) );
  INV_X1 U9679 ( .A(n7813), .ZN(n7816) );
  INV_X1 U9680 ( .A(n7814), .ZN(n7815) );
  NAND2_X1 U9681 ( .A1(n7816), .A2(n7815), .ZN(n7817) );
  NAND2_X1 U9682 ( .A1(n7854), .A2(n9261), .ZN(n9264) );
  NAND2_X1 U9683 ( .A1(n9264), .A2(n7818), .ZN(n7825) );
  INV_X1 U9684 ( .A(n7826), .ZN(n7819) );
  AND2_X1 U9685 ( .A1(n7820), .A2(n7858), .ZN(n7821) );
  NAND2_X1 U9686 ( .A1(n9150), .A2(n7821), .ZN(n7824) );
  INV_X1 U9687 ( .A(n7858), .ZN(n7822) );
  AND2_X1 U9688 ( .A1(n9261), .A2(n7826), .ZN(n7853) );
  OR2_X1 U9689 ( .A1(n7822), .A2(n7853), .ZN(n7823) );
  OAI21_X1 U9690 ( .B1(n7826), .B2(n7825), .A(n7868), .ZN(n7827) );
  NAND2_X1 U9691 ( .A1(n7827), .A2(n9349), .ZN(n7834) );
  NAND2_X1 U9692 ( .A1(n9377), .A2(n9314), .ZN(n7829) );
  NAND2_X1 U9693 ( .A1(n9379), .A2(n9313), .ZN(n7828) );
  NAND2_X1 U9694 ( .A1(n7829), .A2(n7828), .ZN(n9554) );
  INV_X1 U9695 ( .A(n7830), .ZN(n9556) );
  OAI22_X1 U9696 ( .A1(n9556), .A2(n9342), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7831), .ZN(n7832) );
  AOI21_X1 U9697 ( .B1(n9554), .B2(n9356), .A(n7832), .ZN(n7833) );
  OAI211_X1 U9698 ( .C1(n9722), .C2(n9332), .A(n7834), .B(n7833), .ZN(P1_U3225) );
  INV_X1 U9699 ( .A(n7835), .ZN(n7838) );
  MUX2_X1 U9700 ( .A(n9908), .B(n7838), .S(n10323), .Z(n7837) );
  AOI22_X1 U9701 ( .A1(n7841), .A2(n6511), .B1(n8994), .B2(n7840), .ZN(n7836)
         );
  NAND2_X1 U9702 ( .A1(n7837), .A2(n7836), .ZN(P2_U3471) );
  INV_X1 U9703 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7839) );
  MUX2_X1 U9704 ( .A(n7839), .B(n7838), .S(n10308), .Z(n7843) );
  AOI22_X1 U9705 ( .A1(n7841), .A2(n6198), .B1(n6278), .B2(n7840), .ZN(n7842)
         );
  NAND2_X1 U9706 ( .A1(n7843), .A2(n7842), .ZN(P2_U3426) );
  OAI21_X1 U9707 ( .B1(n7852), .B2(n9838), .A(n7848), .ZN(P1_U3518) );
  OAI21_X1 U9708 ( .B1(n7852), .B2(n9773), .A(n7851), .ZN(P1_U3550) );
  INV_X1 U9709 ( .A(n9546), .ZN(n9789) );
  NAND2_X1 U9710 ( .A1(n7854), .A2(n7853), .ZN(n7860) );
  INV_X1 U9711 ( .A(n7855), .ZN(n7856) );
  NAND2_X1 U9712 ( .A1(n7857), .A2(n7856), .ZN(n7866) );
  AND2_X1 U9713 ( .A1(n7858), .A2(n7866), .ZN(n7859) );
  AND2_X1 U9714 ( .A1(n7860), .A2(n7859), .ZN(n7870) );
  NAND2_X1 U9715 ( .A1(n9546), .A2(n9189), .ZN(n7863) );
  NAND2_X1 U9716 ( .A1(n9377), .A2(n7861), .ZN(n7862) );
  NAND2_X1 U9717 ( .A1(n7863), .A2(n7862), .ZN(n7864) );
  XNOR2_X1 U9718 ( .A(n7864), .B(n9192), .ZN(n9110) );
  AND2_X1 U9719 ( .A1(n9377), .A2(n9194), .ZN(n7865) );
  AOI21_X1 U9720 ( .B1(n9546), .B2(n7861), .A(n7865), .ZN(n9108) );
  XNOR2_X1 U9721 ( .A(n9110), .B(n9108), .ZN(n7869) );
  OAI211_X1 U9722 ( .C1(n7870), .C2(n7869), .A(n9349), .B(n9127), .ZN(n7877)
         );
  OR2_X1 U9723 ( .A1(n9116), .A2(n9353), .ZN(n7872) );
  NAND2_X1 U9724 ( .A1(n9378), .A2(n9313), .ZN(n7871) );
  NAND2_X1 U9725 ( .A1(n7872), .A2(n7871), .ZN(n9535) );
  INV_X1 U9726 ( .A(n7873), .ZN(n9541) );
  OAI22_X1 U9727 ( .A1(n9541), .A2(n9342), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7874), .ZN(n7875) );
  AOI21_X1 U9728 ( .B1(n9535), .B2(n9356), .A(n7875), .ZN(n7876) );
  OAI211_X1 U9729 ( .C1(n9789), .C2(n9332), .A(n7877), .B(n7876), .ZN(P1_U3240) );
  INV_X1 U9730 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7879) );
  OAI222_X1 U9731 ( .A1(n9101), .A2(n7879), .B1(n9106), .B2(n7878), .C1(n6194), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  OAI211_X1 U9732 ( .C1(n7882), .C2(n7881), .A(n7880), .B(n6606), .ZN(n7888)
         );
  NAND2_X1 U9733 ( .A1(n8348), .A2(n8622), .ZN(n7884) );
  OAI211_X1 U9734 ( .C1(n8194), .C2(n8350), .A(n7884), .B(n7883), .ZN(n7885)
         );
  AOI21_X1 U9735 ( .B1(n7886), .B2(n8352), .A(n7885), .ZN(n7887) );
  OAI211_X1 U9736 ( .C1(n6176), .C2(n8355), .A(n7888), .B(n7887), .ZN(P2_U3164) );
  NOR2_X1 U9737 ( .A1(n8311), .A2(n10251), .ZN(n7889) );
  OAI21_X1 U9738 ( .B1(n7890), .B2(n7889), .A(n10269), .ZN(n7892) );
  AOI22_X1 U9739 ( .A1(n10272), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8942), .B2(
        n8314), .ZN(n7891) );
  OAI211_X1 U9740 ( .C1(n7893), .C2(n8932), .A(n7892), .B(n7891), .ZN(P2_U3220) );
  NAND2_X1 U9741 ( .A1(n7894), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7899) );
  INV_X1 U9742 ( .A(n7895), .ZN(n7897) );
  INV_X1 U9743 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n7896) );
  NAND4_X1 U9744 ( .A1(n7897), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .A4(n7896), .ZN(n7898) );
  OAI211_X1 U9745 ( .C1(n8361), .C2(n10008), .A(n7899), .B(n7898), .ZN(
        P1_U3324) );
  INV_X1 U9746 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n7901) );
  NAND4_X1 U9747 ( .A1(n4307), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .A4(n7901), .ZN(n7904) );
  NAND2_X1 U9748 ( .A1(n7902), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n7903) );
  OAI211_X1 U9749 ( .C1(n8361), .C2(n9106), .A(n7904), .B(n7903), .ZN(P2_U3264) );
  INV_X1 U9750 ( .A(n9709), .ZN(n7905) );
  NAND2_X1 U9751 ( .A1(n9663), .A2(n7905), .ZN(n9500) );
  NAND2_X1 U9752 ( .A1(n10130), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n7906) );
  OAI211_X1 U9753 ( .C1(n8169), .C2(n9697), .A(n9500), .B(n7906), .ZN(n7907)
         );
  INV_X1 U9754 ( .A(n7907), .ZN(n7908) );
  OAI21_X1 U9755 ( .B1(n7909), .B2(n9667), .A(n7908), .ZN(P1_U3263) );
  INV_X1 U9756 ( .A(n7910), .ZN(n8185) );
  OAI222_X1 U9757 ( .A1(n7913), .A2(n7912), .B1(n10008), .B2(n8185), .C1(n7911), .C2(P1_U3086), .ZN(P1_U3325) );
  NOR2_X1 U9758 ( .A1(n10269), .A2(n7915), .ZN(n7917) );
  NOR2_X1 U9759 ( .A1(n7916), .A2(n10253), .ZN(n8759) );
  AOI211_X1 U9760 ( .C1(n7918), .C2(n8929), .A(n7917), .B(n8759), .ZN(n7921)
         );
  NAND2_X1 U9761 ( .A1(n7919), .A2(n8945), .ZN(n7920) );
  OAI211_X1 U9762 ( .C1(n7914), .C2(n10272), .A(n7921), .B(n7920), .ZN(
        P2_U3204) );
  OAI21_X1 U9763 ( .B1(n8169), .B2(n9374), .A(n9373), .ZN(n8040) );
  NAND2_X1 U9764 ( .A1(n8002), .A2(n8000), .ZN(n8081) );
  INV_X1 U9765 ( .A(n8039), .ZN(n8168) );
  MUX2_X1 U9766 ( .A(n7922), .B(n8081), .S(n8168), .Z(n8005) );
  NAND2_X1 U9767 ( .A1(n8076), .A2(n9680), .ZN(n8131) );
  NAND2_X1 U9768 ( .A1(n8131), .A2(n7925), .ZN(n7933) );
  NAND2_X1 U9769 ( .A1(n9384), .A2(n8039), .ZN(n7932) );
  OAI21_X1 U9770 ( .B1(n7933), .B2(n8168), .A(n7932), .ZN(n7923) );
  AND2_X1 U9771 ( .A1(n7923), .A2(n4810), .ZN(n7935) );
  NAND3_X1 U9772 ( .A1(n8109), .A2(n8168), .A3(n8076), .ZN(n7926) );
  NAND2_X1 U9773 ( .A1(n9340), .A2(n8168), .ZN(n7928) );
  NAND2_X1 U9774 ( .A1(n7926), .A2(n7928), .ZN(n7927) );
  NAND2_X1 U9775 ( .A1(n7927), .A2(n9822), .ZN(n7931) );
  INV_X1 U9776 ( .A(n7928), .ZN(n7929) );
  NAND3_X1 U9777 ( .A1(n8109), .A2(n7929), .A3(n8076), .ZN(n7930) );
  OAI211_X1 U9778 ( .C1(n7933), .C2(n7932), .A(n7931), .B(n7930), .ZN(n7934)
         );
  NAND2_X1 U9779 ( .A1(n10108), .A2(n7953), .ZN(n7939) );
  NAND2_X1 U9780 ( .A1(n7939), .A2(n7938), .ZN(n7944) );
  INV_X1 U9781 ( .A(n7957), .ZN(n7943) );
  NAND2_X1 U9782 ( .A1(n7941), .A2(n7940), .ZN(n7942) );
  AOI21_X1 U9783 ( .B1(n7944), .B2(n7943), .A(n7942), .ZN(n7946) );
  NAND2_X1 U9784 ( .A1(n7947), .A2(n10124), .ZN(n7950) );
  NAND3_X1 U9785 ( .A1(n7950), .A2(n7949), .A3(n7948), .ZN(n7952) );
  NAND3_X1 U9786 ( .A1(n7952), .A2(n8111), .A3(n7951), .ZN(n7955) );
  INV_X1 U9787 ( .A(n7953), .ZN(n7954) );
  AOI21_X1 U9788 ( .B1(n7955), .B2(n8114), .A(n7954), .ZN(n7958) );
  OAI21_X1 U9789 ( .B1(n7958), .B2(n7957), .A(n7956), .ZN(n7961) );
  INV_X1 U9790 ( .A(n7959), .ZN(n7960) );
  NAND2_X1 U9791 ( .A1(n7961), .A2(n7960), .ZN(n7962) );
  NAND3_X1 U9792 ( .A1(n7966), .A2(n8062), .A3(n7973), .ZN(n7967) );
  INV_X1 U9793 ( .A(n8062), .ZN(n7968) );
  AOI21_X1 U9794 ( .B1(n7970), .B2(n7969), .A(n7968), .ZN(n7976) );
  NAND2_X1 U9795 ( .A1(n7972), .A2(n7971), .ZN(n8061) );
  NAND2_X1 U9796 ( .A1(n7974), .A2(n7973), .ZN(n8066) );
  INV_X1 U9797 ( .A(n8066), .ZN(n7975) );
  NOR2_X1 U9798 ( .A1(n9391), .A2(n8039), .ZN(n7979) );
  OAI21_X1 U9799 ( .B1(n7977), .B2(n8168), .A(n9234), .ZN(n7978) );
  OAI21_X1 U9800 ( .B1(n9234), .B2(n7979), .A(n7978), .ZN(n7980) );
  AND2_X1 U9801 ( .A1(n7990), .A2(n7991), .ZN(n8071) );
  NAND3_X1 U9802 ( .A1(n7982), .A2(n8071), .A3(n8068), .ZN(n7984) );
  NAND2_X1 U9803 ( .A1(n7990), .A2(n4553), .ZN(n7983) );
  INV_X1 U9804 ( .A(n7985), .ZN(n8128) );
  NAND2_X1 U9805 ( .A1(n8128), .A2(n8069), .ZN(n7986) );
  AOI21_X1 U9806 ( .B1(n7987), .B2(n8064), .A(n7986), .ZN(n7992) );
  NAND2_X1 U9807 ( .A1(n7989), .A2(n7988), .ZN(n8072) );
  AND2_X1 U9808 ( .A1(n7990), .A2(n8039), .ZN(n7994) );
  OAI211_X1 U9809 ( .C1(n7992), .C2(n8072), .A(n7994), .B(n7991), .ZN(n7999)
         );
  INV_X1 U9810 ( .A(n7993), .ZN(n7997) );
  INV_X1 U9811 ( .A(n7994), .ZN(n7995) );
  OR2_X1 U9812 ( .A1(n7995), .A2(n8075), .ZN(n7996) );
  AND4_X1 U9813 ( .A1(n8077), .A2(n7997), .A3(n4384), .A4(n7996), .ZN(n7998)
         );
  MUX2_X1 U9814 ( .A(n8003), .B(n8002), .S(n8039), .Z(n8004) );
  INV_X1 U9815 ( .A(n9604), .ZN(n8006) );
  NAND2_X1 U9816 ( .A1(n8007), .A2(n8006), .ZN(n8011) );
  AND2_X1 U9817 ( .A1(n9563), .A2(n8008), .ZN(n8085) );
  INV_X1 U9818 ( .A(n8085), .ZN(n8009) );
  NAND2_X1 U9819 ( .A1(n8009), .A2(n8168), .ZN(n8010) );
  NAND2_X1 U9820 ( .A1(n8011), .A2(n8010), .ZN(n8013) );
  AOI21_X1 U9821 ( .B1(n8044), .B2(n9588), .A(n8168), .ZN(n8012) );
  AOI21_X1 U9822 ( .B1(n8013), .B2(n8044), .A(n8012), .ZN(n8018) );
  NOR2_X1 U9823 ( .A1(n9563), .A2(n8168), .ZN(n8014) );
  NAND2_X1 U9824 ( .A1(n9578), .A2(n8015), .ZN(n8086) );
  MUX2_X1 U9825 ( .A(n8086), .B(n9550), .S(n8039), .Z(n8016) );
  NAND2_X1 U9826 ( .A1(n8021), .A2(n8020), .ZN(n8089) );
  OAI21_X1 U9827 ( .B1(n8023), .B2(n8022), .A(n8021), .ZN(n8024) );
  NAND2_X1 U9828 ( .A1(n8027), .A2(n8025), .ZN(n8093) );
  INV_X1 U9829 ( .A(n8093), .ZN(n8026) );
  NAND2_X1 U9830 ( .A1(n8027), .A2(n8168), .ZN(n8028) );
  AOI21_X1 U9831 ( .B1(n8019), .B2(n8047), .A(n8089), .ZN(n8031) );
  NAND3_X1 U9832 ( .A1(n8080), .A2(n8168), .A3(n8079), .ZN(n8030) );
  NAND3_X1 U9833 ( .A1(n9715), .A2(n9116), .A3(n8168), .ZN(n8029) );
  OAI211_X1 U9834 ( .C1(n8031), .C2(n8030), .A(n8029), .B(n8042), .ZN(n8032)
         );
  OAI21_X1 U9835 ( .B1(n8039), .B2(n8042), .A(n8032), .ZN(n8033) );
  NAND3_X1 U9836 ( .A1(n8034), .A2(n9508), .A3(n8033), .ZN(n8036) );
  MUX2_X1 U9837 ( .A(n8043), .B(n8097), .S(n8039), .Z(n8035) );
  INV_X1 U9838 ( .A(n9373), .ZN(n8037) );
  INV_X1 U9839 ( .A(n8169), .ZN(n8147) );
  OAI21_X1 U9840 ( .B1(n8037), .B2(n9374), .A(n8147), .ZN(n8038) );
  AOI21_X1 U9841 ( .B1(n8041), .B2(n8159), .A(n7401), .ZN(n8183) );
  OAI211_X1 U9842 ( .C1(n8045), .C2(n9588), .A(n9550), .B(n8044), .ZN(n8046)
         );
  NAND2_X1 U9843 ( .A1(n8046), .A2(n8086), .ZN(n8048) );
  NAND2_X1 U9844 ( .A1(n8048), .A2(n8047), .ZN(n8088) );
  NOR2_X1 U9845 ( .A1(n8094), .A2(n8088), .ZN(n8145) );
  NAND2_X1 U9846 ( .A1(n9402), .A2(n10168), .ZN(n8049) );
  NAND3_X1 U9847 ( .A1(n8111), .A2(n4312), .A3(n8049), .ZN(n8057) );
  INV_X1 U9848 ( .A(n8050), .ZN(n8053) );
  OAI211_X1 U9849 ( .C1(n8053), .C2(n10147), .A(n8052), .B(n8051), .ZN(n8056)
         );
  INV_X1 U9850 ( .A(n8054), .ZN(n8055) );
  OAI21_X1 U9851 ( .B1(n8057), .B2(n8056), .A(n8055), .ZN(n8058) );
  INV_X1 U9852 ( .A(n8058), .ZN(n8060) );
  OAI21_X1 U9853 ( .B1(n8060), .B2(n8122), .A(n8059), .ZN(n8063) );
  AOI21_X1 U9854 ( .B1(n8063), .B2(n8062), .A(n8061), .ZN(n8067) );
  OAI211_X1 U9855 ( .C1(n8067), .C2(n8066), .A(n8065), .B(n8064), .ZN(n8070)
         );
  AND3_X1 U9856 ( .A1(n8070), .A2(n8069), .A3(n8068), .ZN(n8073) );
  OAI21_X1 U9857 ( .B1(n8073), .B2(n8072), .A(n8071), .ZN(n8074) );
  AOI21_X1 U9858 ( .B1(n8075), .B2(n8074), .A(n8131), .ZN(n8078) );
  OAI211_X1 U9859 ( .C1(n8078), .C2(n8109), .A(n8077), .B(n8076), .ZN(n8082)
         );
  AOI211_X1 U9860 ( .C1(n8083), .C2(n8082), .A(n8081), .B(n8142), .ZN(n8100)
         );
  INV_X1 U9861 ( .A(n9605), .ZN(n8084) );
  AND3_X1 U9862 ( .A1(n8086), .A2(n8085), .A3(n8084), .ZN(n8087) );
  NOR2_X1 U9863 ( .A1(n8088), .A2(n8087), .ZN(n8090) );
  NOR2_X1 U9864 ( .A1(n8090), .A2(n8089), .ZN(n8091) );
  NOR2_X1 U9865 ( .A1(n8142), .A2(n8091), .ZN(n8092) );
  OR2_X1 U9866 ( .A1(n8093), .A2(n8092), .ZN(n8096) );
  INV_X1 U9867 ( .A(n9374), .ZN(n8101) );
  NAND2_X1 U9868 ( .A1(n9503), .A2(n8101), .ZN(n8140) );
  NAND2_X1 U9869 ( .A1(n8099), .A2(n8098), .ZN(n8149) );
  AOI21_X1 U9870 ( .B1(n8145), .B2(n8100), .A(n8149), .ZN(n8103) );
  OR2_X1 U9871 ( .A1(n9503), .A2(n8101), .ZN(n8102) );
  NAND2_X1 U9872 ( .A1(n8169), .A2(n9373), .ZN(n8170) );
  OAI21_X1 U9873 ( .B1(n8103), .B2(n8107), .A(n8170), .ZN(n8104) );
  MUX2_X1 U9874 ( .A(n8106), .B(n8105), .S(n8104), .Z(n8163) );
  INV_X1 U9875 ( .A(n8163), .ZN(n8166) );
  INV_X1 U9876 ( .A(n8162), .ZN(n8152) );
  INV_X1 U9877 ( .A(n8107), .ZN(n8153) );
  INV_X1 U9878 ( .A(n9587), .ZN(n9589) );
  XNOR2_X1 U9879 ( .A(n9816), .B(n8108), .ZN(n9639) );
  INV_X1 U9880 ( .A(n9624), .ZN(n9620) );
  INV_X1 U9881 ( .A(n8109), .ZN(n8133) );
  INV_X1 U9882 ( .A(n8110), .ZN(n8112) );
  NAND4_X1 U9883 ( .A1(n8113), .A2(n8112), .A3(n7401), .A4(n8111), .ZN(n8116)
         );
  INV_X1 U9884 ( .A(n8114), .ZN(n8115) );
  NOR3_X1 U9885 ( .A1(n8116), .A2(n8115), .A3(n10145), .ZN(n8118) );
  INV_X1 U9886 ( .A(n10133), .ZN(n8117) );
  NAND4_X1 U9887 ( .A1(n8120), .A2(n8119), .A3(n8118), .A4(n8117), .ZN(n8121)
         );
  NOR4_X1 U9888 ( .A1(n8124), .A2(n8123), .A3(n8122), .A4(n8121), .ZN(n8125)
         );
  NAND4_X1 U9889 ( .A1(n8128), .A2(n8127), .A3(n8126), .A4(n8125), .ZN(n8129)
         );
  NOR4_X1 U9890 ( .A1(n8131), .A2(n9690), .A3(n8130), .A4(n8129), .ZN(n8132)
         );
  NAND4_X1 U9891 ( .A1(n9620), .A2(n8133), .A3(n9657), .A4(n8132), .ZN(n8134)
         );
  NOR4_X1 U9892 ( .A1(n9589), .A2(n9639), .A3(n9604), .A4(n8134), .ZN(n8136)
         );
  INV_X1 U9893 ( .A(n9571), .ZN(n8135) );
  NAND4_X1 U9894 ( .A1(n9537), .A2(n9552), .A3(n8136), .A4(n8135), .ZN(n8137)
         );
  NOR4_X1 U9895 ( .A1(n8139), .A2(n8138), .A3(n5639), .A4(n8137), .ZN(n8141)
         );
  NAND4_X1 U9896 ( .A1(n8153), .A2(n8141), .A3(n8170), .A4(n8140), .ZN(n8156)
         );
  NAND4_X1 U9897 ( .A1(n8166), .A2(n8175), .A3(n8152), .A4(n8156), .ZN(n8182)
         );
  INV_X1 U9898 ( .A(n8142), .ZN(n8144) );
  INV_X1 U9899 ( .A(n8143), .ZN(n9606) );
  NAND3_X1 U9900 ( .A1(n8145), .A2(n8144), .A3(n9606), .ZN(n8146) );
  OAI211_X1 U9901 ( .C1(n8147), .C2(n9784), .A(n8146), .B(n8170), .ZN(n8150)
         );
  OAI21_X1 U9902 ( .B1(n8150), .B2(n8149), .A(n8148), .ZN(n8155) );
  OAI211_X1 U9903 ( .C1(n8153), .C2(n8169), .A(n8152), .B(n8151), .ZN(n8154)
         );
  AOI21_X1 U9904 ( .B1(n8156), .B2(n8155), .A(n8154), .ZN(n8167) );
  NOR4_X1 U9905 ( .A1(n9351), .A2(n8158), .A3(n10002), .A4(n8157), .ZN(n8161)
         );
  NOR2_X1 U9906 ( .A1(n8162), .A2(n8159), .ZN(n8173) );
  INV_X1 U9907 ( .A(P1_B_REG_SCAN_IN), .ZN(n8160) );
  NOR3_X1 U9908 ( .A1(n8161), .A2(n8173), .A3(n8160), .ZN(n8165) );
  NOR3_X1 U9909 ( .A1(n8163), .A2(n8171), .A3(n8162), .ZN(n8164) );
  NOR3_X1 U9910 ( .A1(n8169), .A2(n8168), .A3(n9373), .ZN(n8178) );
  INV_X1 U9911 ( .A(n8170), .ZN(n8176) );
  NAND3_X1 U9912 ( .A1(n8173), .A2(n4312), .A3(n8171), .ZN(n8174) );
  AOI21_X1 U9913 ( .B1(n8176), .B2(n8175), .A(n8174), .ZN(n8177) );
  OAI211_X1 U9914 ( .C1(n8183), .C2(n8182), .A(n8181), .B(n8180), .ZN(P1_U3242) );
  OAI222_X1 U9915 ( .A1(n9101), .A2(n8357), .B1(n9106), .B2(n8185), .C1(
        P2_U3151), .C2(n8184), .ZN(P2_U3265) );
  INV_X1 U9916 ( .A(n8186), .ZN(n8190) );
  OAI222_X1 U9917 ( .A1(n9106), .A2(n8190), .B1(n6498), .B2(P2_U3151), .C1(
        n8188), .C2(n8187), .ZN(P2_U3267) );
  OAI222_X1 U9918 ( .A1(n10005), .A2(n9842), .B1(n10008), .B2(n8190), .C1(
        n8189), .C2(P1_U3086), .ZN(P1_U3327) );
  XOR2_X1 U9919 ( .A(n8192), .B(n8191), .Z(n8198) );
  NAND2_X1 U9920 ( .A1(n8336), .A2(n8936), .ZN(n8193) );
  NAND2_X1 U9921 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8672) );
  OAI211_X1 U9922 ( .C1(n8194), .C2(n8339), .A(n8193), .B(n8672), .ZN(n8196)
         );
  NOR2_X1 U9923 ( .A1(n8933), .A2(n8355), .ZN(n8195) );
  AOI211_X1 U9924 ( .C1(n8941), .C2(n8352), .A(n8196), .B(n8195), .ZN(n8197)
         );
  OAI21_X1 U9925 ( .B1(n8198), .B2(n8345), .A(n8197), .ZN(P2_U3155) );
  XNOR2_X1 U9926 ( .A(n8278), .B(n8321), .ZN(n8203) );
  NAND2_X1 U9927 ( .A1(n8805), .A2(n8336), .ZN(n8200) );
  AOI22_X1 U9928 ( .A1(n8808), .A2(n8352), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8199) );
  OAI211_X1 U9929 ( .C1(n8243), .C2(n8339), .A(n8200), .B(n8199), .ZN(n8201)
         );
  AOI21_X1 U9930 ( .B1(n9042), .B2(n8341), .A(n8201), .ZN(n8202) );
  OAI21_X1 U9931 ( .B1(n8203), .B2(n8345), .A(n8202), .ZN(P2_U3156) );
  AOI21_X1 U9932 ( .B1(n8205), .B2(n8204), .A(n8345), .ZN(n8207) );
  NAND2_X1 U9933 ( .A1(n8207), .A2(n8206), .ZN(n8216) );
  AOI22_X1 U9934 ( .A1(n8336), .A2(n8626), .B1(n8341), .B2(n8208), .ZN(n8215)
         );
  INV_X1 U9935 ( .A(n8209), .ZN(n8212) );
  NOR2_X1 U9936 ( .A1(n8339), .A2(n8210), .ZN(n8211) );
  AOI211_X1 U9937 ( .C1(n8213), .C2(n8352), .A(n8212), .B(n8211), .ZN(n8214)
         );
  NAND3_X1 U9938 ( .A1(n8216), .A2(n8215), .A3(n8214), .ZN(P2_U3158) );
  INV_X1 U9939 ( .A(n8976), .ZN(n8225) );
  AOI21_X1 U9940 ( .B1(n8217), .B2(n8218), .A(n8345), .ZN(n8220) );
  NAND2_X1 U9941 ( .A1(n8220), .A2(n8219), .ZN(n8224) );
  NAND2_X1 U9942 ( .A1(n8833), .A2(n8336), .ZN(n8221) );
  NAND2_X1 U9943 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8750) );
  OAI211_X1 U9944 ( .C1(n8893), .C2(n8339), .A(n8221), .B(n8750), .ZN(n8222)
         );
  AOI21_X1 U9945 ( .B1(n8863), .B2(n8352), .A(n8222), .ZN(n8223) );
  OAI211_X1 U9946 ( .C1(n8225), .C2(n8355), .A(n8224), .B(n8223), .ZN(P2_U3159) );
  INV_X1 U9947 ( .A(n8226), .ZN(n8227) );
  XNOR2_X1 U9948 ( .A(n8412), .B(n8229), .ZN(n8230) );
  XNOR2_X1 U9949 ( .A(n8231), .B(n8230), .ZN(n8238) );
  NOR2_X1 U9950 ( .A1(n8569), .A2(n8350), .ZN(n8236) );
  AOI22_X1 U9951 ( .A1(n8232), .A2(n8352), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8233) );
  OAI21_X1 U9952 ( .B1(n8234), .B2(n8339), .A(n8233), .ZN(n8235) );
  AOI211_X1 U9953 ( .C1(n8576), .C2(n8341), .A(n8236), .B(n8235), .ZN(n8237)
         );
  OAI21_X1 U9954 ( .B1(n8238), .B2(n8345), .A(n8237), .ZN(P2_U3160) );
  XOR2_X1 U9955 ( .A(n8239), .B(n8240), .Z(n8246) );
  AOI22_X1 U9956 ( .A1(n8833), .A2(n8348), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8242) );
  NAND2_X1 U9957 ( .A1(n8836), .A2(n8352), .ZN(n8241) );
  OAI211_X1 U9958 ( .C1(n8243), .C2(n8350), .A(n8242), .B(n8241), .ZN(n8244)
         );
  AOI21_X1 U9959 ( .B1(n9054), .B2(n8341), .A(n8244), .ZN(n8245) );
  OAI21_X1 U9960 ( .B1(n8246), .B2(n8345), .A(n8245), .ZN(P2_U3163) );
  XOR2_X1 U9961 ( .A(n8248), .B(n8247), .Z(n8253) );
  NAND2_X1 U9962 ( .A1(n8767), .A2(n8336), .ZN(n8250) );
  AOI22_X1 U9963 ( .A1(n8785), .A2(n8352), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8249) );
  OAI211_X1 U9964 ( .C1(n8783), .C2(n8339), .A(n8250), .B(n8249), .ZN(n8251)
         );
  AOI21_X1 U9965 ( .B1(n9030), .B2(n8341), .A(n8251), .ZN(n8252) );
  OAI21_X1 U9966 ( .B1(n8253), .B2(n8345), .A(n8252), .ZN(P2_U3165) );
  XNOR2_X1 U9967 ( .A(n8254), .B(n8924), .ZN(n8259) );
  XNOR2_X1 U9968 ( .A(n8256), .B(n8936), .ZN(n8346) );
  NOR2_X1 U9969 ( .A1(n8255), .A2(n8346), .ZN(n8344) );
  OR2_X1 U9970 ( .A1(n8344), .A2(n8257), .ZN(n8258) );
  NOR2_X1 U9971 ( .A1(n8258), .A2(n8259), .ZN(n8265) );
  AOI21_X1 U9972 ( .B1(n8259), .B2(n8258), .A(n8265), .ZN(n8264) );
  NAND2_X1 U9973 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8707) );
  NAND2_X1 U9974 ( .A1(n8348), .A2(n8936), .ZN(n8260) );
  OAI211_X1 U9975 ( .C1(n8911), .C2(n8350), .A(n8707), .B(n8260), .ZN(n8261)
         );
  AOI21_X1 U9976 ( .B1(n8917), .B2(n8352), .A(n8261), .ZN(n8263) );
  NAND2_X1 U9977 ( .A1(n8986), .A2(n8341), .ZN(n8262) );
  OAI211_X1 U9978 ( .C1(n8264), .C2(n8345), .A(n8263), .B(n8262), .ZN(P2_U3166) );
  INV_X1 U9979 ( .A(n9073), .ZN(n8275) );
  AOI211_X1 U9980 ( .C1(n8892), .C2(n8267), .A(n8266), .B(n8265), .ZN(n8270)
         );
  INV_X1 U9981 ( .A(n8268), .ZN(n8269) );
  OAI21_X1 U9982 ( .B1(n8270), .B2(n8269), .A(n6606), .ZN(n8274) );
  NAND2_X1 U9983 ( .A1(n8924), .A2(n8348), .ZN(n8271) );
  NAND2_X1 U9984 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8726) );
  OAI211_X1 U9985 ( .C1(n8893), .C2(n8350), .A(n8271), .B(n8726), .ZN(n8272)
         );
  AOI21_X1 U9986 ( .B1(n8898), .B2(n8352), .A(n8272), .ZN(n8273) );
  OAI211_X1 U9987 ( .C1(n8275), .C2(n8355), .A(n8274), .B(n8273), .ZN(P2_U3168) );
  XNOR2_X1 U9988 ( .A(n8279), .B(n8783), .ZN(n8280) );
  NAND2_X1 U9989 ( .A1(n4568), .A2(n8336), .ZN(n8282) );
  AOI22_X1 U9990 ( .A1(n8798), .A2(n8352), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8281) );
  OAI211_X1 U9991 ( .C1(n8321), .C2(n8339), .A(n8282), .B(n8281), .ZN(n8283)
         );
  AOI21_X1 U9992 ( .B1(n9036), .B2(n8341), .A(n8283), .ZN(n8284) );
  OAI21_X1 U9993 ( .B1(n8287), .B2(n8286), .A(n8285), .ZN(n8288) );
  NAND2_X1 U9994 ( .A1(n8288), .A2(n6606), .ZN(n8296) );
  AOI22_X1 U9995 ( .A1(n8336), .A2(n8625), .B1(n8341), .B2(n8289), .ZN(n8295)
         );
  INV_X1 U9996 ( .A(n8290), .ZN(n8291) );
  AOI21_X1 U9997 ( .B1(n8348), .B2(n10260), .A(n8291), .ZN(n8294) );
  NAND2_X1 U9998 ( .A1(n8352), .A2(n8292), .ZN(n8293) );
  NAND4_X1 U9999 ( .A1(n8296), .A2(n8295), .A3(n8294), .A4(n8293), .ZN(
        P2_U3170) );
  AOI21_X1 U10000 ( .B1(n8298), .B2(n8297), .A(n4371), .ZN(n8304) );
  AOI22_X1 U10001 ( .A1(n8847), .A2(n8348), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8300) );
  NAND2_X1 U10002 ( .A1(n8850), .A2(n8352), .ZN(n8299) );
  OAI211_X1 U10003 ( .C1(n8301), .C2(n8350), .A(n8300), .B(n8299), .ZN(n8302)
         );
  AOI21_X1 U10004 ( .B1(n9060), .B2(n8341), .A(n8302), .ZN(n8303) );
  OAI21_X1 U10005 ( .B1(n8304), .B2(n8345), .A(n8303), .ZN(P2_U3173) );
  INV_X1 U10006 ( .A(n8305), .ZN(n8306) );
  AOI21_X1 U10007 ( .B1(n8308), .B2(n8307), .A(n8306), .ZN(n8316) );
  NAND2_X1 U10008 ( .A1(n8336), .A2(n8925), .ZN(n8309) );
  NAND2_X1 U10009 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8653) );
  OAI211_X1 U10010 ( .C1(n8310), .C2(n8339), .A(n8309), .B(n8653), .ZN(n8313)
         );
  NOR2_X1 U10011 ( .A1(n8311), .A2(n8355), .ZN(n8312) );
  AOI211_X1 U10012 ( .C1(n8314), .C2(n8352), .A(n8313), .B(n8312), .ZN(n8315)
         );
  OAI21_X1 U10013 ( .B1(n8316), .B2(n8345), .A(n8315), .ZN(P2_U3174) );
  XOR2_X1 U10014 ( .A(n8318), .B(n8317), .Z(n8324) );
  AOI22_X1 U10015 ( .A1(n8846), .A2(n8348), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8320) );
  NAND2_X1 U10016 ( .A1(n8822), .A2(n8352), .ZN(n8319) );
  OAI211_X1 U10017 ( .C1(n8321), .C2(n8350), .A(n8320), .B(n8319), .ZN(n8322)
         );
  AOI21_X1 U10018 ( .B1(n9048), .B2(n8341), .A(n8322), .ZN(n8323) );
  OAI21_X1 U10019 ( .B1(n8324), .B2(n8345), .A(n8323), .ZN(P2_U3175) );
  XOR2_X1 U10020 ( .A(n8326), .B(n8325), .Z(n8333) );
  NAND2_X1 U10021 ( .A1(n8327), .A2(n8348), .ZN(n8329) );
  OAI211_X1 U10022 ( .C1(n8873), .C2(n8350), .A(n8329), .B(n8328), .ZN(n8331)
         );
  NOR2_X1 U10023 ( .A1(n8881), .A2(n8355), .ZN(n8330) );
  AOI211_X1 U10024 ( .C1(n8878), .C2(n8352), .A(n8331), .B(n8330), .ZN(n8332)
         );
  OAI21_X1 U10025 ( .B1(n8333), .B2(n8345), .A(n8332), .ZN(P2_U3178) );
  XOR2_X1 U10026 ( .A(n8335), .B(n8334), .Z(n8343) );
  NAND2_X1 U10027 ( .A1(n8775), .A2(n8336), .ZN(n8338) );
  AOI22_X1 U10028 ( .A1(n8776), .A2(n8352), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8337) );
  OAI211_X1 U10029 ( .C1(n8423), .C2(n8339), .A(n8338), .B(n8337), .ZN(n8340)
         );
  AOI21_X1 U10030 ( .B1(n9024), .B2(n8341), .A(n8340), .ZN(n8342) );
  OAI21_X1 U10031 ( .B1(n8343), .B2(n8345), .A(n8342), .ZN(P2_U3180) );
  INV_X1 U10032 ( .A(n9085), .ZN(n8356) );
  AOI211_X1 U10033 ( .C1(n8346), .C2(n8255), .A(n8345), .B(n8344), .ZN(n8347)
         );
  INV_X1 U10034 ( .A(n8347), .ZN(n8354) );
  NAND2_X1 U10035 ( .A1(n8348), .A2(n8925), .ZN(n8349) );
  NAND2_X1 U10036 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8692) );
  OAI211_X1 U10037 ( .C1(n8892), .C2(n8350), .A(n8349), .B(n8692), .ZN(n8351)
         );
  AOI21_X1 U10038 ( .B1(n8928), .B2(n8352), .A(n8351), .ZN(n8353) );
  OAI211_X1 U10039 ( .C1(n8356), .C2(n8355), .A(n8354), .B(n8353), .ZN(
        P2_U3181) );
  INV_X1 U10040 ( .A(n8586), .ZN(n8377) );
  NAND2_X1 U10041 ( .A1(n7910), .A2(n8563), .ZN(n8359) );
  OR2_X1 U10042 ( .A1(n8363), .A2(n8357), .ZN(n8358) );
  INV_X1 U10043 ( .A(n8619), .ZN(n8379) );
  NAND2_X1 U10044 ( .A1(n8949), .A2(n8379), .ZN(n8592) );
  NAND2_X1 U10045 ( .A1(n8592), .A2(n8360), .ZN(n8421) );
  OR2_X1 U10046 ( .A1(n8361), .A2(n8565), .ZN(n8365) );
  INV_X1 U10047 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8362) );
  OR2_X1 U10048 ( .A1(n8363), .A2(n8362), .ZN(n8364) );
  NAND2_X1 U10049 ( .A1(n9012), .A2(n8949), .ZN(n8374) );
  INV_X1 U10050 ( .A(n9012), .ZN(n8414) );
  NAND2_X1 U10051 ( .A1(n8366), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8371) );
  NAND2_X1 U10052 ( .A1(n4311), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8370) );
  NAND2_X1 U10053 ( .A1(n8368), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8369) );
  AND3_X1 U10054 ( .A1(n8371), .A2(n8370), .A3(n8369), .ZN(n8372) );
  NAND2_X1 U10055 ( .A1(n8374), .A2(n8598), .ZN(n8375) );
  NOR2_X1 U10056 ( .A1(n8421), .A2(n8375), .ZN(n8376) );
  OAI21_X1 U10057 ( .B1(n8378), .B2(n8377), .A(n8376), .ZN(n8382) );
  AOI21_X1 U10058 ( .B1(n8594), .B2(n8758), .A(n9012), .ZN(n8380) );
  NOR2_X1 U10059 ( .A1(n8380), .A2(n8445), .ZN(n8381) );
  NAND2_X1 U10060 ( .A1(n8382), .A2(n8381), .ZN(n8419) );
  INV_X1 U10061 ( .A(n8383), .ZN(n8557) );
  INV_X1 U10062 ( .A(n8794), .ZN(n8408) );
  INV_X1 U10063 ( .A(n8790), .ZN(n8384) );
  NAND3_X1 U10064 ( .A1(n8386), .A2(n8385), .A3(n7034), .ZN(n8390) );
  NAND3_X1 U10065 ( .A1(n8388), .A2(n8387), .A3(n8457), .ZN(n8389) );
  NOR2_X1 U10066 ( .A1(n8390), .A2(n8389), .ZN(n8394) );
  NAND4_X1 U10067 ( .A1(n8394), .A2(n8393), .A3(n8392), .A4(n8391), .ZN(n8395)
         );
  NOR3_X1 U10068 ( .A1(n8397), .A2(n8396), .A3(n8395), .ZN(n8398) );
  NAND4_X1 U10069 ( .A1(n8513), .A2(n8509), .A3(n8399), .A4(n8398), .ZN(n8400)
         );
  NAND2_X1 U10070 ( .A1(n8431), .A2(n8432), .ZN(n8935) );
  NOR2_X1 U10071 ( .A1(n8400), .A2(n8935), .ZN(n8402) );
  INV_X1 U10072 ( .A(n8901), .ZN(n8401) );
  NAND2_X1 U10073 ( .A1(n8401), .A2(n8903), .ZN(n8922) );
  NAND3_X1 U10074 ( .A1(n8915), .A2(n8402), .A3(n8922), .ZN(n8403) );
  NAND2_X1 U10075 ( .A1(n8859), .A2(n8404), .ZN(n8405) );
  OR4_X1 U10076 ( .A1(n8813), .A2(n8844), .A3(n8828), .A4(n8405), .ZN(n8406)
         );
  NOR2_X1 U10077 ( .A1(n8804), .A2(n8406), .ZN(n8407) );
  NAND2_X1 U10078 ( .A1(n8408), .A2(n8407), .ZN(n8409) );
  NOR2_X1 U10079 ( .A1(n8409), .A2(n8786), .ZN(n8410) );
  NAND4_X1 U10080 ( .A1(n8586), .A2(n8764), .A3(n8774), .A4(n8410), .ZN(n8411)
         );
  NOR2_X1 U10081 ( .A1(n8412), .A2(n8411), .ZN(n8415) );
  NAND2_X1 U10082 ( .A1(n8414), .A2(n8413), .ZN(n8593) );
  NAND4_X1 U10083 ( .A1(n8594), .A2(n8415), .A3(n8593), .A4(n8598), .ZN(n8416)
         );
  NOR2_X1 U10084 ( .A1(n8416), .A2(n8421), .ZN(n8417) );
  NAND2_X1 U10085 ( .A1(n8419), .A2(n8418), .ZN(n8611) );
  INV_X1 U10086 ( .A(n8609), .ZN(n8420) );
  NAND2_X1 U10087 ( .A1(n8739), .A2(n8420), .ZN(n8602) );
  OR3_X1 U10088 ( .A1(n8611), .A2(n8613), .A3(n8602), .ZN(n8618) );
  INV_X1 U10089 ( .A(n8421), .ZN(n8585) );
  NAND2_X1 U10090 ( .A1(n8422), .A2(n8584), .ZN(n8549) );
  OR3_X1 U10091 ( .A1(n9030), .A2(n8591), .A3(n8423), .ZN(n8424) );
  OAI211_X1 U10092 ( .C1(n8426), .C2(n8584), .A(n8425), .B(n8424), .ZN(n8427)
         );
  INV_X1 U10093 ( .A(n8786), .ZN(n8780) );
  INV_X1 U10094 ( .A(n8428), .ZN(n8429) );
  OAI21_X1 U10095 ( .B1(n8430), .B2(n8429), .A(n8591), .ZN(n8548) );
  INV_X1 U10096 ( .A(n8521), .ZN(n8525) );
  NAND2_X1 U10097 ( .A1(n8516), .A2(n8431), .ZN(n8434) );
  INV_X1 U10098 ( .A(n8432), .ZN(n8433) );
  MUX2_X1 U10099 ( .A(n8434), .B(n8433), .S(n8591), .Z(n8435) );
  INV_X1 U10100 ( .A(n8435), .ZN(n8515) );
  AND2_X1 U10101 ( .A1(n8436), .A2(n8591), .ZN(n8438) );
  NOR2_X1 U10102 ( .A1(n8436), .A2(n8591), .ZN(n8437) );
  MUX2_X1 U10103 ( .A(n8438), .B(n8437), .S(n8937), .Z(n8439) );
  NAND2_X1 U10104 ( .A1(n8442), .A2(n8440), .ZN(n8441) );
  NAND2_X1 U10105 ( .A1(n8441), .A2(n8584), .ZN(n8444) );
  NAND3_X1 U10106 ( .A1(n8447), .A2(n8442), .A3(n8603), .ZN(n8443) );
  NOR2_X1 U10107 ( .A1(n8447), .A2(n8591), .ZN(n8448) );
  NOR2_X1 U10108 ( .A1(n8448), .A2(n10255), .ZN(n8449) );
  NAND2_X1 U10109 ( .A1(n8491), .A2(n8450), .ZN(n8453) );
  NAND2_X1 U10110 ( .A1(n8459), .A2(n8451), .ZN(n8452) );
  MUX2_X1 U10111 ( .A(n8453), .B(n8452), .S(n8591), .Z(n8454) );
  INV_X1 U10112 ( .A(n8454), .ZN(n8455) );
  NAND2_X1 U10113 ( .A1(n8456), .A2(n8455), .ZN(n8458) );
  NAND2_X1 U10114 ( .A1(n8458), .A2(n8457), .ZN(n8496) );
  INV_X1 U10115 ( .A(n8459), .ZN(n8463) );
  INV_X1 U10116 ( .A(n8460), .ZN(n8462) );
  OAI211_X1 U10117 ( .C1(n8496), .C2(n8463), .A(n8462), .B(n8461), .ZN(n8468)
         );
  NAND2_X1 U10118 ( .A1(n8465), .A2(n8464), .ZN(n8492) );
  NAND2_X1 U10119 ( .A1(n8492), .A2(n8466), .ZN(n8467) );
  AOI21_X1 U10120 ( .B1(n8468), .B2(n8467), .A(n8497), .ZN(n8475) );
  NAND2_X1 U10121 ( .A1(n8470), .A2(n8469), .ZN(n8474) );
  NAND2_X1 U10122 ( .A1(n8477), .A2(n8470), .ZN(n8472) );
  NAND2_X1 U10123 ( .A1(n8503), .A2(n8500), .ZN(n8471) );
  MUX2_X1 U10124 ( .A(n8472), .B(n8471), .S(n8584), .Z(n8473) );
  INV_X1 U10125 ( .A(n8473), .ZN(n8507) );
  OAI21_X1 U10126 ( .B1(n8475), .B2(n8474), .A(n8507), .ZN(n8479) );
  NOR2_X1 U10127 ( .A1(n8476), .A2(n8591), .ZN(n8478) );
  NAND4_X1 U10128 ( .A1(n8479), .A2(n8478), .A3(n8483), .A4(n8477), .ZN(n8490)
         );
  NAND4_X1 U10129 ( .A1(n8505), .A2(n8591), .A3(n8480), .A4(n8623), .ZN(n8489)
         );
  NAND4_X1 U10130 ( .A1(n8483), .A2(n8482), .A3(n8584), .A4(n8481), .ZN(n8488)
         );
  NOR2_X1 U10131 ( .A1(n8484), .A2(n8584), .ZN(n8486) );
  OAI21_X1 U10132 ( .B1(n8591), .B2(n8622), .A(n8997), .ZN(n8485) );
  OAI21_X1 U10133 ( .B1(n8486), .B2(n8997), .A(n8485), .ZN(n8487) );
  INV_X1 U10134 ( .A(n8491), .ZN(n8495) );
  INV_X1 U10135 ( .A(n8492), .ZN(n8494) );
  NAND2_X1 U10136 ( .A1(n10290), .A2(n8626), .ZN(n8493) );
  OAI211_X1 U10137 ( .C1(n8496), .C2(n8495), .A(n8494), .B(n8493), .ZN(n8499)
         );
  AOI21_X1 U10138 ( .B1(n8499), .B2(n8498), .A(n8497), .ZN(n8502) );
  NAND4_X1 U10139 ( .A1(n8505), .A2(n8591), .A3(n8504), .A4(n8503), .ZN(n8506)
         );
  MUX2_X1 U10140 ( .A(n8511), .B(n8510), .S(n8584), .Z(n8512) );
  INV_X1 U10141 ( .A(n8935), .ZN(n8944) );
  OAI211_X1 U10142 ( .C1(n8527), .C2(n8526), .A(n8528), .B(n8516), .ZN(n8517)
         );
  NAND2_X1 U10143 ( .A1(n8521), .A2(n8520), .ZN(n8522) );
  NAND2_X1 U10144 ( .A1(n8522), .A2(n8591), .ZN(n8523) );
  NAND3_X1 U10145 ( .A1(n8531), .A2(n8536), .A3(n8532), .ZN(n8524) );
  NAND2_X1 U10146 ( .A1(n8527), .A2(n4896), .ZN(n8529) );
  NAND3_X1 U10147 ( .A1(n8529), .A2(n8584), .A3(n8528), .ZN(n8530) );
  NAND2_X1 U10148 ( .A1(n8531), .A2(n8530), .ZN(n8533) );
  OAI211_X1 U10149 ( .C1(n8911), .C2(n9073), .A(n8533), .B(n8532), .ZN(n8534)
         );
  AND2_X1 U10150 ( .A1(n8825), .A2(n8535), .ZN(n8539) );
  INV_X1 U10151 ( .A(n8536), .ZN(n8537) );
  NOR2_X1 U10152 ( .A1(n8844), .A2(n8537), .ZN(n8538) );
  MUX2_X1 U10153 ( .A(n8539), .B(n8538), .S(n8584), .Z(n8540) );
  OR2_X1 U10154 ( .A1(n8541), .A2(n8591), .ZN(n8542) );
  AOI21_X1 U10155 ( .B1(n8544), .B2(n8543), .A(n8584), .ZN(n8547) );
  NOR2_X1 U10156 ( .A1(n8545), .A2(n8584), .ZN(n8546) );
  INV_X1 U10157 ( .A(n8549), .ZN(n8551) );
  NAND4_X1 U10158 ( .A1(n8780), .A2(n8552), .A3(n8551), .A4(n8550), .ZN(n8556)
         );
  MUX2_X1 U10159 ( .A(n8558), .B(n8557), .S(n8584), .Z(n8559) );
  NAND3_X1 U10160 ( .A1(n8560), .A2(n8764), .A3(n8559), .ZN(n8575) );
  MUX2_X1 U10161 ( .A(n8562), .B(n8561), .S(n8584), .Z(n8573) );
  NAND2_X1 U10162 ( .A1(n8569), .A2(n8563), .ZN(n8564) );
  OR2_X1 U10163 ( .A1(n10000), .A2(n8564), .ZN(n8572) );
  INV_X1 U10164 ( .A(n8569), .ZN(n8620) );
  NAND3_X1 U10165 ( .A1(n10000), .A2(n8620), .A3(n8566), .ZN(n8571) );
  AND2_X1 U10166 ( .A1(n8566), .A2(n8565), .ZN(n8568) );
  NAND2_X1 U10167 ( .A1(n8569), .A2(n8566), .ZN(n8567) );
  OAI21_X1 U10168 ( .B1(n8569), .B2(n8568), .A(n8567), .ZN(n8570) );
  AND3_X1 U10169 ( .A1(n8572), .A2(n8571), .A3(n8570), .ZN(n8578) );
  AND2_X1 U10170 ( .A1(n8573), .A2(n8578), .ZN(n8574) );
  NAND2_X1 U10171 ( .A1(n8575), .A2(n8574), .ZN(n8581) );
  MUX2_X1 U10172 ( .A(n8766), .B(n8576), .S(n8584), .Z(n8579) );
  INV_X1 U10173 ( .A(n8579), .ZN(n8577) );
  NAND2_X1 U10174 ( .A1(n8579), .A2(n8578), .ZN(n8580) );
  NAND2_X1 U10175 ( .A1(n8581), .A2(n8580), .ZN(n8588) );
  NAND2_X1 U10176 ( .A1(n8588), .A2(n8582), .ZN(n8583) );
  NAND4_X1 U10177 ( .A1(n8585), .A2(n8584), .A3(n8589), .A4(n8583), .ZN(n8601)
         );
  AND2_X1 U10178 ( .A1(n8593), .A2(n8586), .ZN(n8590) );
  NAND2_X1 U10179 ( .A1(n8592), .A2(n8591), .ZN(n8595) );
  NAND3_X1 U10180 ( .A1(n8595), .A2(n8594), .A3(n8593), .ZN(n8596) );
  NAND2_X1 U10181 ( .A1(n8597), .A2(n8596), .ZN(n8600) );
  INV_X1 U10182 ( .A(n8598), .ZN(n8599) );
  NOR2_X1 U10183 ( .A1(n8602), .A2(n8610), .ZN(n8608) );
  NOR2_X1 U10184 ( .A1(n6498), .A2(n8744), .ZN(n8605) );
  OAI21_X1 U10185 ( .B1(n8609), .B2(n8603), .A(P2_B_REG_SCAN_IN), .ZN(n8604)
         );
  AOI21_X1 U10186 ( .B1(n8606), .B2(n8605), .A(n8604), .ZN(n8607) );
  AOI21_X1 U10187 ( .B1(n8612), .B2(n8608), .A(n8607), .ZN(n8617) );
  NOR2_X1 U10188 ( .A1(n8739), .A2(n8609), .ZN(n8614) );
  NAND3_X1 U10189 ( .A1(n8611), .A2(n8610), .A3(n8614), .ZN(n8616) );
  NAND4_X1 U10190 ( .A1(n8618), .A2(n8617), .A3(n8616), .A4(n8615), .ZN(
        P2_U3296) );
  MUX2_X1 U10191 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8758), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10192 ( .A(n8619), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8628), .Z(
        P2_U3521) );
  MUX2_X1 U10193 ( .A(n8620), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8628), .Z(
        P2_U3520) );
  MUX2_X1 U10194 ( .A(n8766), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8628), .Z(
        P2_U3519) );
  MUX2_X1 U10195 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8775), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10196 ( .A(n8767), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8628), .Z(
        P2_U3517) );
  MUX2_X1 U10197 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n4568), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10198 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8805), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10199 ( .A(n8819), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8628), .Z(
        P2_U3514) );
  MUX2_X1 U10200 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8832), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10201 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8846), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10202 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8833), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10203 ( .A(n8924), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8628), .Z(
        P2_U3507) );
  MUX2_X1 U10204 ( .A(n8936), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8628), .Z(
        P2_U3506) );
  MUX2_X1 U10205 ( .A(n8925), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8628), .Z(
        P2_U3505) );
  MUX2_X1 U10206 ( .A(n8937), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8628), .Z(
        P2_U3504) );
  MUX2_X1 U10207 ( .A(n8621), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8628), .Z(
        P2_U3503) );
  MUX2_X1 U10208 ( .A(n8622), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8628), .Z(
        P2_U3502) );
  MUX2_X1 U10209 ( .A(n8623), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8628), .Z(
        P2_U3501) );
  MUX2_X1 U10210 ( .A(n8624), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8628), .Z(
        P2_U3498) );
  MUX2_X1 U10211 ( .A(n8625), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8628), .Z(
        P2_U3496) );
  MUX2_X1 U10212 ( .A(n8626), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8628), .Z(
        P2_U3495) );
  MUX2_X1 U10213 ( .A(n10260), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8628), .Z(
        P2_U3494) );
  MUX2_X1 U10214 ( .A(n8627), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8628), .Z(
        P2_U3493) );
  MUX2_X1 U10215 ( .A(n6168), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8628), .Z(
        P2_U3492) );
  MUX2_X1 U10216 ( .A(n6695), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8628), .Z(
        P2_U3491) );
  OAI21_X1 U10217 ( .B1(n8631), .B2(n8630), .A(n8629), .ZN(n8632) );
  NAND2_X1 U10218 ( .A1(n8632), .A2(n8753), .ZN(n8650) );
  INV_X1 U10219 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n8634) );
  OAI21_X1 U10220 ( .B1(n8654), .B2(n8634), .A(n8633), .ZN(n8635) );
  AOI21_X1 U10221 ( .B1(n8636), .B2(n8663), .A(n8635), .ZN(n8649) );
  AND3_X1 U10222 ( .A1(n6741), .A2(n8638), .A3(n8637), .ZN(n8640) );
  OAI21_X1 U10223 ( .B1(n8641), .B2(n8640), .A(n8639), .ZN(n8648) );
  AND3_X1 U10224 ( .A1(n8642), .A2(n8643), .A3(n8644), .ZN(n8645) );
  OAI21_X1 U10225 ( .B1(n8646), .B2(n8645), .A(n8740), .ZN(n8647) );
  NAND4_X1 U10226 ( .A1(n8650), .A2(n8649), .A3(n8648), .A4(n8647), .ZN(
        P2_U3188) );
  AOI21_X1 U10227 ( .B1(n8652), .B2(n8651), .A(n8676), .ZN(n8667) );
  INV_X1 U10228 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n9856) );
  OAI21_X1 U10229 ( .B1(n8654), .B2(n9856), .A(n8653), .ZN(n8661) );
  NAND2_X1 U10230 ( .A1(n8656), .A2(n8655), .ZN(n8658) );
  AOI21_X1 U10231 ( .B1(n8659), .B2(n8658), .A(n8657), .ZN(n8660) );
  AOI211_X1 U10232 ( .C1(n8663), .C2(n8662), .A(n8661), .B(n8660), .ZN(n8666)
         );
  NOR2_X1 U10233 ( .A1(n4396), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8664) );
  OAI21_X1 U10234 ( .B1(n8664), .B2(n8684), .A(n8740), .ZN(n8665) );
  OAI211_X1 U10235 ( .C1(n8667), .C2(n8756), .A(n8666), .B(n8665), .ZN(
        P2_U3195) );
  OAI21_X1 U10236 ( .B1(n8670), .B2(n8669), .A(n8668), .ZN(n8681) );
  NAND2_X1 U10237 ( .A1(n8748), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n8671) );
  OAI211_X1 U10238 ( .C1(n8751), .C2(n8673), .A(n8672), .B(n8671), .ZN(n8680)
         );
  OR3_X1 U10239 ( .A1(n8676), .A2(n8675), .A3(n8674), .ZN(n8677) );
  AOI21_X1 U10240 ( .B1(n8678), .B2(n8677), .A(n8756), .ZN(n8679) );
  AOI211_X1 U10241 ( .C1(n8753), .C2(n8681), .A(n8680), .B(n8679), .ZN(n8687)
         );
  NOR3_X1 U10242 ( .A1(n8684), .A2(n8683), .A3(n8682), .ZN(n8685) );
  OAI21_X1 U10243 ( .B1(n4400), .B2(n8685), .A(n8740), .ZN(n8686) );
  NAND2_X1 U10244 ( .A1(n8687), .A2(n8686), .ZN(P2_U3196) );
  AOI21_X1 U10245 ( .B1(n8989), .B2(n8688), .A(n4322), .ZN(n8700) );
  XNOR2_X1 U10246 ( .A(n8690), .B(n8689), .ZN(n8698) );
  NAND2_X1 U10247 ( .A1(n8748), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n8691) );
  OAI211_X1 U10248 ( .C1(n8751), .C2(n8693), .A(n8692), .B(n8691), .ZN(n8697)
         );
  AOI21_X1 U10249 ( .B1(n8927), .B2(n8694), .A(n8711), .ZN(n8695) );
  NOR2_X1 U10250 ( .A1(n8695), .A2(n8712), .ZN(n8696) );
  AOI211_X1 U10251 ( .C1(n8753), .C2(n8698), .A(n8697), .B(n8696), .ZN(n8699)
         );
  OAI21_X1 U10252 ( .B1(n8700), .B2(n8756), .A(n8699), .ZN(P2_U3197) );
  NOR3_X1 U10253 ( .A1(n4322), .A2(n8702), .A3(n8701), .ZN(n8703) );
  NOR2_X1 U10254 ( .A1(n4359), .A2(n8703), .ZN(n8719) );
  XNOR2_X1 U10255 ( .A(n8705), .B(n8704), .ZN(n8717) );
  NAND2_X1 U10256 ( .A1(n8748), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8706) );
  OAI211_X1 U10257 ( .C1(n8751), .C2(n8708), .A(n8707), .B(n8706), .ZN(n8716)
         );
  OR3_X1 U10258 ( .A1(n8711), .A2(n8710), .A3(n8709), .ZN(n8713) );
  AOI21_X1 U10259 ( .B1(n8714), .B2(n8713), .A(n8712), .ZN(n8715) );
  AOI211_X1 U10260 ( .C1(n8753), .C2(n8717), .A(n8716), .B(n8715), .ZN(n8718)
         );
  OAI21_X1 U10261 ( .B1(n8719), .B2(n8756), .A(n8718), .ZN(P2_U3198) );
  INV_X1 U10262 ( .A(n8720), .ZN(n8721) );
  AOI21_X1 U10263 ( .B1(n8983), .B2(n8722), .A(n8721), .ZN(n8734) );
  XNOR2_X1 U10264 ( .A(n8724), .B(n8723), .ZN(n8729) );
  NAND2_X1 U10265 ( .A1(n8748), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n8725) );
  OAI211_X1 U10266 ( .C1(n8751), .C2(n8727), .A(n8726), .B(n8725), .ZN(n8728)
         );
  AOI21_X1 U10267 ( .B1(n8729), .B2(n8753), .A(n8728), .ZN(n8733) );
  OAI21_X1 U10268 ( .B1(n4364), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8730), .ZN(
        n8731) );
  NAND2_X1 U10269 ( .A1(n8731), .A2(n8740), .ZN(n8732) );
  OAI211_X1 U10270 ( .C1(n8734), .C2(n8756), .A(n8733), .B(n8732), .ZN(
        P2_U3199) );
  XNOR2_X1 U10271 ( .A(n8739), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8745) );
  MUX2_X1 U10272 ( .A(n4408), .B(n8745), .S(n8744), .Z(n8746) );
  XNOR2_X1 U10273 ( .A(n8747), .B(n8746), .ZN(n8754) );
  NAND2_X1 U10274 ( .A1(n8748), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8749) );
  OAI211_X1 U10275 ( .C1(n8751), .C2(n6194), .A(n8750), .B(n8749), .ZN(n8752)
         );
  AOI21_X1 U10276 ( .B1(n8754), .B2(n8753), .A(n8752), .ZN(n8755) );
  AOI21_X1 U10277 ( .B1(n9010), .B2(n10269), .A(n8759), .ZN(n8762) );
  NAND2_X1 U10278 ( .A1(n10272), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8760) );
  OAI211_X1 U10279 ( .C1(n9012), .C2(n8880), .A(n8762), .B(n8760), .ZN(
        P2_U3202) );
  INV_X1 U10280 ( .A(n8949), .ZN(n9015) );
  NAND2_X1 U10281 ( .A1(n10272), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8761) );
  OAI211_X1 U10282 ( .C1(n9015), .C2(n8880), .A(n8762), .B(n8761), .ZN(
        P2_U3203) );
  XNOR2_X1 U10283 ( .A(n8763), .B(n8764), .ZN(n9021) );
  INV_X1 U10284 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8768) );
  MUX2_X1 U10285 ( .A(n8768), .B(n9016), .S(n10269), .Z(n8771) );
  AOI22_X1 U10286 ( .A1(n9018), .A2(n8929), .B1(n8942), .B2(n8769), .ZN(n8770)
         );
  OAI211_X1 U10287 ( .C1(n9021), .C2(n8932), .A(n8771), .B(n8770), .ZN(
        P2_U3206) );
  XOR2_X1 U10288 ( .A(n8772), .B(n8774), .Z(n9027) );
  MUX2_X1 U10289 ( .A(n9904), .B(n9022), .S(n10269), .Z(n8778) );
  AOI22_X1 U10290 ( .A1(n9024), .A2(n8929), .B1(n8942), .B2(n8776), .ZN(n8777)
         );
  OAI211_X1 U10291 ( .C1(n9027), .C2(n8932), .A(n8778), .B(n8777), .ZN(
        P2_U3207) );
  NOR2_X1 U10292 ( .A1(n4567), .A2(n10251), .ZN(n8784) );
  XNOR2_X1 U10293 ( .A(n8779), .B(n8780), .ZN(n8781) );
  OAI222_X1 U10294 ( .A1(n8908), .A2(n8783), .B1(n8910), .B2(n8782), .C1(n8871), .C2(n8781), .ZN(n8957) );
  AOI211_X1 U10295 ( .C1(n8942), .C2(n8785), .A(n8784), .B(n8957), .ZN(n8789)
         );
  XNOR2_X1 U10296 ( .A(n8787), .B(n8786), .ZN(n9031) );
  AOI22_X1 U10297 ( .A1(n9031), .A2(n8945), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n10272), .ZN(n8788) );
  OAI21_X1 U10298 ( .B1(n8789), .B2(n10272), .A(n8788), .ZN(P2_U3208) );
  NAND2_X1 U10299 ( .A1(n8791), .A2(n8790), .ZN(n8792) );
  XNOR2_X1 U10300 ( .A(n8792), .B(n8794), .ZN(n9039) );
  INV_X1 U10301 ( .A(n9036), .ZN(n8796) );
  XNOR2_X1 U10302 ( .A(n8793), .B(n8794), .ZN(n8795) );
  AOI222_X1 U10303 ( .A1(n10257), .A2(n8795), .B1(n8819), .B2(n10262), .C1(
        n4568), .C2(n10261), .ZN(n9034) );
  OAI21_X1 U10304 ( .B1(n8796), .B2(n10251), .A(n9034), .ZN(n8797) );
  NAND2_X1 U10305 ( .A1(n8797), .A2(n10269), .ZN(n8800) );
  AOI22_X1 U10306 ( .A1(n8798), .A2(n8942), .B1(n10272), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8799) );
  OAI211_X1 U10307 ( .C1(n9039), .C2(n8932), .A(n8800), .B(n8799), .ZN(
        P2_U3209) );
  XNOR2_X1 U10308 ( .A(n8801), .B(n8804), .ZN(n9043) );
  INV_X1 U10309 ( .A(n9043), .ZN(n8811) );
  INV_X1 U10310 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8807) );
  XNOR2_X1 U10311 ( .A(n8803), .B(n8804), .ZN(n8806) );
  AOI222_X1 U10312 ( .A1(n10257), .A2(n8806), .B1(n8832), .B2(n10262), .C1(
        n8805), .C2(n10261), .ZN(n9040) );
  MUX2_X1 U10313 ( .A(n8807), .B(n9040), .S(n10269), .Z(n8810) );
  AOI22_X1 U10314 ( .A1(n9042), .A2(n8929), .B1(n8942), .B2(n8808), .ZN(n8809)
         );
  OAI211_X1 U10315 ( .C1(n8811), .C2(n8932), .A(n8810), .B(n8809), .ZN(
        P2_U3210) );
  XOR2_X1 U10316 ( .A(n8812), .B(n8813), .Z(n9051) );
  INV_X1 U10317 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8821) );
  INV_X1 U10318 ( .A(n8844), .ZN(n8839) );
  OAI21_X1 U10319 ( .B1(n8842), .B2(n8829), .A(n8828), .ZN(n8831) );
  INV_X1 U10320 ( .A(n8813), .ZN(n8816) );
  INV_X1 U10321 ( .A(n8814), .ZN(n8815) );
  NAND3_X1 U10322 ( .A1(n8831), .A2(n8816), .A3(n8815), .ZN(n8818) );
  NAND2_X1 U10323 ( .A1(n8818), .A2(n8817), .ZN(n8820) );
  AOI222_X1 U10324 ( .A1(n10257), .A2(n8820), .B1(n8846), .B2(n10262), .C1(
        n8819), .C2(n10261), .ZN(n9046) );
  MUX2_X1 U10325 ( .A(n8821), .B(n9046), .S(n10269), .Z(n8824) );
  AOI22_X1 U10326 ( .A1(n9048), .A2(n8929), .B1(n8942), .B2(n8822), .ZN(n8823)
         );
  OAI211_X1 U10327 ( .C1(n9051), .C2(n8932), .A(n8824), .B(n8823), .ZN(
        P2_U3211) );
  NAND2_X1 U10328 ( .A1(n8826), .A2(n8825), .ZN(n8827) );
  XNOR2_X1 U10329 ( .A(n8827), .B(n8828), .ZN(n9057) );
  INV_X1 U10330 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8835) );
  OR3_X1 U10331 ( .A1(n8842), .A2(n8829), .A3(n8828), .ZN(n8830) );
  NAND2_X1 U10332 ( .A1(n8831), .A2(n8830), .ZN(n8834) );
  AOI222_X1 U10333 ( .A1(n10257), .A2(n8834), .B1(n8833), .B2(n10262), .C1(
        n8832), .C2(n10261), .ZN(n9052) );
  MUX2_X1 U10334 ( .A(n8835), .B(n9052), .S(n10269), .Z(n8838) );
  AOI22_X1 U10335 ( .A1(n9054), .A2(n8929), .B1(n8942), .B2(n8836), .ZN(n8837)
         );
  OAI211_X1 U10336 ( .C1(n9057), .C2(n8932), .A(n8838), .B(n8837), .ZN(
        P2_U3212) );
  XNOR2_X1 U10337 ( .A(n8840), .B(n8839), .ZN(n9063) );
  INV_X1 U10338 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8849) );
  INV_X1 U10339 ( .A(n8841), .ZN(n8845) );
  INV_X1 U10340 ( .A(n8842), .ZN(n8843) );
  OAI21_X1 U10341 ( .B1(n8845), .B2(n8844), .A(n8843), .ZN(n8848) );
  AOI222_X1 U10342 ( .A1(n10257), .A2(n8848), .B1(n8847), .B2(n10262), .C1(
        n8846), .C2(n10261), .ZN(n9058) );
  MUX2_X1 U10343 ( .A(n8849), .B(n9058), .S(n10269), .Z(n8852) );
  AOI22_X1 U10344 ( .A1(n9060), .A2(n8929), .B1(n8942), .B2(n8850), .ZN(n8851)
         );
  OAI211_X1 U10345 ( .C1(n9063), .C2(n8932), .A(n8852), .B(n8851), .ZN(
        P2_U3213) );
  NAND2_X1 U10346 ( .A1(n8854), .A2(n8853), .ZN(n8856) );
  XNOR2_X1 U10347 ( .A(n8856), .B(n8855), .ZN(n8857) );
  OAI222_X1 U10348 ( .A1(n8910), .A2(n8858), .B1(n8908), .B2(n8893), .C1(n8857), .C2(n8871), .ZN(n8975) );
  OR2_X1 U10349 ( .A1(n8860), .A2(n8859), .ZN(n8861) );
  NAND2_X1 U10350 ( .A1(n8862), .A2(n8861), .ZN(n9067) );
  AOI22_X1 U10351 ( .A1(n8942), .A2(n8863), .B1(n10272), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n8865) );
  NAND2_X1 U10352 ( .A1(n8976), .A2(n8929), .ZN(n8864) );
  OAI211_X1 U10353 ( .C1(n9067), .C2(n8932), .A(n8865), .B(n8864), .ZN(n8866)
         );
  AOI21_X1 U10354 ( .B1(n8975), .B2(n10269), .A(n8866), .ZN(n8867) );
  INV_X1 U10355 ( .A(n8867), .ZN(P2_U3214) );
  NAND2_X1 U10356 ( .A1(n8888), .A2(n8868), .ZN(n8889) );
  NAND2_X1 U10357 ( .A1(n8889), .A2(n8869), .ZN(n8870) );
  XNOR2_X1 U10358 ( .A(n8870), .B(n8876), .ZN(n8872) );
  OAI222_X1 U10359 ( .A1(n8910), .A2(n8873), .B1(n8908), .B2(n8911), .C1(n8872), .C2(n8871), .ZN(n8979) );
  INV_X1 U10360 ( .A(n8979), .ZN(n8885) );
  NAND2_X1 U10361 ( .A1(n8875), .A2(n8876), .ZN(n8877) );
  NAND2_X1 U10362 ( .A1(n8874), .A2(n8877), .ZN(n9071) );
  INV_X1 U10363 ( .A(n9071), .ZN(n8883) );
  AOI22_X1 U10364 ( .A1(n10272), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8942), 
        .B2(n8878), .ZN(n8879) );
  OAI21_X1 U10365 ( .B1(n8881), .B2(n8880), .A(n8879), .ZN(n8882) );
  AOI21_X1 U10366 ( .B1(n8883), .B2(n8945), .A(n8882), .ZN(n8884) );
  OAI21_X1 U10367 ( .B1(n8885), .B2(n10272), .A(n8884), .ZN(P2_U3215) );
  XNOR2_X1 U10368 ( .A(n8886), .B(n8890), .ZN(n9076) );
  AND2_X1 U10369 ( .A1(n8888), .A2(n8887), .ZN(n8891) );
  OAI211_X1 U10370 ( .C1(n8891), .C2(n8890), .A(n8889), .B(n10257), .ZN(n8896)
         );
  OAI22_X1 U10371 ( .A1(n8893), .A2(n8910), .B1(n8892), .B2(n8908), .ZN(n8894)
         );
  INV_X1 U10372 ( .A(n8894), .ZN(n8895) );
  AND2_X1 U10373 ( .A1(n8896), .A2(n8895), .ZN(n9072) );
  MUX2_X1 U10374 ( .A(n9072), .B(n8897), .S(n10272), .Z(n8900) );
  AOI22_X1 U10375 ( .A1(n9073), .A2(n8929), .B1(n8942), .B2(n8898), .ZN(n8899)
         );
  OAI211_X1 U10376 ( .C1(n9076), .C2(n8932), .A(n8900), .B(n8899), .ZN(
        P2_U3216) );
  OR2_X1 U10377 ( .A1(n8923), .A2(n8901), .ZN(n8904) );
  NAND2_X1 U10378 ( .A1(n8904), .A2(n8902), .ZN(n8907) );
  NAND2_X1 U10379 ( .A1(n8904), .A2(n8903), .ZN(n8905) );
  NAND2_X1 U10380 ( .A1(n8905), .A2(n8915), .ZN(n8906) );
  NAND3_X1 U10381 ( .A1(n8907), .A2(n10257), .A3(n8906), .ZN(n8914) );
  OAI22_X1 U10382 ( .A1(n8911), .A2(n8910), .B1(n8909), .B2(n8908), .ZN(n8912)
         );
  INV_X1 U10383 ( .A(n8912), .ZN(n8913) );
  NAND2_X1 U10384 ( .A1(n8914), .A2(n8913), .ZN(n9077) );
  MUX2_X1 U10385 ( .A(n9077), .B(P2_REG2_REG_16__SCAN_IN), .S(n10272), .Z(
        n8920) );
  XNOR2_X1 U10386 ( .A(n4308), .B(n8915), .ZN(n9080) );
  AOI22_X1 U10387 ( .A1(n8986), .A2(n8929), .B1(n8942), .B2(n8917), .ZN(n8918)
         );
  OAI21_X1 U10388 ( .B1(n9080), .B2(n8932), .A(n8918), .ZN(n8919) );
  XOR2_X1 U10389 ( .A(n8921), .B(n8922), .Z(n9089) );
  XNOR2_X1 U10390 ( .A(n8923), .B(n8922), .ZN(n8926) );
  AOI222_X1 U10391 ( .A1(n10257), .A2(n8926), .B1(n8925), .B2(n10262), .C1(
        n8924), .C2(n10261), .ZN(n9083) );
  MUX2_X1 U10392 ( .A(n8927), .B(n9083), .S(n10269), .Z(n8931) );
  AOI22_X1 U10393 ( .A1(n9085), .A2(n8929), .B1(n8942), .B2(n8928), .ZN(n8930)
         );
  OAI211_X1 U10394 ( .C1(n9089), .C2(n8932), .A(n8931), .B(n8930), .ZN(
        P2_U3218) );
  NOR2_X1 U10395 ( .A1(n8933), .A2(n10251), .ZN(n8940) );
  XNOR2_X1 U10396 ( .A(n8934), .B(n8935), .ZN(n8938) );
  AOI222_X1 U10397 ( .A1(n10257), .A2(n8938), .B1(n8937), .B2(n10262), .C1(
        n8936), .C2(n10261), .ZN(n9090) );
  INV_X1 U10398 ( .A(n9090), .ZN(n8939) );
  AOI211_X1 U10399 ( .C1(n8942), .C2(n8941), .A(n8940), .B(n8939), .ZN(n8947)
         );
  XNOR2_X1 U10400 ( .A(n8943), .B(n8944), .ZN(n9093) );
  AOI22_X1 U10401 ( .A1(n9093), .A2(n8945), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n10272), .ZN(n8946) );
  OAI21_X1 U10402 ( .B1(n8947), .B2(n10272), .A(n8946), .ZN(P2_U3219) );
  NAND2_X1 U10403 ( .A1(n9010), .A2(n10323), .ZN(n8950) );
  NAND2_X1 U10404 ( .A1(n10320), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8948) );
  OAI211_X1 U10405 ( .C1(n9012), .C2(n6292), .A(n8950), .B(n8948), .ZN(
        P2_U3490) );
  NAND2_X1 U10406 ( .A1(n8949), .A2(n8994), .ZN(n8951) );
  OAI211_X1 U10407 ( .C1(n10323), .C2(n8952), .A(n8951), .B(n8950), .ZN(
        P2_U3489) );
  INV_X1 U10408 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8954) );
  MUX2_X1 U10409 ( .A(n8954), .B(n9022), .S(n10323), .Z(n8956) );
  NAND2_X1 U10410 ( .A1(n9024), .A2(n8994), .ZN(n8955) );
  OAI211_X1 U10411 ( .C1(n8992), .C2(n9027), .A(n8956), .B(n8955), .ZN(
        P2_U3485) );
  INV_X1 U10412 ( .A(n8957), .ZN(n9028) );
  MUX2_X1 U10413 ( .A(n8958), .B(n9028), .S(n10323), .Z(n8960) );
  AOI22_X1 U10414 ( .A1(n9031), .A2(n6511), .B1(n8994), .B2(n9030), .ZN(n8959)
         );
  NAND2_X1 U10415 ( .A1(n8960), .A2(n8959), .ZN(P2_U3484) );
  MUX2_X1 U10416 ( .A(n8961), .B(n9034), .S(n10323), .Z(n8963) );
  NAND2_X1 U10417 ( .A1(n9036), .A2(n8994), .ZN(n8962) );
  OAI211_X1 U10418 ( .C1(n8992), .C2(n9039), .A(n8963), .B(n8962), .ZN(
        P2_U3483) );
  MUX2_X1 U10419 ( .A(n9952), .B(n9040), .S(n10323), .Z(n8965) );
  AOI22_X1 U10420 ( .A1(n9043), .A2(n6511), .B1(n8994), .B2(n9042), .ZN(n8964)
         );
  NAND2_X1 U10421 ( .A1(n8965), .A2(n8964), .ZN(P2_U3482) );
  MUX2_X1 U10422 ( .A(n8966), .B(n9046), .S(n10323), .Z(n8968) );
  NAND2_X1 U10423 ( .A1(n9048), .A2(n8994), .ZN(n8967) );
  OAI211_X1 U10424 ( .C1(n9051), .C2(n8992), .A(n8968), .B(n8967), .ZN(
        P2_U3481) );
  MUX2_X1 U10425 ( .A(n8969), .B(n9052), .S(n10323), .Z(n8971) );
  NAND2_X1 U10426 ( .A1(n9054), .A2(n8994), .ZN(n8970) );
  OAI211_X1 U10427 ( .C1(n8992), .C2(n9057), .A(n8971), .B(n8970), .ZN(
        P2_U3480) );
  MUX2_X1 U10428 ( .A(n8972), .B(n9058), .S(n10323), .Z(n8974) );
  NAND2_X1 U10429 ( .A1(n9060), .A2(n8994), .ZN(n8973) );
  OAI211_X1 U10430 ( .C1(n9063), .C2(n8992), .A(n8974), .B(n8973), .ZN(
        P2_U3479) );
  AOI21_X1 U10431 ( .B1(n10300), .B2(n8976), .A(n8975), .ZN(n9064) );
  MUX2_X1 U10432 ( .A(n8977), .B(n9064), .S(n10323), .Z(n8978) );
  OAI21_X1 U10433 ( .B1(n8992), .B2(n9067), .A(n8978), .ZN(P2_U3478) );
  AOI21_X1 U10434 ( .B1(n10300), .B2(n8980), .A(n8979), .ZN(n9068) );
  MUX2_X1 U10435 ( .A(n8981), .B(n9068), .S(n10323), .Z(n8982) );
  OAI21_X1 U10436 ( .B1(n8992), .B2(n9071), .A(n8982), .ZN(P2_U3477) );
  MUX2_X1 U10437 ( .A(n8983), .B(n9072), .S(n10323), .Z(n8985) );
  NAND2_X1 U10438 ( .A1(n9073), .A2(n8994), .ZN(n8984) );
  OAI211_X1 U10439 ( .C1(n9076), .C2(n8992), .A(n8985), .B(n8984), .ZN(
        P2_U3476) );
  MUX2_X1 U10440 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9077), .S(n10323), .Z(
        n8988) );
  INV_X1 U10441 ( .A(n8986), .ZN(n9079) );
  OAI22_X1 U10442 ( .A1(n9080), .A2(n8992), .B1(n9079), .B2(n6292), .ZN(n8987)
         );
  MUX2_X1 U10443 ( .A(n8989), .B(n9083), .S(n10323), .Z(n8991) );
  NAND2_X1 U10444 ( .A1(n9085), .A2(n8994), .ZN(n8990) );
  OAI211_X1 U10445 ( .C1(n9089), .C2(n8992), .A(n8991), .B(n8990), .ZN(
        P2_U3474) );
  MUX2_X1 U10446 ( .A(n8993), .B(n9090), .S(n10323), .Z(n8996) );
  AOI22_X1 U10447 ( .A1(n9093), .A2(n6511), .B1(n8994), .B2(n9092), .ZN(n8995)
         );
  NAND2_X1 U10448 ( .A1(n8996), .A2(n8995), .ZN(P2_U3473) );
  INV_X1 U10449 ( .A(n8997), .ZN(n9000) );
  NAND2_X1 U10450 ( .A1(n8998), .A2(n10293), .ZN(n8999) );
  OAI21_X1 U10451 ( .B1(n9000), .B2(n10302), .A(n8999), .ZN(n9001) );
  OR2_X1 U10452 ( .A1(n9002), .A2(n9001), .ZN(n9096) );
  MUX2_X1 U10453 ( .A(n9096), .B(P2_REG1_REG_11__SCAN_IN), .S(n10320), .Z(
        P2_U3470) );
  OAI21_X1 U10454 ( .B1(n10293), .B2(n10257), .A(n9003), .ZN(n9008) );
  NAND2_X1 U10455 ( .A1(n9004), .A2(n10300), .ZN(n9005) );
  AND2_X1 U10456 ( .A1(n9006), .A2(n9005), .ZN(n9007) );
  AND2_X1 U10457 ( .A1(n9008), .A2(n9007), .ZN(n10273) );
  INV_X1 U10458 ( .A(n10273), .ZN(n9009) );
  MUX2_X1 U10459 ( .A(n9009), .B(P2_REG1_REG_0__SCAN_IN), .S(n10320), .Z(
        P2_U3459) );
  NAND2_X1 U10460 ( .A1(n9010), .A2(n10308), .ZN(n9014) );
  NAND2_X1 U10461 ( .A1(n10310), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9011) );
  OAI211_X1 U10462 ( .C1(n9012), .C2(n9078), .A(n9014), .B(n9011), .ZN(
        P2_U3458) );
  NAND2_X1 U10463 ( .A1(n10310), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9013) );
  OAI211_X1 U10464 ( .C1(n9015), .C2(n9078), .A(n9014), .B(n9013), .ZN(
        P2_U3457) );
  INV_X1 U10465 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9017) );
  MUX2_X1 U10466 ( .A(n9017), .B(n9016), .S(n10308), .Z(n9020) );
  NAND2_X1 U10467 ( .A1(n9018), .A2(n6278), .ZN(n9019) );
  OAI211_X1 U10468 ( .C1(n9021), .C2(n9088), .A(n9020), .B(n9019), .ZN(
        P2_U3454) );
  INV_X1 U10469 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9023) );
  MUX2_X1 U10470 ( .A(n9023), .B(n9022), .S(n10308), .Z(n9026) );
  NAND2_X1 U10471 ( .A1(n9024), .A2(n6278), .ZN(n9025) );
  OAI211_X1 U10472 ( .C1(n9027), .C2(n9088), .A(n9026), .B(n9025), .ZN(
        P2_U3453) );
  INV_X1 U10473 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9029) );
  MUX2_X1 U10474 ( .A(n9029), .B(n9028), .S(n10308), .Z(n9033) );
  AOI22_X1 U10475 ( .A1(n9031), .A2(n6198), .B1(n6278), .B2(n9030), .ZN(n9032)
         );
  NAND2_X1 U10476 ( .A1(n9033), .A2(n9032), .ZN(P2_U3452) );
  INV_X1 U10477 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9035) );
  MUX2_X1 U10478 ( .A(n9035), .B(n9034), .S(n10308), .Z(n9038) );
  NAND2_X1 U10479 ( .A1(n9036), .A2(n6278), .ZN(n9037) );
  OAI211_X1 U10480 ( .C1(n9039), .C2(n9088), .A(n9038), .B(n9037), .ZN(
        P2_U3451) );
  INV_X1 U10481 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9041) );
  MUX2_X1 U10482 ( .A(n9041), .B(n9040), .S(n10308), .Z(n9045) );
  AOI22_X1 U10483 ( .A1(n9043), .A2(n6198), .B1(n6278), .B2(n9042), .ZN(n9044)
         );
  NAND2_X1 U10484 ( .A1(n9045), .A2(n9044), .ZN(P2_U3450) );
  INV_X1 U10485 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9047) );
  MUX2_X1 U10486 ( .A(n9047), .B(n9046), .S(n10308), .Z(n9050) );
  NAND2_X1 U10487 ( .A1(n9048), .A2(n6278), .ZN(n9049) );
  OAI211_X1 U10488 ( .C1(n9051), .C2(n9088), .A(n9050), .B(n9049), .ZN(
        P2_U3449) );
  INV_X1 U10489 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9053) );
  MUX2_X1 U10490 ( .A(n9053), .B(n9052), .S(n10308), .Z(n9056) );
  NAND2_X1 U10491 ( .A1(n9054), .A2(n6278), .ZN(n9055) );
  OAI211_X1 U10492 ( .C1(n9057), .C2(n9088), .A(n9056), .B(n9055), .ZN(
        P2_U3448) );
  INV_X1 U10493 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9059) );
  MUX2_X1 U10494 ( .A(n9059), .B(n9058), .S(n10308), .Z(n9062) );
  NAND2_X1 U10495 ( .A1(n9060), .A2(n6278), .ZN(n9061) );
  OAI211_X1 U10496 ( .C1(n9063), .C2(n9088), .A(n9062), .B(n9061), .ZN(
        P2_U3447) );
  INV_X1 U10497 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9065) );
  MUX2_X1 U10498 ( .A(n9065), .B(n9064), .S(n10308), .Z(n9066) );
  OAI21_X1 U10499 ( .B1(n9067), .B2(n9088), .A(n9066), .ZN(P2_U3446) );
  INV_X1 U10500 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9069) );
  MUX2_X1 U10501 ( .A(n9069), .B(n9068), .S(n10308), .Z(n9070) );
  OAI21_X1 U10502 ( .B1(n9071), .B2(n9088), .A(n9070), .ZN(P2_U3444) );
  MUX2_X1 U10503 ( .A(n9072), .B(n9943), .S(n10310), .Z(n9075) );
  NAND2_X1 U10504 ( .A1(n9073), .A2(n6278), .ZN(n9074) );
  OAI211_X1 U10505 ( .C1(n9076), .C2(n9088), .A(n9075), .B(n9074), .ZN(
        P2_U3441) );
  MUX2_X1 U10506 ( .A(n9077), .B(P2_REG0_REG_16__SCAN_IN), .S(n10310), .Z(
        n9082) );
  OAI22_X1 U10507 ( .A1(n9080), .A2(n9088), .B1(n9079), .B2(n9078), .ZN(n9081)
         );
  INV_X1 U10508 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9084) );
  MUX2_X1 U10509 ( .A(n9084), .B(n9083), .S(n10308), .Z(n9087) );
  NAND2_X1 U10510 ( .A1(n9085), .A2(n6278), .ZN(n9086) );
  OAI211_X1 U10511 ( .C1(n9089), .C2(n9088), .A(n9087), .B(n9086), .ZN(
        P2_U3435) );
  INV_X1 U10512 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9091) );
  MUX2_X1 U10513 ( .A(n9091), .B(n9090), .S(n10308), .Z(n9095) );
  AOI22_X1 U10514 ( .A1(n9093), .A2(n6198), .B1(n6278), .B2(n9092), .ZN(n9094)
         );
  NAND2_X1 U10515 ( .A1(n9095), .A2(n9094), .ZN(P2_U3432) );
  MUX2_X1 U10516 ( .A(n9096), .B(P2_REG0_REG_11__SCAN_IN), .S(n10310), .Z(
        P2_U3423) );
  OAI222_X1 U10517 ( .A1(n9101), .A2(n9097), .B1(n5717), .B2(P2_U3151), .C1(
        n9106), .C2(n10000), .ZN(P2_U3266) );
  INV_X1 U10518 ( .A(n9098), .ZN(n10003) );
  OAI222_X1 U10519 ( .A1(n9106), .A2(n10003), .B1(n6472), .B2(P2_U3151), .C1(
        n9099), .C2(n9101), .ZN(P2_U3268) );
  OAI222_X1 U10520 ( .A1(n9106), .A2(n9105), .B1(P2_U3151), .B2(n9103), .C1(
        n9102), .C2(n9101), .ZN(P2_U3269) );
  MUX2_X1 U10521 ( .A(n9107), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10522 ( .A(n9108), .ZN(n9109) );
  NAND2_X1 U10523 ( .A1(n9110), .A2(n9109), .ZN(n9123) );
  NAND2_X1 U10524 ( .A1(n9715), .A2(n9189), .ZN(n9112) );
  OR2_X1 U10525 ( .A1(n9116), .A2(n7791), .ZN(n9111) );
  NAND2_X1 U10526 ( .A1(n9112), .A2(n9111), .ZN(n9114) );
  XNOR2_X1 U10527 ( .A(n9114), .B(n4310), .ZN(n9119) );
  INV_X1 U10528 ( .A(n9119), .ZN(n9121) );
  NOR2_X1 U10529 ( .A1(n9116), .A2(n9115), .ZN(n9117) );
  AOI21_X1 U10530 ( .B1(n9715), .B2(n7861), .A(n9117), .ZN(n9118) );
  INV_X1 U10531 ( .A(n9118), .ZN(n9120) );
  AOI21_X1 U10532 ( .B1(n9121), .B2(n9120), .A(n9204), .ZN(n9122) );
  AOI21_X1 U10533 ( .B1(n9127), .B2(n9123), .A(n9122), .ZN(n9128) );
  INV_X1 U10534 ( .A(n9122), .ZN(n9125) );
  INV_X1 U10535 ( .A(n9123), .ZN(n9124) );
  NOR2_X1 U10536 ( .A1(n9125), .A2(n9124), .ZN(n9126) );
  OAI21_X1 U10537 ( .B1(n9128), .B2(n9197), .A(n9349), .ZN(n9132) );
  AOI22_X1 U10538 ( .A1(n9375), .A2(n9314), .B1(n9313), .B2(n9377), .ZN(n9523)
         );
  AOI22_X1 U10539 ( .A1(n9526), .A2(n9364), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n9129) );
  OAI21_X1 U10540 ( .B1(n9523), .B2(n9366), .A(n9129), .ZN(n9130) );
  AOI21_X1 U10541 ( .B1(n9715), .B2(n9369), .A(n9130), .ZN(n9131) );
  NAND2_X1 U10542 ( .A1(n9132), .A2(n9131), .ZN(P1_U3214) );
  NOR2_X1 U10543 ( .A1(n9133), .A2(n9134), .ZN(n9235) );
  AOI21_X1 U10544 ( .B1(n9134), .B2(n9133), .A(n9235), .ZN(n9135) );
  NAND2_X1 U10545 ( .A1(n9135), .A2(n9136), .ZN(n9237) );
  OAI21_X1 U10546 ( .B1(n9136), .B2(n9135), .A(n9237), .ZN(n9137) );
  NAND2_X1 U10547 ( .A1(n9137), .A2(n9349), .ZN(n9142) );
  NAND2_X1 U10548 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10027)
         );
  OAI21_X1 U10549 ( .B1(n9366), .B2(n9138), .A(n10027), .ZN(n9139) );
  AOI21_X1 U10550 ( .B1(n9140), .B2(n9364), .A(n9139), .ZN(n9141) );
  OAI211_X1 U10551 ( .C1(n9143), .C2(n9332), .A(n9142), .B(n9141), .ZN(
        P1_U3215) );
  INV_X1 U10552 ( .A(n9144), .ZN(n9145) );
  NAND2_X1 U10553 ( .A1(n9146), .A2(n9145), .ZN(n9147) );
  OAI21_X1 U10554 ( .B1(n9146), .B2(n9145), .A(n9147), .ZN(n9311) );
  NOR2_X1 U10555 ( .A1(n9311), .A2(n9312), .ZN(n9310) );
  INV_X1 U10556 ( .A(n9147), .ZN(n9148) );
  NOR3_X1 U10557 ( .A1(n9310), .A2(n9149), .A3(n9148), .ZN(n9151) );
  INV_X1 U10558 ( .A(n9150), .ZN(n9263) );
  OAI21_X1 U10559 ( .B1(n9151), .B2(n9263), .A(n9349), .ZN(n9158) );
  NAND2_X1 U10560 ( .A1(n9379), .A2(n9314), .ZN(n9153) );
  NAND2_X1 U10561 ( .A1(n9381), .A2(n9313), .ZN(n9152) );
  NAND2_X1 U10562 ( .A1(n9153), .A2(n9152), .ZN(n9592) );
  INV_X1 U10563 ( .A(n9595), .ZN(n9155) );
  OAI22_X1 U10564 ( .A1(n9155), .A2(n9342), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9154), .ZN(n9156) );
  AOI21_X1 U10565 ( .B1(n9592), .B2(n9356), .A(n9156), .ZN(n9157) );
  OAI211_X1 U10566 ( .C1(n9598), .C2(n9332), .A(n9158), .B(n9157), .ZN(
        P1_U3216) );
  INV_X1 U10567 ( .A(n9159), .ZN(n9161) );
  NAND2_X1 U10568 ( .A1(n9161), .A2(n9160), .ZN(n9320) );
  OAI21_X1 U10569 ( .B1(n9161), .B2(n9160), .A(n9320), .ZN(n9162) );
  NOR2_X1 U10570 ( .A1(n9162), .A2(n9163), .ZN(n9323) );
  AOI21_X1 U10571 ( .B1(n9163), .B2(n9162), .A(n9323), .ZN(n9171) );
  AOI21_X1 U10572 ( .B1(n9356), .B2(n9165), .A(n9164), .ZN(n9166) );
  OAI21_X1 U10573 ( .B1(n9167), .B2(n9342), .A(n9166), .ZN(n9168) );
  AOI21_X1 U10574 ( .B1(n9169), .B2(n9369), .A(n9168), .ZN(n9170) );
  OAI21_X1 U10575 ( .B1(n9171), .B2(n9371), .A(n9170), .ZN(P1_U3217) );
  OAI21_X1 U10576 ( .B1(n9173), .B2(n9172), .A(n6968), .ZN(n9174) );
  NAND2_X1 U10577 ( .A1(n9174), .A2(n9349), .ZN(n9179) );
  AOI22_X1 U10578 ( .A1(n9356), .A2(n9176), .B1(n9369), .B2(n9175), .ZN(n9178)
         );
  MUX2_X1 U10579 ( .A(n9342), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n9177) );
  NAND3_X1 U10580 ( .A1(n9179), .A2(n9178), .A3(n9177), .ZN(P1_U3218) );
  NOR2_X1 U10581 ( .A1(n9180), .A2(n4395), .ZN(n9181) );
  XNOR2_X1 U10582 ( .A(n9182), .B(n9181), .ZN(n9188) );
  NOR2_X1 U10583 ( .A1(n9342), .A2(n9661), .ZN(n9186) );
  AND2_X1 U10584 ( .A1(n9385), .A2(n9313), .ZN(n9183) );
  AOI21_X1 U10585 ( .B1(n9383), .B2(n9314), .A(n9183), .ZN(n9654) );
  OAI22_X1 U10586 ( .A1(n9654), .A2(n9366), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9184), .ZN(n9185) );
  AOI211_X1 U10587 ( .C1(n9822), .C2(n9369), .A(n9186), .B(n9185), .ZN(n9187)
         );
  OAI21_X1 U10588 ( .B1(n9188), .B2(n9371), .A(n9187), .ZN(P1_U3219) );
  NAND2_X1 U10589 ( .A1(n9203), .A2(n9189), .ZN(n9191) );
  NAND2_X1 U10590 ( .A1(n9375), .A2(n7710), .ZN(n9190) );
  NAND2_X1 U10591 ( .A1(n9191), .A2(n9190), .ZN(n9193) );
  XNOR2_X1 U10592 ( .A(n9193), .B(n9192), .ZN(n9196) );
  AOI22_X1 U10593 ( .A1(n9203), .A2(n7861), .B1(n9194), .B2(n9375), .ZN(n9195)
         );
  XNOR2_X1 U10594 ( .A(n9196), .B(n9195), .ZN(n9205) );
  NOR2_X1 U10595 ( .A1(n9198), .A2(n9366), .ZN(n9202) );
  OAI22_X1 U10596 ( .A1(n9200), .A2(n9342), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9199), .ZN(n9201) );
  AOI211_X1 U10597 ( .C1(n9203), .C2(n9369), .A(n9202), .B(n9201), .ZN(n9206)
         );
  XOR2_X1 U10598 ( .A(n9274), .B(n9275), .Z(n9209) );
  INV_X1 U10599 ( .A(n9207), .ZN(n9208) );
  NAND2_X1 U10600 ( .A1(n9209), .A2(n9208), .ZN(n9273) );
  OAI21_X1 U10601 ( .B1(n9209), .B2(n9208), .A(n9273), .ZN(n9210) );
  NAND2_X1 U10602 ( .A1(n9210), .A2(n9349), .ZN(n9214) );
  OAI22_X1 U10603 ( .A1(n9354), .A2(n9351), .B1(n9211), .B2(n9353), .ZN(n10097) );
  AOI22_X1 U10604 ( .A1(n9356), .A2(n10097), .B1(P1_REG3_REG_8__SCAN_IN), .B2(
        P1_U3086), .ZN(n9213) );
  AOI22_X1 U10605 ( .A1(n9369), .A2(n10101), .B1(n9364), .B2(n10099), .ZN(
        n9212) );
  NAND3_X1 U10606 ( .A1(n9214), .A2(n9213), .A3(n9212), .ZN(P1_U3221) );
  OAI21_X1 U10607 ( .B1(n9217), .B2(n9216), .A(n9215), .ZN(n9218) );
  NAND2_X1 U10608 ( .A1(n9218), .A2(n9349), .ZN(n9222) );
  AOI22_X1 U10609 ( .A1(n9381), .A2(n9314), .B1(n9313), .B2(n9383), .ZN(n9626)
         );
  OAI22_X1 U10610 ( .A1(n9626), .A2(n9366), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9219), .ZN(n9220) );
  AOI21_X1 U10611 ( .B1(n9630), .B2(n9364), .A(n9220), .ZN(n9221) );
  OAI211_X1 U10612 ( .C1(n9813), .C2(n9332), .A(n9222), .B(n9221), .ZN(
        P1_U3223) );
  AND3_X1 U10613 ( .A1(n9223), .A2(n9225), .A3(n9224), .ZN(n9226) );
  OAI21_X1 U10614 ( .B1(n9227), .B2(n9226), .A(n9349), .ZN(n9233) );
  OAI21_X1 U10615 ( .B1(n9366), .B2(n9229), .A(n9228), .ZN(n9230) );
  AOI21_X1 U10616 ( .B1(n9231), .B2(n9364), .A(n9230), .ZN(n9232) );
  OAI211_X1 U10617 ( .C1(n9234), .C2(n9332), .A(n9233), .B(n9232), .ZN(
        P1_U3224) );
  INV_X1 U10618 ( .A(n9764), .ZN(n9698) );
  INV_X1 U10619 ( .A(n9235), .ZN(n9236) );
  NAND2_X1 U10620 ( .A1(n9237), .A2(n9236), .ZN(n9239) );
  NAND2_X1 U10621 ( .A1(n9239), .A2(n9238), .ZN(n9240) );
  OAI21_X1 U10622 ( .B1(n9239), .B2(n9238), .A(n9240), .ZN(n9361) );
  NOR2_X1 U10623 ( .A1(n9361), .A2(n9362), .ZN(n9360) );
  INV_X1 U10624 ( .A(n9240), .ZN(n9241) );
  NOR3_X1 U10625 ( .A1(n9360), .A2(n9242), .A3(n9241), .ZN(n9245) );
  INV_X1 U10626 ( .A(n9243), .ZN(n9244) );
  OAI21_X1 U10627 ( .B1(n9245), .B2(n9244), .A(n9349), .ZN(n9250) );
  INV_X1 U10628 ( .A(n9246), .ZN(n9695) );
  AND2_X1 U10629 ( .A1(n9388), .A2(n9313), .ZN(n9247) );
  AOI21_X1 U10630 ( .B1(n9386), .B2(n9314), .A(n9247), .ZN(n9702) );
  NAND2_X1 U10631 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10054)
         );
  OAI21_X1 U10632 ( .B1(n9366), .B2(n9702), .A(n10054), .ZN(n9248) );
  AOI21_X1 U10633 ( .B1(n9695), .B2(n9364), .A(n9248), .ZN(n9249) );
  OAI211_X1 U10634 ( .C1(n9698), .C2(n9332), .A(n9250), .B(n9249), .ZN(
        P1_U3226) );
  OAI21_X1 U10635 ( .B1(n9253), .B2(n9252), .A(n9251), .ZN(n9254) );
  NAND2_X1 U10636 ( .A1(n9254), .A2(n9349), .ZN(n9259) );
  NAND2_X1 U10637 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10071)
         );
  OAI21_X1 U10638 ( .B1(n9255), .B2(n9366), .A(n10071), .ZN(n9256) );
  AOI21_X1 U10639 ( .B1(n9257), .B2(n9364), .A(n9256), .ZN(n9258) );
  OAI211_X1 U10640 ( .C1(n9260), .C2(n9332), .A(n9259), .B(n9258), .ZN(
        P1_U3228) );
  INV_X1 U10641 ( .A(n9578), .ZN(n9574) );
  NOR3_X1 U10642 ( .A1(n9263), .A2(n9262), .A3(n9261), .ZN(n9266) );
  INV_X1 U10643 ( .A(n9264), .ZN(n9265) );
  OAI21_X1 U10644 ( .B1(n9266), .B2(n9265), .A(n9349), .ZN(n9272) );
  NAND2_X1 U10645 ( .A1(n9378), .A2(n9314), .ZN(n9268) );
  NAND2_X1 U10646 ( .A1(n9380), .A2(n9313), .ZN(n9267) );
  NAND2_X1 U10647 ( .A1(n9268), .A2(n9267), .ZN(n9568) );
  OAI22_X1 U10648 ( .A1(n9576), .A2(n9342), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9269), .ZN(n9270) );
  AOI21_X1 U10649 ( .B1(n9568), .B2(n9356), .A(n9270), .ZN(n9271) );
  OAI211_X1 U10650 ( .C1(n9574), .C2(n9332), .A(n9272), .B(n9271), .ZN(
        P1_U3229) );
  OAI21_X1 U10651 ( .B1(n9275), .B2(n9274), .A(n9273), .ZN(n9279) );
  XNOR2_X1 U10652 ( .A(n9277), .B(n9276), .ZN(n9278) );
  XNOR2_X1 U10653 ( .A(n9279), .B(n9278), .ZN(n9280) );
  NAND2_X1 U10654 ( .A1(n9280), .A2(n9349), .ZN(n9290) );
  NAND2_X1 U10655 ( .A1(n9282), .A2(n9281), .ZN(n9284) );
  AOI21_X1 U10656 ( .B1(n9356), .B2(n9284), .A(n9283), .ZN(n9289) );
  NAND2_X1 U10657 ( .A1(n9369), .A2(n10224), .ZN(n9288) );
  INV_X1 U10658 ( .A(n9285), .ZN(n9286) );
  NAND2_X1 U10659 ( .A1(n9364), .A2(n9286), .ZN(n9287) );
  NAND4_X1 U10660 ( .A1(n9290), .A2(n9289), .A3(n9288), .A4(n9287), .ZN(
        P1_U3231) );
  OAI21_X1 U10661 ( .B1(n9293), .B2(n9292), .A(n9291), .ZN(n9294) );
  NAND2_X1 U10662 ( .A1(n9294), .A2(n9349), .ZN(n9299) );
  INV_X1 U10663 ( .A(n9295), .ZN(n9647) );
  AOI22_X1 U10664 ( .A1(n9382), .A2(n9314), .B1(n9313), .B2(n9384), .ZN(n9641)
         );
  OAI22_X1 U10665 ( .A1(n9641), .A2(n9366), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9296), .ZN(n9297) );
  AOI21_X1 U10666 ( .B1(n9647), .B2(n9364), .A(n9297), .ZN(n9298) );
  OAI211_X1 U10667 ( .C1(n4808), .C2(n9332), .A(n9299), .B(n9298), .ZN(
        P1_U3233) );
  AOI21_X1 U10668 ( .B1(n9301), .B2(n9300), .A(n4397), .ZN(n9309) );
  NAND2_X1 U10669 ( .A1(n9364), .A2(n9302), .ZN(n9304) );
  OAI211_X1 U10670 ( .C1(n9366), .C2(n9305), .A(n9304), .B(n9303), .ZN(n9306)
         );
  AOI21_X1 U10671 ( .B1(n9307), .B2(n9369), .A(n9306), .ZN(n9308) );
  OAI21_X1 U10672 ( .B1(n9309), .B2(n9371), .A(n9308), .ZN(P1_U3234) );
  AOI21_X1 U10673 ( .B1(n9312), .B2(n9311), .A(n9310), .ZN(n9319) );
  NOR2_X1 U10674 ( .A1(n9613), .A2(n9342), .ZN(n9317) );
  AOI22_X1 U10675 ( .A1(n9380), .A2(n9314), .B1(n9382), .B2(n9313), .ZN(n9609)
         );
  OAI22_X1 U10676 ( .A1(n9609), .A2(n9366), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9315), .ZN(n9316) );
  AOI211_X1 U10677 ( .C1(n9806), .C2(n9369), .A(n9317), .B(n9316), .ZN(n9318)
         );
  OAI21_X1 U10678 ( .B1(n9319), .B2(n9371), .A(n9318), .ZN(P1_U3235) );
  INV_X1 U10679 ( .A(n9320), .ZN(n9321) );
  NOR3_X1 U10680 ( .A1(n9323), .A2(n9322), .A3(n9321), .ZN(n9325) );
  INV_X1 U10681 ( .A(n9223), .ZN(n9324) );
  OAI21_X1 U10682 ( .B1(n9325), .B2(n9324), .A(n9349), .ZN(n9331) );
  NOR2_X1 U10683 ( .A1(n9342), .A2(n9326), .ZN(n9327) );
  AOI211_X1 U10684 ( .C1(n9356), .C2(n9329), .A(n9328), .B(n9327), .ZN(n9330)
         );
  OAI211_X1 U10685 ( .C1(n9333), .C2(n9332), .A(n9331), .B(n9330), .ZN(
        P1_U3236) );
  INV_X1 U10686 ( .A(n9334), .ZN(n9336) );
  NAND2_X1 U10687 ( .A1(n9336), .A2(n9335), .ZN(n9337) );
  XNOR2_X1 U10688 ( .A(n9338), .B(n9337), .ZN(n9345) );
  OAI22_X1 U10689 ( .A1(n9340), .A2(n9353), .B1(n9339), .B2(n9351), .ZN(n9684)
         );
  AOI22_X1 U10690 ( .A1(n9684), .A2(n9356), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n9341) );
  OAI21_X1 U10691 ( .B1(n9676), .B2(n9342), .A(n9341), .ZN(n9343) );
  AOI21_X1 U10692 ( .B1(n9754), .B2(n9369), .A(n9343), .ZN(n9344) );
  OAI21_X1 U10693 ( .B1(n9345), .B2(n9371), .A(n9344), .ZN(P1_U3238) );
  OAI21_X1 U10694 ( .B1(n9348), .B2(n9347), .A(n9346), .ZN(n9350) );
  NAND2_X1 U10695 ( .A1(n9350), .A2(n9349), .ZN(n9359) );
  OAI22_X1 U10696 ( .A1(n9354), .A2(n9353), .B1(n9352), .B2(n9351), .ZN(n10109) );
  NAND2_X1 U10697 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9459) );
  INV_X1 U10698 ( .A(n9459), .ZN(n9355) );
  AOI21_X1 U10699 ( .B1(n9356), .B2(n10109), .A(n9355), .ZN(n9358) );
  AOI22_X1 U10700 ( .A1(n9369), .A2(n10116), .B1(n9364), .B2(n10111), .ZN(
        n9357) );
  NAND3_X1 U10701 ( .A1(n9359), .A2(n9358), .A3(n9357), .ZN(P1_U3239) );
  AOI21_X1 U10702 ( .B1(n9362), .B2(n9361), .A(n9360), .ZN(n9372) );
  NAND2_X1 U10703 ( .A1(n9364), .A2(n9363), .ZN(n9365) );
  NAND2_X1 U10704 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10040)
         );
  OAI211_X1 U10705 ( .C1(n9367), .C2(n9366), .A(n9365), .B(n10040), .ZN(n9368)
         );
  AOI21_X1 U10706 ( .B1(n9835), .B2(n9369), .A(n9368), .ZN(n9370) );
  OAI21_X1 U10707 ( .B1(n9372), .B2(n9371), .A(n9370), .ZN(P1_U3241) );
  MUX2_X1 U10708 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9373), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U10709 ( .A(n9374), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9400), .Z(
        P1_U3584) );
  MUX2_X1 U10710 ( .A(n9375), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9400), .Z(
        P1_U3582) );
  MUX2_X1 U10711 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9376), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10712 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9377), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10713 ( .A(n9378), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9400), .Z(
        P1_U3579) );
  MUX2_X1 U10714 ( .A(n9379), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9400), .Z(
        P1_U3578) );
  MUX2_X1 U10715 ( .A(n9380), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9400), .Z(
        P1_U3577) );
  MUX2_X1 U10716 ( .A(n9381), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9400), .Z(
        P1_U3576) );
  MUX2_X1 U10717 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9382), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10718 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9383), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10719 ( .A(n9384), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9400), .Z(
        P1_U3573) );
  MUX2_X1 U10720 ( .A(n9385), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9400), .Z(
        P1_U3572) );
  MUX2_X1 U10721 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9386), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10722 ( .A(n9387), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9400), .Z(
        P1_U3570) );
  MUX2_X1 U10723 ( .A(n9388), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9400), .Z(
        P1_U3569) );
  MUX2_X1 U10724 ( .A(n9389), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9400), .Z(
        P1_U3568) );
  MUX2_X1 U10725 ( .A(n9390), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9400), .Z(
        P1_U3567) );
  MUX2_X1 U10726 ( .A(n9391), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9400), .Z(
        P1_U3566) );
  MUX2_X1 U10727 ( .A(n9392), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9400), .Z(
        P1_U3565) );
  MUX2_X1 U10728 ( .A(n9393), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9400), .Z(
        P1_U3564) );
  MUX2_X1 U10729 ( .A(n9394), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9400), .Z(
        P1_U3563) );
  MUX2_X1 U10730 ( .A(n9395), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9400), .Z(
        P1_U3562) );
  MUX2_X1 U10731 ( .A(n9396), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9400), .Z(
        P1_U3561) );
  MUX2_X1 U10732 ( .A(n9397), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9400), .Z(
        P1_U3560) );
  MUX2_X1 U10733 ( .A(n9398), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9400), .Z(
        P1_U3559) );
  MUX2_X1 U10734 ( .A(n9399), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9400), .Z(
        P1_U3558) );
  MUX2_X1 U10735 ( .A(n9401), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9400), .Z(
        P1_U3557) );
  MUX2_X1 U10736 ( .A(n9402), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9400), .Z(
        P1_U3555) );
  OAI211_X1 U10737 ( .C1(n9405), .C2(n9404), .A(n10081), .B(n9403), .ZN(n9413)
         );
  OAI211_X1 U10738 ( .C1(n9408), .C2(n9407), .A(n10075), .B(n9406), .ZN(n9412)
         );
  AOI22_X1 U10739 ( .A1(n10014), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9411) );
  NAND2_X1 U10740 ( .A1(n10083), .A2(n9409), .ZN(n9410) );
  NAND4_X1 U10741 ( .A1(n9413), .A2(n9412), .A3(n9411), .A4(n9410), .ZN(
        P1_U3244) );
  INV_X1 U10742 ( .A(n9414), .ZN(n9417) );
  INV_X1 U10743 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9889) );
  NAND2_X1 U10744 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9415) );
  OAI21_X1 U10745 ( .B1(n10089), .B2(n9889), .A(n9415), .ZN(n9416) );
  AOI21_X1 U10746 ( .B1(n9417), .B2(n10083), .A(n9416), .ZN(n9426) );
  OAI211_X1 U10747 ( .C1(n9420), .C2(n9419), .A(n10075), .B(n9418), .ZN(n9425)
         );
  OAI211_X1 U10748 ( .C1(n9423), .C2(n9422), .A(n10081), .B(n9421), .ZN(n9424)
         );
  NAND3_X1 U10749 ( .A1(n9426), .A2(n9425), .A3(n9424), .ZN(P1_U3246) );
  AOI21_X1 U10750 ( .B1(n10014), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n9427), .ZN(
        n9428) );
  OAI21_X1 U10751 ( .B1(n9429), .B2(n10069), .A(n9428), .ZN(n9430) );
  INV_X1 U10752 ( .A(n9430), .ZN(n9440) );
  INV_X1 U10753 ( .A(n9431), .ZN(n9432) );
  OAI211_X1 U10754 ( .C1(n9434), .C2(n9433), .A(n10081), .B(n9432), .ZN(n9439)
         );
  OAI211_X1 U10755 ( .C1(n9437), .C2(n9436), .A(n10075), .B(n9435), .ZN(n9438)
         );
  NAND4_X1 U10756 ( .A1(n9441), .A2(n9440), .A3(n9439), .A4(n9438), .ZN(
        P1_U3247) );
  AOI211_X1 U10757 ( .C1(n9444), .C2(n9443), .A(n10030), .B(n9442), .ZN(n9445)
         );
  INV_X1 U10758 ( .A(n9445), .ZN(n9454) );
  INV_X1 U10759 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9941) );
  NAND2_X1 U10760 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9446) );
  OAI21_X1 U10761 ( .B1(n10089), .B2(n9941), .A(n9446), .ZN(n9447) );
  AOI21_X1 U10762 ( .B1(n9448), .B2(n10083), .A(n9447), .ZN(n9453) );
  OAI211_X1 U10763 ( .C1(n9451), .C2(n9450), .A(n10075), .B(n9449), .ZN(n9452)
         );
  NAND3_X1 U10764 ( .A1(n9454), .A2(n9453), .A3(n9452), .ZN(P1_U3248) );
  AOI211_X1 U10765 ( .C1(n9457), .C2(n9456), .A(n10030), .B(n9455), .ZN(n9458)
         );
  INV_X1 U10766 ( .A(n9458), .ZN(n9468) );
  INV_X1 U10767 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9460) );
  OAI21_X1 U10768 ( .B1(n10089), .B2(n9460), .A(n9459), .ZN(n9461) );
  AOI21_X1 U10769 ( .B1(n9462), .B2(n10083), .A(n9461), .ZN(n9467) );
  OAI211_X1 U10770 ( .C1(n9465), .C2(n9464), .A(n10075), .B(n9463), .ZN(n9466)
         );
  NAND3_X1 U10771 ( .A1(n9468), .A2(n9467), .A3(n9466), .ZN(P1_U3249) );
  AOI211_X1 U10772 ( .C1(n9471), .C2(n9470), .A(n10030), .B(n9469), .ZN(n9472)
         );
  INV_X1 U10773 ( .A(n9472), .ZN(n9482) );
  INV_X1 U10774 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9474) );
  NAND2_X1 U10775 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9473) );
  OAI21_X1 U10776 ( .B1(n10089), .B2(n9474), .A(n9473), .ZN(n9475) );
  AOI21_X1 U10777 ( .B1(n9476), .B2(n10083), .A(n9475), .ZN(n9481) );
  OAI211_X1 U10778 ( .C1(n9479), .C2(n9478), .A(n9477), .B(n10075), .ZN(n9480)
         );
  NAND3_X1 U10779 ( .A1(n9482), .A2(n9481), .A3(n9480), .ZN(P1_U3250) );
  AOI211_X1 U10780 ( .C1(n9485), .C2(n9484), .A(n10030), .B(n9483), .ZN(n9486)
         );
  INV_X1 U10781 ( .A(n9486), .ZN(n9496) );
  INV_X1 U10782 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9488) );
  NAND2_X1 U10783 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n9487) );
  OAI21_X1 U10784 ( .B1(n10089), .B2(n9488), .A(n9487), .ZN(n9489) );
  AOI21_X1 U10785 ( .B1(n9490), .B2(n10083), .A(n9489), .ZN(n9495) );
  OAI211_X1 U10786 ( .C1(n9493), .C2(n9492), .A(n9491), .B(n10075), .ZN(n9494)
         );
  NAND3_X1 U10787 ( .A1(n9496), .A2(n9495), .A3(n9494), .ZN(P1_U3251) );
  AOI21_X1 U10788 ( .B1(n9503), .B2(n9497), .A(n9693), .ZN(n9499) );
  NAND2_X1 U10789 ( .A1(n9499), .A2(n9498), .ZN(n9710) );
  OAI21_X1 U10790 ( .B1(n9663), .B2(n9501), .A(n9500), .ZN(n9502) );
  AOI21_X1 U10791 ( .B1(n9503), .B2(n10142), .A(n9502), .ZN(n9504) );
  OAI21_X1 U10792 ( .B1(n9710), .B2(n9667), .A(n9504), .ZN(P1_U3264) );
  XNOR2_X1 U10793 ( .A(n9509), .B(n9508), .ZN(n9519) );
  NOR2_X1 U10794 ( .A1(n9510), .A2(n9697), .ZN(n9514) );
  OAI22_X1 U10795 ( .A1(n9512), .A2(n9660), .B1(n9511), .B2(n9663), .ZN(n9513)
         );
  AOI211_X1 U10796 ( .C1(n9515), .C2(n10153), .A(n9514), .B(n9513), .ZN(n9518)
         );
  NAND2_X1 U10797 ( .A1(n9516), .A2(n9663), .ZN(n9517) );
  OAI211_X1 U10798 ( .C1(n9519), .C2(n9708), .A(n9518), .B(n9517), .ZN(
        P1_U3356) );
  XOR2_X2 U10799 ( .A(n9520), .B(n5639), .Z(n9788) );
  XNOR2_X1 U10800 ( .A(n9521), .B(n5640), .ZN(n9522) );
  NAND2_X1 U10801 ( .A1(n9522), .A2(n10140), .ZN(n9524) );
  NAND2_X1 U10802 ( .A1(n9524), .A2(n9523), .ZN(n9714) );
  INV_X1 U10803 ( .A(n9715), .ZN(n9529) );
  AOI211_X1 U10804 ( .C1(n9715), .C2(n9542), .A(n9693), .B(n4342), .ZN(n9713)
         );
  NAND2_X1 U10805 ( .A1(n9713), .A2(n10153), .ZN(n9528) );
  AOI22_X1 U10806 ( .A1(n9526), .A2(n10143), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10130), .ZN(n9527) );
  OAI211_X1 U10807 ( .C1(n9529), .C2(n9697), .A(n9528), .B(n9527), .ZN(n9530)
         );
  AOI21_X1 U10808 ( .B1(n9663), .B2(n9714), .A(n9530), .ZN(n9531) );
  OAI21_X1 U10809 ( .B1(n9788), .B2(n9708), .A(n9531), .ZN(P1_U3266) );
  NAND2_X1 U10810 ( .A1(n9532), .A2(n8047), .ZN(n9534) );
  INV_X1 U10811 ( .A(n9537), .ZN(n9533) );
  XNOR2_X1 U10812 ( .A(n9534), .B(n9533), .ZN(n9536) );
  AOI21_X1 U10813 ( .B1(n9536), .B2(n10140), .A(n9535), .ZN(n9718) );
  XOR2_X1 U10814 ( .A(n9538), .B(n9537), .Z(n9790) );
  INV_X1 U10815 ( .A(n9790), .ZN(n9539) );
  NAND2_X1 U10816 ( .A1(n9539), .A2(n10154), .ZN(n9548) );
  OAI22_X1 U10817 ( .A1(n9541), .A2(n9660), .B1(n9540), .B2(n9663), .ZN(n9545)
         );
  INV_X1 U10818 ( .A(n9557), .ZN(n9543) );
  OAI211_X1 U10819 ( .C1(n9789), .C2(n9543), .A(n9542), .B(n10148), .ZN(n9717)
         );
  NOR2_X1 U10820 ( .A1(n9717), .A2(n9667), .ZN(n9544) );
  AOI211_X1 U10821 ( .C1(n10142), .C2(n9546), .A(n9545), .B(n9544), .ZN(n9547)
         );
  OAI211_X1 U10822 ( .C1(n10130), .C2(n9718), .A(n9548), .B(n9547), .ZN(
        P1_U3267) );
  XNOR2_X1 U10823 ( .A(n9549), .B(n9552), .ZN(n9796) );
  INV_X1 U10824 ( .A(n9550), .ZN(n9551) );
  NOR2_X1 U10825 ( .A1(n9552), .A2(n9551), .ZN(n9553) );
  AOI21_X1 U10826 ( .B1(n9553), .B2(n9567), .A(n9642), .ZN(n9555) );
  AOI21_X1 U10827 ( .B1(n9555), .B2(n9532), .A(n9554), .ZN(n9721) );
  OAI21_X1 U10828 ( .B1(n9556), .B2(n9660), .A(n9721), .ZN(n9561) );
  OAI211_X1 U10829 ( .C1(n9722), .C2(n9581), .A(n10148), .B(n9557), .ZN(n9720)
         );
  AOI22_X1 U10830 ( .A1(n9558), .A2(n10142), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10130), .ZN(n9559) );
  OAI21_X1 U10831 ( .B1(n9720), .B2(n9667), .A(n9559), .ZN(n9560) );
  AOI21_X1 U10832 ( .B1(n9561), .B2(n9663), .A(n9560), .ZN(n9562) );
  OAI21_X1 U10833 ( .B1(n9796), .B2(n9708), .A(n9562), .ZN(P1_U3268) );
  NAND2_X1 U10834 ( .A1(n9564), .A2(n9563), .ZN(n9565) );
  NAND2_X1 U10835 ( .A1(n9565), .A2(n9571), .ZN(n9566) );
  NAND3_X1 U10836 ( .A1(n9567), .A2(n10140), .A3(n9566), .ZN(n9570) );
  INV_X1 U10837 ( .A(n9568), .ZN(n9569) );
  AND2_X1 U10838 ( .A1(n9570), .A2(n9569), .ZN(n9726) );
  XNOR2_X1 U10839 ( .A(n9572), .B(n9571), .ZN(n9800) );
  INV_X1 U10840 ( .A(n9800), .ZN(n9573) );
  NAND2_X1 U10841 ( .A1(n9573), .A2(n10154), .ZN(n9585) );
  OAI22_X1 U10842 ( .A1(n9576), .A2(n9660), .B1(n9575), .B2(n9663), .ZN(n9583)
         );
  NAND2_X1 U10843 ( .A1(n9578), .A2(n9577), .ZN(n9579) );
  NAND2_X1 U10844 ( .A1(n9579), .A2(n10148), .ZN(n9580) );
  OR2_X1 U10845 ( .A1(n9581), .A2(n9580), .ZN(n9725) );
  NOR2_X1 U10846 ( .A1(n9725), .A2(n9667), .ZN(n9582) );
  AOI211_X1 U10847 ( .C1(n10142), .C2(n9578), .A(n9583), .B(n9582), .ZN(n9584)
         );
  OAI211_X1 U10848 ( .C1(n10130), .C2(n9726), .A(n9585), .B(n9584), .ZN(
        P1_U3269) );
  XNOR2_X1 U10849 ( .A(n9586), .B(n9587), .ZN(n9803) );
  NAND2_X1 U10850 ( .A1(n9607), .A2(n9588), .ZN(n9590) );
  XNOR2_X1 U10851 ( .A(n9590), .B(n9589), .ZN(n9591) );
  NAND2_X1 U10852 ( .A1(n9591), .A2(n10140), .ZN(n9594) );
  INV_X1 U10853 ( .A(n9592), .ZN(n9593) );
  NAND2_X1 U10854 ( .A1(n9594), .A2(n9593), .ZN(n9729) );
  AOI211_X1 U10855 ( .C1(n9731), .C2(n9611), .A(n9693), .B(n5609), .ZN(n9730)
         );
  NAND2_X1 U10856 ( .A1(n9730), .A2(n10153), .ZN(n9597) );
  AOI22_X1 U10857 ( .A1(n9595), .A2(n10143), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10130), .ZN(n9596) );
  OAI211_X1 U10858 ( .C1(n9598), .C2(n9697), .A(n9597), .B(n9596), .ZN(n9599)
         );
  AOI21_X1 U10859 ( .B1(n9663), .B2(n9729), .A(n9599), .ZN(n9600) );
  OAI21_X1 U10860 ( .B1(n9803), .B2(n9708), .A(n9600), .ZN(P1_U3270) );
  NAND2_X1 U10861 ( .A1(n9602), .A2(n9601), .ZN(n9603) );
  XNOR2_X1 U10862 ( .A(n9603), .B(n9604), .ZN(n9808) );
  OAI21_X1 U10863 ( .B1(n9606), .B2(n9605), .A(n9604), .ZN(n9608) );
  NAND3_X1 U10864 ( .A1(n9608), .A2(n10140), .A3(n9607), .ZN(n9610) );
  AND2_X1 U10865 ( .A1(n9610), .A2(n9609), .ZN(n9735) );
  INV_X1 U10866 ( .A(n9735), .ZN(n9618) );
  OAI211_X1 U10867 ( .C1(n9612), .C2(n9628), .A(n10148), .B(n9611), .ZN(n9734)
         );
  INV_X1 U10868 ( .A(n9613), .ZN(n9614) );
  AOI22_X1 U10869 ( .A1(n9614), .A2(n10143), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10130), .ZN(n9616) );
  NAND2_X1 U10870 ( .A1(n9806), .A2(n10142), .ZN(n9615) );
  OAI211_X1 U10871 ( .C1(n9734), .C2(n9667), .A(n9616), .B(n9615), .ZN(n9617)
         );
  AOI21_X1 U10872 ( .B1(n9618), .B2(n9663), .A(n9617), .ZN(n9619) );
  OAI21_X1 U10873 ( .B1(n9808), .B2(n9708), .A(n9619), .ZN(P1_U3271) );
  XNOR2_X1 U10874 ( .A(n4422), .B(n9620), .ZN(n9740) );
  INV_X1 U10875 ( .A(n9740), .ZN(n9635) );
  NAND2_X1 U10876 ( .A1(n9623), .A2(n9622), .ZN(n9625) );
  XNOR2_X1 U10877 ( .A(n9625), .B(n9624), .ZN(n9627) );
  OAI21_X1 U10878 ( .B1(n9627), .B2(n9642), .A(n9626), .ZN(n9738) );
  OAI21_X1 U10879 ( .B1(n9813), .B2(n9646), .A(n10148), .ZN(n9629) );
  NOR2_X1 U10880 ( .A1(n9629), .A2(n9628), .ZN(n9739) );
  NAND2_X1 U10881 ( .A1(n9739), .A2(n10153), .ZN(n9632) );
  AOI22_X1 U10882 ( .A1(n9630), .A2(n10143), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n10130), .ZN(n9631) );
  OAI211_X1 U10883 ( .C1(n9813), .C2(n9697), .A(n9632), .B(n9631), .ZN(n9633)
         );
  AOI21_X1 U10884 ( .B1(n9738), .B2(n9663), .A(n9633), .ZN(n9634) );
  OAI21_X1 U10885 ( .B1(n9635), .B2(n9708), .A(n9634), .ZN(P1_U3272) );
  NAND2_X1 U10886 ( .A1(n9637), .A2(n9636), .ZN(n9638) );
  XOR2_X1 U10887 ( .A(n9639), .B(n9638), .Z(n9819) );
  XNOR2_X1 U10888 ( .A(n9640), .B(n9639), .ZN(n9643) );
  OAI21_X1 U10889 ( .B1(n9643), .B2(n9642), .A(n9641), .ZN(n9745) );
  NAND2_X1 U10890 ( .A1(n9665), .A2(n9816), .ZN(n9644) );
  NAND2_X1 U10891 ( .A1(n9644), .A2(n10148), .ZN(n9645) );
  NOR2_X1 U10892 ( .A1(n9646), .A2(n9645), .ZN(n9744) );
  NAND2_X1 U10893 ( .A1(n9744), .A2(n10153), .ZN(n9649) );
  AOI22_X1 U10894 ( .A1(n9647), .A2(n10143), .B1(P1_REG2_REG_20__SCAN_IN), 
        .B2(n10130), .ZN(n9648) );
  OAI211_X1 U10895 ( .C1(n4808), .C2(n9697), .A(n9649), .B(n9648), .ZN(n9650)
         );
  AOI21_X1 U10896 ( .B1(n9745), .B2(n9663), .A(n9650), .ZN(n9651) );
  OAI21_X1 U10897 ( .B1(n9819), .B2(n9708), .A(n9651), .ZN(P1_U3273) );
  OAI21_X1 U10898 ( .B1(n9657), .B2(n9653), .A(n9652), .ZN(n9656) );
  INV_X1 U10899 ( .A(n9654), .ZN(n9655) );
  AOI21_X1 U10900 ( .B1(n9656), .B2(n10140), .A(n9655), .ZN(n9750) );
  XOR2_X1 U10901 ( .A(n9657), .B(n9658), .Z(n9824) );
  INV_X1 U10902 ( .A(n9824), .ZN(n9659) );
  NAND2_X1 U10903 ( .A1(n9659), .A2(n10154), .ZN(n9671) );
  OAI22_X1 U10904 ( .A1(n9663), .A2(n9662), .B1(n9661), .B2(n9660), .ZN(n9669)
         );
  AOI21_X1 U10905 ( .B1(n9664), .B2(n9822), .A(n9693), .ZN(n9666) );
  NAND2_X1 U10906 ( .A1(n9666), .A2(n9665), .ZN(n9749) );
  NOR2_X1 U10907 ( .A1(n9749), .A2(n9667), .ZN(n9668) );
  AOI211_X1 U10908 ( .C1(n10142), .C2(n9822), .A(n9669), .B(n9668), .ZN(n9670)
         );
  OAI211_X1 U10909 ( .C1(n10130), .C2(n9750), .A(n9671), .B(n9670), .ZN(
        P1_U3274) );
  XNOR2_X1 U10910 ( .A(n9672), .B(n4384), .ZN(n9757) );
  INV_X1 U10911 ( .A(n9673), .ZN(n9675) );
  INV_X1 U10912 ( .A(n9664), .ZN(n9674) );
  AOI211_X1 U10913 ( .C1(n9754), .C2(n9675), .A(n9693), .B(n9674), .ZN(n9753)
         );
  INV_X1 U10914 ( .A(n9676), .ZN(n9677) );
  AOI22_X1 U10915 ( .A1(n10130), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9677), 
        .B2(n10143), .ZN(n9678) );
  OAI21_X1 U10916 ( .B1(n9679), .B2(n9697), .A(n9678), .ZN(n9687) );
  AND2_X1 U10917 ( .A1(n9681), .A2(n9680), .ZN(n9683) );
  OAI21_X1 U10918 ( .B1(n9683), .B2(n4384), .A(n9682), .ZN(n9685) );
  AOI21_X1 U10919 ( .B1(n9685), .B2(n10140), .A(n9684), .ZN(n9756) );
  NOR2_X1 U10920 ( .A1(n9756), .A2(n10130), .ZN(n9686) );
  AOI211_X1 U10921 ( .C1(n9753), .C2(n10153), .A(n9687), .B(n9686), .ZN(n9688)
         );
  OAI21_X1 U10922 ( .B1(n9757), .B2(n9708), .A(n9688), .ZN(P1_U3275) );
  XNOR2_X1 U10923 ( .A(n9689), .B(n9690), .ZN(n9767) );
  INV_X1 U10924 ( .A(n9691), .ZN(n9692) );
  AOI211_X1 U10925 ( .C1(n9764), .C2(n9694), .A(n9693), .B(n9692), .ZN(n9763)
         );
  AOI22_X1 U10926 ( .A1(n10130), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9695), 
        .B2(n10143), .ZN(n9696) );
  OAI21_X1 U10927 ( .B1(n9698), .B2(n9697), .A(n9696), .ZN(n9706) );
  OAI21_X1 U10928 ( .B1(n9701), .B2(n9700), .A(n9699), .ZN(n9704) );
  INV_X1 U10929 ( .A(n9702), .ZN(n9703) );
  AOI21_X1 U10930 ( .B1(n9704), .B2(n10140), .A(n9703), .ZN(n9766) );
  NOR2_X1 U10931 ( .A1(n9766), .A2(n10130), .ZN(n9705) );
  AOI211_X1 U10932 ( .C1(n9763), .C2(n10153), .A(n9706), .B(n9705), .ZN(n9707)
         );
  OAI21_X1 U10933 ( .B1(n9708), .B2(n9767), .A(n9707), .ZN(P1_U3277) );
  INV_X1 U10934 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9711) );
  MUX2_X1 U10935 ( .A(n9711), .B(n9781), .S(n10248), .Z(n9712) );
  OAI21_X1 U10936 ( .B1(n9784), .B2(n9743), .A(n9712), .ZN(P1_U3552) );
  INV_X1 U10937 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9716) );
  NAND2_X1 U10938 ( .A1(n9718), .A2(n9717), .ZN(n9791) );
  MUX2_X1 U10939 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9791), .S(n10248), .Z(
        n9719) );
  OAI211_X1 U10940 ( .C1(n9722), .C2(n10213), .A(n9721), .B(n9720), .ZN(n9793)
         );
  MUX2_X1 U10941 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9793), .S(n10248), .Z(
        n9723) );
  INV_X1 U10942 ( .A(n9723), .ZN(n9724) );
  OAI21_X1 U10943 ( .B1(n9796), .B2(n9773), .A(n9724), .ZN(P1_U3547) );
  NAND2_X1 U10944 ( .A1(n9726), .A2(n9725), .ZN(n9797) );
  MUX2_X1 U10945 ( .A(n9797), .B(P1_REG1_REG_24__SCAN_IN), .S(n10245), .Z(
        n9727) );
  AOI21_X1 U10946 ( .B1(n9771), .B2(n9578), .A(n9727), .ZN(n9728) );
  OAI21_X1 U10947 ( .B1(n9800), .B2(n9773), .A(n9728), .ZN(P1_U3546) );
  INV_X1 U10948 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9732) );
  AOI211_X1 U10949 ( .C1(n10223), .C2(n9731), .A(n9730), .B(n9729), .ZN(n9801)
         );
  MUX2_X1 U10950 ( .A(n9732), .B(n9801), .S(n10248), .Z(n9733) );
  OAI21_X1 U10951 ( .B1(n9803), .B2(n9773), .A(n9733), .ZN(P1_U3545) );
  NAND2_X1 U10952 ( .A1(n9735), .A2(n9734), .ZN(n9804) );
  MUX2_X1 U10953 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9804), .S(n10248), .Z(
        n9736) );
  AOI21_X1 U10954 ( .B1(n9771), .B2(n9806), .A(n9736), .ZN(n9737) );
  OAI21_X1 U10955 ( .B1(n9773), .B2(n9808), .A(n9737), .ZN(P1_U3544) );
  INV_X1 U10956 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9741) );
  AOI211_X1 U10957 ( .C1(n9740), .C2(n10221), .A(n9739), .B(n9738), .ZN(n9809)
         );
  MUX2_X1 U10958 ( .A(n9741), .B(n9809), .S(n10248), .Z(n9742) );
  OAI21_X1 U10959 ( .B1(n9813), .B2(n9743), .A(n9742), .ZN(P1_U3543) );
  INV_X1 U10960 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9746) );
  NOR2_X1 U10961 ( .A1(n9745), .A2(n9744), .ZN(n9814) );
  MUX2_X1 U10962 ( .A(n9746), .B(n9814), .S(n10248), .Z(n9748) );
  NAND2_X1 U10963 ( .A1(n9816), .A2(n9771), .ZN(n9747) );
  OAI211_X1 U10964 ( .C1(n9819), .C2(n9773), .A(n9748), .B(n9747), .ZN(
        P1_U3542) );
  NAND2_X1 U10965 ( .A1(n9750), .A2(n9749), .ZN(n9820) );
  MUX2_X1 U10966 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9820), .S(n10248), .Z(
        n9751) );
  AOI21_X1 U10967 ( .B1(n9771), .B2(n9822), .A(n9751), .ZN(n9752) );
  OAI21_X1 U10968 ( .B1(n9773), .B2(n9824), .A(n9752), .ZN(P1_U3541) );
  AOI21_X1 U10969 ( .B1(n10223), .B2(n9754), .A(n9753), .ZN(n9755) );
  OAI211_X1 U10970 ( .C1(n9757), .C2(n10195), .A(n9756), .B(n9755), .ZN(n9825)
         );
  MUX2_X1 U10971 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9825), .S(n10248), .Z(
        P1_U3540) );
  NOR2_X1 U10972 ( .A1(n9759), .A2(n9758), .ZN(n9826) );
  MUX2_X1 U10973 ( .A(n9760), .B(n9826), .S(n10248), .Z(n9762) );
  NAND2_X1 U10974 ( .A1(n9828), .A2(n9771), .ZN(n9761) );
  OAI211_X1 U10975 ( .C1(n9773), .C2(n9831), .A(n9762), .B(n9761), .ZN(
        P1_U3539) );
  AOI21_X1 U10976 ( .B1(n10223), .B2(n9764), .A(n9763), .ZN(n9765) );
  OAI211_X1 U10977 ( .C1(n9767), .C2(n10195), .A(n9766), .B(n9765), .ZN(n9832)
         );
  MUX2_X1 U10978 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9832), .S(n10248), .Z(
        P1_U3538) );
  NAND2_X1 U10979 ( .A1(n9769), .A2(n9768), .ZN(n9833) );
  MUX2_X1 U10980 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9833), .S(n10248), .Z(
        n9770) );
  AOI21_X1 U10981 ( .B1(n9771), .B2(n9835), .A(n9770), .ZN(n9772) );
  OAI21_X1 U10982 ( .B1(n9839), .B2(n9773), .A(n9772), .ZN(P1_U3537) );
  INV_X1 U10983 ( .A(n9774), .ZN(n9780) );
  AOI21_X1 U10984 ( .B1(n10223), .B2(n9776), .A(n9775), .ZN(n9777) );
  OAI211_X1 U10985 ( .C1(n9780), .C2(n9779), .A(n9778), .B(n9777), .ZN(n9840)
         );
  MUX2_X1 U10986 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9840), .S(n10248), .Z(
        P1_U3536) );
  INV_X1 U10987 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9782) );
  MUX2_X1 U10988 ( .A(n9782), .B(n9781), .S(n10232), .Z(n9783) );
  OAI21_X1 U10989 ( .B1(n9784), .B2(n9812), .A(n9783), .ZN(P1_U3520) );
  INV_X1 U10990 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9786) );
  OAI21_X1 U10991 ( .B1(n9788), .B2(n9838), .A(n9787), .ZN(P1_U3517) );
  MUX2_X1 U10992 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9791), .S(n10232), .Z(
        n9792) );
  INV_X1 U10993 ( .A(n9793), .ZN(n9794) );
  MUX2_X1 U10994 ( .A(n9915), .B(n9794), .S(n10232), .Z(n9795) );
  OAI21_X1 U10995 ( .B1(n9796), .B2(n9838), .A(n9795), .ZN(P1_U3515) );
  MUX2_X1 U10996 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9797), .S(n10232), .Z(
        n9798) );
  AOI21_X1 U10997 ( .B1(n9836), .B2(n9578), .A(n9798), .ZN(n9799) );
  OAI21_X1 U10998 ( .B1(n9800), .B2(n9838), .A(n9799), .ZN(P1_U3514) );
  MUX2_X1 U10999 ( .A(n9940), .B(n9801), .S(n10232), .Z(n9802) );
  OAI21_X1 U11000 ( .B1(n9803), .B2(n9838), .A(n9802), .ZN(P1_U3513) );
  MUX2_X1 U11001 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9804), .S(n10232), .Z(
        n9805) );
  AOI21_X1 U11002 ( .B1(n9836), .B2(n9806), .A(n9805), .ZN(n9807) );
  OAI21_X1 U11003 ( .B1(n9838), .B2(n9808), .A(n9807), .ZN(P1_U3512) );
  INV_X1 U11004 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9810) );
  MUX2_X1 U11005 ( .A(n9810), .B(n9809), .S(n10232), .Z(n9811) );
  OAI21_X1 U11006 ( .B1(n9813), .B2(n9812), .A(n9811), .ZN(P1_U3511) );
  INV_X1 U11007 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9815) );
  MUX2_X1 U11008 ( .A(n9815), .B(n9814), .S(n10232), .Z(n9818) );
  NAND2_X1 U11009 ( .A1(n9816), .A2(n9836), .ZN(n9817) );
  OAI211_X1 U11010 ( .C1(n9819), .C2(n9838), .A(n9818), .B(n9817), .ZN(
        P1_U3510) );
  MUX2_X1 U11011 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9820), .S(n10232), .Z(
        n9821) );
  AOI21_X1 U11012 ( .B1(n9836), .B2(n9822), .A(n9821), .ZN(n9823) );
  OAI21_X1 U11013 ( .B1(n9838), .B2(n9824), .A(n9823), .ZN(P1_U3509) );
  MUX2_X1 U11014 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9825), .S(n10232), .Z(
        P1_U3507) );
  INV_X1 U11015 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9827) );
  MUX2_X1 U11016 ( .A(n9827), .B(n9826), .S(n10232), .Z(n9830) );
  NAND2_X1 U11017 ( .A1(n9828), .A2(n9836), .ZN(n9829) );
  OAI211_X1 U11018 ( .C1(n9831), .C2(n9838), .A(n9830), .B(n9829), .ZN(
        P1_U3504) );
  MUX2_X1 U11019 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9832), .S(n10232), .Z(
        P1_U3501) );
  MUX2_X1 U11020 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9833), .S(n10232), .Z(
        n9834) );
  AOI21_X1 U11021 ( .B1(n9836), .B2(n9835), .A(n9834), .ZN(n9837) );
  OAI21_X1 U11022 ( .B1(n9839), .B2(n9838), .A(n9837), .ZN(P1_U3498) );
  MUX2_X1 U11023 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9840), .S(n10232), .Z(
        n9994) );
  AOI22_X1 U11024 ( .A1(n5147), .A2(keyinput6), .B1(keyinput29), .B2(n9842), 
        .ZN(n9841) );
  OAI221_X1 U11025 ( .B1(n5147), .B2(keyinput6), .C1(n9842), .C2(keyinput29), 
        .A(n9841), .ZN(n9852) );
  INV_X1 U11026 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9844) );
  INV_X1 U11027 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10056) );
  AOI22_X1 U11028 ( .A1(n9844), .A2(keyinput42), .B1(keyinput58), .B2(n10056), 
        .ZN(n9843) );
  OAI221_X1 U11029 ( .B1(n9844), .B2(keyinput42), .C1(n10056), .C2(keyinput58), 
        .A(n9843), .ZN(n9851) );
  AOI22_X1 U11030 ( .A1(n9928), .A2(keyinput30), .B1(keyinput37), .B2(n9846), 
        .ZN(n9845) );
  OAI221_X1 U11031 ( .B1(n9928), .B2(keyinput30), .C1(n9846), .C2(keyinput37), 
        .A(n9845), .ZN(n9850) );
  INV_X1 U11032 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10158) );
  AOI22_X1 U11033 ( .A1(n10158), .A2(keyinput8), .B1(keyinput61), .B2(n9848), 
        .ZN(n9847) );
  OAI221_X1 U11034 ( .B1(n10158), .B2(keyinput8), .C1(n9848), .C2(keyinput61), 
        .A(n9847), .ZN(n9849) );
  NOR4_X1 U11035 ( .A1(n9852), .A2(n9851), .A3(n9850), .A4(n9849), .ZN(n9992)
         );
  AOI22_X1 U11036 ( .A1(n9854), .A2(keyinput32), .B1(keyinput41), .B2(n6221), 
        .ZN(n9853) );
  OAI221_X1 U11037 ( .B1(n9854), .B2(keyinput32), .C1(n6221), .C2(keyinput41), 
        .A(n9853), .ZN(n9865) );
  INV_X1 U11038 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9857) );
  AOI22_X1 U11039 ( .A1(n9857), .A2(keyinput56), .B1(keyinput45), .B2(n9856), 
        .ZN(n9855) );
  OAI221_X1 U11040 ( .B1(n9857), .B2(keyinput56), .C1(n9856), .C2(keyinput45), 
        .A(n9855), .ZN(n9864) );
  INV_X1 U11041 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9860) );
  AOI22_X1 U11042 ( .A1(n9860), .A2(keyinput23), .B1(keyinput16), .B2(n9859), 
        .ZN(n9858) );
  OAI221_X1 U11043 ( .B1(n9860), .B2(keyinput23), .C1(n9859), .C2(keyinput16), 
        .A(n9858), .ZN(n9863) );
  INV_X1 U11044 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9909) );
  AOI22_X1 U11045 ( .A1(n9908), .A2(keyinput46), .B1(n9909), .B2(keyinput24), 
        .ZN(n9861) );
  OAI221_X1 U11046 ( .B1(n9908), .B2(keyinput46), .C1(n9909), .C2(keyinput24), 
        .A(n9861), .ZN(n9862) );
  NOR4_X1 U11047 ( .A1(n9865), .A2(n9864), .A3(n9863), .A4(n9862), .ZN(n9991)
         );
  AOI22_X1 U11048 ( .A1(n9867), .A2(keyinput35), .B1(n9904), .B2(keyinput38), 
        .ZN(n9866) );
  OAI221_X1 U11049 ( .B1(n9867), .B2(keyinput35), .C1(n9904), .C2(keyinput38), 
        .A(n9866), .ZN(n9873) );
  XNOR2_X1 U11050 ( .A(P1_REG3_REG_0__SCAN_IN), .B(keyinput10), .ZN(n9871) );
  XNOR2_X1 U11051 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(keyinput0), .ZN(n9870) );
  XNOR2_X1 U11052 ( .A(P1_REG3_REG_10__SCAN_IN), .B(keyinput44), .ZN(n9869) );
  XNOR2_X1 U11053 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput48), .ZN(n9868) );
  NAND4_X1 U11054 ( .A1(n9871), .A2(n9870), .A3(n9869), .A4(n9868), .ZN(n9872)
         );
  NOR2_X1 U11055 ( .A1(n9873), .A2(n9872), .ZN(n9887) );
  XNOR2_X1 U11056 ( .A(keyinput21), .B(n9874), .ZN(n9876) );
  XNOR2_X1 U11057 ( .A(keyinput27), .B(n7462), .ZN(n9875) );
  NOR2_X1 U11058 ( .A1(n9876), .A2(n9875), .ZN(n9886) );
  AOI22_X1 U11059 ( .A1(n9914), .A2(keyinput36), .B1(n9878), .B2(keyinput60), 
        .ZN(n9877) );
  OAI221_X1 U11060 ( .B1(n9914), .B2(keyinput36), .C1(n9878), .C2(keyinput60), 
        .A(n9877), .ZN(n9879) );
  INV_X1 U11061 ( .A(n9879), .ZN(n9885) );
  INV_X1 U11062 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9881) );
  AOI22_X1 U11063 ( .A1(n9882), .A2(keyinput15), .B1(n9881), .B2(keyinput34), 
        .ZN(n9880) );
  OAI221_X1 U11064 ( .B1(n9882), .B2(keyinput15), .C1(n9881), .C2(keyinput34), 
        .A(n9880), .ZN(n9883) );
  INV_X1 U11065 ( .A(n9883), .ZN(n9884) );
  AND4_X1 U11066 ( .A1(n9887), .A2(n9886), .A3(n9885), .A4(n9884), .ZN(n9938)
         );
  INV_X1 U11067 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10204) );
  AOI22_X1 U11068 ( .A1(n10204), .A2(keyinput26), .B1(keyinput28), .B2(n9889), 
        .ZN(n9888) );
  OAI221_X1 U11069 ( .B1(n10204), .B2(keyinput26), .C1(n9889), .C2(keyinput28), 
        .A(n9888), .ZN(n9892) );
  INV_X1 U11070 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9912) );
  AOI22_X1 U11071 ( .A1(n5332), .A2(keyinput40), .B1(keyinput18), .B2(n9912), 
        .ZN(n9890) );
  OAI221_X1 U11072 ( .B1(n5332), .B2(keyinput40), .C1(n9912), .C2(keyinput18), 
        .A(n9890), .ZN(n9891) );
  NOR2_X1 U11073 ( .A1(n9892), .A2(n9891), .ZN(n9937) );
  INV_X1 U11074 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10172) );
  AOI22_X1 U11075 ( .A1(n9894), .A2(keyinput11), .B1(keyinput12), .B2(n10172), 
        .ZN(n9893) );
  OAI221_X1 U11076 ( .B1(n9894), .B2(keyinput11), .C1(n10172), .C2(keyinput12), 
        .A(n9893), .ZN(n9898) );
  INV_X1 U11077 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9896) );
  AOI22_X1 U11078 ( .A1(n5701), .A2(keyinput22), .B1(keyinput51), .B2(n9896), 
        .ZN(n9895) );
  OAI221_X1 U11079 ( .B1(n5701), .B2(keyinput22), .C1(n9896), .C2(keyinput51), 
        .A(n9895), .ZN(n9897) );
  NOR2_X1 U11080 ( .A1(n9898), .A2(n9897), .ZN(n9936) );
  NOR4_X1 U11081 ( .A1(P1_REG1_REG_13__SCAN_IN), .A2(P2_REG3_REG_23__SCAN_IN), 
        .A3(P2_D_REG_11__SCAN_IN), .A4(P2_ADDR_REG_13__SCAN_IN), .ZN(n9934) );
  NAND4_X1 U11082 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), 
        .A3(P2_D_REG_14__SCAN_IN), .A4(n10172), .ZN(n9902) );
  NAND3_X1 U11083 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P2_REG3_REG_8__SCAN_IN), 
        .A3(P1_ADDR_REG_5__SCAN_IN), .ZN(n9901) );
  INV_X1 U11084 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9899) );
  NAND4_X1 U11085 ( .A1(n9899), .A2(n9940), .A3(P1_REG0_REG_31__SCAN_IN), .A4(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n9900) );
  NOR3_X1 U11086 ( .A1(n9902), .A2(n9901), .A3(n9900), .ZN(n9933) );
  NAND4_X1 U11087 ( .A1(n9904), .A2(n9903), .A3(n9952), .A4(
        P2_REG3_REG_24__SCAN_IN), .ZN(n9906) );
  NAND4_X1 U11088 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), 
        .A3(P1_REG3_REG_4__SCAN_IN), .A4(P1_B_REG_SCAN_IN), .ZN(n9905) );
  NOR2_X1 U11089 ( .A1(n9906), .A2(n9905), .ZN(n9925) );
  NAND4_X1 U11090 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(P1_DATAO_REG_8__SCAN_IN), .A3(P1_DATAO_REG_4__SCAN_IN), .A4(P2_REG2_REG_29__SCAN_IN), .ZN(n9907) );
  NOR2_X1 U11091 ( .A1(n5701), .A2(n9907), .ZN(n9913) );
  NOR4_X1 U11092 ( .A1(P1_REG1_REG_22__SCAN_IN), .A2(P1_REG2_REG_18__SCAN_IN), 
        .A3(P1_REG2_REG_11__SCAN_IN), .A4(P2_IR_REG_11__SCAN_IN), .ZN(n9911)
         );
  NOR4_X1 U11093 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(SI_31_), .A3(n9909), 
        .A4(n9908), .ZN(n9910) );
  NAND4_X1 U11094 ( .A1(n9913), .A2(n9912), .A3(n9911), .A4(n9910), .ZN(n9920)
         );
  AND4_X1 U11095 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(SI_23_), .A3(
        P2_REG0_REG_17__SCAN_IN), .A4(n9914), .ZN(n9918) );
  AND4_X1 U11096 ( .A1(SI_0_), .A2(P1_REG0_REG_6__SCAN_IN), .A3(
        P1_REG3_REG_0__SCAN_IN), .A4(n9948), .ZN(n9917) );
  AND4_X1 U11097 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_REG1_REG_16__SCAN_IN), 
        .A3(P1_REG2_REG_16__SCAN_IN), .A4(n9915), .ZN(n9916) );
  NAND4_X1 U11098 ( .A1(n9918), .A2(n9917), .A3(n9916), .A4(n5332), .ZN(n9919)
         );
  NOR2_X1 U11099 ( .A1(n9920), .A2(n9919), .ZN(n9921) );
  AND4_X1 U11100 ( .A1(n9923), .A2(n9922), .A3(P2_IR_REG_26__SCAN_IN), .A4(
        n9921), .ZN(n9924) );
  NAND4_X1 U11101 ( .A1(n9925), .A2(P1_ADDR_REG_3__SCAN_IN), .A3(n9924), .A4(
        n9896), .ZN(n9927) );
  NAND4_X1 U11102 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(P2_REG0_REG_6__SCAN_IN), 
        .A3(n5147), .A4(n10056), .ZN(n9926) );
  NOR2_X1 U11103 ( .A1(n9927), .A2(n9926), .ZN(n9932) );
  NOR3_X1 U11104 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .A3(n9928), .ZN(n9929) );
  AND2_X1 U11105 ( .A1(n9930), .A2(n9929), .ZN(n9931) );
  NAND4_X1 U11106 ( .A1(n9934), .A2(n9933), .A3(n9932), .A4(n9931), .ZN(n9935)
         );
  AND4_X1 U11107 ( .A1(n9938), .A2(n9937), .A3(n9936), .A4(n9935), .ZN(n9990)
         );
  AOI22_X1 U11108 ( .A1(n9941), .A2(keyinput52), .B1(n9940), .B2(keyinput63), 
        .ZN(n9939) );
  OAI221_X1 U11109 ( .B1(n9941), .B2(keyinput52), .C1(n9940), .C2(keyinput63), 
        .A(n9939), .ZN(n9946) );
  AOI22_X1 U11110 ( .A1(n9944), .A2(keyinput4), .B1(keyinput1), .B2(n9943), 
        .ZN(n9942) );
  OAI221_X1 U11111 ( .B1(n9944), .B2(keyinput4), .C1(n9943), .C2(keyinput1), 
        .A(n9942), .ZN(n9945) );
  NOR2_X1 U11112 ( .A1(n9946), .A2(n9945), .ZN(n9978) );
  INV_X1 U11113 ( .A(SI_0_), .ZN(n9949) );
  AOI22_X1 U11114 ( .A1(n9949), .A2(keyinput57), .B1(n9948), .B2(keyinput47), 
        .ZN(n9947) );
  OAI221_X1 U11115 ( .B1(n9949), .B2(keyinput57), .C1(n9948), .C2(keyinput47), 
        .A(n9947), .ZN(n9954) );
  INV_X1 U11116 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9951) );
  AOI22_X1 U11117 ( .A1(n9952), .A2(keyinput49), .B1(n9951), .B2(keyinput50), 
        .ZN(n9950) );
  OAI221_X1 U11118 ( .B1(n9952), .B2(keyinput49), .C1(n9951), .C2(keyinput50), 
        .A(n9950), .ZN(n9953) );
  NOR2_X1 U11119 ( .A1(n9954), .A2(n9953), .ZN(n9977) );
  XNOR2_X1 U11120 ( .A(SI_6_), .B(keyinput54), .ZN(n9958) );
  XNOR2_X1 U11121 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput14), .ZN(n9957) );
  XNOR2_X1 U11122 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput9), .ZN(n9956) );
  XNOR2_X1 U11123 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput31), .ZN(n9955)
         );
  NAND4_X1 U11124 ( .A1(n9958), .A2(n9957), .A3(n9956), .A4(n9955), .ZN(n9964)
         );
  XNOR2_X1 U11125 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput5), .ZN(n9962) );
  XNOR2_X1 U11126 ( .A(P1_REG0_REG_12__SCAN_IN), .B(keyinput59), .ZN(n9961) );
  XNOR2_X1 U11127 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(keyinput25), .ZN(n9960) );
  XNOR2_X1 U11128 ( .A(P1_REG3_REG_4__SCAN_IN), .B(keyinput3), .ZN(n9959) );
  NAND4_X1 U11129 ( .A1(n9962), .A2(n9961), .A3(n9960), .A4(n9959), .ZN(n9963)
         );
  NOR2_X1 U11130 ( .A1(n9964), .A2(n9963), .ZN(n9976) );
  XNOR2_X1 U11131 ( .A(P1_B_REG_SCAN_IN), .B(keyinput19), .ZN(n9968) );
  XNOR2_X1 U11132 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput13), .ZN(n9967) );
  XNOR2_X1 U11133 ( .A(P2_IR_REG_5__SCAN_IN), .B(keyinput43), .ZN(n9966) );
  XNOR2_X1 U11134 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput62), .ZN(n9965) );
  NAND4_X1 U11135 ( .A1(n9968), .A2(n9967), .A3(n9966), .A4(n9965), .ZN(n9974)
         );
  XNOR2_X1 U11136 ( .A(P2_REG2_REG_29__SCAN_IN), .B(keyinput55), .ZN(n9972) );
  XNOR2_X1 U11137 ( .A(P2_IR_REG_26__SCAN_IN), .B(keyinput20), .ZN(n9971) );
  XNOR2_X1 U11138 ( .A(P1_REG0_REG_25__SCAN_IN), .B(keyinput2), .ZN(n9970) );
  XNOR2_X1 U11139 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput7), .ZN(n9969) );
  NAND4_X1 U11140 ( .A1(n9972), .A2(n9971), .A3(n9970), .A4(n9969), .ZN(n9973)
         );
  NOR2_X1 U11141 ( .A1(n9974), .A2(n9973), .ZN(n9975) );
  NAND4_X1 U11142 ( .A1(n9978), .A2(n9977), .A3(n9976), .A4(n9975), .ZN(n9988)
         );
  INV_X1 U11143 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10162) );
  INV_X1 U11144 ( .A(keyinput53), .ZN(n9979) );
  XNOR2_X1 U11145 ( .A(n10162), .B(n9979), .ZN(n9986) );
  INV_X1 U11146 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10161) );
  INV_X1 U11147 ( .A(keyinput33), .ZN(n9980) );
  XNOR2_X1 U11148 ( .A(n10161), .B(n9980), .ZN(n9985) );
  INV_X1 U11149 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10157) );
  INV_X1 U11150 ( .A(keyinput39), .ZN(n9981) );
  XNOR2_X1 U11151 ( .A(n10157), .B(n9981), .ZN(n9984) );
  INV_X1 U11152 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10159) );
  INV_X1 U11153 ( .A(keyinput17), .ZN(n9982) );
  XNOR2_X1 U11154 ( .A(n10159), .B(n9982), .ZN(n9983) );
  NAND4_X1 U11155 ( .A1(n9986), .A2(n9985), .A3(n9984), .A4(n9983), .ZN(n9987)
         );
  NOR2_X1 U11156 ( .A1(n9988), .A2(n9987), .ZN(n9989) );
  NAND4_X1 U11157 ( .A1(n9992), .A2(n9991), .A3(n9990), .A4(n9989), .ZN(n9993)
         );
  XNOR2_X1 U11158 ( .A(n9994), .B(n9993), .ZN(P1_U3495) );
  MUX2_X1 U11159 ( .A(P1_D_REG_1__SCAN_IN), .B(n9997), .S(n10163), .Z(P1_U3440) );
  MUX2_X1 U11160 ( .A(P1_D_REG_0__SCAN_IN), .B(n9998), .S(n10163), .Z(P1_U3439) );
  OAI222_X1 U11161 ( .A1(n10005), .A2(n10001), .B1(n10008), .B2(n10000), .C1(
        n9999), .C2(P1_U3086), .ZN(P1_U3326) );
  OAI222_X1 U11162 ( .A1(n10005), .A2(n10004), .B1(n10008), .B2(n10003), .C1(
        n10002), .C2(P1_U3086), .ZN(P1_U3328) );
  OAI222_X1 U11163 ( .A1(n10009), .A2(P1_U3086), .B1(n10008), .B2(n10007), 
        .C1(n10006), .C2(n10005), .ZN(P1_U3330) );
  MUX2_X1 U11164 ( .A(n10010), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U11165 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11166 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  OAI21_X1 U11167 ( .B1(n10012), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10011), .ZN(
        n10013) );
  XOR2_X1 U11168 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10013), .Z(n10017) );
  AOI22_X1 U11169 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n10014), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n10015) );
  OAI21_X1 U11170 ( .B1(n10017), .B2(n10016), .A(n10015), .ZN(P1_U3243) );
  INV_X1 U11171 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10029) );
  AOI211_X1 U11172 ( .C1(n10020), .C2(n10019), .A(n10047), .B(n10018), .ZN(
        n10025) );
  AOI211_X1 U11173 ( .C1(n10023), .C2(n10022), .A(n10030), .B(n10021), .ZN(
        n10024) );
  AOI211_X1 U11174 ( .C1(n10083), .C2(n10026), .A(n10025), .B(n10024), .ZN(
        n10028) );
  OAI211_X1 U11175 ( .C1(n10089), .C2(n10029), .A(n10028), .B(n10027), .ZN(
        P1_U3257) );
  INV_X1 U11176 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10042) );
  AOI211_X1 U11177 ( .C1(n10033), .C2(n10032), .A(n10031), .B(n10030), .ZN(
        n10038) );
  AOI211_X1 U11178 ( .C1(n10036), .C2(n10035), .A(n10034), .B(n10047), .ZN(
        n10037) );
  AOI211_X1 U11179 ( .C1(n10083), .C2(n10039), .A(n10038), .B(n10037), .ZN(
        n10041) );
  OAI211_X1 U11180 ( .C1(n10089), .C2(n10042), .A(n10041), .B(n10040), .ZN(
        P1_U3258) );
  OAI21_X1 U11181 ( .B1(n10045), .B2(n10044), .A(n10043), .ZN(n10053) );
  NOR2_X1 U11182 ( .A1(n10069), .A2(n10046), .ZN(n10052) );
  AOI211_X1 U11183 ( .C1(n10050), .C2(n10049), .A(n10048), .B(n10047), .ZN(
        n10051) );
  AOI211_X1 U11184 ( .C1(n10081), .C2(n10053), .A(n10052), .B(n10051), .ZN(
        n10055) );
  OAI211_X1 U11185 ( .C1(n10056), .C2(n10089), .A(n10055), .B(n10054), .ZN(
        P1_U3259) );
  INV_X1 U11186 ( .A(n10057), .ZN(n10068) );
  OAI21_X1 U11187 ( .B1(n10060), .B2(n10059), .A(n10058), .ZN(n10061) );
  NAND2_X1 U11188 ( .A1(n10075), .A2(n10061), .ZN(n10067) );
  OAI21_X1 U11189 ( .B1(n10064), .B2(n10063), .A(n10062), .ZN(n10065) );
  NAND2_X1 U11190 ( .A1(n10081), .A2(n10065), .ZN(n10066) );
  OAI211_X1 U11191 ( .C1(n10069), .C2(n10068), .A(n10067), .B(n10066), .ZN(
        n10070) );
  INV_X1 U11192 ( .A(n10070), .ZN(n10072) );
  OAI211_X1 U11193 ( .C1(n10089), .C2(n10073), .A(n10072), .B(n10071), .ZN(
        P1_U3260) );
  OAI211_X1 U11194 ( .C1(n10076), .C2(n4339), .A(n10075), .B(n10074), .ZN(
        n10086) );
  NAND2_X1 U11195 ( .A1(n10078), .A2(n10077), .ZN(n10079) );
  NAND3_X1 U11196 ( .A1(n10081), .A2(n10080), .A3(n10079), .ZN(n10085) );
  NAND2_X1 U11197 ( .A1(n10083), .A2(n10082), .ZN(n10084) );
  AND3_X1 U11198 ( .A1(n10086), .A2(n10085), .A3(n10084), .ZN(n10088) );
  NAND2_X1 U11199 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n10087)
         );
  OAI211_X1 U11200 ( .C1(n10089), .C2(n10330), .A(n10088), .B(n10087), .ZN(
        P1_U3261) );
  INV_X1 U11201 ( .A(n10090), .ZN(n10091) );
  OR2_X1 U11202 ( .A1(n10092), .A2(n10091), .ZN(n10094) );
  XNOR2_X1 U11203 ( .A(n10093), .B(n10094), .ZN(n10098) );
  XNOR2_X1 U11204 ( .A(n7277), .B(n10094), .ZN(n10100) );
  NOR2_X1 U11205 ( .A1(n10100), .A2(n10095), .ZN(n10096) );
  AOI211_X1 U11206 ( .C1(n10140), .C2(n10098), .A(n10097), .B(n10096), .ZN(
        n10215) );
  AOI222_X1 U11207 ( .A1(n10101), .A2(n10142), .B1(P1_REG2_REG_8__SCAN_IN), 
        .B2(n10130), .C1(n10143), .C2(n10099), .ZN(n10107) );
  INV_X1 U11208 ( .A(n10100), .ZN(n10218) );
  INV_X1 U11209 ( .A(n7318), .ZN(n10103) );
  INV_X1 U11210 ( .A(n10101), .ZN(n10214) );
  OAI211_X1 U11211 ( .C1(n10103), .C2(n10214), .A(n10148), .B(n10102), .ZN(
        n10212) );
  INV_X1 U11212 ( .A(n10212), .ZN(n10104) );
  AOI22_X1 U11213 ( .A1(n10218), .A2(n10105), .B1(n10153), .B2(n10104), .ZN(
        n10106) );
  OAI211_X1 U11214 ( .C1(n10130), .C2(n10215), .A(n10107), .B(n10106), .ZN(
        P1_U3285) );
  XOR2_X1 U11215 ( .A(n10108), .B(n10114), .Z(n10110) );
  AOI21_X1 U11216 ( .B1(n10110), .B2(n10140), .A(n10109), .ZN(n10200) );
  AOI222_X1 U11217 ( .A1(n10116), .A2(n10142), .B1(n10111), .B2(n10143), .C1(
        P1_REG2_REG_6__SCAN_IN), .C2(n10130), .ZN(n10123) );
  NAND2_X1 U11218 ( .A1(n10113), .A2(n10112), .ZN(n10115) );
  XNOR2_X1 U11219 ( .A(n10114), .B(n10115), .ZN(n10203) );
  NAND2_X1 U11220 ( .A1(n10117), .A2(n10116), .ZN(n10118) );
  NAND2_X1 U11221 ( .A1(n10118), .A2(n10148), .ZN(n10120) );
  OR2_X1 U11222 ( .A1(n10120), .A2(n10119), .ZN(n10199) );
  INV_X1 U11223 ( .A(n10199), .ZN(n10121) );
  AOI22_X1 U11224 ( .A1(n10203), .A2(n10154), .B1(n10153), .B2(n10121), .ZN(
        n10122) );
  OAI211_X1 U11225 ( .C1(n10130), .C2(n10200), .A(n10123), .B(n10122), .ZN(
        P1_U3287) );
  NAND2_X1 U11226 ( .A1(n10125), .A2(n10124), .ZN(n10126) );
  XNOR2_X1 U11227 ( .A(n10126), .B(n10133), .ZN(n10128) );
  AOI21_X1 U11228 ( .B1(n10128), .B2(n10140), .A(n10127), .ZN(n10186) );
  AOI222_X1 U11229 ( .A1(n10131), .A2(n10142), .B1(P1_REG2_REG_4__SCAN_IN), 
        .B2(n10130), .C1(n10129), .C2(n10143), .ZN(n10136) );
  XNOR2_X1 U11230 ( .A(n10132), .B(n10133), .ZN(n10189) );
  OAI211_X1 U11231 ( .C1(n4803), .C2(n10185), .A(n10148), .B(n4334), .ZN(
        n10184) );
  INV_X1 U11232 ( .A(n10184), .ZN(n10134) );
  AOI22_X1 U11233 ( .A1(n10189), .A2(n10154), .B1(n10153), .B2(n10134), .ZN(
        n10135) );
  OAI211_X1 U11234 ( .C1(n10130), .C2(n10186), .A(n10136), .B(n10135), .ZN(
        P1_U3289) );
  XNOR2_X1 U11235 ( .A(n10138), .B(n10137), .ZN(n10141) );
  AOI21_X1 U11236 ( .B1(n10141), .B2(n10140), .A(n10139), .ZN(n10174) );
  AOI222_X1 U11237 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n10130), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10143), .C1(n10147), .C2(n10142), .ZN(
        n10156) );
  XNOR2_X1 U11238 ( .A(n10145), .B(n10144), .ZN(n10177) );
  NAND2_X1 U11239 ( .A1(n10147), .A2(n10146), .ZN(n10149) );
  NAND2_X1 U11240 ( .A1(n10149), .A2(n10148), .ZN(n10150) );
  OR2_X1 U11241 ( .A1(n10151), .A2(n10150), .ZN(n10173) );
  INV_X1 U11242 ( .A(n10173), .ZN(n10152) );
  AOI22_X1 U11243 ( .A1(n10177), .A2(n10154), .B1(n10153), .B2(n10152), .ZN(
        n10155) );
  OAI211_X1 U11244 ( .C1(n10130), .C2(n10174), .A(n10156), .B(n10155), .ZN(
        P1_U3291) );
  AND2_X1 U11245 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10160), .ZN(P1_U3294) );
  AND2_X1 U11246 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10160), .ZN(P1_U3295) );
  AND2_X1 U11247 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10160), .ZN(P1_U3296) );
  NOR2_X1 U11248 ( .A1(n10163), .A2(n10157), .ZN(P1_U3297) );
  AND2_X1 U11249 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10160), .ZN(P1_U3298) );
  AND2_X1 U11250 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10160), .ZN(P1_U3299) );
  AND2_X1 U11251 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10160), .ZN(P1_U3300) );
  AND2_X1 U11252 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10160), .ZN(P1_U3301) );
  NOR2_X1 U11253 ( .A1(n10163), .A2(n10158), .ZN(P1_U3302) );
  AND2_X1 U11254 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10160), .ZN(P1_U3303) );
  AND2_X1 U11255 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10160), .ZN(P1_U3304) );
  AND2_X1 U11256 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10160), .ZN(P1_U3305) );
  AND2_X1 U11257 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10160), .ZN(P1_U3306) );
  AND2_X1 U11258 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10160), .ZN(P1_U3307) );
  NOR2_X1 U11259 ( .A1(n10163), .A2(n10159), .ZN(P1_U3308) );
  AND2_X1 U11260 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10160), .ZN(P1_U3309) );
  AND2_X1 U11261 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10160), .ZN(P1_U3310) );
  AND2_X1 U11262 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10160), .ZN(P1_U3311) );
  AND2_X1 U11263 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10160), .ZN(P1_U3312) );
  AND2_X1 U11264 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10160), .ZN(P1_U3313) );
  AND2_X1 U11265 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10160), .ZN(P1_U3314) );
  AND2_X1 U11266 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10160), .ZN(P1_U3315) );
  AND2_X1 U11267 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10160), .ZN(P1_U3316) );
  AND2_X1 U11268 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10160), .ZN(P1_U3317) );
  AND2_X1 U11269 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10160), .ZN(P1_U3318) );
  AND2_X1 U11270 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10160), .ZN(P1_U3319) );
  AND2_X1 U11271 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10160), .ZN(P1_U3320) );
  AND2_X1 U11272 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10160), .ZN(P1_U3321) );
  NOR2_X1 U11273 ( .A1(n10163), .A2(n10161), .ZN(P1_U3322) );
  NOR2_X1 U11274 ( .A1(n10163), .A2(n10162), .ZN(P1_U3323) );
  INV_X1 U11275 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10164) );
  AOI22_X1 U11276 ( .A1(n10232), .A2(n10165), .B1(n10164), .B2(n10230), .ZN(
        P1_U3453) );
  INV_X1 U11277 ( .A(n10166), .ZN(n10171) );
  OAI21_X1 U11278 ( .B1(n10168), .B2(n10213), .A(n10167), .ZN(n10170) );
  AOI211_X1 U11279 ( .C1(n10219), .C2(n10171), .A(n10170), .B(n10169), .ZN(
        n10234) );
  AOI22_X1 U11280 ( .A1(n10232), .A2(n10234), .B1(n10172), .B2(n10230), .ZN(
        P1_U3456) );
  OAI21_X1 U11281 ( .B1(n5614), .B2(n10213), .A(n10173), .ZN(n10176) );
  INV_X1 U11282 ( .A(n10174), .ZN(n10175) );
  AOI211_X1 U11283 ( .C1(n10177), .C2(n10221), .A(n10176), .B(n10175), .ZN(
        n10236) );
  INV_X1 U11284 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10178) );
  AOI22_X1 U11285 ( .A1(n10232), .A2(n10236), .B1(n10178), .B2(n10230), .ZN(
        P1_U3459) );
  OAI21_X1 U11286 ( .B1(n10180), .B2(n10213), .A(n10179), .ZN(n10182) );
  AOI211_X1 U11287 ( .C1(n10221), .C2(n10183), .A(n10182), .B(n10181), .ZN(
        n10237) );
  AOI22_X1 U11288 ( .A1(n10232), .A2(n10237), .B1(n5022), .B2(n10230), .ZN(
        P1_U3462) );
  OAI21_X1 U11289 ( .B1(n10185), .B2(n10213), .A(n10184), .ZN(n10188) );
  INV_X1 U11290 ( .A(n10186), .ZN(n10187) );
  AOI211_X1 U11291 ( .C1(n10189), .C2(n10221), .A(n10188), .B(n10187), .ZN(
        n10238) );
  INV_X1 U11292 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10190) );
  AOI22_X1 U11293 ( .A1(n10232), .A2(n10238), .B1(n10190), .B2(n10230), .ZN(
        P1_U3465) );
  AOI21_X1 U11294 ( .B1(n10223), .B2(n10192), .A(n10191), .ZN(n10193) );
  OAI211_X1 U11295 ( .C1(n10196), .C2(n10195), .A(n10194), .B(n10193), .ZN(
        n10197) );
  INV_X1 U11296 ( .A(n10197), .ZN(n10239) );
  INV_X1 U11297 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10198) );
  AOI22_X1 U11298 ( .A1(n10232), .A2(n10239), .B1(n10198), .B2(n10230), .ZN(
        P1_U3468) );
  OAI211_X1 U11299 ( .C1(n10201), .C2(n10213), .A(n10200), .B(n10199), .ZN(
        n10202) );
  AOI21_X1 U11300 ( .B1(n10221), .B2(n10203), .A(n10202), .ZN(n10241) );
  AOI22_X1 U11301 ( .A1(n10232), .A2(n10241), .B1(n10204), .B2(n10230), .ZN(
        P1_U3471) );
  AND2_X1 U11302 ( .A1(n10205), .A2(n10219), .ZN(n10209) );
  OAI21_X1 U11303 ( .B1(n10207), .B2(n10213), .A(n10206), .ZN(n10208) );
  NOR3_X1 U11304 ( .A1(n10210), .A2(n10209), .A3(n10208), .ZN(n10242) );
  INV_X1 U11305 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10211) );
  AOI22_X1 U11306 ( .A1(n10232), .A2(n10242), .B1(n10211), .B2(n10230), .ZN(
        P1_U3474) );
  OAI21_X1 U11307 ( .B1(n10214), .B2(n10213), .A(n10212), .ZN(n10217) );
  INV_X1 U11308 ( .A(n10215), .ZN(n10216) );
  AOI211_X1 U11309 ( .C1(n10219), .C2(n10218), .A(n10217), .B(n10216), .ZN(
        n10244) );
  INV_X1 U11310 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10220) );
  AOI22_X1 U11311 ( .A1(n10232), .A2(n10244), .B1(n10220), .B2(n10230), .ZN(
        P1_U3477) );
  AND2_X1 U11312 ( .A1(n10222), .A2(n10221), .ZN(n10229) );
  NAND2_X1 U11313 ( .A1(n10224), .A2(n10223), .ZN(n10225) );
  NAND2_X1 U11314 ( .A1(n10226), .A2(n10225), .ZN(n10227) );
  NOR3_X1 U11315 ( .A1(n10229), .A2(n10228), .A3(n10227), .ZN(n10247) );
  INV_X1 U11316 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10231) );
  AOI22_X1 U11317 ( .A1(n10232), .A2(n10247), .B1(n10231), .B2(n10230), .ZN(
        P1_U3480) );
  AOI22_X1 U11318 ( .A1(n10248), .A2(n10234), .B1(n10233), .B2(n10245), .ZN(
        P1_U3523) );
  AOI22_X1 U11319 ( .A1(n10248), .A2(n10236), .B1(n10235), .B2(n10245), .ZN(
        P1_U3524) );
  AOI22_X1 U11320 ( .A1(n10248), .A2(n10237), .B1(n6318), .B2(n10245), .ZN(
        P1_U3525) );
  AOI22_X1 U11321 ( .A1(n10248), .A2(n10238), .B1(n6320), .B2(n10245), .ZN(
        P1_U3526) );
  AOI22_X1 U11322 ( .A1(n10248), .A2(n10239), .B1(n6321), .B2(n10245), .ZN(
        P1_U3527) );
  INV_X1 U11323 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10240) );
  AOI22_X1 U11324 ( .A1(n10248), .A2(n10241), .B1(n10240), .B2(n10245), .ZN(
        P1_U3528) );
  AOI22_X1 U11325 ( .A1(n10248), .A2(n10242), .B1(n6322), .B2(n10245), .ZN(
        P1_U3529) );
  INV_X1 U11326 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10243) );
  AOI22_X1 U11327 ( .A1(n10248), .A2(n10244), .B1(n10243), .B2(n10245), .ZN(
        P1_U3530) );
  INV_X1 U11328 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10246) );
  AOI22_X1 U11329 ( .A1(n10248), .A2(n10247), .B1(n10246), .B2(n10245), .ZN(
        P1_U3531) );
  OAI21_X1 U11330 ( .B1(n10250), .B2(n8385), .A(n10249), .ZN(n10281) );
  INV_X1 U11331 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10252) );
  OAI22_X1 U11332 ( .A1(n10253), .A2(n10252), .B1(n10278), .B2(n10251), .ZN(
        n10267) );
  INV_X1 U11333 ( .A(n10281), .ZN(n10266) );
  AOI211_X1 U11334 ( .C1(n6522), .C2(n10256), .A(n10255), .B(n10254), .ZN(
        n10259) );
  INV_X1 U11335 ( .A(n6983), .ZN(n10258) );
  OAI21_X1 U11336 ( .B1(n10259), .B2(n10258), .A(n10257), .ZN(n10264) );
  AOI22_X1 U11337 ( .A1(n6168), .A2(n10262), .B1(n10261), .B2(n10260), .ZN(
        n10263) );
  OAI211_X1 U11338 ( .C1(n10266), .C2(n10265), .A(n10264), .B(n10263), .ZN(
        n10279) );
  AOI211_X1 U11339 ( .C1(n10268), .C2(n10281), .A(n10267), .B(n10279), .ZN(
        n10270) );
  AOI22_X1 U11340 ( .A1(n10272), .A2(n10271), .B1(n10270), .B2(n10269), .ZN(
        P2_U3231) );
  INV_X1 U11341 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10274) );
  AOI22_X1 U11342 ( .A1(n10310), .A2(n10274), .B1(n10273), .B2(n10308), .ZN(
        P2_U3390) );
  NOR2_X1 U11343 ( .A1(n6522), .A2(n10302), .ZN(n10276) );
  AOI211_X1 U11344 ( .C1(n10282), .C2(n10277), .A(n10276), .B(n10275), .ZN(
        n10312) );
  AOI22_X1 U11345 ( .A1(n10310), .A2(n5730), .B1(n10312), .B2(n10308), .ZN(
        P2_U3393) );
  INV_X1 U11346 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10283) );
  NOR2_X1 U11347 ( .A1(n10278), .A2(n10302), .ZN(n10280) );
  AOI211_X1 U11348 ( .C1(n10282), .C2(n10281), .A(n10280), .B(n10279), .ZN(
        n10314) );
  AOI22_X1 U11349 ( .A1(n10310), .A2(n10283), .B1(n10314), .B2(n10308), .ZN(
        P2_U3396) );
  INV_X1 U11350 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10288) );
  OAI21_X1 U11351 ( .B1(n10285), .B2(n10302), .A(n10284), .ZN(n10286) );
  AOI21_X1 U11352 ( .B1(n10293), .B2(n10287), .A(n10286), .ZN(n10315) );
  AOI22_X1 U11353 ( .A1(n10310), .A2(n10288), .B1(n10315), .B2(n10308), .ZN(
        P2_U3399) );
  INV_X1 U11354 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10294) );
  OAI21_X1 U11355 ( .B1(n10290), .B2(n10302), .A(n10289), .ZN(n10291) );
  AOI21_X1 U11356 ( .B1(n10293), .B2(n10292), .A(n10291), .ZN(n10317) );
  AOI22_X1 U11357 ( .A1(n10310), .A2(n10294), .B1(n10317), .B2(n10308), .ZN(
        P2_U3402) );
  INV_X1 U11358 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10301) );
  NOR2_X1 U11359 ( .A1(n10296), .A2(n10295), .ZN(n10297) );
  AOI211_X1 U11360 ( .C1(n10300), .C2(n10299), .A(n10298), .B(n10297), .ZN(
        n10319) );
  AOI22_X1 U11361 ( .A1(n10310), .A2(n10301), .B1(n10319), .B2(n10308), .ZN(
        P2_U3405) );
  INV_X1 U11362 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10309) );
  OAI22_X1 U11363 ( .A1(n10305), .A2(n10304), .B1(n10303), .B2(n10302), .ZN(
        n10306) );
  NOR2_X1 U11364 ( .A1(n10307), .A2(n10306), .ZN(n10322) );
  AOI22_X1 U11365 ( .A1(n10310), .A2(n10309), .B1(n10322), .B2(n10308), .ZN(
        P2_U3411) );
  AOI22_X1 U11366 ( .A1(n10323), .A2(n10312), .B1(n10311), .B2(n10320), .ZN(
        P2_U3460) );
  AOI22_X1 U11367 ( .A1(n10323), .A2(n10314), .B1(n10313), .B2(n10320), .ZN(
        P2_U3461) );
  AOI22_X1 U11368 ( .A1(n10323), .A2(n10315), .B1(n4761), .B2(n10320), .ZN(
        P2_U3462) );
  AOI22_X1 U11369 ( .A1(n10323), .A2(n10317), .B1(n10316), .B2(n10320), .ZN(
        P2_U3463) );
  INV_X1 U11370 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10318) );
  AOI22_X1 U11371 ( .A1(n10323), .A2(n10319), .B1(n10318), .B2(n10320), .ZN(
        P2_U3464) );
  AOI22_X1 U11372 ( .A1(n10323), .A2(n10322), .B1(n10321), .B2(n10320), .ZN(
        P2_U3466) );
  OAI222_X1 U11373 ( .A1(n10328), .A2(n10327), .B1(n10328), .B2(n10326), .C1(
        n10325), .C2(n10324), .ZN(ADD_1068_U5) );
  XOR2_X1 U11374 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI21_X1 U11375 ( .B1(n10331), .B2(n10330), .A(n10329), .ZN(n10332) );
  XNOR2_X1 U11376 ( .A(n10332), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1068_U55)
         );
  OAI21_X1 U11377 ( .B1(n10335), .B2(n10334), .A(n10333), .ZN(ADD_1068_U56) );
  OAI21_X1 U11378 ( .B1(n10338), .B2(n10337), .A(n10336), .ZN(ADD_1068_U57) );
  OAI21_X1 U11379 ( .B1(n10341), .B2(n10340), .A(n10339), .ZN(ADD_1068_U58) );
  OAI21_X1 U11380 ( .B1(n10344), .B2(n10343), .A(n10342), .ZN(ADD_1068_U59) );
  OAI21_X1 U11381 ( .B1(n10347), .B2(n10346), .A(n10345), .ZN(ADD_1068_U60) );
  OAI21_X1 U11382 ( .B1(n10350), .B2(n10349), .A(n10348), .ZN(ADD_1068_U61) );
  OAI21_X1 U11383 ( .B1(n10353), .B2(n10352), .A(n10351), .ZN(ADD_1068_U62) );
  OAI21_X1 U11384 ( .B1(n10356), .B2(n10355), .A(n10354), .ZN(ADD_1068_U63) );
  OAI21_X1 U11385 ( .B1(n10359), .B2(n10358), .A(n10357), .ZN(ADD_1068_U50) );
  OAI21_X1 U11386 ( .B1(n10362), .B2(n10361), .A(n10360), .ZN(ADD_1068_U51) );
  OAI21_X1 U11387 ( .B1(n10365), .B2(n10364), .A(n10363), .ZN(ADD_1068_U47) );
  OAI21_X1 U11388 ( .B1(n10368), .B2(n10367), .A(n10366), .ZN(ADD_1068_U49) );
  OAI21_X1 U11389 ( .B1(n10371), .B2(n10370), .A(n10369), .ZN(ADD_1068_U48) );
  AOI21_X1 U11390 ( .B1(n10374), .B2(n10373), .A(n10372), .ZN(ADD_1068_U54) );
  AOI21_X1 U11391 ( .B1(n10377), .B2(n10376), .A(n10375), .ZN(ADD_1068_U53) );
  OAI21_X1 U11392 ( .B1(n10380), .B2(n10379), .A(n10378), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4827 ( .A(n5914), .Z(n6103) );
endmodule

