

module b20_C_AntiSAT_k_128_5 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, 
        ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, 
        ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, 
        ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, 
        U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, 
        P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, 
        P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, 
        P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, 
        P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, 
        P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, 
        P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, 
        P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, 
        P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, 
        P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, 
        P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, 
        P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, 
        P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, 
        P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, 
        P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, 
        P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, 
        P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, 
        P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, 
        P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, 
        P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, 
        P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, 
        P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, 
        P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, 
        P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, 
        P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, 
        P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, 
        P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, 
        P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, 
        P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, 
        P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4329, n4330, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323;

  INV_X1 U4835 ( .A(n8293), .ZN(n6412) );
  CLKBUF_X2 U4836 ( .A(n6088), .Z(n4335) );
  NAND2_X1 U4837 ( .A1(n9087), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4478) );
  INV_X1 U4838 ( .A(n6305), .ZN(n6103) );
  AOI21_X1 U4840 ( .B1(n8851), .B2(n8516), .A(n5614), .ZN(n8832) );
  NAND2_X1 U4841 ( .A1(n5575), .A2(n5574), .ZN(n8892) );
  INV_X1 U4842 ( .A(n5358), .ZN(n5788) );
  NAND2_X2 U4843 ( .A1(n6046), .A2(n6653), .ZN(n6546) );
  INV_X1 U4844 ( .A(n6546), .ZN(n6587) );
  INV_X1 U4845 ( .A(n6570), .ZN(n6584) );
  NAND2_X1 U4846 ( .A1(n7553), .A2(n7703), .ZN(n7663) );
  NOR2_X1 U4847 ( .A1(n7485), .A2(n7145), .ZN(n7213) );
  AOI21_X1 U4848 ( .B1(n7767), .B2(n7768), .A(n7766), .ZN(n7808) );
  INV_X1 U4849 ( .A(n5787), .ZN(n5314) );
  INV_X1 U4850 ( .A(n8628), .ZN(n7595) );
  INV_X1 U4851 ( .A(n6062), .ZN(n6411) );
  AND3_X1 U4853 ( .A1(n6099), .A2(n6098), .A3(n6097), .ZN(n9864) );
  OAI21_X1 U4854 ( .B1(n6051), .B2(P1_IR_REG_27__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n4510) );
  AND4_X1 U4855 ( .A1(n4400), .A2(n5270), .A3(n5268), .A4(n5269), .ZN(n7074)
         );
  INV_X1 U4857 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6044) );
  NAND4_X2 U4858 ( .A1(n5634), .A2(n5633), .A3(n5632), .A4(n5631), .ZN(n8833)
         );
  OAI21_X2 U4860 ( .B1(n5082), .B2(n4334), .A(n8334), .ZN(n8288) );
  OAI211_X2 U4861 ( .C1(n5314), .C2(n6670), .A(n5277), .B(n5276), .ZN(n6988)
         );
  NOR2_X1 U4862 ( .A1(n7678), .A2(n7763), .ZN(n7679) );
  OR2_X2 U4863 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5225) );
  OAI21_X1 U4864 ( .B1(n6972), .B2(n6971), .A(n4526), .ZN(n4527) );
  NAND2_X2 U4865 ( .A1(n4361), .A2(n4808), .ZN(n7140) );
  OAI211_X2 U4866 ( .C1(n4780), .C2(n6206), .A(n4778), .B(n6226), .ZN(n9120)
         );
  AND2_X1 U4867 ( .A1(n5263), .A2(n6662), .ZN(n4330) );
  BUF_X2 U4868 ( .A(n5280), .Z(n5745) );
  AOI211_X1 U4871 ( .C1(n9709), .C2(n9398), .A(n9595), .B(n4357), .ZN(n9634)
         );
  NAND2_X1 U4872 ( .A1(n7763), .A2(n7672), .ZN(n8239) );
  NAND2_X1 U4873 ( .A1(n7211), .A2(n8390), .ZN(n8394) );
  AND2_X1 U4874 ( .A1(n7510), .A2(n9875), .ZN(n7530) );
  INV_X2 U4875 ( .A(n6305), .ZN(n6286) );
  INV_X1 U4876 ( .A(n8381), .ZN(n4334) );
  INV_X1 U4877 ( .A(n4527), .ZN(n8488) );
  INV_X2 U4878 ( .A(n8632), .ZN(n7359) );
  INV_X1 U4879 ( .A(n8631), .ZN(n5700) );
  INV_X1 U4880 ( .A(n8629), .ZN(n7475) );
  INV_X1 U4881 ( .A(n8634), .ZN(n10029) );
  INV_X4 U4882 ( .A(n6656), .ZN(n5986) );
  NAND2_X2 U4883 ( .A1(n6062), .A2(n6661), .ZN(n6271) );
  XNOR2_X1 U4884 ( .A(n6045), .B(n6044), .ZN(n6047) );
  NAND2_X1 U4885 ( .A1(n6026), .A2(n6021), .ZN(n8372) );
  AND3_X1 U4886 ( .A1(n6017), .A2(n6044), .A3(n4785), .ZN(n6004) );
  INV_X1 U4887 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4785) );
  NOR2_X1 U4888 ( .A1(n8441), .A2(n4736), .ZN(n8449) );
  OR2_X1 U4889 ( .A1(n9708), .A2(n4699), .ZN(n4825) );
  OAI21_X1 U4890 ( .B1(n8379), .B2(n4735), .A(n4733), .ZN(n4736) );
  AND2_X1 U4891 ( .A1(n9375), .A2(n4700), .ZN(n8189) );
  AOI21_X1 U4892 ( .B1(n4606), .B2(n4792), .A(n9377), .ZN(n9380) );
  OAI21_X1 U4893 ( .B1(n8156), .B2(n4930), .A(n4925), .ZN(n4494) );
  INV_X1 U4894 ( .A(n4818), .ZN(n6645) );
  NAND2_X1 U4895 ( .A1(n4817), .A2(n4816), .ZN(n4818) );
  OR2_X1 U4896 ( .A1(n4898), .A2(n4539), .ZN(n4537) );
  AND2_X1 U4897 ( .A1(n8486), .A2(n4899), .ZN(n4898) );
  NOR2_X1 U4898 ( .A1(n9484), .A2(n4506), .ZN(n8148) );
  NAND2_X1 U4899 ( .A1(n4507), .A2(n4416), .ZN(n9484) );
  AND2_X1 U4900 ( .A1(n4509), .A2(n4508), .ZN(n9504) );
  INV_X1 U4901 ( .A(n4623), .ZN(n4622) );
  OAI21_X1 U4902 ( .B1(n4343), .B2(n4358), .A(n6473), .ZN(n4623) );
  AND2_X1 U4903 ( .A1(n9024), .A2(n8482), .ZN(n5928) );
  AOI21_X1 U4904 ( .B1(n4564), .B2(n4565), .A(n4563), .ZN(n4562) );
  NAND2_X1 U4905 ( .A1(n5618), .A2(n5617), .ZN(n9030) );
  OAI21_X1 U4906 ( .B1(n4918), .B2(n4544), .A(n4542), .ZN(n4550) );
  OR2_X1 U4907 ( .A1(n8472), .A2(n8620), .ZN(n8473) );
  OR2_X1 U4908 ( .A1(n9739), .A2(n8165), .ZN(n8304) );
  OAI21_X1 U4909 ( .B1(n10076), .B2(n4401), .A(n4349), .ZN(n8037) );
  NAND2_X1 U4910 ( .A1(n7868), .A2(n7867), .ZN(n7911) );
  CLKBUF_X1 U4911 ( .A(n7857), .Z(n4598) );
  OAI21_X1 U4912 ( .B1(n4569), .B2(n8625), .A(n7876), .ZN(n4568) );
  NAND2_X1 U4913 ( .A1(n6437), .A2(n6436), .ZN(n9744) );
  NAND2_X1 U4914 ( .A1(n6397), .A2(n6396), .ZN(n9528) );
  OR2_X1 U4915 ( .A1(n7898), .A2(n7897), .ZN(n10076) );
  NAND2_X1 U4916 ( .A1(n4434), .A2(n4432), .ZN(n5579) );
  AOI21_X1 U4917 ( .B1(n8250), .B2(n4693), .A(n4386), .ZN(n4690) );
  AND2_X1 U4918 ( .A1(n7777), .A2(n8242), .ZN(n7778) );
  NAND2_X1 U4919 ( .A1(n6352), .A2(n6351), .ZN(n9761) );
  NAND2_X1 U4920 ( .A1(n7675), .A2(n7674), .ZN(n7783) );
  AND2_X1 U4921 ( .A1(n4777), .A2(n8401), .ZN(n7669) );
  AND2_X1 U4922 ( .A1(n7591), .A2(n8627), .ZN(n7766) );
  OR2_X1 U4923 ( .A1(n6155), .A2(n6154), .ZN(n5078) );
  NAND2_X1 U4924 ( .A1(n6337), .A2(n6336), .ZN(n9766) );
  NAND2_X1 U4925 ( .A1(n8137), .A2(n8138), .ZN(n9604) );
  AND4_X1 U4926 ( .A1(n5623), .A2(n5622), .A3(n5621), .A4(n5620), .ZN(n8823)
         );
  AND2_X1 U4927 ( .A1(n4431), .A2(n5009), .ZN(n5490) );
  OR2_X1 U4928 ( .A1(n8203), .A2(n8381), .ZN(n4760) );
  NAND2_X1 U4929 ( .A1(n8394), .A2(n8207), .ZN(n8203) );
  NAND2_X1 U4930 ( .A1(n5384), .A2(n5383), .ZN(n10062) );
  NAND2_X1 U4931 ( .A1(n6192), .A2(n6191), .ZN(n7697) );
  NAND2_X1 U4932 ( .A1(n6212), .A2(n6211), .ZN(n7763) );
  NAND2_X1 U4933 ( .A1(n5369), .A2(n5368), .ZN(n7560) );
  OR2_X1 U4934 ( .A1(n9990), .A2(n9989), .ZN(n4459) );
  NAND2_X1 U4935 ( .A1(n5325), .A2(n5128), .ZN(n5338) );
  NAND2_X1 U4936 ( .A1(n5323), .A2(n5083), .ZN(n5325) );
  NAND2_X4 U4937 ( .A1(n6546), .A2(n6570), .ZN(n6131) );
  NOR2_X1 U4938 ( .A1(n7318), .A2(n4453), .ZN(n9947) );
  NAND4_X1 U4939 ( .A1(n6078), .A2(n6077), .A3(n6076), .A4(n6075), .ZN(n9293)
         );
  CLKBUF_X3 U4940 ( .A(n8488), .Z(n8491) );
  AND2_X1 U4941 ( .A1(n4456), .A2(n4455), .ZN(n7318) );
  NAND2_X1 U4942 ( .A1(n6395), .A2(n8372), .ZN(n7162) );
  OAI211_X2 U4943 ( .C1(n6659), .C2(n8293), .A(n4512), .B(n6065), .ZN(n4511)
         );
  CLKBUF_X1 U4944 ( .A(n6395), .Z(n8383) );
  AND2_X1 U4945 ( .A1(n6047), .A2(n8372), .ZN(n8437) );
  OR2_X1 U4946 ( .A1(n8338), .A2(n6899), .ZN(n4636) );
  OR2_X1 U4947 ( .A1(n6271), .A2(n6663), .ZN(n4512) );
  NOR2_X2 U4948 ( .A1(n5953), .A2(n5986), .ZN(n5656) );
  NAND2_X1 U4949 ( .A1(n4637), .A2(n6610), .ZN(n8193) );
  NAND4_X1 U4950 ( .A1(n5287), .A2(n5286), .A3(n5285), .A4(n5284), .ZN(n8634)
         );
  NOR2_X1 U4951 ( .A1(n4781), .A2(n9777), .ZN(n6011) );
  NAND2_X2 U4952 ( .A1(n6062), .A2(n6662), .ZN(n8293) );
  NAND2_X1 U4953 ( .A1(n4937), .A2(n4784), .ZN(n8500) );
  NAND2_X1 U4954 ( .A1(n6410), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6045) );
  XNOR2_X1 U4955 ( .A(n6022), .B(n4785), .ZN(n8338) );
  OAI21_X1 U4956 ( .B1(n4351), .B2(n4975), .A(n5084), .ZN(n4974) );
  NAND2_X1 U4957 ( .A1(n6021), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6022) );
  OAI21_X1 U4958 ( .B1(n6038), .B2(n6029), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6030) );
  CLKBUF_X1 U4959 ( .A(n5256), .Z(n5607) );
  INV_X2 U4960 ( .A(n5263), .ZN(n5551) );
  NOR2_X1 U4961 ( .A1(n5364), .A2(n4688), .ZN(n4687) );
  NAND2_X2 U4962 ( .A1(n5655), .A2(n6702), .ZN(n5263) );
  NAND2_X1 U4963 ( .A1(n5670), .A2(n5669), .ZN(n5689) );
  NAND2_X1 U4964 ( .A1(n9087), .A2(n4826), .ZN(n5239) );
  NOR2_X1 U4965 ( .A1(n6041), .A2(n6019), .ZN(n6023) );
  NAND2_X1 U4966 ( .A1(n6041), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6377) );
  AND2_X1 U4967 ( .A1(n5672), .A2(n5664), .ZN(n8029) );
  MUX2_X1 U4968 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5668), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n5670) );
  INV_X2 U4969 ( .A(n7905), .ZN(n4336) );
  NAND2_X1 U4970 ( .A1(n4595), .A2(n10124), .ZN(n9087) );
  INV_X1 U4971 ( .A(n5237), .ZN(n4595) );
  AND2_X1 U4972 ( .A1(n5366), .A2(n5095), .ZN(n5667) );
  INV_X1 U4973 ( .A(n5111), .ZN(n6662) );
  XNOR2_X1 U4974 ( .A(n4448), .B(P2_IR_REG_2__SCAN_IN), .ZN(n4602) );
  NOR2_X1 U4975 ( .A1(n4499), .A2(n4501), .ZN(n4496) );
  NAND2_X1 U4976 ( .A1(n5254), .A2(n5253), .ZN(n6807) );
  NAND2_X2 U4977 ( .A1(n5006), .A2(n5005), .ZN(n5111) );
  NAND3_X1 U4978 ( .A1(n4436), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5005) );
  AND4_X1 U4979 ( .A1(n5094), .A2(n5093), .A3(n5092), .A4(n5091), .ZN(n5095)
         );
  NAND3_X1 U4980 ( .A1(n8770), .A2(n5008), .A3(n5007), .ZN(n5006) );
  NOR2_X2 U4981 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5252) );
  INV_X2 U4982 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X1 U4983 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n6018) );
  INV_X1 U4984 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5995) );
  NOR2_X1 U4985 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n4877) );
  INV_X1 U4986 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4436) );
  INV_X1 U4987 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4477) );
  INV_X1 U4988 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5534) );
  NOR2_X1 U4989 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5223) );
  INV_X4 U4990 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X2 U4991 ( .A1(n5443), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5462) );
  XNOR2_X1 U4992 ( .A(n4510), .B(n6050), .ZN(n6617) );
  INV_X1 U4993 ( .A(n5256), .ZN(n4338) );
  NOR2_X2 U4994 ( .A1(n4352), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5509) );
  OR2_X2 U4995 ( .A1(n5481), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n4352) );
  INV_X2 U4996 ( .A(n4511), .ZN(n7636) );
  XNOR2_X1 U4997 ( .A(n7140), .B(n4511), .ZN(n7122) );
  OR2_X2 U4998 ( .A1(n5298), .A2(n8826), .ZN(n5634) );
  OR2_X1 U4999 ( .A1(n9709), .A2(n9397), .ZN(n8358) );
  AND2_X1 U5000 ( .A1(n4879), .A2(n4878), .ZN(n4706) );
  NOR2_X1 U5001 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n4879) );
  NOR2_X1 U5002 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4878) );
  OAI21_X1 U5003 ( .B1(n5024), .B2(n5022), .A(n5961), .ZN(n5021) );
  INV_X1 U5004 ( .A(n5960), .ZN(n5022) );
  OR2_X1 U5005 ( .A1(n9047), .A2(n8877), .ZN(n5894) );
  OAI21_X1 U5006 ( .B1(n5500), .B2(n4415), .A(n5163), .ZN(n5518) );
  INV_X1 U5007 ( .A(n5501), .ZN(n5162) );
  INV_X1 U5008 ( .A(n5151), .ZN(n4979) );
  BUF_X1 U5009 ( .A(n5301), .Z(n5763) );
  BUF_X1 U5010 ( .A(n5282), .Z(n5760) );
  INV_X1 U5011 ( .A(n5256), .ZN(n5298) );
  NAND2_X1 U5012 ( .A1(n5238), .A2(n5239), .ZN(n5282) );
  NAND2_X1 U5013 ( .A1(n9090), .A2(n5239), .ZN(n5301) );
  AND2_X1 U5014 ( .A1(n9094), .A2(n5238), .ZN(n5280) );
  NOR2_X1 U5015 ( .A1(n5238), .A2(n5239), .ZN(n5256) );
  XNOR2_X1 U5016 ( .A(n7313), .B(n9983), .ZN(n9977) );
  AND2_X1 U5017 ( .A1(n6583), .A2(n6582), .ZN(n9397) );
  OAI21_X1 U5018 ( .B1(n8148), .B2(n4942), .A(n4940), .ZN(n4605) );
  AOI21_X1 U5019 ( .B1(n4941), .B2(n8151), .A(n4950), .ZN(n4940) );
  NAND2_X1 U5020 ( .A1(n4943), .A2(n8151), .ZN(n4942) );
  NAND2_X1 U5021 ( .A1(n6900), .A2(n8382), .ZN(n9608) );
  NAND2_X1 U5022 ( .A1(n5874), .A2(n5986), .ZN(n4732) );
  NAND2_X1 U5023 ( .A1(n4442), .A2(n8274), .ZN(n4441) );
  NAND2_X1 U5024 ( .A1(n4443), .A2(n8331), .ZN(n4442) );
  AND2_X1 U5025 ( .A1(n4741), .A2(n4334), .ZN(n4738) );
  AND2_X1 U5026 ( .A1(n8356), .A2(n8351), .ZN(n4741) );
  NOR2_X1 U5027 ( .A1(n4405), .A2(n4907), .ZN(n4906) );
  INV_X1 U5028 ( .A(n8471), .ZN(n4907) );
  NAND2_X1 U5029 ( .A1(n4392), .A2(n4471), .ZN(n4844) );
  NAND2_X1 U5030 ( .A1(n5965), .A2(n5933), .ZN(n4471) );
  NAND2_X1 U5031 ( .A1(n8961), .A2(n8784), .ZN(n4845) );
  OR2_X1 U5032 ( .A1(n7337), .A2(n9939), .ZN(n4892) );
  NAND2_X1 U5033 ( .A1(n7337), .A2(n4893), .ZN(n4891) );
  NOR2_X1 U5034 ( .A1(n4895), .A2(n7338), .ZN(n4893) );
  NAND2_X1 U5035 ( .A1(n4685), .A2(n4684), .ZN(n7337) );
  INV_X1 U5036 ( .A(n6747), .ZN(n4684) );
  AND2_X1 U5037 ( .A1(n9967), .A2(n7312), .ZN(n7313) );
  NAND2_X1 U5038 ( .A1(n4873), .A2(n4872), .ZN(n9997) );
  INV_X1 U5039 ( .A(n9999), .ZN(n4872) );
  XNOR2_X1 U5040 ( .A(n4463), .B(P2_IR_REG_27__SCAN_IN), .ZN(n5655) );
  AOI21_X1 U5041 ( .B1(n4836), .B2(n4372), .A(n9086), .ZN(n4463) );
  INV_X1 U5042 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4834) );
  NAND2_X1 U5043 ( .A1(n5004), .A2(n5002), .ZN(n5933) );
  NOR2_X1 U5044 ( .A1(n8619), .A2(n5003), .ZN(n5002) );
  INV_X1 U5045 ( .A(n5759), .ZN(n5003) );
  NAND2_X1 U5046 ( .A1(n5028), .A2(n5030), .ZN(n5024) );
  NAND2_X1 U5047 ( .A1(n5956), .A2(n5029), .ZN(n5028) );
  OR2_X1 U5048 ( .A1(n8816), .A2(n8824), .ZN(n5935) );
  NAND2_X1 U5049 ( .A1(n7101), .A2(n10027), .ZN(n5806) );
  NOR2_X1 U5050 ( .A1(n5239), .A2(n6817), .ZN(n5015) );
  NAND2_X1 U5051 ( .A1(n4607), .A2(n4345), .ZN(n5018) );
  NOR2_X1 U5052 ( .A1(n5928), .A2(n5925), .ZN(n4861) );
  INV_X1 U5053 ( .A(n9042), .ZN(n8477) );
  NAND2_X1 U5054 ( .A1(n4389), .A2(n5075), .ZN(n5067) );
  NAND2_X1 U5055 ( .A1(n8477), .A2(n8848), .ZN(n5916) );
  OR2_X1 U5056 ( .A1(n8534), .A2(n8893), .ZN(n5893) );
  NAND2_X1 U5057 ( .A1(n5036), .A2(n8903), .ZN(n5035) );
  AND2_X1 U5058 ( .A1(n5044), .A2(n5043), .ZN(n5042) );
  NAND2_X1 U5059 ( .A1(n4342), .A2(n4840), .ZN(n4837) );
  INV_X1 U5060 ( .A(n7695), .ZN(n5980) );
  OR2_X1 U5061 ( .A1(n5326), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5340) );
  AND2_X1 U5062 ( .A1(n4636), .A2(n6896), .ZN(n6046) );
  NAND2_X1 U5063 ( .A1(n7292), .A2(n6140), .ZN(n6155) );
  OR2_X1 U5064 ( .A1(n9352), .A2(n9355), .ZN(n8434) );
  OR2_X1 U5065 ( .A1(n9734), .A2(n9491), .ZN(n9454) );
  NAND2_X1 U5066 ( .A1(n9560), .A2(n9548), .ZN(n9547) );
  NAND2_X1 U5067 ( .A1(n4587), .A2(n4966), .ZN(n7537) );
  AOI21_X1 U5068 ( .B1(n7541), .B2(n4967), .A(n4382), .ZN(n4966) );
  NAND2_X1 U5069 ( .A1(n7220), .A2(n4367), .ZN(n4587) );
  INV_X1 U5070 ( .A(n7507), .ZN(n4967) );
  INV_X1 U5071 ( .A(n6886), .ZN(n6890) );
  OAI21_X1 U5072 ( .B1(n5758), .B2(SI_29_), .A(n5731), .ZN(n5750) );
  INV_X1 U5073 ( .A(n6005), .ZN(n4498) );
  NOR2_X1 U5074 ( .A1(n4500), .A2(n6157), .ZN(n4497) );
  NAND2_X1 U5075 ( .A1(n6000), .A2(n6033), .ZN(n4500) );
  INV_X1 U5076 ( .A(n5012), .ZN(n5009) );
  AOI21_X1 U5077 ( .B1(n7971), .B2(n7970), .A(n4412), .ZN(n7974) );
  INV_X1 U5078 ( .A(n8476), .ZN(n4558) );
  INV_X1 U5079 ( .A(n5760), .ZN(n5753) );
  INV_X1 U5080 ( .A(n5745), .ZN(n5761) );
  OR2_X1 U5081 ( .A1(n5282), .A2(n5257), .ZN(n5259) );
  OAI21_X1 U5082 ( .B1(n9911), .B2(n9912), .A(n4457), .ZN(n9930) );
  OR2_X1 U5083 ( .A1(n6720), .A2(n4602), .ZN(n4457) );
  OR2_X1 U5084 ( .A1(n9930), .A2(n9931), .ZN(n4456) );
  NOR2_X1 U5085 ( .A1(n9937), .A2(n10087), .ZN(n9936) );
  NAND2_X1 U5086 ( .A1(n4488), .A2(n4601), .ZN(n9967) );
  INV_X1 U5087 ( .A(n9969), .ZN(n4601) );
  OR2_X1 U5088 ( .A1(n9977), .A2(n7317), .ZN(n4599) );
  OR2_X1 U5089 ( .A1(n7316), .A2(n10121), .ZN(n4597) );
  NAND2_X1 U5090 ( .A1(n4888), .A2(n4887), .ZN(n7747) );
  OR2_X1 U5091 ( .A1(n7830), .A2(n7829), .ZN(n4658) );
  OR2_X1 U5092 ( .A1(n5457), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5458) );
  NOR2_X1 U5093 ( .A1(n7951), .A2(n5465), .ZN(n8656) );
  AND4_X1 U5094 ( .A1(n5654), .A2(n5653), .A3(n5652), .A4(n5651), .ZN(n8505)
         );
  OR2_X1 U5095 ( .A1(n9058), .A2(n8904), .ZN(n5890) );
  AND2_X1 U5096 ( .A1(n5598), .A2(n5597), .ZN(n8877) );
  NAND2_X1 U5097 ( .A1(n4468), .A2(n5885), .ZN(n5709) );
  INV_X1 U5098 ( .A(n8935), .ZN(n4468) );
  NAND2_X1 U5099 ( .A1(n7817), .A2(n7816), .ZN(n5434) );
  NAND2_X1 U5100 ( .A1(n5263), .A2(n6661), .ZN(n5358) );
  NAND2_X1 U5101 ( .A1(n8842), .A2(n5913), .ZN(n5712) );
  INV_X1 U5102 ( .A(n5358), .ZN(n5601) );
  INV_X1 U5103 ( .A(n5656), .ZN(n10028) );
  AND2_X1 U5104 ( .A1(n5953), .A2(n6656), .ZN(n8949) );
  NAND2_X1 U5105 ( .A1(n5667), .A2(n4381), .ZN(n5645) );
  XNOR2_X1 U5106 ( .A(n5550), .B(n5549), .ZN(n8763) );
  XNOR2_X1 U5107 ( .A(n5360), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9983) );
  INV_X1 U5108 ( .A(n5252), .ZN(n5253) );
  NAND2_X1 U5109 ( .A1(n6522), .A2(n8451), .ZN(n4633) );
  NAND2_X1 U5110 ( .A1(n6491), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6506) );
  INV_X1 U5111 ( .A(n9734), .ZN(n9479) );
  AND2_X1 U5112 ( .A1(n6566), .A2(n6565), .ZN(n9251) );
  AND4_X1 U5113 ( .A1(n6360), .A2(n6359), .A3(n6358), .A4(n6357), .ZN(n9261)
         );
  AND2_X1 U5114 ( .A1(n6011), .A2(n8500), .ZN(n6088) );
  AND2_X1 U5115 ( .A1(n8500), .A2(n9785), .ZN(n6089) );
  AND2_X1 U5116 ( .A1(n9785), .A2(n6012), .ZN(n6074) );
  NOR2_X1 U5117 ( .A1(n9785), .A2(n8500), .ZN(n6114) );
  INV_X1 U5118 ( .A(n8500), .ZN(n6012) );
  AND2_X1 U5119 ( .A1(n6011), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n4748) );
  OR2_X1 U5120 ( .A1(n8105), .A2(n8106), .ZN(n4524) );
  NAND2_X1 U5121 ( .A1(n4524), .A2(n4523), .ZN(n9325) );
  INV_X1 U5122 ( .A(n9327), .ZN(n4523) );
  INV_X1 U5123 ( .A(n9541), .ZN(n4815) );
  NAND2_X1 U5124 ( .A1(n4954), .A2(n4957), .ZN(n9584) );
  AND2_X1 U5125 ( .A1(n8142), .A2(n4958), .ZN(n4957) );
  NAND2_X1 U5126 ( .A1(n4394), .A2(n4951), .ZN(n4944) );
  AND2_X1 U5127 ( .A1(n9739), .A2(n9277), .ZN(n4506) );
  INV_X2 U5128 ( .A(n6271), .ZN(n8291) );
  INV_X1 U5129 ( .A(n6051), .ZN(n4764) );
  NAND2_X1 U5130 ( .A1(n4433), .A2(n5180), .ZN(n4432) );
  NAND2_X1 U5131 ( .A1(n5565), .A2(n5562), .ZN(n4434) );
  OAI21_X1 U5132 ( .B1(n5579), .B2(n4997), .A(n4995), .ZN(n5600) );
  INV_X1 U5133 ( .A(n4998), .ZN(n4997) );
  AOI21_X1 U5134 ( .B1(n4998), .B2(n4996), .A(n5599), .ZN(n4995) );
  INV_X1 U5135 ( .A(n5000), .ZN(n4996) );
  NAND2_X1 U5136 ( .A1(n4976), .A2(n4369), .ZN(n5438) );
  INV_X1 U5137 ( .A(n5435), .ZN(n4983) );
  NAND2_X1 U5138 ( .A1(n5338), .A2(n4351), .ZN(n5339) );
  AND2_X1 U5139 ( .A1(n7027), .A2(n7025), .ZN(n4901) );
  INV_X1 U5140 ( .A(n8848), .ZN(n8868) );
  INV_X1 U5141 ( .A(n5958), .ZN(n8965) );
  AOI21_X1 U5142 ( .B1(n8185), .B2(n9608), .A(n8184), .ZN(n9375) );
  AOI21_X1 U5143 ( .B1(n5812), .B2(n5813), .A(n4722), .ZN(n4721) );
  NAND2_X1 U5144 ( .A1(n4724), .A2(n4723), .ZN(n4722) );
  NAND2_X1 U5145 ( .A1(n4718), .A2(n7185), .ZN(n5828) );
  NAND2_X1 U5146 ( .A1(n4720), .A2(n4719), .ZN(n4718) );
  INV_X1 U5147 ( .A(n5818), .ZN(n4719) );
  NAND2_X1 U5148 ( .A1(n4725), .A2(n4721), .ZN(n4720) );
  MUX2_X1 U5149 ( .A(n5839), .B(n5843), .S(n5986), .Z(n5840) );
  NAND2_X1 U5150 ( .A1(n4730), .A2(n4727), .ZN(n4726) );
  NOR2_X1 U5151 ( .A1(n5883), .A2(n5986), .ZN(n4727) );
  NAND2_X1 U5152 ( .A1(n4440), .A2(n4370), .ZN(n8282) );
  INV_X1 U5153 ( .A(n4740), .ZN(n4739) );
  NOR2_X1 U5154 ( .A1(n5956), .A2(n5791), .ZN(n4590) );
  OR2_X1 U5155 ( .A1(n6742), .A2(n6741), .ZN(n4883) );
  NAND2_X1 U5156 ( .A1(n6742), .A2(n6741), .ZN(n4880) );
  NAND2_X1 U5157 ( .A1(n8816), .A2(n8798), .ZN(n5030) );
  INV_X1 U5158 ( .A(n6293), .ZN(n4797) );
  INV_X1 U5159 ( .A(n8220), .ZN(n4694) );
  NOR2_X1 U5160 ( .A1(n5546), .A2(n4646), .ZN(n4645) );
  INV_X1 U5161 ( .A(n5172), .ZN(n4646) );
  NAND2_X1 U5162 ( .A1(n6001), .A2(n4635), .ZN(n6041) );
  AND2_X1 U5163 ( .A1(n6000), .A2(n6017), .ZN(n4635) );
  NAND2_X1 U5164 ( .A1(n5166), .A2(n5165), .ZN(n5169) );
  NOR2_X1 U5165 ( .A1(n5012), .A2(n5011), .ZN(n5010) );
  NOR2_X1 U5166 ( .A1(n5471), .A2(SI_14_), .ZN(n5012) );
  NAND2_X1 U5167 ( .A1(n5456), .A2(n5013), .ZN(n4431) );
  AND2_X1 U5168 ( .A1(n5159), .A2(n5014), .ZN(n5013) );
  NAND2_X1 U5169 ( .A1(n5471), .A2(SI_14_), .ZN(n5014) );
  INV_X1 U5170 ( .A(n4545), .ZN(n4544) );
  AND2_X1 U5171 ( .A1(n4919), .A2(n4549), .ZN(n4548) );
  INV_X1 U5172 ( .A(n8544), .ZN(n4549) );
  OR2_X1 U5173 ( .A1(n6807), .A2(n6737), .ZN(n4661) );
  NAND2_X1 U5174 ( .A1(n5252), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6738) );
  NAND2_X1 U5175 ( .A1(n4883), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4881) );
  NAND2_X1 U5176 ( .A1(n4868), .A2(n9902), .ZN(n4869) );
  AND2_X1 U5177 ( .A1(n9924), .A2(n6728), .ZN(n4868) );
  NAND2_X1 U5178 ( .A1(n4881), .A2(n4880), .ZN(n4685) );
  AND2_X1 U5179 ( .A1(n4894), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4890) );
  INV_X1 U5180 ( .A(n9956), .ZN(n4671) );
  AND2_X1 U5181 ( .A1(n4452), .A2(n4451), .ZN(n8687) );
  NAND2_X1 U5182 ( .A1(n8681), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4451) );
  AND3_X1 U5183 ( .A1(n4678), .A2(n4677), .A3(n4428), .ZN(n8743) );
  NAND2_X1 U5184 ( .A1(n8965), .A2(n5959), .ZN(n5960) );
  NAND2_X1 U5185 ( .A1(n9024), .A2(n8833), .ZN(n5031) );
  INV_X1 U5186 ( .A(n5837), .ZN(n4848) );
  INV_X1 U5187 ( .A(n5058), .ZN(n5054) );
  OAI21_X1 U5188 ( .B1(n5090), .B2(n5060), .A(n8633), .ZN(n5059) );
  INV_X1 U5189 ( .A(n5090), .ZN(n5053) );
  NAND2_X1 U5190 ( .A1(n7110), .A2(n5297), .ZN(n5058) );
  NAND2_X1 U5191 ( .A1(n7074), .A2(n6988), .ZN(n5815) );
  OR2_X1 U5192 ( .A1(n9030), .A2(n8823), .ZN(n5713) );
  NOR2_X1 U5193 ( .A1(n5067), .A2(n5074), .ZN(n5062) );
  OR2_X1 U5194 ( .A1(n9047), .A2(n8860), .ZN(n5075) );
  INV_X1 U5195 ( .A(n5897), .ZN(n4830) );
  INV_X1 U5196 ( .A(n8909), .ZN(n5034) );
  OR2_X1 U5197 ( .A1(n8922), .A2(n5545), .ZN(n5037) );
  INV_X1 U5198 ( .A(n5779), .ZN(n5043) );
  OR2_X1 U5199 ( .A1(n9080), .A2(n8604), .ZN(n5882) );
  AND2_X1 U5200 ( .A1(n5666), .A2(n4464), .ZN(n4836) );
  AND2_X1 U5201 ( .A1(n5095), .A2(n5077), .ZN(n4464) );
  AND2_X1 U5202 ( .A1(n5252), .A2(n4877), .ZN(n4705) );
  INV_X1 U5203 ( .A(n7047), .ZN(n4613) );
  NAND2_X1 U5204 ( .A1(n4621), .A2(n4801), .ZN(n6203) );
  AND2_X1 U5205 ( .A1(n4802), .A2(n7440), .ZN(n4801) );
  NAND2_X1 U5206 ( .A1(n4803), .A2(n7439), .ZN(n4802) );
  AND2_X1 U5207 ( .A1(n7756), .A2(n7699), .ZN(n4779) );
  NOR2_X1 U5208 ( .A1(n6523), .A2(n6503), .ZN(n4634) );
  NAND2_X1 U5209 ( .A1(n6371), .A2(n6370), .ZN(n9181) );
  OR2_X1 U5210 ( .A1(n9725), .A2(n9172), .ZN(n8340) );
  OR2_X1 U5211 ( .A1(n8186), .A2(n9250), .ZN(n8343) );
  INV_X1 U5212 ( .A(n6089), .ZN(n6542) );
  NOR2_X1 U5213 ( .A1(n9606), .A2(n8228), .ZN(n8250) );
  NAND2_X1 U5214 ( .A1(n7856), .A2(n8236), .ZN(n7857) );
  NOR2_X1 U5215 ( .A1(n7864), .A2(n7909), .ZN(n4770) );
  OR2_X1 U5216 ( .A1(n7864), .A2(n7863), .ZN(n8236) );
  NAND2_X1 U5217 ( .A1(n6212), .A2(n4695), .ZN(n8224) );
  NOR2_X1 U5218 ( .A1(n7672), .A2(n4696), .ZN(n4695) );
  INV_X1 U5219 ( .A(n6211), .ZN(n4696) );
  OR2_X1 U5220 ( .A1(n9716), .A2(n9173), .ZN(n8345) );
  NAND2_X1 U5221 ( .A1(n9731), .A2(n8164), .ZN(n4951) );
  INV_X1 U5222 ( .A(n6008), .ZN(n4783) );
  AOI21_X1 U5223 ( .B1(n4990), .B2(n4993), .A(n4989), .ZN(n4988) );
  AND2_X1 U5224 ( .A1(n5215), .A2(n5214), .ZN(n5624) );
  AND2_X1 U5225 ( .A1(n5209), .A2(n5208), .ZN(n5615) );
  NAND2_X1 U5226 ( .A1(n6027), .A2(n4785), .ZN(n6038) );
  AND2_X1 U5227 ( .A1(n5202), .A2(n5201), .ZN(n5233) );
  INV_X1 U5228 ( .A(n5532), .ZN(n5173) );
  OAI21_X1 U5229 ( .B1(n5518), .B2(n5517), .A(n5169), .ZN(n5533) );
  NAND2_X1 U5230 ( .A1(n5454), .A2(n4354), .ZN(n5456) );
  AND2_X1 U5231 ( .A1(n5150), .A2(n5398), .ZN(n5151) );
  OAI21_X1 U5232 ( .B1(n5338), .B2(n4686), .A(n4651), .ZN(n4445) );
  AOI21_X1 U5233 ( .B1(n4974), .B2(n4687), .A(n4388), .ZN(n4651) );
  NAND2_X1 U5234 ( .A1(n5132), .A2(n4687), .ZN(n4686) );
  INV_X1 U5235 ( .A(n4445), .ZN(n4981) );
  OAI21_X1 U5236 ( .B1(n6661), .B2(n4573), .A(n4572), .ZN(n5129) );
  NAND2_X1 U5237 ( .A1(n6661), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n4572) );
  OAI21_X1 U5238 ( .B1(n5111), .B2(n5113), .A(n5112), .ZN(n5116) );
  NAND2_X1 U5239 ( .A1(n5101), .A2(SI_1_), .ZN(n5107) );
  NAND2_X1 U5240 ( .A1(n8597), .A2(n8482), .ZN(n8487) );
  OR2_X1 U5241 ( .A1(n8492), .A2(n4540), .ZN(n4539) );
  INV_X1 U5242 ( .A(n8490), .ZN(n4540) );
  XNOR2_X1 U5243 ( .A(n8808), .B(n8491), .ZN(n8492) );
  AND2_X1 U5244 ( .A1(n4911), .A2(n4557), .ZN(n4556) );
  NAND2_X1 U5245 ( .A1(n4559), .A2(n8476), .ZN(n4557) );
  AND2_X1 U5246 ( .A1(n8561), .A2(n4912), .ZN(n4911) );
  NAND2_X1 U5247 ( .A1(n4556), .A2(n4558), .ZN(n4554) );
  NAND2_X1 U5248 ( .A1(n4920), .A2(n4924), .ZN(n4919) );
  INV_X1 U5249 ( .A(n4922), .ZN(n4920) );
  AND2_X1 U5250 ( .A1(n7973), .A2(n4924), .ZN(n4921) );
  NOR2_X1 U5251 ( .A1(n8554), .A2(n4546), .ZN(n4545) );
  INV_X1 U5252 ( .A(n4551), .ZN(n4546) );
  OR2_X1 U5253 ( .A1(n8511), .A2(n8868), .ZN(n4912) );
  AND2_X1 U5254 ( .A1(n8511), .A2(n8868), .ZN(n4913) );
  XNOR2_X1 U5255 ( .A(n4329), .B(n7190), .ZN(n7105) );
  AOI21_X1 U5256 ( .B1(n4914), .B2(n4531), .A(n4348), .ZN(n4530) );
  INV_X1 U5257 ( .A(n4914), .ZN(n4535) );
  INV_X1 U5258 ( .A(n7173), .ZN(n4531) );
  OR2_X1 U5259 ( .A1(n7806), .A2(n7769), .ZN(n4569) );
  NOR2_X1 U5260 ( .A1(n5985), .A2(n7061), .ZN(n6931) );
  INV_X1 U5261 ( .A(n5949), .ZN(n4710) );
  INV_X1 U5262 ( .A(n5950), .ZN(n4712) );
  NAND2_X1 U5263 ( .A1(n4844), .A2(n4843), .ZN(n4842) );
  NAND2_X1 U5264 ( .A1(n5799), .A2(n5980), .ZN(n4841) );
  AOI21_X1 U5265 ( .B1(n5797), .B2(n9010), .A(n5980), .ZN(n4843) );
  OAI21_X1 U5266 ( .B1(n8643), .B2(P2_REG2_REG_0__SCAN_IN), .A(n4462), .ZN(
        n4461) );
  NAND2_X1 U5267 ( .A1(n8643), .A2(n6704), .ZN(n4462) );
  OAI21_X1 U5268 ( .B1(n4602), .B2(P2_REG1_REG_2__SCAN_IN), .A(n4447), .ZN(
        n9904) );
  NAND2_X1 U5269 ( .A1(n4602), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4447) );
  NOR2_X1 U5270 ( .A1(n6722), .A2(n6723), .ZN(n4455) );
  OR2_X1 U5271 ( .A1(n9936), .A2(n7310), .ZN(n4488) );
  OAI211_X1 U5272 ( .C1(n9957), .C2(n4668), .A(n4665), .B(n4664), .ZN(n9979)
         );
  NAND2_X1 U5273 ( .A1(n4671), .A2(n7341), .ZN(n4668) );
  INV_X1 U5274 ( .A(n4666), .ZN(n4665) );
  NAND2_X1 U5275 ( .A1(n9957), .A2(n4669), .ZN(n4664) );
  NOR2_X1 U5276 ( .A1(n9963), .A2(n4460), .ZN(n9990) );
  AND2_X1 U5277 ( .A1(n7324), .A2(n7325), .ZN(n4460) );
  NOR2_X1 U5278 ( .A1(n9979), .A2(n7376), .ZN(n9978) );
  NAND2_X1 U5279 ( .A1(n4663), .A2(n4671), .ZN(n9954) );
  INV_X1 U5280 ( .A(n9957), .ZN(n4663) );
  NAND2_X1 U5281 ( .A1(n4599), .A2(n4366), .ZN(n4873) );
  NAND3_X1 U5282 ( .A1(n4672), .A2(n4676), .A3(n4673), .ZN(n4889) );
  AND2_X1 U5283 ( .A1(n4674), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4673) );
  NAND2_X1 U5284 ( .A1(n4597), .A2(n4360), .ZN(n4871) );
  NAND2_X1 U5285 ( .A1(n4871), .A2(n4870), .ZN(n7737) );
  INV_X1 U5286 ( .A(n7424), .ZN(n4870) );
  NAND2_X1 U5287 ( .A1(n7740), .A2(n7741), .ZN(n7742) );
  NAND2_X1 U5288 ( .A1(n7742), .A2(n7743), .ZN(n7847) );
  OR2_X1 U5289 ( .A1(n7839), .A2(n7838), .ZN(n4876) );
  NAND2_X1 U5290 ( .A1(n7747), .A2(n7746), .ZN(n7824) );
  NAND2_X1 U5291 ( .A1(n4876), .A2(n4875), .ZN(n4874) );
  NAND2_X1 U5292 ( .A1(n7949), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4875) );
  INV_X1 U5293 ( .A(n4902), .ZN(n8654) );
  OR2_X1 U5294 ( .A1(n8660), .A2(n8659), .ZN(n4452) );
  NOR2_X1 U5295 ( .A1(n8665), .A2(n4422), .ZN(n8698) );
  XNOR2_X1 U5296 ( .A(n8687), .B(n8699), .ZN(n8682) );
  NOR2_X1 U5297 ( .A1(n8693), .A2(n8694), .ZN(n8714) );
  AND2_X1 U5298 ( .A1(n4486), .A2(n4427), .ZN(n8729) );
  OR2_X1 U5299 ( .A1(n8711), .A2(n4866), .ZN(n4864) );
  OR2_X1 U5300 ( .A1(n8731), .A2(n9002), .ZN(n4866) );
  OR2_X1 U5301 ( .A1(n4353), .A2(n8731), .ZN(n4865) );
  NAND2_X1 U5302 ( .A1(n8805), .A2(n5796), .ZN(n5965) );
  AOI21_X1 U5303 ( .B1(n4858), .B2(n4860), .A(n4857), .ZN(n4856) );
  OR2_X1 U5304 ( .A1(n5649), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8781) );
  AND2_X1 U5305 ( .A1(n5790), .A2(n5789), .ZN(n5958) );
  OR2_X1 U5306 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n5606), .ZN(n5079) );
  NOR2_X2 U5307 ( .A1(n5079), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5628) );
  NAND2_X1 U5308 ( .A1(n5072), .A2(n5076), .ZN(n5071) );
  NAND2_X1 U5309 ( .A1(n7815), .A2(n5778), .ZN(n5702) );
  OAI21_X1 U5310 ( .B1(n7616), .B2(n5394), .A(n5038), .ZN(n7727) );
  OR2_X1 U5311 ( .A1(n10062), .A2(n8628), .ZN(n5038) );
  NOR2_X2 U5312 ( .A1(n5350), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5371) );
  NAND2_X1 U5313 ( .A1(n5698), .A2(n7065), .ZN(n7016) );
  INV_X1 U5314 ( .A(n8952), .ZN(n10026) );
  NAND2_X1 U5315 ( .A1(n5004), .A2(n5759), .ZN(n5973) );
  AOI21_X1 U5316 ( .B1(n4859), .B2(n4861), .A(n4383), .ZN(n4858) );
  INV_X1 U5317 ( .A(n4863), .ZN(n4859) );
  INV_X1 U5318 ( .A(n4861), .ZN(n4860) );
  NOR2_X1 U5319 ( .A1(n5926), .A2(n5912), .ZN(n4863) );
  AND2_X1 U5320 ( .A1(n5713), .A2(n5924), .ZN(n8831) );
  OR2_X1 U5321 ( .A1(n8856), .A2(n5711), .ZN(n8842) );
  NOR2_X1 U5322 ( .A1(n8870), .A2(n5069), .ZN(n5068) );
  INV_X1 U5323 ( .A(n5071), .ZN(n5069) );
  INV_X1 U5324 ( .A(n5075), .ZN(n5064) );
  AOI21_X1 U5325 ( .B1(n5910), .B2(n4833), .A(n4832), .ZN(n4831) );
  INV_X1 U5326 ( .A(n5890), .ZN(n4833) );
  INV_X1 U5327 ( .A(n5893), .ZN(n4832) );
  AND2_X1 U5328 ( .A1(n5894), .A2(n5897), .ZN(n8870) );
  AND3_X1 U5329 ( .A1(n5587), .A2(n5586), .A3(n5585), .ZN(n8893) );
  NAND2_X1 U5330 ( .A1(n5710), .A2(n5907), .ZN(n8888) );
  NAND2_X1 U5331 ( .A1(n8920), .A2(n4346), .ZN(n5710) );
  NAND2_X1 U5332 ( .A1(n5709), .A2(n4853), .ZN(n8920) );
  NOR2_X1 U5333 ( .A1(n8921), .A2(n4854), .ZN(n4853) );
  INV_X1 U5334 ( .A(n5901), .ZN(n4854) );
  OR2_X1 U5335 ( .A1(n8931), .A2(n8903), .ZN(n5904) );
  AND2_X1 U5336 ( .A1(n5903), .A2(n5907), .ZN(n8909) );
  INV_X1 U5337 ( .A(n8949), .ZN(n10030) );
  NAND2_X1 U5338 ( .A1(n5553), .A2(n5552), .ZN(n8520) );
  NAND2_X1 U5339 ( .A1(n8037), .A2(n5801), .ZN(n5707) );
  AOI21_X1 U5340 ( .B1(n5046), .B2(n5045), .A(n4380), .ZN(n5044) );
  INV_X1 U5341 ( .A(n5050), .ZN(n5045) );
  INV_X1 U5342 ( .A(n5877), .ZN(n8036) );
  NAND2_X1 U5343 ( .A1(n5049), .A2(n5769), .ZN(n7989) );
  NAND2_X1 U5344 ( .A1(n5453), .A2(n5050), .ZN(n5049) );
  INV_X1 U5345 ( .A(n5704), .ZN(n4840) );
  NAND2_X1 U5346 ( .A1(n5704), .A2(n4839), .ZN(n4838) );
  INV_X1 U5347 ( .A(n5862), .ZN(n4839) );
  AND2_X1 U5348 ( .A1(n10051), .A2(n10063), .ZN(n10068) );
  INV_X1 U5349 ( .A(n5238), .ZN(n9090) );
  AOI21_X1 U5350 ( .B1(n5237), .B2(n4377), .A(n4827), .ZN(n4826) );
  NOR2_X1 U5351 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n4827) );
  NAND2_X1 U5352 ( .A1(n4596), .A2(n4593), .ZN(n6702) );
  NOR2_X1 U5353 ( .A1(n4595), .A2(n4594), .ZN(n4593) );
  OR2_X1 U5354 ( .A1(n5229), .A2(n10246), .ZN(n4596) );
  NOR2_X1 U5355 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4594) );
  XNOR2_X1 U5356 ( .A(n5663), .B(n5662), .ZN(n6922) );
  INV_X1 U5357 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5662) );
  OAI21_X1 U5358 ( .B1(n5661), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5663) );
  OAI21_X1 U5359 ( .B1(n5504), .B2(n4904), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5644) );
  AND2_X1 U5360 ( .A1(n5422), .A2(n5457), .ZN(n7834) );
  INV_X1 U5361 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U5362 ( .A1(n5089), .A2(n6333), .ZN(n4618) );
  NAND2_X1 U5363 ( .A1(n4793), .A2(n4619), .ZN(n5089) );
  NOR2_X1 U5364 ( .A1(n4620), .A2(n6329), .ZN(n4619) );
  INV_X1 U5365 ( .A(n4364), .ZN(n4620) );
  OR2_X1 U5366 ( .A1(n6506), .A2(n8457), .ZN(n6526) );
  INV_X1 U5367 ( .A(n7294), .ZN(n4615) );
  INV_X1 U5368 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6233) );
  AND2_X1 U5369 ( .A1(n4633), .A2(n4631), .ZN(n4630) );
  INV_X1 U5370 ( .A(n9170), .ZN(n4631) );
  INV_X1 U5371 ( .A(n8439), .ZN(n4737) );
  NAND2_X1 U5372 ( .A1(n6941), .A2(n6942), .ZN(n6940) );
  AOI21_X1 U5373 ( .B1(n6960), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6954), .ZN(
        n6955) );
  NAND2_X1 U5374 ( .A1(n6955), .A2(n6956), .ZN(n7083) );
  OR2_X1 U5375 ( .A1(n7084), .A2(n7085), .ZN(n4514) );
  NOR2_X1 U5376 ( .A1(n8158), .A2(n4932), .ZN(n4931) );
  INV_X1 U5377 ( .A(n8155), .ZN(n4932) );
  NAND2_X1 U5378 ( .A1(n8334), .A2(n4339), .ZN(n4930) );
  OAI21_X1 U5379 ( .B1(n4927), .B2(n4933), .A(n4926), .ZN(n4925) );
  NAND2_X1 U5380 ( .A1(n4933), .A2(n4339), .ZN(n4926) );
  NAND2_X1 U5381 ( .A1(n4702), .A2(n4341), .ZN(n9381) );
  NAND2_X1 U5382 ( .A1(n4703), .A2(n8346), .ZN(n4702) );
  NAND2_X1 U5383 ( .A1(n9428), .A2(n9413), .ZN(n9412) );
  INV_X1 U5384 ( .A(n8196), .ZN(n4704) );
  NAND2_X1 U5385 ( .A1(n4949), .A2(n8149), .ZN(n4948) );
  INV_X1 U5386 ( .A(n4953), .ZN(n4949) );
  NAND2_X1 U5387 ( .A1(n9734), .A2(n9276), .ZN(n4952) );
  AND2_X1 U5388 ( .A1(n8197), .A2(n8196), .ZN(n9456) );
  NAND2_X1 U5389 ( .A1(n6476), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6493) );
  NOR2_X1 U5390 ( .A1(n9751), .A2(n9522), .ZN(n8147) );
  OR2_X1 U5391 ( .A1(n9548), .A2(n9137), .ZN(n5080) );
  NOR2_X1 U5392 ( .A1(n9554), .A2(n4814), .ZN(n4813) );
  INV_X1 U5393 ( .A(n8417), .ZN(n4814) );
  OR2_X1 U5394 ( .A1(n9770), .A2(n8167), .ZN(n9586) );
  NAND2_X1 U5395 ( .A1(n7911), .A2(n7910), .ZN(n7912) );
  NAND2_X1 U5396 ( .A1(n8408), .A2(n9604), .ZN(n8324) );
  NAND2_X1 U5397 ( .A1(n7783), .A2(n7782), .ZN(n7785) );
  OR2_X1 U5398 ( .A1(n9128), .A2(n9286), .ZN(n7782) );
  NAND2_X1 U5399 ( .A1(n7520), .A2(n7569), .ZN(n7567) );
  AND4_X1 U5400 ( .A1(n6146), .A2(n6145), .A3(n6144), .A4(n6143), .ZN(n7506)
         );
  INV_X1 U5401 ( .A(n7216), .ZN(n4492) );
  AOI21_X1 U5402 ( .B1(n4491), .B2(n7216), .A(n4490), .ZN(n4489) );
  INV_X1 U5403 ( .A(n8308), .ZN(n4491) );
  NAND2_X1 U5404 ( .A1(n4946), .A2(n4951), .ZN(n4945) );
  INV_X1 U5405 ( .A(n4948), .ZN(n4946) );
  NAND2_X1 U5406 ( .A1(n6490), .A2(n6489), .ZN(n9462) );
  NAND2_X1 U5407 ( .A1(n9504), .A2(n4968), .ZN(n4507) );
  OR2_X1 U5408 ( .A1(n9744), .A2(n9525), .ZN(n4968) );
  NAND2_X1 U5409 ( .A1(n6379), .A2(n6378), .ZN(n9561) );
  NAND2_X1 U5410 ( .A1(n7912), .A2(n8324), .ZN(n8140) );
  NAND2_X1 U5411 ( .A1(n7220), .A2(n8306), .ZN(n7508) );
  XNOR2_X1 U5412 ( .A(n9293), .B(n7247), .ZN(n8308) );
  NAND2_X1 U5413 ( .A1(n6594), .A2(n6606), .ZN(n6886) );
  XNOR2_X1 U5414 ( .A(n5742), .B(n5741), .ZN(n9085) );
  NAND2_X1 U5415 ( .A1(n5738), .A2(n5737), .ZN(n5742) );
  OAI21_X1 U5416 ( .B1(n6008), .B2(n4935), .A(n4390), .ZN(n4934) );
  NAND2_X1 U5417 ( .A1(n4936), .A2(n6010), .ZN(n4935) );
  INV_X1 U5418 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4936) );
  XNOR2_X1 U5419 ( .A(n5750), .B(n5749), .ZN(n8498) );
  INV_X1 U5420 ( .A(n6031), .ZN(n6007) );
  XNOR2_X1 U5421 ( .A(n5720), .B(n5719), .ZN(n9099) );
  XNOR2_X1 U5422 ( .A(n4437), .B(n5624), .ZN(n8043) );
  OAI21_X1 U5423 ( .B1(n5203), .B2(n4993), .A(n4990), .ZN(n4437) );
  XNOR2_X1 U5424 ( .A(n5232), .B(n5233), .ZN(n7982) );
  NOR2_X1 U5425 ( .A1(n5588), .A2(n5001), .ZN(n5000) );
  INV_X1 U5426 ( .A(n5183), .ZN(n5001) );
  AOI21_X1 U5427 ( .B1(n5000), .B2(n5184), .A(n4999), .ZN(n4998) );
  INV_X1 U5428 ( .A(n5190), .ZN(n4999) );
  OAI21_X1 U5429 ( .B1(n5579), .B2(n5184), .A(n5183), .ZN(n5589) );
  NAND2_X1 U5430 ( .A1(n4435), .A2(n4641), .ZN(n5565) );
  INV_X1 U5431 ( .A(n4643), .ZN(n4641) );
  XNOR2_X1 U5432 ( .A(n5500), .B(n5502), .ZN(n7245) );
  AOI21_X1 U5433 ( .B1(n4982), .B2(n4978), .A(n4350), .ZN(n4977) );
  INV_X1 U5434 ( .A(SI_11_), .ZN(n4984) );
  NAND2_X1 U5435 ( .A1(n4445), .A2(n4978), .ZN(n4976) );
  OAI21_X1 U5436 ( .B1(n5338), .B2(n4975), .A(n4973), .ZN(n5357) );
  INV_X1 U5437 ( .A(n4974), .ZN(n4973) );
  NAND2_X1 U5438 ( .A1(n5291), .A2(n5118), .ZN(n5307) );
  NAND2_X1 U5439 ( .A1(n5307), .A2(n5306), .ZN(n5309) );
  NAND2_X1 U5440 ( .A1(n5289), .A2(n5288), .ZN(n5291) );
  INV_X1 U5441 ( .A(n8859), .ZN(n8516) );
  AOI21_X1 U5442 ( .B1(n8579), .B2(n8578), .A(n4558), .ZN(n4555) );
  AND3_X1 U5443 ( .A1(n5573), .A2(n5572), .A3(n5571), .ZN(n8904) );
  NAND2_X1 U5444 ( .A1(n7005), .A2(n7004), .ZN(n7026) );
  NAND2_X1 U5445 ( .A1(n5613), .A2(n5612), .ZN(n8848) );
  INV_X1 U5446 ( .A(n8877), .ZN(n8860) );
  NAND2_X1 U5447 ( .A1(n4885), .A2(n4884), .ZN(n9996) );
  AND2_X1 U5448 ( .A1(n5406), .A2(n5421), .ZN(n7429) );
  NOR2_X1 U5449 ( .A1(n7738), .A2(n5425), .ZN(n7835) );
  XNOR2_X1 U5450 ( .A(n4874), .B(n7950), .ZN(n7935) );
  NOR2_X1 U5451 ( .A1(n7935), .A2(n8012), .ZN(n8637) );
  XNOR2_X1 U5452 ( .A(n8698), .B(n8699), .ZN(n8666) );
  OR2_X1 U5453 ( .A1(n8711), .A2(n9002), .ZN(n4867) );
  NAND2_X1 U5454 ( .A1(n4585), .A2(n4582), .ZN(n8752) );
  NOR2_X1 U5455 ( .A1(n4584), .A2(n4583), .ZN(n4582) );
  NAND2_X1 U5456 ( .A1(n8740), .A2(n4586), .ZN(n4585) );
  INV_X1 U5457 ( .A(n8741), .ZN(n4583) );
  NAND2_X1 U5458 ( .A1(n4864), .A2(n4865), .ZN(n8757) );
  NAND2_X1 U5459 ( .A1(n4683), .A2(n10009), .ZN(n4581) );
  XNOR2_X1 U5460 ( .A(n8774), .B(n8775), .ZN(n4683) );
  INV_X1 U5461 ( .A(n8776), .ZN(n4682) );
  AND3_X1 U5462 ( .A1(n4865), .A2(n4864), .A3(n8756), .ZN(n8759) );
  NAND2_X1 U5463 ( .A1(n5970), .A2(n5969), .ZN(n8788) );
  INV_X1 U5464 ( .A(n5968), .ZN(n5969) );
  AOI21_X1 U5465 ( .B1(n8802), .B2(n8952), .A(n8801), .ZN(n8968) );
  NAND2_X1 U5466 ( .A1(n8800), .A2(n8799), .ZN(n8801) );
  NAND2_X1 U5467 ( .A1(n5441), .A2(n5440), .ZN(n10079) );
  OAI21_X1 U5468 ( .B1(n6676), .B2(n5314), .A(n4570), .ZN(n7363) );
  INV_X1 U5469 ( .A(n5346), .ZN(n4570) );
  INV_X1 U5470 ( .A(n10021), .ZN(n8955) );
  INV_X1 U5471 ( .A(n5973), .ZN(n8789) );
  NOR2_X1 U5472 ( .A1(n8788), .A2(n5972), .ZN(n5993) );
  NOR2_X1 U5473 ( .A1(n8795), .A2(n10063), .ZN(n5972) );
  NAND2_X1 U5474 ( .A1(n5603), .A2(n5602), .ZN(n9042) );
  NAND2_X1 U5475 ( .A1(n10081), .A2(n10080), .ZN(n9070) );
  AND3_X1 U5476 ( .A1(n5255), .A2(n4529), .A3(n4528), .ZN(n7101) );
  NAND2_X1 U5477 ( .A1(n5263), .A2(n4376), .ZN(n4529) );
  NAND2_X1 U5478 ( .A1(n5551), .A2(n6807), .ZN(n4528) );
  AND2_X1 U5479 ( .A1(n6606), .A2(n6035), .ZN(n6036) );
  AOI21_X1 U5480 ( .B1(n4363), .B2(n9170), .A(n4819), .ZN(n4816) );
  OR2_X1 U5481 ( .A1(n6642), .A2(n6641), .ZN(n4819) );
  INV_X1 U5482 ( .A(n9725), .ZN(n9445) );
  AOI21_X1 U5483 ( .B1(n9230), .B2(n9229), .A(n9226), .ZN(n9231) );
  NOR2_X2 U5484 ( .A1(n6614), .A2(n6612), .ZN(n9809) );
  NAND3_X1 U5485 ( .A1(n6653), .A2(n6693), .A3(P1_STATE_REG_SCAN_IN), .ZN(
        n8444) );
  NAND4_X1 U5486 ( .A1(n6093), .A2(n6092), .A3(n6091), .A4(n6090), .ZN(n9292)
         );
  AND2_X1 U5487 ( .A1(n6058), .A2(n6061), .ZN(n4808) );
  NAND2_X1 U5488 ( .A1(n6012), .A2(n4748), .ZN(n6058) );
  OR2_X1 U5489 ( .A1(n6849), .A2(n6848), .ZN(n4516) );
  NOR2_X1 U5490 ( .A1(n6827), .A2(n4517), .ZN(n6849) );
  AND2_X1 U5491 ( .A1(n6828), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4517) );
  NOR2_X1 U5492 ( .A1(n7964), .A2(n7965), .ZN(n8105) );
  AND2_X1 U5493 ( .A1(n9325), .A2(n8110), .ZN(n9842) );
  OR2_X1 U5494 ( .A1(n9827), .A2(n6763), .ZN(n9847) );
  OR2_X1 U5495 ( .A1(n9344), .A2(n8115), .ZN(n8117) );
  OR2_X1 U5496 ( .A1(n6577), .A2(n6576), .ZN(n9368) );
  NAND2_X1 U5497 ( .A1(n9392), .A2(n4786), .ZN(n4790) );
  AND2_X1 U5498 ( .A1(n4604), .A2(n9396), .ZN(n4603) );
  INV_X1 U5499 ( .A(n9369), .ZN(n4701) );
  NAND2_X1 U5500 ( .A1(n8162), .A2(n8161), .ZN(n9372) );
  OAI21_X1 U5501 ( .B1(n9380), .B2(n9379), .A(n9378), .ZN(n9710) );
  NAND2_X1 U5502 ( .A1(n9380), .A2(n9379), .ZN(n9378) );
  AOI21_X1 U5503 ( .B1(n9709), .B2(n9769), .A(n4823), .ZN(n4822) );
  NOR2_X1 U5504 ( .A1(n9890), .A2(n4824), .ZN(n4823) );
  INV_X1 U5505 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n4824) );
  AND2_X1 U5506 ( .A1(n9890), .A2(n7135), .ZN(n9769) );
  AND2_X1 U5507 ( .A1(n4764), .A2(n4762), .ZN(n9777) );
  AND2_X1 U5508 ( .A1(n4763), .A2(n6010), .ZN(n4762) );
  NAND2_X1 U5509 ( .A1(n5810), .A2(n6656), .ZN(n4723) );
  NAND2_X1 U5510 ( .A1(n5809), .A2(n5986), .ZN(n4725) );
  NOR2_X1 U5511 ( .A1(n4717), .A2(n4716), .ZN(n4715) );
  INV_X1 U5512 ( .A(n5820), .ZN(n4716) );
  NAND2_X1 U5513 ( .A1(n4746), .A2(n4745), .ZN(n4744) );
  OAI21_X1 U5514 ( .B1(n8206), .B2(n8398), .A(n4334), .ZN(n4747) );
  MUX2_X1 U5515 ( .A(n5848), .B(n5847), .S(n6656), .Z(n5849) );
  NAND2_X1 U5516 ( .A1(n5904), .A2(n5885), .ZN(n4729) );
  AOI21_X1 U5517 ( .B1(n8268), .B2(n8269), .A(n8267), .ZN(n4758) );
  NAND2_X1 U5518 ( .A1(n4653), .A2(n6656), .ZN(n4652) );
  NAND2_X1 U5519 ( .A1(n5916), .A2(n5894), .ZN(n4653) );
  NOR2_X1 U5520 ( .A1(n5891), .A2(n4656), .ZN(n4655) );
  NOR2_X1 U5521 ( .A1(n5897), .A2(n6656), .ZN(n4656) );
  NAND2_X1 U5522 ( .A1(n5892), .A2(n5897), .ZN(n4654) );
  AND2_X1 U5523 ( .A1(n9456), .A2(n8329), .ZN(n4754) );
  AOI21_X1 U5524 ( .B1(n4589), .B2(n4588), .A(n4391), .ZN(n5931) );
  NOR2_X1 U5525 ( .A1(n5921), .A2(n5920), .ZN(n4588) );
  OAI22_X1 U5526 ( .A1(n8381), .A2(n8345), .B1(n8356), .B2(n4334), .ZN(n4740)
         );
  NAND2_X1 U5527 ( .A1(n4738), .A2(n8275), .ZN(n4438) );
  NAND2_X1 U5528 ( .A1(n9897), .A2(n6740), .ZN(n6742) );
  INV_X1 U5529 ( .A(n7336), .ZN(n4895) );
  NOR2_X1 U5530 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n4835) );
  NOR2_X1 U5531 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n5077) );
  INV_X1 U5532 ( .A(n6172), .ZN(n4803) );
  NOR2_X1 U5533 ( .A1(n4804), .A2(n6173), .ZN(n4799) );
  INV_X1 U5534 ( .A(n7439), .ZN(n4804) );
  OR2_X1 U5535 ( .A1(n8279), .A2(n8278), .ZN(n8280) );
  OR2_X1 U5536 ( .A1(n9372), .A2(n8163), .ZN(n8359) );
  NOR2_X1 U5537 ( .A1(n9716), .A2(n9399), .ZN(n4775) );
  NAND2_X1 U5538 ( .A1(n5727), .A2(n5726), .ZN(n5730) );
  INV_X1 U5539 ( .A(n5624), .ZN(n4989) );
  INV_X1 U5540 ( .A(n5577), .ZN(n5182) );
  INV_X1 U5541 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5164) );
  INV_X1 U5542 ( .A(n5136), .ZN(n4688) );
  INV_X1 U5543 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5007) );
  XNOR2_X1 U5544 ( .A(n7378), .B(n8491), .ZN(n7400) );
  NAND2_X1 U5545 ( .A1(n8464), .A2(n8948), .ZN(n4924) );
  NOR2_X1 U5546 ( .A1(n4714), .A2(n4647), .ZN(n4713) );
  NOR2_X1 U5547 ( .A1(n5943), .A2(n5986), .ZN(n4714) );
  INV_X1 U5548 ( .A(n8821), .ZN(n4592) );
  NAND2_X1 U5549 ( .A1(n5252), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6727) );
  OR2_X1 U5550 ( .A1(n6808), .A2(n7019), .ZN(n6810) );
  INV_X1 U5551 ( .A(n4883), .ZN(n4882) );
  INV_X1 U5552 ( .A(n4880), .ZN(n6743) );
  NAND2_X1 U5553 ( .A1(n7338), .A2(n4895), .ZN(n4894) );
  AND2_X1 U5554 ( .A1(n7308), .A2(n4600), .ZN(n7309) );
  NAND2_X1 U5555 ( .A1(n7319), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4600) );
  AND2_X1 U5556 ( .A1(n7340), .A2(n9983), .ZN(n4669) );
  OAI21_X1 U5557 ( .B1(n4671), .B2(n4667), .A(n4670), .ZN(n4666) );
  OR2_X1 U5558 ( .A1(n9983), .A2(n7340), .ZN(n4670) );
  INV_X1 U5559 ( .A(n4669), .ZN(n4667) );
  NAND2_X1 U5560 ( .A1(n4658), .A2(n4423), .ZN(n4902) );
  INV_X1 U5561 ( .A(n8733), .ZN(n8734) );
  INV_X1 U5562 ( .A(n5934), .ZN(n4857) );
  INV_X1 U5563 ( .A(n5843), .ZN(n4851) );
  INV_X1 U5564 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7109) );
  NOR2_X2 U5565 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5316) );
  NAND2_X1 U5566 ( .A1(n6913), .A2(n7020), .ZN(n5807) );
  NAND2_X1 U5567 ( .A1(n9093), .A2(n5787), .ZN(n5004) );
  NOR2_X1 U5568 ( .A1(n5867), .A2(n5051), .ZN(n5050) );
  INV_X1 U5569 ( .A(n5452), .ZN(n5051) );
  NOR2_X2 U5570 ( .A1(n5226), .A2(n5225), .ZN(n5666) );
  INV_X1 U5571 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5222) );
  NAND2_X1 U5572 ( .A1(n4905), .A2(n5096), .ZN(n4904) );
  NOR2_X1 U5573 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5096) );
  INV_X1 U5574 ( .A(n5225), .ZN(n4905) );
  NAND2_X1 U5575 ( .A1(n9217), .A2(n4797), .ZN(n4796) );
  NOR2_X1 U5576 ( .A1(n4798), .A2(n4795), .ZN(n4794) );
  INV_X1 U5577 ( .A(n9162), .ZN(n4795) );
  INV_X1 U5578 ( .A(n9217), .ZN(n4798) );
  NAND2_X1 U5579 ( .A1(n6334), .A2(n4618), .ZN(n6368) );
  AND2_X1 U5580 ( .A1(n6516), .A2(n6515), .ZN(n6518) );
  INV_X1 U5581 ( .A(n6454), .ZN(n4624) );
  XNOR2_X1 U5582 ( .A(n6068), .B(n6546), .ZN(n6070) );
  OR2_X1 U5583 ( .A1(n9198), .A2(n4812), .ZN(n4811) );
  INV_X1 U5584 ( .A(n6394), .ZN(n4812) );
  AND2_X1 U5585 ( .A1(n6394), .A2(n9187), .ZN(n4810) );
  INV_X1 U5586 ( .A(n6157), .ZN(n4972) );
  NOR2_X1 U5587 ( .A1(n9709), .A2(n4774), .ZN(n4773) );
  INV_X1 U5588 ( .A(n4775), .ZN(n4774) );
  AND2_X1 U5589 ( .A1(n4339), .A2(n4928), .ZN(n4927) );
  INV_X1 U5590 ( .A(n4931), .ZN(n4928) );
  INV_X1 U5591 ( .A(n4945), .ZN(n4943) );
  INV_X1 U5592 ( .A(n4944), .ZN(n4941) );
  NOR2_X1 U5593 ( .A1(n4960), .A2(n4956), .ZN(n4955) );
  INV_X1 U5594 ( .A(n8141), .ZN(n4960) );
  INV_X1 U5595 ( .A(n8324), .ZN(n4956) );
  NAND2_X1 U5596 ( .A1(n8141), .A2(n4959), .ZN(n4958) );
  INV_X1 U5597 ( .A(n8139), .ZN(n4959) );
  INV_X1 U5598 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6319) );
  OR2_X1 U5599 ( .A1(n8316), .A2(n7666), .ZN(n7667) );
  INV_X1 U5600 ( .A(n7572), .ZN(n4965) );
  INV_X1 U5601 ( .A(n4963), .ZN(n4503) );
  AOI21_X1 U5602 ( .B1(n7572), .B2(n4964), .A(n4385), .ZN(n4963) );
  INV_X1 U5603 ( .A(n7566), .ZN(n4964) );
  INV_X1 U5604 ( .A(n7519), .ZN(n4504) );
  NAND2_X1 U5605 ( .A1(n7207), .A2(n8386), .ZN(n7235) );
  INV_X1 U5606 ( .A(n8309), .ZN(n4490) );
  INV_X1 U5607 ( .A(n6047), .ZN(n6395) );
  NAND2_X1 U5608 ( .A1(n9290), .A2(n7629), .ZN(n8400) );
  AND2_X1 U5609 ( .A1(n5737), .A2(n5736), .ZN(n5749) );
  XNOR2_X1 U5610 ( .A(n5730), .B(n5729), .ZN(n5758) );
  AND2_X1 U5611 ( .A1(n5721), .A2(n5221), .ZN(n5719) );
  AOI21_X1 U5612 ( .B1(n5615), .B2(n4992), .A(n4991), .ZN(n4990) );
  INV_X1 U5613 ( .A(n5209), .ZN(n4991) );
  INV_X1 U5614 ( .A(n5202), .ZN(n4992) );
  INV_X1 U5615 ( .A(n5615), .ZN(n4993) );
  NOR2_X1 U5616 ( .A1(n4643), .A2(n5562), .ZN(n4642) );
  NAND2_X1 U5617 ( .A1(n6038), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6040) );
  INV_X1 U5618 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6020) );
  NAND2_X1 U5619 ( .A1(n4644), .A2(n5179), .ZN(n4643) );
  NAND2_X1 U5620 ( .A1(n4645), .A2(n5173), .ZN(n4644) );
  NAND2_X1 U5621 ( .A1(n5533), .A2(n4645), .ZN(n4435) );
  NAND2_X1 U5622 ( .A1(n6043), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6408) );
  INV_X1 U5623 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6407) );
  INV_X1 U5624 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5161) );
  NAND2_X1 U5625 ( .A1(n4430), .A2(n5160), .ZN(n4429) );
  NAND2_X1 U5626 ( .A1(n4431), .A2(n5010), .ZN(n4430) );
  INV_X1 U5627 ( .A(n5152), .ZN(n4985) );
  NOR2_X2 U5628 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6079) );
  AND2_X1 U5629 ( .A1(n7259), .A2(n7257), .ZN(n4914) );
  INV_X1 U5630 ( .A(n8501), .ZN(n4899) );
  NAND2_X1 U5631 ( .A1(n8465), .A2(n8938), .ZN(n4551) );
  NAND2_X1 U5632 ( .A1(n4918), .A2(n4548), .ZN(n4547) );
  INV_X1 U5633 ( .A(n8530), .ZN(n4563) );
  AOI21_X1 U5634 ( .B1(n4906), .B2(n8521), .A(n4344), .ZN(n4564) );
  INV_X1 U5635 ( .A(n4906), .ZN(n4565) );
  NAND2_X1 U5636 ( .A1(n4566), .A2(n7819), .ZN(n7767) );
  INV_X1 U5637 ( .A(n7591), .ZN(n4566) );
  AND2_X1 U5638 ( .A1(n6973), .A2(n6970), .ZN(n4526) );
  NAND2_X1 U5639 ( .A1(n4550), .A2(n8586), .ZN(n8585) );
  INV_X1 U5640 ( .A(n4543), .ZN(n4542) );
  OAI21_X1 U5641 ( .B1(n4548), .B2(n4544), .A(n8467), .ZN(n4543) );
  XNOR2_X1 U5642 ( .A(n7363), .B(n4329), .ZN(n7255) );
  NOR2_X1 U5643 ( .A1(n4923), .A2(n8612), .ZN(n4922) );
  INV_X1 U5644 ( .A(n8462), .ZN(n4923) );
  OR2_X1 U5645 ( .A1(n8461), .A2(n8623), .ZN(n8462) );
  NAND2_X1 U5646 ( .A1(n7974), .A2(n7973), .ZN(n8463) );
  INV_X1 U5647 ( .A(n6973), .ZN(n4639) );
  AND4_X1 U5648 ( .A1(n5767), .A2(n5766), .A3(n5765), .A4(n5764), .ZN(n8619)
         );
  NAND2_X1 U5649 ( .A1(n4661), .A2(n4659), .ZN(n6813) );
  NOR2_X1 U5650 ( .A1(n4660), .A2(n7100), .ZN(n4659) );
  INV_X1 U5651 ( .A(n6738), .ZN(n4660) );
  NAND2_X1 U5652 ( .A1(n4661), .A2(n6738), .ZN(n4662) );
  NAND2_X1 U5653 ( .A1(n6810), .A2(n6727), .ZN(n9903) );
  NAND2_X1 U5654 ( .A1(n6813), .A2(n6738), .ZN(n9898) );
  NAND2_X1 U5655 ( .A1(n9898), .A2(n9899), .ZN(n9897) );
  OR2_X1 U5656 ( .A1(n4882), .A2(n6743), .ZN(n9920) );
  NOR2_X1 U5657 ( .A1(n6743), .A2(n4881), .ZN(n9919) );
  INV_X1 U5658 ( .A(n4483), .ZN(n4480) );
  INV_X1 U5659 ( .A(n4685), .ZN(n6746) );
  NAND2_X1 U5660 ( .A1(n4449), .A2(n6729), .ZN(n7308) );
  NAND2_X1 U5661 ( .A1(n6730), .A2(n6732), .ZN(n4449) );
  NOR2_X1 U5662 ( .A1(n4454), .A2(n6744), .ZN(n4453) );
  INV_X1 U5663 ( .A(n7320), .ZN(n4454) );
  AND2_X1 U5664 ( .A1(n4897), .A2(n4896), .ZN(n9957) );
  AOI21_X1 U5665 ( .B1(n7337), .B2(n7336), .A(n9939), .ZN(n7339) );
  AND2_X1 U5666 ( .A1(n4459), .A2(n4458), .ZN(n10012) );
  NAND2_X1 U5667 ( .A1(n7326), .A2(n9983), .ZN(n4458) );
  NOR2_X1 U5668 ( .A1(n10012), .A2(n10011), .ZN(n10010) );
  NAND2_X1 U5669 ( .A1(n9996), .A2(n4410), .ZN(n4676) );
  OR2_X1 U5670 ( .A1(n9996), .A2(n7421), .ZN(n4672) );
  NAND2_X1 U5671 ( .A1(n4675), .A2(n7330), .ZN(n4674) );
  INV_X1 U5672 ( .A(n7345), .ZN(n4675) );
  AND2_X1 U5673 ( .A1(n9997), .A2(n7315), .ZN(n7420) );
  NAND2_X1 U5674 ( .A1(n7417), .A2(n7416), .ZN(n7740) );
  NAND2_X1 U5675 ( .A1(n4886), .A2(n4889), .ZN(n4888) );
  INV_X1 U5676 ( .A(n7408), .ZN(n4886) );
  AOI21_X1 U5677 ( .B1(n9996), .B2(n7345), .A(n7421), .ZN(n7408) );
  NAND2_X1 U5678 ( .A1(n7737), .A2(n7736), .ZN(n7832) );
  NAND2_X1 U5679 ( .A1(n7847), .A2(n7848), .ZN(n7939) );
  XNOR2_X1 U5680 ( .A(n4902), .B(n7950), .ZN(n7951) );
  NAND2_X1 U5681 ( .A1(n4450), .A2(n4425), .ZN(n4677) );
  INV_X1 U5682 ( .A(n8682), .ZN(n4450) );
  NAND2_X1 U5683 ( .A1(n8689), .A2(n4679), .ZN(n4678) );
  INV_X1 U5684 ( .A(n8691), .ZN(n4679) );
  OAI21_X1 U5685 ( .B1(n8714), .B2(n8715), .A(n8713), .ZN(n8717) );
  NAND2_X1 U5686 ( .A1(n8717), .A2(n8716), .ZN(n8733) );
  AND2_X1 U5687 ( .A1(n9949), .A2(n8747), .ZN(n4586) );
  NOR2_X1 U5688 ( .A1(n10017), .A2(n8742), .ZN(n4584) );
  NOR2_X1 U5689 ( .A1(n8722), .A2(n8941), .ZN(n8746) );
  OAI21_X1 U5690 ( .B1(n5504), .B2(n5225), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5535) );
  OAI21_X1 U5691 ( .B1(n8722), .B2(n4916), .A(n4915), .ZN(n8773) );
  NAND2_X1 U5692 ( .A1(n4917), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4916) );
  NAND2_X1 U5693 ( .A1(n8745), .A2(n4917), .ZN(n4915) );
  INV_X1 U5694 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8770) );
  NOR2_X1 U5695 ( .A1(n8737), .A2(n8736), .ZN(n8760) );
  OAI21_X1 U5696 ( .B1(n5025), .B2(n5023), .A(n5020), .ZN(n5962) );
  NAND2_X1 U5697 ( .A1(n5026), .A2(n5960), .ZN(n5023) );
  INV_X1 U5698 ( .A(n5021), .ZN(n5020) );
  OAI21_X1 U5699 ( .B1(n8795), .B2(n10051), .A(n5967), .ZN(n5968) );
  NAND2_X1 U5700 ( .A1(n4472), .A2(n4591), .ZN(n8805) );
  INV_X1 U5701 ( .A(n8807), .ZN(n4472) );
  OAI21_X1 U5702 ( .B1(n5025), .B2(n5027), .A(n5024), .ZN(n8796) );
  OR2_X1 U5703 ( .A1(n5604), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5606) );
  OR2_X1 U5704 ( .A1(n5592), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5604) );
  INV_X1 U5705 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U5706 ( .A1(n5583), .A2(n5582), .ZN(n5592) );
  AND2_X1 U5707 ( .A1(n5569), .A2(n5568), .ZN(n5583) );
  INV_X1 U5708 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5523) );
  NAND2_X1 U5709 ( .A1(n5524), .A2(n5523), .ZN(n5539) );
  INV_X1 U5710 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5508) );
  AND2_X1 U5711 ( .A1(n5509), .A2(n5508), .ZN(n5524) );
  AND4_X1 U5712 ( .A1(n5432), .A2(n5431), .A3(n5430), .A4(n5429), .ZN(n7894)
         );
  OR2_X1 U5713 ( .A1(n5426), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5443) );
  NAND2_X1 U5714 ( .A1(n4469), .A2(n5853), .ZN(n7815) );
  OAI21_X1 U5715 ( .B1(n7366), .B2(n4849), .A(n4846), .ZN(n4469) );
  INV_X1 U5716 ( .A(n4850), .ZN(n4849) );
  AND2_X1 U5717 ( .A1(n4847), .A2(n5841), .ZN(n4846) );
  OAI21_X1 U5718 ( .B1(n7727), .B2(n5416), .A(n5417), .ZN(n7817) );
  OR2_X1 U5719 ( .A1(n5409), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5426) );
  AND2_X1 U5720 ( .A1(n5852), .A2(n5853), .ZN(n7726) );
  AND2_X1 U5721 ( .A1(n5371), .A2(n5370), .ZN(n5386) );
  INV_X1 U5722 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U5723 ( .A1(n5386), .A2(n5385), .ZN(n5409) );
  NAND2_X1 U5724 ( .A1(n7366), .A2(n5837), .ZN(n4852) );
  NAND2_X1 U5725 ( .A1(n4852), .A2(n4850), .ZN(n7724) );
  OAI21_X1 U5726 ( .B1(n7493), .B2(n5379), .A(n5378), .ZN(n7616) );
  AND4_X1 U5727 ( .A1(n5355), .A2(n5354), .A3(n5353), .A4(n5352), .ZN(n7495)
         );
  AND2_X1 U5728 ( .A1(n5056), .A2(n5058), .ZN(n5055) );
  AOI22_X1 U5729 ( .A1(n5059), .A2(n5315), .B1(n5054), .B2(n5053), .ZN(n5052)
         );
  NAND2_X1 U5730 ( .A1(n5297), .A2(n5315), .ZN(n5056) );
  OR2_X1 U5731 ( .A1(n5301), .A2(n5267), .ZN(n5269) );
  AND2_X1 U5732 ( .A1(n5824), .A2(n5819), .ZN(n7071) );
  NAND2_X1 U5733 ( .A1(n7014), .A2(n5806), .ZN(n10020) );
  NAND2_X1 U5734 ( .A1(n5807), .A2(n5806), .ZN(n5770) );
  OR2_X1 U5735 ( .A1(n5770), .A2(n7016), .ZN(n7014) );
  AND4_X1 U5736 ( .A1(n5019), .A2(n5018), .A3(n5017), .A4(n5016), .ZN(n10027)
         );
  AND4_X1 U5737 ( .A1(n5643), .A2(n5642), .A3(n5641), .A4(n5640), .ZN(n8824)
         );
  OAI21_X1 U5738 ( .B1(n6972), .B2(n5695), .A(n5694), .ZN(n7057) );
  AND2_X1 U5739 ( .A1(n8780), .A2(n8779), .ZN(n9011) );
  INV_X1 U5740 ( .A(n5066), .ZN(n5065) );
  OAI22_X1 U5741 ( .A1(n5068), .A2(n5067), .B1(n8477), .B2(n8868), .ZN(n5066)
         );
  NAND2_X1 U5742 ( .A1(n4470), .A2(n5894), .ZN(n8856) );
  NAND2_X1 U5743 ( .A1(n4828), .A2(n4829), .ZN(n4470) );
  AOI21_X1 U5744 ( .B1(n4831), .B2(n5895), .A(n4830), .ZN(n4829) );
  NAND2_X1 U5745 ( .A1(n5032), .A2(n5033), .ZN(n8890) );
  AOI21_X1 U5746 ( .B1(n4340), .B2(n5545), .A(n4384), .ZN(n5033) );
  AND2_X1 U5747 ( .A1(n5890), .A2(n8880), .ZN(n8889) );
  NAND2_X1 U5748 ( .A1(n5037), .A2(n5035), .ZN(n8900) );
  NAND2_X1 U5749 ( .A1(n5037), .A2(n4340), .ZN(n8902) );
  NAND2_X1 U5750 ( .A1(n5708), .A2(n5882), .ZN(n8935) );
  AOI21_X1 U5751 ( .B1(n5041), .B2(n5044), .A(n4374), .ZN(n5040) );
  AND2_X1 U5752 ( .A1(n5047), .A2(n5043), .ZN(n5041) );
  OR2_X1 U5753 ( .A1(n4401), .A2(n4342), .ZN(n4467) );
  OR2_X1 U5754 ( .A1(n5986), .A2(n6973), .ZN(n5982) );
  OR2_X1 U5755 ( .A1(n5645), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n5661) );
  INV_X1 U5756 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n10273) );
  INV_X1 U5757 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5381) );
  NAND2_X1 U5758 ( .A1(n5253), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4448) );
  AND2_X1 U5759 ( .A1(n6555), .A2(n6554), .ZN(n6641) );
  NAND2_X1 U5760 ( .A1(n6113), .A2(n4613), .ZN(n4612) );
  AND2_X1 U5761 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6141) );
  NAND2_X1 U5762 ( .A1(n7700), .A2(n7699), .ZN(n7698) );
  NAND2_X1 U5763 ( .A1(n7700), .A2(n4779), .ZN(n4778) );
  AND2_X1 U5764 ( .A1(n4809), .A2(n4811), .ZN(n9131) );
  AND2_X1 U5765 ( .A1(n6141), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6161) );
  AND2_X1 U5766 ( .A1(n9180), .A2(n9181), .ZN(n9259) );
  OR2_X1 U5767 ( .A1(n6628), .A2(n8444), .ZN(n6614) );
  OR2_X1 U5768 ( .A1(n6320), .A2(n6319), .ZN(n6340) );
  NAND2_X1 U5769 ( .A1(n6338), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6355) );
  INV_X1 U5770 ( .A(n6340), .ZN(n6338) );
  AND2_X1 U5771 ( .A1(n6545), .A2(n6544), .ZN(n9173) );
  OR2_X1 U5772 ( .A1(n9414), .A2(n6561), .ZN(n6545) );
  AND2_X1 U5773 ( .A1(n6513), .A2(n6512), .ZN(n9172) );
  INV_X1 U5774 ( .A(n4335), .ZN(n6620) );
  AND4_X1 U5775 ( .A1(n6238), .A2(n6237), .A3(n6236), .A4(n6235), .ZN(n7863)
         );
  NAND2_X1 U5776 ( .A1(n6871), .A2(n4362), .ZN(n9315) );
  AND2_X1 U5777 ( .A1(n6940), .A2(n4525), .ZN(n6769) );
  NAND2_X1 U5778 ( .A1(n6767), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4525) );
  NOR2_X1 U5779 ( .A1(n6769), .A2(n6768), .ZN(n6792) );
  OR2_X1 U5780 ( .A1(n7716), .A2(n4521), .ZN(n4520) );
  AND2_X1 U5781 ( .A1(n7717), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4521) );
  NOR2_X1 U5782 ( .A1(n7962), .A2(n4518), .ZN(n8104) );
  AND2_X1 U5783 ( .A1(n7963), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4518) );
  NAND2_X1 U5784 ( .A1(n9428), .A2(n4771), .ZN(n9360) );
  NOR2_X1 U5785 ( .A1(n9372), .A2(n4772), .ZN(n4771) );
  INV_X1 U5786 ( .A(n4773), .ZN(n4772) );
  NOR2_X1 U5787 ( .A1(n9382), .A2(n8278), .ZN(n4786) );
  NAND2_X1 U5788 ( .A1(n4792), .A2(n8346), .ZN(n4791) );
  NAND2_X1 U5789 ( .A1(n4789), .A2(n9608), .ZN(n4788) );
  NAND2_X1 U5790 ( .A1(n4341), .A2(n8278), .ZN(n4789) );
  NAND2_X1 U5791 ( .A1(n8156), .A2(n8155), .ZN(n9376) );
  NAND2_X1 U5792 ( .A1(n9394), .A2(n9393), .ZN(n9392) );
  OR2_X1 U5793 ( .A1(n9394), .A2(n9393), .ZN(n4580) );
  OR2_X1 U5794 ( .A1(n9397), .A2(n9490), .ZN(n4604) );
  AND2_X1 U5795 ( .A1(n6538), .A2(n6527), .ZN(n9430) );
  AND2_X1 U5796 ( .A1(n8343), .A2(n8351), .ZN(n9423) );
  OR2_X1 U5797 ( .A1(n6459), .A2(n6458), .ZN(n6478) );
  NOR2_X1 U5798 ( .A1(n9739), .A2(n9510), .ZN(n9494) );
  AND2_X1 U5799 ( .A1(n6485), .A2(n6484), .ZN(n9491) );
  NAND2_X1 U5800 ( .A1(n4766), .A2(n4765), .ZN(n9510) );
  NAND2_X1 U5801 ( .A1(n8173), .A2(n8423), .ZN(n9506) );
  AND2_X1 U5802 ( .A1(n8263), .A2(n8423), .ZN(n9520) );
  OAI21_X1 U5803 ( .B1(n4693), .B2(n4598), .A(n4418), .ZN(n9609) );
  NAND2_X1 U5804 ( .A1(n7914), .A2(n7867), .ZN(n4689) );
  NOR2_X1 U5805 ( .A1(n9770), .A2(n4769), .ZN(n4767) );
  NAND2_X1 U5806 ( .A1(n7915), .A2(n7914), .ZN(n9605) );
  INV_X1 U5807 ( .A(n6280), .ZN(n6278) );
  NAND2_X1 U5808 ( .A1(n4598), .A2(n8322), .ZN(n7915) );
  NAND2_X1 U5809 ( .A1(n7788), .A2(n4770), .ZN(n7921) );
  NAND2_X1 U5810 ( .A1(n7788), .A2(n9801), .ZN(n7862) );
  NAND2_X1 U5811 ( .A1(n7778), .A2(n8320), .ZN(n7856) );
  NAND2_X1 U5812 ( .A1(n7785), .A2(n7784), .ZN(n7866) );
  OAI21_X1 U5813 ( .B1(n7536), .B2(n4505), .A(n4502), .ZN(n7675) );
  INV_X1 U5814 ( .A(n4961), .ZN(n4505) );
  AOI21_X1 U5815 ( .B1(n4961), .B2(n4504), .A(n4503), .ZN(n4502) );
  NOR2_X1 U5816 ( .A1(n4965), .A2(n4962), .ZN(n4961) );
  NAND2_X1 U5817 ( .A1(n7536), .A2(n7519), .ZN(n7520) );
  AND2_X1 U5818 ( .A1(n7119), .A2(n8372), .ZN(n9613) );
  INV_X1 U5819 ( .A(n9289), .ZN(n7545) );
  INV_X1 U5820 ( .A(n9608), .ZN(n9592) );
  NAND2_X1 U5821 ( .A1(n7230), .A2(n7218), .ZN(n7270) );
  INV_X1 U5822 ( .A(n9524), .ZN(n9490) );
  INV_X1 U5823 ( .A(n9523), .ZN(n9488) );
  NAND2_X1 U5824 ( .A1(n7636), .A2(n7164), .ZN(n7145) );
  INV_X1 U5825 ( .A(n9613), .ZN(n9595) );
  OR2_X1 U5826 ( .A1(n7157), .A2(n7156), .ZN(n7165) );
  NAND2_X1 U5827 ( .A1(n8295), .A2(n8294), .ZN(n9352) );
  NAND2_X1 U5828 ( .A1(n8290), .A2(n8289), .ZN(n9361) );
  AND2_X1 U5829 ( .A1(n8358), .A2(n8283), .ZN(n9382) );
  INV_X1 U5830 ( .A(n9376), .ZN(n4606) );
  NAND2_X1 U5831 ( .A1(n6525), .A2(n6524), .ZN(n8186) );
  NOR2_X1 U5832 ( .A1(n9739), .A2(n9277), .ZN(n4953) );
  AND2_X1 U5833 ( .A1(n8304), .A2(n8303), .ZN(n9486) );
  NAND2_X1 U5834 ( .A1(n9750), .A2(n8200), .ZN(n4508) );
  NAND2_X1 U5835 ( .A1(n4970), .A2(n4969), .ZN(n4509) );
  NAND2_X1 U5836 ( .A1(n9528), .A2(n9278), .ZN(n4969) );
  NOR2_X1 U5837 ( .A1(n9766), .A2(n9281), .ZN(n8143) );
  NAND2_X1 U5838 ( .A1(n7866), .A2(n7865), .ZN(n7868) );
  OR2_X1 U5839 ( .A1(n7864), .A2(n9285), .ZN(n7865) );
  AND2_X1 U5840 ( .A1(n6160), .A2(n6159), .ZN(n9875) );
  NAND2_X1 U5841 ( .A1(n8193), .A2(n8338), .ZN(n7163) );
  NOR2_X1 U5842 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n4763) );
  NAND2_X1 U5843 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), 
        .ZN(n4782) );
  XNOR2_X1 U5844 ( .A(n6032), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6606) );
  XNOR2_X1 U5845 ( .A(n5616), .B(n5615), .ZN(n8028) );
  NAND2_X1 U5846 ( .A1(n5203), .A2(n5202), .ZN(n5616) );
  OR2_X1 U5847 ( .A1(n6040), .A2(n6039), .ZN(n4637) );
  NAND2_X1 U5848 ( .A1(n6040), .A2(n6039), .ZN(n6610) );
  INV_X1 U5849 ( .A(SI_20_), .ZN(n5562) );
  OAI21_X1 U5850 ( .B1(n5533), .B2(n5173), .A(n5172), .ZN(n5547) );
  AND2_X1 U5851 ( .A1(n6294), .A2(n6275), .ZN(n7466) );
  NAND2_X1 U5852 ( .A1(n4980), .A2(n5151), .ZN(n5419) );
  NAND2_X1 U5853 ( .A1(n4981), .A2(n4986), .ZN(n4980) );
  INV_X1 U5854 ( .A(n5395), .ZN(n4446) );
  AND2_X1 U5855 ( .A1(n5117), .A2(n5118), .ZN(n5288) );
  NAND2_X1 U5856 ( .A1(n4522), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6123) );
  INV_X1 U5857 ( .A(n6079), .ZN(n4522) );
  OR2_X1 U5858 ( .A1(n5101), .A2(SI_1_), .ZN(n4640) );
  NOR2_X1 U5859 ( .A1(n5106), .A2(n5105), .ZN(n5246) );
  OAI21_X1 U5860 ( .B1(n5111), .B2(P1_DATAO_REG_0__SCAN_IN), .A(n5104), .ZN(
        n5106) );
  NAND2_X1 U5861 ( .A1(n5111), .A2(n5103), .ZN(n5104) );
  INV_X4 U5862 ( .A(n6662), .ZN(n6661) );
  AND2_X1 U5863 ( .A1(n6700), .A2(n6657), .ZN(n6703) );
  INV_X1 U5864 ( .A(n7378), .ZN(n10053) );
  NAND2_X1 U5865 ( .A1(n8487), .A2(n8486), .ZN(n4900) );
  NAND2_X1 U5866 ( .A1(n8487), .A2(n4898), .ZN(n8502) );
  AND2_X1 U5867 ( .A1(n6977), .A2(n6976), .ZN(n8606) );
  NAND2_X1 U5868 ( .A1(n4610), .A2(n4609), .ZN(n8523) );
  NOR2_X1 U5869 ( .A1(n4539), .A2(n8833), .ZN(n4536) );
  NAND2_X1 U5870 ( .A1(n8492), .A2(n4540), .ZN(n4538) );
  NAND2_X1 U5871 ( .A1(n4561), .A2(n4564), .ZN(n8529) );
  OR2_X1 U5872 ( .A1(n4610), .A2(n4565), .ZN(n4561) );
  NAND2_X1 U5873 ( .A1(n5581), .A2(n5580), .ZN(n8534) );
  INV_X1 U5874 ( .A(n4569), .ZN(n7878) );
  AOI21_X1 U5875 ( .B1(n8579), .B2(n4556), .A(n4553), .ZN(n4552) );
  NAND2_X1 U5876 ( .A1(n4554), .A2(n4908), .ZN(n4553) );
  AOI21_X1 U5877 ( .B1(n4911), .B2(n4913), .A(n4387), .ZN(n4908) );
  NAND2_X1 U5878 ( .A1(n4918), .A2(n4919), .ZN(n8545) );
  INV_X1 U5879 ( .A(n4913), .ZN(n4909) );
  NAND2_X1 U5880 ( .A1(n8513), .A2(n4912), .ZN(n4910) );
  NAND2_X1 U5881 ( .A1(n8523), .A2(n8471), .ZN(n8570) );
  NAND2_X1 U5882 ( .A1(n4568), .A2(n4567), .ZN(n7971) );
  NAND2_X1 U5883 ( .A1(n4569), .A2(n8625), .ZN(n4567) );
  AND3_X1 U5884 ( .A1(n5561), .A2(n5560), .A3(n5559), .ZN(n8925) );
  NAND2_X1 U5885 ( .A1(n4532), .A2(n4533), .ZN(n7174) );
  NAND2_X1 U5886 ( .A1(n4534), .A2(n4359), .ZN(n4533) );
  NAND2_X1 U5887 ( .A1(n4393), .A2(n7107), .ZN(n4532) );
  INV_X1 U5888 ( .A(n7171), .ZN(n4534) );
  NAND2_X1 U5889 ( .A1(n7173), .A2(n7174), .ZN(n7258) );
  NAND2_X1 U5890 ( .A1(n8463), .A2(n8462), .ZN(n8611) );
  AND2_X1 U5891 ( .A1(n6933), .A2(n6932), .ZN(n8608) );
  OAI211_X1 U5892 ( .C1(n5951), .C2(n6969), .A(n4638), .B(n4475), .ZN(n4474)
         );
  INV_X1 U5893 ( .A(n8824), .ZN(n8798) );
  INV_X1 U5894 ( .A(n8823), .ZN(n8847) );
  INV_X1 U5895 ( .A(n8925), .ZN(n8622) );
  NAND4_X1 U5896 ( .A1(n5337), .A2(n5336), .A3(n5335), .A4(n5334), .ZN(n8631)
         );
  INV_X1 U5897 ( .A(n7074), .ZN(n8635) );
  NAND2_X1 U5898 ( .A1(n5256), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5261) );
  INV_X1 U5899 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6736) );
  NAND2_X1 U5900 ( .A1(n6805), .A2(n4426), .ZN(n6705) );
  NAND2_X1 U5901 ( .A1(n4461), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6805) );
  INV_X1 U5902 ( .A(n4456), .ZN(n9929) );
  INV_X1 U5903 ( .A(n4488), .ZN(n9970) );
  INV_X1 U5904 ( .A(n4599), .ZN(n9976) );
  INV_X1 U5905 ( .A(n4459), .ZN(n9988) );
  AOI21_X1 U5906 ( .B1(n9954), .B2(n7340), .A(n9983), .ZN(n7342) );
  INV_X1 U5907 ( .A(n4873), .ZN(n10000) );
  XNOR2_X1 U5908 ( .A(n7420), .B(n7421), .ZN(n7316) );
  INV_X1 U5909 ( .A(n4597), .ZN(n7422) );
  INV_X1 U5910 ( .A(n4871), .ZN(n7425) );
  INV_X1 U5911 ( .A(n4888), .ZN(n7412) );
  INV_X1 U5912 ( .A(n4876), .ZN(n7934) );
  INV_X1 U5913 ( .A(n7824), .ZN(n7825) );
  INV_X1 U5914 ( .A(n4658), .ZN(n7948) );
  INV_X1 U5915 ( .A(n4874), .ZN(n8636) );
  INV_X1 U5916 ( .A(n4452), .ZN(n8680) );
  OR2_X1 U5917 ( .A1(n8682), .A2(n8049), .ZN(n4681) );
  INV_X1 U5918 ( .A(n4486), .ZN(n8710) );
  NAND2_X1 U5919 ( .A1(n4678), .A2(n4677), .ZN(n8720) );
  NAND2_X1 U5920 ( .A1(n5752), .A2(n5751), .ZN(n8784) );
  AND2_X1 U5921 ( .A1(n8781), .A2(n5650), .ZN(n8803) );
  AND2_X1 U5922 ( .A1(n5649), .A2(n5639), .ZN(n8813) );
  OAI21_X1 U5923 ( .B1(n5660), .B2(n10026), .A(n5659), .ZN(n8812) );
  NOR2_X1 U5924 ( .A1(n5658), .A2(n5657), .ZN(n5659) );
  NOR2_X1 U5925 ( .A1(n8505), .A2(n10030), .ZN(n5658) );
  NAND2_X1 U5926 ( .A1(n5231), .A2(n5230), .ZN(n8816) );
  AND2_X1 U5927 ( .A1(n5638), .A2(n5630), .ZN(n8826) );
  NAND2_X1 U5928 ( .A1(n5070), .A2(n5071), .ZN(n8866) );
  NAND2_X1 U5929 ( .A1(n8888), .A2(n5890), .ZN(n8881) );
  NAND2_X1 U5930 ( .A1(n8892), .A2(n5576), .ZN(n8876) );
  NAND2_X1 U5931 ( .A1(n5709), .A2(n5901), .ZN(n8918) );
  NAND2_X1 U5932 ( .A1(n5057), .A2(n5297), .ZN(n7186) );
  NAND2_X1 U5933 ( .A1(n5296), .A2(n5090), .ZN(n5057) );
  NAND2_X1 U5934 ( .A1(n8926), .A2(n10032), .ZN(n8959) );
  NAND2_X1 U5935 ( .A1(n6918), .A2(n6917), .ZN(n10021) );
  INV_X1 U5936 ( .A(n8912), .ZN(n8956) );
  OAI211_X2 U5937 ( .C1(n5314), .C2(n6668), .A(n5295), .B(n5294), .ZN(n7077)
         );
  INV_X1 U5938 ( .A(n9001), .ZN(n9006) );
  INV_X1 U5939 ( .A(n7101), .ZN(n7020) );
  NAND2_X1 U5940 ( .A1(n5744), .A2(n5743), .ZN(n9010) );
  AND2_X1 U5941 ( .A1(n5087), .A2(n8966), .ZN(n8967) );
  OAI21_X1 U5942 ( .B1(n5712), .B2(n4860), .A(n4858), .ZN(n5794) );
  NAND2_X1 U5943 ( .A1(n4862), .A2(n5924), .ZN(n8819) );
  NAND2_X1 U5944 ( .A1(n5712), .A2(n4863), .ZN(n4862) );
  NAND2_X1 U5945 ( .A1(n5712), .A2(n5917), .ZN(n8830) );
  NAND2_X1 U5946 ( .A1(n5235), .A2(n5234), .ZN(n9036) );
  INV_X1 U5947 ( .A(n5063), .ZN(n8858) );
  AOI21_X1 U5948 ( .B1(n5070), .B2(n5068), .A(n5064), .ZN(n5063) );
  NAND2_X1 U5949 ( .A1(n5591), .A2(n5590), .ZN(n9047) );
  OAI21_X1 U5950 ( .B1(n8888), .B2(n5895), .A(n4831), .ZN(n8872) );
  NAND2_X1 U5951 ( .A1(n5567), .A2(n5566), .ZN(n9058) );
  NAND2_X1 U5952 ( .A1(n8920), .A2(n5904), .ZN(n8910) );
  NAND2_X1 U5953 ( .A1(n5522), .A2(n5521), .ZN(n9073) );
  NAND2_X1 U5954 ( .A1(n5507), .A2(n5506), .ZN(n9080) );
  NAND2_X1 U5955 ( .A1(n5494), .A2(n5493), .ZN(n8616) );
  OAI21_X1 U5956 ( .B1(n5453), .B2(n5047), .A(n5044), .ZN(n8034) );
  AND2_X1 U5957 ( .A1(n7992), .A2(n7991), .ZN(n8023) );
  NAND2_X1 U5958 ( .A1(n5480), .A2(n5479), .ZN(n8024) );
  OAI21_X1 U5959 ( .B1(n10076), .B2(n4840), .A(n4342), .ZN(n7996) );
  NAND2_X1 U5960 ( .A1(n5453), .A2(n5452), .ZN(n8002) );
  NAND2_X1 U5961 ( .A1(n5460), .A2(n5459), .ZN(n8016) );
  NAND2_X1 U5962 ( .A1(n10076), .A2(n5862), .ZN(n8008) );
  INV_X1 U5963 ( .A(n9070), .ZN(n9079) );
  AND2_X1 U5964 ( .A1(n6681), .A2(n6923), .ZN(n6918) );
  CLKBUF_X1 U5965 ( .A(n9090), .Z(n4607) );
  XNOR2_X1 U5966 ( .A(n5665), .B(P2_IR_REG_26__SCAN_IN), .ZN(n8044) );
  XNOR2_X1 U5967 ( .A(n5097), .B(P2_IR_REG_22__SCAN_IN), .ZN(n7813) );
  NAND2_X1 U5968 ( .A1(n5661), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5097) );
  INV_X1 U5969 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10244) );
  INV_X1 U5970 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7284) );
  INV_X1 U5971 ( .A(n8702), .ZN(n8721) );
  NAND2_X1 U5972 ( .A1(n5491), .A2(n5478), .ZN(n8681) );
  INV_X1 U5973 ( .A(n8655), .ZN(n7950) );
  INV_X1 U5974 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6759) );
  INV_X1 U5975 ( .A(n7429), .ZN(n7745) );
  AND2_X1 U5976 ( .A1(n6661), .A2(P2_U3151), .ZN(n9100) );
  INV_X1 U5977 ( .A(n10002), .ZN(n7344) );
  OR2_X1 U5978 ( .A1(n5345), .A2(n5344), .ZN(n9959) );
  NAND2_X1 U5979 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5251) );
  NAND2_X1 U5980 ( .A1(n4800), .A2(n6172), .ZN(n7442) );
  OR2_X1 U5981 ( .A1(n4806), .A2(n4805), .ZN(n4800) );
  INV_X1 U5982 ( .A(n5078), .ZN(n4805) );
  NAND2_X1 U5983 ( .A1(n6156), .A2(n4807), .ZN(n4806) );
  INV_X1 U5984 ( .A(n4618), .ZN(n4617) );
  AND4_X1 U5985 ( .A1(n6183), .A2(n6182), .A3(n6181), .A4(n6180), .ZN(n7703)
         );
  INV_X1 U5986 ( .A(n9525), .ZN(n9489) );
  NAND2_X1 U5987 ( .A1(n4625), .A2(n6454), .ZN(n9154) );
  NAND2_X1 U5988 ( .A1(n6435), .A2(n4343), .ZN(n4625) );
  NAND2_X1 U5989 ( .A1(n4632), .A2(n4633), .ZN(n9171) );
  NAND2_X1 U5990 ( .A1(n9197), .A2(n9198), .ZN(n9196) );
  AOI21_X1 U5991 ( .B1(n8450), .B2(n8452), .A(n8451), .ZN(n8454) );
  INV_X1 U5992 ( .A(n4616), .ZN(n7291) );
  NAND2_X1 U5993 ( .A1(n9160), .A2(n6293), .ZN(n9216) );
  AND4_X1 U5994 ( .A1(n6256), .A2(n6255), .A3(n6254), .A4(n6253), .ZN(n9804)
         );
  NAND2_X1 U5995 ( .A1(n9144), .A2(n6073), .ZN(n7046) );
  INV_X1 U5996 ( .A(n9809), .ZN(n9245) );
  NAND2_X1 U5997 ( .A1(n8043), .A2(n8291), .ZN(n6536) );
  INV_X1 U5998 ( .A(n9265), .ZN(n9254) );
  AND2_X1 U5999 ( .A1(n6632), .A2(n8448), .ZN(n9814) );
  NAND2_X1 U6000 ( .A1(n4629), .A2(n4363), .ZN(n4628) );
  INV_X1 U6001 ( .A(n4630), .ZN(n4629) );
  AOI21_X1 U6002 ( .B1(n8378), .B2(n8383), .A(n8377), .ZN(n8441) );
  INV_X1 U6003 ( .A(n8376), .ZN(n8377) );
  OAI21_X1 U6004 ( .B1(n8379), .B2(n8338), .A(n8369), .ZN(n8378) );
  AOI21_X1 U6005 ( .B1(n8375), .B2(n6047), .A(n8374), .ZN(n8376) );
  INV_X1 U6006 ( .A(n8440), .ZN(n4735) );
  AND2_X1 U6007 ( .A1(n4737), .A2(n4734), .ZN(n4733) );
  NAND2_X1 U6008 ( .A1(n8440), .A2(n4378), .ZN(n4734) );
  INV_X1 U6009 ( .A(n9251), .ZN(n9272) );
  INV_X1 U6010 ( .A(n9173), .ZN(n9395) );
  INV_X1 U6011 ( .A(n9172), .ZN(n9274) );
  INV_X1 U6012 ( .A(n7703), .ZN(n7518) );
  INV_X1 U6013 ( .A(n7506), .ZN(n9290) );
  OR2_X1 U6014 ( .A1(n6423), .A2(n6116), .ZN(n6117) );
  NOR2_X1 U6015 ( .A1(n6832), .A2(n6831), .ZN(n6954) );
  AND2_X1 U6016 ( .A1(n4516), .A2(n4515), .ZN(n6832) );
  NAND2_X1 U6017 ( .A1(n6851), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4515) );
  NAND2_X1 U6018 ( .A1(n7083), .A2(n4408), .ZN(n7084) );
  INV_X1 U6019 ( .A(n4514), .ZN(n7194) );
  AND2_X1 U6020 ( .A1(n4514), .A2(n4513), .ZN(n7198) );
  NAND2_X1 U6021 ( .A1(n7200), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4513) );
  NOR2_X1 U6022 ( .A1(n7467), .A2(n7468), .ZN(n7716) );
  AND2_X1 U6023 ( .A1(n4520), .A2(n4519), .ZN(n7962) );
  INV_X1 U6024 ( .A(n7718), .ZN(n4519) );
  INV_X1 U6025 ( .A(n4520), .ZN(n7719) );
  INV_X1 U6026 ( .A(n4524), .ZN(n9328) );
  AND2_X1 U6027 ( .A1(n6695), .A2(n6762), .ZN(n9824) );
  NAND2_X1 U6028 ( .A1(n4929), .A2(n4493), .ZN(n9366) );
  NAND2_X1 U6029 ( .A1(n8156), .A2(n4375), .ZN(n4929) );
  AND2_X1 U6030 ( .A1(n9368), .A2(n6578), .ZN(n9386) );
  AND2_X1 U6031 ( .A1(n4947), .A2(n4952), .ZN(n9453) );
  OR2_X1 U6032 ( .A1(n8148), .A2(n4948), .ZN(n4947) );
  NAND2_X1 U6033 ( .A1(n9557), .A2(n8257), .ZN(n9536) );
  NAND2_X1 U6034 ( .A1(n8170), .A2(n8417), .ZN(n9555) );
  INV_X1 U6035 ( .A(n9766), .ZN(n9599) );
  NAND2_X1 U6036 ( .A1(n7568), .A2(n7572), .ZN(n7673) );
  NAND2_X1 U6037 ( .A1(n7567), .A2(n7566), .ZN(n7568) );
  NAND2_X1 U6038 ( .A1(n7509), .A2(n7541), .ZN(n7517) );
  NAND2_X1 U6039 ( .A1(n7508), .A2(n7507), .ZN(n7509) );
  NAND2_X1 U6040 ( .A1(n7217), .A2(n7216), .ZN(n7231) );
  OR2_X1 U6041 ( .A1(n9617), .A2(n8383), .ZN(n9621) );
  NOR2_X1 U6042 ( .A1(n9617), .A2(n7482), .ZN(n9868) );
  INV_X1 U6043 ( .A(n9621), .ZN(n9858) );
  OR2_X1 U6044 ( .A1(n6615), .A2(n8444), .ZN(n9544) );
  NAND2_X1 U6045 ( .A1(n6248), .A2(n6247), .ZN(n9128) );
  AND2_X1 U6046 ( .A1(n9896), .A2(n7135), .ZN(n9695) );
  INV_X1 U6047 ( .A(n9352), .ZN(n9703) );
  INV_X1 U6048 ( .A(n9361), .ZN(n9707) );
  INV_X1 U6049 ( .A(n8186), .ZN(n9722) );
  NAND2_X1 U6050 ( .A1(n6505), .A2(n6504), .ZN(n9725) );
  OR2_X1 U6051 ( .A1(n8148), .A2(n4945), .ZN(n4939) );
  INV_X1 U6052 ( .A(n9462), .ZN(n9731) );
  NAND2_X1 U6053 ( .A1(n6475), .A2(n6474), .ZN(n9734) );
  NAND2_X1 U6054 ( .A1(n6414), .A2(n6413), .ZN(n9751) );
  INV_X1 U6055 ( .A(n9561), .ZN(n9760) );
  NAND2_X1 U6056 ( .A1(n8140), .A2(n8139), .ZN(n9603) );
  INV_X1 U6057 ( .A(n7214), .ZN(n7629) );
  AND3_X1 U6058 ( .A1(n6130), .A2(n6129), .A3(n6128), .ZN(n7290) );
  AND2_X1 U6059 ( .A1(n7986), .A2(n8055), .ZN(n6715) );
  INV_X1 U6060 ( .A(n9871), .ZN(n9872) );
  OR2_X1 U6061 ( .A1(n9777), .A2(n4938), .ZN(n4937) );
  INV_X1 U6062 ( .A(n4934), .ZN(n4784) );
  NAND2_X1 U6063 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_30__SCAN_IN), 
        .ZN(n4938) );
  INV_X1 U6064 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U6065 ( .A1(n6051), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4776) );
  XNOR2_X1 U6066 ( .A(n6034), .B(n6033), .ZN(n8032) );
  NOR2_X1 U6067 ( .A1(n6005), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n4971) );
  INV_X1 U6068 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7908) );
  NAND2_X1 U6069 ( .A1(n4657), .A2(n5600), .ZN(n7906) );
  INV_X1 U6070 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7855) );
  INV_X1 U6071 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7707) );
  INV_X1 U6072 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8058) );
  INV_X1 U6073 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7438) );
  INV_X1 U6074 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10271) );
  NAND2_X1 U6075 ( .A1(n6001), .A2(n6000), .ZN(n6349) );
  NAND2_X1 U6076 ( .A1(n4976), .A2(n4977), .ZN(n5436) );
  OAI21_X1 U6077 ( .B1(n5356), .B2(n5084), .A(n5357), .ZN(n6683) );
  OAI21_X1 U6078 ( .B1(n4351), .B2(n5338), .A(n5339), .ZN(n6676) );
  XNOR2_X1 U6079 ( .A(n6064), .B(n6063), .ZN(n9299) );
  NAND2_X1 U6080 ( .A1(n7107), .A2(n7106), .ZN(n7172) );
  NAND2_X1 U6081 ( .A1(n7026), .A2(n7025), .ZN(n7029) );
  AND2_X1 U6082 ( .A1(n4867), .A2(n4353), .ZN(n8732) );
  OAI21_X1 U6083 ( .B1(n8778), .B2(n10005), .A(n4465), .ZN(P2_U3201) );
  AOI21_X1 U6084 ( .B1(n8777), .B2(n9949), .A(n4466), .ZN(n4465) );
  NAND2_X1 U6085 ( .A1(n4581), .A2(n4682), .ZN(n4466) );
  OAI21_X1 U6086 ( .B1(n8789), .B2(n9001), .A(n5975), .ZN(n5976) );
  OAI21_X1 U6087 ( .B1(n8789), .B2(n9070), .A(n5990), .ZN(n5991) );
  NAND2_X1 U6088 ( .A1(n4818), .A2(n4365), .ZN(n6640) );
  INV_X1 U6089 ( .A(n4516), .ZN(n6847) );
  MUX2_X1 U6090 ( .A(n8133), .B(n8132), .S(n6047), .Z(n8136) );
  INV_X1 U6091 ( .A(n4577), .ZN(n4576) );
  OAI22_X1 U6092 ( .A1(n9713), .A2(n9686), .B1(n9896), .B2(n9642), .ZN(n4577)
         );
  OAI21_X1 U6093 ( .B1(n8189), .B2(n4699), .A(n4697), .ZN(P1_U3519) );
  NOR2_X1 U6094 ( .A1(n4698), .A2(n4411), .ZN(n4697) );
  NOR2_X1 U6095 ( .A1(n9890), .A2(n8188), .ZN(n4698) );
  INV_X1 U6096 ( .A(n4821), .ZN(n4820) );
  OAI21_X1 U6097 ( .B1(n9710), .B2(n9774), .A(n4822), .ZN(n4821) );
  NOR2_X1 U6098 ( .A1(n4417), .A2(n4575), .ZN(n4574) );
  NOR2_X1 U6099 ( .A1(n9890), .A2(n9712), .ZN(n4575) );
  AND2_X2 U6100 ( .A1(n6037), .A2(n6653), .ZN(n6305) );
  OAI211_X1 U6101 ( .C1(n5314), .C2(n6667), .A(n5313), .B(n5312), .ZN(n7190)
         );
  NAND2_X1 U6102 ( .A1(n8160), .A2(n8159), .ZN(n4339) );
  AND2_X1 U6103 ( .A1(n5034), .A2(n5035), .ZN(n4340) );
  AND2_X1 U6104 ( .A1(n9382), .A2(n4791), .ZN(n4341) );
  AND2_X1 U6105 ( .A1(n5705), .A2(n4838), .ZN(n4342) );
  NAND2_X1 U6106 ( .A1(n4972), .A2(n5995), .ZN(n6174) );
  NOR2_X1 U6107 ( .A1(n5146), .A2(n5145), .ZN(n4986) );
  NOR2_X1 U6108 ( .A1(n4626), .A2(n6455), .ZN(n4343) );
  INV_X1 U6109 ( .A(n5132), .ZN(n4975) );
  NAND2_X1 U6110 ( .A1(n5031), .A2(n5030), .ZN(n5027) );
  INV_X1 U6111 ( .A(n4555), .ZN(n8513) );
  INV_X1 U6112 ( .A(n9744), .ZN(n4765) );
  AND2_X1 U6113 ( .A1(n8568), .A2(n8904), .ZN(n4344) );
  INV_X1 U6114 ( .A(n5655), .ZN(n6734) );
  AND2_X1 U6115 ( .A1(n5239), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4345) );
  NAND2_X1 U6116 ( .A1(n6318), .A2(n6317), .ZN(n9770) );
  AND2_X1 U6117 ( .A1(n5903), .A2(n5904), .ZN(n4346) );
  AND4_X1 U6118 ( .A1(n5252), .A2(n4877), .A3(n4706), .A4(n10246), .ZN(n4347)
         );
  INV_X1 U6119 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6033) );
  INV_X1 U6120 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5227) );
  AND2_X1 U6121 ( .A1(n7401), .A2(n7495), .ZN(n4348) );
  AND2_X1 U6122 ( .A1(n4467), .A2(n5876), .ZN(n4349) );
  AND2_X1 U6123 ( .A1(n4985), .A2(n4984), .ZN(n4350) );
  XNOR2_X1 U6124 ( .A(n5786), .B(n5785), .ZN(n9096) );
  NAND2_X1 U6125 ( .A1(n7258), .A2(n4914), .ZN(n7402) );
  INV_X1 U6126 ( .A(n6074), .ZN(n6423) );
  AND2_X1 U6127 ( .A1(n4571), .A2(n5132), .ZN(n4351) );
  NAND2_X1 U6128 ( .A1(n8892), .A2(n5073), .ZN(n5070) );
  AND2_X2 U6129 ( .A1(n4705), .A2(n4706), .ZN(n5366) );
  INV_X1 U6130 ( .A(n8633), .ZN(n7110) );
  OR2_X1 U6131 ( .A1(n8744), .A2(n8729), .ZN(n4353) );
  AND2_X1 U6132 ( .A1(n5159), .A2(n5158), .ZN(n4354) );
  OAI21_X1 U6133 ( .B1(n6683), .B2(n5314), .A(n5361), .ZN(n7378) );
  NAND2_X1 U6134 ( .A1(n5366), .A2(n4836), .ZN(n5664) );
  AND2_X1 U6135 ( .A1(n4632), .A2(n4630), .ZN(n4355) );
  AND2_X1 U6136 ( .A1(n4627), .A2(n4628), .ZN(n4356) );
  AND2_X1 U6137 ( .A1(n9428), .A2(n4773), .ZN(n4357) );
  OR2_X1 U6138 ( .A1(n9153), .A2(n4624), .ZN(n4358) );
  NAND2_X1 U6139 ( .A1(n7359), .A2(n7170), .ZN(n4359) );
  XNOR2_X1 U6140 ( .A(n8505), .B(n8965), .ZN(n8808) );
  INV_X1 U6141 ( .A(n8808), .ZN(n4591) );
  OR2_X1 U6142 ( .A1(n7421), .A2(n7420), .ZN(n4360) );
  NAND2_X1 U6143 ( .A1(n5626), .A2(n5625), .ZN(n9024) );
  AND2_X1 U6144 ( .A1(n6023), .A2(n6020), .ZN(n6027) );
  AND2_X1 U6145 ( .A1(n6060), .A2(n6059), .ZN(n4361) );
  OR2_X1 U6146 ( .A1(n6876), .A2(n6765), .ZN(n4362) );
  NAND2_X1 U6147 ( .A1(n4939), .A2(n4944), .ZN(n9436) );
  NOR2_X1 U6148 ( .A1(n9247), .A2(n9248), .ZN(n4363) );
  AND2_X1 U6149 ( .A1(n4796), .A2(n6310), .ZN(n4364) );
  NAND2_X1 U6150 ( .A1(n4910), .A2(n4909), .ZN(n8560) );
  INV_X1 U6151 ( .A(n5047), .ZN(n5046) );
  OR2_X1 U6152 ( .A1(n5487), .A2(n5048), .ZN(n5047) );
  AND3_X1 U6153 ( .A1(n6635), .A2(n9809), .A3(n6634), .ZN(n4365) );
  OR2_X1 U6154 ( .A1(n9983), .A2(n7313), .ZN(n4366) );
  XNOR2_X1 U6155 ( .A(n5327), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9939) );
  AND2_X1 U6156 ( .A1(n7541), .A2(n8306), .ZN(n4367) );
  OR2_X1 U6157 ( .A1(n9010), .A2(n5768), .ZN(n4368) );
  INV_X1 U6158 ( .A(n5769), .ZN(n5048) );
  INV_X1 U6159 ( .A(n8521), .ZN(n4609) );
  NAND2_X1 U6160 ( .A1(n6232), .A2(n6231), .ZN(n7864) );
  AND2_X1 U6161 ( .A1(n4977), .A2(n4983), .ZN(n4369) );
  AND3_X1 U6162 ( .A1(n4439), .A2(n4739), .A3(n4438), .ZN(n4370) );
  NOR2_X1 U6163 ( .A1(n8700), .A2(n8701), .ZN(n4371) );
  OR2_X1 U6164 ( .A1(n9036), .A2(n8516), .ZN(n5917) );
  AND2_X1 U6165 ( .A1(n5366), .A2(n4834), .ZN(n4372) );
  NOR2_X1 U6166 ( .A1(n4742), .A2(n4334), .ZN(n4373) );
  INV_X1 U6167 ( .A(n9225), .ZN(n8137) );
  AND2_X1 U6168 ( .A1(n6297), .A2(n6296), .ZN(n9225) );
  OR2_X1 U6169 ( .A1(n9399), .A2(n9251), .ZN(n8346) );
  AND2_X1 U6170 ( .A1(n8616), .A2(n8948), .ZN(n4374) );
  AND2_X1 U6171 ( .A1(n4933), .A2(n4931), .ZN(n4375) );
  NAND2_X1 U6172 ( .A1(n5932), .A2(n5933), .ZN(n5964) );
  NOR2_X1 U6173 ( .A1(n4979), .A2(n5418), .ZN(n4978) );
  NAND2_X1 U6174 ( .A1(n5600), .A2(n5196), .ZN(n5232) );
  AND2_X1 U6175 ( .A1(n6661), .A2(n5100), .ZN(n4376) );
  AND2_X1 U6176 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n4377) );
  NAND2_X1 U6177 ( .A1(n6575), .A2(n6574), .ZN(n9709) );
  AND2_X1 U6178 ( .A1(n8299), .A2(n4334), .ZN(n4378) );
  AND4_X1 U6179 ( .A1(n6218), .A2(n6217), .A3(n6216), .A4(n6215), .ZN(n7672)
         );
  AND4_X1 U6180 ( .A1(n6198), .A2(n6197), .A3(n6196), .A4(n6195), .ZN(n7760)
         );
  OR2_X1 U6181 ( .A1(n7131), .A2(n6112), .ZN(n4379) );
  INV_X1 U6182 ( .A(n8331), .ZN(n9438) );
  AND2_X1 U6183 ( .A1(n8340), .A2(n8347), .ZN(n8331) );
  OR2_X1 U6184 ( .A1(n9073), .A2(n8924), .ZN(n5885) );
  NOR2_X1 U6185 ( .A1(n8024), .A2(n8623), .ZN(n4380) );
  NOR2_X1 U6186 ( .A1(n4904), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n4381) );
  AND2_X1 U6187 ( .A1(n9875), .A2(n7545), .ZN(n4382) );
  INV_X1 U6188 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6010) );
  NOR2_X1 U6189 ( .A1(n9024), .A2(n8482), .ZN(n4383) );
  AND2_X1 U6190 ( .A1(n8520), .A2(n8622), .ZN(n4384) );
  NOR2_X1 U6191 ( .A1(n9287), .A2(n7763), .ZN(n4385) );
  AND2_X1 U6192 ( .A1(n8346), .A2(n8281), .ZN(n9393) );
  INV_X1 U6193 ( .A(n9393), .ZN(n4792) );
  OR2_X1 U6194 ( .A1(n9590), .A2(n8169), .ZN(n4386) );
  INV_X1 U6195 ( .A(n5074), .ZN(n5073) );
  NAND2_X1 U6196 ( .A1(n5076), .A2(n5576), .ZN(n5074) );
  INV_X1 U6197 ( .A(n4769), .ZN(n4768) );
  NAND2_X1 U6198 ( .A1(n4770), .A2(n9225), .ZN(n4769) );
  INV_X1 U6199 ( .A(n5297), .ZN(n5060) );
  AND2_X1 U6200 ( .A1(n8479), .A2(n8516), .ZN(n4387) );
  AND2_X1 U6201 ( .A1(n5139), .A2(n5138), .ZN(n4388) );
  OR2_X1 U6202 ( .A1(n9042), .A2(n8848), .ZN(n4389) );
  OR2_X1 U6203 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_30__SCAN_IN), .ZN(
        n4390) );
  OR2_X1 U6204 ( .A1(n8821), .A2(n5927), .ZN(n4391) );
  INV_X1 U6205 ( .A(n8334), .ZN(n4933) );
  AND2_X1 U6206 ( .A1(n8359), .A2(n8364), .ZN(n8334) );
  AND2_X1 U6207 ( .A1(n5798), .A2(n4845), .ZN(n4392) );
  INV_X1 U6208 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9086) );
  AND2_X1 U6209 ( .A1(n4359), .A2(n7106), .ZN(n4393) );
  INV_X1 U6210 ( .A(n4986), .ZN(n4982) );
  INV_X1 U6211 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6000) );
  OR2_X1 U6212 ( .A1(n8520), .A2(n8925), .ZN(n5903) );
  INV_X1 U6213 ( .A(n5027), .ZN(n5026) );
  NAND2_X1 U6214 ( .A1(n4952), .A2(n8150), .ZN(n4394) );
  NOR2_X1 U6215 ( .A1(n8148), .A2(n4953), .ZN(n4395) );
  OR2_X1 U6216 ( .A1(n8255), .A2(n8254), .ZN(n4396) );
  OR2_X1 U6217 ( .A1(n5944), .A2(n5945), .ZN(n4397) );
  AND2_X1 U6218 ( .A1(n6429), .A2(n4811), .ZN(n4398) );
  AND2_X1 U6219 ( .A1(n5946), .A2(n5932), .ZN(n4399) );
  OR2_X1 U6220 ( .A1(n4338), .A2(n10022), .ZN(n4400) );
  NAND2_X1 U6221 ( .A1(n5871), .A2(n4837), .ZN(n4401) );
  AND2_X1 U6222 ( .A1(n9456), .A2(n9454), .ZN(n4402) );
  AND2_X1 U6223 ( .A1(n4815), .A2(n8257), .ZN(n4403) );
  AND2_X1 U6224 ( .A1(n4363), .A2(n4634), .ZN(n4404) );
  NOR2_X1 U6225 ( .A1(n8568), .A2(n8904), .ZN(n4405) );
  AND2_X1 U6226 ( .A1(n5252), .A2(n10279), .ZN(n5292) );
  NAND2_X1 U6227 ( .A1(n6001), .A2(n4971), .ZN(n4406) );
  NAND2_X1 U6228 ( .A1(n8597), .A2(n4536), .ZN(n4407) );
  XNOR2_X1 U6229 ( .A(n6030), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6592) );
  AND2_X1 U6230 ( .A1(n4547), .A2(n4545), .ZN(n8552) );
  XNOR2_X1 U6231 ( .A(n5758), .B(SI_29_), .ZN(n9093) );
  INV_X1 U6232 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n4573) );
  NOR2_X1 U6233 ( .A1(n9547), .A2(n9528), .ZN(n4766) );
  INV_X1 U6234 ( .A(n4495), .ZN(n6001) );
  NAND2_X1 U6235 ( .A1(n4972), .A2(n4496), .ZN(n4495) );
  INV_X1 U6236 ( .A(n8882), .ZN(n5072) );
  OAI22_X1 U6237 ( .A1(n9584), .A2(n8143), .B1(n8168), .B2(n9599), .ZN(n9568)
         );
  OR2_X1 U6238 ( .A1(n7087), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4408) );
  INV_X1 U6239 ( .A(n8627), .ZN(n7819) );
  NAND2_X1 U6240 ( .A1(n9161), .A2(n9162), .ZN(n9160) );
  NAND2_X1 U6241 ( .A1(n9216), .A2(n9217), .ZN(n9215) );
  INV_X1 U6242 ( .A(n8578), .ZN(n4559) );
  AND2_X1 U6243 ( .A1(n4617), .A2(n6334), .ZN(n4409) );
  AND2_X1 U6244 ( .A1(n7345), .A2(n7421), .ZN(n4410) );
  AND2_X1 U6245 ( .A1(n9372), .A2(n9769), .ZN(n4411) );
  AND4_X1 U6246 ( .A1(n5514), .A2(n5513), .A3(n5512), .A4(n5511), .ZN(n8604)
         );
  INV_X1 U6247 ( .A(n8833), .ZN(n8482) );
  AND2_X1 U6248 ( .A1(n7969), .A2(n8624), .ZN(n4412) );
  NAND2_X1 U6249 ( .A1(n10079), .A2(n8625), .ZN(n4413) );
  AND2_X1 U6250 ( .A1(n8463), .A2(n4922), .ZN(n4414) );
  INV_X1 U6251 ( .A(n9399), .ZN(n9713) );
  NAND2_X1 U6252 ( .A1(n6557), .A2(n6556), .ZN(n9399) );
  NOR2_X1 U6253 ( .A1(n5162), .A2(SI_16_), .ZN(n4415) );
  OR2_X1 U6254 ( .A1(n4765), .A2(n9489), .ZN(n4416) );
  INV_X1 U6255 ( .A(n9169), .ZN(n7909) );
  AND2_X1 U6256 ( .A1(n6277), .A2(n6276), .ZN(n9169) );
  NOR2_X1 U6257 ( .A1(n9713), .A2(n9759), .ZN(n4417) );
  AND2_X1 U6258 ( .A1(n8250), .A2(n4689), .ZN(n4418) );
  AND2_X1 U6259 ( .A1(n4681), .A2(n4680), .ZN(n4419) );
  INV_X1 U6260 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6039) );
  AND2_X1 U6261 ( .A1(n5682), .A2(n8044), .ZN(n5688) );
  NAND2_X1 U6262 ( .A1(n5538), .A2(n5537), .ZN(n8931) );
  INV_X1 U6263 ( .A(n8931), .ZN(n5036) );
  NAND2_X1 U6264 ( .A1(n7368), .A2(n7367), .ZN(n7366) );
  NOR2_X1 U6265 ( .A1(n5838), .A2(n4851), .ZN(n4850) );
  AND2_X1 U6266 ( .A1(n7788), .A2(n4768), .ZN(n4420) );
  NAND2_X1 U6267 ( .A1(n7269), .A2(n7219), .ZN(n7220) );
  XNOR2_X1 U6268 ( .A(n7255), .B(n8631), .ZN(n7173) );
  INV_X1 U6269 ( .A(n7569), .ZN(n4962) );
  NAND2_X1 U6270 ( .A1(n4616), .A2(n4615), .ZN(n7292) );
  AND2_X1 U6271 ( .A1(n4852), .A2(n5843), .ZN(n4421) );
  AND2_X1 U6272 ( .A1(n8681), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4422) );
  NAND2_X1 U6273 ( .A1(n7949), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4423) );
  INV_X1 U6274 ( .A(SI_15_), .ZN(n5011) );
  AND2_X1 U6275 ( .A1(n7258), .A2(n7257), .ZN(n4424) );
  AND4_X2 U6276 ( .A1(n7058), .A2(n5979), .A3(n6916), .A4(n7057), .ZN(n10096)
         );
  AND2_X2 U6277 ( .A1(n6905), .A2(n6904), .ZN(n9890) );
  INV_X1 U6278 ( .A(n9890), .ZN(n4699) );
  AND2_X2 U6279 ( .A1(n6904), .A2(n7156), .ZN(n9896) );
  NAND2_X1 U6280 ( .A1(n7149), .A2(n8308), .ZN(n7217) );
  NOR2_X1 U6281 ( .A1(n8691), .A2(n8049), .ZN(n4425) );
  OR2_X1 U6282 ( .A1(n4461), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n4426) );
  NAND2_X1 U6283 ( .A1(n7026), .A2(n4901), .ZN(n7107) );
  AND2_X2 U6284 ( .A1(n7695), .A2(n7813), .ZN(n6656) );
  INV_X1 U6285 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6028) );
  OR2_X1 U6286 ( .A1(n9978), .A2(n7342), .ZN(n4885) );
  NAND2_X1 U6287 ( .A1(n8721), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4427) );
  NAND2_X1 U6288 ( .A1(n8721), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4428) );
  XNOR2_X1 U6289 ( .A(n5098), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7695) );
  INV_X1 U6290 ( .A(n9995), .ZN(n4884) );
  INV_X1 U6291 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5008) );
  MUX2_X1 U6292 ( .A(n8339), .B(n8198), .S(n8381), .Z(n8273) );
  NAND2_X1 U6293 ( .A1(n8251), .A2(n8381), .ZN(n4750) );
  AND2_X1 U6294 ( .A1(n8210), .A2(n8381), .ZN(n4745) );
  NAND2_X1 U6295 ( .A1(n8204), .A2(n8381), .ZN(n4761) );
  XNOR2_X1 U6296 ( .A(n8729), .B(n8744), .ZN(n8711) );
  AOI21_X1 U6297 ( .B1(n8735), .B2(n8744), .A(n8734), .ZN(n8737) );
  XNOR2_X1 U6298 ( .A(n8743), .B(n8744), .ZN(n8722) );
  NAND2_X1 U6299 ( .A1(n5274), .A2(n5110), .ZN(n5289) );
  OAI21_X2 U6300 ( .B1(n5490), .B2(SI_15_), .A(n4429), .ZN(n5500) );
  NAND2_X1 U6301 ( .A1(n4435), .A2(n4642), .ZN(n4433) );
  NAND2_X1 U6302 ( .A1(n4373), .A2(n8276), .ZN(n4439) );
  OAI21_X1 U6303 ( .B1(n4738), .B2(n4373), .A(n4441), .ZN(n4440) );
  NAND2_X1 U6304 ( .A1(n8272), .A2(n8273), .ZN(n4443) );
  NAND2_X1 U6305 ( .A1(n5250), .A2(n5107), .ZN(n5271) );
  NAND2_X1 U6306 ( .A1(n4444), .A2(n5246), .ZN(n5250) );
  INV_X1 U6307 ( .A(n5248), .ZN(n4444) );
  NAND2_X1 U6308 ( .A1(n4640), .A2(n5107), .ZN(n5248) );
  NAND2_X1 U6309 ( .A1(n4445), .A2(n5395), .ZN(n5397) );
  XNOR2_X1 U6310 ( .A(n4981), .B(n4446), .ZN(n6709) );
  NOR2_X1 U6311 ( .A1(n7835), .A2(n7836), .ZN(n7839) );
  NAND3_X1 U6312 ( .A1(n4479), .A2(n4480), .A3(n4869), .ZN(n6730) );
  NOR2_X1 U6313 ( .A1(n7826), .A2(n7827), .ZN(n7830) );
  NOR2_X1 U6314 ( .A1(n8746), .A2(n8745), .ZN(n8749) );
  XNOR2_X1 U6315 ( .A(n4602), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n9899) );
  NAND2_X1 U6316 ( .A1(n4473), .A2(n5955), .ZN(P2_U3296) );
  NAND2_X1 U6317 ( .A1(n4474), .A2(n5952), .ZN(n4473) );
  NAND2_X1 U6318 ( .A1(n4476), .A2(n7097), .ZN(n4475) );
  INV_X1 U6319 ( .A(n4708), .ZN(n4476) );
  XNOR2_X2 U6320 ( .A(n4478), .B(n4477), .ZN(n5238) );
  NAND2_X1 U6321 ( .A1(n5814), .A2(n5815), .ZN(n5811) );
  NAND2_X1 U6322 ( .A1(n4482), .A2(n6741), .ZN(n4479) );
  NAND2_X1 U6323 ( .A1(n4481), .A2(n6741), .ZN(n6732) );
  NAND2_X1 U6324 ( .A1(n9902), .A2(n6728), .ZN(n4481) );
  INV_X1 U6325 ( .A(n9902), .ZN(n4482) );
  OAI21_X1 U6326 ( .B1(n6728), .B2(n9924), .A(P2_REG1_REG_3__SCAN_IN), .ZN(
        n4483) );
  NOR2_X1 U6327 ( .A1(n8666), .A2(n8667), .ZN(n8700) );
  OAI211_X1 U6328 ( .C1(n8701), .C2(n4485), .A(n4484), .B(n4487), .ZN(n4486)
         );
  OR2_X1 U6329 ( .A1(n8701), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4484) );
  INV_X1 U6330 ( .A(n8666), .ZN(n4485) );
  INV_X1 U6331 ( .A(n8703), .ZN(n4487) );
  OAI21_X1 U6332 ( .B1(n7149), .B2(n4492), .A(n4489), .ZN(n7230) );
  AOI21_X1 U6333 ( .B1(n9366), .B2(n9878), .A(n4701), .ZN(n4700) );
  INV_X1 U6334 ( .A(n4494), .ZN(n4493) );
  NAND2_X1 U6335 ( .A1(n9407), .A2(n8154), .ZN(n8156) );
  NAND3_X1 U6336 ( .A1(n4498), .A2(n4497), .A3(n4496), .ZN(n6031) );
  NAND4_X1 U6337 ( .A1(n6004), .A2(n6018), .A3(n6003), .A4(n6002), .ZN(n6005)
         );
  NAND3_X1 U6338 ( .A1(n5999), .A2(n5997), .A3(n5995), .ZN(n4499) );
  NAND2_X1 U6339 ( .A1(n5996), .A2(n5998), .ZN(n4501) );
  INV_X1 U6340 ( .A(n7122), .ZN(n7117) );
  NAND2_X1 U6341 ( .A1(n9316), .A2(n9315), .ZN(n9314) );
  NAND2_X1 U6342 ( .A1(n6872), .A2(n6873), .ZN(n6871) );
  XNOR2_X1 U6343 ( .A(n6876), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6873) );
  NAND2_X1 U6344 ( .A1(n5691), .A2(n6679), .ZN(n6972) );
  XNOR2_X1 U6345 ( .A(n8488), .B(n7101), .ZN(n6984) );
  OAI21_X1 U6346 ( .B1(n7174), .B2(n4535), .A(n4530), .ZN(n7590) );
  NAND4_X1 U6347 ( .A1(n4541), .A2(n4407), .A3(n4538), .A4(n4537), .ZN(n8497)
         );
  NAND3_X1 U6348 ( .A1(n8487), .A2(n8492), .A3(n4898), .ZN(n4541) );
  NAND2_X1 U6349 ( .A1(n4547), .A2(n4551), .ZN(n8553) );
  INV_X1 U6350 ( .A(n4552), .ZN(n8537) );
  NAND2_X1 U6351 ( .A1(n4560), .A2(n4562), .ZN(n8474) );
  NAND2_X1 U6352 ( .A1(n4610), .A2(n4564), .ZN(n4560) );
  AOI21_X1 U6353 ( .B1(n8537), .B2(n8538), .A(n8481), .ZN(n8485) );
  OAI21_X1 U6354 ( .B1(n7590), .B2(n7589), .A(n7588), .ZN(n7591) );
  NOR2_X1 U6355 ( .A1(n7808), .A2(n7807), .ZN(n7806) );
  NAND2_X1 U6356 ( .A1(n6982), .A2(n6983), .ZN(n6987) );
  XNOR2_X1 U6357 ( .A(n6984), .B(n10027), .ZN(n6982) );
  AND2_X4 U6358 ( .A1(n5263), .A2(n6662), .ZN(n5787) );
  NAND2_X1 U6359 ( .A1(n6007), .A2(n6006), .ZN(n6051) );
  NAND2_X1 U6360 ( .A1(n5131), .A2(n5130), .ZN(n4571) );
  NAND2_X1 U6361 ( .A1(n4579), .A2(n4603), .ZN(n9639) );
  NAND2_X1 U6362 ( .A1(n9571), .A2(n9570), .ZN(n8170) );
  AOI21_X1 U6363 ( .B1(n9472), .B2(n4402), .A(n4704), .ZN(n9437) );
  INV_X1 U6364 ( .A(n4703), .ZN(n9394) );
  OAI21_X1 U6365 ( .B1(n9711), .B2(n4699), .A(n4574), .ZN(P1_U3517) );
  NAND2_X1 U6366 ( .A1(n7669), .A2(n8319), .ZN(n7777) );
  NAND2_X1 U6367 ( .A1(n4578), .A2(n4576), .ZN(P1_U3549) );
  OR2_X1 U6368 ( .A1(n9711), .A2(n9893), .ZN(n4578) );
  OAI21_X1 U6369 ( .B1(n9409), .B2(n9408), .A(n8356), .ZN(n4703) );
  OR2_X2 U6370 ( .A1(n7697), .A2(n7760), .ZN(n8214) );
  INV_X1 U6371 ( .A(n8318), .ZN(n8397) );
  INV_X1 U6372 ( .A(n7857), .ZN(n4691) );
  NAND3_X1 U6373 ( .A1(n9392), .A2(n9608), .A3(n4580), .ZN(n4579) );
  NAND2_X1 U6374 ( .A1(n5271), .A2(n5109), .ZN(n5274) );
  XOR2_X1 U6375 ( .A(n6807), .B(n6718), .Z(n6806) );
  OAI21_X1 U6376 ( .B1(n7940), .B2(n7939), .A(n7938), .ZN(n7944) );
  NOR2_X1 U6377 ( .A1(n7329), .A2(n10010), .ZN(n7414) );
  NOR2_X1 U6378 ( .A1(n8647), .A2(n8646), .ZN(n8648) );
  NAND2_X1 U6379 ( .A1(n4648), .A2(n4397), .ZN(n4647) );
  AOI21_X1 U6380 ( .B1(n5875), .B2(n6656), .A(n5881), .ZN(n4731) );
  INV_X1 U6381 ( .A(n5831), .ZN(n4717) );
  NAND2_X1 U6382 ( .A1(n4713), .A2(n5986), .ZN(n4711) );
  NAND2_X1 U6383 ( .A1(n4650), .A2(n4399), .ZN(n4649) );
  AOI21_X1 U6384 ( .B1(n5868), .B2(n5867), .A(n5866), .ZN(n5869) );
  OAI21_X1 U6385 ( .B1(n5828), .B2(n5821), .A(n4715), .ZN(n5822) );
  AOI21_X1 U6386 ( .B1(n4730), .B2(n5884), .A(n4729), .ZN(n4728) );
  OAI22_X1 U6387 ( .A1(n5872), .A2(n7995), .B1(n6656), .B2(n5871), .ZN(n5879)
         );
  NAND2_X1 U6388 ( .A1(n5922), .A2(n5923), .ZN(n4589) );
  MUX2_X2 U6389 ( .A(n8190), .B(n8189), .S(n9896), .Z(n8192) );
  NAND2_X1 U6390 ( .A1(n4649), .A2(n5986), .ZN(n4648) );
  NAND2_X1 U6391 ( .A1(n5942), .A2(n8505), .ZN(n4650) );
  OAI21_X1 U6392 ( .B1(n4728), .B2(n6656), .A(n4726), .ZN(n5906) );
  AOI21_X1 U6393 ( .B1(n4732), .B2(n4731), .A(n5880), .ZN(n4730) );
  INV_X1 U6394 ( .A(n9518), .ZN(n4970) );
  NAND3_X1 U6395 ( .A1(n4592), .A2(n4591), .A3(n4590), .ZN(n5792) );
  NOR2_X2 U6396 ( .A1(n5554), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U6397 ( .A1(n4842), .A2(n4841), .ZN(n5800) );
  INV_X1 U6398 ( .A(n4605), .ZN(n9421) );
  AOI211_X1 U6399 ( .C1(n9641), .C2(n9878), .A(n9640), .B(n9639), .ZN(n9711)
         );
  AND2_X1 U6400 ( .A1(n7664), .A2(n8239), .ZN(n8318) );
  NAND2_X1 U6401 ( .A1(n5357), .A2(n5136), .ZN(n5365) );
  NAND2_X1 U6402 ( .A1(n8763), .A2(n6969), .ZN(n6973) );
  NAND2_X1 U6403 ( .A1(n6987), .A2(n6986), .ZN(n6997) );
  OR2_X2 U6404 ( .A1(n9470), .A2(n9474), .ZN(n9472) );
  NAND2_X1 U6405 ( .A1(n8174), .A2(n8270), .ZN(n9470) );
  NAND2_X1 U6406 ( .A1(n9437), .A2(n8331), .ZN(n9441) );
  OAI21_X1 U6407 ( .B1(n5111), .B2(n5100), .A(n5099), .ZN(n5101) );
  NAND2_X1 U6408 ( .A1(n5111), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5099) );
  NAND2_X1 U6409 ( .A1(n5339), .A2(n5132), .ZN(n5356) );
  NAND2_X1 U6410 ( .A1(n5667), .A2(n5666), .ZN(n4608) );
  XNOR2_X1 U6411 ( .A(n8488), .B(n6988), .ZN(n6998) );
  NAND4_X1 U6412 ( .A1(n5366), .A2(n4707), .A3(n5095), .A4(n5666), .ZN(n5228)
         );
  NAND2_X1 U6413 ( .A1(n7001), .A2(n7000), .ZN(n7002) );
  NAND2_X1 U6414 ( .A1(n7912), .A2(n4955), .ZN(n4954) );
  NAND2_X1 U6415 ( .A1(n4825), .A2(n4820), .ZN(P1_U3518) );
  OR2_X1 U6416 ( .A1(n8277), .A2(n8279), .ZN(n5082) );
  MUX2_X2 U6417 ( .A(n8297), .B(n4334), .S(n9361), .Z(n8300) );
  AOI21_X2 U6418 ( .B1(n8300), .B2(n5086), .A(n8299), .ZN(n8301) );
  OAI21_X1 U6419 ( .B1(n4783), .B2(n4782), .A(n6009), .ZN(n4781) );
  NAND2_X1 U6420 ( .A1(n4749), .A2(n8256), .ZN(n8264) );
  NAND2_X1 U6421 ( .A1(n4755), .A2(n4754), .ZN(n8272) );
  NAND2_X1 U6422 ( .A1(n4752), .A2(n4334), .ZN(n4751) );
  AOI21_X1 U6423 ( .B1(n8266), .B2(n4334), .A(n4757), .ZN(n4756) );
  INV_X1 U6424 ( .A(n8265), .ZN(n4759) );
  NOR3_X1 U6425 ( .A1(n8231), .A2(n9606), .A3(n8230), .ZN(n4753) );
  NAND2_X1 U6426 ( .A1(n4608), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U6427 ( .A1(n5309), .A2(n5123), .ZN(n5323) );
  NAND2_X1 U6428 ( .A1(n8585), .A2(n8469), .ZN(n8522) );
  INV_X1 U6429 ( .A(n8522), .ZN(n4610) );
  NAND2_X1 U6430 ( .A1(n8474), .A2(n8473), .ZN(n8579) );
  NAND3_X1 U6431 ( .A1(n4611), .A2(n6376), .A3(n4810), .ZN(n4809) );
  NAND3_X1 U6432 ( .A1(n4611), .A2(n6376), .A3(n9187), .ZN(n9197) );
  AND2_X1 U6433 ( .A1(n9183), .A2(n4611), .ZN(n9185) );
  NAND2_X1 U6434 ( .A1(n6366), .A2(n9188), .ZN(n4611) );
  NAND3_X1 U6435 ( .A1(n6113), .A2(n6073), .A3(n9144), .ZN(n4614) );
  NAND3_X1 U6436 ( .A1(n4379), .A2(n4614), .A3(n4612), .ZN(n4616) );
  NAND2_X1 U6437 ( .A1(n7046), .A2(n7047), .ZN(n7129) );
  NAND2_X1 U6438 ( .A1(n4793), .A2(n4364), .ZN(n6330) );
  XNOR2_X2 U6439 ( .A(n6203), .B(n6204), .ZN(n7700) );
  NAND3_X1 U6440 ( .A1(n5078), .A2(n4799), .A3(n6156), .ZN(n4621) );
  OAI21_X2 U6441 ( .B1(n6435), .B2(n4358), .A(n4622), .ZN(n6488) );
  NAND2_X1 U6442 ( .A1(n6435), .A2(n6434), .ZN(n9208) );
  INV_X1 U6443 ( .A(n6434), .ZN(n4626) );
  NOR2_X1 U6444 ( .A1(n6488), .A2(n6487), .ZN(n9226) );
  NAND2_X1 U6445 ( .A1(n8450), .A2(n4404), .ZN(n4627) );
  NAND2_X1 U6446 ( .A1(n8450), .A2(n4634), .ZN(n4632) );
  NAND3_X1 U6447 ( .A1(n4637), .A2(n6047), .A3(n6610), .ZN(n6896) );
  INV_X1 U6448 ( .A(n4636), .ZN(n6037) );
  NAND2_X1 U6449 ( .A1(n4708), .A2(n4639), .ZN(n4638) );
  NAND4_X1 U6450 ( .A1(n4655), .A2(n4654), .A3(n5896), .A4(n4652), .ZN(n5898)
         );
  NAND3_X1 U6451 ( .A1(n4994), .A2(n4998), .A3(n5599), .ZN(n4657) );
  NAND2_X1 U6452 ( .A1(n4662), .A2(n7100), .ZN(n6812) );
  NAND3_X1 U6453 ( .A1(n4676), .A2(n4674), .A3(n4672), .ZN(n7346) );
  INV_X1 U6454 ( .A(n4681), .ZN(n8688) );
  INV_X1 U6455 ( .A(n8689), .ZN(n4680) );
  NAND2_X1 U6456 ( .A1(n8250), .A2(n8322), .ZN(n4692) );
  INV_X1 U6457 ( .A(n7914), .ZN(n4693) );
  OAI21_X1 U6458 ( .B1(n4692), .B2(n4691), .A(n4690), .ZN(n9587) );
  NAND2_X1 U6459 ( .A1(n8214), .A2(n8224), .ZN(n8220) );
  NAND2_X1 U6460 ( .A1(n7665), .A2(n4694), .ZN(n8316) );
  NAND4_X1 U6461 ( .A1(n4707), .A2(n5666), .A3(n5095), .A4(n4347), .ZN(n5237)
         );
  AND2_X1 U6462 ( .A1(n4835), .A2(n5077), .ZN(n4707) );
  NAND2_X1 U6463 ( .A1(n4709), .A2(n4368), .ZN(n4708) );
  OAI211_X1 U6464 ( .C1(n4713), .C2(n4712), .A(n4711), .B(n4710), .ZN(n4709)
         );
  INV_X1 U6465 ( .A(n5811), .ZN(n4724) );
  NAND2_X1 U6466 ( .A1(n7142), .A2(n7141), .ZN(n7207) );
  NAND2_X1 U6467 ( .A1(n7122), .A2(n7121), .ZN(n7142) );
  NAND2_X1 U6468 ( .A1(n8345), .A2(n8343), .ZN(n4742) );
  AOI21_X2 U6469 ( .B1(n4743), .B2(n8223), .A(n8222), .ZN(n8235) );
  NAND3_X1 U6470 ( .A1(n4747), .A2(n4744), .A3(n8213), .ZN(n4743) );
  OR2_X1 U6471 ( .A1(n8212), .A2(n8211), .ZN(n4746) );
  NAND3_X1 U6472 ( .A1(n4751), .A2(n4750), .A3(n4396), .ZN(n4749) );
  OAI21_X1 U6473 ( .B1(n4753), .B2(n8385), .A(n8252), .ZN(n4752) );
  OAI22_X1 U6474 ( .A1(n4756), .A2(n8271), .B1(n4334), .B2(n8303), .ZN(n4755)
         );
  OAI21_X1 U6475 ( .B1(n4759), .B2(n4334), .A(n4758), .ZN(n4757) );
  NAND2_X1 U6476 ( .A1(n4760), .A2(n4761), .ZN(n8209) );
  NAND2_X1 U6477 ( .A1(n4764), .A2(n4763), .ZN(n6008) );
  NOR2_X2 U6478 ( .A1(n9576), .A2(n9561), .ZN(n9560) );
  NAND2_X1 U6479 ( .A1(n7788), .A2(n4767), .ZN(n9614) );
  AND2_X1 U6480 ( .A1(n9428), .A2(n4775), .ZN(n9385) );
  NAND2_X2 U6481 ( .A1(n6617), .A2(n9817), .ZN(n6062) );
  XNOR2_X2 U6482 ( .A(n4776), .B(n6052), .ZN(n9817) );
  OR2_X1 U6483 ( .A1(n7668), .A2(n8397), .ZN(n4777) );
  INV_X1 U6484 ( .A(n7756), .ZN(n4780) );
  NAND2_X1 U6485 ( .A1(n7698), .A2(n6206), .ZN(n7755) );
  AOI21_X1 U6486 ( .B1(n9394), .B2(n4341), .A(n4788), .ZN(n4787) );
  NAND2_X1 U6487 ( .A1(n4790), .A2(n4787), .ZN(n9384) );
  NAND2_X1 U6488 ( .A1(n9161), .A2(n4794), .ZN(n4793) );
  NAND2_X1 U6489 ( .A1(n5078), .A2(n6156), .ZN(n7381) );
  INV_X1 U6490 ( .A(n6173), .ZN(n4807) );
  NAND2_X1 U6491 ( .A1(n5089), .A2(n6334), .ZN(n9105) );
  NAND2_X1 U6492 ( .A1(n4809), .A2(n4398), .ZN(n6435) );
  OAI21_X1 U6493 ( .B1(n8203), .B2(n8306), .A(n8400), .ZN(n7542) );
  NAND2_X1 U6494 ( .A1(n8170), .A2(n4813), .ZN(n9557) );
  NAND2_X1 U6495 ( .A1(n9557), .A2(n4403), .ZN(n8172) );
  NAND2_X1 U6496 ( .A1(n9171), .A2(n4363), .ZN(n4817) );
  NAND2_X1 U6497 ( .A1(n8888), .A2(n4831), .ZN(n4828) );
  NAND2_X1 U6498 ( .A1(n4850), .A2(n4848), .ZN(n4847) );
  NAND2_X1 U6499 ( .A1(n5712), .A2(n4858), .ZN(n4855) );
  NAND2_X1 U6500 ( .A1(n4855), .A2(n4856), .ZN(n5795) );
  NAND2_X1 U6501 ( .A1(n10020), .A2(n4724), .ZN(n10019) );
  NAND2_X1 U6502 ( .A1(n5699), .A2(n5820), .ZN(n7391) );
  NAND2_X1 U6503 ( .A1(n5702), .A2(n5856), .ZN(n7898) );
  NAND2_X1 U6504 ( .A1(n10019), .A2(n5815), .ZN(n7070) );
  NAND4_X1 U6505 ( .A1(n5261), .A2(n5260), .A3(n5259), .A4(n5258), .ZN(n5697)
         );
  INV_X1 U6506 ( .A(n4867), .ZN(n8730) );
  NAND2_X1 U6507 ( .A1(n6732), .A2(n4869), .ZN(n9918) );
  INV_X1 U6508 ( .A(n6730), .ZN(n9916) );
  MUX2_X1 U6509 ( .A(n9104), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  MUX2_X1 U6510 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9104), .S(n5263), .Z(n7065) );
  INV_X1 U6511 ( .A(n4889), .ZN(n7409) );
  INV_X1 U6512 ( .A(n7411), .ZN(n4887) );
  NAND3_X1 U6513 ( .A1(n4892), .A2(n4890), .A3(n4891), .ZN(n4896) );
  NAND3_X1 U6514 ( .A1(n4892), .A2(n4894), .A3(n4891), .ZN(n9941) );
  INV_X1 U6515 ( .A(n4896), .ZN(n9940) );
  INV_X1 U6516 ( .A(n7339), .ZN(n4897) );
  AOI21_X1 U6517 ( .B1(n4900), .B2(n8501), .A(n8610), .ZN(n8503) );
  NAND2_X1 U6519 ( .A1(n5645), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5098) );
  INV_X1 U6520 ( .A(n8748), .ZN(n4917) );
  NAND2_X1 U6521 ( .A1(n7974), .A2(n4921), .ZN(n4918) );
  AND2_X1 U6522 ( .A1(n9725), .A2(n9274), .ZN(n4950) );
  NAND2_X1 U6523 ( .A1(n5203), .A2(n4990), .ZN(n4987) );
  NAND2_X1 U6524 ( .A1(n4987), .A2(n4988), .ZN(n5216) );
  NAND2_X1 U6525 ( .A1(n5579), .A2(n5000), .ZN(n4994) );
  NAND2_X1 U6526 ( .A1(n5456), .A2(n5159), .ZN(n5470) );
  NAND3_X1 U6527 ( .A1(n5238), .A2(n5239), .A3(P2_REG0_REG_1__SCAN_IN), .ZN(
        n5017) );
  NAND3_X1 U6528 ( .A1(n9094), .A2(n5238), .A3(P2_REG1_REG_1__SCAN_IN), .ZN(
        n5016) );
  INV_X1 U6529 ( .A(n5239), .ZN(n9094) );
  NAND2_X1 U6530 ( .A1(n4607), .A2(n5015), .ZN(n5019) );
  INV_X1 U6531 ( .A(n8820), .ZN(n5025) );
  OAI21_X1 U6532 ( .B1(n8820), .B2(n5635), .A(n5031), .ZN(n5957) );
  NAND2_X1 U6533 ( .A1(n5031), .A2(n5635), .ZN(n5029) );
  NAND2_X1 U6534 ( .A1(n8922), .A2(n4340), .ZN(n5032) );
  INV_X1 U6535 ( .A(n8890), .ZN(n5575) );
  NAND2_X1 U6536 ( .A1(n5453), .A2(n5042), .ZN(n5039) );
  NAND2_X1 U6537 ( .A1(n5039), .A2(n5040), .ZN(n8947) );
  OAI21_X1 U6538 ( .B1(n5296), .B2(n5055), .A(n5052), .ZN(n7392) );
  NAND2_X1 U6539 ( .A1(n8892), .A2(n5062), .ZN(n5061) );
  NAND2_X1 U6540 ( .A1(n5061), .A2(n5065), .ZN(n8846) );
  NAND2_X1 U6541 ( .A1(n9055), .A2(n8893), .ZN(n5076) );
  NAND4_X1 U6542 ( .A1(n5366), .A2(n5666), .A3(n5095), .A4(n5227), .ZN(n5669)
         );
  NOR2_X2 U6543 ( .A1(n9360), .A2(n9361), .ZN(n9359) );
  INV_X1 U6544 ( .A(n6368), .ZN(n6371) );
  NAND2_X1 U6545 ( .A1(n6089), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6013) );
  NOR2_X1 U6546 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5994) );
  INV_X1 U6547 ( .A(n10027), .ZN(n6913) );
  INV_X2 U6548 ( .A(n10082), .ZN(n10081) );
  AND2_X1 U6549 ( .A1(n7064), .A2(n10021), .ZN(n10034) );
  INV_X2 U6550 ( .A(n10034), .ZN(n8926) );
  INV_X1 U6551 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5100) );
  OR2_X1 U6552 ( .A1(n8285), .A2(n8284), .ZN(n5081) );
  AND3_X1 U6553 ( .A1(n8180), .A2(n8179), .A3(n8178), .ZN(n8335) );
  AND2_X1 U6554 ( .A1(n5692), .A2(n7097), .ZN(n5971) );
  INV_X1 U6555 ( .A(n5971), .ZN(n10063) );
  AND2_X1 U6556 ( .A1(n5128), .A2(n5127), .ZN(n5083) );
  INV_X1 U6557 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5113) );
  AND2_X1 U6558 ( .A1(n5136), .A2(n5135), .ZN(n5084) );
  AND3_X1 U6559 ( .A1(n6757), .A2(n6756), .A3(n6755), .ZN(n9355) );
  INV_X1 U6560 ( .A(n8505), .ZN(n5959) );
  NOR2_X1 U6561 ( .A1(n6213), .A2(n6194), .ZN(n5085) );
  AND2_X1 U6562 ( .A1(n8434), .A2(n8298), .ZN(n5086) );
  INV_X1 U6563 ( .A(n8380), .ZN(n8299) );
  INV_X1 U6564 ( .A(n9382), .ZN(n9379) );
  OR2_X1 U6565 ( .A1(n8964), .A2(n10068), .ZN(n5087) );
  OR2_X1 U6566 ( .A1(n9478), .A2(n9462), .ZN(n5088) );
  INV_X1 U6567 ( .A(n9939), .ZN(n7338) );
  OR2_X1 U6568 ( .A1(n8634), .A2(n7077), .ZN(n5090) );
  AND2_X1 U6569 ( .A1(n6616), .A2(n9544), .ZN(n9800) );
  AND2_X2 U6570 ( .A1(n7165), .A2(n9544), .ZN(n9617) );
  OAI21_X1 U6571 ( .B1(n8235), .B2(n8225), .A(n8242), .ZN(n8226) );
  INV_X1 U6572 ( .A(n5945), .ZN(n5939) );
  NAND2_X1 U6573 ( .A1(n5937), .A2(n5939), .ZN(n5940) );
  NAND2_X1 U6574 ( .A1(n8362), .A2(n9270), .ZN(n8298) );
  INV_X1 U6575 ( .A(n7190), .ZN(n5315) );
  INV_X1 U6576 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5191) );
  NAND2_X1 U6577 ( .A1(n7695), .A2(n6969), .ZN(n6970) );
  INV_X1 U6578 ( .A(n9983), .ZN(n7341) );
  NAND2_X1 U6579 ( .A1(n5958), .A2(n8505), .ZN(n5961) );
  AOI21_X1 U6580 ( .B1(n4334), .B2(n8389), .A(n8372), .ZN(n8373) );
  INV_X1 U6581 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n5174) );
  NAND2_X1 U6582 ( .A1(n5111), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5112) );
  INV_X1 U6583 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5370) );
  INV_X1 U6584 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5461) );
  INV_X1 U6585 ( .A(n8889), .ZN(n5574) );
  INV_X1 U6586 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n10246) );
  INV_X1 U6587 ( .A(n9106), .ZN(n6333) );
  NOR2_X1 U6588 ( .A1(n6262), .A2(n6261), .ZN(n6263) );
  INV_X1 U6589 ( .A(n8373), .ZN(n8374) );
  INV_X1 U6590 ( .A(n6440), .ZN(n6438) );
  INV_X1 U6591 ( .A(n6478), .ZN(n6476) );
  INV_X1 U6592 ( .A(n6416), .ZN(n6398) );
  NOR2_X1 U6593 ( .A1(n6178), .A2(n6857), .ZN(n6193) );
  NAND2_X1 U6594 ( .A1(n9615), .A2(n8167), .ZN(n8142) );
  INV_X1 U6595 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6006) );
  NAND2_X1 U6596 ( .A1(n6028), .A2(n6039), .ZN(n6029) );
  INV_X1 U6597 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n5181) );
  INV_X1 U6598 ( .A(SI_17_), .ZN(n5165) );
  OR2_X1 U6599 ( .A1(n8468), .A2(n8939), .ZN(n8469) );
  INV_X1 U6600 ( .A(n5763), .ZN(n5608) );
  XNOR2_X1 U6601 ( .A(n7824), .B(n7845), .ZN(n7748) );
  NAND2_X1 U6602 ( .A1(n5637), .A2(n5636), .ZN(n5649) );
  NOR2_X1 U6603 ( .A1(n8482), .A2(n10028), .ZN(n5657) );
  INV_X1 U6604 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5568) );
  INV_X1 U6605 ( .A(n5916), .ZN(n5711) );
  INV_X1 U6606 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5404) );
  AND2_X1 U6607 ( .A1(n6193), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6213) );
  INV_X1 U6608 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6298) );
  AND2_X1 U6609 ( .A1(n6213), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6250) );
  OR2_X1 U6610 ( .A1(n6526), .A2(n9174), .ZN(n6538) );
  NAND2_X1 U6611 ( .A1(n6438), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6459) );
  INV_X1 U6612 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6857) );
  NAND2_X1 U6613 ( .A1(n6398), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6418) );
  INV_X1 U6614 ( .A(n9385), .ZN(n9398) );
  NAND2_X1 U6615 ( .A1(n9760), .A2(n8171), .ZN(n8145) );
  INV_X1 U6616 ( .A(n9283), .ZN(n8138) );
  NAND2_X1 U6617 ( .A1(n9169), .A2(n9805), .ZN(n7910) );
  NAND2_X1 U6618 ( .A1(n5176), .A2(n5175), .ZN(n5179) );
  AND2_X1 U6619 ( .A1(n6245), .A2(n6229), .ZN(n6273) );
  OR2_X1 U6620 ( .A1(n8475), .A2(n8860), .ZN(n8476) );
  INV_X1 U6621 ( .A(n8606), .ZN(n8574) );
  OR2_X1 U6622 ( .A1(n5539), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5554) );
  OR2_X1 U6623 ( .A1(n6914), .A2(n6976), .ZN(n8603) );
  OR2_X1 U6624 ( .A1(n5282), .A2(n5266), .ZN(n5270) );
  NOR2_X1 U6625 ( .A1(n8657), .A2(n8656), .ZN(n8660) );
  AND2_X1 U6626 ( .A1(n6969), .A2(n8767), .ZN(n7097) );
  OR2_X1 U6627 ( .A1(n7097), .A2(n10052), .ZN(n10023) );
  OR2_X1 U6628 ( .A1(n10081), .A2(n5989), .ZN(n5990) );
  INV_X1 U6629 ( .A(n8625), .ZN(n7877) );
  OR2_X1 U6630 ( .A1(n5421), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5457) );
  AND2_X1 U6631 ( .A1(n6864), .A2(n6057), .ZN(n9145) );
  NAND2_X1 U6632 ( .A1(n6353), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6381) );
  OR2_X1 U6633 ( .A1(n6381), .A2(n6380), .ZN(n6416) );
  OR2_X1 U6634 ( .A1(n6299), .A2(n6298), .ZN(n6320) );
  OR2_X1 U6635 ( .A1(n9400), .A2(n6561), .ZN(n6566) );
  OR2_X1 U6636 ( .A1(n6418), .A2(n8134), .ZN(n6440) );
  INV_X1 U6637 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8134) );
  NAND2_X1 U6638 ( .A1(n6278), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6299) );
  OR2_X1 U6639 ( .A1(n8193), .A2(n8338), .ZN(n8367) );
  INV_X1 U6640 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6609) );
  INV_X1 U6641 ( .A(n9584), .ZN(n9585) );
  NAND2_X1 U6642 ( .A1(n9225), .A2(n8138), .ZN(n8139) );
  INV_X1 U6643 ( .A(n9881), .ZN(n7135) );
  OR2_X1 U6644 ( .A1(n7163), .A2(n8437), .ZN(n9881) );
  NOR2_X2 U6645 ( .A1(n7271), .A2(n7214), .ZN(n7510) );
  XNOR2_X1 U6646 ( .A(n9291), .B(n7290), .ZN(n8310) );
  INV_X1 U6647 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6050) );
  AND2_X1 U6648 ( .A1(n5122), .A2(n5123), .ZN(n5306) );
  INV_X1 U6649 ( .A(n8603), .ZN(n8571) );
  NAND2_X1 U6650 ( .A1(n6919), .A2(n10021), .ZN(n8615) );
  INV_X1 U6651 ( .A(n7902), .ZN(n5952) );
  AND4_X1 U6652 ( .A1(n5529), .A2(n5528), .A3(n5527), .A4(n5526), .ZN(n8924)
         );
  NOR2_X1 U6653 ( .A1(P2_U3150), .A2(n6701), .ZN(n9962) );
  AND2_X1 U6654 ( .A1(P2_U3893), .A2(n6702), .ZN(n9949) );
  NAND2_X1 U6655 ( .A1(n5981), .A2(n5647), .ZN(n8952) );
  AND2_X1 U6656 ( .A1(n8920), .A2(n8919), .ZN(n8998) );
  INV_X1 U6657 ( .A(n8959), .ZN(n8914) );
  INV_X1 U6658 ( .A(n10052), .ZN(n10080) );
  INV_X1 U6659 ( .A(n10068), .ZN(n10075) );
  AND2_X1 U6660 ( .A1(n5687), .A2(n5686), .ZN(n7061) );
  INV_X1 U6661 ( .A(n8763), .ZN(n8767) );
  INV_X1 U6662 ( .A(n9800), .ZN(n6649) );
  OR2_X1 U6663 ( .A1(n6252), .A2(n6233), .ZN(n6280) );
  INV_X1 U6664 ( .A(n9814), .ZN(n9267) );
  INV_X1 U6665 ( .A(n4333), .ZN(n6561) );
  OR2_X1 U6666 ( .A1(n9827), .A2(n8442), .ZN(n9343) );
  INV_X1 U6667 ( .A(n9343), .ZN(n9853) );
  INV_X1 U6668 ( .A(n7290), .ZN(n7607) );
  AOI21_X1 U6669 ( .B1(n6890), .B2(n6609), .A(n6715), .ZN(n7156) );
  NAND2_X1 U6670 ( .A1(n7781), .A2(n7116), .ZN(n9878) );
  AND3_X1 U6671 ( .A1(n6893), .A2(n6892), .A3(n6891), .ZN(n6904) );
  INV_X1 U6672 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10288) );
  OR2_X1 U6673 ( .A1(n6923), .A2(n6655), .ZN(n6700) );
  INV_X1 U6674 ( .A(n8520), .ZN(n9063) );
  INV_X1 U6675 ( .A(n8615), .ZN(n8596) );
  NAND2_X1 U6676 ( .A1(n5244), .A2(n5243), .ZN(n8859) );
  INV_X1 U6677 ( .A(n8604), .ZN(n8938) );
  INV_X1 U6678 ( .A(n10003), .ZN(n9958) );
  INV_X1 U6679 ( .A(n9962), .ZN(n10017) );
  NAND2_X1 U6680 ( .A1(n6735), .A2(n8643), .ZN(n10005) );
  INV_X1 U6681 ( .A(n5976), .ZN(n5977) );
  NAND2_X1 U6682 ( .A1(n10096), .A2(n10080), .ZN(n9001) );
  INV_X1 U6683 ( .A(n10096), .ZN(n10094) );
  INV_X1 U6684 ( .A(n8534), .ZN(n9055) );
  OR2_X1 U6685 ( .A1(n10082), .A2(n10068), .ZN(n9083) );
  AND2_X1 U6686 ( .A1(n5988), .A2(n5987), .ZN(n10082) );
  INV_X1 U6687 ( .A(n10119), .ZN(n6690) );
  NAND2_X1 U6688 ( .A1(n6918), .A2(n6678), .ZN(n10119) );
  INV_X1 U6689 ( .A(n8762), .ZN(n8747) );
  INV_X1 U6690 ( .A(n7834), .ZN(n7845) );
  INV_X1 U6691 ( .A(n9924), .ZN(n6741) );
  XNOR2_X1 U6692 ( .A(n6611), .B(n6028), .ZN(n6693) );
  INV_X1 U6693 ( .A(n9397), .ZN(n9271) );
  NAND2_X1 U6694 ( .A1(n6532), .A2(n6531), .ZN(n9273) );
  OR2_X1 U6695 ( .A1(n9827), .A2(n8181), .ZN(n9849) );
  INV_X1 U6696 ( .A(n9618), .ZN(n9865) );
  INV_X1 U6697 ( .A(n9868), .ZN(n9626) );
  INV_X1 U6698 ( .A(n9695), .ZN(n9686) );
  INV_X2 U6699 ( .A(n9896), .ZN(n9893) );
  INV_X1 U6700 ( .A(n9528), .ZN(n9750) );
  NAND2_X1 U6701 ( .A1(n9890), .A2(n9878), .ZN(n9774) );
  INV_X1 U6702 ( .A(n9890), .ZN(n9888) );
  AND2_X1 U6703 ( .A1(n6886), .A2(n6713), .ZN(n9871) );
  INV_X1 U6704 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9787) );
  INV_X1 U6705 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7985) );
  NOR2_X2 U6706 ( .A1(n6700), .A2(P2_U3151), .ZN(P2_U3893) );
  AND2_X1 U6707 ( .A1(n6654), .A2(n6693), .ZN(P1_U3973) );
  INV_X1 U6708 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n5696) );
  NOR2_X1 U6709 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5094) );
  NOR2_X1 U6710 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5093) );
  NOR2_X1 U6711 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5092) );
  NOR2_X1 U6712 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5091) );
  INV_X1 U6713 ( .A(n5667), .ZN(n5504) );
  INV_X1 U6714 ( .A(n7813), .ZN(n5692) );
  NAND2_X1 U6715 ( .A1(n5692), .A2(n5980), .ZN(n10052) );
  INV_X1 U6716 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5102) );
  INV_X1 U6717 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5103) );
  INV_X1 U6718 ( .A(SI_0_), .ZN(n5105) );
  MUX2_X1 U6719 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5111), .Z(n5108) );
  NAND2_X1 U6720 ( .A1(n5108), .A2(SI_2_), .ZN(n5110) );
  OAI21_X1 U6721 ( .B1(n5108), .B2(SI_2_), .A(n5110), .ZN(n5272) );
  INV_X1 U6722 ( .A(n5272), .ZN(n5109) );
  INV_X1 U6723 ( .A(n5116), .ZN(n5115) );
  INV_X1 U6724 ( .A(SI_3_), .ZN(n5114) );
  NAND2_X1 U6725 ( .A1(n5115), .A2(n5114), .ZN(n5117) );
  NAND2_X1 U6726 ( .A1(n5116), .A2(SI_3_), .ZN(n5118) );
  MUX2_X1 U6727 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5111), .Z(n5121) );
  INV_X1 U6728 ( .A(n5121), .ZN(n5120) );
  INV_X1 U6729 ( .A(SI_4_), .ZN(n5119) );
  NAND2_X1 U6730 ( .A1(n5120), .A2(n5119), .ZN(n5122) );
  NAND2_X1 U6731 ( .A1(n5121), .A2(SI_4_), .ZN(n5123) );
  MUX2_X1 U6732 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n6661), .Z(n5124) );
  NAND2_X1 U6733 ( .A1(n5124), .A2(SI_5_), .ZN(n5128) );
  INV_X1 U6734 ( .A(n5124), .ZN(n5126) );
  INV_X1 U6735 ( .A(SI_5_), .ZN(n5125) );
  NAND2_X1 U6736 ( .A1(n5126), .A2(n5125), .ZN(n5127) );
  NAND2_X1 U6737 ( .A1(n5129), .A2(SI_6_), .ZN(n5132) );
  INV_X1 U6738 ( .A(n5129), .ZN(n5131) );
  INV_X1 U6739 ( .A(SI_6_), .ZN(n5130) );
  MUX2_X1 U6740 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6661), .Z(n5133) );
  NAND2_X1 U6741 ( .A1(n5133), .A2(SI_7_), .ZN(n5136) );
  INV_X1 U6742 ( .A(n5133), .ZN(n5134) );
  INV_X1 U6743 ( .A(SI_7_), .ZN(n10287) );
  NAND2_X1 U6744 ( .A1(n5134), .A2(n10287), .ZN(n5135) );
  MUX2_X1 U6745 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n6661), .Z(n5137) );
  XNOR2_X1 U6746 ( .A(n5137), .B(SI_8_), .ZN(n5364) );
  INV_X1 U6747 ( .A(n5137), .ZN(n5139) );
  INV_X1 U6748 ( .A(SI_8_), .ZN(n5138) );
  INV_X1 U6749 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5141) );
  INV_X1 U6750 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5140) );
  MUX2_X1 U6751 ( .A(n5141), .B(n5140), .S(n6661), .Z(n5380) );
  INV_X1 U6752 ( .A(SI_9_), .ZN(n5142) );
  NAND2_X1 U6753 ( .A1(n5380), .A2(n5142), .ZN(n5396) );
  INV_X1 U6754 ( .A(n5396), .ZN(n5146) );
  INV_X1 U6755 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5143) );
  MUX2_X1 U6756 ( .A(n6759), .B(n5143), .S(n6661), .Z(n5148) );
  INV_X1 U6757 ( .A(SI_10_), .ZN(n5144) );
  NAND2_X1 U6758 ( .A1(n5148), .A2(n5144), .ZN(n5399) );
  INV_X1 U6759 ( .A(n5399), .ZN(n5145) );
  INV_X1 U6760 ( .A(n5380), .ZN(n5147) );
  NAND3_X1 U6761 ( .A1(n5399), .A2(n5147), .A3(SI_9_), .ZN(n5150) );
  INV_X1 U6762 ( .A(n5148), .ZN(n5149) );
  NAND2_X1 U6763 ( .A1(n5149), .A2(SI_10_), .ZN(n5398) );
  MUX2_X1 U6764 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6661), .Z(n5152) );
  XNOR2_X1 U6765 ( .A(n5152), .B(SI_11_), .ZN(n5418) );
  MUX2_X1 U6766 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6661), .Z(n5153) );
  NAND2_X1 U6767 ( .A1(n5153), .A2(SI_12_), .ZN(n5154) );
  OAI21_X1 U6768 ( .B1(n5153), .B2(SI_12_), .A(n5154), .ZN(n5435) );
  NAND2_X1 U6769 ( .A1(n5438), .A2(n5154), .ZN(n5454) );
  MUX2_X1 U6770 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6661), .Z(n5155) );
  NAND2_X1 U6771 ( .A1(n5155), .A2(SI_13_), .ZN(n5159) );
  INV_X1 U6772 ( .A(n5155), .ZN(n5157) );
  INV_X1 U6773 ( .A(SI_13_), .ZN(n5156) );
  NAND2_X1 U6774 ( .A1(n5157), .A2(n5156), .ZN(n5158) );
  MUX2_X1 U6775 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6661), .Z(n5471) );
  MUX2_X1 U6776 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6661), .Z(n5488) );
  INV_X1 U6777 ( .A(n5488), .ZN(n5160) );
  MUX2_X1 U6778 ( .A(n7284), .B(n5161), .S(n6661), .Z(n5501) );
  NAND2_X1 U6779 ( .A1(n5162), .A2(SI_16_), .ZN(n5163) );
  MUX2_X1 U6780 ( .A(n5164), .B(n10271), .S(n6661), .Z(n5166) );
  INV_X1 U6781 ( .A(n5166), .ZN(n5167) );
  NAND2_X1 U6782 ( .A1(n5167), .A2(SI_17_), .ZN(n5168) );
  NAND2_X1 U6783 ( .A1(n5169), .A2(n5168), .ZN(n5517) );
  MUX2_X1 U6784 ( .A(n10244), .B(n7438), .S(n6661), .Z(n5170) );
  XNOR2_X1 U6785 ( .A(n5170), .B(SI_18_), .ZN(n5532) );
  INV_X1 U6786 ( .A(n5170), .ZN(n5171) );
  NAND2_X1 U6787 ( .A1(n5171), .A2(SI_18_), .ZN(n5172) );
  MUX2_X1 U6788 ( .A(n5174), .B(n8058), .S(n6661), .Z(n5176) );
  INV_X1 U6789 ( .A(SI_19_), .ZN(n5175) );
  INV_X1 U6790 ( .A(n5176), .ZN(n5177) );
  NAND2_X1 U6791 ( .A1(n5177), .A2(SI_19_), .ZN(n5178) );
  NAND2_X1 U6792 ( .A1(n5179), .A2(n5178), .ZN(n5546) );
  MUX2_X1 U6793 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6661), .Z(n5563) );
  INV_X1 U6794 ( .A(n5563), .ZN(n5180) );
  MUX2_X1 U6795 ( .A(n5181), .B(n7707), .S(n6661), .Z(n5577) );
  NOR2_X1 U6796 ( .A1(n5182), .A2(SI_21_), .ZN(n5184) );
  NAND2_X1 U6797 ( .A1(n5182), .A2(SI_21_), .ZN(n5183) );
  INV_X1 U6798 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n5185) );
  MUX2_X1 U6799 ( .A(n5185), .B(n7855), .S(n6661), .Z(n5187) );
  INV_X1 U6800 ( .A(SI_22_), .ZN(n5186) );
  NAND2_X1 U6801 ( .A1(n5187), .A2(n5186), .ZN(n5190) );
  INV_X1 U6802 ( .A(n5187), .ZN(n5188) );
  NAND2_X1 U6803 ( .A1(n5188), .A2(SI_22_), .ZN(n5189) );
  NAND2_X1 U6804 ( .A1(n5190), .A2(n5189), .ZN(n5588) );
  MUX2_X1 U6805 ( .A(n5191), .B(n7908), .S(n6661), .Z(n5193) );
  INV_X1 U6806 ( .A(SI_23_), .ZN(n5192) );
  NAND2_X1 U6807 ( .A1(n5193), .A2(n5192), .ZN(n5196) );
  INV_X1 U6808 ( .A(n5193), .ZN(n5194) );
  NAND2_X1 U6809 ( .A1(n5194), .A2(SI_23_), .ZN(n5195) );
  NAND2_X1 U6810 ( .A1(n5196), .A2(n5195), .ZN(n5599) );
  INV_X1 U6811 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n5197) );
  MUX2_X1 U6812 ( .A(n5197), .B(n7985), .S(n6661), .Z(n5199) );
  INV_X1 U6813 ( .A(SI_24_), .ZN(n5198) );
  NAND2_X1 U6814 ( .A1(n5199), .A2(n5198), .ZN(n5202) );
  INV_X1 U6815 ( .A(n5199), .ZN(n5200) );
  NAND2_X1 U6816 ( .A1(n5200), .A2(SI_24_), .ZN(n5201) );
  NAND2_X1 U6817 ( .A1(n5232), .A2(n5233), .ZN(n5203) );
  INV_X1 U6818 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n5204) );
  INV_X1 U6819 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8031) );
  MUX2_X1 U6820 ( .A(n5204), .B(n8031), .S(n6661), .Z(n5206) );
  INV_X1 U6821 ( .A(SI_25_), .ZN(n5205) );
  NAND2_X1 U6822 ( .A1(n5206), .A2(n5205), .ZN(n5209) );
  INV_X1 U6823 ( .A(n5206), .ZN(n5207) );
  NAND2_X1 U6824 ( .A1(n5207), .A2(SI_25_), .ZN(n5208) );
  INV_X1 U6825 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n5210) );
  INV_X1 U6826 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8054) );
  MUX2_X1 U6827 ( .A(n5210), .B(n8054), .S(n6661), .Z(n5212) );
  INV_X1 U6828 ( .A(SI_26_), .ZN(n5211) );
  NAND2_X1 U6829 ( .A1(n5212), .A2(n5211), .ZN(n5215) );
  INV_X1 U6830 ( .A(n5212), .ZN(n5213) );
  NAND2_X1 U6831 ( .A1(n5213), .A2(SI_26_), .ZN(n5214) );
  NAND2_X1 U6832 ( .A1(n5216), .A2(n5215), .ZN(n5720) );
  INV_X1 U6833 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5217) );
  INV_X1 U6834 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9790) );
  MUX2_X1 U6835 ( .A(n5217), .B(n9790), .S(n6661), .Z(n5219) );
  INV_X1 U6836 ( .A(SI_27_), .ZN(n5218) );
  NAND2_X1 U6837 ( .A1(n5219), .A2(n5218), .ZN(n5721) );
  INV_X1 U6838 ( .A(n5219), .ZN(n5220) );
  NAND2_X1 U6839 ( .A1(n5220), .A2(SI_27_), .ZN(n5221) );
  NOR2_X1 U6840 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5224) );
  NAND4_X1 U6841 ( .A1(n5224), .A2(n5223), .A3(n5534), .A4(n5222), .ZN(n5226)
         );
  NAND2_X1 U6842 ( .A1(n5228), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5229) );
  NAND2_X1 U6843 ( .A1(n9099), .A2(n5787), .ZN(n5231) );
  NAND2_X1 U6844 ( .A1(n5788), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5230) );
  NAND2_X1 U6845 ( .A1(n7982), .A2(n5787), .ZN(n5235) );
  NAND2_X1 U6846 ( .A1(n5788), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5234) );
  INV_X1 U6847 ( .A(n9036), .ZN(n8851) );
  NAND2_X1 U6848 ( .A1(n5316), .A2(n7109), .ZN(n5331) );
  OR2_X2 U6849 ( .A1(n5331), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5350) );
  NAND2_X1 U6850 ( .A1(n5462), .A2(n5461), .ZN(n5481) );
  NAND2_X1 U6851 ( .A1(n5606), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5236) );
  NAND2_X1 U6852 ( .A1(n5236), .A2(n5079), .ZN(n8562) );
  NAND2_X1 U6853 ( .A1(n8562), .A2(n5607), .ZN(n5244) );
  INV_X1 U6854 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8976) );
  NAND2_X1 U6855 ( .A1(n5608), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5241) );
  NAND2_X1 U6856 ( .A1(n5753), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5240) );
  OAI211_X1 U6857 ( .C1(n5761), .C2(n8976), .A(n5241), .B(n5240), .ZN(n5242)
         );
  INV_X1 U6858 ( .A(n5242), .ZN(n5243) );
  INV_X1 U6859 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6817) );
  INV_X1 U6860 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7100) );
  INV_X1 U6861 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5245) );
  INV_X1 U6862 ( .A(n5246), .ZN(n5247) );
  NAND2_X1 U6863 ( .A1(n5248), .A2(n5247), .ZN(n5249) );
  NAND2_X1 U6864 ( .A1(n5250), .A2(n5249), .ZN(n6663) );
  NAND2_X1 U6865 ( .A1(n4330), .A2(n6663), .ZN(n5255) );
  MUX2_X1 U6866 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5251), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5254) );
  NAND2_X1 U6867 ( .A1(n5280), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5260) );
  INV_X1 U6868 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5257) );
  INV_X1 U6869 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7063) );
  OR2_X1 U6870 ( .A1(n5301), .A2(n7063), .ZN(n5258) );
  NAND2_X1 U6871 ( .A1(n6662), .A2(SI_0_), .ZN(n5262) );
  XNOR2_X1 U6872 ( .A(n5262), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9104) );
  NAND2_X1 U6873 ( .A1(n5697), .A2(n7065), .ZN(n7017) );
  NAND2_X1 U6874 ( .A1(n5770), .A2(n7017), .ZN(n5265) );
  NAND2_X1 U6875 ( .A1(n10027), .A2(n7020), .ZN(n5264) );
  NAND2_X1 U6876 ( .A1(n5265), .A2(n5264), .ZN(n10024) );
  INV_X1 U6877 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5266) );
  INV_X1 U6878 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10022) );
  INV_X1 U6879 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5267) );
  NAND2_X1 U6880 ( .A1(n5280), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5268) );
  INV_X1 U6881 ( .A(n5271), .ZN(n5273) );
  NAND2_X1 U6882 ( .A1(n5273), .A2(n5272), .ZN(n5275) );
  NAND2_X1 U6883 ( .A1(n5275), .A2(n5274), .ZN(n6670) );
  NAND2_X1 U6884 ( .A1(n5601), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5277) );
  NAND2_X1 U6885 ( .A1(n5551), .A2(n4602), .ZN(n5276) );
  INV_X1 U6886 ( .A(n6988), .ZN(n10035) );
  NAND2_X1 U6887 ( .A1(n8635), .A2(n10035), .ZN(n5814) );
  NAND2_X1 U6888 ( .A1(n10024), .A2(n5811), .ZN(n5279) );
  NAND2_X1 U6889 ( .A1(n7074), .A2(n10035), .ZN(n5278) );
  NAND2_X1 U6890 ( .A1(n5279), .A2(n5278), .ZN(n7072) );
  INV_X1 U6891 ( .A(n7072), .ZN(n5296) );
  OR2_X1 U6892 ( .A1(n5298), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5287) );
  NAND2_X1 U6893 ( .A1(n5280), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5286) );
  INV_X1 U6894 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5281) );
  OR2_X1 U6895 ( .A1(n5282), .A2(n5281), .ZN(n5285) );
  INV_X1 U6896 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5283) );
  OR2_X1 U6897 ( .A1(n5301), .A2(n5283), .ZN(n5284) );
  OR2_X1 U6898 ( .A1(n5289), .A2(n5288), .ZN(n5290) );
  NAND2_X1 U6899 ( .A1(n5291), .A2(n5290), .ZN(n6668) );
  NAND2_X1 U6900 ( .A1(n5601), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5295) );
  OR2_X1 U6901 ( .A1(n5292), .A2(n9086), .ZN(n5293) );
  XNOR2_X1 U6902 ( .A(n5293), .B(P2_IR_REG_3__SCAN_IN), .ZN(n9924) );
  NAND2_X1 U6903 ( .A1(n5551), .A2(n9924), .ZN(n5294) );
  NAND2_X1 U6904 ( .A1(n8634), .A2(n7077), .ZN(n5297) );
  AND2_X1 U6905 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5299) );
  NOR2_X1 U6906 ( .A1(n5316), .A2(n5299), .ZN(n7031) );
  OR2_X1 U6907 ( .A1(n5298), .A2(n7031), .ZN(n5305) );
  NAND2_X1 U6908 ( .A1(n5745), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5304) );
  INV_X1 U6909 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5300) );
  OR2_X1 U6910 ( .A1(n5282), .A2(n5300), .ZN(n5303) );
  INV_X1 U6911 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7188) );
  OR2_X1 U6912 ( .A1(n5301), .A2(n7188), .ZN(n5302) );
  NAND4_X1 U6913 ( .A1(n5305), .A2(n5304), .A3(n5303), .A4(n5302), .ZN(n8633)
         );
  OR2_X1 U6914 ( .A1(n5307), .A2(n5306), .ZN(n5308) );
  NAND2_X1 U6915 ( .A1(n5309), .A2(n5308), .ZN(n6667) );
  NAND2_X1 U6916 ( .A1(n5601), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5313) );
  INV_X1 U6917 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5310) );
  NAND2_X1 U6918 ( .A1(n5292), .A2(n5310), .ZN(n5326) );
  NAND2_X1 U6919 ( .A1(n5326), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5311) );
  XNOR2_X1 U6920 ( .A(n5311), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6744) );
  NAND2_X1 U6921 ( .A1(n5551), .A2(n6744), .ZN(n5312) );
  OR2_X1 U6922 ( .A1(n5316), .A2(n7109), .ZN(n5317) );
  AND2_X1 U6923 ( .A1(n5331), .A2(n5317), .ZN(n7108) );
  OR2_X1 U6924 ( .A1(n5298), .A2(n7108), .ZN(n5322) );
  NAND2_X1 U6925 ( .A1(n5745), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5321) );
  INV_X1 U6926 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5318) );
  OR2_X1 U6927 ( .A1(n5760), .A2(n5318), .ZN(n5320) );
  INV_X1 U6928 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7395) );
  OR2_X1 U6929 ( .A1(n5763), .A2(n7395), .ZN(n5319) );
  NAND4_X1 U6930 ( .A1(n5322), .A2(n5321), .A3(n5320), .A4(n5319), .ZN(n8632)
         );
  OR2_X1 U6931 ( .A1(n5323), .A2(n5083), .ZN(n5324) );
  NAND2_X1 U6932 ( .A1(n5325), .A2(n5324), .ZN(n6672) );
  NAND2_X1 U6933 ( .A1(n5601), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5329) );
  NAND2_X1 U6934 ( .A1(n5340), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U6935 ( .A1(n5551), .A2(n9939), .ZN(n5328) );
  OAI211_X1 U6936 ( .C1(n5314), .C2(n6672), .A(n5329), .B(n5328), .ZN(n7397)
         );
  NAND2_X1 U6937 ( .A1(n8632), .A2(n7397), .ZN(n5773) );
  NAND2_X1 U6938 ( .A1(n7392), .A2(n5773), .ZN(n5330) );
  INV_X1 U6939 ( .A(n7397), .ZN(n10043) );
  NAND2_X1 U6940 ( .A1(n7359), .A2(n10043), .ZN(n5774) );
  NAND2_X1 U6941 ( .A1(n5330), .A2(n5774), .ZN(n7356) );
  NAND2_X1 U6942 ( .A1(n5331), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5332) );
  AND2_X1 U6943 ( .A1(n5350), .A2(n5332), .ZN(n7360) );
  OR2_X1 U6944 ( .A1(n5298), .A2(n7360), .ZN(n5337) );
  NAND2_X1 U6945 ( .A1(n5745), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5336) );
  INV_X1 U6946 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5333) );
  OR2_X1 U6947 ( .A1(n5760), .A2(n5333), .ZN(n5335) );
  INV_X1 U6948 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7361) );
  OR2_X1 U6949 ( .A1(n5763), .A2(n7361), .ZN(n5334) );
  NOR2_X1 U6950 ( .A1(n5340), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5343) );
  NOR2_X1 U6951 ( .A1(n5343), .A2(n9086), .ZN(n5341) );
  MUX2_X1 U6952 ( .A(n9086), .B(n5341), .S(P2_IR_REG_6__SCAN_IN), .Z(n5345) );
  NAND2_X1 U6953 ( .A1(n5343), .A2(n5342), .ZN(n5359) );
  INV_X1 U6954 ( .A(n5359), .ZN(n5344) );
  OAI22_X1 U6955 ( .A1(n5358), .A2(n4573), .B1(n5263), .B2(n9959), .ZN(n5346)
         );
  NAND2_X1 U6956 ( .A1(n8631), .A2(n7363), .ZN(n5347) );
  NAND2_X1 U6957 ( .A1(n7356), .A2(n5347), .ZN(n5349) );
  INV_X1 U6958 ( .A(n7363), .ZN(n10047) );
  NAND2_X1 U6959 ( .A1(n5700), .A2(n10047), .ZN(n5348) );
  NAND2_X1 U6960 ( .A1(n5349), .A2(n5348), .ZN(n7370) );
  NAND2_X1 U6961 ( .A1(n5753), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5355) );
  INV_X1 U6962 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7317) );
  OR2_X1 U6963 ( .A1(n5761), .A2(n7317), .ZN(n5354) );
  AND2_X1 U6964 ( .A1(n5350), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5351) );
  NOR2_X1 U6965 ( .A1(n5371), .A2(n5351), .ZN(n7375) );
  OR2_X1 U6966 ( .A1(n5298), .A2(n7375), .ZN(n5353) );
  INV_X1 U6967 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7376) );
  OR2_X1 U6968 ( .A1(n5763), .A2(n7376), .ZN(n5352) );
  NAND2_X1 U6969 ( .A1(n5359), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5360) );
  AOI22_X1 U6970 ( .A1(n5788), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5551), .B2(
        n9983), .ZN(n5361) );
  NAND2_X1 U6971 ( .A1(n7495), .A2(n7378), .ZN(n5842) );
  INV_X1 U6972 ( .A(n7495), .ZN(n8630) );
  NAND2_X1 U6973 ( .A1(n10053), .A2(n8630), .ZN(n7496) );
  NAND2_X1 U6974 ( .A1(n5842), .A2(n7496), .ZN(n7371) );
  NAND2_X1 U6975 ( .A1(n7370), .A2(n7371), .ZN(n5363) );
  NAND2_X1 U6976 ( .A1(n7495), .A2(n10053), .ZN(n5362) );
  NAND2_X1 U6977 ( .A1(n5363), .A2(n5362), .ZN(n7493) );
  XNOR2_X1 U6978 ( .A(n5365), .B(n5364), .ZN(n6685) );
  NAND2_X1 U6979 ( .A1(n6685), .A2(n5787), .ZN(n5369) );
  OR2_X1 U6980 ( .A1(n5366), .A2(n9086), .ZN(n5367) );
  XNOR2_X1 U6981 ( .A(n5367), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10002) );
  AOI22_X1 U6982 ( .A1(n5788), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5551), .B2(
        n10002), .ZN(n5368) );
  NAND2_X1 U6983 ( .A1(n5745), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5377) );
  NOR2_X1 U6984 ( .A1(n5371), .A2(n5370), .ZN(n5372) );
  OR2_X1 U6985 ( .A1(n5386), .A2(n5372), .ZN(n7499) );
  NAND2_X1 U6986 ( .A1(n5607), .A2(n7499), .ZN(n5376) );
  INV_X1 U6987 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5373) );
  OR2_X1 U6988 ( .A1(n5760), .A2(n5373), .ZN(n5375) );
  INV_X1 U6989 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7343) );
  OR2_X1 U6990 ( .A1(n5763), .A2(n7343), .ZN(n5374) );
  NAND4_X1 U6991 ( .A1(n5377), .A2(n5376), .A3(n5375), .A4(n5374), .ZN(n8629)
         );
  NOR2_X1 U6992 ( .A1(n7560), .A2(n8629), .ZN(n5379) );
  NAND2_X1 U6993 ( .A1(n7560), .A2(n8629), .ZN(n5378) );
  XNOR2_X1 U6994 ( .A(n5380), .B(SI_9_), .ZN(n5395) );
  NAND2_X1 U6995 ( .A1(n6709), .A2(n5787), .ZN(n5384) );
  NAND2_X1 U6996 ( .A1(n5366), .A2(n5381), .ZN(n5402) );
  NAND2_X1 U6997 ( .A1(n5402), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5382) );
  XNOR2_X1 U6998 ( .A(n5382), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7421) );
  AOI22_X1 U6999 ( .A1(n5788), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5551), .B2(
        n7421), .ZN(n5383) );
  OR2_X1 U7000 ( .A1(n5386), .A2(n5385), .ZN(n5387) );
  AND2_X1 U7001 ( .A1(n5409), .A2(n5387), .ZN(n7621) );
  OR2_X1 U7002 ( .A1(n4338), .A2(n7621), .ZN(n5393) );
  NAND2_X1 U7003 ( .A1(n5745), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5392) );
  INV_X1 U7004 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5388) );
  OR2_X1 U7005 ( .A1(n5760), .A2(n5388), .ZN(n5391) );
  INV_X1 U7006 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5389) );
  OR2_X1 U7007 ( .A1(n5763), .A2(n5389), .ZN(n5390) );
  NAND4_X1 U7008 ( .A1(n5393), .A2(n5392), .A3(n5391), .A4(n5390), .ZN(n8628)
         );
  AND2_X1 U7009 ( .A1(n10062), .A2(n8628), .ZN(n5394) );
  NAND2_X1 U7010 ( .A1(n5397), .A2(n5396), .ZN(n5401) );
  AND2_X1 U7011 ( .A1(n5399), .A2(n5398), .ZN(n5400) );
  XNOR2_X1 U7012 ( .A(n5401), .B(n5400), .ZN(n6716) );
  NAND2_X1 U7013 ( .A1(n6716), .A2(n5787), .ZN(n5408) );
  NOR2_X1 U7014 ( .A1(n5402), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5405) );
  OR2_X1 U7015 ( .A1(n5405), .A2(n9086), .ZN(n5403) );
  MUX2_X1 U7016 ( .A(n5403), .B(P2_IR_REG_31__SCAN_IN), .S(n5404), .Z(n5406)
         );
  NAND2_X1 U7017 ( .A1(n5405), .A2(n5404), .ZN(n5421) );
  AOI22_X1 U7018 ( .A1(n5788), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5551), .B2(
        n7429), .ZN(n5407) );
  NAND2_X1 U7019 ( .A1(n5408), .A2(n5407), .ZN(n10067) );
  NAND2_X1 U7020 ( .A1(n5409), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5410) );
  AND2_X1 U7021 ( .A1(n5426), .A2(n5410), .ZN(n7731) );
  OR2_X1 U7022 ( .A1(n5298), .A2(n7731), .ZN(n5415) );
  NAND2_X1 U7023 ( .A1(n5745), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5414) );
  INV_X1 U7024 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5411) );
  OR2_X1 U7025 ( .A1(n5760), .A2(n5411), .ZN(n5413) );
  INV_X1 U7026 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7732) );
  OR2_X1 U7027 ( .A1(n5763), .A2(n7732), .ZN(n5412) );
  NAND4_X1 U7028 ( .A1(n5415), .A2(n5414), .A3(n5413), .A4(n5412), .ZN(n8627)
         );
  NOR2_X1 U7029 ( .A1(n10067), .A2(n8627), .ZN(n5416) );
  NAND2_X1 U7030 ( .A1(n10067), .A2(n8627), .ZN(n5417) );
  XNOR2_X1 U7031 ( .A(n5419), .B(n5418), .ZN(n6822) );
  NAND2_X1 U7032 ( .A1(n6822), .A2(n5787), .ZN(n5424) );
  NAND2_X1 U7033 ( .A1(n5421), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5420) );
  MUX2_X1 U7034 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5420), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n5422) );
  AOI22_X1 U7035 ( .A1(n5788), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5551), .B2(
        n7834), .ZN(n5423) );
  NAND2_X1 U7036 ( .A1(n5424), .A2(n5423), .ZN(n10072) );
  NAND2_X1 U7037 ( .A1(n5753), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5432) );
  INV_X1 U7038 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5425) );
  OR2_X1 U7039 ( .A1(n5761), .A2(n5425), .ZN(n5431) );
  NAND2_X1 U7040 ( .A1(n5426), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5427) );
  AND2_X1 U7041 ( .A1(n5443), .A2(n5427), .ZN(n7820) );
  OR2_X1 U7042 ( .A1(n5298), .A2(n7820), .ZN(n5430) );
  INV_X1 U7043 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5428) );
  OR2_X1 U7044 ( .A1(n5763), .A2(n5428), .ZN(n5429) );
  OR2_X1 U7045 ( .A1(n10072), .A2(n7894), .ZN(n5857) );
  NAND2_X1 U7046 ( .A1(n10072), .A2(n7894), .ZN(n5856) );
  NAND2_X1 U7047 ( .A1(n5857), .A2(n5856), .ZN(n7816) );
  INV_X1 U7048 ( .A(n7894), .ZN(n8626) );
  NAND2_X1 U7049 ( .A1(n10072), .A2(n8626), .ZN(n5433) );
  NAND2_X1 U7050 ( .A1(n5434), .A2(n5433), .ZN(n7891) );
  INV_X1 U7051 ( .A(n7891), .ZN(n5451) );
  NAND2_X1 U7052 ( .A1(n5436), .A2(n5435), .ZN(n5437) );
  NAND2_X1 U7053 ( .A1(n5438), .A2(n5437), .ZN(n6846) );
  OR2_X1 U7054 ( .A1(n6846), .A2(n5314), .ZN(n5441) );
  NAND2_X1 U7055 ( .A1(n5457), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5439) );
  XNOR2_X1 U7056 ( .A(n5439), .B(n10273), .ZN(n7949) );
  INV_X1 U7057 ( .A(n7949), .ZN(n7843) );
  AOI22_X1 U7058 ( .A1(n5788), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5551), .B2(
        n7843), .ZN(n5440) );
  INV_X1 U7059 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n5442) );
  OR2_X1 U7060 ( .A1(n5761), .A2(n5442), .ZN(n5450) );
  AND2_X1 U7061 ( .A1(n5443), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5444) );
  NOR2_X1 U7062 ( .A1(n5462), .A2(n5444), .ZN(n7895) );
  OR2_X1 U7063 ( .A1(n4338), .A2(n7895), .ZN(n5449) );
  INV_X1 U7064 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n5445) );
  OR2_X1 U7065 ( .A1(n5760), .A2(n5445), .ZN(n5448) );
  INV_X1 U7066 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n5446) );
  OR2_X1 U7067 ( .A1(n5763), .A2(n5446), .ZN(n5447) );
  NAND4_X1 U7068 ( .A1(n5450), .A2(n5449), .A3(n5448), .A4(n5447), .ZN(n8625)
         );
  NAND2_X1 U7069 ( .A1(n5451), .A2(n4413), .ZN(n5453) );
  INV_X1 U7070 ( .A(n10079), .ZN(n5703) );
  NAND2_X1 U7071 ( .A1(n5703), .A2(n7877), .ZN(n5452) );
  OR2_X1 U7072 ( .A1(n5454), .A2(n4354), .ZN(n5455) );
  AND2_X1 U7073 ( .A1(n5455), .A2(n5456), .ZN(n6994) );
  NAND2_X1 U7074 ( .A1(n6994), .A2(n5787), .ZN(n5460) );
  NAND2_X1 U7075 ( .A1(n5458), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5474) );
  XNOR2_X1 U7076 ( .A(n5474), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8655) );
  AOI22_X1 U7077 ( .A1(n5788), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5551), .B2(
        n8655), .ZN(n5459) );
  OR2_X1 U7078 ( .A1(n5462), .A2(n5461), .ZN(n5463) );
  AND2_X1 U7079 ( .A1(n5463), .A2(n5481), .ZN(n8004) );
  OR2_X1 U7080 ( .A1(n4338), .A2(n8004), .ZN(n5469) );
  NAND2_X1 U7081 ( .A1(n5745), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5468) );
  INV_X1 U7082 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n5464) );
  OR2_X1 U7083 ( .A1(n5760), .A2(n5464), .ZN(n5467) );
  INV_X1 U7084 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5465) );
  OR2_X1 U7085 ( .A1(n5763), .A2(n5465), .ZN(n5466) );
  NAND4_X1 U7086 ( .A1(n5469), .A2(n5468), .A3(n5467), .A4(n5466), .ZN(n8624)
         );
  NOR2_X1 U7087 ( .A1(n8016), .A2(n8624), .ZN(n5867) );
  NAND2_X1 U7088 ( .A1(n8016), .A2(n8624), .ZN(n5769) );
  XNOR2_X1 U7089 ( .A(n5471), .B(SI_14_), .ZN(n5472) );
  XNOR2_X1 U7090 ( .A(n5470), .B(n5472), .ZN(n7043) );
  NAND2_X1 U7091 ( .A1(n7043), .A2(n5787), .ZN(n5480) );
  INV_X1 U7092 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U7093 ( .A1(n5474), .A2(n5473), .ZN(n5475) );
  NAND2_X1 U7094 ( .A1(n5475), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5477) );
  INV_X1 U7095 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5476) );
  NAND2_X1 U7096 ( .A1(n5477), .A2(n5476), .ZN(n5491) );
  OR2_X1 U7097 ( .A1(n5477), .A2(n5476), .ZN(n5478) );
  INV_X1 U7098 ( .A(n8681), .ZN(n8653) );
  AOI22_X1 U7099 ( .A1(n5788), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5551), .B2(
        n8653), .ZN(n5479) );
  INV_X1 U7100 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10138) );
  OR2_X1 U7101 ( .A1(n5761), .A2(n10138), .ZN(n5486) );
  NAND2_X1 U7102 ( .A1(n5481), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5482) );
  AND2_X1 U7103 ( .A1(n4352), .A2(n5482), .ZN(n7997) );
  OR2_X1 U7104 ( .A1(n5298), .A2(n7997), .ZN(n5485) );
  INV_X1 U7105 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8020) );
  OR2_X1 U7106 ( .A1(n5760), .A2(n8020), .ZN(n5484) );
  INV_X1 U7107 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7998) );
  OR2_X1 U7108 ( .A1(n5763), .A2(n7998), .ZN(n5483) );
  NAND4_X1 U7109 ( .A1(n5486), .A2(n5485), .A3(n5484), .A4(n5483), .ZN(n8623)
         );
  AND2_X1 U7110 ( .A1(n8024), .A2(n8623), .ZN(n5487) );
  XNOR2_X1 U7111 ( .A(n5488), .B(SI_15_), .ZN(n5489) );
  XNOR2_X1 U7112 ( .A(n5490), .B(n5489), .ZN(n7180) );
  NAND2_X1 U7113 ( .A1(n7180), .A2(n5787), .ZN(n5494) );
  NAND2_X1 U7114 ( .A1(n5491), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5492) );
  XNOR2_X1 U7115 ( .A(n5492), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8699) );
  AOI22_X1 U7116 ( .A1(n5788), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5551), .B2(
        n8699), .ZN(n5493) );
  INV_X1 U7117 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8667) );
  OR2_X1 U7118 ( .A1(n5761), .A2(n8667), .ZN(n5499) );
  AND2_X1 U7119 ( .A1(n4352), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5495) );
  NOR2_X1 U7120 ( .A1(n5509), .A2(n5495), .ZN(n8609) );
  OR2_X1 U7121 ( .A1(n5298), .A2(n8609), .ZN(n5498) );
  INV_X1 U7122 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8040) );
  OR2_X1 U7123 ( .A1(n5760), .A2(n8040), .ZN(n5497) );
  INV_X1 U7124 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8049) );
  OR2_X1 U7125 ( .A1(n5763), .A2(n8049), .ZN(n5496) );
  NAND4_X1 U7126 ( .A1(n5499), .A2(n5498), .A3(n5497), .A4(n5496), .ZN(n8948)
         );
  NOR2_X1 U7127 ( .A1(n8616), .A2(n8948), .ZN(n5779) );
  XNOR2_X1 U7128 ( .A(n5501), .B(SI_16_), .ZN(n5502) );
  NAND2_X1 U7129 ( .A1(n7245), .A2(n5787), .ZN(n5507) );
  NAND2_X1 U7130 ( .A1(n5504), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5503) );
  MUX2_X1 U7131 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5503), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5505) );
  OR2_X1 U7132 ( .A1(n5504), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5519) );
  AND2_X1 U7133 ( .A1(n5505), .A2(n5519), .ZN(n8702) );
  AOI22_X1 U7134 ( .A1(n5788), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5551), .B2(
        n8702), .ZN(n5506) );
  NAND2_X1 U7135 ( .A1(n5753), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5514) );
  INV_X1 U7136 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9005) );
  OR2_X1 U7137 ( .A1(n5761), .A2(n9005), .ZN(n5513) );
  NOR2_X1 U7138 ( .A1(n5509), .A2(n5508), .ZN(n5510) );
  OR2_X1 U7139 ( .A1(n5524), .A2(n5510), .ZN(n8954) );
  INV_X1 U7140 ( .A(n8954), .ZN(n8548) );
  OR2_X1 U7141 ( .A1(n4338), .A2(n8548), .ZN(n5512) );
  INV_X1 U7142 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8953) );
  OR2_X1 U7143 ( .A1(n5763), .A2(n8953), .ZN(n5511) );
  NAND2_X1 U7144 ( .A1(n9080), .A2(n8604), .ZN(n5884) );
  NAND2_X1 U7145 ( .A1(n5882), .A2(n5884), .ZN(n8946) );
  NAND2_X1 U7146 ( .A1(n8947), .A2(n8946), .ZN(n5516) );
  NAND2_X1 U7147 ( .A1(n9080), .A2(n8938), .ZN(n5515) );
  NAND2_X1 U7148 ( .A1(n5516), .A2(n5515), .ZN(n8937) );
  XNOR2_X1 U7149 ( .A(n5518), .B(n5517), .ZN(n7267) );
  NAND2_X1 U7150 ( .A1(n7267), .A2(n5787), .ZN(n5522) );
  NAND2_X1 U7151 ( .A1(n5519), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5520) );
  XNOR2_X1 U7152 ( .A(n5520), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8744) );
  AOI22_X1 U7153 ( .A1(n5788), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5551), .B2(
        n8744), .ZN(n5521) );
  OR2_X1 U7154 ( .A1(n5524), .A2(n5523), .ZN(n5525) );
  NAND2_X1 U7155 ( .A1(n5539), .A2(n5525), .ZN(n8942) );
  NAND2_X1 U7156 ( .A1(n5607), .A2(n8942), .ZN(n5529) );
  INV_X1 U7157 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9002) );
  OR2_X1 U7158 ( .A1(n5761), .A2(n9002), .ZN(n5528) );
  INV_X1 U7159 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9072) );
  OR2_X1 U7160 ( .A1(n5760), .A2(n9072), .ZN(n5527) );
  INV_X1 U7161 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8941) );
  OR2_X1 U7162 ( .A1(n5763), .A2(n8941), .ZN(n5526) );
  NAND2_X1 U7163 ( .A1(n9073), .A2(n8924), .ZN(n5901) );
  NAND2_X1 U7164 ( .A1(n5885), .A2(n5901), .ZN(n5880) );
  NAND2_X1 U7165 ( .A1(n8937), .A2(n5880), .ZN(n5531) );
  INV_X1 U7166 ( .A(n8924), .ZN(n8950) );
  NAND2_X1 U7167 ( .A1(n9073), .A2(n8950), .ZN(n5530) );
  NAND2_X1 U7168 ( .A1(n5531), .A2(n5530), .ZN(n8922) );
  XNOR2_X1 U7169 ( .A(n5533), .B(n5532), .ZN(n7433) );
  NAND2_X1 U7170 ( .A1(n7433), .A2(n5787), .ZN(n5538) );
  NAND2_X1 U7171 ( .A1(n5535), .A2(n5534), .ZN(n5548) );
  OR2_X1 U7172 ( .A1(n5535), .A2(n5534), .ZN(n5536) );
  AND2_X1 U7173 ( .A1(n5548), .A2(n5536), .ZN(n8762) );
  AOI22_X1 U7174 ( .A1(n5788), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5551), .B2(
        n8762), .ZN(n5537) );
  NAND2_X1 U7175 ( .A1(n5745), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U7176 ( .A1(n5539), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5540) );
  NAND2_X1 U7177 ( .A1(n5554), .A2(n5540), .ZN(n8927) );
  NAND2_X1 U7178 ( .A1(n5607), .A2(n8927), .ZN(n5543) );
  INV_X1 U7179 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9068) );
  OR2_X1 U7180 ( .A1(n5760), .A2(n9068), .ZN(n5542) );
  INV_X1 U7181 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8929) );
  OR2_X1 U7182 ( .A1(n5763), .A2(n8929), .ZN(n5541) );
  NAND4_X1 U7183 ( .A1(n5544), .A2(n5543), .A3(n5542), .A4(n5541), .ZN(n8939)
         );
  AND2_X1 U7184 ( .A1(n8931), .A2(n8939), .ZN(n5545) );
  XNOR2_X1 U7185 ( .A(n5547), .B(n5546), .ZN(n7435) );
  NAND2_X1 U7186 ( .A1(n7435), .A2(n5787), .ZN(n5553) );
  NAND2_X1 U7187 ( .A1(n5548), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5550) );
  INV_X1 U7188 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5549) );
  AOI22_X1 U7189 ( .A1(n5788), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8767), .B2(
        n5551), .ZN(n5552) );
  AND2_X1 U7190 ( .A1(n5554), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5555) );
  OR2_X1 U7191 ( .A1(n5555), .A2(n5569), .ZN(n8908) );
  NAND2_X1 U7192 ( .A1(n8908), .A2(n5607), .ZN(n5561) );
  INV_X1 U7193 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n10291) );
  OR2_X1 U7194 ( .A1(n5761), .A2(n10291), .ZN(n5558) );
  INV_X1 U7195 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n5556) );
  OR2_X1 U7196 ( .A1(n5760), .A2(n5556), .ZN(n5557) );
  AND2_X1 U7197 ( .A1(n5558), .A2(n5557), .ZN(n5560) );
  INV_X1 U7198 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8911) );
  OR2_X1 U7199 ( .A1(n5763), .A2(n8911), .ZN(n5559) );
  NAND2_X1 U7200 ( .A1(n8520), .A2(n8925), .ZN(n5907) );
  XNOR2_X1 U7201 ( .A(n5563), .B(n5562), .ZN(n5564) );
  XNOR2_X1 U7202 ( .A(n5565), .B(n5564), .ZN(n7601) );
  NAND2_X1 U7203 ( .A1(n7601), .A2(n5787), .ZN(n5567) );
  NAND2_X1 U7204 ( .A1(n5788), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5566) );
  NOR2_X1 U7205 ( .A1(n5569), .A2(n5568), .ZN(n5570) );
  OR2_X1 U7206 ( .A1(n5583), .A2(n5570), .ZN(n8897) );
  NAND2_X1 U7207 ( .A1(n8897), .A2(n5607), .ZN(n5573) );
  AOI22_X1 U7208 ( .A1(n5745), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n5753), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U7209 ( .A1(n5608), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5571) );
  NAND2_X1 U7210 ( .A1(n9058), .A2(n8904), .ZN(n8880) );
  INV_X1 U7211 ( .A(n8904), .ZN(n8621) );
  OR2_X1 U7212 ( .A1(n9058), .A2(n8621), .ZN(n5576) );
  XNOR2_X1 U7213 ( .A(n5577), .B(SI_21_), .ZN(n5578) );
  XNOR2_X1 U7214 ( .A(n5579), .B(n5578), .ZN(n7694) );
  NAND2_X1 U7215 ( .A1(n7694), .A2(n5787), .ZN(n5581) );
  NAND2_X1 U7216 ( .A1(n5788), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5580) );
  OR2_X1 U7217 ( .A1(n5583), .A2(n5582), .ZN(n5584) );
  NAND2_X1 U7218 ( .A1(n5592), .A2(n5584), .ZN(n8884) );
  NAND2_X1 U7219 ( .A1(n8884), .A2(n5607), .ZN(n5587) );
  AOI22_X1 U7220 ( .A1(n5745), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n5753), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n5586) );
  NAND2_X1 U7221 ( .A1(n5608), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U7222 ( .A1(n8534), .A2(n8893), .ZN(n5888) );
  NAND2_X1 U7223 ( .A1(n5893), .A2(n5888), .ZN(n8882) );
  XNOR2_X1 U7224 ( .A(n5589), .B(n5588), .ZN(n7812) );
  NAND2_X1 U7225 ( .A1(n7812), .A2(n5787), .ZN(n5591) );
  NAND2_X1 U7226 ( .A1(n5788), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5590) );
  NAND2_X1 U7227 ( .A1(n5592), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U7228 ( .A1(n5604), .A2(n5593), .ZN(n8869) );
  NAND2_X1 U7229 ( .A1(n8869), .A2(n5607), .ZN(n5598) );
  INV_X1 U7230 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n10158) );
  NAND2_X1 U7231 ( .A1(n5608), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U7232 ( .A1(n5745), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5594) );
  OAI211_X1 U7233 ( .C1(n5760), .C2(n10158), .A(n5595), .B(n5594), .ZN(n5596)
         );
  INV_X1 U7234 ( .A(n5596), .ZN(n5597) );
  NAND2_X1 U7235 ( .A1(n9047), .A2(n8877), .ZN(n5897) );
  NAND2_X1 U7236 ( .A1(n7906), .A2(n5787), .ZN(n5603) );
  NAND2_X1 U7237 ( .A1(n5601), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5602) );
  NAND2_X1 U7238 ( .A1(n5604), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U7239 ( .A1(n5606), .A2(n5605), .ZN(n8863) );
  NAND2_X1 U7240 ( .A1(n8863), .A2(n5607), .ZN(n5613) );
  INV_X1 U7241 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8979) );
  NAND2_X1 U7242 ( .A1(n5608), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5610) );
  NAND2_X1 U7243 ( .A1(n5753), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5609) );
  OAI211_X1 U7244 ( .C1(n5761), .C2(n8979), .A(n5610), .B(n5609), .ZN(n5611)
         );
  INV_X1 U7245 ( .A(n5611), .ZN(n5612) );
  AOI21_X1 U7246 ( .B1(n8859), .B2(n9036), .A(n8846), .ZN(n5614) );
  NAND2_X1 U7247 ( .A1(n8028), .A2(n5787), .ZN(n5618) );
  NAND2_X1 U7248 ( .A1(n5788), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U7249 ( .A1(n5745), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5623) );
  INV_X1 U7250 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9029) );
  OR2_X1 U7251 ( .A1(n5760), .A2(n9029), .ZN(n5622) );
  AOI21_X1 U7252 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n5079), .A(n5628), .ZN(
        n8835) );
  OR2_X1 U7253 ( .A1(n5298), .A2(n8835), .ZN(n5621) );
  INV_X1 U7254 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n5619) );
  OR2_X1 U7255 ( .A1(n5763), .A2(n5619), .ZN(n5620) );
  NAND2_X1 U7256 ( .A1(n9030), .A2(n8823), .ZN(n5924) );
  OAI22_X1 U7257 ( .A1(n8832), .A2(n8831), .B1(n8847), .B2(n9030), .ZN(n8820)
         );
  NAND2_X1 U7258 ( .A1(n8043), .A2(n5787), .ZN(n5626) );
  NAND2_X1 U7259 ( .A1(n5788), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5625) );
  INV_X1 U7260 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U7261 ( .A1(n5627), .A2(n5628), .ZN(n5638) );
  INV_X1 U7262 ( .A(n5628), .ZN(n5629) );
  NAND2_X1 U7263 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(n5629), .ZN(n5630) );
  NAND2_X1 U7264 ( .A1(n5745), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5633) );
  INV_X1 U7265 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9023) );
  OR2_X1 U7266 ( .A1(n5760), .A2(n9023), .ZN(n5632) );
  INV_X1 U7267 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8825) );
  OR2_X1 U7268 ( .A1(n5763), .A2(n8825), .ZN(n5631) );
  NOR2_X1 U7269 ( .A1(n9024), .A2(n8833), .ZN(n5635) );
  INV_X1 U7270 ( .A(n9024), .ZN(n8970) );
  NAND2_X1 U7271 ( .A1(n5745), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5643) );
  INV_X1 U7272 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9019) );
  OR2_X1 U7273 ( .A1(n5760), .A2(n9019), .ZN(n5642) );
  INV_X1 U7274 ( .A(n5638), .ZN(n5637) );
  INV_X1 U7275 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5636) );
  NAND2_X1 U7276 ( .A1(n5638), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5639) );
  OR2_X1 U7277 ( .A1(n4338), .A2(n8813), .ZN(n5641) );
  INV_X1 U7278 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8814) );
  OR2_X1 U7279 ( .A1(n5763), .A2(n8814), .ZN(n5640) );
  NAND2_X1 U7280 ( .A1(n8816), .A2(n8824), .ZN(n5934) );
  NAND2_X1 U7281 ( .A1(n5935), .A2(n5934), .ZN(n5956) );
  XNOR2_X1 U7282 ( .A(n5957), .B(n5956), .ZN(n5660) );
  NAND2_X1 U7283 ( .A1(n7813), .A2(n8767), .ZN(n5981) );
  MUX2_X1 U7284 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5644), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n5646) );
  NAND2_X1 U7285 ( .A1(n5646), .A2(n5645), .ZN(n6969) );
  INV_X1 U7286 ( .A(n6969), .ZN(n7563) );
  NAND2_X1 U7287 ( .A1(n7695), .A2(n7563), .ZN(n5647) );
  NAND2_X1 U7288 ( .A1(n5745), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5654) );
  INV_X1 U7289 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5648) );
  OR2_X1 U7290 ( .A1(n5760), .A2(n5648), .ZN(n5653) );
  NAND2_X1 U7291 ( .A1(n5649), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5650) );
  OR2_X1 U7292 ( .A1(n5298), .A2(n8803), .ZN(n5652) );
  INV_X1 U7293 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8804) );
  OR2_X1 U7294 ( .A1(n5763), .A2(n8804), .ZN(n5651) );
  OAI21_X1 U7295 ( .B1(n6702), .B2(n8643), .A(n5263), .ZN(n5953) );
  AOI21_X1 U7296 ( .B1(n10080), .B2(n8816), .A(n8812), .ZN(n9018) );
  AND2_X1 U7297 ( .A1(n6922), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6681) );
  NAND2_X1 U7298 ( .A1(n5664), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5665) );
  INV_X1 U7299 ( .A(n5689), .ZN(n7983) );
  NAND2_X1 U7300 ( .A1(n5669), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5671) );
  MUX2_X1 U7301 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5671), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5672) );
  NAND3_X1 U7302 ( .A1(n8044), .A2(n7983), .A3(n8029), .ZN(n6923) );
  NOR2_X1 U7303 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .ZN(
        n5676) );
  NOR4_X1 U7304 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n5675) );
  NOR4_X1 U7305 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_31__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n5674) );
  NOR4_X1 U7306 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5673) );
  NAND4_X1 U7307 ( .A1(n5676), .A2(n5675), .A3(n5674), .A4(n5673), .ZN(n5684)
         );
  NOR4_X1 U7308 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n5680) );
  NOR4_X1 U7309 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5679) );
  NOR4_X1 U7310 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5678) );
  NOR4_X1 U7311 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n5677) );
  NAND4_X1 U7312 ( .A1(n5680), .A2(n5679), .A3(n5678), .A4(n5677), .ZN(n5683)
         );
  XNOR2_X1 U7313 ( .A(n5689), .B(P2_B_REG_SCAN_IN), .ZN(n5681) );
  INV_X1 U7314 ( .A(n8029), .ZN(n5685) );
  NAND2_X1 U7315 ( .A1(n5681), .A2(n5685), .ZN(n5682) );
  OAI21_X1 U7316 ( .B1(n5684), .B2(n5683), .A(n5688), .ZN(n5984) );
  NAND2_X1 U7317 ( .A1(n6656), .A2(n6973), .ZN(n6924) );
  AND3_X1 U7318 ( .A1(n6918), .A2(n5984), .A3(n6924), .ZN(n7058) );
  INV_X1 U7319 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6675) );
  NAND2_X1 U7320 ( .A1(n5688), .A2(n6675), .ZN(n5687) );
  INV_X1 U7321 ( .A(n8044), .ZN(n5690) );
  NAND2_X1 U7322 ( .A1(n5690), .A2(n5685), .ZN(n5686) );
  INV_X1 U7323 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6682) );
  NAND2_X1 U7324 ( .A1(n5688), .A2(n6682), .ZN(n5691) );
  NAND2_X1 U7325 ( .A1(n5690), .A2(n5689), .ZN(n6679) );
  INV_X1 U7326 ( .A(n6972), .ZN(n7060) );
  NAND2_X1 U7327 ( .A1(n7061), .A2(n7060), .ZN(n5979) );
  NAND2_X1 U7328 ( .A1(n5971), .A2(n5980), .ZN(n6916) );
  NAND2_X1 U7329 ( .A1(n7813), .A2(n8763), .ZN(n5714) );
  OR2_X1 U7330 ( .A1(n5714), .A2(n6969), .ZN(n5693) );
  NAND2_X1 U7331 ( .A1(n5693), .A2(n5986), .ZN(n5695) );
  NAND2_X1 U7332 ( .A1(n7061), .A2(n5695), .ZN(n5694) );
  MUX2_X1 U7333 ( .A(n5696), .B(n9018), .S(n10096), .Z(n5718) );
  INV_X1 U7334 ( .A(n5697), .ZN(n5698) );
  NAND2_X1 U7335 ( .A1(n10029), .A2(n7077), .ZN(n5824) );
  INV_X1 U7336 ( .A(n7077), .ZN(n7224) );
  NAND2_X1 U7337 ( .A1(n8634), .A2(n7224), .ZN(n5819) );
  NAND2_X1 U7338 ( .A1(n7070), .A2(n7071), .ZN(n7069) );
  NAND2_X1 U7339 ( .A1(n7069), .A2(n5824), .ZN(n7184) );
  NAND2_X1 U7340 ( .A1(n8633), .A2(n5315), .ZN(n5826) );
  NAND2_X1 U7341 ( .A1(n7184), .A2(n5826), .ZN(n5699) );
  NAND2_X1 U7342 ( .A1(n7110), .A2(n7190), .ZN(n5820) );
  NAND2_X1 U7343 ( .A1(n8632), .A2(n10043), .ZN(n5825) );
  NAND2_X1 U7344 ( .A1(n7391), .A2(n5825), .ZN(n7354) );
  NAND2_X1 U7345 ( .A1(n5700), .A2(n7363), .ZN(n5802) );
  NAND2_X1 U7346 ( .A1(n7359), .A2(n7397), .ZN(n7353) );
  AND2_X1 U7347 ( .A1(n5802), .A2(n7353), .ZN(n5831) );
  NAND2_X1 U7348 ( .A1(n7354), .A2(n5831), .ZN(n5701) );
  NAND2_X1 U7349 ( .A1(n8631), .A2(n10047), .ZN(n5829) );
  NAND2_X1 U7350 ( .A1(n5701), .A2(n5829), .ZN(n7368) );
  INV_X1 U7351 ( .A(n7371), .ZN(n7367) );
  OR2_X1 U7352 ( .A1(n7560), .A2(n7475), .ZN(n5839) );
  AND2_X1 U7353 ( .A1(n5839), .A2(n7496), .ZN(n5837) );
  NAND2_X1 U7354 ( .A1(n7560), .A2(n7475), .ZN(n5843) );
  OR2_X1 U7355 ( .A1(n10062), .A2(n7595), .ZN(n7723) );
  NAND2_X1 U7356 ( .A1(n10062), .A2(n7595), .ZN(n5844) );
  NAND2_X1 U7357 ( .A1(n7723), .A2(n5844), .ZN(n5838) );
  OR2_X1 U7358 ( .A1(n10067), .A2(n7819), .ZN(n5852) );
  AND2_X1 U7359 ( .A1(n5852), .A2(n7723), .ZN(n5841) );
  NAND2_X1 U7360 ( .A1(n10067), .A2(n7819), .ZN(n5853) );
  INV_X1 U7361 ( .A(n7816), .ZN(n5778) );
  XNOR2_X1 U7362 ( .A(n10079), .B(n7877), .ZN(n7897) );
  NAND2_X1 U7363 ( .A1(n5703), .A2(n8625), .ZN(n5862) );
  INV_X1 U7364 ( .A(n8624), .ZN(n7893) );
  NAND2_X1 U7365 ( .A1(n8016), .A2(n7893), .ZN(n5704) );
  INV_X1 U7366 ( .A(n8016), .ZN(n8005) );
  NAND2_X1 U7367 ( .A1(n8005), .A2(n8624), .ZN(n5705) );
  INV_X1 U7368 ( .A(n8623), .ZN(n7972) );
  NAND2_X1 U7369 ( .A1(n8024), .A2(n7972), .ZN(n5871) );
  OR2_X1 U7370 ( .A1(n8024), .A2(n7972), .ZN(n5876) );
  INV_X1 U7371 ( .A(n8948), .ZN(n5706) );
  NAND2_X1 U7372 ( .A1(n8616), .A2(n5706), .ZN(n5801) );
  OR2_X1 U7373 ( .A1(n8616), .A2(n5706), .ZN(n5873) );
  NAND2_X1 U7374 ( .A1(n5707), .A2(n5873), .ZN(n8945) );
  NAND2_X1 U7375 ( .A1(n8945), .A2(n5884), .ZN(n5708) );
  INV_X1 U7376 ( .A(n8939), .ZN(n8903) );
  NAND2_X1 U7377 ( .A1(n8931), .A2(n8903), .ZN(n5902) );
  NAND2_X1 U7378 ( .A1(n5904), .A2(n5902), .ZN(n8921) );
  AND2_X1 U7379 ( .A1(n5888), .A2(n8880), .ZN(n5910) );
  NAND2_X1 U7380 ( .A1(n9036), .A2(n8516), .ZN(n5914) );
  NAND2_X1 U7381 ( .A1(n9042), .A2(n8868), .ZN(n8841) );
  AND2_X1 U7382 ( .A1(n5914), .A2(n8841), .ZN(n5913) );
  INV_X1 U7383 ( .A(n5713), .ZN(n5926) );
  INV_X1 U7384 ( .A(n5956), .ZN(n5929) );
  XNOR2_X1 U7385 ( .A(n5794), .B(n5929), .ZN(n9021) );
  INV_X1 U7386 ( .A(n9021), .ZN(n5716) );
  NAND2_X1 U7387 ( .A1(n5714), .A2(n6973), .ZN(n5715) );
  NAND3_X1 U7388 ( .A1(n5982), .A2(n10052), .A3(n5715), .ZN(n10051) );
  NAND2_X1 U7389 ( .A1(n10096), .A2(n10075), .ZN(n9009) );
  NAND2_X1 U7390 ( .A1(n5716), .A2(n8984), .ZN(n5717) );
  NAND2_X1 U7391 ( .A1(n5718), .A2(n5717), .ZN(P2_U3486) );
  NAND2_X1 U7392 ( .A1(n5720), .A2(n5719), .ZN(n5722) );
  NAND2_X1 U7393 ( .A1(n5722), .A2(n5721), .ZN(n5786) );
  INV_X1 U7394 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5723) );
  MUX2_X1 U7395 ( .A(n5723), .B(n9787), .S(n6661), .Z(n5725) );
  XNOR2_X1 U7396 ( .A(n5725), .B(SI_28_), .ZN(n5785) );
  NAND2_X1 U7397 ( .A1(n5786), .A2(n5785), .ZN(n5727) );
  INV_X1 U7398 ( .A(SI_28_), .ZN(n5724) );
  NAND2_X1 U7399 ( .A1(n5725), .A2(n5724), .ZN(n5726) );
  INV_X1 U7400 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n5728) );
  INV_X1 U7401 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9784) );
  MUX2_X1 U7402 ( .A(n5728), .B(n9784), .S(n6661), .Z(n5729) );
  NAND2_X1 U7403 ( .A1(n5730), .A2(n5729), .ZN(n5731) );
  INV_X1 U7404 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n5732) );
  INV_X1 U7405 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8499) );
  MUX2_X1 U7406 ( .A(n5732), .B(n8499), .S(n6661), .Z(n5734) );
  INV_X1 U7407 ( .A(SI_30_), .ZN(n5733) );
  NAND2_X1 U7408 ( .A1(n5734), .A2(n5733), .ZN(n5737) );
  INV_X1 U7409 ( .A(n5734), .ZN(n5735) );
  NAND2_X1 U7410 ( .A1(n5735), .A2(SI_30_), .ZN(n5736) );
  NAND2_X1 U7411 ( .A1(n5750), .A2(n5749), .ZN(n5738) );
  INV_X1 U7412 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5739) );
  INV_X1 U7413 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n8292) );
  MUX2_X1 U7414 ( .A(n5739), .B(n8292), .S(n6661), .Z(n5740) );
  XNOR2_X1 U7415 ( .A(n5740), .B(SI_31_), .ZN(n5741) );
  NAND2_X1 U7416 ( .A1(n9085), .A2(n5787), .ZN(n5744) );
  NAND2_X1 U7417 ( .A1(n5788), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n5743) );
  OR2_X1 U7418 ( .A1(n5298), .A2(n8781), .ZN(n5767) );
  NAND2_X1 U7419 ( .A1(n5745), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5748) );
  INV_X1 U7420 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9013) );
  OR2_X1 U7421 ( .A1(n5760), .A2(n9013), .ZN(n5747) );
  INV_X1 U7422 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8783) );
  OR2_X1 U7423 ( .A1(n5763), .A2(n8783), .ZN(n5746) );
  NAND4_X1 U7424 ( .A1(n5767), .A2(n5748), .A3(n5747), .A4(n5746), .ZN(n8780)
         );
  INV_X1 U7425 ( .A(n8780), .ZN(n5768) );
  NAND2_X1 U7426 ( .A1(n8498), .A2(n5787), .ZN(n5752) );
  NAND2_X1 U7427 ( .A1(n5788), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n5751) );
  NAND2_X1 U7428 ( .A1(n5745), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U7429 ( .A1(n5753), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5755) );
  INV_X1 U7430 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8787) );
  OR2_X1 U7431 ( .A1(n5763), .A2(n8787), .ZN(n5754) );
  NAND4_X1 U7432 ( .A1(n5767), .A2(n5756), .A3(n5755), .A4(n5754), .ZN(n8618)
         );
  INV_X1 U7433 ( .A(n8618), .ZN(n5757) );
  NAND2_X1 U7434 ( .A1(n8784), .A2(n5757), .ZN(n5946) );
  NAND2_X1 U7435 ( .A1(n5788), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5759) );
  INV_X1 U7436 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5989) );
  OR2_X1 U7437 ( .A1(n5760), .A2(n5989), .ZN(n5766) );
  INV_X1 U7438 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5974) );
  OR2_X1 U7439 ( .A1(n5761), .A2(n5974), .ZN(n5765) );
  INV_X1 U7440 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n5762) );
  OR2_X1 U7441 ( .A1(n5763), .A2(n5762), .ZN(n5764) );
  NAND2_X1 U7442 ( .A1(n5973), .A2(n8619), .ZN(n5932) );
  AND2_X1 U7443 ( .A1(n4368), .A2(n4399), .ZN(n5798) );
  INV_X1 U7444 ( .A(n5798), .ZN(n5793) );
  AND2_X1 U7445 ( .A1(n9010), .A2(n5768), .ZN(n5949) );
  INV_X1 U7446 ( .A(n8784), .ZN(n9016) );
  NAND2_X1 U7447 ( .A1(n9016), .A2(n8618), .ZN(n5947) );
  NAND2_X1 U7448 ( .A1(n5947), .A2(n5933), .ZN(n5941) );
  OR2_X2 U7449 ( .A1(n4383), .A2(n5928), .ZN(n8821) );
  NAND2_X1 U7450 ( .A1(n5917), .A2(n5914), .ZN(n8843) );
  INV_X1 U7451 ( .A(n8843), .ZN(n8845) );
  NAND2_X1 U7452 ( .A1(n5916), .A2(n8841), .ZN(n8857) );
  OR2_X1 U7453 ( .A1(n5867), .A2(n5048), .ZN(n8009) );
  INV_X1 U7454 ( .A(n7071), .ZN(n5772) );
  AND2_X1 U7455 ( .A1(n5820), .A2(n5826), .ZN(n7185) );
  INV_X1 U7456 ( .A(n7185), .ZN(n5771) );
  NOR4_X1 U7457 ( .A1(n5772), .A2(n5771), .A3(n5811), .A4(n5770), .ZN(n5775)
         );
  AND2_X1 U7458 ( .A1(n5802), .A2(n5829), .ZN(n7357) );
  INV_X1 U7459 ( .A(n7016), .ZN(n5804) );
  INV_X1 U7460 ( .A(n7065), .ZN(n6974) );
  AND2_X1 U7461 ( .A1(n5697), .A2(n6974), .ZN(n5803) );
  NOR2_X1 U7462 ( .A1(n5804), .A2(n5803), .ZN(n7054) );
  NAND2_X1 U7463 ( .A1(n5774), .A2(n5773), .ZN(n7393) );
  NAND4_X1 U7464 ( .A1(n5775), .A2(n7357), .A3(n7054), .A4(n7393), .ZN(n5776)
         );
  NAND2_X1 U7465 ( .A1(n5839), .A2(n5843), .ZN(n7497) );
  NOR4_X1 U7466 ( .A1(n5838), .A2(n5776), .A3(n7371), .A4(n7497), .ZN(n5777)
         );
  NAND4_X1 U7467 ( .A1(n8009), .A2(n5778), .A3(n7726), .A4(n5777), .ZN(n5780)
         );
  OR2_X1 U7468 ( .A1(n5779), .A2(n4374), .ZN(n5877) );
  NAND2_X1 U7469 ( .A1(n5876), .A2(n5871), .ZN(n7995) );
  OR4_X1 U7470 ( .A1(n5780), .A2(n8036), .A3(n7897), .A4(n7995), .ZN(n5781) );
  NOR4_X1 U7471 ( .A1(n8921), .A2(n5880), .A3(n8946), .A4(n5781), .ZN(n5782)
         );
  NAND3_X1 U7472 ( .A1(n8889), .A2(n8909), .A3(n5782), .ZN(n5783) );
  NOR3_X1 U7473 ( .A1(n8857), .A2(n8882), .A3(n5783), .ZN(n5784) );
  NAND4_X1 U7474 ( .A1(n8831), .A2(n8870), .A3(n8845), .A4(n5784), .ZN(n5791)
         );
  NAND2_X1 U7475 ( .A1(n9096), .A2(n5787), .ZN(n5790) );
  NAND2_X1 U7476 ( .A1(n5788), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5789) );
  NOR4_X1 U7477 ( .A1(n5793), .A2(n5949), .A3(n5941), .A4(n5792), .ZN(n5799)
         );
  NAND2_X1 U7478 ( .A1(n5795), .A2(n5935), .ZN(n8807) );
  NAND2_X1 U7479 ( .A1(n8965), .A2(n8505), .ZN(n5796) );
  INV_X1 U7480 ( .A(n9010), .ZN(n8961) );
  NAND2_X1 U7481 ( .A1(n5947), .A2(n8780), .ZN(n5797) );
  XNOR2_X1 U7482 ( .A(n5800), .B(n8767), .ZN(n5951) );
  MUX2_X1 U7483 ( .A(n8505), .B(n5958), .S(n5986), .Z(n5945) );
  INV_X1 U7484 ( .A(n5801), .ZN(n5875) );
  INV_X1 U7485 ( .A(n5802), .ZN(n5823) );
  NOR2_X1 U7486 ( .A1(n5770), .A2(n5803), .ZN(n5813) );
  NOR2_X1 U7487 ( .A1(n5803), .A2(n7813), .ZN(n5805) );
  MUX2_X1 U7488 ( .A(n5805), .B(n5804), .S(n5980), .Z(n5808) );
  INV_X1 U7489 ( .A(n5808), .ZN(n5812) );
  INV_X1 U7490 ( .A(n5806), .ZN(n5810) );
  AOI21_X1 U7491 ( .B1(n5808), .B2(n5807), .A(n5810), .ZN(n5809) );
  NAND2_X1 U7492 ( .A1(n5819), .A2(n5814), .ZN(n5817) );
  NAND2_X1 U7493 ( .A1(n5824), .A2(n5815), .ZN(n5816) );
  MUX2_X1 U7494 ( .A(n5817), .B(n5816), .S(n5986), .Z(n5818) );
  INV_X1 U7495 ( .A(n5819), .ZN(n5821) );
  OAI211_X1 U7496 ( .C1(n5823), .C2(n5825), .A(n5822), .B(n5829), .ZN(n5834)
         );
  INV_X1 U7497 ( .A(n5824), .ZN(n5827) );
  OAI211_X1 U7498 ( .C1(n5828), .C2(n5827), .A(n5826), .B(n5825), .ZN(n5832)
         );
  INV_X1 U7499 ( .A(n5829), .ZN(n5830) );
  AOI21_X1 U7500 ( .B1(n5832), .B2(n5831), .A(n5830), .ZN(n5833) );
  MUX2_X1 U7501 ( .A(n5834), .B(n5833), .S(n6656), .Z(n5835) );
  NAND2_X1 U7502 ( .A1(n5835), .A2(n7367), .ZN(n5836) );
  OAI21_X1 U7503 ( .B1(n6656), .B2(n5837), .A(n5836), .ZN(n5851) );
  INV_X1 U7504 ( .A(n5838), .ZN(n7617) );
  NAND2_X1 U7505 ( .A1(n7617), .A2(n5840), .ZN(n5846) );
  INV_X1 U7506 ( .A(n5846), .ZN(n5850) );
  INV_X1 U7507 ( .A(n5841), .ZN(n5848) );
  AND2_X1 U7508 ( .A1(n5843), .A2(n5842), .ZN(n5845) );
  OAI211_X1 U7509 ( .C1(n5846), .C2(n5845), .A(n5853), .B(n5844), .ZN(n5847)
         );
  AOI21_X1 U7510 ( .B1(n5851), .B2(n5850), .A(n5849), .ZN(n5861) );
  NAND2_X1 U7511 ( .A1(n5857), .A2(n5852), .ZN(n5855) );
  NAND2_X1 U7512 ( .A1(n5856), .A2(n5853), .ZN(n5854) );
  MUX2_X1 U7513 ( .A(n5855), .B(n5854), .S(n5986), .Z(n5860) );
  MUX2_X1 U7514 ( .A(n5857), .B(n5856), .S(n6656), .Z(n5859) );
  INV_X1 U7515 ( .A(n7897), .ZN(n5858) );
  OAI211_X1 U7516 ( .C1(n5861), .C2(n5860), .A(n5859), .B(n5858), .ZN(n5865)
         );
  NAND2_X1 U7517 ( .A1(n10079), .A2(n7877), .ZN(n5863) );
  MUX2_X1 U7518 ( .A(n5863), .B(n5862), .S(n6656), .Z(n5864) );
  AND2_X1 U7519 ( .A1(n5865), .A2(n5864), .ZN(n5868) );
  INV_X1 U7520 ( .A(n5868), .ZN(n5870) );
  MUX2_X1 U7521 ( .A(n8016), .B(n8624), .S(n5986), .Z(n5866) );
  AOI21_X1 U7522 ( .B1(n5048), .B2(n5870), .A(n5869), .ZN(n5872) );
  OAI211_X1 U7523 ( .C1(n5879), .C2(n8036), .A(n5873), .B(n5882), .ZN(n5874)
         );
  NAND2_X1 U7524 ( .A1(n5877), .A2(n5876), .ZN(n5878) );
  OAI21_X1 U7525 ( .B1(n5879), .B2(n5878), .A(n5884), .ZN(n5881) );
  INV_X1 U7526 ( .A(n5880), .ZN(n8936) );
  INV_X1 U7527 ( .A(n5882), .ZN(n5883) );
  NAND3_X1 U7528 ( .A1(n5906), .A2(n5902), .A3(n5907), .ZN(n5900) );
  INV_X1 U7529 ( .A(n5894), .ZN(n5887) );
  NAND4_X1 U7530 ( .A1(n5893), .A2(n5986), .A3(n5903), .A4(n5890), .ZN(n5886)
         );
  NOR2_X1 U7531 ( .A1(n5887), .A2(n5886), .ZN(n5899) );
  INV_X1 U7532 ( .A(n5888), .ZN(n5889) );
  AOI211_X1 U7533 ( .C1(n5893), .C2(n5890), .A(n5986), .B(n5889), .ZN(n5892)
         );
  INV_X1 U7534 ( .A(n8841), .ZN(n5891) );
  INV_X1 U7535 ( .A(n5910), .ZN(n5895) );
  NAND4_X1 U7536 ( .A1(n5895), .A2(n5986), .A3(n5894), .A4(n5893), .ZN(n5896)
         );
  AOI211_X1 U7537 ( .C1(n5900), .C2(n5899), .A(n8843), .B(n5898), .ZN(n5923)
         );
  NAND2_X1 U7538 ( .A1(n5902), .A2(n5901), .ZN(n5905) );
  OAI211_X1 U7539 ( .C1(n5906), .C2(n5905), .A(n5904), .B(n5903), .ZN(n5911)
         );
  INV_X1 U7540 ( .A(n5907), .ZN(n5908) );
  NOR2_X1 U7541 ( .A1(n5908), .A2(n5986), .ZN(n5909) );
  NAND4_X1 U7542 ( .A1(n5911), .A2(n8870), .A3(n5910), .A4(n5909), .ZN(n5922)
         );
  INV_X1 U7543 ( .A(n5917), .ZN(n5912) );
  NOR2_X1 U7544 ( .A1(n5913), .A2(n5912), .ZN(n5919) );
  INV_X1 U7545 ( .A(n5914), .ZN(n5915) );
  AOI21_X1 U7546 ( .B1(n5917), .B2(n5916), .A(n5915), .ZN(n5918) );
  MUX2_X1 U7547 ( .A(n5919), .B(n5918), .S(n5986), .Z(n5921) );
  INV_X1 U7548 ( .A(n8831), .ZN(n5920) );
  INV_X1 U7549 ( .A(n5924), .ZN(n5925) );
  MUX2_X1 U7550 ( .A(n5926), .B(n5925), .S(n5986), .Z(n5927) );
  MUX2_X1 U7551 ( .A(n4383), .B(n5928), .S(n6656), .Z(n5930) );
  OAI21_X1 U7552 ( .B1(n5931), .B2(n5930), .A(n5929), .ZN(n5938) );
  INV_X1 U7553 ( .A(n5964), .ZN(n5937) );
  MUX2_X1 U7554 ( .A(n5935), .B(n5934), .S(n6656), .Z(n5936) );
  NAND3_X1 U7555 ( .A1(n5938), .A2(n5937), .A3(n5936), .ZN(n5944) );
  NAND2_X1 U7556 ( .A1(n5944), .A2(n5940), .ZN(n5942) );
  AOI21_X1 U7557 ( .B1(n5942), .B2(n5958), .A(n5941), .ZN(n5943) );
  INV_X1 U7558 ( .A(n5946), .ZN(n5948) );
  OAI21_X1 U7559 ( .B1(n5948), .B2(n5986), .A(n5947), .ZN(n5950) );
  OR2_X1 U7560 ( .A1(n6922), .A2(P2_U3151), .ZN(n7902) );
  INV_X1 U7561 ( .A(n5953), .ZN(n6976) );
  INV_X1 U7562 ( .A(n5982), .ZN(n7053) );
  AND2_X1 U7563 ( .A1(n6918), .A2(n7053), .ZN(n6929) );
  NAND3_X1 U7564 ( .A1(n6976), .A2(n6929), .A3(n8643), .ZN(n5954) );
  OAI211_X1 U7565 ( .C1(n7813), .C2(n7902), .A(n5954), .B(P2_B_REG_SCAN_IN), 
        .ZN(n5955) );
  XNOR2_X1 U7566 ( .A(n5964), .B(n5962), .ZN(n5963) );
  NAND2_X1 U7567 ( .A1(n5963), .A2(n8952), .ZN(n5970) );
  XNOR2_X1 U7568 ( .A(n5965), .B(n5964), .ZN(n8795) );
  NAND2_X1 U7569 ( .A1(n5263), .A2(P2_B_REG_SCAN_IN), .ZN(n5966) );
  AND2_X1 U7570 ( .A1(n8949), .A2(n5966), .ZN(n8779) );
  AOI22_X1 U7571 ( .A1(n8779), .A2(n8618), .B1(n5959), .B2(n5656), .ZN(n5967)
         );
  OR2_X1 U7572 ( .A1(n10096), .A2(n5974), .ZN(n5975) );
  OAI21_X1 U7573 ( .B1(n5993), .B2(n10094), .A(n5977), .ZN(P2_U3488) );
  INV_X1 U7574 ( .A(n5984), .ZN(n5978) );
  NOR2_X1 U7575 ( .A1(n5979), .A2(n5978), .ZN(n6921) );
  NAND2_X1 U7576 ( .A1(n6921), .A2(n6918), .ZN(n6915) );
  NAND2_X1 U7577 ( .A1(n5980), .A2(n7563), .ZN(n6971) );
  OR2_X1 U7578 ( .A1(n5981), .A2(n6971), .ZN(n6927) );
  AND2_X1 U7579 ( .A1(n6927), .A2(n5982), .ZN(n5983) );
  OR2_X1 U7580 ( .A1(n6915), .A2(n5983), .ZN(n5988) );
  NAND2_X1 U7581 ( .A1(n6972), .A2(n5984), .ZN(n5985) );
  NAND2_X1 U7582 ( .A1(n6931), .A2(n6918), .ZN(n6910) );
  NAND3_X1 U7583 ( .A1(n5986), .A2(n6927), .A3(n10052), .ZN(n6909) );
  AND2_X1 U7584 ( .A1(n6909), .A2(n10023), .ZN(n6920) );
  OR2_X1 U7585 ( .A1(n6910), .A2(n6920), .ZN(n5987) );
  INV_X1 U7586 ( .A(n5991), .ZN(n5992) );
  OAI21_X1 U7587 ( .B1(n5993), .B2(n10082), .A(n5992), .ZN(P2_U3456) );
  NOR2_X2 U7588 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6121) );
  NAND3_X1 U7589 ( .A1(n6079), .A2(n6121), .A3(n5994), .ZN(n6157) );
  NOR2_X1 U7590 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5999) );
  NOR2_X1 U7591 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5998) );
  NOR2_X1 U7592 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5997) );
  NOR2_X1 U7593 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5996) );
  NOR2_X1 U7594 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n6003) );
  NOR2_X1 U7595 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n6002) );
  NAND2_X1 U7596 ( .A1(n6010), .A2(n6244), .ZN(n6009) );
  NAND2_X1 U7597 ( .A1(n6114), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U7598 ( .A1(n6088), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6015) );
  INV_X1 U7599 ( .A(n6011), .ZN(n9785) );
  NAND2_X1 U7600 ( .A1(n6074), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6014) );
  NAND4_X1 U7601 ( .A1(n6016), .A2(n6015), .A3(n6014), .A4(n6013), .ZN(n6901)
         );
  INV_X1 U7602 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7603 ( .A1(n6018), .A2(n6044), .ZN(n6019) );
  INV_X1 U7604 ( .A(n6027), .ZN(n6021) );
  INV_X1 U7605 ( .A(n6023), .ZN(n6024) );
  NAND2_X1 U7606 ( .A1(n6024), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6025) );
  MUX2_X1 U7607 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6025), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n6026) );
  INV_X1 U7608 ( .A(n8372), .ZN(n6899) );
  NAND2_X1 U7609 ( .A1(n6031), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6032) );
  NAND2_X1 U7610 ( .A1(n4406), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6034) );
  INV_X1 U7611 ( .A(n8032), .ZN(n6035) );
  NAND2_X2 U7612 ( .A1(n6592), .A2(n6036), .ZN(n6653) );
  NAND2_X1 U7613 ( .A1(n6901), .A2(n6305), .ZN(n6054) );
  INV_X1 U7614 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6042) );
  NAND2_X1 U7615 ( .A1(n6377), .A2(n6042), .ZN(n6043) );
  NAND2_X1 U7616 ( .A1(n6408), .A2(n6407), .ZN(n6410) );
  OR2_X1 U7617 ( .A1(n7162), .A2(n8338), .ZN(n7529) );
  NAND2_X1 U7618 ( .A1(n8437), .A2(n8193), .ZN(n6048) );
  NAND3_X2 U7619 ( .A1(n7529), .A2(n6653), .A3(n6048), .ZN(n6570) );
  NAND2_X1 U7620 ( .A1(n6661), .A2(SI_0_), .ZN(n6049) );
  XNOR2_X1 U7621 ( .A(n6049), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9792) );
  MUX2_X1 U7622 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9792), .S(n6062), .Z(n8387) );
  INV_X1 U7623 ( .A(n6653), .ZN(n6631) );
  AOI22_X1 U7624 ( .A1(n6131), .A2(n8387), .B1(n6631), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7625 ( .A1(n6054), .A2(n6053), .ZN(n6865) );
  NAND2_X1 U7626 ( .A1(n6901), .A2(n6584), .ZN(n6056) );
  AOI22_X1 U7627 ( .A1(n8387), .A2(n6305), .B1(n6631), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U7628 ( .A1(n6056), .A2(n6055), .ZN(n6866) );
  NAND2_X1 U7629 ( .A1(n6865), .A2(n6866), .ZN(n6864) );
  OR2_X1 U7630 ( .A1(n6546), .A2(n8387), .ZN(n6057) );
  NAND2_X1 U7631 ( .A1(n6088), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7632 ( .A1(n6074), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7633 ( .A1(n6089), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U7634 ( .A1(n7140), .A2(n6305), .ZN(n6067) );
  INV_X1 U7635 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6659) );
  INV_X1 U7636 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7637 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6063) );
  OR2_X1 U7638 ( .A1(n6062), .A2(n9299), .ZN(n6065) );
  NAND2_X1 U7639 ( .A1(n4511), .A2(n6131), .ZN(n6066) );
  NAND2_X1 U7640 ( .A1(n6067), .A2(n6066), .ZN(n6068) );
  NOR2_X1 U7641 ( .A1(n7636), .A2(n6103), .ZN(n6069) );
  AOI21_X1 U7642 ( .B1(n7140), .B2(n6584), .A(n6069), .ZN(n6071) );
  XNOR2_X1 U7643 ( .A(n6070), .B(n6071), .ZN(n9146) );
  NAND2_X1 U7644 ( .A1(n9145), .A2(n9146), .ZN(n9144) );
  INV_X1 U7645 ( .A(n6070), .ZN(n6072) );
  NAND2_X1 U7646 ( .A1(n6072), .A2(n6071), .ZN(n6073) );
  NAND2_X1 U7647 ( .A1(n6114), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6078) );
  NAND2_X1 U7648 ( .A1(n6088), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U7649 ( .A1(n6074), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7650 ( .A1(n6089), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7651 ( .A1(n9293), .A2(n6305), .ZN(n6085) );
  OR2_X1 U7652 ( .A1(n6271), .A2(n6670), .ZN(n6083) );
  INV_X1 U7653 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6660) );
  OR2_X1 U7654 ( .A1(n8293), .A2(n6660), .ZN(n6082) );
  INV_X1 U7655 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7656 ( .A1(n6123), .A2(n6080), .ZN(n6094) );
  OAI21_X1 U7657 ( .B1(n6123), .B2(n6080), .A(n6094), .ZN(n6876) );
  OR2_X1 U7658 ( .A1(n6062), .A2(n6876), .ZN(n6081) );
  AND3_X2 U7659 ( .A1(n6083), .A2(n6082), .A3(n6081), .ZN(n7247) );
  INV_X1 U7660 ( .A(n7247), .ZN(n7485) );
  NAND2_X1 U7661 ( .A1(n7485), .A2(n6131), .ZN(n6084) );
  NAND2_X1 U7662 ( .A1(n6085), .A2(n6084), .ZN(n6086) );
  XNOR2_X1 U7663 ( .A(n6086), .B(n6546), .ZN(n6106) );
  NOR2_X1 U7664 ( .A1(n7247), .A2(n6286), .ZN(n6087) );
  AOI21_X1 U7665 ( .B1(n9293), .B2(n6584), .A(n6087), .ZN(n6107) );
  XNOR2_X1 U7666 ( .A(n6106), .B(n6107), .ZN(n7047) );
  NAND2_X1 U7667 ( .A1(n6088), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6093) );
  NAND2_X1 U7668 ( .A1(n6089), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6092) );
  INV_X1 U7669 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9860) );
  NAND2_X1 U7670 ( .A1(n6114), .A2(n9860), .ZN(n6091) );
  NAND2_X1 U7671 ( .A1(n6074), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U7672 ( .A1(n9292), .A2(n6305), .ZN(n6101) );
  OR2_X1 U7673 ( .A1(n6271), .A2(n6668), .ZN(n6099) );
  INV_X1 U7674 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6664) );
  OR2_X1 U7675 ( .A1(n8293), .A2(n6664), .ZN(n6098) );
  NAND2_X1 U7676 ( .A1(n6094), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6096) );
  INV_X1 U7677 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n6095) );
  XNOR2_X1 U7678 ( .A(n6096), .B(n6095), .ZN(n6776) );
  OR2_X1 U7679 ( .A1(n6062), .A2(n6776), .ZN(n6097) );
  INV_X1 U7680 ( .A(n9864), .ZN(n7242) );
  NAND2_X1 U7681 ( .A1(n7242), .A2(n6131), .ZN(n6100) );
  NAND2_X1 U7682 ( .A1(n6101), .A2(n6100), .ZN(n6102) );
  XNOR2_X1 U7683 ( .A(n6102), .B(n6546), .ZN(n6110) );
  INV_X1 U7684 ( .A(n6110), .ZN(n6105) );
  NOR2_X1 U7685 ( .A1(n9864), .A2(n6103), .ZN(n6104) );
  AOI21_X1 U7686 ( .B1(n9292), .B2(n6584), .A(n6104), .ZN(n6109) );
  NAND2_X1 U7687 ( .A1(n6105), .A2(n6109), .ZN(n6111) );
  INV_X1 U7688 ( .A(n6106), .ZN(n6108) );
  NAND2_X1 U7689 ( .A1(n6108), .A2(n6107), .ZN(n7128) );
  AND2_X1 U7690 ( .A1(n6111), .A2(n7128), .ZN(n6113) );
  XNOR2_X1 U7691 ( .A(n6110), .B(n6109), .ZN(n7131) );
  INV_X1 U7692 ( .A(n6111), .ZN(n6112) );
  NAND2_X1 U7693 ( .A1(n6089), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7694 ( .A1(n4335), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6119) );
  NOR2_X1 U7695 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6115) );
  NOR2_X1 U7696 ( .A1(n6141), .A2(n6115), .ZN(n7606) );
  NAND2_X1 U7697 ( .A1(n6114), .A2(n7606), .ZN(n6118) );
  INV_X1 U7698 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6116) );
  NAND4_X1 U7699 ( .A1(n6120), .A2(n6119), .A3(n6118), .A4(n6117), .ZN(n9291)
         );
  NAND2_X1 U7700 ( .A1(n9291), .A2(n6305), .ZN(n6133) );
  OR2_X1 U7701 ( .A1(n6667), .A2(n6271), .ZN(n6130) );
  INV_X1 U7702 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6665) );
  OR2_X1 U7703 ( .A1(n8293), .A2(n6665), .ZN(n6129) );
  INV_X1 U7704 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6244) );
  OR2_X1 U7705 ( .A1(n6121), .A2(n6244), .ZN(n6122) );
  AND2_X1 U7706 ( .A1(n6123), .A2(n6122), .ZN(n6125) );
  INV_X1 U7707 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U7708 ( .A1(n6125), .A2(n6124), .ZN(n6147) );
  INV_X1 U7709 ( .A(n6125), .ZN(n6126) );
  NAND2_X1 U7710 ( .A1(n6126), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U7711 ( .A1(n6147), .A2(n6127), .ZN(n6937) );
  OR2_X1 U7712 ( .A1(n6062), .A2(n6937), .ZN(n6128) );
  INV_X1 U7713 ( .A(n6131), .ZN(n6249) );
  NAND2_X1 U7714 ( .A1(n7607), .A2(n6131), .ZN(n6132) );
  NAND2_X1 U7715 ( .A1(n6133), .A2(n6132), .ZN(n6134) );
  XNOR2_X1 U7716 ( .A(n6134), .B(n6587), .ZN(n6136) );
  NOR2_X1 U7717 ( .A1(n7290), .A2(n6286), .ZN(n6135) );
  AOI21_X1 U7718 ( .B1(n9291), .B2(n6584), .A(n6135), .ZN(n6137) );
  XNOR2_X1 U7719 ( .A(n6136), .B(n6137), .ZN(n7294) );
  INV_X1 U7720 ( .A(n6136), .ZN(n6139) );
  INV_X1 U7721 ( .A(n6137), .ZN(n6138) );
  NAND2_X1 U7722 ( .A1(n6139), .A2(n6138), .ZN(n6140) );
  NAND2_X1 U7723 ( .A1(n8177), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7724 ( .A1(n4335), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6145) );
  NOR2_X1 U7725 ( .A1(n6141), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6142) );
  NOR2_X1 U7726 ( .A1(n6161), .A2(n6142), .ZN(n7627) );
  NAND2_X1 U7727 ( .A1(n4333), .A2(n7627), .ZN(n6144) );
  NAND2_X1 U7728 ( .A1(n6074), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6143) );
  OR2_X1 U7729 ( .A1(n6672), .A2(n6271), .ZN(n6150) );
  NAND2_X1 U7730 ( .A1(n6147), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6148) );
  XNOR2_X1 U7731 ( .A(n6148), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6795) );
  AOI22_X1 U7732 ( .A1(n6412), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6411), .B2(
        n6795), .ZN(n6149) );
  NAND2_X1 U7733 ( .A1(n6150), .A2(n6149), .ZN(n7214) );
  OAI22_X1 U7734 ( .A1(n7506), .A2(n6286), .B1(n7629), .B2(n6249), .ZN(n6151)
         );
  XNOR2_X1 U7735 ( .A(n6151), .B(n6546), .ZN(n6154) );
  NAND2_X1 U7736 ( .A1(n6155), .A2(n6154), .ZN(n7298) );
  OR2_X1 U7737 ( .A1(n7506), .A2(n6570), .ZN(n6153) );
  NAND2_X1 U7738 ( .A1(n7214), .A2(n6305), .ZN(n6152) );
  AND2_X1 U7739 ( .A1(n6153), .A2(n6152), .ZN(n7299) );
  NAND2_X1 U7740 ( .A1(n7298), .A2(n7299), .ZN(n6156) );
  OR2_X1 U7741 ( .A1(n6676), .A2(n6271), .ZN(n6160) );
  NAND2_X1 U7742 ( .A1(n6157), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6158) );
  XNOR2_X1 U7743 ( .A(n6158), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6828) );
  AOI22_X1 U7744 ( .A1(n6412), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6411), .B2(
        n6828), .ZN(n6159) );
  NAND2_X1 U7745 ( .A1(n4335), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6165) );
  INV_X2 U7746 ( .A(n6423), .ZN(n8176) );
  NAND2_X1 U7747 ( .A1(n8176), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6164) );
  NAND2_X1 U7748 ( .A1(n6161), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6178) );
  OAI21_X1 U7749 ( .B1(n6161), .B2(P1_REG3_REG_6__SCAN_IN), .A(n6178), .ZN(
        n7387) );
  INV_X1 U7750 ( .A(n7387), .ZN(n7511) );
  NAND2_X1 U7751 ( .A1(n4332), .A2(n7511), .ZN(n6163) );
  INV_X2 U7752 ( .A(n6542), .ZN(n8177) );
  NAND2_X1 U7753 ( .A1(n8177), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6162) );
  NAND4_X1 U7754 ( .A1(n6165), .A2(n6164), .A3(n6163), .A4(n6162), .ZN(n9289)
         );
  NAND2_X1 U7755 ( .A1(n9289), .A2(n6305), .ZN(n6166) );
  OAI21_X1 U7756 ( .B1(n9875), .B2(n6249), .A(n6166), .ZN(n6167) );
  XNOR2_X1 U7757 ( .A(n6167), .B(n6587), .ZN(n7383) );
  OR2_X1 U7758 ( .A1(n9875), .A2(n6103), .ZN(n6169) );
  NAND2_X1 U7759 ( .A1(n9289), .A2(n6584), .ZN(n6168) );
  NAND2_X1 U7760 ( .A1(n6169), .A2(n6168), .ZN(n7382) );
  INV_X1 U7761 ( .A(n7382), .ZN(n6170) );
  AND2_X1 U7762 ( .A1(n7383), .A2(n6170), .ZN(n6173) );
  INV_X1 U7763 ( .A(n7383), .ZN(n6171) );
  NAND2_X1 U7764 ( .A1(n6171), .A2(n7382), .ZN(n6172) );
  OR2_X1 U7765 ( .A1(n6683), .A2(n6271), .ZN(n6177) );
  NAND2_X1 U7766 ( .A1(n6174), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6175) );
  XNOR2_X1 U7767 ( .A(n6175), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6851) );
  AOI22_X1 U7768 ( .A1(n6412), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6411), .B2(
        n6851), .ZN(n6176) );
  NAND2_X1 U7769 ( .A1(n6177), .A2(n6176), .ZN(n7553) );
  NAND2_X1 U7770 ( .A1(n7553), .A2(n6131), .ZN(n6185) );
  NAND2_X1 U7771 ( .A1(n8177), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7772 ( .A1(n4335), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6182) );
  AND2_X1 U7773 ( .A1(n6178), .A2(n6857), .ZN(n6179) );
  NOR2_X1 U7774 ( .A1(n6193), .A2(n6179), .ZN(n7644) );
  NAND2_X1 U7775 ( .A1(n4332), .A2(n7644), .ZN(n6181) );
  NAND2_X1 U7776 ( .A1(n8176), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6180) );
  OR2_X1 U7777 ( .A1(n7703), .A2(n6286), .ZN(n6184) );
  NAND2_X1 U7778 ( .A1(n6185), .A2(n6184), .ZN(n6186) );
  XNOR2_X1 U7779 ( .A(n6186), .B(n6587), .ZN(n6187) );
  AOI22_X1 U7780 ( .A1(n7553), .A2(n6305), .B1(n7518), .B2(n6584), .ZN(n6188)
         );
  NAND2_X1 U7781 ( .A1(n6187), .A2(n6188), .ZN(n7439) );
  INV_X1 U7782 ( .A(n6187), .ZN(n6190) );
  INV_X1 U7783 ( .A(n6188), .ZN(n6189) );
  NAND2_X1 U7784 ( .A1(n6190), .A2(n6189), .ZN(n7440) );
  NAND2_X1 U7785 ( .A1(n6685), .A2(n8291), .ZN(n6192) );
  NOR2_X1 U7786 ( .A1(n6174), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n6228) );
  OR2_X1 U7787 ( .A1(n6228), .A2(n6244), .ZN(n6208) );
  XNOR2_X1 U7788 ( .A(n6208), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6960) );
  AOI22_X1 U7789 ( .A1(n6412), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6411), .B2(
        n6960), .ZN(n6191) );
  NAND2_X1 U7790 ( .A1(n7697), .A2(n6131), .ZN(n6200) );
  NAND2_X1 U7791 ( .A1(n4335), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7792 ( .A1(n8176), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6197) );
  NOR2_X1 U7793 ( .A1(n6193), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7794 ( .A1(n4332), .A2(n5085), .ZN(n6196) );
  NAND2_X1 U7795 ( .A1(n8177), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6195) );
  OR2_X1 U7796 ( .A1(n7760), .A2(n6286), .ZN(n6199) );
  NAND2_X1 U7797 ( .A1(n6200), .A2(n6199), .ZN(n6201) );
  XNOR2_X1 U7798 ( .A(n6201), .B(n6587), .ZN(n6204) );
  NOR2_X1 U7799 ( .A1(n7760), .A2(n6570), .ZN(n6202) );
  AOI21_X1 U7800 ( .B1(n7697), .B2(n6305), .A(n6202), .ZN(n7699) );
  INV_X1 U7801 ( .A(n6203), .ZN(n6205) );
  NAND2_X1 U7802 ( .A1(n6205), .A2(n6204), .ZN(n6206) );
  NAND2_X1 U7803 ( .A1(n6709), .A2(n8291), .ZN(n6212) );
  INV_X1 U7804 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U7805 ( .A1(n6208), .A2(n6207), .ZN(n6209) );
  NAND2_X1 U7806 ( .A1(n6209), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6210) );
  XNOR2_X1 U7807 ( .A(n6210), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7087) );
  AOI22_X1 U7808 ( .A1(n6412), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6411), .B2(
        n7087), .ZN(n6211) );
  NAND2_X1 U7809 ( .A1(n7763), .A2(n6131), .ZN(n6220) );
  NAND2_X1 U7810 ( .A1(n4335), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U7811 ( .A1(n8177), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6217) );
  NOR2_X1 U7812 ( .A1(n6213), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6214) );
  OR2_X1 U7813 ( .A1(n6250), .A2(n6214), .ZN(n7757) );
  INV_X1 U7814 ( .A(n7757), .ZN(n7655) );
  NAND2_X1 U7815 ( .A1(n4333), .A2(n7655), .ZN(n6216) );
  NAND2_X1 U7816 ( .A1(n8176), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6215) );
  OR2_X1 U7817 ( .A1(n7672), .A2(n6286), .ZN(n6219) );
  NAND2_X1 U7818 ( .A1(n6220), .A2(n6219), .ZN(n6221) );
  XNOR2_X1 U7819 ( .A(n6221), .B(n6546), .ZN(n6223) );
  NOR2_X1 U7820 ( .A1(n7672), .A2(n6570), .ZN(n6222) );
  AOI21_X1 U7821 ( .B1(n7763), .B2(n6305), .A(n6222), .ZN(n6224) );
  XNOR2_X1 U7822 ( .A(n6223), .B(n6224), .ZN(n7756) );
  INV_X1 U7823 ( .A(n6223), .ZN(n6225) );
  NAND2_X1 U7824 ( .A1(n6225), .A2(n6224), .ZN(n6226) );
  NAND2_X1 U7825 ( .A1(n6822), .A2(n8291), .ZN(n6232) );
  NOR2_X1 U7826 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n6227) );
  AND2_X1 U7827 ( .A1(n6228), .A2(n6227), .ZN(n6245) );
  INV_X1 U7828 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6229) );
  OR2_X1 U7829 ( .A1(n6273), .A2(n6244), .ZN(n6230) );
  XNOR2_X1 U7830 ( .A(n6230), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7465) );
  AOI22_X1 U7831 ( .A1(n6412), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6411), .B2(
        n7465), .ZN(n6231) );
  NAND2_X1 U7832 ( .A1(n7864), .A2(n6131), .ZN(n6240) );
  NAND2_X1 U7833 ( .A1(n6250), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6252) );
  NAND2_X1 U7834 ( .A1(n6252), .A2(n6233), .ZN(n6234) );
  NAND2_X1 U7835 ( .A1(n6280), .A2(n6234), .ZN(n9813) );
  INV_X1 U7836 ( .A(n9813), .ZN(n7791) );
  NAND2_X1 U7837 ( .A1(n4332), .A2(n7791), .ZN(n6238) );
  NAND2_X1 U7838 ( .A1(n4335), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U7839 ( .A1(n8176), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7840 ( .A1(n8177), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6235) );
  OR2_X1 U7841 ( .A1(n7863), .A2(n6103), .ZN(n6239) );
  NAND2_X1 U7842 ( .A1(n6240), .A2(n6239), .ZN(n6241) );
  XNOR2_X1 U7843 ( .A(n6241), .B(n6546), .ZN(n9796) );
  NAND2_X1 U7844 ( .A1(n7864), .A2(n6305), .ZN(n6243) );
  OR2_X1 U7845 ( .A1(n7863), .A2(n6570), .ZN(n6242) );
  NAND2_X1 U7846 ( .A1(n6243), .A2(n6242), .ZN(n9797) );
  NAND2_X1 U7847 ( .A1(n9796), .A2(n9797), .ZN(n9795) );
  INV_X1 U7848 ( .A(n9795), .ZN(n6262) );
  NAND2_X1 U7849 ( .A1(n6716), .A2(n8291), .ZN(n6248) );
  OR2_X1 U7850 ( .A1(n6245), .A2(n6244), .ZN(n6246) );
  XNOR2_X1 U7851 ( .A(n6246), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7200) );
  AOI22_X1 U7852 ( .A1(n6412), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6411), .B2(
        n7200), .ZN(n6247) );
  NAND2_X1 U7853 ( .A1(n9128), .A2(n6131), .ZN(n6258) );
  OR2_X1 U7854 ( .A1(n6250), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6251) );
  AND2_X1 U7855 ( .A1(n6252), .A2(n6251), .ZN(n7676) );
  NAND2_X1 U7856 ( .A1(n4333), .A2(n7676), .ZN(n6256) );
  NAND2_X1 U7857 ( .A1(n4335), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U7858 ( .A1(n8176), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U7859 ( .A1(n8177), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6253) );
  OR2_X1 U7860 ( .A1(n9804), .A2(n6103), .ZN(n6257) );
  NAND2_X1 U7861 ( .A1(n6258), .A2(n6257), .ZN(n6259) );
  XNOR2_X1 U7862 ( .A(n6259), .B(n6587), .ZN(n9794) );
  NOR2_X1 U7863 ( .A1(n9804), .A2(n6570), .ZN(n6260) );
  AOI21_X1 U7864 ( .B1(n9128), .B2(n6305), .A(n6260), .ZN(n9121) );
  NOR2_X1 U7865 ( .A1(n9794), .A2(n9121), .ZN(n6261) );
  NAND2_X1 U7866 ( .A1(n9120), .A2(n6263), .ZN(n6270) );
  INV_X1 U7867 ( .A(n9796), .ZN(n6268) );
  NAND2_X1 U7868 ( .A1(n9794), .A2(n9121), .ZN(n6264) );
  NAND2_X1 U7869 ( .A1(n6264), .A2(n9797), .ZN(n6267) );
  INV_X1 U7870 ( .A(n6264), .ZN(n6266) );
  INV_X1 U7871 ( .A(n9797), .ZN(n6265) );
  AOI22_X1 U7872 ( .A1(n6268), .A2(n6267), .B1(n6266), .B2(n6265), .ZN(n6269)
         );
  NAND2_X1 U7873 ( .A1(n6270), .A2(n6269), .ZN(n9161) );
  OR2_X1 U7874 ( .A1(n6846), .A2(n6271), .ZN(n6277) );
  INV_X1 U7875 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6272) );
  NAND2_X1 U7876 ( .A1(n6273), .A2(n6272), .ZN(n6314) );
  NAND2_X1 U7877 ( .A1(n6314), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6274) );
  INV_X1 U7878 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6312) );
  NAND2_X1 U7879 ( .A1(n6274), .A2(n6312), .ZN(n6294) );
  OR2_X1 U7880 ( .A1(n6274), .A2(n6312), .ZN(n6275) );
  AOI22_X1 U7881 ( .A1(n6412), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6411), .B2(
        n7466), .ZN(n6276) );
  NAND2_X1 U7882 ( .A1(n8177), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U7883 ( .A1(n4335), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6284) );
  INV_X1 U7884 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U7885 ( .A1(n6280), .A2(n6279), .ZN(n6281) );
  AND2_X1 U7886 ( .A1(n6299), .A2(n6281), .ZN(n9166) );
  NAND2_X1 U7887 ( .A1(n4333), .A2(n9166), .ZN(n6283) );
  NAND2_X1 U7888 ( .A1(n8176), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6282) );
  NAND4_X1 U7889 ( .A1(n6285), .A2(n6284), .A3(n6283), .A4(n6282), .ZN(n9284)
         );
  INV_X1 U7890 ( .A(n9284), .ZN(n9805) );
  OAI22_X1 U7891 ( .A1(n9169), .A2(n6249), .B1(n9805), .B2(n6286), .ZN(n6287)
         );
  XNOR2_X1 U7892 ( .A(n6287), .B(n6587), .ZN(n6289) );
  OAI22_X1 U7893 ( .A1(n9169), .A2(n6286), .B1(n9805), .B2(n6570), .ZN(n6290)
         );
  INV_X1 U7894 ( .A(n6290), .ZN(n6288) );
  NAND2_X1 U7895 ( .A1(n6289), .A2(n6288), .ZN(n6293) );
  INV_X1 U7896 ( .A(n6289), .ZN(n6291) );
  NAND2_X1 U7897 ( .A1(n6291), .A2(n6290), .ZN(n6292) );
  AND2_X1 U7898 ( .A1(n6293), .A2(n6292), .ZN(n9162) );
  NAND2_X1 U7899 ( .A1(n6994), .A2(n8291), .ZN(n6297) );
  NAND2_X1 U7900 ( .A1(n6294), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6295) );
  XNOR2_X1 U7901 ( .A(n6295), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7717) );
  AOI22_X1 U7902 ( .A1(n6412), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6411), .B2(
        n7717), .ZN(n6296) );
  NAND2_X1 U7903 ( .A1(n8177), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6304) );
  NAND2_X1 U7904 ( .A1(n4335), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U7905 ( .A1(n6299), .A2(n6298), .ZN(n6300) );
  AND2_X1 U7906 ( .A1(n6320), .A2(n6300), .ZN(n9222) );
  NAND2_X1 U7907 ( .A1(n4333), .A2(n9222), .ZN(n6302) );
  NAND2_X1 U7908 ( .A1(n8176), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6301) );
  NAND4_X1 U7909 ( .A1(n6304), .A2(n6303), .A3(n6302), .A4(n6301), .ZN(n9283)
         );
  OAI22_X1 U7910 ( .A1(n9225), .A2(n6249), .B1(n8138), .B2(n6103), .ZN(n6306)
         );
  XNOR2_X1 U7911 ( .A(n6306), .B(n6587), .ZN(n6307) );
  OAI22_X1 U7912 ( .A1(n9225), .A2(n6286), .B1(n8138), .B2(n6570), .ZN(n6308)
         );
  XNOR2_X1 U7913 ( .A(n6307), .B(n6308), .ZN(n9217) );
  INV_X1 U7914 ( .A(n6307), .ZN(n6309) );
  OR2_X1 U7915 ( .A1(n6309), .A2(n6308), .ZN(n6310) );
  NAND2_X1 U7916 ( .A1(n7043), .A2(n8291), .ZN(n6318) );
  INV_X1 U7917 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6311) );
  NAND2_X1 U7918 ( .A1(n6312), .A2(n6311), .ZN(n6313) );
  OAI21_X1 U7919 ( .B1(n6314), .B2(n6313), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6315) );
  MUX2_X1 U7920 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6315), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n6316) );
  AND2_X1 U7921 ( .A1(n4495), .A2(n6316), .ZN(n7963) );
  AOI22_X1 U7922 ( .A1(n6412), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6411), .B2(
        n7963), .ZN(n6317) );
  NAND2_X1 U7923 ( .A1(n9770), .A2(n6131), .ZN(n6327) );
  NAND2_X1 U7924 ( .A1(n8177), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6325) );
  NAND2_X1 U7925 ( .A1(n4335), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6324) );
  NAND2_X1 U7926 ( .A1(n6320), .A2(n6319), .ZN(n6321) );
  AND2_X1 U7927 ( .A1(n6340), .A2(n6321), .ZN(n9616) );
  NAND2_X1 U7928 ( .A1(n4332), .A2(n9616), .ZN(n6323) );
  NAND2_X1 U7929 ( .A1(n8176), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6322) );
  NAND4_X1 U7930 ( .A1(n6325), .A2(n6324), .A3(n6323), .A4(n6322), .ZN(n9282)
         );
  NAND2_X1 U7931 ( .A1(n9282), .A2(n6305), .ZN(n6326) );
  NAND2_X1 U7932 ( .A1(n6327), .A2(n6326), .ZN(n6328) );
  XNOR2_X1 U7933 ( .A(n6328), .B(n6587), .ZN(n6329) );
  NAND2_X1 U7934 ( .A1(n6330), .A2(n6329), .ZN(n6334) );
  NAND2_X1 U7935 ( .A1(n9770), .A2(n6305), .ZN(n6332) );
  NAND2_X1 U7936 ( .A1(n9282), .A2(n6584), .ZN(n6331) );
  NAND2_X1 U7937 ( .A1(n6332), .A2(n6331), .ZN(n9106) );
  NAND2_X1 U7938 ( .A1(n7180), .A2(n8291), .ZN(n6337) );
  NAND2_X1 U7939 ( .A1(n4495), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6335) );
  XNOR2_X1 U7940 ( .A(n6335), .B(P1_IR_REG_15__SCAN_IN), .ZN(n8119) );
  AOI22_X1 U7941 ( .A1(n6412), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6411), .B2(
        n8119), .ZN(n6336) );
  NAND2_X1 U7942 ( .A1(n9766), .A2(n6131), .ZN(n6347) );
  NAND2_X1 U7943 ( .A1(n4335), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6345) );
  NAND2_X1 U7944 ( .A1(n8176), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6344) );
  INV_X1 U7945 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6339) );
  NAND2_X1 U7946 ( .A1(n6340), .A2(n6339), .ZN(n6341) );
  AND2_X1 U7947 ( .A1(n6355), .A2(n6341), .ZN(n9596) );
  NAND2_X1 U7948 ( .A1(n4332), .A2(n9596), .ZN(n6343) );
  NAND2_X1 U7949 ( .A1(n8177), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6342) );
  NAND4_X1 U7950 ( .A1(n6345), .A2(n6344), .A3(n6343), .A4(n6342), .ZN(n9281)
         );
  NAND2_X1 U7951 ( .A1(n9281), .A2(n6305), .ZN(n6346) );
  NAND2_X1 U7952 ( .A1(n6347), .A2(n6346), .ZN(n6348) );
  XNOR2_X1 U7953 ( .A(n6348), .B(n6587), .ZN(n6369) );
  NAND2_X1 U7954 ( .A1(n6368), .A2(n6369), .ZN(n9180) );
  INV_X1 U7955 ( .A(n9180), .ZN(n6366) );
  NAND2_X1 U7956 ( .A1(n7245), .A2(n8291), .ZN(n6352) );
  NAND2_X1 U7957 ( .A1(n6349), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6350) );
  XNOR2_X1 U7958 ( .A(n6350), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9331) );
  AOI22_X1 U7959 ( .A1(n6412), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6411), .B2(
        n9331), .ZN(n6351) );
  NAND2_X1 U7960 ( .A1(n9761), .A2(n6131), .ZN(n6362) );
  NAND2_X1 U7961 ( .A1(n8177), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6360) );
  NAND2_X1 U7962 ( .A1(n4335), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6359) );
  INV_X1 U7963 ( .A(n6355), .ZN(n6353) );
  INV_X1 U7964 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6354) );
  NAND2_X1 U7965 ( .A1(n6355), .A2(n6354), .ZN(n6356) );
  AND2_X1 U7966 ( .A1(n6381), .A2(n6356), .ZN(n9578) );
  NAND2_X1 U7967 ( .A1(n4332), .A2(n9578), .ZN(n6358) );
  NAND2_X1 U7968 ( .A1(n8176), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6357) );
  OR2_X1 U7969 ( .A1(n9261), .A2(n6103), .ZN(n6361) );
  NAND2_X1 U7970 ( .A1(n6362), .A2(n6361), .ZN(n6363) );
  XNOR2_X1 U7971 ( .A(n6363), .B(n6546), .ZN(n6372) );
  NAND2_X1 U7972 ( .A1(n9761), .A2(n6305), .ZN(n6365) );
  OR2_X1 U7973 ( .A1(n9261), .A2(n6570), .ZN(n6364) );
  NAND2_X1 U7974 ( .A1(n6365), .A2(n6364), .ZN(n6373) );
  NAND2_X1 U7975 ( .A1(n6372), .A2(n6373), .ZN(n9188) );
  AND2_X1 U7976 ( .A1(n9281), .A2(n6584), .ZN(n6367) );
  AOI21_X1 U7977 ( .B1(n9766), .B2(n6305), .A(n6367), .ZN(n9258) );
  AND2_X1 U7978 ( .A1(n9258), .A2(n9188), .ZN(n9182) );
  INV_X1 U7979 ( .A(n6369), .ZN(n6370) );
  NAND2_X1 U7980 ( .A1(n9182), .A2(n9181), .ZN(n6376) );
  INV_X1 U7981 ( .A(n6372), .ZN(n6375) );
  INV_X1 U7982 ( .A(n6373), .ZN(n6374) );
  NAND2_X1 U7983 ( .A1(n6375), .A2(n6374), .ZN(n9187) );
  NAND2_X1 U7984 ( .A1(n7267), .A2(n8291), .ZN(n6379) );
  XNOR2_X1 U7985 ( .A(n6377), .B(P1_IR_REG_17__SCAN_IN), .ZN(n8125) );
  AOI22_X1 U7986 ( .A1(n6412), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6411), .B2(
        n8125), .ZN(n6378) );
  NAND2_X1 U7987 ( .A1(n9561), .A2(n6131), .ZN(n6388) );
  INV_X1 U7988 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6380) );
  NAND2_X1 U7989 ( .A1(n6381), .A2(n6380), .ZN(n6382) );
  AND2_X1 U7990 ( .A1(n6416), .A2(n6382), .ZN(n9562) );
  NAND2_X1 U7991 ( .A1(n9562), .A2(n4332), .ZN(n6386) );
  NAND2_X1 U7992 ( .A1(n4335), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6385) );
  NAND2_X1 U7993 ( .A1(n8177), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6384) );
  NAND2_X1 U7994 ( .A1(n8176), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6383) );
  NAND4_X1 U7995 ( .A1(n6386), .A2(n6385), .A3(n6384), .A4(n6383), .ZN(n9279)
         );
  NAND2_X1 U7996 ( .A1(n9279), .A2(n6305), .ZN(n6387) );
  NAND2_X1 U7997 ( .A1(n6388), .A2(n6387), .ZN(n6389) );
  XNOR2_X1 U7998 ( .A(n6389), .B(n6546), .ZN(n6391) );
  AND2_X1 U7999 ( .A1(n9279), .A2(n6584), .ZN(n6390) );
  AOI21_X1 U8000 ( .B1(n9561), .B2(n6305), .A(n6390), .ZN(n6392) );
  XNOR2_X1 U8001 ( .A(n6391), .B(n6392), .ZN(n9198) );
  INV_X1 U8002 ( .A(n6391), .ZN(n6393) );
  NAND2_X1 U8003 ( .A1(n6393), .A2(n6392), .ZN(n6394) );
  NAND2_X1 U8004 ( .A1(n7435), .A2(n8291), .ZN(n6397) );
  AOI22_X1 U8005 ( .A1(n6412), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8383), .B2(
        n6411), .ZN(n6396) );
  NAND2_X1 U8006 ( .A1(n9528), .A2(n6131), .ZN(n6403) );
  NAND2_X1 U8007 ( .A1(n6418), .A2(n8134), .ZN(n6399) );
  NAND2_X1 U8008 ( .A1(n6440), .A2(n6399), .ZN(n9529) );
  AOI22_X1 U8009 ( .A1(n4335), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n8177), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n6401) );
  NAND2_X1 U8010 ( .A1(n8176), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6400) );
  OAI211_X1 U8011 ( .C1(n9529), .C2(n6561), .A(n6401), .B(n6400), .ZN(n9278)
         );
  NAND2_X1 U8012 ( .A1(n9278), .A2(n6305), .ZN(n6402) );
  NAND2_X1 U8013 ( .A1(n6403), .A2(n6402), .ZN(n6404) );
  XNOR2_X1 U8014 ( .A(n6404), .B(n6546), .ZN(n6430) );
  NAND2_X1 U8015 ( .A1(n9528), .A2(n6305), .ZN(n6406) );
  NAND2_X1 U8016 ( .A1(n9278), .A2(n6584), .ZN(n6405) );
  NAND2_X1 U8017 ( .A1(n6406), .A2(n6405), .ZN(n9133) );
  NAND2_X1 U8018 ( .A1(n7433), .A2(n8291), .ZN(n6414) );
  OR2_X1 U8019 ( .A1(n6408), .A2(n6407), .ZN(n6409) );
  AND2_X1 U8020 ( .A1(n6410), .A2(n6409), .ZN(n8126) );
  AOI22_X1 U8021 ( .A1(n6412), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6411), .B2(
        n8126), .ZN(n6413) );
  NAND2_X1 U8022 ( .A1(n9751), .A2(n6305), .ZN(n6425) );
  INV_X1 U8023 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9546) );
  INV_X1 U8024 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6415) );
  NAND2_X1 U8025 ( .A1(n6416), .A2(n6415), .ZN(n6417) );
  NAND2_X1 U8026 ( .A1(n6418), .A2(n6417), .ZN(n9545) );
  OR2_X1 U8027 ( .A1(n9545), .A2(n6561), .ZN(n6422) );
  NAND2_X1 U8028 ( .A1(n4335), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6420) );
  NAND2_X1 U8029 ( .A1(n8177), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6419) );
  AND2_X1 U8030 ( .A1(n6420), .A2(n6419), .ZN(n6421) );
  OAI211_X1 U8031 ( .C1(n6423), .C2(n9546), .A(n6422), .B(n6421), .ZN(n9522)
         );
  NAND2_X1 U8032 ( .A1(n9522), .A2(n6584), .ZN(n6424) );
  NAND2_X1 U8033 ( .A1(n6425), .A2(n6424), .ZN(n9239) );
  NAND2_X1 U8034 ( .A1(n9751), .A2(n6131), .ZN(n6427) );
  NAND2_X1 U8035 ( .A1(n9522), .A2(n6305), .ZN(n6426) );
  NAND2_X1 U8036 ( .A1(n6427), .A2(n6426), .ZN(n6428) );
  XNOR2_X1 U8037 ( .A(n6428), .B(n6546), .ZN(n6431) );
  AOI22_X1 U8038 ( .A1(n6430), .A2(n9133), .B1(n9239), .B2(n6431), .ZN(n6429)
         );
  INV_X1 U8039 ( .A(n6430), .ZN(n9134) );
  OAI21_X1 U8040 ( .B1(n6431), .B2(n9239), .A(n9133), .ZN(n6433) );
  NOR2_X1 U8041 ( .A1(n9133), .A2(n9239), .ZN(n6432) );
  INV_X1 U8042 ( .A(n6431), .ZN(n9132) );
  AOI22_X1 U8043 ( .A1(n9134), .A2(n6433), .B1(n6432), .B2(n9132), .ZN(n6434)
         );
  NAND2_X1 U8044 ( .A1(n7601), .A2(n8291), .ZN(n6437) );
  INV_X1 U8045 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7604) );
  OR2_X1 U8046 ( .A1(n8293), .A2(n7604), .ZN(n6436) );
  NAND2_X1 U8047 ( .A1(n9744), .A2(n6131), .ZN(n6449) );
  INV_X1 U8048 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U8049 ( .A1(n6440), .A2(n6439), .ZN(n6441) );
  NAND2_X1 U8050 ( .A1(n6459), .A2(n6441), .ZN(n9511) );
  OR2_X1 U8051 ( .A1(n9511), .A2(n6561), .ZN(n6447) );
  INV_X1 U8052 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n6444) );
  NAND2_X1 U8053 ( .A1(n8177), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6443) );
  NAND2_X1 U8054 ( .A1(n8176), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6442) );
  OAI211_X1 U8055 ( .C1(n6620), .C2(n6444), .A(n6443), .B(n6442), .ZN(n6445)
         );
  INV_X1 U8056 ( .A(n6445), .ZN(n6446) );
  NAND2_X1 U8057 ( .A1(n6447), .A2(n6446), .ZN(n9525) );
  NAND2_X1 U8058 ( .A1(n9525), .A2(n6305), .ZN(n6448) );
  NAND2_X1 U8059 ( .A1(n6449), .A2(n6448), .ZN(n6450) );
  XNOR2_X1 U8060 ( .A(n6450), .B(n6587), .ZN(n9206) );
  AND2_X1 U8061 ( .A1(n9525), .A2(n6584), .ZN(n6451) );
  AOI21_X1 U8062 ( .B1(n9744), .B2(n6305), .A(n6451), .ZN(n9205) );
  AND2_X1 U8063 ( .A1(n9206), .A2(n9205), .ZN(n6455) );
  INV_X1 U8064 ( .A(n9206), .ZN(n6453) );
  INV_X1 U8065 ( .A(n9205), .ZN(n6452) );
  NAND2_X1 U8066 ( .A1(n6453), .A2(n6452), .ZN(n6454) );
  NAND2_X1 U8067 ( .A1(n7694), .A2(n8291), .ZN(n6457) );
  OR2_X1 U8068 ( .A1(n8293), .A2(n7707), .ZN(n6456) );
  NAND2_X2 U8069 ( .A1(n6457), .A2(n6456), .ZN(n9739) );
  NAND2_X1 U8070 ( .A1(n9739), .A2(n6131), .ZN(n6468) );
  INV_X1 U8071 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U8072 ( .A1(n6459), .A2(n6458), .ZN(n6460) );
  AND2_X1 U8073 ( .A1(n6478), .A2(n6460), .ZN(n9498) );
  NAND2_X1 U8074 ( .A1(n9498), .A2(n4333), .ZN(n6466) );
  INV_X1 U8075 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U8076 ( .A1(n8177), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6462) );
  NAND2_X1 U8077 ( .A1(n8176), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6461) );
  OAI211_X1 U8078 ( .C1(n6620), .C2(n6463), .A(n6462), .B(n6461), .ZN(n6464)
         );
  INV_X1 U8079 ( .A(n6464), .ZN(n6465) );
  NAND2_X1 U8080 ( .A1(n6466), .A2(n6465), .ZN(n9277) );
  NAND2_X1 U8081 ( .A1(n9277), .A2(n6305), .ZN(n6467) );
  NAND2_X1 U8082 ( .A1(n6468), .A2(n6467), .ZN(n6469) );
  XNOR2_X1 U8083 ( .A(n6469), .B(n6587), .ZN(n6472) );
  AND2_X1 U8084 ( .A1(n9277), .A2(n6584), .ZN(n6470) );
  AOI21_X1 U8085 ( .B1(n9739), .B2(n6305), .A(n6470), .ZN(n6471) );
  XNOR2_X1 U8086 ( .A(n6472), .B(n6471), .ZN(n9153) );
  NAND2_X1 U8087 ( .A1(n6472), .A2(n6471), .ZN(n6473) );
  NAND2_X1 U8088 ( .A1(n7812), .A2(n8291), .ZN(n6475) );
  OR2_X1 U8089 ( .A1(n8293), .A2(n7855), .ZN(n6474) );
  INV_X1 U8090 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6477) );
  NAND2_X1 U8091 ( .A1(n6478), .A2(n6477), .ZN(n6479) );
  NAND2_X1 U8092 ( .A1(n6493), .A2(n6479), .ZN(n9476) );
  OR2_X1 U8093 ( .A1(n9476), .A2(n6561), .ZN(n6485) );
  INV_X1 U8094 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n6482) );
  NAND2_X1 U8095 ( .A1(n4335), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6481) );
  NAND2_X1 U8096 ( .A1(n8176), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6480) );
  OAI211_X1 U8097 ( .C1(n6542), .C2(n6482), .A(n6481), .B(n6480), .ZN(n6483)
         );
  INV_X1 U8098 ( .A(n6483), .ZN(n6484) );
  OAI22_X1 U8099 ( .A1(n9479), .A2(n6249), .B1(n9491), .B2(n6103), .ZN(n6486)
         );
  XNOR2_X1 U8100 ( .A(n6486), .B(n6587), .ZN(n6487) );
  NAND2_X1 U8101 ( .A1(n6488), .A2(n6487), .ZN(n9230) );
  OAI22_X1 U8102 ( .A1(n9479), .A2(n6286), .B1(n9491), .B2(n6570), .ZN(n9229)
         );
  NAND2_X1 U8103 ( .A1(n7906), .A2(n8291), .ZN(n6490) );
  OR2_X1 U8104 ( .A1(n8293), .A2(n7908), .ZN(n6489) );
  INV_X1 U8105 ( .A(n6493), .ZN(n6491) );
  INV_X1 U8106 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6492) );
  NAND2_X1 U8107 ( .A1(n6493), .A2(n6492), .ZN(n6494) );
  NAND2_X1 U8108 ( .A1(n6506), .A2(n6494), .ZN(n9463) );
  OR2_X1 U8109 ( .A1(n9463), .A2(n6561), .ZN(n6499) );
  INV_X1 U8110 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9659) );
  NAND2_X1 U8111 ( .A1(n8177), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6496) );
  NAND2_X1 U8112 ( .A1(n8176), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6495) );
  OAI211_X1 U8113 ( .C1(n6620), .C2(n9659), .A(n6496), .B(n6495), .ZN(n6497)
         );
  INV_X1 U8114 ( .A(n6497), .ZN(n6498) );
  NAND2_X1 U8115 ( .A1(n6499), .A2(n6498), .ZN(n9275) );
  AOI22_X1 U8116 ( .A1(n9462), .A2(n6131), .B1(n6305), .B2(n9275), .ZN(n6500)
         );
  XOR2_X1 U8117 ( .A(n6546), .B(n6500), .Z(n6502) );
  INV_X1 U8118 ( .A(n9275), .ZN(n8164) );
  OAI22_X1 U8119 ( .A1(n9731), .A2(n6286), .B1(n8164), .B2(n6570), .ZN(n6501)
         );
  NOR2_X1 U8120 ( .A1(n6502), .A2(n6501), .ZN(n6503) );
  AOI21_X1 U8121 ( .B1(n6502), .B2(n6501), .A(n6503), .ZN(n9114) );
  NAND2_X1 U8122 ( .A1(n9231), .A2(n9114), .ZN(n8450) );
  INV_X1 U8123 ( .A(n6503), .ZN(n8452) );
  NAND2_X1 U8124 ( .A1(n7982), .A2(n8291), .ZN(n6505) );
  OR2_X1 U8125 ( .A1(n8293), .A2(n7985), .ZN(n6504) );
  INV_X1 U8126 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8457) );
  NAND2_X1 U8127 ( .A1(n6506), .A2(n8457), .ZN(n6507) );
  NAND2_X1 U8128 ( .A1(n6526), .A2(n6507), .ZN(n9446) );
  OR2_X1 U8129 ( .A1(n9446), .A2(n6561), .ZN(n6513) );
  INV_X1 U8130 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n6510) );
  NAND2_X1 U8131 ( .A1(n4335), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U8132 ( .A1(n8176), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6508) );
  OAI211_X1 U8133 ( .C1(n6542), .C2(n6510), .A(n6509), .B(n6508), .ZN(n6511)
         );
  INV_X1 U8134 ( .A(n6511), .ZN(n6512) );
  OAI22_X1 U8135 ( .A1(n9445), .A2(n6249), .B1(n9172), .B2(n6286), .ZN(n6514)
         );
  XNOR2_X1 U8136 ( .A(n6514), .B(n6587), .ZN(n6517) );
  OR2_X1 U8137 ( .A1(n9445), .A2(n6103), .ZN(n6516) );
  NAND2_X1 U8138 ( .A1(n9274), .A2(n6584), .ZN(n6515) );
  NAND2_X1 U8139 ( .A1(n6517), .A2(n6518), .ZN(n6522) );
  INV_X1 U8140 ( .A(n6517), .ZN(n6520) );
  INV_X1 U8141 ( .A(n6518), .ZN(n6519) );
  NAND2_X1 U8142 ( .A1(n6520), .A2(n6519), .ZN(n6521) );
  NAND2_X1 U8143 ( .A1(n6522), .A2(n6521), .ZN(n8451) );
  INV_X1 U8144 ( .A(n6522), .ZN(n6523) );
  NAND2_X1 U8145 ( .A1(n8028), .A2(n8291), .ZN(n6525) );
  OR2_X1 U8146 ( .A1(n8293), .A2(n8031), .ZN(n6524) );
  INV_X1 U8147 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9174) );
  NAND2_X1 U8148 ( .A1(n6526), .A2(n9174), .ZN(n6527) );
  NAND2_X1 U8149 ( .A1(n9430), .A2(n4332), .ZN(n6532) );
  INV_X1 U8150 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9650) );
  NAND2_X1 U8151 ( .A1(n6089), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U8152 ( .A1(n8176), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6528) );
  OAI211_X1 U8153 ( .C1(n6620), .C2(n9650), .A(n6529), .B(n6528), .ZN(n6530)
         );
  INV_X1 U8154 ( .A(n6530), .ZN(n6531) );
  AOI22_X1 U8155 ( .A1(n8186), .A2(n6131), .B1(n6305), .B2(n9273), .ZN(n6533)
         );
  XNOR2_X1 U8156 ( .A(n6533), .B(n6546), .ZN(n6550) );
  AND2_X1 U8157 ( .A1(n9273), .A2(n6584), .ZN(n6534) );
  AOI21_X1 U8158 ( .B1(n8186), .B2(n6305), .A(n6534), .ZN(n6551) );
  XNOR2_X1 U8159 ( .A(n6550), .B(n6551), .ZN(n9170) );
  OR2_X1 U8160 ( .A1(n8293), .A2(n8054), .ZN(n6535) );
  AND2_X2 U8161 ( .A1(n6536), .A2(n6535), .ZN(n9413) );
  INV_X1 U8162 ( .A(n6538), .ZN(n6537) );
  NAND2_X1 U8163 ( .A1(n6537), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6559) );
  INV_X1 U8164 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9252) );
  NAND2_X1 U8165 ( .A1(n6538), .A2(n9252), .ZN(n6539) );
  NAND2_X1 U8166 ( .A1(n6559), .A2(n6539), .ZN(n9414) );
  INV_X1 U8167 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10159) );
  NAND2_X1 U8168 ( .A1(n4335), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6541) );
  NAND2_X1 U8169 ( .A1(n8176), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6540) );
  OAI211_X1 U8170 ( .C1(n6542), .C2(n10159), .A(n6541), .B(n6540), .ZN(n6543)
         );
  INV_X1 U8171 ( .A(n6543), .ZN(n6544) );
  OAI22_X1 U8172 ( .A1(n9413), .A2(n6249), .B1(n9173), .B2(n6286), .ZN(n6547)
         );
  XNOR2_X1 U8173 ( .A(n6547), .B(n6546), .ZN(n6555) );
  OR2_X1 U8174 ( .A1(n9413), .A2(n6103), .ZN(n6549) );
  NAND2_X1 U8175 ( .A1(n9395), .A2(n6584), .ZN(n6548) );
  NAND2_X1 U8176 ( .A1(n6549), .A2(n6548), .ZN(n6554) );
  XNOR2_X1 U8177 ( .A(n6555), .B(n6554), .ZN(n9247) );
  INV_X1 U8178 ( .A(n6550), .ZN(n6553) );
  INV_X1 U8179 ( .A(n6551), .ZN(n6552) );
  NOR2_X1 U8180 ( .A1(n6553), .A2(n6552), .ZN(n9248) );
  NAND2_X1 U8181 ( .A1(n9099), .A2(n8291), .ZN(n6557) );
  OR2_X1 U8182 ( .A1(n8293), .A2(n9790), .ZN(n6556) );
  NAND2_X1 U8183 ( .A1(n9399), .A2(n6131), .ZN(n6568) );
  INV_X1 U8184 ( .A(n6559), .ZN(n6558) );
  NAND2_X1 U8185 ( .A1(n6558), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6577) );
  INV_X1 U8186 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n10145) );
  NAND2_X1 U8187 ( .A1(n6559), .A2(n10145), .ZN(n6560) );
  NAND2_X1 U8188 ( .A1(n6577), .A2(n6560), .ZN(n9400) );
  INV_X1 U8189 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9642) );
  NAND2_X1 U8190 ( .A1(n8177), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6563) );
  NAND2_X1 U8191 ( .A1(n8176), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6562) );
  OAI211_X1 U8192 ( .C1(n6620), .C2(n9642), .A(n6563), .B(n6562), .ZN(n6564)
         );
  INV_X1 U8193 ( .A(n6564), .ZN(n6565) );
  NAND2_X1 U8194 ( .A1(n9272), .A2(n6305), .ZN(n6567) );
  NAND2_X1 U8195 ( .A1(n6568), .A2(n6567), .ZN(n6569) );
  XNOR2_X1 U8196 ( .A(n6569), .B(n6587), .ZN(n6573) );
  NOR2_X1 U8197 ( .A1(n9251), .A2(n6570), .ZN(n6571) );
  AOI21_X1 U8198 ( .B1(n9399), .B2(n6305), .A(n6571), .ZN(n6572) );
  NAND2_X1 U8199 ( .A1(n6573), .A2(n6572), .ZN(n6634) );
  OAI21_X1 U8200 ( .B1(n6573), .B2(n6572), .A(n6634), .ZN(n6642) );
  NAND2_X1 U8201 ( .A1(n9096), .A2(n8291), .ZN(n6575) );
  OR2_X1 U8202 ( .A1(n8293), .A2(n9787), .ZN(n6574) );
  NAND2_X1 U8203 ( .A1(n9709), .A2(n6305), .ZN(n6586) );
  INV_X1 U8204 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6576) );
  NAND2_X1 U8205 ( .A1(n6577), .A2(n6576), .ZN(n6578) );
  NAND2_X1 U8206 ( .A1(n9386), .A2(n4333), .ZN(n6583) );
  INV_X1 U8207 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9636) );
  NAND2_X1 U8208 ( .A1(n6089), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6580) );
  NAND2_X1 U8209 ( .A1(n8176), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6579) );
  OAI211_X1 U8210 ( .C1(n6620), .C2(n9636), .A(n6580), .B(n6579), .ZN(n6581)
         );
  INV_X1 U8211 ( .A(n6581), .ZN(n6582) );
  NAND2_X1 U8212 ( .A1(n9271), .A2(n6584), .ZN(n6585) );
  NAND2_X1 U8213 ( .A1(n6586), .A2(n6585), .ZN(n6588) );
  XNOR2_X1 U8214 ( .A(n6588), .B(n6587), .ZN(n6591) );
  NAND2_X1 U8215 ( .A1(n9709), .A2(n6131), .ZN(n6589) );
  OAI21_X1 U8216 ( .B1(n9397), .B2(n6286), .A(n6589), .ZN(n6590) );
  XNOR2_X1 U8217 ( .A(n6591), .B(n6590), .ZN(n6613) );
  INV_X1 U8218 ( .A(n6613), .ZN(n6635) );
  NAND2_X1 U8219 ( .A1(n8032), .A2(P1_B_REG_SCAN_IN), .ZN(n6593) );
  MUX2_X1 U8220 ( .A(n6593), .B(P1_B_REG_SCAN_IN), .S(n6592), .Z(n6594) );
  NOR4_X1 U8221 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n6598) );
  NOR4_X1 U8222 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n6597) );
  NOR4_X1 U8223 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6596) );
  NOR4_X1 U8224 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n6595) );
  AND4_X1 U8225 ( .A1(n6598), .A2(n6597), .A3(n6596), .A4(n6595), .ZN(n6604)
         );
  NOR2_X1 U8226 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n6602) );
  NOR4_X1 U8227 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6601) );
  NOR4_X1 U8228 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6600) );
  NOR4_X1 U8229 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n6599) );
  AND4_X1 U8230 ( .A1(n6602), .A2(n6601), .A3(n6600), .A4(n6599), .ZN(n6603)
         );
  NAND2_X1 U8231 ( .A1(n6604), .A2(n6603), .ZN(n6889) );
  INV_X1 U8232 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6605) );
  OR2_X1 U8233 ( .A1(n6889), .A2(n6605), .ZN(n6608) );
  INV_X1 U8234 ( .A(n6606), .ZN(n8055) );
  NAND2_X1 U8235 ( .A1(n8055), .A2(n8032), .ZN(n9776) );
  INV_X1 U8236 ( .A(n9776), .ZN(n6607) );
  AOI21_X1 U8237 ( .B1(n6890), .B2(n6608), .A(n6607), .ZN(n7155) );
  INV_X1 U8238 ( .A(n6592), .ZN(n7986) );
  NAND2_X1 U8239 ( .A1(n7155), .A2(n7156), .ZN(n6628) );
  NAND2_X1 U8240 ( .A1(n6610), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6611) );
  NAND2_X1 U8241 ( .A1(n9881), .A2(n8367), .ZN(n6612) );
  NAND3_X1 U8242 ( .A1(n6645), .A2(n6613), .A3(n9809), .ZN(n6639) );
  INV_X1 U8243 ( .A(n6614), .ZN(n6626) );
  NOR2_X1 U8244 ( .A1(n7163), .A2(n8372), .ZN(n7483) );
  NAND2_X1 U8245 ( .A1(n6626), .A2(n7483), .ZN(n6616) );
  NOR2_X1 U8246 ( .A1(n7163), .A2(n7162), .ZN(n6888) );
  INV_X1 U8247 ( .A(n6888), .ZN(n6615) );
  NOR2_X2 U8248 ( .A1(n8367), .A2(n4337), .ZN(n9523) );
  NAND2_X1 U8249 ( .A1(n9272), .A2(n9523), .ZN(n6625) );
  INV_X1 U8250 ( .A(n9368), .ZN(n6623) );
  INV_X1 U8251 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n8190) );
  NAND2_X1 U8252 ( .A1(n8177), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6619) );
  NAND2_X1 U8253 ( .A1(n8176), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6618) );
  OAI211_X1 U8254 ( .C1(n6620), .C2(n8190), .A(n6619), .B(n6618), .ZN(n6621)
         );
  AOI21_X1 U8255 ( .B1(n6623), .B2(n4332), .A(n6621), .ZN(n8163) );
  INV_X1 U8256 ( .A(n4337), .ZN(n6763) );
  NOR2_X2 U8257 ( .A1(n8367), .A2(n6763), .ZN(n9524) );
  OR2_X1 U8258 ( .A1(n8163), .A2(n9490), .ZN(n6624) );
  AND2_X1 U8259 ( .A1(n6625), .A2(n6624), .ZN(n9383) );
  NAND2_X1 U8260 ( .A1(n6626), .A2(n8437), .ZN(n9265) );
  OR2_X1 U8261 ( .A1(n8372), .A2(P1_U3086), .ZN(n7602) );
  NAND2_X1 U8262 ( .A1(n7135), .A2(n7602), .ZN(n6627) );
  NAND2_X1 U8263 ( .A1(n6628), .A2(n6627), .ZN(n6630) );
  NOR2_X1 U8264 ( .A1(n8367), .A2(n8437), .ZN(n6887) );
  INV_X1 U8265 ( .A(n6887), .ZN(n6629) );
  NAND2_X1 U8266 ( .A1(n6630), .A2(n6629), .ZN(n7039) );
  OAI21_X1 U8267 ( .B1(n7039), .B2(n6631), .A(P1_STATE_REG_SCAN_IN), .ZN(n6632) );
  OR2_X1 U8268 ( .A1(n6693), .A2(P1_U3086), .ZN(n8448) );
  AOI22_X1 U8269 ( .A1(n9386), .A2(n9267), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6633) );
  OAI21_X1 U8270 ( .B1(n9383), .B2(n9265), .A(n6633), .ZN(n6637) );
  NOR3_X1 U8271 ( .A1(n6635), .A2(n6634), .A3(n9245), .ZN(n6636) );
  AOI211_X1 U8272 ( .C1(n9709), .C2(n6649), .A(n6637), .B(n6636), .ZN(n6638)
         );
  NAND3_X1 U8273 ( .A1(n6640), .A2(n6639), .A3(n6638), .ZN(P1_U3220) );
  INV_X1 U8274 ( .A(n6641), .ZN(n6644) );
  INV_X1 U8275 ( .A(n6642), .ZN(n6643) );
  AOI21_X1 U8276 ( .B1(n4356), .B2(n6644), .A(n6643), .ZN(n6646) );
  OAI21_X1 U8277 ( .B1(n6646), .B2(n6645), .A(n9809), .ZN(n6652) );
  AND2_X1 U8278 ( .A1(n9254), .A2(n9524), .ZN(n9802) );
  NOR2_X1 U8279 ( .A1(n9400), .A2(n9814), .ZN(n6648) );
  OR2_X1 U8280 ( .A1(n9265), .A2(n9488), .ZN(n9803) );
  OAI22_X1 U8281 ( .A1(n9173), .A2(n9803), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10145), .ZN(n6647) );
  AOI211_X1 U8282 ( .C1(n9271), .C2(n9802), .A(n6648), .B(n6647), .ZN(n6651)
         );
  NAND2_X1 U8283 ( .A1(n9399), .A2(n6649), .ZN(n6650) );
  NAND3_X1 U8284 ( .A1(n6652), .A2(n6651), .A3(n6650), .ZN(P1_U3214) );
  NOR2_X1 U8285 ( .A1(n6653), .A2(P1_U3086), .ZN(n6654) );
  INV_X1 U8286 ( .A(n6922), .ZN(n6655) );
  NAND2_X1 U8287 ( .A1(n6656), .A2(n6922), .ZN(n6657) );
  NAND2_X1 U8288 ( .A1(n6703), .A2(n5263), .ZN(n6658) );
  NAND2_X1 U8289 ( .A1(n6658), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NOR2_X1 U8290 ( .A1(n6661), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9781) );
  INV_X2 U8291 ( .A(n9781), .ZN(n9789) );
  AND2_X1 U8292 ( .A1(n6661), .A2(P1_U3086), .ZN(n7905) );
  OAI222_X1 U8293 ( .A1(n9789), .A2(n6659), .B1(n9299), .B2(P1_U3086), .C1(
        n4336), .C2(n6663), .ZN(P1_U3354) );
  OAI222_X1 U8294 ( .A1(n9789), .A2(n6660), .B1(n6876), .B2(P1_U3086), .C1(
        n4336), .C2(n6670), .ZN(P1_U3353) );
  INV_X1 U8295 ( .A(n9100), .ZN(n7434) );
  NAND2_X1 U8296 ( .A1(n6662), .A2(P2_U3151), .ZN(n8046) );
  OAI222_X1 U8297 ( .A1(n6807), .A2(P2_U3151), .B1(n7434), .B2(n5100), .C1(
        n8046), .C2(n6663), .ZN(P2_U3294) );
  OAI222_X1 U8298 ( .A1(n9789), .A2(n6664), .B1(n6776), .B2(P1_U3086), .C1(
        n4336), .C2(n6668), .ZN(P1_U3352) );
  OAI222_X1 U8299 ( .A1(n9789), .A2(n6665), .B1(n6937), .B2(P1_U3086), .C1(
        n4336), .C2(n6667), .ZN(P1_U3351) );
  INV_X1 U8300 ( .A(n6744), .ZN(n7319) );
  CLKBUF_X1 U8301 ( .A(n8046), .Z(n9103) );
  INV_X1 U8302 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6666) );
  OAI222_X1 U8303 ( .A1(P2_U3151), .A2(n7319), .B1(n9103), .B2(n6667), .C1(
        n6666), .C2(n7434), .ZN(P2_U3291) );
  OAI222_X1 U8304 ( .A1(P2_U3151), .A2(n6741), .B1(n9103), .B2(n6668), .C1(
        n5113), .C2(n7434), .ZN(P2_U3292) );
  INV_X1 U8305 ( .A(n4602), .ZN(n6739) );
  INV_X1 U8306 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6669) );
  OAI222_X1 U8307 ( .A1(P2_U3151), .A2(n6739), .B1(n9103), .B2(n6670), .C1(
        n6669), .C2(n7434), .ZN(P2_U3293) );
  INV_X1 U8308 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6671) );
  OAI222_X1 U8309 ( .A1(P2_U3151), .A2(n7338), .B1(n9103), .B2(n6672), .C1(
        n6671), .C2(n7434), .ZN(P2_U3290) );
  INV_X1 U8310 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6673) );
  INV_X1 U8311 ( .A(n6795), .ZN(n6789) );
  OAI222_X1 U8312 ( .A1(n9789), .A2(n6673), .B1(n6789), .B2(P1_U3086), .C1(
        n4336), .C2(n6672), .ZN(P1_U3350) );
  NAND2_X1 U8313 ( .A1(n6918), .A2(n7061), .ZN(n6674) );
  OAI21_X1 U8314 ( .B1(n6918), .B2(n6675), .A(n6674), .ZN(P2_U3377) );
  OAI222_X1 U8315 ( .A1(P2_U3151), .A2(n9959), .B1(n9103), .B2(n6676), .C1(
        n4573), .C2(n7434), .ZN(P2_U3289) );
  INV_X1 U8316 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6677) );
  INV_X1 U8317 ( .A(n6828), .ZN(n6833) );
  OAI222_X1 U8318 ( .A1(n9789), .A2(n6677), .B1(n6833), .B2(P1_U3086), .C1(
        n4336), .C2(n6676), .ZN(P1_U3349) );
  INV_X1 U8319 ( .A(n5688), .ZN(n6678) );
  AND2_X1 U8320 ( .A1(n10119), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8321 ( .A1(n10119), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8322 ( .A1(n10119), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8323 ( .A1(n10119), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8324 ( .A1(n10119), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8325 ( .A1(n10119), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8326 ( .A1(n10119), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8327 ( .A1(n10119), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8328 ( .A1(n10119), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8329 ( .A1(n10119), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8330 ( .A1(n10119), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8331 ( .A1(n10119), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8332 ( .A1(n10119), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8333 ( .A1(n10119), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8334 ( .A1(n10119), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8335 ( .A1(n10119), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8336 ( .A1(n10119), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8337 ( .A1(n10119), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8338 ( .A1(n10119), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8339 ( .A1(n10119), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8340 ( .A1(n10119), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8341 ( .A1(n10119), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  INV_X1 U8342 ( .A(n6679), .ZN(n6680) );
  AOI22_X1 U8343 ( .A1(n10119), .A2(n6682), .B1(n6681), .B2(n6680), .ZN(
        P2_U3376) );
  INV_X1 U8344 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6791) );
  OAI222_X1 U8345 ( .A1(n7341), .A2(P2_U3151), .B1(n7434), .B2(n6791), .C1(
        n6683), .C2(n8046), .ZN(P2_U3288) );
  INV_X1 U8346 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6684) );
  INV_X1 U8347 ( .A(n6851), .ZN(n6861) );
  OAI222_X1 U8348 ( .A1(n9789), .A2(n6684), .B1(n6861), .B2(P1_U3086), .C1(
        n4336), .C2(n6683), .ZN(P1_U3348) );
  INV_X1 U8349 ( .A(n6685), .ZN(n6692) );
  AOI22_X1 U8350 ( .A1(n6960), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9781), .ZN(n6686) );
  OAI21_X1 U8351 ( .B1(n6692), .B2(n4336), .A(n6686), .ZN(P1_U3347) );
  INV_X1 U8352 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10280) );
  NOR2_X1 U8353 ( .A1(n6690), .A2(n10280), .ZN(P2_U3260) );
  INV_X1 U8354 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n10255) );
  NOR2_X1 U8355 ( .A1(n6690), .A2(n10255), .ZN(P2_U3236) );
  INV_X1 U8356 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n10251) );
  NOR2_X1 U8357 ( .A1(n6690), .A2(n10251), .ZN(P2_U3244) );
  INV_X1 U8358 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n6687) );
  NOR2_X1 U8359 ( .A1(n6690), .A2(n6687), .ZN(P2_U3253) );
  INV_X1 U8360 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n6688) );
  NOR2_X1 U8361 ( .A1(n6690), .A2(n6688), .ZN(P2_U3251) );
  INV_X1 U8362 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n10162) );
  NOR2_X1 U8363 ( .A1(n6690), .A2(n10162), .ZN(P2_U3237) );
  INV_X1 U8364 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n6689) );
  NOR2_X1 U8365 ( .A1(n6690), .A2(n6689), .ZN(P2_U3255) );
  INV_X1 U8366 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6691) );
  OAI222_X1 U8367 ( .A1(n7344), .A2(P2_U3151), .B1(n9103), .B2(n6692), .C1(
        n6691), .C2(n7434), .ZN(P2_U3287) );
  INV_X1 U8368 ( .A(n8367), .ZN(n6894) );
  NAND2_X1 U8369 ( .A1(n6693), .A2(n6894), .ZN(n6694) );
  AND2_X1 U8370 ( .A1(n6694), .A2(n6062), .ZN(n6761) );
  INV_X1 U8371 ( .A(n6761), .ZN(n6695) );
  NAND2_X1 U8372 ( .A1(n8444), .A2(n8448), .ZN(n6762) );
  NOR2_X1 U8373 ( .A1(n9824), .A2(P1_U3973), .ZN(P1_U3085) );
  NAND2_X1 U8374 ( .A1(n6901), .A2(P1_U3973), .ZN(n6696) );
  OAI21_X1 U8375 ( .B1(P1_U3973), .B2(n5102), .A(n6696), .ZN(P1_U3554) );
  INV_X1 U8376 ( .A(n6703), .ZN(n6697) );
  INV_X2 U8377 ( .A(n6734), .ZN(n8643) );
  OR2_X1 U8378 ( .A1(n8643), .A2(P2_U3151), .ZN(n9102) );
  NOR2_X1 U8379 ( .A1(n6697), .A2(n9102), .ZN(n6699) );
  INV_X1 U8380 ( .A(n6702), .ZN(n6698) );
  MUX2_X1 U8381 ( .A(n6699), .B(P2_U3893), .S(n6698), .Z(n10003) );
  INV_X1 U8382 ( .A(n6700), .ZN(n6701) );
  INV_X1 U8383 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7068) );
  NOR2_X1 U8384 ( .A1(n6702), .A2(P2_U3151), .ZN(n9097) );
  AND2_X1 U8385 ( .A1(n9097), .A2(n6703), .ZN(n6735) );
  INV_X1 U8386 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6704) );
  OAI21_X1 U8387 ( .B1(n9949), .B2(n6735), .A(n6705), .ZN(n6706) );
  OAI21_X1 U8388 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n7068), .A(n6706), .ZN(n6707) );
  AOI21_X1 U8389 ( .B1(n9962), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n6707), .ZN(
        n6708) );
  OAI21_X1 U8390 ( .B1(n6736), .B2(n9958), .A(n6708), .ZN(P2_U3182) );
  INV_X1 U8391 ( .A(n6709), .ZN(n6712) );
  AOI22_X1 U8392 ( .A1(n7421), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n9100), .ZN(n6710) );
  OAI21_X1 U8393 ( .B1(n6712), .B2(n9103), .A(n6710), .ZN(P2_U3286) );
  AOI22_X1 U8394 ( .A1(n7087), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9781), .ZN(n6711) );
  OAI21_X1 U8395 ( .B1(n6712), .B2(n4336), .A(n6711), .ZN(P1_U3346) );
  INV_X1 U8396 ( .A(n8444), .ZN(n6713) );
  NAND2_X1 U8397 ( .A1(n9872), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6714) );
  OAI21_X1 U8398 ( .B1(n9872), .B2(n6715), .A(n6714), .ZN(P1_U3439) );
  INV_X1 U8399 ( .A(n6716), .ZN(n6760) );
  AOI22_X1 U8400 ( .A1(n7200), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9781), .ZN(n6717) );
  OAI21_X1 U8401 ( .B1(n6760), .B2(n4336), .A(n6717), .ZN(P1_U3345) );
  MUX2_X1 U8402 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8643), .Z(n6718) );
  AOI22_X1 U8403 ( .A1(n6806), .A2(n6805), .B1(n6718), .B2(n6807), .ZN(n9911)
         );
  MUX2_X1 U8404 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8643), .Z(n6719) );
  XNOR2_X1 U8405 ( .A(n6719), .B(n6739), .ZN(n9912) );
  INV_X1 U8406 ( .A(n6719), .ZN(n6720) );
  MUX2_X1 U8407 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8643), .Z(n6721) );
  XOR2_X1 U8408 ( .A(n9924), .B(n6721), .Z(n9931) );
  NOR2_X1 U8409 ( .A1(n6721), .A2(n6741), .ZN(n6723) );
  MUX2_X1 U8410 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8643), .Z(n7320) );
  XNOR2_X1 U8411 ( .A(n7320), .B(n7319), .ZN(n6722) );
  INV_X1 U8412 ( .A(n7318), .ZN(n6725) );
  OAI21_X1 U8413 ( .B1(n9929), .B2(n6723), .A(n6722), .ZN(n6724) );
  NAND3_X1 U8414 ( .A1(n6725), .A2(n9949), .A3(n6724), .ZN(n6754) );
  INV_X1 U8415 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10083) );
  AND2_X1 U8416 ( .A1(n6736), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6726) );
  OAI21_X1 U8417 ( .B1(n6807), .B2(n6726), .A(n6727), .ZN(n6808) );
  INV_X1 U8418 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7019) );
  NAND2_X1 U8419 ( .A1(n9904), .A2(n9903), .ZN(n9902) );
  NAND2_X1 U8420 ( .A1(n6739), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6728) );
  INV_X1 U8421 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9917) );
  XNOR2_X1 U8422 ( .A(n6744), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n6729) );
  INV_X1 U8423 ( .A(n6729), .ZN(n6731) );
  NAND3_X1 U8424 ( .A1(n6732), .A2(n6731), .A3(n6730), .ZN(n6733) );
  AND2_X1 U8425 ( .A1(n7308), .A2(n6733), .ZN(n6751) );
  NAND2_X1 U8426 ( .A1(n6735), .A2(n6734), .ZN(n9980) );
  INV_X1 U8427 ( .A(n9980), .ZN(n10009) );
  AND2_X1 U8428 ( .A1(n6736), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6737) );
  NAND2_X1 U8429 ( .A1(n6739), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6740) );
  OR2_X1 U8430 ( .A1(n6744), .A2(n7188), .ZN(n7336) );
  NAND2_X1 U8431 ( .A1(n6744), .A2(n7188), .ZN(n6745) );
  NAND2_X1 U8432 ( .A1(n7336), .A2(n6745), .ZN(n6747) );
  NAND2_X1 U8433 ( .A1(n6747), .A2(n6746), .ZN(n6748) );
  NAND2_X1 U8434 ( .A1(n7337), .A2(n6748), .ZN(n6749) );
  NAND2_X1 U8435 ( .A1(n10009), .A2(n6749), .ZN(n6750) );
  NAND2_X1 U8436 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7032) );
  OAI211_X1 U8437 ( .C1(n6751), .C2(n10005), .A(n6750), .B(n7032), .ZN(n6752)
         );
  AOI21_X1 U8438 ( .B1(n9962), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6752), .ZN(
        n6753) );
  OAI211_X1 U8439 ( .C1(n9958), .C2(n7319), .A(n6754), .B(n6753), .ZN(P2_U3186) );
  NAND2_X1 U8440 ( .A1(n4335), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6757) );
  NAND2_X1 U8441 ( .A1(n8176), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6756) );
  NAND2_X1 U8442 ( .A1(n8177), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6755) );
  INV_X1 U8443 ( .A(n9355), .ZN(n8362) );
  NAND2_X1 U8444 ( .A1(n8362), .A2(P1_U3973), .ZN(n6758) );
  OAI21_X1 U8445 ( .B1(P1_U3973), .B2(n5739), .A(n6758), .ZN(P1_U3585) );
  OAI222_X1 U8446 ( .A1(P2_U3151), .A2(n7745), .B1(n9103), .B2(n6760), .C1(
        n6759), .C2(n7434), .ZN(P2_U3285) );
  NAND2_X1 U8447 ( .A1(n6762), .A2(n6761), .ZN(n9827) );
  INV_X1 U8448 ( .A(n6937), .ZN(n6767) );
  INV_X1 U8449 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6766) );
  INV_X1 U8450 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6765) );
  XNOR2_X1 U8451 ( .A(n9299), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9305) );
  NAND2_X1 U8452 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6868) );
  INV_X1 U8453 ( .A(n6868), .ZN(n9304) );
  NAND2_X1 U8454 ( .A1(n9305), .A2(n9304), .ZN(n9303) );
  INV_X1 U8455 ( .A(n9299), .ZN(n9298) );
  NAND2_X1 U8456 ( .A1(n9298), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6764) );
  NAND2_X1 U8457 ( .A1(n9303), .A2(n6764), .ZN(n6872) );
  XNOR2_X1 U8458 ( .A(n6776), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9316) );
  OAI21_X1 U8459 ( .B1(n6766), .B2(n6776), .A(n9314), .ZN(n6941) );
  MUX2_X1 U8460 ( .A(n6116), .B(P1_REG2_REG_4__SCAN_IN), .S(n6937), .Z(n6942)
         );
  XNOR2_X1 U8461 ( .A(n6795), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n6768) );
  OR2_X1 U8462 ( .A1(n4337), .A2(n9817), .ZN(n8442) );
  AOI211_X1 U8463 ( .C1(n6769), .C2(n6768), .A(n6792), .B(n9343), .ZN(n6785)
         );
  INV_X1 U8464 ( .A(n6776), .ZN(n9313) );
  INV_X1 U8465 ( .A(n6876), .ZN(n6874) );
  INV_X1 U8466 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6770) );
  MUX2_X1 U8467 ( .A(n6770), .B(P1_REG1_REG_2__SCAN_IN), .S(n6876), .Z(n6775)
         );
  INV_X1 U8468 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6773) );
  MUX2_X1 U8469 ( .A(n6773), .B(P1_REG1_REG_1__SCAN_IN), .S(n9299), .Z(n6772)
         );
  AND2_X1 U8470 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6771) );
  NAND2_X1 U8471 ( .A1(n6772), .A2(n6771), .ZN(n9302) );
  OR2_X1 U8472 ( .A1(n9299), .A2(n6773), .ZN(n6877) );
  NAND2_X1 U8473 ( .A1(n9302), .A2(n6877), .ZN(n6774) );
  AND2_X1 U8474 ( .A1(n6775), .A2(n6774), .ZN(n6875) );
  AOI21_X1 U8475 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(n6874), .A(n6875), .ZN(
        n9311) );
  INV_X1 U8476 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6777) );
  MUX2_X1 U8477 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6777), .S(n6776), .Z(n9310)
         );
  NOR2_X1 U8478 ( .A1(n9311), .A2(n9310), .ZN(n9309) );
  AOI21_X1 U8479 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n9313), .A(n9309), .ZN(
        n6939) );
  INV_X1 U8480 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6778) );
  MUX2_X1 U8481 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6778), .S(n6937), .Z(n6938)
         );
  OAI22_X1 U8482 ( .A1(n6939), .A2(n6938), .B1(n6778), .B2(n6937), .ZN(n6780)
         );
  INV_X1 U8483 ( .A(n6780), .ZN(n6783) );
  INV_X1 U8484 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7251) );
  MUX2_X1 U8485 ( .A(n7251), .B(P1_REG1_REG_5__SCAN_IN), .S(n6795), .Z(n6782)
         );
  MUX2_X1 U8486 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n7251), .S(n6795), .Z(n6779)
         );
  NAND2_X1 U8487 ( .A1(n6780), .A2(n6779), .ZN(n6798) );
  INV_X1 U8488 ( .A(n6798), .ZN(n6781) );
  INV_X1 U8489 ( .A(n9817), .ZN(n8181) );
  AOI211_X1 U8490 ( .C1(n6783), .C2(n6782), .A(n6781), .B(n9849), .ZN(n6784)
         );
  NOR2_X1 U8491 ( .A1(n6785), .A2(n6784), .ZN(n6788) );
  NAND2_X1 U8492 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n7301) );
  INV_X1 U8493 ( .A(n7301), .ZN(n6786) );
  AOI21_X1 U8494 ( .B1(n9824), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n6786), .ZN(
        n6787) );
  OAI211_X1 U8495 ( .C1(n6789), .C2(n9847), .A(n6788), .B(n6787), .ZN(P1_U3248) );
  NAND2_X1 U8496 ( .A1(n7518), .A2(P1_U3973), .ZN(n6790) );
  OAI21_X1 U8497 ( .B1(P1_U3973), .B2(n6791), .A(n6790), .ZN(P1_U3561) );
  AOI21_X1 U8498 ( .B1(n6795), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6792), .ZN(
        n6794) );
  XNOR2_X1 U8499 ( .A(n6828), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n6793) );
  NOR2_X1 U8500 ( .A1(n6794), .A2(n6793), .ZN(n6827) );
  AOI211_X1 U8501 ( .C1(n6794), .C2(n6793), .A(n9343), .B(n6827), .ZN(n6801)
         );
  NAND2_X1 U8502 ( .A1(n6795), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6797) );
  INV_X1 U8503 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9891) );
  MUX2_X1 U8504 ( .A(n9891), .B(P1_REG1_REG_6__SCAN_IN), .S(n6828), .Z(n6796)
         );
  AOI21_X1 U8505 ( .B1(n6798), .B2(n6797), .A(n6796), .ZN(n6856) );
  AND3_X1 U8506 ( .A1(n6798), .A2(n6797), .A3(n6796), .ZN(n6799) );
  NOR3_X1 U8507 ( .A1(n9849), .A2(n6856), .A3(n6799), .ZN(n6800) );
  NOR2_X1 U8508 ( .A1(n6801), .A2(n6800), .ZN(n6804) );
  AND2_X1 U8509 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6802) );
  AOI21_X1 U8510 ( .B1(n9824), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n6802), .ZN(
        n6803) );
  OAI211_X1 U8511 ( .C1(n6833), .C2(n9847), .A(n6804), .B(n6803), .ZN(P1_U3249) );
  INV_X1 U8512 ( .A(n9949), .ZN(n10013) );
  XNOR2_X1 U8513 ( .A(n6806), .B(n6805), .ZN(n6821) );
  NOR2_X1 U8514 ( .A1(n9958), .A2(n6807), .ZN(n6819) );
  INV_X1 U8515 ( .A(n10005), .ZN(n9906) );
  NAND2_X1 U8516 ( .A1(n6808), .A2(n7019), .ZN(n6809) );
  NAND2_X1 U8517 ( .A1(n6810), .A2(n6809), .ZN(n6811) );
  NAND2_X1 U8518 ( .A1(n9906), .A2(n6811), .ZN(n6816) );
  NAND2_X1 U8519 ( .A1(n6813), .A2(n6812), .ZN(n6814) );
  NAND2_X1 U8520 ( .A1(n10009), .A2(n6814), .ZN(n6815) );
  OAI211_X1 U8521 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6817), .A(n6816), .B(n6815), .ZN(n6818) );
  AOI211_X1 U8522 ( .C1(n9962), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n6819), .B(
        n6818), .ZN(n6820) );
  OAI21_X1 U8523 ( .B1(n10013), .B2(n6821), .A(n6820), .ZN(P2_U3183) );
  INV_X1 U8524 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6823) );
  INV_X1 U8525 ( .A(n6822), .ZN(n6825) );
  INV_X1 U8526 ( .A(n7465), .ZN(n7453) );
  OAI222_X1 U8527 ( .A1(n9789), .A2(n6823), .B1(n4336), .B2(n6825), .C1(
        P1_U3086), .C2(n7453), .ZN(P1_U3344) );
  INV_X1 U8528 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6824) );
  OAI222_X1 U8529 ( .A1(n7845), .A2(P2_U3151), .B1(n8046), .B2(n6825), .C1(
        n6824), .C2(n7434), .ZN(P2_U3284) );
  INV_X1 U8530 ( .A(n7466), .ZN(n9834) );
  INV_X1 U8531 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6826) );
  OAI222_X1 U8532 ( .A1(n4336), .A2(n6846), .B1(n9834), .B2(P1_U3086), .C1(
        n6826), .C2(n9789), .ZN(P1_U3343) );
  INV_X1 U8533 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6829) );
  MUX2_X1 U8534 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n6829), .S(n6851), .Z(n6830)
         );
  INV_X1 U8535 ( .A(n6830), .ZN(n6848) );
  XNOR2_X1 U8536 ( .A(n6960), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n6831) );
  AOI211_X1 U8537 ( .C1(n6832), .C2(n6831), .A(n9343), .B(n6954), .ZN(n6844)
         );
  NOR2_X1 U8538 ( .A1(n6833), .A2(n9891), .ZN(n6850) );
  INV_X1 U8539 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6834) );
  MUX2_X1 U8540 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6834), .S(n6851), .Z(n6835)
         );
  OAI21_X1 U8541 ( .B1(n6856), .B2(n6850), .A(n6835), .ZN(n6854) );
  NAND2_X1 U8542 ( .A1(n6851), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6837) );
  INV_X1 U8543 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9894) );
  MUX2_X1 U8544 ( .A(n9894), .B(P1_REG1_REG_8__SCAN_IN), .S(n6960), .Z(n6836)
         );
  AOI21_X1 U8545 ( .B1(n6854), .B2(n6837), .A(n6836), .ZN(n6959) );
  AND3_X1 U8546 ( .A1(n6854), .A2(n6837), .A3(n6836), .ZN(n6838) );
  NOR3_X1 U8547 ( .A1(n6959), .A2(n6838), .A3(n9849), .ZN(n6843) );
  INV_X1 U8548 ( .A(n6960), .ZN(n6841) );
  AND2_X1 U8549 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6839) );
  AOI21_X1 U8550 ( .B1(n9824), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n6839), .ZN(
        n6840) );
  OAI21_X1 U8551 ( .B1(n6841), .B2(n9847), .A(n6840), .ZN(n6842) );
  OR3_X1 U8552 ( .A1(n6844), .A2(n6843), .A3(n6842), .ZN(P1_U3251) );
  INV_X1 U8553 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6845) );
  OAI222_X1 U8554 ( .A1(P2_U3151), .A2(n7949), .B1(n8046), .B2(n6846), .C1(
        n6845), .C2(n7434), .ZN(P2_U3283) );
  AOI211_X1 U8555 ( .C1(n6849), .C2(n6848), .A(n9343), .B(n6847), .ZN(n6863)
         );
  INV_X1 U8556 ( .A(n6850), .ZN(n6853) );
  MUX2_X1 U8557 ( .A(n6834), .B(P1_REG1_REG_7__SCAN_IN), .S(n6851), .Z(n6852)
         );
  NAND2_X1 U8558 ( .A1(n6853), .A2(n6852), .ZN(n6855) );
  INV_X1 U8559 ( .A(n9849), .ZN(n9340) );
  OAI211_X1 U8560 ( .C1(n6856), .C2(n6855), .A(n6854), .B(n9340), .ZN(n6860)
         );
  NOR2_X1 U8561 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6857), .ZN(n6858) );
  AOI21_X1 U8562 ( .B1(n9824), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n6858), .ZN(
        n6859) );
  OAI211_X1 U8563 ( .C1(n9847), .C2(n6861), .A(n6860), .B(n6859), .ZN(n6862)
         );
  OR2_X1 U8564 ( .A1(n6863), .A2(n6862), .ZN(P1_U3250) );
  OAI21_X1 U8565 ( .B1(n6866), .B2(n6865), .A(n6864), .ZN(n7042) );
  NOR2_X1 U8566 ( .A1(n4337), .A2(n8181), .ZN(n6870) );
  NOR2_X1 U8567 ( .A1(n9817), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6867) );
  OR2_X1 U8568 ( .A1(n6867), .A2(n4337), .ZN(n9815) );
  INV_X1 U8569 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9819) );
  NAND2_X1 U8570 ( .A1(n9815), .A2(n9819), .ZN(n9822) );
  OAI211_X1 U8571 ( .C1(n6868), .C2(n8442), .A(P1_U3973), .B(n9822), .ZN(n6869) );
  AOI21_X1 U8572 ( .B1(n7042), .B2(n6870), .A(n6869), .ZN(n6947) );
  OAI211_X1 U8573 ( .C1(n6873), .C2(n6872), .A(n9853), .B(n6871), .ZN(n6884)
         );
  AOI22_X1 U8574 ( .A1(n9824), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6883) );
  INV_X1 U8575 ( .A(n9847), .ZN(n9332) );
  NAND2_X1 U8576 ( .A1(n9332), .A2(n6874), .ZN(n6882) );
  INV_X1 U8577 ( .A(n6875), .ZN(n6880) );
  MUX2_X1 U8578 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6770), .S(n6876), .Z(n6878)
         );
  NAND3_X1 U8579 ( .A1(n6878), .A2(n9302), .A3(n6877), .ZN(n6879) );
  NAND3_X1 U8580 ( .A1(n9340), .A2(n6880), .A3(n6879), .ZN(n6881) );
  NAND4_X1 U8581 ( .A1(n6884), .A2(n6883), .A3(n6882), .A4(n6881), .ZN(n6885)
         );
  OR2_X1 U8582 ( .A1(n6947), .A2(n6885), .ZN(P1_U3245) );
  OAI21_X1 U8583 ( .B1(n6886), .B2(P1_D_REG_1__SCAN_IN), .A(n9776), .ZN(n6893)
         );
  OR2_X1 U8584 ( .A1(n8444), .A2(n6887), .ZN(n7153) );
  NOR2_X1 U8585 ( .A1(n7153), .A2(n6888), .ZN(n6892) );
  NAND2_X1 U8586 ( .A1(n6890), .A2(n6889), .ZN(n6891) );
  INV_X1 U8587 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9816) );
  INV_X1 U8588 ( .A(n8387), .ZN(n7164) );
  NAND2_X1 U8589 ( .A1(n6894), .A2(n8437), .ZN(n8443) );
  INV_X1 U8590 ( .A(n8437), .ZN(n6895) );
  NAND2_X1 U8591 ( .A1(n6896), .A2(n6895), .ZN(n6897) );
  AND2_X1 U8592 ( .A1(n6897), .A2(n7163), .ZN(n6898) );
  NAND2_X1 U8593 ( .A1(n8443), .A2(n6898), .ZN(n7781) );
  INV_X1 U8594 ( .A(n8193), .ZN(n8445) );
  OR2_X1 U8595 ( .A1(n8445), .A2(n7162), .ZN(n7116) );
  OR2_X1 U8596 ( .A1(n8193), .A2(n6047), .ZN(n6900) );
  INV_X1 U8597 ( .A(n8338), .ZN(n8389) );
  NAND2_X1 U8598 ( .A1(n8389), .A2(n6899), .ZN(n8382) );
  NAND2_X1 U8599 ( .A1(n6901), .A2(n8387), .ZN(n7118) );
  OAI21_X1 U8600 ( .B1(n6901), .B2(n8387), .A(n7118), .ZN(n8305) );
  INV_X1 U8601 ( .A(n8305), .ZN(n7158) );
  OAI21_X1 U8602 ( .B1(n9878), .B2(n9608), .A(n7158), .ZN(n6902) );
  NAND2_X1 U8603 ( .A1(n7140), .A2(n9524), .ZN(n7159) );
  OAI211_X1 U8604 ( .C1(n7163), .C2(n7164), .A(n6902), .B(n7159), .ZN(n6906)
         );
  NAND2_X1 U8605 ( .A1(n6906), .A2(n9896), .ZN(n6903) );
  OAI21_X1 U8606 ( .B1(n9896), .B2(n9816), .A(n6903), .ZN(P1_U3522) );
  INV_X1 U8607 ( .A(n7156), .ZN(n6905) );
  INV_X1 U8608 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6908) );
  NAND2_X1 U8609 ( .A1(n6906), .A2(n9890), .ZN(n6907) );
  OAI21_X1 U8610 ( .B1(n9890), .B2(n6908), .A(n6907), .ZN(P1_U3453) );
  OR2_X1 U8611 ( .A1(n6915), .A2(n6909), .ZN(n6912) );
  OR2_X1 U8612 ( .A1(n6910), .A2(n6927), .ZN(n6911) );
  AND2_X2 U8613 ( .A1(n6912), .A2(n6911), .ZN(n8610) );
  AND2_X1 U8614 ( .A1(n6931), .A2(n6929), .ZN(n6977) );
  INV_X1 U8615 ( .A(n6977), .ZN(n6914) );
  OR2_X1 U8616 ( .A1(n6915), .A2(n10052), .ZN(n6919) );
  INV_X1 U8617 ( .A(n6916), .ZN(n6917) );
  AOI22_X1 U8618 ( .A1(n6913), .A2(n8571), .B1(n7065), .B2(n8615), .ZN(n6935)
         );
  OR2_X1 U8619 ( .A1(n6921), .A2(n6920), .ZN(n6926) );
  AND3_X1 U8620 ( .A1(n6924), .A2(n6923), .A3(n6922), .ZN(n6925) );
  OAI211_X1 U8621 ( .C1(n6931), .C2(n6927), .A(n6926), .B(n6925), .ZN(n6928)
         );
  NAND2_X1 U8622 ( .A1(n6928), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6933) );
  INV_X1 U8623 ( .A(n6929), .ZN(n6930) );
  OR2_X1 U8624 ( .A1(n6931), .A2(n6930), .ZN(n6932) );
  NAND2_X1 U8625 ( .A1(n8608), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6991) );
  NAND2_X1 U8626 ( .A1(n6991), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6934) );
  OAI211_X1 U8627 ( .C1(n7054), .C2(n8610), .A(n6935), .B(n6934), .ZN(P2_U3172) );
  NAND2_X1 U8628 ( .A1(n9824), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n6936) );
  NAND2_X1 U8629 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7288) );
  OAI211_X1 U8630 ( .C1(n9847), .C2(n6937), .A(n6936), .B(n7288), .ZN(n6946)
         );
  XNOR2_X1 U8631 ( .A(n6939), .B(n6938), .ZN(n6944) );
  OAI211_X1 U8632 ( .C1(n6942), .C2(n6941), .A(n9853), .B(n6940), .ZN(n6943)
         );
  OAI21_X1 U8633 ( .B1(n9849), .B2(n6944), .A(n6943), .ZN(n6945) );
  OR3_X1 U8634 ( .A1(n6947), .A2(n6946), .A3(n6945), .ZN(P1_U3247) );
  INV_X1 U8635 ( .A(n7054), .ZN(n6948) );
  OAI21_X1 U8636 ( .B1(n8952), .B2(n10075), .A(n6948), .ZN(n6950) );
  NOR2_X1 U8637 ( .A1(n10027), .A2(n10030), .ZN(n7055) );
  INV_X1 U8638 ( .A(n7055), .ZN(n6949) );
  OAI211_X1 U8639 ( .C1(n6974), .C2(n10052), .A(n6950), .B(n6949), .ZN(n6952)
         );
  NAND2_X1 U8640 ( .A1(n6952), .A2(n10096), .ZN(n6951) );
  OAI21_X1 U8641 ( .B1(n10096), .B2(n6704), .A(n6951), .ZN(P2_U3459) );
  NAND2_X1 U8642 ( .A1(n6952), .A2(n10081), .ZN(n6953) );
  OAI21_X1 U8643 ( .B1(n5257), .B2(n10081), .A(n6953), .ZN(P2_U3390) );
  XOR2_X1 U8644 ( .A(n7087), .B(P1_REG2_REG_9__SCAN_IN), .Z(n6956) );
  OAI21_X1 U8645 ( .B1(n6956), .B2(n6955), .A(n7083), .ZN(n6957) );
  NAND2_X1 U8646 ( .A1(n6957), .A2(n9853), .ZN(n6968) );
  INV_X1 U8647 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6958) );
  MUX2_X1 U8648 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n6958), .S(n7087), .Z(n6962)
         );
  AOI21_X1 U8649 ( .B1(n6960), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6959), .ZN(
        n6961) );
  NAND2_X1 U8650 ( .A1(n6961), .A2(n6962), .ZN(n7086) );
  OAI21_X1 U8651 ( .B1(n6962), .B2(n6961), .A(n7086), .ZN(n6966) );
  INV_X1 U8652 ( .A(n7087), .ZN(n6964) );
  NAND2_X1 U8653 ( .A1(n9824), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n6963) );
  NAND2_X1 U8654 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7758) );
  OAI211_X1 U8655 ( .C1(n9847), .C2(n6964), .A(n6963), .B(n7758), .ZN(n6965)
         );
  AOI21_X1 U8656 ( .B1(n6966), .B2(n9340), .A(n6965), .ZN(n6967) );
  NAND2_X1 U8657 ( .A1(n6968), .A2(n6967), .ZN(P1_U3252) );
  NAND2_X1 U8658 ( .A1(n8491), .A2(n6974), .ZN(n6975) );
  NAND2_X1 U8659 ( .A1(n7016), .A2(n6975), .ZN(n6983) );
  XOR2_X1 U8660 ( .A(n6982), .B(n6983), .Z(n6981) );
  AOI22_X1 U8661 ( .A1(n8635), .A2(n8571), .B1(n8606), .B2(n5697), .ZN(n6978)
         );
  OAI21_X1 U8662 ( .B1(n8596), .B2(n7020), .A(n6978), .ZN(n6979) );
  AOI21_X1 U8663 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n6991), .A(n6979), .ZN(
        n6980) );
  OAI21_X1 U8664 ( .B1(n6981), .B2(n8610), .A(n6980), .ZN(P2_U3162) );
  INV_X1 U8665 ( .A(n6984), .ZN(n6985) );
  NAND2_X1 U8666 ( .A1(n6985), .A2(n10027), .ZN(n6986) );
  XNOR2_X1 U8667 ( .A(n6998), .B(n7074), .ZN(n6996) );
  XOR2_X1 U8668 ( .A(n6997), .B(n6996), .Z(n6993) );
  AOI22_X1 U8669 ( .A1(n6913), .A2(n8606), .B1(n8571), .B2(n8634), .ZN(n6989)
         );
  OAI21_X1 U8670 ( .B1(n10035), .B2(n8596), .A(n6989), .ZN(n6990) );
  AOI21_X1 U8671 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n6991), .A(n6990), .ZN(
        n6992) );
  OAI21_X1 U8672 ( .B1(n6993), .B2(n8610), .A(n6992), .ZN(P2_U3177) );
  INV_X1 U8673 ( .A(n6994), .ZN(n7013) );
  INV_X1 U8674 ( .A(n7717), .ZN(n7711) );
  INV_X1 U8675 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6995) );
  OAI222_X1 U8676 ( .A1(n4336), .A2(n7013), .B1(n7711), .B2(P1_U3086), .C1(
        n6995), .C2(n9789), .ZN(P1_U3342) );
  NAND2_X1 U8677 ( .A1(n6997), .A2(n6996), .ZN(n7001) );
  INV_X1 U8678 ( .A(n6998), .ZN(n6999) );
  NAND2_X1 U8679 ( .A1(n6999), .A2(n7074), .ZN(n7000) );
  XNOR2_X1 U8680 ( .A(n4329), .B(n7077), .ZN(n7023) );
  XNOR2_X1 U8681 ( .A(n7023), .B(n10029), .ZN(n7003) );
  AOI21_X1 U8682 ( .B1(n7002), .B2(n7003), .A(n8610), .ZN(n7006) );
  INV_X1 U8683 ( .A(n7002), .ZN(n7005) );
  INV_X1 U8684 ( .A(n7003), .ZN(n7004) );
  NAND2_X1 U8685 ( .A1(n7006), .A2(n7026), .ZN(n7011) );
  NAND2_X1 U8686 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9921) );
  NAND2_X1 U8687 ( .A1(n8633), .A2(n8571), .ZN(n7007) );
  OAI211_X1 U8688 ( .C1(n7074), .C2(n8574), .A(n9921), .B(n7007), .ZN(n7009)
         );
  NOR2_X1 U8689 ( .A1(n8608), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7008) );
  AOI211_X1 U8690 ( .C1(n7077), .C2(n8615), .A(n7009), .B(n7008), .ZN(n7010)
         );
  NAND2_X1 U8691 ( .A1(n7011), .A2(n7010), .ZN(P2_U3158) );
  INV_X1 U8692 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7012) );
  OAI222_X1 U8693 ( .A1(P2_U3151), .A2(n7950), .B1(n9103), .B2(n7013), .C1(
        n7012), .C2(n7434), .ZN(P2_U3282) );
  INV_X1 U8694 ( .A(n7014), .ZN(n7015) );
  AOI21_X1 U8695 ( .B1(n7016), .B2(n5770), .A(n7015), .ZN(n7104) );
  XNOR2_X1 U8696 ( .A(n5770), .B(n7017), .ZN(n7018) );
  AOI222_X1 U8697 ( .A1(n8952), .A2(n7018), .B1(n5697), .B2(n5656), .C1(n8635), 
        .C2(n8949), .ZN(n7099) );
  OAI21_X1 U8698 ( .B1(n10068), .B2(n7104), .A(n7099), .ZN(n7080) );
  OAI22_X1 U8699 ( .A1(n9001), .A2(n7020), .B1(n10096), .B2(n7019), .ZN(n7021)
         );
  AOI21_X1 U8700 ( .B1(n7080), .B2(n10096), .A(n7021), .ZN(n7022) );
  INV_X1 U8701 ( .A(n7022), .ZN(P2_U3460) );
  XNOR2_X1 U8702 ( .A(n7105), .B(n7110), .ZN(n7030) );
  INV_X1 U8703 ( .A(n7023), .ZN(n7024) );
  NAND2_X1 U8704 ( .A1(n7024), .A2(n8634), .ZN(n7025) );
  INV_X1 U8705 ( .A(n7030), .ZN(n7027) );
  INV_X1 U8706 ( .A(n7107), .ZN(n7028) );
  AOI21_X1 U8707 ( .B1(n7030), .B2(n7029), .A(n7028), .ZN(n7038) );
  INV_X1 U8708 ( .A(n8608), .ZN(n8593) );
  INV_X1 U8709 ( .A(n7031), .ZN(n7189) );
  NAND2_X1 U8710 ( .A1(n8615), .A2(n7190), .ZN(n7035) );
  NAND2_X1 U8711 ( .A1(n8632), .A2(n8571), .ZN(n7034) );
  NAND2_X1 U8712 ( .A1(n8634), .A2(n8606), .ZN(n7033) );
  NAND4_X1 U8713 ( .A1(n7035), .A2(n7034), .A3(n7033), .A4(n7032), .ZN(n7036)
         );
  AOI21_X1 U8714 ( .B1(n8593), .B2(n7189), .A(n7036), .ZN(n7037) );
  OAI21_X1 U8715 ( .B1(n7038), .B2(n8610), .A(n7037), .ZN(P2_U3170) );
  AOI22_X1 U8716 ( .A1(n6649), .A2(n8387), .B1(n9802), .B2(n7140), .ZN(n7041)
         );
  OR2_X1 U8717 ( .A1(n7039), .A2(n8444), .ZN(n9149) );
  NAND2_X1 U8718 ( .A1(n9149), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7040) );
  OAI211_X1 U8719 ( .C1(n9245), .C2(n7042), .A(n7041), .B(n7040), .ZN(P1_U3232) );
  INV_X1 U8720 ( .A(n7043), .ZN(n7044) );
  INV_X1 U8721 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10161) );
  OAI222_X1 U8722 ( .A1(n8681), .A2(P2_U3151), .B1(n8046), .B2(n7044), .C1(
        n10161), .C2(n7434), .ZN(P2_U3281) );
  INV_X1 U8723 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7045) );
  INV_X1 U8724 ( .A(n7963), .ZN(n7958) );
  OAI222_X1 U8725 ( .A1(n9789), .A2(n7045), .B1(n4336), .B2(n7044), .C1(
        P1_U3086), .C2(n7958), .ZN(P1_U3341) );
  XNOR2_X1 U8726 ( .A(n7046), .B(n7047), .ZN(n7048) );
  NAND2_X1 U8727 ( .A1(n7048), .A2(n9809), .ZN(n7052) );
  NAND2_X1 U8728 ( .A1(n7140), .A2(n9523), .ZN(n7050) );
  NAND2_X1 U8729 ( .A1(n9292), .A2(n9524), .ZN(n7049) );
  NAND2_X1 U8730 ( .A1(n7050), .A2(n7049), .ZN(n7143) );
  AOI22_X1 U8731 ( .A1(n9254), .A2(n7143), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n9149), .ZN(n7051) );
  OAI211_X1 U8732 ( .C1(n7247), .C2(n9800), .A(n7052), .B(n7051), .ZN(P1_U3237) );
  NOR3_X1 U8733 ( .A1(n7054), .A2(n10080), .A3(n7053), .ZN(n7056) );
  NOR2_X1 U8734 ( .A1(n7056), .A2(n7055), .ZN(n7062) );
  INV_X1 U8735 ( .A(n7057), .ZN(n7059) );
  OAI211_X1 U8736 ( .C1(n7061), .C2(n7060), .A(n7059), .B(n7058), .ZN(n7064)
         );
  MUX2_X1 U8737 ( .A(n7063), .B(n7062), .S(n8926), .Z(n7067) );
  OR2_X1 U8738 ( .A1(n7064), .A2(n10023), .ZN(n8912) );
  NAND2_X1 U8739 ( .A1(n8956), .A2(n7065), .ZN(n7066) );
  OAI211_X1 U8740 ( .C1(n10021), .C2(n7068), .A(n7067), .B(n7066), .ZN(
        P2_U3233) );
  OAI21_X1 U8741 ( .B1(n7070), .B2(n7071), .A(n7069), .ZN(n7228) );
  XNOR2_X1 U8742 ( .A(n7072), .B(n7071), .ZN(n7073) );
  OAI222_X1 U8743 ( .A1(n10030), .A2(n7110), .B1(n10028), .B2(n7074), .C1(
        n10026), .C2(n7073), .ZN(n7225) );
  AOI21_X1 U8744 ( .B1(n10075), .B2(n7228), .A(n7225), .ZN(n7079) );
  OAI22_X1 U8745 ( .A1(n9070), .A2(n7224), .B1(n5281), .B2(n10081), .ZN(n7075)
         );
  INV_X1 U8746 ( .A(n7075), .ZN(n7076) );
  OAI21_X1 U8747 ( .B1(n7079), .B2(n10082), .A(n7076), .ZN(P2_U3399) );
  AOI22_X1 U8748 ( .A1(n9006), .A2(n7077), .B1(n10094), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n7078) );
  OAI21_X1 U8749 ( .B1(n7079), .B2(n10094), .A(n7078), .ZN(P2_U3462) );
  INV_X1 U8750 ( .A(n7080), .ZN(n7082) );
  AOI22_X1 U8751 ( .A1(n9079), .A2(n7101), .B1(n10082), .B2(
        P2_REG0_REG_1__SCAN_IN), .ZN(n7081) );
  OAI21_X1 U8752 ( .B1(n7082), .B2(n10082), .A(n7081), .ZN(P2_U3393) );
  XNOR2_X1 U8753 ( .A(n7200), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n7085) );
  AOI211_X1 U8754 ( .C1(n7085), .C2(n7084), .A(n9343), .B(n7194), .ZN(n7096)
         );
  OAI21_X1 U8755 ( .B1(n7087), .B2(P1_REG1_REG_9__SCAN_IN), .A(n7086), .ZN(
        n7090) );
  INV_X1 U8756 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7088) );
  MUX2_X1 U8757 ( .A(n7088), .B(P1_REG1_REG_10__SCAN_IN), .S(n7200), .Z(n7089)
         );
  NOR2_X1 U8758 ( .A1(n7090), .A2(n7089), .ZN(n7199) );
  AOI211_X1 U8759 ( .C1(n7090), .C2(n7089), .A(n9849), .B(n7199), .ZN(n7095)
         );
  INV_X1 U8760 ( .A(n7200), .ZN(n7093) );
  AND2_X1 U8761 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7091) );
  AOI21_X1 U8762 ( .B1(n9824), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n7091), .ZN(
        n7092) );
  OAI21_X1 U8763 ( .B1(n7093), .B2(n9847), .A(n7092), .ZN(n7094) );
  OR3_X1 U8764 ( .A1(n7096), .A2(n7095), .A3(n7094), .ZN(P1_U3253) );
  AND2_X1 U8765 ( .A1(n7097), .A2(n7695), .ZN(n7615) );
  INV_X1 U8766 ( .A(n7615), .ZN(n7098) );
  NAND2_X1 U8767 ( .A1(n10051), .A2(n7098), .ZN(n10032) );
  MUX2_X1 U8768 ( .A(n7100), .B(n7099), .S(n8926), .Z(n7103) );
  AOI22_X1 U8769 ( .A1(n8956), .A2(n7101), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8955), .ZN(n7102) );
  OAI211_X1 U8770 ( .C1(n7104), .C2(n8959), .A(n7103), .B(n7102), .ZN(P2_U3232) );
  XNOR2_X1 U8771 ( .A(n4329), .B(n7397), .ZN(n7170) );
  XNOR2_X1 U8772 ( .A(n7170), .B(n8632), .ZN(n7171) );
  NAND2_X1 U8773 ( .A1(n7105), .A2(n7110), .ZN(n7106) );
  XOR2_X1 U8774 ( .A(n7172), .B(n7171), .Z(n7115) );
  INV_X1 U8775 ( .A(n7108), .ZN(n7396) );
  NOR2_X1 U8776 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7109), .ZN(n9938) );
  NOR2_X1 U8777 ( .A1(n7110), .A2(n8574), .ZN(n7111) );
  AOI211_X1 U8778 ( .C1(n8571), .C2(n8631), .A(n9938), .B(n7111), .ZN(n7112)
         );
  OAI21_X1 U8779 ( .B1(n10043), .B2(n8596), .A(n7112), .ZN(n7113) );
  AOI21_X1 U8780 ( .B1(n7396), .B2(n8593), .A(n7113), .ZN(n7114) );
  OAI21_X1 U8781 ( .B1(n7115), .B2(n8610), .A(n7114), .ZN(P2_U3167) );
  INV_X1 U8782 ( .A(n7116), .ZN(n9884) );
  NAND2_X1 U8783 ( .A1(n7118), .A2(n7117), .ZN(n7148) );
  OAI21_X1 U8784 ( .B1(n7117), .B2(n7118), .A(n7148), .ZN(n7126) );
  INV_X1 U8785 ( .A(n7163), .ZN(n7119) );
  INV_X1 U8786 ( .A(n7145), .ZN(n7120) );
  AOI211_X1 U8787 ( .C1(n8387), .C2(n4511), .A(n9595), .B(n7120), .ZN(n7638)
         );
  INV_X1 U8788 ( .A(n7126), .ZN(n7642) );
  NOR2_X1 U8789 ( .A1(n6901), .A2(n7164), .ZN(n7121) );
  OAI21_X1 U8790 ( .B1(n7122), .B2(n7121), .A(n7142), .ZN(n7124) );
  INV_X1 U8791 ( .A(n6901), .ZN(n8388) );
  INV_X1 U8792 ( .A(n9293), .ZN(n7215) );
  OAI22_X1 U8793 ( .A1(n8388), .A2(n9488), .B1(n7215), .B2(n9490), .ZN(n7123)
         );
  AOI21_X1 U8794 ( .B1(n7124), .B2(n9608), .A(n7123), .ZN(n7125) );
  OAI21_X1 U8795 ( .B1(n7642), .B2(n7781), .A(n7125), .ZN(n7639) );
  AOI211_X1 U8796 ( .C1(n9884), .C2(n7126), .A(n7638), .B(n7639), .ZN(n7139)
         );
  AOI22_X1 U8797 ( .A1(n9695), .A2(n4511), .B1(n9893), .B2(
        P1_REG1_REG_1__SCAN_IN), .ZN(n7127) );
  OAI21_X1 U8798 ( .B1(n7139), .B2(n9893), .A(n7127), .ZN(P1_U3523) );
  NAND2_X1 U8799 ( .A1(n7129), .A2(n7128), .ZN(n7130) );
  XOR2_X1 U8800 ( .A(n7131), .B(n7130), .Z(n7134) );
  INV_X1 U8801 ( .A(n9291), .ZN(n7303) );
  OAI22_X1 U8802 ( .A1(n7303), .A2(n9490), .B1(n7215), .B2(n9488), .ZN(n7236)
         );
  AOI22_X1 U8803 ( .A1(n6649), .A2(n7242), .B1(n9254), .B2(n7236), .ZN(n7133)
         );
  MUX2_X1 U8804 ( .A(P1_STATE_REG_SCAN_IN), .B(n9814), .S(n9860), .Z(n7132) );
  OAI211_X1 U8805 ( .C1(n7134), .C2(n9245), .A(n7133), .B(n7132), .ZN(P1_U3218) );
  INV_X1 U8806 ( .A(n9769), .ZN(n9759) );
  INV_X1 U8807 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7136) );
  OAI22_X1 U8808 ( .A1(n9759), .A2(n7636), .B1(n9890), .B2(n7136), .ZN(n7137)
         );
  INV_X1 U8809 ( .A(n7137), .ZN(n7138) );
  OAI21_X1 U8810 ( .B1(n7139), .B2(n9888), .A(n7138), .ZN(P1_U3456) );
  INV_X1 U8811 ( .A(n7140), .ZN(n8391) );
  NAND2_X1 U8812 ( .A1(n8391), .A2(n4511), .ZN(n7141) );
  XOR2_X1 U8813 ( .A(n8308), .B(n7207), .Z(n7144) );
  AOI21_X1 U8814 ( .B1(n7144), .B2(n9608), .A(n7143), .ZN(n7492) );
  INV_X1 U8815 ( .A(n7213), .ZN(n7233) );
  AOI21_X1 U8816 ( .B1(n7485), .B2(n7145), .A(n9595), .ZN(n7146) );
  NAND2_X1 U8817 ( .A1(n7233), .A2(n7146), .ZN(n7488) );
  AND2_X1 U8818 ( .A1(n7492), .A2(n7488), .ZN(n7250) );
  INV_X1 U8819 ( .A(n9774), .ZN(n7869) );
  NAND2_X1 U8820 ( .A1(n8391), .A2(n7636), .ZN(n7147) );
  NAND2_X1 U8821 ( .A1(n7148), .A2(n7147), .ZN(n7149) );
  OAI21_X1 U8822 ( .B1(n7149), .B2(n8308), .A(n7217), .ZN(n7490) );
  INV_X1 U8823 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7150) );
  OAI22_X1 U8824 ( .A1(n9759), .A2(n7247), .B1(n9890), .B2(n7150), .ZN(n7151)
         );
  AOI21_X1 U8825 ( .B1(n7869), .B2(n7490), .A(n7151), .ZN(n7152) );
  OAI21_X1 U8826 ( .B1(n7250), .B2(n9888), .A(n7152), .ZN(P1_U3459) );
  INV_X1 U8827 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7169) );
  INV_X1 U8828 ( .A(n7153), .ZN(n7154) );
  NAND2_X1 U8829 ( .A1(n7155), .A2(n7154), .ZN(n7157) );
  INV_X2 U8830 ( .A(n9617), .ZN(n9623) );
  INV_X1 U8831 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7161) );
  NAND3_X1 U8832 ( .A1(n7158), .A2(n8443), .A3(n7163), .ZN(n7160) );
  OAI211_X1 U8833 ( .C1(n9544), .C2(n7161), .A(n7160), .B(n7159), .ZN(n7167)
         );
  INV_X1 U8834 ( .A(n7162), .ZN(n8438) );
  NOR4_X1 U8835 ( .A1(n7165), .A2(n8438), .A3(n7164), .A4(n7163), .ZN(n7166)
         );
  AOI21_X1 U8836 ( .B1(n9623), .B2(n7167), .A(n7166), .ZN(n7168) );
  OAI21_X1 U8837 ( .B1(n7169), .B2(n9623), .A(n7168), .ZN(P1_U3293) );
  INV_X1 U8838 ( .A(n8610), .ZN(n8588) );
  OAI211_X1 U8839 ( .C1(n7174), .C2(n7173), .A(n7258), .B(n8588), .ZN(n7179)
         );
  NAND2_X1 U8840 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3151), .ZN(n9974) );
  NAND2_X1 U8841 ( .A1(n8632), .A2(n8606), .ZN(n7175) );
  OAI211_X1 U8842 ( .C1(n7495), .C2(n8603), .A(n9974), .B(n7175), .ZN(n7177)
         );
  NOR2_X1 U8843 ( .A1(n8608), .A2(n7360), .ZN(n7176) );
  AOI211_X1 U8844 ( .C1(n7363), .C2(n8615), .A(n7177), .B(n7176), .ZN(n7178)
         );
  NAND2_X1 U8845 ( .A1(n7179), .A2(n7178), .ZN(P2_U3179) );
  INV_X1 U8846 ( .A(n8699), .ZN(n8670) );
  INV_X1 U8847 ( .A(n7180), .ZN(n7182) );
  INV_X1 U8848 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7181) );
  OAI222_X1 U8849 ( .A1(n8670), .A2(P2_U3151), .B1(n9103), .B2(n7182), .C1(
        n7181), .C2(n7434), .ZN(P2_U3280) );
  INV_X1 U8850 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7183) );
  INV_X1 U8851 ( .A(n8119), .ZN(n8103) );
  OAI222_X1 U8852 ( .A1(n9789), .A2(n7183), .B1(n4336), .B2(n7182), .C1(
        P1_U3086), .C2(n8103), .ZN(P1_U3340) );
  XNOR2_X1 U8853 ( .A(n7184), .B(n7185), .ZN(n10041) );
  INV_X1 U8854 ( .A(n10041), .ZN(n7193) );
  XNOR2_X1 U8855 ( .A(n7186), .B(n7185), .ZN(n7187) );
  AOI222_X1 U8856 ( .A1(n8952), .A2(n7187), .B1(n8634), .B2(n5656), .C1(n8632), 
        .C2(n8949), .ZN(n10039) );
  MUX2_X1 U8857 ( .A(n7188), .B(n10039), .S(n8926), .Z(n7192) );
  AOI22_X1 U8858 ( .A1(n8956), .A2(n7190), .B1(n8955), .B2(n7189), .ZN(n7191)
         );
  OAI211_X1 U8859 ( .C1(n8959), .C2(n7193), .A(n7192), .B(n7191), .ZN(P2_U3229) );
  INV_X1 U8860 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7195) );
  MUX2_X1 U8861 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n7195), .S(n7465), .Z(n7196)
         );
  INV_X1 U8862 ( .A(n7196), .ZN(n7197) );
  NOR2_X1 U8863 ( .A1(n7198), .A2(n7197), .ZN(n7464) );
  AOI211_X1 U8864 ( .C1(n7198), .C2(n7197), .A(n9343), .B(n7464), .ZN(n7206)
         );
  AOI21_X1 U8865 ( .B1(n7200), .B2(P1_REG1_REG_10__SCAN_IN), .A(n7199), .ZN(
        n7451) );
  XNOR2_X1 U8866 ( .A(n7465), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n7450) );
  XNOR2_X1 U8867 ( .A(n7451), .B(n7450), .ZN(n7204) );
  NAND2_X1 U8868 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9811) );
  INV_X1 U8869 ( .A(n9811), .ZN(n7201) );
  AOI21_X1 U8870 ( .B1(n9824), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n7201), .ZN(
        n7203) );
  NAND2_X1 U8871 ( .A1(n9332), .A2(n7465), .ZN(n7202) );
  OAI211_X1 U8872 ( .C1(n7204), .C2(n9849), .A(n7203), .B(n7202), .ZN(n7205)
         );
  OR2_X1 U8873 ( .A1(n7206), .A2(n7205), .ZN(P1_U3254) );
  NAND2_X1 U8874 ( .A1(n9293), .A2(n7247), .ZN(n8386) );
  NAND2_X1 U8875 ( .A1(n7215), .A2(n7485), .ZN(n7234) );
  INV_X1 U8876 ( .A(n9292), .ZN(n7278) );
  NAND2_X1 U8877 ( .A1(n7278), .A2(n7242), .ZN(n7274) );
  AND2_X1 U8878 ( .A1(n7234), .A2(n7274), .ZN(n7208) );
  NAND2_X1 U8879 ( .A1(n7235), .A2(n7208), .ZN(n7211) );
  NAND2_X1 U8880 ( .A1(n9291), .A2(n7290), .ZN(n7210) );
  NAND2_X1 U8881 ( .A1(n9292), .A2(n9864), .ZN(n7209) );
  AND2_X1 U8882 ( .A1(n7210), .A2(n7209), .ZN(n8390) );
  NAND2_X1 U8883 ( .A1(n7303), .A2(n7607), .ZN(n8207) );
  NAND2_X1 U8884 ( .A1(n7506), .A2(n7214), .ZN(n8208) );
  NAND2_X1 U8885 ( .A1(n8208), .A2(n8400), .ZN(n8306) );
  XNOR2_X1 U8886 ( .A(n8203), .B(n8306), .ZN(n7212) );
  OAI222_X1 U8887 ( .A1(n9490), .A2(n7545), .B1(n9488), .B2(n7303), .C1(n7212), 
        .C2(n9592), .ZN(n7626) );
  NAND2_X1 U8888 ( .A1(n7213), .A2(n9864), .ZN(n7273) );
  OR2_X2 U8889 ( .A1(n7273), .A2(n7607), .ZN(n7271) );
  AOI211_X1 U8890 ( .C1(n7214), .C2(n7271), .A(n9595), .B(n7510), .ZN(n7631)
         );
  NOR2_X1 U8891 ( .A1(n7626), .A2(n7631), .ZN(n7254) );
  NAND2_X1 U8892 ( .A1(n7215), .A2(n7247), .ZN(n7216) );
  XNOR2_X1 U8893 ( .A(n9292), .B(n9864), .ZN(n8309) );
  NAND2_X1 U8894 ( .A1(n7278), .A2(n9864), .ZN(n7218) );
  NAND2_X1 U8895 ( .A1(n7270), .A2(n8310), .ZN(n7269) );
  NAND2_X1 U8896 ( .A1(n7303), .A2(n7290), .ZN(n7219) );
  OAI21_X1 U8897 ( .B1(n7220), .B2(n8306), .A(n7508), .ZN(n7625) );
  INV_X1 U8898 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7221) );
  OAI22_X1 U8899 ( .A1(n9759), .A2(n7629), .B1(n9890), .B2(n7221), .ZN(n7222)
         );
  AOI21_X1 U8900 ( .B1(n7625), .B2(n7869), .A(n7222), .ZN(n7223) );
  OAI21_X1 U8901 ( .B1(n7254), .B2(n9888), .A(n7223), .ZN(P1_U3468) );
  OAI22_X1 U8902 ( .A1(n8912), .A2(n7224), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n10021), .ZN(n7227) );
  MUX2_X1 U8903 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7225), .S(n8926), .Z(n7226)
         );
  AOI211_X1 U8904 ( .C1(n8914), .C2(n7228), .A(n7227), .B(n7226), .ZN(n7229)
         );
  INV_X1 U8905 ( .A(n7229), .ZN(P2_U3230) );
  OAI21_X1 U8906 ( .B1(n7231), .B2(n8309), .A(n7230), .ZN(n9867) );
  INV_X1 U8907 ( .A(n7273), .ZN(n7232) );
  AOI211_X1 U8908 ( .C1(n7242), .C2(n7233), .A(n9595), .B(n7232), .ZN(n9859)
         );
  AND2_X1 U8909 ( .A1(n7235), .A2(n7234), .ZN(n7275) );
  XNOR2_X1 U8910 ( .A(n7275), .B(n8309), .ZN(n7237) );
  AOI21_X1 U8911 ( .B1(n7237), .B2(n9608), .A(n7236), .ZN(n9870) );
  INV_X1 U8912 ( .A(n9870), .ZN(n7238) );
  AOI211_X1 U8913 ( .C1(n9878), .C2(n9867), .A(n9859), .B(n7238), .ZN(n7244)
         );
  INV_X1 U8914 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7239) );
  OAI22_X1 U8915 ( .A1(n9759), .A2(n9864), .B1(n9890), .B2(n7239), .ZN(n7240)
         );
  INV_X1 U8916 ( .A(n7240), .ZN(n7241) );
  OAI21_X1 U8917 ( .B1(n7244), .B2(n9888), .A(n7241), .ZN(P1_U3462) );
  AOI22_X1 U8918 ( .A1(n9695), .A2(n7242), .B1(n9893), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n7243) );
  OAI21_X1 U8919 ( .B1(n7244), .B2(n9893), .A(n7243), .ZN(P1_U3525) );
  INV_X1 U8920 ( .A(n7245), .ZN(n7285) );
  AOI22_X1 U8921 ( .A1(n9331), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9781), .ZN(n7246) );
  OAI21_X1 U8922 ( .B1(n7285), .B2(n4336), .A(n7246), .ZN(P1_U3339) );
  NAND2_X1 U8923 ( .A1(n9896), .A2(n9878), .ZN(n9700) );
  INV_X1 U8924 ( .A(n9700), .ZN(n7872) );
  OAI22_X1 U8925 ( .A1(n9686), .A2(n7247), .B1(n9896), .B2(n6770), .ZN(n7248)
         );
  AOI21_X1 U8926 ( .B1(n7872), .B2(n7490), .A(n7248), .ZN(n7249) );
  OAI21_X1 U8927 ( .B1(n7250), .B2(n9893), .A(n7249), .ZN(P1_U3524) );
  OAI22_X1 U8928 ( .A1(n9686), .A2(n7629), .B1(n9896), .B2(n7251), .ZN(n7252)
         );
  AOI21_X1 U8929 ( .B1(n7625), .B2(n7872), .A(n7252), .ZN(n7253) );
  OAI21_X1 U8930 ( .B1(n7254), .B2(n9893), .A(n7253), .ZN(P1_U3527) );
  INV_X1 U8931 ( .A(n7255), .ZN(n7256) );
  NAND2_X1 U8932 ( .A1(n7256), .A2(n8631), .ZN(n7257) );
  XNOR2_X1 U8933 ( .A(n7400), .B(n7495), .ZN(n7259) );
  OAI21_X1 U8934 ( .B1(n4424), .B2(n7259), .A(n7402), .ZN(n7260) );
  NAND2_X1 U8935 ( .A1(n7260), .A2(n8588), .ZN(n7266) );
  INV_X1 U8936 ( .A(n7375), .ZN(n7264) );
  INV_X1 U8937 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7261) );
  NOR2_X1 U8938 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7261), .ZN(n9982) );
  AOI21_X1 U8939 ( .B1(n8631), .B2(n8606), .A(n9982), .ZN(n7262) );
  OAI21_X1 U8940 ( .B1(n7475), .B2(n8603), .A(n7262), .ZN(n7263) );
  AOI21_X1 U8941 ( .B1(n7264), .B2(n8593), .A(n7263), .ZN(n7265) );
  OAI211_X1 U8942 ( .C1(n10053), .C2(n8596), .A(n7266), .B(n7265), .ZN(
        P2_U3153) );
  INV_X1 U8943 ( .A(n7267), .ZN(n7287) );
  AOI22_X1 U8944 ( .A1(n8744), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n9100), .ZN(n7268) );
  OAI21_X1 U8945 ( .B1(n7287), .B2(n9103), .A(n7268), .ZN(P2_U3278) );
  OAI21_X1 U8946 ( .B1(n7270), .B2(n8310), .A(n7269), .ZN(n7613) );
  INV_X1 U8947 ( .A(n7271), .ZN(n7272) );
  AOI211_X1 U8948 ( .C1(n7607), .C2(n7273), .A(n9595), .B(n7272), .ZN(n7605)
         );
  OAI21_X1 U8949 ( .B1(n7275), .B2(n8309), .A(n7274), .ZN(n7276) );
  XNOR2_X1 U8950 ( .A(n7276), .B(n8310), .ZN(n7277) );
  OAI222_X1 U8951 ( .A1(n9490), .A2(n7506), .B1(n9488), .B2(n7278), .C1(n9592), 
        .C2(n7277), .ZN(n7610) );
  AOI211_X1 U8952 ( .C1(n9878), .C2(n7613), .A(n7605), .B(n7610), .ZN(n7283)
         );
  INV_X1 U8953 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7279) );
  OAI22_X1 U8954 ( .A1(n9759), .A2(n7290), .B1(n9890), .B2(n7279), .ZN(n7280)
         );
  INV_X1 U8955 ( .A(n7280), .ZN(n7281) );
  OAI21_X1 U8956 ( .B1(n7283), .B2(n9888), .A(n7281), .ZN(P1_U3465) );
  AOI22_X1 U8957 ( .A1(n9695), .A2(n7607), .B1(n9893), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n7282) );
  OAI21_X1 U8958 ( .B1(n7283), .B2(n9893), .A(n7282), .ZN(P1_U3526) );
  OAI222_X1 U8959 ( .A1(P2_U3151), .A2(n8721), .B1(n9103), .B2(n7285), .C1(
        n7284), .C2(n7434), .ZN(P2_U3279) );
  INV_X2 U8960 ( .A(P1_U3973), .ZN(n9294) );
  NAND2_X1 U8961 ( .A1(n9294), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7286) );
  OAI21_X1 U8962 ( .B1(n8163), .B2(n9294), .A(n7286), .ZN(P1_U3583) );
  INV_X1 U8963 ( .A(n8125), .ZN(n9848) );
  OAI222_X1 U8964 ( .A1(n9789), .A2(n10271), .B1(n4336), .B2(n7287), .C1(
        P1_U3086), .C2(n9848), .ZN(P1_U3338) );
  INV_X1 U8965 ( .A(n9803), .ZN(n9148) );
  AOI22_X1 U8966 ( .A1(n9148), .A2(n9292), .B1(n9802), .B2(n9290), .ZN(n7289)
         );
  OAI211_X1 U8967 ( .C1(n7290), .C2(n9800), .A(n7289), .B(n7288), .ZN(n7296)
         );
  INV_X1 U8968 ( .A(n7292), .ZN(n7293) );
  AOI211_X1 U8969 ( .C1(n7294), .C2(n7291), .A(n9245), .B(n7293), .ZN(n7295)
         );
  AOI211_X1 U8970 ( .C1(n7606), .C2(n9267), .A(n7296), .B(n7295), .ZN(n7297)
         );
  INV_X1 U8971 ( .A(n7297), .ZN(P1_U3230) );
  NAND2_X1 U8972 ( .A1(n5078), .A2(n7298), .ZN(n7300) );
  XNOR2_X1 U8973 ( .A(n7300), .B(n7299), .ZN(n7307) );
  OAI21_X1 U8974 ( .B1(n9800), .B2(n7629), .A(n7301), .ZN(n7305) );
  NAND2_X1 U8975 ( .A1(n9802), .A2(n9289), .ZN(n7302) );
  OAI21_X1 U8976 ( .B1(n7303), .B2(n9803), .A(n7302), .ZN(n7304) );
  AOI211_X1 U8977 ( .C1(n7627), .C2(n9267), .A(n7305), .B(n7304), .ZN(n7306)
         );
  OAI21_X1 U8978 ( .B1(n7307), .B2(n9245), .A(n7306), .ZN(P1_U3227) );
  NOR2_X1 U8979 ( .A1(n9939), .A2(n7309), .ZN(n7310) );
  INV_X1 U8980 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10087) );
  XNOR2_X1 U8981 ( .A(n9939), .B(n7309), .ZN(n9937) );
  INV_X1 U8982 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7311) );
  MUX2_X1 U8983 ( .A(n7311), .B(P2_REG1_REG_6__SCAN_IN), .S(n9959), .Z(n9969)
         );
  NAND2_X1 U8984 ( .A1(n9959), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7312) );
  INV_X1 U8985 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7314) );
  MUX2_X1 U8986 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7314), .S(n10002), .Z(n9999)
         );
  NAND2_X1 U8987 ( .A1(n7344), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7315) );
  INV_X1 U8988 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10121) );
  AOI21_X1 U8989 ( .B1(n7316), .B2(n10121), .A(n7422), .ZN(n7352) );
  MUX2_X1 U8990 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8643), .Z(n7327) );
  NOR2_X1 U8991 ( .A1(n7327), .A2(n7344), .ZN(n7329) );
  MUX2_X1 U8992 ( .A(n7376), .B(n7317), .S(n8643), .Z(n7326) );
  INV_X1 U8993 ( .A(n9959), .ZN(n7325) );
  MUX2_X1 U8994 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8643), .Z(n7323) );
  INV_X1 U8995 ( .A(n7323), .ZN(n7324) );
  MUX2_X1 U8996 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8643), .Z(n7321) );
  XNOR2_X1 U8997 ( .A(n7321), .B(n7338), .ZN(n9948) );
  INV_X1 U8998 ( .A(n7321), .ZN(n7322) );
  OAI22_X1 U8999 ( .A1(n9947), .A2(n9948), .B1(n9939), .B2(n7322), .ZN(n9964)
         );
  XNOR2_X1 U9000 ( .A(n7323), .B(n9959), .ZN(n9965) );
  NOR2_X1 U9001 ( .A1(n9964), .A2(n9965), .ZN(n9963) );
  XNOR2_X1 U9002 ( .A(n7326), .B(n9983), .ZN(n9989) );
  AOI21_X1 U9003 ( .B1(n7327), .B2(n7344), .A(n7329), .ZN(n7328) );
  INV_X1 U9004 ( .A(n7328), .ZN(n10011) );
  MUX2_X1 U9005 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8643), .Z(n7331) );
  INV_X1 U9006 ( .A(n7421), .ZN(n7330) );
  OR2_X1 U9007 ( .A1(n7331), .A2(n7330), .ZN(n7413) );
  AND2_X1 U9008 ( .A1(n7331), .A2(n7330), .ZN(n7415) );
  INV_X1 U9009 ( .A(n7415), .ZN(n7332) );
  NAND2_X1 U9010 ( .A1(n7413), .A2(n7332), .ZN(n7333) );
  XNOR2_X1 U9011 ( .A(n7414), .B(n7333), .ZN(n7334) );
  NAND2_X1 U9012 ( .A1(n7334), .A2(n9949), .ZN(n7351) );
  INV_X1 U9013 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n8075) );
  AND2_X1 U9014 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7477) );
  INV_X1 U9015 ( .A(n7477), .ZN(n7335) );
  OAI21_X1 U9016 ( .B1(n10017), .B2(n8075), .A(n7335), .ZN(n7349) );
  MUX2_X1 U9017 ( .A(n7361), .B(P2_REG2_REG_6__SCAN_IN), .S(n9959), .Z(n9956)
         );
  NAND2_X1 U9018 ( .A1(n9959), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7340) );
  MUX2_X1 U9019 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7343), .S(n10002), .Z(n9995)
         );
  NAND2_X1 U9020 ( .A1(n7344), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7345) );
  AOI21_X1 U9021 ( .B1(n5389), .B2(n7346), .A(n7409), .ZN(n7347) );
  NOR2_X1 U9022 ( .A1(n7347), .A2(n9980), .ZN(n7348) );
  AOI211_X1 U9023 ( .C1(n10003), .C2(n7421), .A(n7349), .B(n7348), .ZN(n7350)
         );
  OAI211_X1 U9024 ( .C1(n7352), .C2(n10005), .A(n7351), .B(n7350), .ZN(
        P2_U3191) );
  NAND2_X1 U9025 ( .A1(n7354), .A2(n7353), .ZN(n7355) );
  XOR2_X1 U9026 ( .A(n7357), .B(n7355), .Z(n10048) );
  XNOR2_X1 U9027 ( .A(n7356), .B(n7357), .ZN(n7358) );
  OAI222_X1 U9028 ( .A1(n10030), .A2(n7495), .B1(n10028), .B2(n7359), .C1(
        n10026), .C2(n7358), .ZN(n10050) );
  NAND2_X1 U9029 ( .A1(n10050), .A2(n8926), .ZN(n7365) );
  OAI22_X1 U9030 ( .A1(n8926), .A2(n7361), .B1(n7360), .B2(n10021), .ZN(n7362)
         );
  AOI21_X1 U9031 ( .B1(n8956), .B2(n7363), .A(n7362), .ZN(n7364) );
  OAI211_X1 U9032 ( .C1(n10048), .C2(n8959), .A(n7365), .B(n7364), .ZN(
        P2_U3227) );
  OR2_X1 U9033 ( .A1(n7368), .A2(n7367), .ZN(n7369) );
  NAND2_X1 U9034 ( .A1(n7366), .A2(n7369), .ZN(n10054) );
  XNOR2_X1 U9035 ( .A(n7370), .B(n7371), .ZN(n7372) );
  NAND2_X1 U9036 ( .A1(n7372), .A2(n8952), .ZN(n7374) );
  AOI22_X1 U9037 ( .A1(n8949), .A2(n8629), .B1(n8631), .B2(n5656), .ZN(n7373)
         );
  NAND2_X1 U9038 ( .A1(n7374), .A2(n7373), .ZN(n10057) );
  NAND2_X1 U9039 ( .A1(n10057), .A2(n8926), .ZN(n7380) );
  OAI22_X1 U9040 ( .A1(n8926), .A2(n7376), .B1(n7375), .B2(n10021), .ZN(n7377)
         );
  AOI21_X1 U9041 ( .B1(n8956), .B2(n7378), .A(n7377), .ZN(n7379) );
  OAI211_X1 U9042 ( .C1(n8959), .C2(n10054), .A(n7380), .B(n7379), .ZN(
        P2_U3226) );
  XNOR2_X1 U9043 ( .A(n7383), .B(n7382), .ZN(n7384) );
  XNOR2_X1 U9044 ( .A(n7381), .B(n7384), .ZN(n7389) );
  AOI22_X1 U9045 ( .A1(n9148), .A2(n9290), .B1(n9802), .B2(n7518), .ZN(n7386)
         );
  INV_X1 U9046 ( .A(n9875), .ZN(n7512) );
  AOI22_X1 U9047 ( .A1(n6649), .A2(n7512), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n7385) );
  OAI211_X1 U9048 ( .C1(n9814), .C2(n7387), .A(n7386), .B(n7385), .ZN(n7388)
         );
  AOI21_X1 U9049 ( .B1(n7389), .B2(n9809), .A(n7388), .ZN(n7390) );
  INV_X1 U9050 ( .A(n7390), .ZN(P1_U3239) );
  XOR2_X1 U9051 ( .A(n7391), .B(n7393), .Z(n10044) );
  XOR2_X1 U9052 ( .A(n7392), .B(n7393), .Z(n7394) );
  AOI222_X1 U9053 ( .A1(n8952), .A2(n7394), .B1(n8631), .B2(n8949), .C1(n8633), 
        .C2(n5656), .ZN(n10042) );
  MUX2_X1 U9054 ( .A(n7395), .B(n10042), .S(n8926), .Z(n7399) );
  AOI22_X1 U9055 ( .A1(n8956), .A2(n7397), .B1(n8955), .B2(n7396), .ZN(n7398)
         );
  OAI211_X1 U9056 ( .C1(n10044), .C2(n8959), .A(n7399), .B(n7398), .ZN(
        P2_U3228) );
  INV_X1 U9057 ( .A(n7400), .ZN(n7401) );
  XNOR2_X1 U9058 ( .A(n7560), .B(n8491), .ZN(n7583) );
  XNOR2_X1 U9059 ( .A(n7590), .B(n7583), .ZN(n7472) );
  XNOR2_X1 U9060 ( .A(n7472), .B(n8629), .ZN(n7407) );
  AND2_X1 U9061 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n10001) );
  AOI21_X1 U9062 ( .B1(n8630), .B2(n8606), .A(n10001), .ZN(n7404) );
  NAND2_X1 U9063 ( .A1(n8593), .A2(n7499), .ZN(n7403) );
  OAI211_X1 U9064 ( .C1(n7595), .C2(n8603), .A(n7404), .B(n7403), .ZN(n7405)
         );
  AOI21_X1 U9065 ( .B1(n7560), .B2(n8615), .A(n7405), .ZN(n7406) );
  OAI21_X1 U9066 ( .B1(n7407), .B2(n8610), .A(n7406), .ZN(P2_U3161) );
  MUX2_X1 U9067 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7732), .S(n7429), .Z(n7411)
         );
  INV_X1 U9068 ( .A(n7747), .ZN(n7410) );
  AOI21_X1 U9069 ( .B1(n7412), .B2(n7411), .A(n7410), .ZN(n7432) );
  OAI21_X1 U9070 ( .B1(n7415), .B2(n7414), .A(n7413), .ZN(n7417) );
  MUX2_X1 U9071 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8643), .Z(n7739) );
  XNOR2_X1 U9072 ( .A(n7739), .B(n7429), .ZN(n7416) );
  OAI21_X1 U9073 ( .B1(n7417), .B2(n7416), .A(n7740), .ZN(n7418) );
  NAND2_X1 U9074 ( .A1(n7418), .A2(n9949), .ZN(n7431) );
  INV_X1 U9075 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8079) );
  INV_X1 U9076 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7419) );
  OR2_X1 U9077 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7419), .ZN(n7594) );
  OAI21_X1 U9078 ( .B1(n10017), .B2(n8079), .A(n7594), .ZN(n7428) );
  INV_X1 U9079 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7423) );
  MUX2_X1 U9080 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7423), .S(n7429), .Z(n7424)
         );
  NAND2_X1 U9081 ( .A1(n7425), .A2(n7424), .ZN(n7426) );
  AOI21_X1 U9082 ( .B1(n7737), .B2(n7426), .A(n10005), .ZN(n7427) );
  AOI211_X1 U9083 ( .C1(n10003), .C2(n7429), .A(n7428), .B(n7427), .ZN(n7430)
         );
  OAI211_X1 U9084 ( .C1(n7432), .C2(n9980), .A(n7431), .B(n7430), .ZN(P2_U3192) );
  INV_X1 U9085 ( .A(n7433), .ZN(n7437) );
  OAI222_X1 U9086 ( .A1(n7434), .A2(n10244), .B1(n9103), .B2(n7437), .C1(
        P2_U3151), .C2(n8747), .ZN(P2_U3277) );
  INV_X1 U9087 ( .A(n7435), .ZN(n8057) );
  AOI22_X1 U9088 ( .A1(n8767), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n9100), .ZN(n7436) );
  OAI21_X1 U9089 ( .B1(n8057), .B2(n9103), .A(n7436), .ZN(P2_U3276) );
  INV_X1 U9090 ( .A(n8126), .ZN(n9351) );
  OAI222_X1 U9091 ( .A1(n9789), .A2(n7438), .B1(n9351), .B2(P1_U3086), .C1(
        n4336), .C2(n7437), .ZN(P1_U3337) );
  NAND2_X1 U9092 ( .A1(n7440), .A2(n7439), .ZN(n7441) );
  XNOR2_X1 U9093 ( .A(n7442), .B(n7441), .ZN(n7448) );
  INV_X1 U9094 ( .A(n7644), .ZN(n7446) );
  INV_X1 U9095 ( .A(n7553), .ZN(n7646) );
  OAI22_X1 U9096 ( .A1(n7646), .A2(n9800), .B1(n9803), .B2(n7545), .ZN(n7443)
         );
  INV_X1 U9097 ( .A(n7443), .ZN(n7445) );
  INV_X1 U9098 ( .A(n7760), .ZN(n9288) );
  AOI22_X1 U9099 ( .A1(n9802), .A2(n9288), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n7444) );
  OAI211_X1 U9100 ( .C1(n9814), .C2(n7446), .A(n7445), .B(n7444), .ZN(n7447)
         );
  AOI21_X1 U9101 ( .B1(n7448), .B2(n9809), .A(n7447), .ZN(n7449) );
  INV_X1 U9102 ( .A(n7449), .ZN(P1_U3213) );
  INV_X1 U9103 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7454) );
  OR2_X1 U9104 ( .A1(n7451), .A2(n7450), .ZN(n7452) );
  OAI21_X1 U9105 ( .B1(n7454), .B2(n7453), .A(n7452), .ZN(n9833) );
  INV_X1 U9106 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7455) );
  AOI22_X1 U9107 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n9834), .B1(n7466), .B2(
        n7455), .ZN(n9832) );
  NOR2_X1 U9108 ( .A1(n9833), .A2(n9832), .ZN(n9831) );
  NOR2_X1 U9109 ( .A1(n7466), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7456) );
  NOR2_X1 U9110 ( .A1(n9831), .A2(n7456), .ZN(n7458) );
  INV_X1 U9111 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7710) );
  XNOR2_X1 U9112 ( .A(n7717), .B(n7710), .ZN(n7457) );
  NAND2_X1 U9113 ( .A1(n7457), .A2(n7458), .ZN(n7709) );
  OAI211_X1 U9114 ( .C1(n7458), .C2(n7457), .A(n7709), .B(n9340), .ZN(n7461)
         );
  NAND2_X1 U9115 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9219) );
  INV_X1 U9116 ( .A(n9219), .ZN(n7459) );
  AOI21_X1 U9117 ( .B1(n9824), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n7459), .ZN(
        n7460) );
  OAI211_X1 U9118 ( .C1(n9847), .C2(n7711), .A(n7461), .B(n7460), .ZN(n7470)
         );
  INV_X1 U9119 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7462) );
  AOI22_X1 U9120 ( .A1(n7717), .A2(n7462), .B1(P1_REG2_REG_13__SCAN_IN), .B2(
        n7711), .ZN(n7468) );
  INV_X1 U9121 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7463) );
  AOI22_X1 U9122 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7466), .B1(n9834), .B2(
        n7463), .ZN(n9830) );
  AOI21_X1 U9123 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7465), .A(n7464), .ZN(
        n9829) );
  NAND2_X1 U9124 ( .A1(n9830), .A2(n9829), .ZN(n9828) );
  OAI21_X1 U9125 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7466), .A(n9828), .ZN(
        n7467) );
  AOI211_X1 U9126 ( .C1(n7468), .C2(n7467), .A(n7716), .B(n9343), .ZN(n7469)
         );
  OR2_X1 U9127 ( .A1(n7470), .A2(n7469), .ZN(P1_U3256) );
  INV_X1 U9128 ( .A(n7583), .ZN(n7471) );
  AOI22_X1 U9129 ( .A1(n7472), .A2(n7475), .B1(n7590), .B2(n7471), .ZN(n7474)
         );
  XNOR2_X1 U9130 ( .A(n10062), .B(n4329), .ZN(n7584) );
  XNOR2_X1 U9131 ( .A(n7584), .B(n8628), .ZN(n7473) );
  XNOR2_X1 U9132 ( .A(n7474), .B(n7473), .ZN(n7481) );
  NOR2_X1 U9133 ( .A1(n7475), .A2(n8574), .ZN(n7476) );
  AOI211_X1 U9134 ( .C1(n8571), .C2(n8627), .A(n7477), .B(n7476), .ZN(n7478)
         );
  OAI21_X1 U9135 ( .B1(n7621), .B2(n8608), .A(n7478), .ZN(n7479) );
  AOI21_X1 U9136 ( .B1(n10062), .B2(n8615), .A(n7479), .ZN(n7480) );
  OAI21_X1 U9137 ( .B1(n7481), .B2(n8610), .A(n7480), .ZN(P2_U3171) );
  AND2_X1 U9138 ( .A1(n7781), .A2(n7529), .ZN(n7482) );
  INV_X1 U9139 ( .A(n7483), .ZN(n7484) );
  NOR2_X2 U9140 ( .A1(n9617), .A2(n7484), .ZN(n9618) );
  NAND2_X1 U9141 ( .A1(n9618), .A2(n7485), .ZN(n7487) );
  INV_X2 U9142 ( .A(n9544), .ZN(n9861) );
  AOI22_X1 U9143 ( .A1(n9617), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9861), .ZN(n7486) );
  OAI211_X1 U9144 ( .C1(n7488), .C2(n9621), .A(n7487), .B(n7486), .ZN(n7489)
         );
  AOI21_X1 U9145 ( .B1(n9868), .B2(n7490), .A(n7489), .ZN(n7491) );
  OAI21_X1 U9146 ( .B1(n7492), .B2(n9617), .A(n7491), .ZN(P1_U3291) );
  XOR2_X1 U9147 ( .A(n7497), .B(n7493), .Z(n7494) );
  OAI222_X1 U9148 ( .A1(n10028), .A2(n7495), .B1(n10030), .B2(n7595), .C1(
        n10026), .C2(n7494), .ZN(n7556) );
  INV_X1 U9149 ( .A(n7556), .ZN(n7504) );
  NAND2_X1 U9150 ( .A1(n7366), .A2(n7496), .ZN(n7498) );
  XNOR2_X1 U9151 ( .A(n7498), .B(n7497), .ZN(n7557) );
  INV_X1 U9152 ( .A(n7560), .ZN(n7501) );
  AOI22_X1 U9153 ( .A1(n10034), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n8955), .B2(
        n7499), .ZN(n7500) );
  OAI21_X1 U9154 ( .B1(n7501), .B2(n8912), .A(n7500), .ZN(n7502) );
  AOI21_X1 U9155 ( .B1(n7557), .B2(n8914), .A(n7502), .ZN(n7503) );
  OAI21_X1 U9156 ( .B1(n7504), .B2(n10034), .A(n7503), .ZN(P2_U3225) );
  NAND2_X1 U9157 ( .A1(n9875), .A2(n9289), .ZN(n8205) );
  NAND2_X1 U9158 ( .A1(n7545), .A2(n7512), .ZN(n8210) );
  NAND2_X1 U9159 ( .A1(n8205), .A2(n8210), .ZN(n7541) );
  XNOR2_X1 U9160 ( .A(n7542), .B(n7541), .ZN(n7505) );
  AOI222_X1 U9161 ( .A1(n9608), .A2(n7505), .B1(n7518), .B2(n9524), .C1(n9290), 
        .C2(n9523), .ZN(n9874) );
  NAND2_X1 U9162 ( .A1(n7506), .A2(n7629), .ZN(n7507) );
  OAI21_X1 U9163 ( .B1(n7509), .B2(n7541), .A(n7517), .ZN(n9877) );
  INV_X1 U9164 ( .A(n7530), .ZN(n7540) );
  OAI211_X1 U9165 ( .C1(n9875), .C2(n7510), .A(n7540), .B(n9613), .ZN(n9873)
         );
  AOI22_X1 U9166 ( .A1(n9617), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7511), .B2(
        n9861), .ZN(n7514) );
  NAND2_X1 U9167 ( .A1(n9618), .A2(n7512), .ZN(n7513) );
  OAI211_X1 U9168 ( .C1(n9873), .C2(n9621), .A(n7514), .B(n7513), .ZN(n7515)
         );
  AOI21_X1 U9169 ( .B1(n9877), .B2(n9868), .A(n7515), .ZN(n7516) );
  OAI21_X1 U9170 ( .B1(n9874), .B2(n9617), .A(n7516), .ZN(P1_U3287) );
  OR2_X1 U9171 ( .A1(n7553), .A2(n7703), .ZN(n7665) );
  NAND2_X1 U9172 ( .A1(n7665), .A2(n7663), .ZN(n7543) );
  NAND2_X1 U9173 ( .A1(n7537), .A2(n7543), .ZN(n7536) );
  OR2_X1 U9174 ( .A1(n7553), .A2(n7518), .ZN(n7519) );
  NAND2_X1 U9175 ( .A1(n7697), .A2(n7760), .ZN(n8219) );
  NAND2_X1 U9176 ( .A1(n8214), .A2(n8219), .ZN(n7569) );
  OR2_X1 U9177 ( .A1(n7520), .A2(n7569), .ZN(n7521) );
  NAND2_X1 U9178 ( .A1(n7567), .A2(n7521), .ZN(n9885) );
  INV_X1 U9179 ( .A(n7781), .ZN(n7528) );
  NAND2_X1 U9180 ( .A1(n7542), .A2(n8210), .ZN(n7668) );
  INV_X1 U9181 ( .A(n8205), .ZN(n7666) );
  NOR2_X1 U9182 ( .A1(n7543), .A2(n7666), .ZN(n7522) );
  NAND2_X1 U9183 ( .A1(n7668), .A2(n7522), .ZN(n7570) );
  NAND2_X1 U9184 ( .A1(n7570), .A2(n7663), .ZN(n7523) );
  XNOR2_X1 U9185 ( .A(n7523), .B(n7569), .ZN(n7526) );
  OAI22_X1 U9186 ( .A1(n7703), .A2(n9488), .B1(n7672), .B2(n9490), .ZN(n7524)
         );
  INV_X1 U9187 ( .A(n7524), .ZN(n7525) );
  OAI21_X1 U9188 ( .B1(n7526), .B2(n9592), .A(n7525), .ZN(n7527) );
  AOI21_X1 U9189 ( .B1(n9885), .B2(n7528), .A(n7527), .ZN(n9887) );
  NOR2_X1 U9190 ( .A1(n9617), .A2(n7529), .ZN(n7787) );
  NAND2_X1 U9191 ( .A1(n7530), .A2(n7646), .ZN(n7538) );
  AOI21_X1 U9192 ( .B1(n7538), .B2(n7697), .A(n9595), .ZN(n7531) );
  OR2_X1 U9193 ( .A1(n7538), .A2(n7697), .ZN(n7678) );
  NAND2_X1 U9194 ( .A1(n7531), .A2(n7678), .ZN(n9880) );
  AOI22_X1 U9195 ( .A1(n9617), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n5085), .B2(
        n9861), .ZN(n7533) );
  NAND2_X1 U9196 ( .A1(n9618), .A2(n7697), .ZN(n7532) );
  OAI211_X1 U9197 ( .C1(n9880), .C2(n9621), .A(n7533), .B(n7532), .ZN(n7534)
         );
  AOI21_X1 U9198 ( .B1(n9885), .B2(n7787), .A(n7534), .ZN(n7535) );
  OAI21_X1 U9199 ( .B1(n9887), .B2(n9617), .A(n7535), .ZN(P1_U3285) );
  OAI21_X1 U9200 ( .B1(n7537), .B2(n7543), .A(n7536), .ZN(n7549) );
  INV_X1 U9201 ( .A(n7538), .ZN(n7539) );
  AOI211_X1 U9202 ( .C1(n7553), .C2(n7540), .A(n9595), .B(n7539), .ZN(n7648)
         );
  INV_X1 U9203 ( .A(n7549), .ZN(n7652) );
  INV_X1 U9204 ( .A(n7541), .ZN(n8313) );
  AOI21_X1 U9205 ( .B1(n7542), .B2(n8313), .A(n7666), .ZN(n7544) );
  INV_X1 U9206 ( .A(n7543), .ZN(n8213) );
  OAI21_X1 U9207 ( .B1(n7544), .B2(n8213), .A(n7570), .ZN(n7547) );
  OAI22_X1 U9208 ( .A1(n7545), .A2(n9488), .B1(n7760), .B2(n9490), .ZN(n7546)
         );
  AOI21_X1 U9209 ( .B1(n7547), .B2(n9608), .A(n7546), .ZN(n7548) );
  OAI21_X1 U9210 ( .B1(n7652), .B2(n7781), .A(n7548), .ZN(n7643) );
  AOI211_X1 U9211 ( .C1(n9884), .C2(n7549), .A(n7648), .B(n7643), .ZN(n7555)
         );
  INV_X1 U9212 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7550) );
  OAI22_X1 U9213 ( .A1(n9759), .A2(n7646), .B1(n9890), .B2(n7550), .ZN(n7551)
         );
  INV_X1 U9214 ( .A(n7551), .ZN(n7552) );
  OAI21_X1 U9215 ( .B1(n7555), .B2(n9888), .A(n7552), .ZN(P1_U3474) );
  AOI22_X1 U9216 ( .A1(n9695), .A2(n7553), .B1(n9893), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7554) );
  OAI21_X1 U9217 ( .B1(n7555), .B2(n9893), .A(n7554), .ZN(P1_U3529) );
  AOI21_X1 U9218 ( .B1(n10075), .B2(n7557), .A(n7556), .ZN(n7562) );
  AOI22_X1 U9219 ( .A1(n7560), .A2(n9006), .B1(n10094), .B2(
        P2_REG1_REG_8__SCAN_IN), .ZN(n7558) );
  OAI21_X1 U9220 ( .B1(n7562), .B2(n10094), .A(n7558), .ZN(P2_U3467) );
  NOR2_X1 U9221 ( .A1(n10081), .A2(n5373), .ZN(n7559) );
  AOI21_X1 U9222 ( .B1(n9079), .B2(n7560), .A(n7559), .ZN(n7561) );
  OAI21_X1 U9223 ( .B1(n7562), .B2(n10082), .A(n7561), .ZN(P2_U3414) );
  INV_X1 U9224 ( .A(n7601), .ZN(n7565) );
  AOI22_X1 U9225 ( .A1(n7563), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n9100), .ZN(n7564) );
  OAI21_X1 U9226 ( .B1(n7565), .B2(n8046), .A(n7564), .ZN(P2_U3275) );
  NAND2_X1 U9227 ( .A1(n7760), .A2(n9882), .ZN(n7566) );
  NAND2_X1 U9228 ( .A1(n8224), .A2(n8239), .ZN(n7572) );
  OAI21_X1 U9229 ( .B1(n7568), .B2(n7572), .A(n7673), .ZN(n7653) );
  NAND3_X1 U9230 ( .A1(n7570), .A2(n4962), .A3(n7663), .ZN(n7571) );
  NAND2_X1 U9231 ( .A1(n7571), .A2(n8214), .ZN(n7573) );
  XNOR2_X1 U9232 ( .A(n7573), .B(n7572), .ZN(n7574) );
  NAND2_X1 U9233 ( .A1(n7574), .A2(n9608), .ZN(n7576) );
  OR2_X1 U9234 ( .A1(n7760), .A2(n9488), .ZN(n7575) );
  NAND2_X1 U9235 ( .A1(n7576), .A2(n7575), .ZN(n7660) );
  XNOR2_X1 U9236 ( .A(n7678), .B(n7763), .ZN(n7577) );
  OAI22_X1 U9237 ( .A1(n7577), .A2(n9595), .B1(n9804), .B2(n9490), .ZN(n7654)
         );
  AOI211_X1 U9238 ( .C1(n7653), .C2(n9878), .A(n7660), .B(n7654), .ZN(n7582)
         );
  INV_X1 U9239 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7578) );
  NOR2_X1 U9240 ( .A1(n9890), .A2(n7578), .ZN(n7579) );
  AOI21_X1 U9241 ( .B1(n7763), .B2(n9769), .A(n7579), .ZN(n7580) );
  OAI21_X1 U9242 ( .B1(n7582), .B2(n9888), .A(n7580), .ZN(P1_U3480) );
  AOI22_X1 U9243 ( .A1(n7763), .A2(n9695), .B1(n9893), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n7581) );
  OAI21_X1 U9244 ( .B1(n7582), .B2(n9893), .A(n7581), .ZN(P1_U3531) );
  NAND2_X1 U9245 ( .A1(n7584), .A2(n7595), .ZN(n7587) );
  OAI21_X1 U9246 ( .B1(n7583), .B2(n8629), .A(n7587), .ZN(n7589) );
  AND2_X1 U9247 ( .A1(n7583), .A2(n8629), .ZN(n7586) );
  INV_X1 U9248 ( .A(n7584), .ZN(n7585) );
  AOI22_X1 U9249 ( .A1(n7587), .A2(n7586), .B1(n7585), .B2(n8628), .ZN(n7588)
         );
  INV_X1 U9250 ( .A(n7767), .ZN(n7592) );
  NOR2_X1 U9251 ( .A1(n7766), .A2(n7592), .ZN(n7593) );
  XNOR2_X1 U9252 ( .A(n10067), .B(n8491), .ZN(n7768) );
  XNOR2_X1 U9253 ( .A(n7593), .B(n7768), .ZN(n7600) );
  OAI21_X1 U9254 ( .B1(n7595), .B2(n8574), .A(n7594), .ZN(n7596) );
  AOI21_X1 U9255 ( .B1(n8571), .B2(n8626), .A(n7596), .ZN(n7597) );
  OAI21_X1 U9256 ( .B1(n7731), .B2(n8608), .A(n7597), .ZN(n7598) );
  AOI21_X1 U9257 ( .B1(n10067), .B2(n8615), .A(n7598), .ZN(n7599) );
  OAI21_X1 U9258 ( .B1(n7600), .B2(n8610), .A(n7599), .ZN(P2_U3157) );
  NAND2_X1 U9259 ( .A1(n7601), .A2(n7905), .ZN(n7603) );
  OAI211_X1 U9260 ( .C1(n7604), .C2(n9789), .A(n7603), .B(n7602), .ZN(P1_U3335) );
  INV_X1 U9261 ( .A(n7605), .ZN(n7609) );
  AOI22_X1 U9262 ( .A1(n9618), .A2(n7607), .B1(n9861), .B2(n7606), .ZN(n7608)
         );
  OAI21_X1 U9263 ( .B1(n7609), .B2(n9621), .A(n7608), .ZN(n7612) );
  MUX2_X1 U9264 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7610), .S(n9623), .Z(n7611)
         );
  AOI211_X1 U9265 ( .C1(n9868), .C2(n7613), .A(n7612), .B(n7611), .ZN(n7614)
         );
  INV_X1 U9266 ( .A(n7614), .ZN(P1_U3289) );
  OAI21_X1 U9267 ( .B1(n4421), .B2(n7617), .A(n7724), .ZN(n10059) );
  NAND2_X1 U9268 ( .A1(n8926), .A2(n7615), .ZN(n8794) );
  AOI22_X1 U9269 ( .A1(n5656), .A2(n8629), .B1(n8627), .B2(n8949), .ZN(n7620)
         );
  XNOR2_X1 U9270 ( .A(n7616), .B(n7617), .ZN(n7618) );
  NAND2_X1 U9271 ( .A1(n7618), .A2(n8952), .ZN(n7619) );
  OAI211_X1 U9272 ( .C1(n10059), .C2(n10051), .A(n7620), .B(n7619), .ZN(n10060) );
  NAND2_X1 U9273 ( .A1(n10060), .A2(n8926), .ZN(n7624) );
  OAI22_X1 U9274 ( .A1(n8926), .A2(n5389), .B1(n7621), .B2(n10021), .ZN(n7622)
         );
  AOI21_X1 U9275 ( .B1(n10062), .B2(n8956), .A(n7622), .ZN(n7623) );
  OAI211_X1 U9276 ( .C1(n10059), .C2(n8794), .A(n7624), .B(n7623), .ZN(
        P2_U3224) );
  INV_X1 U9277 ( .A(n7625), .ZN(n7634) );
  NAND2_X1 U9278 ( .A1(n7626), .A2(n9623), .ZN(n7633) );
  AOI22_X1 U9279 ( .A1(n9617), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7627), .B2(
        n9861), .ZN(n7628) );
  OAI21_X1 U9280 ( .B1(n9865), .B2(n7629), .A(n7628), .ZN(n7630) );
  AOI21_X1 U9281 ( .B1(n7631), .B2(n9858), .A(n7630), .ZN(n7632) );
  OAI211_X1 U9282 ( .C1(n7634), .C2(n9626), .A(n7633), .B(n7632), .ZN(P1_U3288) );
  INV_X1 U9283 ( .A(n7787), .ZN(n7651) );
  AOI22_X1 U9284 ( .A1(n9617), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n9861), .ZN(n7635) );
  OAI21_X1 U9285 ( .B1(n9865), .B2(n7636), .A(n7635), .ZN(n7637) );
  AOI21_X1 U9286 ( .B1(n9858), .B2(n7638), .A(n7637), .ZN(n7641) );
  NAND2_X1 U9287 ( .A1(n7639), .A2(n9623), .ZN(n7640) );
  OAI211_X1 U9288 ( .C1(n7642), .C2(n7651), .A(n7641), .B(n7640), .ZN(P1_U3292) );
  NAND2_X1 U9289 ( .A1(n7643), .A2(n9623), .ZN(n7650) );
  AOI22_X1 U9290 ( .A1(n9617), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7644), .B2(
        n9861), .ZN(n7645) );
  OAI21_X1 U9291 ( .B1(n9865), .B2(n7646), .A(n7645), .ZN(n7647) );
  AOI21_X1 U9292 ( .B1(n7648), .B2(n9858), .A(n7647), .ZN(n7649) );
  OAI211_X1 U9293 ( .C1(n7652), .C2(n7651), .A(n7650), .B(n7649), .ZN(P1_U3286) );
  INV_X1 U9294 ( .A(n7653), .ZN(n7662) );
  INV_X1 U9295 ( .A(n7763), .ZN(n7658) );
  NAND2_X1 U9296 ( .A1(n7654), .A2(n9858), .ZN(n7657) );
  AOI22_X1 U9297 ( .A1(n9617), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7655), .B2(
        n9861), .ZN(n7656) );
  OAI211_X1 U9298 ( .C1(n7658), .C2(n9865), .A(n7657), .B(n7656), .ZN(n7659)
         );
  AOI21_X1 U9299 ( .B1(n7660), .B2(n9623), .A(n7659), .ZN(n7661) );
  OAI21_X1 U9300 ( .B1(n7662), .B2(n9626), .A(n7661), .ZN(P1_U3284) );
  OR2_X1 U9301 ( .A1(n9128), .A2(n9804), .ZN(n8238) );
  NAND2_X1 U9302 ( .A1(n9128), .A2(n9804), .ZN(n8242) );
  NAND2_X1 U9303 ( .A1(n8238), .A2(n8242), .ZN(n7674) );
  INV_X1 U9304 ( .A(n7674), .ZN(n8319) );
  AND2_X1 U9305 ( .A1(n8219), .A2(n7663), .ZN(n8217) );
  OR2_X1 U9306 ( .A1(n8220), .A2(n8217), .ZN(n7664) );
  INV_X1 U9307 ( .A(n7665), .ZN(n8215) );
  NAND2_X1 U9308 ( .A1(n8318), .A2(n7667), .ZN(n8401) );
  OAI21_X1 U9309 ( .B1(n8319), .B2(n7669), .A(n7777), .ZN(n7671) );
  OR2_X1 U9310 ( .A1(n7863), .A2(n9490), .ZN(n7670) );
  OAI21_X1 U9311 ( .B1(n7672), .B2(n9488), .A(n7670), .ZN(n9124) );
  AOI21_X1 U9312 ( .B1(n7671), .B2(n9608), .A(n9124), .ZN(n7685) );
  INV_X1 U9313 ( .A(n7672), .ZN(n9287) );
  OAI21_X1 U9314 ( .B1(n7675), .B2(n7674), .A(n7783), .ZN(n7687) );
  NAND2_X1 U9315 ( .A1(n7687), .A2(n9868), .ZN(n7683) );
  INV_X1 U9316 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7677) );
  INV_X1 U9317 ( .A(n7676), .ZN(n9126) );
  OAI22_X1 U9318 ( .A1(n9623), .A2(n7677), .B1(n9126), .B2(n9544), .ZN(n7681)
         );
  INV_X1 U9319 ( .A(n9128), .ZN(n7689) );
  AND2_X2 U9320 ( .A1(n7679), .A2(n7689), .ZN(n7788) );
  INV_X1 U9321 ( .A(n7788), .ZN(n7790) );
  OAI211_X1 U9322 ( .C1(n7689), .C2(n7679), .A(n7790), .B(n9613), .ZN(n7684)
         );
  NOR2_X1 U9323 ( .A1(n7684), .A2(n9621), .ZN(n7680) );
  AOI211_X1 U9324 ( .C1(n9618), .C2(n9128), .A(n7681), .B(n7680), .ZN(n7682)
         );
  OAI211_X1 U9325 ( .C1(n9617), .C2(n7685), .A(n7683), .B(n7682), .ZN(P1_U3283) );
  NAND2_X1 U9326 ( .A1(n7685), .A2(n7684), .ZN(n7686) );
  AOI21_X1 U9327 ( .B1(n7687), .B2(n9878), .A(n7686), .ZN(n7693) );
  INV_X1 U9328 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7688) );
  OAI22_X1 U9329 ( .A1(n7689), .A2(n9759), .B1(n9890), .B2(n7688), .ZN(n7690)
         );
  INV_X1 U9330 ( .A(n7690), .ZN(n7691) );
  OAI21_X1 U9331 ( .B1(n7693), .B2(n9888), .A(n7691), .ZN(P1_U3483) );
  AOI22_X1 U9332 ( .A1(n9128), .A2(n9695), .B1(n9893), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7692) );
  OAI21_X1 U9333 ( .B1(n7693), .B2(n9893), .A(n7692), .ZN(P1_U3532) );
  INV_X1 U9334 ( .A(n7694), .ZN(n7708) );
  AOI22_X1 U9335 ( .A1(n7695), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n9100), .ZN(n7696) );
  OAI21_X1 U9336 ( .B1(n7708), .B2(n9103), .A(n7696), .ZN(P2_U3274) );
  INV_X1 U9337 ( .A(n7697), .ZN(n9882) );
  OAI21_X1 U9338 ( .B1(n7700), .B2(n7699), .A(n7698), .ZN(n7701) );
  NAND2_X1 U9339 ( .A1(n7701), .A2(n9809), .ZN(n7706) );
  AOI22_X1 U9340 ( .A1(n9802), .A2(n9287), .B1(P1_REG3_REG_8__SCAN_IN), .B2(
        P1_U3086), .ZN(n7702) );
  OAI21_X1 U9341 ( .B1(n7703), .B2(n9803), .A(n7702), .ZN(n7704) );
  AOI21_X1 U9342 ( .B1(n5085), .B2(n9267), .A(n7704), .ZN(n7705) );
  OAI211_X1 U9343 ( .C1(n9882), .C2(n9800), .A(n7706), .B(n7705), .ZN(P1_U3221) );
  OAI222_X1 U9344 ( .A1(n4336), .A2(n7708), .B1(n8338), .B2(P1_U3086), .C1(
        n7707), .C2(n9789), .ZN(P1_U3334) );
  INV_X1 U9345 ( .A(n9824), .ZN(n9857) );
  INV_X1 U9346 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7715) );
  XNOR2_X1 U9347 ( .A(n7958), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n7713) );
  OAI21_X1 U9348 ( .B1(n7711), .B2(n7710), .A(n7709), .ZN(n7712) );
  NAND2_X1 U9349 ( .A1(n7713), .A2(n7712), .ZN(n7956) );
  OAI211_X1 U9350 ( .C1(n7713), .C2(n7712), .A(n9340), .B(n7956), .ZN(n7714)
         );
  NAND2_X1 U9351 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9109) );
  OAI211_X1 U9352 ( .C1(n9857), .C2(n7715), .A(n7714), .B(n9109), .ZN(n7721)
         );
  INV_X1 U9353 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10122) );
  AOI22_X1 U9354 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n7958), .B1(n7963), .B2(
        n10122), .ZN(n7718) );
  AOI211_X1 U9355 ( .C1(n7719), .C2(n7718), .A(n7962), .B(n9343), .ZN(n7720)
         );
  AOI211_X1 U9356 ( .C1(n9332), .C2(n7963), .A(n7721), .B(n7720), .ZN(n7722)
         );
  INV_X1 U9357 ( .A(n7722), .ZN(P1_U3257) );
  NAND2_X1 U9358 ( .A1(n7724), .A2(n7723), .ZN(n7725) );
  XNOR2_X1 U9359 ( .A(n7725), .B(n7726), .ZN(n10064) );
  XOR2_X1 U9360 ( .A(n7727), .B(n7726), .Z(n7728) );
  NAND2_X1 U9361 ( .A1(n7728), .A2(n8952), .ZN(n7730) );
  AOI22_X1 U9362 ( .A1(n8626), .A2(n8949), .B1(n5656), .B2(n8628), .ZN(n7729)
         );
  OAI211_X1 U9363 ( .C1(n10064), .C2(n10051), .A(n7730), .B(n7729), .ZN(n10065) );
  NAND2_X1 U9364 ( .A1(n10065), .A2(n8926), .ZN(n7735) );
  OAI22_X1 U9365 ( .A1(n8926), .A2(n7732), .B1(n7731), .B2(n10021), .ZN(n7733)
         );
  AOI21_X1 U9366 ( .B1(n10067), .B2(n8956), .A(n7733), .ZN(n7734) );
  OAI211_X1 U9367 ( .C1(n10064), .C2(n8794), .A(n7735), .B(n7734), .ZN(
        P2_U3223) );
  NAND2_X1 U9368 ( .A1(n7745), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7736) );
  XNOR2_X1 U9369 ( .A(n7832), .B(n7845), .ZN(n7738) );
  AOI21_X1 U9370 ( .B1(n7738), .B2(n5425), .A(n7835), .ZN(n7754) );
  MUX2_X1 U9371 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8643), .Z(n7846) );
  XNOR2_X1 U9372 ( .A(n7846), .B(n7834), .ZN(n7743) );
  OR2_X1 U9373 ( .A1(n7739), .A2(n7745), .ZN(n7741) );
  OAI21_X1 U9374 ( .B1(n7743), .B2(n7742), .A(n7847), .ZN(n7752) );
  AND2_X1 U9375 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7804) );
  AOI21_X1 U9376 ( .B1(n9962), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7804), .ZN(
        n7744) );
  OAI21_X1 U9377 ( .B1(n7845), .B2(n9958), .A(n7744), .ZN(n7751) );
  NAND2_X1 U9378 ( .A1(n7745), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7746) );
  NOR2_X1 U9379 ( .A1(n5428), .A2(n7748), .ZN(n7826) );
  AOI21_X1 U9380 ( .B1(n5428), .B2(n7748), .A(n7826), .ZN(n7749) );
  NOR2_X1 U9381 ( .A1(n7749), .A2(n9980), .ZN(n7750) );
  AOI211_X1 U9382 ( .C1(n9949), .C2(n7752), .A(n7751), .B(n7750), .ZN(n7753)
         );
  OAI21_X1 U9383 ( .B1(n7754), .B2(n10005), .A(n7753), .ZN(P2_U3193) );
  XOR2_X1 U9384 ( .A(n7755), .B(n7756), .Z(n7765) );
  NOR2_X1 U9385 ( .A1(n9814), .A2(n7757), .ZN(n7762) );
  INV_X1 U9386 ( .A(n9804), .ZN(n9286) );
  NAND2_X1 U9387 ( .A1(n9802), .A2(n9286), .ZN(n7759) );
  OAI211_X1 U9388 ( .C1(n7760), .C2(n9803), .A(n7759), .B(n7758), .ZN(n7761)
         );
  AOI211_X1 U9389 ( .C1(n7763), .C2(n6649), .A(n7762), .B(n7761), .ZN(n7764)
         );
  OAI21_X1 U9390 ( .B1(n7765), .B2(n9245), .A(n7764), .ZN(P1_U3231) );
  XNOR2_X1 U9391 ( .A(n7816), .B(n4329), .ZN(n7807) );
  AND2_X1 U9392 ( .A1(n7807), .A2(n8626), .ZN(n7769) );
  XNOR2_X1 U9393 ( .A(n10079), .B(n8491), .ZN(n7876) );
  XNOR2_X1 U9394 ( .A(n7876), .B(n8625), .ZN(n7770) );
  XNOR2_X1 U9395 ( .A(n7878), .B(n7770), .ZN(n7776) );
  INV_X1 U9396 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7771) );
  OR2_X1 U9397 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7771), .ZN(n7831) );
  OAI21_X1 U9398 ( .B1(n7894), .B2(n8574), .A(n7831), .ZN(n7772) );
  AOI21_X1 U9399 ( .B1(n8571), .B2(n8624), .A(n7772), .ZN(n7773) );
  OAI21_X1 U9400 ( .B1(n7895), .B2(n8608), .A(n7773), .ZN(n7774) );
  AOI21_X1 U9401 ( .B1(n10079), .B2(n8615), .A(n7774), .ZN(n7775) );
  OAI21_X1 U9402 ( .B1(n7776), .B2(n8610), .A(n7775), .ZN(P2_U3164) );
  NAND2_X1 U9403 ( .A1(n7864), .A2(n7863), .ZN(n8243) );
  NAND2_X1 U9404 ( .A1(n8236), .A2(n8243), .ZN(n7784) );
  INV_X1 U9405 ( .A(n7784), .ZN(n8320) );
  OAI211_X1 U9406 ( .C1(n7778), .C2(n8320), .A(n7856), .B(n9608), .ZN(n7780)
         );
  AOI22_X1 U9407 ( .A1(n9286), .A2(n9523), .B1(n9524), .B2(n9284), .ZN(n7779)
         );
  NAND2_X1 U9408 ( .A1(n7780), .A2(n7779), .ZN(n7797) );
  INV_X1 U9409 ( .A(n7797), .ZN(n7796) );
  NOR2_X1 U9410 ( .A1(n9617), .A2(n7781), .ZN(n7786) );
  OAI21_X1 U9411 ( .B1(n7785), .B2(n7784), .A(n7866), .ZN(n7799) );
  OAI21_X1 U9412 ( .B1(n7787), .B2(n7786), .A(n7799), .ZN(n7795) );
  INV_X1 U9413 ( .A(n7864), .ZN(n9801) );
  INV_X1 U9414 ( .A(n7862), .ZN(n7789) );
  AOI211_X1 U9415 ( .C1(n7864), .C2(n7790), .A(n9595), .B(n7789), .ZN(n7798)
         );
  AOI22_X1 U9416 ( .A1(n9617), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7791), .B2(
        n9861), .ZN(n7792) );
  OAI21_X1 U9417 ( .B1(n9801), .B2(n9865), .A(n7792), .ZN(n7793) );
  AOI21_X1 U9418 ( .B1(n7798), .B2(n9858), .A(n7793), .ZN(n7794) );
  OAI211_X1 U9419 ( .C1(n9617), .C2(n7796), .A(n7795), .B(n7794), .ZN(P1_U3282) );
  AOI211_X1 U9420 ( .C1(n7799), .C2(n9878), .A(n7798), .B(n7797), .ZN(n7802)
         );
  AOI22_X1 U9421 ( .A1(n7864), .A2(n9695), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n9893), .ZN(n7800) );
  OAI21_X1 U9422 ( .B1(n7802), .B2(n9893), .A(n7800), .ZN(P1_U3533) );
  AOI22_X1 U9423 ( .A1(n7864), .A2(n9769), .B1(P1_REG0_REG_11__SCAN_IN), .B2(
        n9888), .ZN(n7801) );
  OAI21_X1 U9424 ( .B1(n7802), .B2(n9888), .A(n7801), .ZN(P1_U3486) );
  NOR2_X1 U9425 ( .A1(n7877), .A2(n8603), .ZN(n7803) );
  AOI211_X1 U9426 ( .C1(n8606), .C2(n8627), .A(n7804), .B(n7803), .ZN(n7805)
         );
  OAI21_X1 U9427 ( .B1(n7820), .B2(n8608), .A(n7805), .ZN(n7810) );
  AOI211_X1 U9428 ( .C1(n7808), .C2(n7807), .A(n8610), .B(n7806), .ZN(n7809)
         );
  AOI211_X1 U9429 ( .C1(n10072), .C2(n8615), .A(n7810), .B(n7809), .ZN(n7811)
         );
  INV_X1 U9430 ( .A(n7811), .ZN(P2_U3176) );
  INV_X1 U9431 ( .A(n7812), .ZN(n7854) );
  AOI22_X1 U9432 ( .A1(n7813), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n9100), .ZN(n7814) );
  OAI21_X1 U9433 ( .B1(n7854), .B2(n8046), .A(n7814), .ZN(P2_U3273) );
  XNOR2_X1 U9434 ( .A(n7815), .B(n7816), .ZN(n10069) );
  XNOR2_X1 U9435 ( .A(n7817), .B(n7816), .ZN(n7818) );
  OAI222_X1 U9436 ( .A1(n10030), .A2(n7877), .B1(n10028), .B2(n7819), .C1(
        n7818), .C2(n10026), .ZN(n10070) );
  NAND2_X1 U9437 ( .A1(n10070), .A2(n8926), .ZN(n7823) );
  OAI22_X1 U9438 ( .A1(n8926), .A2(n5428), .B1(n7820), .B2(n10021), .ZN(n7821)
         );
  AOI21_X1 U9439 ( .B1(n10072), .B2(n8956), .A(n7821), .ZN(n7822) );
  OAI211_X1 U9440 ( .C1(n8959), .C2(n10069), .A(n7823), .B(n7822), .ZN(
        P2_U3222) );
  NOR2_X1 U9441 ( .A1(n7834), .A2(n7825), .ZN(n7827) );
  NAND2_X1 U9442 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n7949), .ZN(n7828) );
  OAI21_X1 U9443 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7949), .A(n7828), .ZN(
        n7829) );
  AOI21_X1 U9444 ( .B1(n7830), .B2(n7829), .A(n7948), .ZN(n7853) );
  INV_X1 U9445 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n8086) );
  OAI21_X1 U9446 ( .B1(n10017), .B2(n8086), .A(n7831), .ZN(n7842) );
  INV_X1 U9447 ( .A(n7832), .ZN(n7833) );
  NOR2_X1 U9448 ( .A1(n7834), .A2(n7833), .ZN(n7836) );
  NAND2_X1 U9449 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n7949), .ZN(n7837) );
  OAI21_X1 U9450 ( .B1(n7949), .B2(P2_REG1_REG_12__SCAN_IN), .A(n7837), .ZN(
        n7838) );
  AOI21_X1 U9451 ( .B1(n7839), .B2(n7838), .A(n7934), .ZN(n7840) );
  NOR2_X1 U9452 ( .A1(n7840), .A2(n10005), .ZN(n7841) );
  AOI211_X1 U9453 ( .C1(n10003), .C2(n7843), .A(n7842), .B(n7841), .ZN(n7852)
         );
  MUX2_X1 U9454 ( .A(n5446), .B(n5442), .S(n8643), .Z(n7844) );
  NOR2_X1 U9455 ( .A1(n7844), .A2(n7843), .ZN(n7937) );
  AND2_X1 U9456 ( .A1(n7844), .A2(n7843), .ZN(n7940) );
  NOR2_X1 U9457 ( .A1(n7937), .A2(n7940), .ZN(n7849) );
  OR2_X1 U9458 ( .A1(n7846), .A2(n7845), .ZN(n7848) );
  XNOR2_X1 U9459 ( .A(n7849), .B(n7939), .ZN(n7850) );
  NAND2_X1 U9460 ( .A1(n7850), .A2(n9949), .ZN(n7851) );
  OAI211_X1 U9461 ( .C1(n7853), .C2(n9980), .A(n7852), .B(n7851), .ZN(P2_U3194) );
  OAI222_X1 U9462 ( .A1(n9789), .A2(n7855), .B1(n4336), .B2(n7854), .C1(
        P1_U3086), .C2(n8193), .ZN(P1_U3333) );
  NAND2_X1 U9463 ( .A1(n9169), .A2(n9284), .ZN(n8237) );
  NAND2_X1 U9464 ( .A1(n7909), .A2(n9805), .ZN(n8244) );
  NAND2_X1 U9465 ( .A1(n8237), .A2(n8244), .ZN(n7867) );
  INV_X1 U9466 ( .A(n7867), .ZN(n8322) );
  OAI211_X1 U9467 ( .C1(n8322), .C2(n4598), .A(n7915), .B(n9608), .ZN(n7860)
         );
  OR2_X1 U9468 ( .A1(n7863), .A2(n9488), .ZN(n7859) );
  NAND2_X1 U9469 ( .A1(n9283), .A2(n9524), .ZN(n7858) );
  AND2_X1 U9470 ( .A1(n7859), .A2(n7858), .ZN(n9164) );
  NAND2_X1 U9471 ( .A1(n7860), .A2(n9164), .ZN(n7884) );
  INV_X1 U9472 ( .A(n7921), .ZN(n7861) );
  AOI211_X1 U9473 ( .C1(n7909), .C2(n7862), .A(n9595), .B(n7861), .ZN(n7887)
         );
  NOR2_X1 U9474 ( .A1(n7884), .A2(n7887), .ZN(n7875) );
  INV_X1 U9475 ( .A(n7863), .ZN(n9285) );
  OAI21_X1 U9476 ( .B1(n7868), .B2(n7867), .A(n7911), .ZN(n7885) );
  NAND2_X1 U9477 ( .A1(n7885), .A2(n7869), .ZN(n7871) );
  AOI22_X1 U9478 ( .A1(n7909), .A2(n9769), .B1(P1_REG0_REG_12__SCAN_IN), .B2(
        n9888), .ZN(n7870) );
  OAI211_X1 U9479 ( .C1(n7875), .C2(n9888), .A(n7871), .B(n7870), .ZN(P1_U3489) );
  NAND2_X1 U9480 ( .A1(n7885), .A2(n7872), .ZN(n7874) );
  AOI22_X1 U9481 ( .A1(n7909), .A2(n9695), .B1(P1_REG1_REG_12__SCAN_IN), .B2(
        n9893), .ZN(n7873) );
  OAI211_X1 U9482 ( .C1(n7875), .C2(n9893), .A(n7874), .B(n7873), .ZN(P1_U3534) );
  XNOR2_X1 U9483 ( .A(n8016), .B(n8491), .ZN(n7969) );
  XNOR2_X1 U9484 ( .A(n7969), .B(n7893), .ZN(n7970) );
  XNOR2_X1 U9485 ( .A(n7971), .B(n7970), .ZN(n7883) );
  NAND2_X1 U9486 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7936) );
  OAI21_X1 U9487 ( .B1(n7972), .B2(n8603), .A(n7936), .ZN(n7879) );
  AOI21_X1 U9488 ( .B1(n8606), .B2(n8625), .A(n7879), .ZN(n7880) );
  OAI21_X1 U9489 ( .B1(n8004), .B2(n8608), .A(n7880), .ZN(n7881) );
  AOI21_X1 U9490 ( .B1(n8016), .B2(n8615), .A(n7881), .ZN(n7882) );
  OAI21_X1 U9491 ( .B1(n7883), .B2(n8610), .A(n7882), .ZN(P2_U3174) );
  AOI21_X1 U9492 ( .B1(n9166), .B2(n9861), .A(n7884), .ZN(n7890) );
  NAND2_X1 U9493 ( .A1(n7885), .A2(n9868), .ZN(n7889) );
  OAI22_X1 U9494 ( .A1(n9169), .A2(n9865), .B1(n7463), .B2(n9623), .ZN(n7886)
         );
  AOI21_X1 U9495 ( .B1(n7887), .B2(n9858), .A(n7886), .ZN(n7888) );
  OAI211_X1 U9496 ( .C1(n9617), .C2(n7890), .A(n7889), .B(n7888), .ZN(P1_U3281) );
  XNOR2_X1 U9497 ( .A(n7891), .B(n7897), .ZN(n7892) );
  OAI222_X1 U9498 ( .A1(n10028), .A2(n7894), .B1(n10030), .B2(n7893), .C1(
        n10026), .C2(n7892), .ZN(n10077) );
  INV_X1 U9499 ( .A(n10077), .ZN(n7901) );
  OAI22_X1 U9500 ( .A1(n8926), .A2(n5446), .B1(n7895), .B2(n10021), .ZN(n7896)
         );
  AOI21_X1 U9501 ( .B1(n10079), .B2(n8956), .A(n7896), .ZN(n7900) );
  NAND2_X1 U9502 ( .A1(n7898), .A2(n7897), .ZN(n10074) );
  NAND3_X1 U9503 ( .A1(n10076), .A2(n10074), .A3(n8914), .ZN(n7899) );
  OAI211_X1 U9504 ( .C1(n7901), .C2(n10034), .A(n7900), .B(n7899), .ZN(
        P2_U3221) );
  INV_X1 U9505 ( .A(n7906), .ZN(n7904) );
  NAND2_X1 U9506 ( .A1(n9100), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7903) );
  OAI211_X1 U9507 ( .C1(n7904), .C2(n9103), .A(n7903), .B(n7902), .ZN(P2_U3272) );
  NAND2_X1 U9508 ( .A1(n7906), .A2(n7905), .ZN(n7907) );
  OAI211_X1 U9509 ( .C1(n7908), .C2(n9789), .A(n7907), .B(n8448), .ZN(P1_U3332) );
  NAND2_X1 U9510 ( .A1(n9225), .A2(n9283), .ZN(n8408) );
  OAI21_X1 U9511 ( .B1(n7912), .B2(n8324), .A(n8140), .ZN(n7929) );
  INV_X1 U9512 ( .A(n7929), .ZN(n7926) );
  NAND2_X1 U9513 ( .A1(n7915), .A2(n8237), .ZN(n7917) );
  INV_X1 U9514 ( .A(n8237), .ZN(n7913) );
  NOR2_X1 U9515 ( .A1(n8324), .A2(n7913), .ZN(n7914) );
  INV_X1 U9516 ( .A(n9605), .ZN(n7916) );
  AOI21_X1 U9517 ( .B1(n8324), .B2(n7917), .A(n7916), .ZN(n7920) );
  NAND2_X1 U9518 ( .A1(n9284), .A2(n9523), .ZN(n7919) );
  NAND2_X1 U9519 ( .A1(n9282), .A2(n9524), .ZN(n7918) );
  AND2_X1 U9520 ( .A1(n7919), .A2(n7918), .ZN(n9220) );
  OAI21_X1 U9521 ( .B1(n7920), .B2(n9592), .A(n9220), .ZN(n7927) );
  AOI211_X1 U9522 ( .C1(n8137), .C2(n7921), .A(n9595), .B(n4420), .ZN(n7928)
         );
  NAND2_X1 U9523 ( .A1(n7928), .A2(n9858), .ZN(n7923) );
  AOI22_X1 U9524 ( .A1(n9617), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9222), .B2(
        n9861), .ZN(n7922) );
  OAI211_X1 U9525 ( .C1(n9225), .C2(n9865), .A(n7923), .B(n7922), .ZN(n7924)
         );
  AOI21_X1 U9526 ( .B1(n7927), .B2(n9623), .A(n7924), .ZN(n7925) );
  OAI21_X1 U9527 ( .B1(n7926), .B2(n9626), .A(n7925), .ZN(P1_U3280) );
  AOI211_X1 U9528 ( .C1(n7929), .C2(n9878), .A(n7928), .B(n7927), .ZN(n7933)
         );
  AOI22_X1 U9529 ( .A1(n8137), .A2(n9769), .B1(P1_REG0_REG_13__SCAN_IN), .B2(
        n9888), .ZN(n7930) );
  OAI21_X1 U9530 ( .B1(n7933), .B2(n9888), .A(n7930), .ZN(P1_U3492) );
  NAND2_X1 U9531 ( .A1(n9893), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7932) );
  NAND2_X1 U9532 ( .A1(n8137), .A2(n9695), .ZN(n7931) );
  OAI211_X1 U9533 ( .C1(n7933), .C2(n9893), .A(n7932), .B(n7931), .ZN(P1_U3535) );
  INV_X1 U9534 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8012) );
  AOI21_X1 U9535 ( .B1(n8012), .B2(n7935), .A(n8637), .ZN(n7955) );
  INV_X1 U9536 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8089) );
  OAI21_X1 U9537 ( .B1(n10017), .B2(n8089), .A(n7936), .ZN(n7947) );
  INV_X1 U9538 ( .A(n7937), .ZN(n7938) );
  MUX2_X1 U9539 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8643), .Z(n7941) );
  NOR2_X1 U9540 ( .A1(n7941), .A2(n7950), .ZN(n8647) );
  AOI21_X1 U9541 ( .B1(n7941), .B2(n7950), .A(n8647), .ZN(n7942) );
  INV_X1 U9542 ( .A(n7942), .ZN(n7943) );
  NOR2_X1 U9543 ( .A1(n7944), .A2(n7943), .ZN(n8646) );
  AOI21_X1 U9544 ( .B1(n7944), .B2(n7943), .A(n8646), .ZN(n7945) );
  NOR2_X1 U9545 ( .A1(n7945), .A2(n10013), .ZN(n7946) );
  AOI211_X1 U9546 ( .C1(n10003), .C2(n8655), .A(n7947), .B(n7946), .ZN(n7954)
         );
  AOI21_X1 U9547 ( .B1(n5465), .B2(n7951), .A(n8656), .ZN(n7952) );
  OR2_X1 U9548 ( .A1(n7952), .A2(n9980), .ZN(n7953) );
  OAI211_X1 U9549 ( .C1(n7955), .C2(n10005), .A(n7954), .B(n7953), .ZN(
        P2_U3195) );
  INV_X1 U9550 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7961) );
  INV_X1 U9551 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7957) );
  OAI21_X1 U9552 ( .B1(n7958), .B2(n7957), .A(n7956), .ZN(n8118) );
  XNOR2_X1 U9553 ( .A(n8103), .B(n8118), .ZN(n7959) );
  NAND2_X1 U9554 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n7959), .ZN(n8120) );
  OAI211_X1 U9555 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n7959), .A(n9340), .B(
        n8120), .ZN(n7960) );
  NAND2_X1 U9556 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9264) );
  OAI211_X1 U9557 ( .C1(n9857), .C2(n7961), .A(n7960), .B(n9264), .ZN(n7967)
         );
  INV_X1 U9558 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7965) );
  XOR2_X1 U9559 ( .A(n8119), .B(n8104), .Z(n7964) );
  AOI211_X1 U9560 ( .C1(n7965), .C2(n7964), .A(n8105), .B(n9343), .ZN(n7966)
         );
  AOI211_X1 U9561 ( .C1(n9332), .C2(n8119), .A(n7967), .B(n7966), .ZN(n7968)
         );
  INV_X1 U9562 ( .A(n7968), .ZN(P1_U3258) );
  INV_X1 U9563 ( .A(n8024), .ZN(n7981) );
  XNOR2_X1 U9564 ( .A(n8491), .B(n8024), .ZN(n8461) );
  XNOR2_X1 U9565 ( .A(n8461), .B(n7972), .ZN(n7973) );
  OAI21_X1 U9566 ( .B1(n7974), .B2(n7973), .A(n8463), .ZN(n7975) );
  NAND2_X1 U9567 ( .A1(n7975), .A2(n8588), .ZN(n7980) );
  NAND2_X1 U9568 ( .A1(n8948), .A2(n8571), .ZN(n7976) );
  NAND2_X1 U9569 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8642) );
  NAND2_X1 U9570 ( .A1(n7976), .A2(n8642), .ZN(n7978) );
  NOR2_X1 U9571 ( .A1(n8608), .A2(n7997), .ZN(n7977) );
  AOI211_X1 U9572 ( .C1(n8606), .C2(n8624), .A(n7978), .B(n7977), .ZN(n7979)
         );
  OAI211_X1 U9573 ( .C1(n7981), .C2(n8596), .A(n7980), .B(n7979), .ZN(P2_U3155) );
  INV_X1 U9574 ( .A(n7982), .ZN(n7987) );
  AOI22_X1 U9575 ( .A1(n7983), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n9100), .ZN(n7984) );
  OAI21_X1 U9576 ( .B1(n7987), .B2(n8046), .A(n7984), .ZN(P2_U3271) );
  OAI222_X1 U9577 ( .A1(n4336), .A2(n7987), .B1(n7986), .B2(P1_U3086), .C1(
        n7985), .C2(n9789), .ZN(P1_U3331) );
  INV_X1 U9578 ( .A(n10023), .ZN(n7994) );
  INV_X1 U9579 ( .A(n7995), .ZN(n7988) );
  XNOR2_X1 U9580 ( .A(n7989), .B(n7988), .ZN(n7990) );
  NAND2_X1 U9581 ( .A1(n7990), .A2(n8952), .ZN(n7992) );
  AOI22_X1 U9582 ( .A1(n5656), .A2(n8624), .B1(n8948), .B2(n8949), .ZN(n7991)
         );
  INV_X1 U9583 ( .A(n8023), .ZN(n7993) );
  AOI21_X1 U9584 ( .B1(n7994), .B2(n8024), .A(n7993), .ZN(n8001) );
  XNOR2_X1 U9585 ( .A(n7996), .B(n7995), .ZN(n8025) );
  OAI22_X1 U9586 ( .A1(n8926), .A2(n7998), .B1(n7997), .B2(n10021), .ZN(n7999)
         );
  AOI21_X1 U9587 ( .B1(n8025), .B2(n8914), .A(n7999), .ZN(n8000) );
  OAI21_X1 U9588 ( .B1(n8001), .B2(n10034), .A(n8000), .ZN(P2_U3219) );
  XOR2_X1 U9589 ( .A(n8009), .B(n8002), .Z(n8003) );
  AOI222_X1 U9590 ( .A1(n8952), .A2(n8003), .B1(n8623), .B2(n8949), .C1(n8625), 
        .C2(n5656), .ZN(n8015) );
  INV_X1 U9591 ( .A(n8015), .ZN(n8007) );
  OAI22_X1 U9592 ( .A1(n8005), .A2(n10023), .B1(n8004), .B2(n10021), .ZN(n8006) );
  OAI21_X1 U9593 ( .B1(n8007), .B2(n8006), .A(n8926), .ZN(n8011) );
  XOR2_X1 U9594 ( .A(n8009), .B(n8008), .Z(n8017) );
  AOI22_X1 U9595 ( .A1(n8017), .A2(n8914), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n10034), .ZN(n8010) );
  NAND2_X1 U9596 ( .A1(n8011), .A2(n8010), .ZN(P2_U3220) );
  MUX2_X1 U9597 ( .A(n8012), .B(n8015), .S(n10096), .Z(n8014) );
  INV_X1 U9598 ( .A(n9009), .ZN(n8984) );
  AOI22_X1 U9599 ( .A1(n8017), .A2(n8984), .B1(n9006), .B2(n8016), .ZN(n8013)
         );
  NAND2_X1 U9600 ( .A1(n8014), .A2(n8013), .ZN(P2_U3472) );
  MUX2_X1 U9601 ( .A(n5464), .B(n8015), .S(n10081), .Z(n8019) );
  INV_X1 U9602 ( .A(n9083), .ZN(n9048) );
  AOI22_X1 U9603 ( .A1(n8017), .A2(n9048), .B1(n9079), .B2(n8016), .ZN(n8018)
         );
  NAND2_X1 U9604 ( .A1(n8019), .A2(n8018), .ZN(P2_U3429) );
  MUX2_X1 U9605 ( .A(n8020), .B(n8023), .S(n10081), .Z(n8022) );
  AOI22_X1 U9606 ( .A1(n8025), .A2(n9048), .B1(n9079), .B2(n8024), .ZN(n8021)
         );
  NAND2_X1 U9607 ( .A1(n8022), .A2(n8021), .ZN(P2_U3432) );
  MUX2_X1 U9608 ( .A(n10138), .B(n8023), .S(n10096), .Z(n8027) );
  AOI22_X1 U9609 ( .A1(n8025), .A2(n8984), .B1(n9006), .B2(n8024), .ZN(n8026)
         );
  NAND2_X1 U9610 ( .A1(n8027), .A2(n8026), .ZN(P2_U3473) );
  INV_X1 U9611 ( .A(n8028), .ZN(n8033) );
  AOI22_X1 U9612 ( .A1(n8029), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n9100), .ZN(n8030) );
  OAI21_X1 U9613 ( .B1(n8033), .B2(n8046), .A(n8030), .ZN(P2_U3270) );
  OAI222_X1 U9614 ( .A1(n4336), .A2(n8033), .B1(n8032), .B2(P1_U3086), .C1(
        n8031), .C2(n9789), .ZN(P1_U3330) );
  XNOR2_X1 U9615 ( .A(n8034), .B(n8036), .ZN(n8035) );
  AOI222_X1 U9616 ( .A1(n8952), .A2(n8035), .B1(n8623), .B2(n5656), .C1(n8938), 
        .C2(n8949), .ZN(n8048) );
  MUX2_X1 U9617 ( .A(n8667), .B(n8048), .S(n10096), .Z(n8039) );
  XNOR2_X1 U9618 ( .A(n8037), .B(n8036), .ZN(n8047) );
  AOI22_X1 U9619 ( .A1(n8047), .A2(n8984), .B1(n9006), .B2(n8616), .ZN(n8038)
         );
  NAND2_X1 U9620 ( .A1(n8039), .A2(n8038), .ZN(P2_U3474) );
  MUX2_X1 U9621 ( .A(n8040), .B(n8048), .S(n10081), .Z(n8042) );
  AOI22_X1 U9622 ( .A1(n8047), .A2(n9048), .B1(n9079), .B2(n8616), .ZN(n8041)
         );
  NAND2_X1 U9623 ( .A1(n8042), .A2(n8041), .ZN(P2_U3435) );
  INV_X1 U9624 ( .A(n8043), .ZN(n8056) );
  AOI22_X1 U9625 ( .A1(n8044), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n9100), .ZN(n8045) );
  OAI21_X1 U9626 ( .B1(n8056), .B2(n8046), .A(n8045), .ZN(P2_U3269) );
  INV_X1 U9627 ( .A(n8047), .ZN(n8053) );
  MUX2_X1 U9628 ( .A(n8049), .B(n8048), .S(n8926), .Z(n8052) );
  INV_X1 U9629 ( .A(n8609), .ZN(n8050) );
  AOI22_X1 U9630 ( .A1(n8616), .A2(n8956), .B1(n8955), .B2(n8050), .ZN(n8051)
         );
  OAI211_X1 U9631 ( .C1(n8053), .C2(n8959), .A(n8052), .B(n8051), .ZN(P2_U3218) );
  OAI222_X1 U9632 ( .A1(n4336), .A2(n8056), .B1(n8055), .B2(P1_U3086), .C1(
        n8054), .C2(n9789), .ZN(P1_U3329) );
  OAI222_X1 U9633 ( .A1(n9789), .A2(n8058), .B1(n4336), .B2(n8057), .C1(
        P1_U3086), .C2(n6047), .ZN(P1_U3336) );
  INV_X1 U9634 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n10278) );
  INV_X1 U9635 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9856) );
  NOR2_X1 U9636 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n8097) );
  INV_X1 U9637 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8669) );
  NOR2_X1 U9638 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n8094) );
  NOR2_X1 U9639 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n8092) );
  NOR2_X1 U9640 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n8088) );
  NOR2_X1 U9641 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n8085) );
  NOR2_X1 U9642 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n8082) );
  NOR2_X1 U9643 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n8078) );
  NOR2_X1 U9644 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n8074) );
  INV_X1 U9645 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9994) );
  NOR2_X1 U9646 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n8070) );
  NOR2_X1 U9647 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n8068) );
  NOR2_X1 U9648 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n8066) );
  NAND2_X1 U9649 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n8064) );
  XOR2_X1 U9650 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10321) );
  NAND2_X1 U9651 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n8062) );
  AOI21_X1 U9652 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10098) );
  INV_X1 U9653 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9296) );
  NAND2_X1 U9654 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n8059) );
  NOR2_X1 U9655 ( .A1(n9296), .A2(n8059), .ZN(n10097) );
  NOR2_X1 U9656 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10097), .ZN(n8060) );
  NOR2_X1 U9657 ( .A1(n10098), .A2(n8060), .ZN(n10319) );
  XOR2_X1 U9658 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10318) );
  NAND2_X1 U9659 ( .A1(n10319), .A2(n10318), .ZN(n8061) );
  NAND2_X1 U9660 ( .A1(n8062), .A2(n8061), .ZN(n10320) );
  NAND2_X1 U9661 ( .A1(n10321), .A2(n10320), .ZN(n8063) );
  NAND2_X1 U9662 ( .A1(n8064), .A2(n8063), .ZN(n10323) );
  XNOR2_X1 U9663 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10322) );
  NOR2_X1 U9664 ( .A1(n10323), .A2(n10322), .ZN(n8065) );
  NOR2_X1 U9665 ( .A1(n8066), .A2(n8065), .ZN(n10311) );
  XNOR2_X1 U9666 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10310) );
  NOR2_X1 U9667 ( .A1(n10311), .A2(n10310), .ZN(n8067) );
  NOR2_X1 U9668 ( .A1(n8068), .A2(n8067), .ZN(n10309) );
  XNOR2_X1 U9669 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10308) );
  NOR2_X1 U9670 ( .A1(n10309), .A2(n10308), .ZN(n8069) );
  NOR2_X1 U9671 ( .A1(n8070), .A2(n8069), .ZN(n10315) );
  AOI22_X1 U9672 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10288), .B1(
        P1_ADDR_REG_7__SCAN_IN), .B2(n9994), .ZN(n10314) );
  NOR2_X1 U9673 ( .A1(n10315), .A2(n10314), .ZN(n8071) );
  AOI21_X1 U9674 ( .B1(n9994), .B2(n10288), .A(n8071), .ZN(n10317) );
  INV_X1 U9675 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n8072) );
  INV_X1 U9676 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10018) );
  AOI22_X1 U9677 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n8072), .B1(
        P1_ADDR_REG_8__SCAN_IN), .B2(n10018), .ZN(n10316) );
  NOR2_X1 U9678 ( .A1(n10317), .A2(n10316), .ZN(n8073) );
  NOR2_X1 U9679 ( .A1(n8074), .A2(n8073), .ZN(n10313) );
  INV_X1 U9680 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n8076) );
  AOI22_X1 U9681 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n8076), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n8075), .ZN(n10312) );
  NOR2_X1 U9682 ( .A1(n10313), .A2(n10312), .ZN(n8077) );
  NOR2_X1 U9683 ( .A1(n8078), .A2(n8077), .ZN(n10118) );
  INV_X1 U9684 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n8080) );
  AOI22_X1 U9685 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n8080), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n8079), .ZN(n10117) );
  NOR2_X1 U9686 ( .A1(n10118), .A2(n10117), .ZN(n8081) );
  NOR2_X1 U9687 ( .A1(n8082), .A2(n8081), .ZN(n10116) );
  INV_X1 U9688 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n8083) );
  INV_X1 U9689 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10252) );
  AOI22_X1 U9690 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n8083), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n10252), .ZN(n10115) );
  NOR2_X1 U9691 ( .A1(n10116), .A2(n10115), .ZN(n8084) );
  NOR2_X1 U9692 ( .A1(n8085), .A2(n8084), .ZN(n10114) );
  INV_X1 U9693 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9840) );
  AOI22_X1 U9694 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n9840), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n8086), .ZN(n10113) );
  NOR2_X1 U9695 ( .A1(n10114), .A2(n10113), .ZN(n8087) );
  NOR2_X1 U9696 ( .A1(n8088), .A2(n8087), .ZN(n10112) );
  INV_X1 U9697 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n8090) );
  AOI22_X1 U9698 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n8090), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n8089), .ZN(n10111) );
  NOR2_X1 U9699 ( .A1(n10112), .A2(n10111), .ZN(n8091) );
  NOR2_X1 U9700 ( .A1(n8092), .A2(n8091), .ZN(n10110) );
  INV_X1 U9701 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n10269) );
  AOI22_X1 U9702 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n7715), .B1(
        P1_ADDR_REG_14__SCAN_IN), .B2(n10269), .ZN(n10109) );
  NOR2_X1 U9703 ( .A1(n10110), .A2(n10109), .ZN(n8093) );
  NOR2_X1 U9704 ( .A1(n8094), .A2(n8093), .ZN(n10108) );
  AOI22_X1 U9705 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n7961), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n8669), .ZN(n10107) );
  NOR2_X1 U9706 ( .A1(n10108), .A2(n10107), .ZN(n8095) );
  AOI21_X1 U9707 ( .B1(n8669), .B2(n7961), .A(n8095), .ZN(n10106) );
  XNOR2_X1 U9708 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10105) );
  NOR2_X1 U9709 ( .A1(n10106), .A2(n10105), .ZN(n8096) );
  NOR2_X1 U9710 ( .A1(n8097), .A2(n8096), .ZN(n10104) );
  AOI22_X1 U9711 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n9856), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n10278), .ZN(n10103) );
  NOR2_X1 U9712 ( .A1(n10104), .A2(n10103), .ZN(n8098) );
  AOI21_X1 U9713 ( .B1(n10278), .B2(n9856), .A(n8098), .ZN(n8099) );
  AND2_X1 U9714 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n8099), .ZN(n10100) );
  NOR2_X1 U9715 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10100), .ZN(n8100) );
  NOR2_X1 U9716 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n8099), .ZN(n10101) );
  NOR2_X1 U9717 ( .A1(n8100), .A2(n10101), .ZN(n8102) );
  XNOR2_X1 U9718 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n8101) );
  XNOR2_X1 U9719 ( .A(n8102), .B(n8101), .ZN(ADD_1068_U4) );
  NOR2_X1 U9720 ( .A1(n8104), .A2(n8103), .ZN(n8106) );
  INV_X1 U9721 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n8107) );
  OR2_X1 U9722 ( .A1(n9331), .A2(n8107), .ZN(n8109) );
  NAND2_X1 U9723 ( .A1(n9331), .A2(n8107), .ZN(n8108) );
  AND2_X1 U9724 ( .A1(n8109), .A2(n8108), .ZN(n9327) );
  NAND2_X1 U9725 ( .A1(n9331), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8110) );
  INV_X1 U9726 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8111) );
  XNOR2_X1 U9727 ( .A(n8125), .B(n8111), .ZN(n9843) );
  NAND2_X1 U9728 ( .A1(n9842), .A2(n9843), .ZN(n9841) );
  OR2_X1 U9729 ( .A1(n8125), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8112) );
  NAND2_X1 U9730 ( .A1(n9841), .A2(n8112), .ZN(n9346) );
  NAND2_X1 U9731 ( .A1(n9351), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8114) );
  NAND2_X1 U9732 ( .A1(n8126), .A2(n9546), .ZN(n8113) );
  AND2_X1 U9733 ( .A1(n8114), .A2(n8113), .ZN(n9345) );
  NOR2_X1 U9734 ( .A1(n9346), .A2(n9345), .ZN(n9344) );
  AND2_X1 U9735 ( .A1(n8126), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8115) );
  INV_X1 U9736 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n8116) );
  XNOR2_X1 U9737 ( .A(n8117), .B(n8116), .ZN(n8131) );
  INV_X1 U9738 ( .A(n8131), .ZN(n8129) );
  NAND2_X1 U9739 ( .A1(n8119), .A2(n8118), .ZN(n8121) );
  NAND2_X1 U9740 ( .A1(n8121), .A2(n8120), .ZN(n9323) );
  OR2_X1 U9741 ( .A1(n9331), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8123) );
  NAND2_X1 U9742 ( .A1(n9331), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8122) );
  NAND2_X1 U9743 ( .A1(n8123), .A2(n8122), .ZN(n9322) );
  NOR2_X1 U9744 ( .A1(n9323), .A2(n9322), .ZN(n9321) );
  INV_X1 U9745 ( .A(n8123), .ZN(n8124) );
  NOR2_X1 U9746 ( .A1(n9321), .A2(n8124), .ZN(n9846) );
  XNOR2_X1 U9747 ( .A(n8125), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9845) );
  NOR2_X1 U9748 ( .A1(n9846), .A2(n9845), .ZN(n9844) );
  NOR2_X1 U9749 ( .A1(n8125), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9338) );
  XNOR2_X1 U9750 ( .A(n8126), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9337) );
  NOR3_X1 U9751 ( .A1(n9844), .A2(n9338), .A3(n9337), .ZN(n9336) );
  AOI21_X1 U9752 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n8126), .A(n9336), .ZN(
        n8127) );
  XNOR2_X1 U9753 ( .A(n8127), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n8130) );
  OAI21_X1 U9754 ( .B1(n8130), .B2(n9849), .A(n9847), .ZN(n8128) );
  AOI21_X1 U9755 ( .B1(n8129), .B2(n9853), .A(n8128), .ZN(n8133) );
  AOI22_X1 U9756 ( .A1(n8131), .A2(n9853), .B1(n9340), .B2(n8130), .ZN(n8132)
         );
  NOR2_X1 U9757 ( .A1(n8134), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9139) );
  INV_X1 U9758 ( .A(n9139), .ZN(n8135) );
  OAI211_X1 U9759 ( .C1(n5008), .C2(n9857), .A(n8136), .B(n8135), .ZN(P1_U3262) );
  INV_X1 U9760 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8188) );
  INV_X1 U9761 ( .A(n9277), .ZN(n8165) );
  INV_X1 U9762 ( .A(n9739), .ZN(n9497) );
  INV_X1 U9763 ( .A(n9278), .ZN(n8200) );
  NAND2_X1 U9764 ( .A1(n9770), .A2(n9282), .ZN(n8141) );
  INV_X1 U9765 ( .A(n9770), .ZN(n9615) );
  INV_X1 U9766 ( .A(n9282), .ZN(n8167) );
  INV_X1 U9767 ( .A(n9281), .ZN(n8168) );
  OR2_X1 U9768 ( .A1(n9761), .A2(n9261), .ZN(n8252) );
  NAND2_X1 U9769 ( .A1(n9761), .A2(n9261), .ZN(n8417) );
  NAND2_X1 U9770 ( .A1(n8252), .A2(n8417), .ZN(n9569) );
  INV_X1 U9771 ( .A(n9261), .ZN(n9280) );
  AOI22_X1 U9772 ( .A1(n9568), .A2(n9569), .B1(n9761), .B2(n9280), .ZN(n9553)
         );
  NAND2_X1 U9773 ( .A1(n9561), .A2(n9279), .ZN(n8144) );
  NAND2_X1 U9774 ( .A1(n9553), .A2(n8144), .ZN(n8146) );
  INV_X1 U9775 ( .A(n9279), .ZN(n8171) );
  NAND2_X1 U9776 ( .A1(n8146), .A2(n8145), .ZN(n9540) );
  INV_X1 U9777 ( .A(n9751), .ZN(n9548) );
  INV_X1 U9778 ( .A(n9522), .ZN(n9137) );
  OAI21_X1 U9779 ( .B1(n9540), .B2(n8147), .A(n5080), .ZN(n9518) );
  NAND2_X1 U9780 ( .A1(n9479), .A2(n9491), .ZN(n8149) );
  INV_X1 U9781 ( .A(n9491), .ZN(n9276) );
  NAND2_X1 U9782 ( .A1(n9462), .A2(n9275), .ZN(n8150) );
  NAND2_X1 U9783 ( .A1(n9445), .A2(n9172), .ZN(n8151) );
  NAND2_X1 U9784 ( .A1(n8186), .A2(n9273), .ZN(n8153) );
  NOR2_X1 U9785 ( .A1(n8186), .A2(n9273), .ZN(n8152) );
  AOI21_X1 U9786 ( .B1(n9421), .B2(n8153), .A(n8152), .ZN(n9407) );
  NAND2_X1 U9787 ( .A1(n9413), .A2(n9173), .ZN(n8154) );
  INV_X2 U9788 ( .A(n9413), .ZN(n9716) );
  NAND2_X1 U9789 ( .A1(n9716), .A2(n9395), .ZN(n8155) );
  NAND2_X1 U9790 ( .A1(n9399), .A2(n9251), .ZN(n8281) );
  NAND2_X1 U9791 ( .A1(n9709), .A2(n9271), .ZN(n8160) );
  INV_X1 U9792 ( .A(n8160), .ZN(n8157) );
  OR2_X1 U9793 ( .A1(n9393), .A2(n8157), .ZN(n8158) );
  NAND2_X1 U9794 ( .A1(n9709), .A2(n9397), .ZN(n8283) );
  AND2_X1 U9795 ( .A1(n9713), .A2(n9251), .ZN(n9377) );
  OR2_X1 U9796 ( .A1(n9382), .A2(n9377), .ZN(n8159) );
  NAND2_X1 U9797 ( .A1(n9093), .A2(n8291), .ZN(n8162) );
  OR2_X1 U9798 ( .A1(n8293), .A2(n9784), .ZN(n8161) );
  NAND2_X1 U9799 ( .A1(n9372), .A2(n8163), .ZN(n8364) );
  NAND2_X1 U9800 ( .A1(n9731), .A2(n9275), .ZN(n8197) );
  NAND2_X1 U9801 ( .A1(n9462), .A2(n8164), .ZN(n8196) );
  NAND2_X1 U9802 ( .A1(n9734), .A2(n9491), .ZN(n8195) );
  NAND2_X1 U9803 ( .A1(n9454), .A2(n8195), .ZN(n9474) );
  NAND2_X1 U9804 ( .A1(n9739), .A2(n8165), .ZN(n8303) );
  NAND2_X1 U9805 ( .A1(n9744), .A2(n9489), .ZN(n8201) );
  NAND2_X1 U9806 ( .A1(n8303), .A2(n8201), .ZN(n8166) );
  NAND2_X1 U9807 ( .A1(n8166), .A2(n8304), .ZN(n8270) );
  OR2_X1 U9808 ( .A1(n9528), .A2(n8200), .ZN(n8263) );
  NAND2_X1 U9809 ( .A1(n9528), .A2(n8200), .ZN(n8423) );
  NAND2_X1 U9810 ( .A1(n9770), .A2(n8167), .ZN(n8233) );
  NAND2_X1 U9811 ( .A1(n9586), .A2(n8233), .ZN(n9606) );
  INV_X1 U9812 ( .A(n9604), .ZN(n8228) );
  OR2_X1 U9813 ( .A1(n9766), .A2(n8168), .ZN(n8248) );
  NAND2_X1 U9814 ( .A1(n9766), .A2(n8168), .ZN(n8232) );
  NAND2_X1 U9815 ( .A1(n8248), .A2(n8232), .ZN(n9590) );
  INV_X1 U9816 ( .A(n9586), .ZN(n8169) );
  NAND2_X1 U9817 ( .A1(n9587), .A2(n8232), .ZN(n9571) );
  INV_X1 U9818 ( .A(n9569), .ZN(n9570) );
  OR2_X1 U9819 ( .A1(n9561), .A2(n8171), .ZN(n8257) );
  NAND2_X1 U9820 ( .A1(n9561), .A2(n8171), .ZN(n8260) );
  NAND2_X1 U9821 ( .A1(n8257), .A2(n8260), .ZN(n9554) );
  OR2_X1 U9822 ( .A1(n9751), .A2(n9137), .ZN(n8262) );
  NAND2_X1 U9823 ( .A1(n9751), .A2(n9137), .ZN(n8261) );
  NAND2_X1 U9824 ( .A1(n8262), .A2(n8261), .ZN(n9541) );
  NAND2_X1 U9825 ( .A1(n8172), .A2(n8261), .ZN(n9519) );
  NAND2_X1 U9826 ( .A1(n9520), .A2(n9519), .ZN(n8173) );
  OR2_X1 U9827 ( .A1(n9744), .A2(n9489), .ZN(n9485) );
  NAND3_X1 U9828 ( .A1(n8304), .A2(n9506), .A3(n9485), .ZN(n8174) );
  NAND2_X1 U9829 ( .A1(n9725), .A2(n9172), .ZN(n8347) );
  NAND2_X1 U9830 ( .A1(n9441), .A2(n8340), .ZN(n9424) );
  INV_X1 U9831 ( .A(n9273), .ZN(n9250) );
  NAND2_X1 U9832 ( .A1(n8186), .A2(n9250), .ZN(n8351) );
  NAND2_X1 U9833 ( .A1(n9424), .A2(n9423), .ZN(n9422) );
  NAND2_X1 U9834 ( .A1(n9422), .A2(n8343), .ZN(n9409) );
  NAND2_X1 U9835 ( .A1(n9716), .A2(n9173), .ZN(n8356) );
  NAND2_X1 U9836 ( .A1(n8345), .A2(n8356), .ZN(n9408) );
  NAND2_X1 U9837 ( .A1(n9381), .A2(n8358), .ZN(n8175) );
  XNOR2_X1 U9838 ( .A(n8175), .B(n4933), .ZN(n8185) );
  NAND2_X1 U9839 ( .A1(n4335), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8180) );
  NAND2_X1 U9840 ( .A1(n8176), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8179) );
  NAND2_X1 U9841 ( .A1(n8177), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8178) );
  NAND2_X1 U9842 ( .A1(n8181), .A2(P1_B_REG_SCAN_IN), .ZN(n8182) );
  NAND2_X1 U9843 ( .A1(n9524), .A2(n8182), .ZN(n9354) );
  NAND2_X1 U9844 ( .A1(n9271), .A2(n9523), .ZN(n8183) );
  OAI21_X1 U9845 ( .B1(n8335), .B2(n9354), .A(n8183), .ZN(n8184) );
  INV_X1 U9846 ( .A(n9372), .ZN(n8187) );
  OR2_X1 U9847 ( .A1(n9766), .A2(n9614), .ZN(n9575) );
  OR2_X2 U9848 ( .A1(n9761), .A2(n9575), .ZN(n9576) );
  NAND2_X1 U9849 ( .A1(n9479), .A2(n9494), .ZN(n9478) );
  NOR2_X2 U9850 ( .A1(n5088), .A2(n9725), .ZN(n9443) );
  AND2_X2 U9851 ( .A1(n9722), .A2(n9443), .ZN(n9428) );
  OAI211_X1 U9852 ( .C1(n8187), .C2(n4357), .A(n9613), .B(n9360), .ZN(n9369)
         );
  NAND2_X1 U9853 ( .A1(n9372), .A2(n9695), .ZN(n8191) );
  NAND2_X1 U9854 ( .A1(n8192), .A2(n8191), .ZN(P1_U3551) );
  NAND2_X1 U9855 ( .A1(n8383), .A2(n8193), .ZN(n8381) );
  NAND2_X1 U9856 ( .A1(n8197), .A2(n9454), .ZN(n8194) );
  NAND2_X1 U9857 ( .A1(n8194), .A2(n8196), .ZN(n8339) );
  NAND2_X1 U9858 ( .A1(n8196), .A2(n8195), .ZN(n8348) );
  NAND2_X1 U9859 ( .A1(n8348), .A2(n8197), .ZN(n8198) );
  NAND3_X1 U9860 ( .A1(n9485), .A2(n4334), .A3(n8263), .ZN(n8269) );
  NAND3_X1 U9861 ( .A1(n9485), .A2(n9750), .A3(n8263), .ZN(n8199) );
  OAI21_X1 U9862 ( .B1(n8200), .B2(n4334), .A(n8199), .ZN(n8202) );
  NAND2_X1 U9863 ( .A1(n8202), .A2(n8201), .ZN(n8268) );
  INV_X1 U9864 ( .A(n8304), .ZN(n8267) );
  INV_X1 U9865 ( .A(n8394), .ZN(n8204) );
  NAND2_X1 U9866 ( .A1(n8205), .A2(n8400), .ZN(n8211) );
  AOI21_X1 U9867 ( .B1(n8209), .B2(n8208), .A(n8211), .ZN(n8206) );
  INV_X1 U9868 ( .A(n8210), .ZN(n8398) );
  NAND2_X1 U9869 ( .A1(n8208), .A2(n8207), .ZN(n8392) );
  NOR2_X1 U9870 ( .A1(n8209), .A2(n8392), .ZN(n8212) );
  INV_X1 U9871 ( .A(n8214), .ZN(n8216) );
  NOR2_X1 U9872 ( .A1(n8216), .A2(n8215), .ZN(n8218) );
  MUX2_X1 U9873 ( .A(n8218), .B(n8217), .S(n8381), .Z(n8223) );
  NAND2_X1 U9874 ( .A1(n8239), .A2(n8219), .ZN(n8221) );
  MUX2_X1 U9875 ( .A(n8221), .B(n8220), .S(n8381), .Z(n8222) );
  INV_X1 U9876 ( .A(n8224), .ZN(n8225) );
  NAND3_X1 U9877 ( .A1(n8226), .A2(n8236), .A3(n8238), .ZN(n8227) );
  NAND3_X1 U9878 ( .A1(n8227), .A2(n8243), .A3(n8244), .ZN(n8229) );
  AOI21_X1 U9879 ( .B1(n8229), .B2(n8237), .A(n8228), .ZN(n8231) );
  INV_X1 U9880 ( .A(n8408), .ZN(n8230) );
  NAND2_X1 U9881 ( .A1(n8417), .A2(n8232), .ZN(n8253) );
  INV_X1 U9882 ( .A(n8233), .ZN(n8234) );
  OR2_X1 U9883 ( .A1(n8253), .A2(n8234), .ZN(n8385) );
  INV_X1 U9884 ( .A(n8235), .ZN(n8240) );
  AND2_X1 U9885 ( .A1(n8237), .A2(n8236), .ZN(n8241) );
  NAND2_X1 U9886 ( .A1(n8241), .A2(n8238), .ZN(n8402) );
  AOI21_X1 U9887 ( .B1(n8240), .B2(n8239), .A(n8402), .ZN(n8247) );
  INV_X1 U9888 ( .A(n8241), .ZN(n8246) );
  AND2_X1 U9889 ( .A1(n8243), .A2(n8242), .ZN(n8245) );
  OAI21_X1 U9890 ( .B1(n8246), .B2(n8245), .A(n8244), .ZN(n8405) );
  OAI21_X1 U9891 ( .B1(n8247), .B2(n8405), .A(n8408), .ZN(n8249) );
  AND2_X1 U9892 ( .A1(n8252), .A2(n8248), .ZN(n8416) );
  NAND2_X1 U9893 ( .A1(n8416), .A2(n9586), .ZN(n8407) );
  AOI21_X1 U9894 ( .B1(n8250), .B2(n8249), .A(n8407), .ZN(n8251) );
  AOI22_X1 U9895 ( .A1(n8253), .A2(n8252), .B1(n4334), .B2(n9599), .ZN(n8255)
         );
  AOI21_X1 U9896 ( .B1(n8417), .B2(n9281), .A(n8381), .ZN(n8254) );
  INV_X1 U9897 ( .A(n9554), .ZN(n8256) );
  AND2_X1 U9898 ( .A1(n8262), .A2(n8257), .ZN(n8412) );
  INV_X1 U9899 ( .A(n8423), .ZN(n8259) );
  INV_X1 U9900 ( .A(n8261), .ZN(n8258) );
  AOI211_X1 U9901 ( .C1(n8264), .C2(n8412), .A(n8259), .B(n8258), .ZN(n8266)
         );
  AND2_X1 U9902 ( .A1(n8261), .A2(n8260), .ZN(n8419) );
  NAND2_X1 U9903 ( .A1(n8263), .A2(n8262), .ZN(n8424) );
  AOI21_X1 U9904 ( .B1(n8264), .B2(n8419), .A(n8424), .ZN(n8265) );
  INV_X1 U9905 ( .A(n8270), .ZN(n8349) );
  NAND2_X1 U9906 ( .A1(n8304), .A2(n9485), .ZN(n8344) );
  MUX2_X1 U9907 ( .A(n8349), .B(n8344), .S(n8381), .Z(n8271) );
  INV_X1 U9908 ( .A(n9474), .ZN(n8329) );
  MUX2_X1 U9909 ( .A(n8340), .B(n8347), .S(n8381), .Z(n8274) );
  INV_X1 U9910 ( .A(n8343), .ZN(n8275) );
  INV_X1 U9911 ( .A(n8351), .ZN(n8276) );
  NAND2_X1 U9912 ( .A1(n8283), .A2(n8281), .ZN(n8354) );
  AOI21_X1 U9913 ( .B1(n8282), .B2(n8346), .A(n8354), .ZN(n8277) );
  INV_X1 U9914 ( .A(n8358), .ZN(n8279) );
  INV_X1 U9915 ( .A(n8346), .ZN(n8278) );
  AOI21_X1 U9916 ( .B1(n8282), .B2(n8281), .A(n8280), .ZN(n8285) );
  INV_X1 U9917 ( .A(n8283), .ZN(n8284) );
  NOR2_X1 U9918 ( .A1(n5081), .A2(n8381), .ZN(n8287) );
  MUX2_X1 U9919 ( .A(n8364), .B(n8359), .S(n8381), .Z(n8286) );
  OAI21_X1 U9920 ( .B1(n8288), .B2(n8287), .A(n8286), .ZN(n8297) );
  NAND2_X1 U9921 ( .A1(n8498), .A2(n8291), .ZN(n8290) );
  OR2_X1 U9922 ( .A1(n8293), .A2(n8499), .ZN(n8289) );
  MUX2_X1 U9923 ( .A(n8381), .B(n8297), .S(n9361), .Z(n8296) );
  NAND2_X1 U9924 ( .A1(n9085), .A2(n8291), .ZN(n8295) );
  OR2_X1 U9925 ( .A1(n8293), .A2(n8292), .ZN(n8294) );
  INV_X1 U9926 ( .A(n8335), .ZN(n9270) );
  NAND3_X1 U9927 ( .A1(n8296), .A2(n9352), .A3(n9270), .ZN(n8302) );
  NAND2_X1 U9928 ( .A1(n9352), .A2(n9355), .ZN(n8380) );
  NAND2_X1 U9929 ( .A1(n8302), .A2(n8301), .ZN(n8379) );
  XNOR2_X1 U9930 ( .A(n9744), .B(n9489), .ZN(n9505) );
  NAND2_X1 U9931 ( .A1(n8305), .A2(n8338), .ZN(n8307) );
  NOR2_X1 U9932 ( .A1(n8307), .A2(n8306), .ZN(n8314) );
  NOR2_X1 U9933 ( .A1(n8308), .A2(n7117), .ZN(n8312) );
  NOR2_X1 U9934 ( .A1(n8310), .A2(n8309), .ZN(n8311) );
  NAND4_X1 U9935 ( .A1(n8314), .A2(n8313), .A3(n8312), .A4(n8311), .ZN(n8315)
         );
  NOR2_X1 U9936 ( .A1(n8316), .A2(n8315), .ZN(n8317) );
  AND2_X1 U9937 ( .A1(n8318), .A2(n8317), .ZN(n8321) );
  NAND4_X1 U9938 ( .A1(n8322), .A2(n8321), .A3(n8320), .A4(n8319), .ZN(n8323)
         );
  OR4_X1 U9939 ( .A1(n9590), .A2(n9606), .A3(n8324), .A4(n8323), .ZN(n8325) );
  NOR2_X1 U9940 ( .A1(n9569), .A2(n8325), .ZN(n8326) );
  NAND4_X1 U9941 ( .A1(n9520), .A2(n8419), .A3(n8412), .A4(n8326), .ZN(n8327)
         );
  NOR2_X1 U9942 ( .A1(n9505), .A2(n8327), .ZN(n8328) );
  AND4_X1 U9943 ( .A1(n9456), .A2(n8329), .A3(n9486), .A4(n8328), .ZN(n8330)
         );
  NAND3_X1 U9944 ( .A1(n9423), .A2(n8331), .A3(n8330), .ZN(n8332) );
  NOR2_X1 U9945 ( .A1(n9408), .A2(n8332), .ZN(n8333) );
  AND4_X1 U9946 ( .A1(n8334), .A2(n9382), .A3(n9393), .A4(n8333), .ZN(n8337)
         );
  OR2_X1 U9947 ( .A1(n9361), .A2(n8335), .ZN(n8431) );
  NAND2_X1 U9948 ( .A1(n9361), .A2(n8335), .ZN(n8365) );
  AND2_X1 U9949 ( .A1(n8431), .A2(n8365), .ZN(n8336) );
  NAND4_X1 U9950 ( .A1(n8337), .A2(n8434), .A3(n8336), .A4(n8380), .ZN(n8369)
         );
  NAND2_X1 U9951 ( .A1(n8340), .A2(n8339), .ZN(n8341) );
  NAND2_X1 U9952 ( .A1(n8341), .A2(n8347), .ZN(n8342) );
  NAND2_X1 U9953 ( .A1(n8343), .A2(n8342), .ZN(n8352) );
  NOR2_X1 U9954 ( .A1(n8352), .A2(n8344), .ZN(n8428) );
  AND2_X1 U9955 ( .A1(n8346), .A2(n8345), .ZN(n8361) );
  INV_X1 U9956 ( .A(n8347), .ZN(n8350) );
  NOR3_X1 U9957 ( .A1(n8350), .A2(n8349), .A3(n8348), .ZN(n8353) );
  OAI21_X1 U9958 ( .B1(n8353), .B2(n8352), .A(n8351), .ZN(n8355) );
  AOI21_X1 U9959 ( .B1(n8361), .B2(n8355), .A(n8354), .ZN(n8357) );
  NAND2_X1 U9960 ( .A1(n8357), .A2(n8356), .ZN(n8426) );
  AOI21_X1 U9961 ( .B1(n8428), .B2(n9506), .A(n8426), .ZN(n8363) );
  INV_X1 U9962 ( .A(n8357), .ZN(n8360) );
  OAI211_X1 U9963 ( .C1(n8361), .C2(n8360), .A(n8359), .B(n8358), .ZN(n8429)
         );
  OAI22_X1 U9964 ( .A1(n8363), .A2(n8429), .B1(n9707), .B2(n8362), .ZN(n8366)
         );
  NAND2_X1 U9965 ( .A1(n8365), .A2(n8364), .ZN(n8432) );
  OAI22_X1 U9966 ( .A1(n8366), .A2(n8432), .B1(n9355), .B2(n8431), .ZN(n8368)
         );
  AOI211_X1 U9967 ( .C1(n8368), .C2(n8434), .A(n8299), .B(n8367), .ZN(n8371)
         );
  INV_X1 U9968 ( .A(n8369), .ZN(n8370) );
  NOR2_X1 U9969 ( .A1(n8371), .A2(n8370), .ZN(n8375) );
  INV_X1 U9970 ( .A(n8434), .ZN(n8384) );
  AOI211_X1 U9971 ( .C1(n8384), .C2(n8383), .A(n8445), .B(n8382), .ZN(n8440)
         );
  INV_X1 U9972 ( .A(n8385), .ZN(n8415) );
  OAI21_X1 U9973 ( .B1(n8388), .B2(n8387), .A(n8386), .ZN(n8396) );
  OAI211_X1 U9974 ( .C1(n8391), .C2(n4511), .A(n8390), .B(n8389), .ZN(n8395)
         );
  INV_X1 U9975 ( .A(n8392), .ZN(n8393) );
  OAI211_X1 U9976 ( .C1(n8396), .C2(n8395), .A(n8394), .B(n8393), .ZN(n8399)
         );
  AOI211_X1 U9977 ( .C1(n8400), .C2(n8399), .A(n8398), .B(n8397), .ZN(n8404)
         );
  INV_X1 U9978 ( .A(n8401), .ZN(n8403) );
  NOR3_X1 U9979 ( .A1(n8404), .A2(n8403), .A3(n8402), .ZN(n8411) );
  INV_X1 U9980 ( .A(n8405), .ZN(n8406) );
  NAND2_X1 U9981 ( .A1(n8406), .A2(n9604), .ZN(n8410) );
  INV_X1 U9982 ( .A(n8407), .ZN(n8409) );
  OAI211_X1 U9983 ( .C1(n8411), .C2(n8410), .A(n8409), .B(n8408), .ZN(n8414)
         );
  INV_X1 U9984 ( .A(n8412), .ZN(n8413) );
  AOI21_X1 U9985 ( .B1(n8415), .B2(n8414), .A(n8413), .ZN(n8422) );
  INV_X1 U9986 ( .A(n8416), .ZN(n8418) );
  NAND2_X1 U9987 ( .A1(n8418), .A2(n8417), .ZN(n8421) );
  INV_X1 U9988 ( .A(n8419), .ZN(n8420) );
  AOI21_X1 U9989 ( .B1(n8422), .B2(n8421), .A(n8420), .ZN(n8425) );
  OAI21_X1 U9990 ( .B1(n8425), .B2(n8424), .A(n8423), .ZN(n8427) );
  AOI21_X1 U9991 ( .B1(n8428), .B2(n8427), .A(n8426), .ZN(n8430) );
  NOR2_X1 U9992 ( .A1(n8430), .A2(n8429), .ZN(n8433) );
  OAI21_X1 U9993 ( .B1(n8433), .B2(n8432), .A(n8431), .ZN(n8435) );
  AOI21_X1 U9994 ( .B1(n8435), .B2(n8434), .A(n8299), .ZN(n8436) );
  MUX2_X1 U9995 ( .A(n8438), .B(n8437), .S(n8436), .Z(n8439) );
  NOR3_X1 U9996 ( .A1(n8444), .A2(n8443), .A3(n8442), .ZN(n8447) );
  OAI21_X1 U9997 ( .B1(n8448), .B2(n8445), .A(P1_B_REG_SCAN_IN), .ZN(n8446) );
  OAI22_X1 U9998 ( .A1(n8449), .A2(n8448), .B1(n8447), .B2(n8446), .ZN(
        P1_U3242) );
  AND3_X1 U9999 ( .A1(n8450), .A2(n8452), .A3(n8451), .ZN(n8453) );
  OAI21_X1 U10000 ( .B1(n8454), .B2(n8453), .A(n9809), .ZN(n8460) );
  NAND2_X1 U10001 ( .A1(n9273), .A2(n9524), .ZN(n8456) );
  NAND2_X1 U10002 ( .A1(n9275), .A2(n9523), .ZN(n8455) );
  NAND2_X1 U10003 ( .A1(n8456), .A2(n8455), .ZN(n9440) );
  OAI22_X1 U10004 ( .A1(n9446), .A2(n9814), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8457), .ZN(n8458) );
  AOI21_X1 U10005 ( .B1(n9440), .B2(n9254), .A(n8458), .ZN(n8459) );
  OAI211_X1 U10006 ( .C1(n9445), .C2(n9800), .A(n8460), .B(n8459), .ZN(
        P1_U3229) );
  XNOR2_X1 U10007 ( .A(n8616), .B(n8491), .ZN(n8464) );
  XNOR2_X1 U10008 ( .A(n8464), .B(n8948), .ZN(n8612) );
  XNOR2_X1 U10009 ( .A(n9080), .B(n8491), .ZN(n8465) );
  XNOR2_X1 U10010 ( .A(n8465), .B(n8938), .ZN(n8544) );
  XNOR2_X1 U10011 ( .A(n9073), .B(n4329), .ZN(n8466) );
  NAND2_X1 U10012 ( .A1(n8466), .A2(n8924), .ZN(n8467) );
  OAI21_X1 U10013 ( .B1(n8466), .B2(n8924), .A(n8467), .ZN(n8554) );
  INV_X1 U10014 ( .A(n8467), .ZN(n8587) );
  XNOR2_X1 U10015 ( .A(n8931), .B(n8491), .ZN(n8468) );
  XNOR2_X1 U10016 ( .A(n8468), .B(n8903), .ZN(n8586) );
  XNOR2_X1 U10017 ( .A(n8520), .B(n8491), .ZN(n8470) );
  XNOR2_X1 U10018 ( .A(n8470), .B(n8622), .ZN(n8521) );
  NAND2_X1 U10019 ( .A1(n8470), .A2(n8622), .ZN(n8471) );
  XOR2_X1 U10020 ( .A(n8491), .B(n9058), .Z(n8568) );
  XNOR2_X1 U10021 ( .A(n8534), .B(n8491), .ZN(n8472) );
  XNOR2_X1 U10022 ( .A(n8472), .B(n8893), .ZN(n8530) );
  INV_X1 U10023 ( .A(n8893), .ZN(n8620) );
  XNOR2_X1 U10024 ( .A(n9047), .B(n8491), .ZN(n8475) );
  XNOR2_X1 U10025 ( .A(n8475), .B(n8877), .ZN(n8578) );
  XNOR2_X1 U10026 ( .A(n8477), .B(n8491), .ZN(n8511) );
  XNOR2_X1 U10027 ( .A(n9036), .B(n8491), .ZN(n8478) );
  XNOR2_X1 U10028 ( .A(n8478), .B(n8516), .ZN(n8561) );
  INV_X1 U10029 ( .A(n8478), .ZN(n8479) );
  XNOR2_X1 U10030 ( .A(n9030), .B(n8491), .ZN(n8480) );
  XNOR2_X1 U10031 ( .A(n8480), .B(n8823), .ZN(n8538) );
  NOR2_X1 U10032 ( .A1(n8480), .A2(n8847), .ZN(n8481) );
  XNOR2_X1 U10033 ( .A(n9024), .B(n4329), .ZN(n8483) );
  XNOR2_X1 U10034 ( .A(n8485), .B(n8483), .ZN(n8597) );
  INV_X1 U10035 ( .A(n8483), .ZN(n8484) );
  OR2_X1 U10036 ( .A1(n8485), .A2(n8484), .ZN(n8486) );
  XNOR2_X1 U10037 ( .A(n8816), .B(n8491), .ZN(n8489) );
  NAND2_X1 U10038 ( .A1(n8489), .A2(n8798), .ZN(n8490) );
  OAI21_X1 U10039 ( .B1(n8489), .B2(n8798), .A(n8490), .ZN(n8501) );
  NOR2_X1 U10040 ( .A1(n8608), .A2(n8803), .ZN(n8495) );
  AOI22_X1 U10041 ( .A1(n8798), .A2(n8606), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8493) );
  OAI21_X1 U10042 ( .B1(n8619), .B2(n8603), .A(n8493), .ZN(n8494) );
  AOI211_X1 U10043 ( .C1(n8965), .C2(n8615), .A(n8495), .B(n8494), .ZN(n8496)
         );
  OAI21_X1 U10044 ( .B1(n8497), .B2(n8610), .A(n8496), .ZN(P2_U3160) );
  INV_X1 U10045 ( .A(n8498), .ZN(n9092) );
  OAI222_X1 U10046 ( .A1(n4336), .A2(n9092), .B1(n8500), .B2(P1_U3086), .C1(
        n8499), .C2(n9789), .ZN(P1_U3325) );
  INV_X1 U10047 ( .A(n8816), .ZN(n8510) );
  NAND2_X1 U10048 ( .A1(n8503), .A2(n8502), .ZN(n8509) );
  INV_X1 U10049 ( .A(n8813), .ZN(n8507) );
  AOI22_X1 U10050 ( .A1(n8833), .A2(n8606), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8504) );
  OAI21_X1 U10051 ( .B1(n8505), .B2(n8603), .A(n8504), .ZN(n8506) );
  AOI21_X1 U10052 ( .B1(n8507), .B2(n8593), .A(n8506), .ZN(n8508) );
  OAI211_X1 U10053 ( .C1(n8510), .C2(n8596), .A(n8509), .B(n8508), .ZN(
        P2_U3154) );
  XNOR2_X1 U10054 ( .A(n8511), .B(n8868), .ZN(n8512) );
  XNOR2_X1 U10055 ( .A(n8513), .B(n8512), .ZN(n8519) );
  AOI22_X1 U10056 ( .A1(n8860), .A2(n8606), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8515) );
  NAND2_X1 U10057 ( .A1(n8863), .A2(n8593), .ZN(n8514) );
  OAI211_X1 U10058 ( .C1(n8516), .C2(n8603), .A(n8515), .B(n8514), .ZN(n8517)
         );
  AOI21_X1 U10059 ( .B1(n9042), .B2(n8615), .A(n8517), .ZN(n8518) );
  OAI21_X1 U10060 ( .B1(n8519), .B2(n8610), .A(n8518), .ZN(P2_U3156) );
  AOI21_X1 U10061 ( .B1(n8522), .B2(n8521), .A(n8610), .ZN(n8524) );
  NAND2_X1 U10062 ( .A1(n8524), .A2(n8523), .ZN(n8528) );
  NAND2_X1 U10063 ( .A1(n8939), .A2(n8606), .ZN(n8525) );
  NAND2_X1 U10064 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8769) );
  OAI211_X1 U10065 ( .C1(n8904), .C2(n8603), .A(n8525), .B(n8769), .ZN(n8526)
         );
  AOI21_X1 U10066 ( .B1(n8908), .B2(n8593), .A(n8526), .ZN(n8527) );
  OAI211_X1 U10067 ( .C1(n9063), .C2(n8596), .A(n8528), .B(n8527), .ZN(
        P2_U3159) );
  XOR2_X1 U10068 ( .A(n8529), .B(n8530), .Z(n8536) );
  AOI22_X1 U10069 ( .A1(n8860), .A2(n8571), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8532) );
  NAND2_X1 U10070 ( .A1(n8593), .A2(n8884), .ZN(n8531) );
  OAI211_X1 U10071 ( .C1(n8904), .C2(n8574), .A(n8532), .B(n8531), .ZN(n8533)
         );
  AOI21_X1 U10072 ( .B1(n8534), .B2(n8615), .A(n8533), .ZN(n8535) );
  OAI21_X1 U10073 ( .B1(n8536), .B2(n8610), .A(n8535), .ZN(P2_U3163) );
  XOR2_X1 U10074 ( .A(n8538), .B(n8537), .Z(n8543) );
  NAND2_X1 U10075 ( .A1(n8859), .A2(n8606), .ZN(n8540) );
  AOI22_X1 U10076 ( .A1(n8833), .A2(n8571), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8539) );
  OAI211_X1 U10077 ( .C1(n8835), .C2(n8608), .A(n8540), .B(n8539), .ZN(n8541)
         );
  AOI21_X1 U10078 ( .B1(n9030), .B2(n8615), .A(n8541), .ZN(n8542) );
  OAI21_X1 U10079 ( .B1(n8543), .B2(n8610), .A(n8542), .ZN(P2_U3165) );
  XNOR2_X1 U10080 ( .A(n8545), .B(n8544), .ZN(n8551) );
  NAND2_X1 U10081 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3151), .ZN(n8696) );
  OAI21_X1 U10082 ( .B1(n8924), .B2(n8603), .A(n8696), .ZN(n8546) );
  AOI21_X1 U10083 ( .B1(n8606), .B2(n8948), .A(n8546), .ZN(n8547) );
  OAI21_X1 U10084 ( .B1(n8548), .B2(n8608), .A(n8547), .ZN(n8549) );
  AOI21_X1 U10085 ( .B1(n9080), .B2(n8615), .A(n8549), .ZN(n8550) );
  OAI21_X1 U10086 ( .B1(n8551), .B2(n8610), .A(n8550), .ZN(P2_U3166) );
  AOI21_X1 U10087 ( .B1(n8554), .B2(n8553), .A(n8552), .ZN(n8559) );
  NAND2_X1 U10088 ( .A1(n8939), .A2(n8571), .ZN(n8555) );
  NAND2_X1 U10089 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8719) );
  OAI211_X1 U10090 ( .C1(n8604), .C2(n8574), .A(n8555), .B(n8719), .ZN(n8556)
         );
  AOI21_X1 U10091 ( .B1(n8942), .B2(n8593), .A(n8556), .ZN(n8558) );
  NAND2_X1 U10092 ( .A1(n9073), .A2(n8615), .ZN(n8557) );
  OAI211_X1 U10093 ( .C1(n8559), .C2(n8610), .A(n8558), .B(n8557), .ZN(
        P2_U3168) );
  XOR2_X1 U10094 ( .A(n8560), .B(n8561), .Z(n8567) );
  INV_X1 U10095 ( .A(n8562), .ZN(n8850) );
  NAND2_X1 U10096 ( .A1(n8848), .A2(n8606), .ZN(n8564) );
  AOI22_X1 U10097 ( .A1(n8847), .A2(n8571), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8563) );
  OAI211_X1 U10098 ( .C1(n8850), .C2(n8608), .A(n8564), .B(n8563), .ZN(n8565)
         );
  AOI21_X1 U10099 ( .B1(n9036), .B2(n8615), .A(n8565), .ZN(n8566) );
  OAI21_X1 U10100 ( .B1(n8567), .B2(n8610), .A(n8566), .ZN(P2_U3169) );
  XNOR2_X1 U10101 ( .A(n8568), .B(n8621), .ZN(n8569) );
  XNOR2_X1 U10102 ( .A(n8570), .B(n8569), .ZN(n8577) );
  AOI22_X1 U10103 ( .A1(n8620), .A2(n8571), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8573) );
  NAND2_X1 U10104 ( .A1(n8593), .A2(n8897), .ZN(n8572) );
  OAI211_X1 U10105 ( .C1(n8925), .C2(n8574), .A(n8573), .B(n8572), .ZN(n8575)
         );
  AOI21_X1 U10106 ( .B1(n9058), .B2(n8615), .A(n8575), .ZN(n8576) );
  OAI21_X1 U10107 ( .B1(n8577), .B2(n8610), .A(n8576), .ZN(P2_U3173) );
  XOR2_X1 U10108 ( .A(n8579), .B(n8578), .Z(n8584) );
  AOI22_X1 U10109 ( .A1(n8620), .A2(n8606), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8581) );
  NAND2_X1 U10110 ( .A1(n8593), .A2(n8869), .ZN(n8580) );
  OAI211_X1 U10111 ( .C1(n8868), .C2(n8603), .A(n8581), .B(n8580), .ZN(n8582)
         );
  AOI21_X1 U10112 ( .B1(n9047), .B2(n8615), .A(n8582), .ZN(n8583) );
  OAI21_X1 U10113 ( .B1(n8584), .B2(n8610), .A(n8583), .ZN(P2_U3175) );
  INV_X1 U10114 ( .A(n8585), .ZN(n8590) );
  NOR3_X1 U10115 ( .A1(n8552), .A2(n8587), .A3(n8586), .ZN(n8589) );
  OAI21_X1 U10116 ( .B1(n8590), .B2(n8589), .A(n8588), .ZN(n8595) );
  NAND2_X1 U10117 ( .A1(n8950), .A2(n8606), .ZN(n8591) );
  NAND2_X1 U10118 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8741) );
  OAI211_X1 U10119 ( .C1(n8925), .C2(n8603), .A(n8591), .B(n8741), .ZN(n8592)
         );
  AOI21_X1 U10120 ( .B1(n8927), .B2(n8593), .A(n8592), .ZN(n8594) );
  OAI211_X1 U10121 ( .C1(n5036), .C2(n8596), .A(n8595), .B(n8594), .ZN(
        P2_U3178) );
  XNOR2_X1 U10122 ( .A(n8597), .B(n8833), .ZN(n8602) );
  NOR2_X1 U10123 ( .A1(n8608), .A2(n8826), .ZN(n8600) );
  AOI22_X1 U10124 ( .A1(n8847), .A2(n8606), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8598) );
  OAI21_X1 U10125 ( .B1(n8824), .B2(n8603), .A(n8598), .ZN(n8599) );
  AOI211_X1 U10126 ( .C1(n9024), .C2(n8615), .A(n8600), .B(n8599), .ZN(n8601)
         );
  OAI21_X1 U10127 ( .B1(n8602), .B2(n8610), .A(n8601), .ZN(P2_U3180) );
  NAND2_X1 U10128 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8668) );
  OAI21_X1 U10129 ( .B1(n8604), .B2(n8603), .A(n8668), .ZN(n8605) );
  AOI21_X1 U10130 ( .B1(n8606), .B2(n8623), .A(n8605), .ZN(n8607) );
  OAI21_X1 U10131 ( .B1(n8609), .B2(n8608), .A(n8607), .ZN(n8614) );
  AOI211_X1 U10132 ( .C1(n8612), .C2(n8611), .A(n8610), .B(n4414), .ZN(n8613)
         );
  AOI211_X1 U10133 ( .C1(n8616), .C2(n8615), .A(n8614), .B(n8613), .ZN(n8617)
         );
  INV_X1 U10134 ( .A(n8617), .ZN(P2_U3181) );
  INV_X2 U10135 ( .A(P2_U3893), .ZN(n8739) );
  MUX2_X1 U10136 ( .A(n8780), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8739), .Z(
        P2_U3522) );
  MUX2_X1 U10137 ( .A(n8618), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8739), .Z(
        P2_U3521) );
  INV_X1 U10138 ( .A(n8619), .ZN(n8797) );
  MUX2_X1 U10139 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8797), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10140 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n5959), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10141 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8798), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10142 ( .A(n8833), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8739), .Z(
        P2_U3517) );
  MUX2_X1 U10143 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8847), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10144 ( .A(n8859), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8739), .Z(
        P2_U3515) );
  MUX2_X1 U10145 ( .A(n8848), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8739), .Z(
        P2_U3514) );
  MUX2_X1 U10146 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8860), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10147 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8620), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10148 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8621), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10149 ( .A(n8622), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8739), .Z(
        P2_U3510) );
  MUX2_X1 U10150 ( .A(n8939), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8739), .Z(
        P2_U3509) );
  MUX2_X1 U10151 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8950), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10152 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8938), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10153 ( .A(n8948), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8739), .Z(
        P2_U3506) );
  MUX2_X1 U10154 ( .A(n8623), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8739), .Z(
        P2_U3505) );
  MUX2_X1 U10155 ( .A(n8624), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8739), .Z(
        P2_U3504) );
  MUX2_X1 U10156 ( .A(n8625), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8739), .Z(
        P2_U3503) );
  MUX2_X1 U10157 ( .A(n8626), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8739), .Z(
        P2_U3502) );
  MUX2_X1 U10158 ( .A(n8627), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8739), .Z(
        P2_U3501) );
  MUX2_X1 U10159 ( .A(n8628), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8739), .Z(
        P2_U3500) );
  MUX2_X1 U10160 ( .A(n8629), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8739), .Z(
        P2_U3499) );
  MUX2_X1 U10161 ( .A(n8630), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8739), .Z(
        P2_U3498) );
  MUX2_X1 U10162 ( .A(n8631), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8739), .Z(
        P2_U3497) );
  MUX2_X1 U10163 ( .A(n8632), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8739), .Z(
        P2_U3496) );
  MUX2_X1 U10164 ( .A(n8633), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8739), .Z(
        P2_U3495) );
  MUX2_X1 U10165 ( .A(n8634), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8739), .Z(
        P2_U3494) );
  MUX2_X1 U10166 ( .A(n8635), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8739), .Z(
        P2_U3493) );
  MUX2_X1 U10167 ( .A(n6913), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8739), .Z(
        P2_U3492) );
  MUX2_X1 U10168 ( .A(n5697), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8739), .Z(
        P2_U3491) );
  NOR2_X1 U10169 ( .A1(n8655), .A2(n8636), .ZN(n8638) );
  NOR2_X1 U10170 ( .A1(n8638), .A2(n8637), .ZN(n8641) );
  NAND2_X1 U10171 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8681), .ZN(n8639) );
  OAI21_X1 U10172 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n8681), .A(n8639), .ZN(
        n8640) );
  NOR2_X1 U10173 ( .A1(n8641), .A2(n8640), .ZN(n8665) );
  AOI21_X1 U10174 ( .B1(n8641), .B2(n8640), .A(n8665), .ZN(n8664) );
  OAI21_X1 U10175 ( .B1(n10017), .B2(n10269), .A(n8642), .ZN(n8652) );
  MUX2_X1 U10176 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8643), .Z(n8644) );
  NOR2_X1 U10177 ( .A1(n8644), .A2(n8681), .ZN(n8674) );
  AOI21_X1 U10178 ( .B1(n8644), .B2(n8681), .A(n8674), .ZN(n8645) );
  INV_X1 U10179 ( .A(n8645), .ZN(n8649) );
  NOR2_X1 U10180 ( .A1(n8648), .A2(n8649), .ZN(n8673) );
  AOI21_X1 U10181 ( .B1(n8649), .B2(n8648), .A(n8673), .ZN(n8650) );
  NOR2_X1 U10182 ( .A1(n8650), .A2(n10013), .ZN(n8651) );
  AOI211_X1 U10183 ( .C1(n10003), .C2(n8653), .A(n8652), .B(n8651), .ZN(n8663)
         );
  NOR2_X1 U10184 ( .A1(n8655), .A2(n8654), .ZN(n8657) );
  NAND2_X1 U10185 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8681), .ZN(n8658) );
  OAI21_X1 U10186 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8681), .A(n8658), .ZN(
        n8659) );
  AOI21_X1 U10187 ( .B1(n8660), .B2(n8659), .A(n8680), .ZN(n8661) );
  OR2_X1 U10188 ( .A1(n8661), .A2(n9980), .ZN(n8662) );
  OAI211_X1 U10189 ( .C1(n8664), .C2(n10005), .A(n8663), .B(n8662), .ZN(
        P2_U3196) );
  AOI21_X1 U10190 ( .B1(n8667), .B2(n8666), .A(n8700), .ZN(n8686) );
  OAI21_X1 U10191 ( .B1(n10017), .B2(n8669), .A(n8668), .ZN(n8679) );
  MUX2_X1 U10192 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8643), .Z(n8671) );
  NOR2_X1 U10193 ( .A1(n8671), .A2(n8670), .ZN(n8694) );
  AOI21_X1 U10194 ( .B1(n8671), .B2(n8670), .A(n8694), .ZN(n8672) );
  INV_X1 U10195 ( .A(n8672), .ZN(n8676) );
  NOR2_X1 U10196 ( .A1(n8674), .A2(n8673), .ZN(n8675) );
  NOR2_X1 U10197 ( .A1(n8675), .A2(n8676), .ZN(n8693) );
  AOI21_X1 U10198 ( .B1(n8676), .B2(n8675), .A(n8693), .ZN(n8677) );
  NOR2_X1 U10199 ( .A1(n8677), .A2(n10013), .ZN(n8678) );
  AOI211_X1 U10200 ( .C1(n10003), .C2(n8699), .A(n8679), .B(n8678), .ZN(n8685)
         );
  AOI21_X1 U10201 ( .B1(n8049), .B2(n8682), .A(n8688), .ZN(n8683) );
  OR2_X1 U10202 ( .A1(n8683), .A2(n9980), .ZN(n8684) );
  OAI211_X1 U10203 ( .C1(n8686), .C2(n10005), .A(n8685), .B(n8684), .ZN(
        P2_U3197) );
  NOR2_X1 U10204 ( .A1(n8699), .A2(n8687), .ZN(n8689) );
  NAND2_X1 U10205 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8721), .ZN(n8690) );
  OAI21_X1 U10206 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8721), .A(n8690), .ZN(
        n8691) );
  AOI21_X1 U10207 ( .B1(n4419), .B2(n8691), .A(n8720), .ZN(n8709) );
  MUX2_X1 U10208 ( .A(n8953), .B(n9005), .S(n8643), .Z(n8692) );
  AND2_X1 U10209 ( .A1(n8692), .A2(n8702), .ZN(n8712) );
  NOR2_X1 U10210 ( .A1(n8692), .A2(n8702), .ZN(n8715) );
  NOR2_X1 U10211 ( .A1(n8712), .A2(n8715), .ZN(n8695) );
  XOR2_X1 U10212 ( .A(n8695), .B(n8714), .Z(n8707) );
  NAND2_X1 U10213 ( .A1(n9962), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8697) );
  OAI211_X1 U10214 ( .C1(n9958), .C2(n8721), .A(n8697), .B(n8696), .ZN(n8706)
         );
  NOR2_X1 U10215 ( .A1(n8699), .A2(n8698), .ZN(n8701) );
  AOI22_X1 U10216 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8702), .B1(n8721), .B2(
        n9005), .ZN(n8703) );
  AOI21_X1 U10217 ( .B1(n4371), .B2(n8703), .A(n8710), .ZN(n8704) );
  NOR2_X1 U10218 ( .A1(n8704), .A2(n10005), .ZN(n8705) );
  AOI211_X1 U10219 ( .C1(n9949), .C2(n8707), .A(n8706), .B(n8705), .ZN(n8708)
         );
  OAI21_X1 U10220 ( .B1(n8709), .B2(n9980), .A(n8708), .ZN(P2_U3198) );
  AOI21_X1 U10221 ( .B1(n8711), .B2(n9002), .A(n8730), .ZN(n8728) );
  INV_X1 U10222 ( .A(n8712), .ZN(n8713) );
  MUX2_X1 U10223 ( .A(n8941), .B(n9002), .S(n8643), .Z(n8735) );
  XOR2_X1 U10224 ( .A(n8744), .B(n8735), .Z(n8716) );
  OAI21_X1 U10225 ( .B1(n8717), .B2(n8716), .A(n8733), .ZN(n8726) );
  NAND2_X1 U10226 ( .A1(n10003), .A2(n8744), .ZN(n8718) );
  OAI211_X1 U10227 ( .C1(n10017), .C2(n10278), .A(n8719), .B(n8718), .ZN(n8725) );
  AOI21_X1 U10228 ( .B1(n8941), .B2(n8722), .A(n8746), .ZN(n8723) );
  NOR2_X1 U10229 ( .A1(n8723), .A2(n9980), .ZN(n8724) );
  AOI211_X1 U10230 ( .C1(n9949), .C2(n8726), .A(n8725), .B(n8724), .ZN(n8727)
         );
  OAI21_X1 U10231 ( .B1(n8728), .B2(n10005), .A(n8727), .ZN(P2_U3199) );
  NAND2_X1 U10232 ( .A1(n8747), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8756) );
  OAI21_X1 U10233 ( .B1(n8747), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8756), .ZN(
        n8731) );
  AOI21_X1 U10234 ( .B1(n8732), .B2(n8731), .A(n8757), .ZN(n8755) );
  MUX2_X1 U10235 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8643), .Z(n8736) );
  INV_X1 U10236 ( .A(n8760), .ZN(n8738) );
  NAND2_X1 U10237 ( .A1(n8737), .A2(n8736), .ZN(n8761) );
  NAND2_X1 U10238 ( .A1(n8738), .A2(n8761), .ZN(n8740) );
  OAI21_X1 U10239 ( .B1(n8740), .B2(n8739), .A(n9958), .ZN(n8753) );
  INV_X1 U10240 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8742) );
  NOR2_X1 U10241 ( .A1(n8744), .A2(n8743), .ZN(n8745) );
  NAND2_X1 U10242 ( .A1(n8747), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8771) );
  OAI21_X1 U10243 ( .B1(n8747), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8771), .ZN(
        n8748) );
  AOI21_X1 U10244 ( .B1(n8749), .B2(n8748), .A(n8773), .ZN(n8750) );
  NOR2_X1 U10245 ( .A1(n8750), .A2(n9980), .ZN(n8751) );
  AOI211_X1 U10246 ( .C1(n8762), .C2(n8753), .A(n8752), .B(n8751), .ZN(n8754)
         );
  OAI21_X1 U10247 ( .B1(n8755), .B2(n10005), .A(n8754), .ZN(P2_U3200) );
  XNOR2_X1 U10248 ( .A(n8763), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8764) );
  INV_X1 U10249 ( .A(n8764), .ZN(n8758) );
  XNOR2_X1 U10250 ( .A(n8759), .B(n8758), .ZN(n8778) );
  AOI21_X1 U10251 ( .B1(n8762), .B2(n8761), .A(n8760), .ZN(n8766) );
  MUX2_X1 U10252 ( .A(n8911), .B(P2_REG2_REG_19__SCAN_IN), .S(n8763), .Z(n8775) );
  MUX2_X1 U10253 ( .A(n8775), .B(n8764), .S(n8643), .Z(n8765) );
  XNOR2_X1 U10254 ( .A(n8766), .B(n8765), .ZN(n8777) );
  NAND2_X1 U10255 ( .A1(n10003), .A2(n8767), .ZN(n8768) );
  OAI211_X1 U10256 ( .C1(n10017), .C2(n8770), .A(n8769), .B(n8768), .ZN(n8776)
         );
  INV_X1 U10257 ( .A(n8771), .ZN(n8772) );
  NOR2_X1 U10258 ( .A1(n8773), .A2(n8772), .ZN(n8774) );
  NAND2_X1 U10259 ( .A1(n9010), .A2(n8956), .ZN(n8782) );
  NOR2_X1 U10260 ( .A1(n10021), .A2(n8781), .ZN(n8791) );
  OAI21_X1 U10261 ( .B1(n9011), .B2(n8791), .A(n8926), .ZN(n8785) );
  OAI211_X1 U10262 ( .C1(n8926), .C2(n8783), .A(n8782), .B(n8785), .ZN(
        P2_U3202) );
  NAND2_X1 U10263 ( .A1(n8784), .A2(n8956), .ZN(n8786) );
  OAI211_X1 U10264 ( .C1(n8926), .C2(n8787), .A(n8786), .B(n8785), .ZN(
        P2_U3203) );
  NAND2_X1 U10265 ( .A1(n8788), .A2(n8926), .ZN(n8793) );
  NOR2_X1 U10266 ( .A1(n8789), .A2(n8912), .ZN(n8790) );
  AOI211_X1 U10267 ( .C1(n10034), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8791), .B(
        n8790), .ZN(n8792) );
  OAI211_X1 U10268 ( .C1(n8795), .C2(n8794), .A(n8793), .B(n8792), .ZN(
        P2_U3204) );
  XNOR2_X1 U10269 ( .A(n8796), .B(n8808), .ZN(n8802) );
  NAND2_X1 U10270 ( .A1(n8797), .A2(n8949), .ZN(n8800) );
  NAND2_X1 U10271 ( .A1(n8798), .A2(n5656), .ZN(n8799) );
  OAI22_X1 U10272 ( .A1(n8926), .A2(n8804), .B1(n8803), .B2(n10021), .ZN(n8810) );
  INV_X1 U10273 ( .A(n8805), .ZN(n8806) );
  AOI21_X1 U10274 ( .B1(n8808), .B2(n8807), .A(n8806), .ZN(n8964) );
  NOR2_X1 U10275 ( .A1(n8964), .A2(n8959), .ZN(n8809) );
  AOI211_X1 U10276 ( .C1(n8956), .C2(n8965), .A(n8810), .B(n8809), .ZN(n8811)
         );
  OAI21_X1 U10277 ( .B1(n8968), .B2(n10034), .A(n8811), .ZN(P2_U3205) );
  NAND2_X1 U10278 ( .A1(n8812), .A2(n8926), .ZN(n8818) );
  OAI22_X1 U10279 ( .A1(n8926), .A2(n8814), .B1(n8813), .B2(n10021), .ZN(n8815) );
  AOI21_X1 U10280 ( .B1(n8816), .B2(n8956), .A(n8815), .ZN(n8817) );
  OAI211_X1 U10281 ( .C1(n9021), .C2(n8959), .A(n8818), .B(n8817), .ZN(
        P2_U3206) );
  XNOR2_X1 U10282 ( .A(n8819), .B(n8821), .ZN(n9027) );
  XOR2_X1 U10283 ( .A(n8821), .B(n8820), .Z(n8822) );
  OAI222_X1 U10284 ( .A1(n10030), .A2(n8824), .B1(n10028), .B2(n8823), .C1(
        n10026), .C2(n8822), .ZN(n8969) );
  INV_X1 U10285 ( .A(n8969), .ZN(n9022) );
  MUX2_X1 U10286 ( .A(n8825), .B(n9022), .S(n8926), .Z(n8829) );
  INV_X1 U10287 ( .A(n8826), .ZN(n8827) );
  AOI22_X1 U10288 ( .A1(n9024), .A2(n8956), .B1(n8955), .B2(n8827), .ZN(n8828)
         );
  OAI211_X1 U10289 ( .C1(n9027), .C2(n8959), .A(n8829), .B(n8828), .ZN(
        P2_U3207) );
  XNOR2_X1 U10290 ( .A(n8830), .B(n8831), .ZN(n9033) );
  XNOR2_X1 U10291 ( .A(n8832), .B(n8831), .ZN(n8834) );
  AOI222_X1 U10292 ( .A1(n8952), .A2(n8834), .B1(n8833), .B2(n8949), .C1(n8859), .C2(n5656), .ZN(n9028) );
  INV_X1 U10293 ( .A(n9028), .ZN(n8838) );
  INV_X1 U10294 ( .A(n9030), .ZN(n8836) );
  OAI22_X1 U10295 ( .A1(n8836), .A2(n10023), .B1(n8835), .B2(n10021), .ZN(
        n8837) );
  OAI21_X1 U10296 ( .B1(n8838), .B2(n8837), .A(n8926), .ZN(n8840) );
  NAND2_X1 U10297 ( .A1(n10034), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8839) );
  OAI211_X1 U10298 ( .C1(n9033), .C2(n8959), .A(n8840), .B(n8839), .ZN(
        P2_U3208) );
  NAND2_X1 U10299 ( .A1(n8842), .A2(n8841), .ZN(n8844) );
  XNOR2_X1 U10300 ( .A(n8844), .B(n8843), .ZN(n9039) );
  XNOR2_X1 U10301 ( .A(n8846), .B(n8845), .ZN(n8849) );
  AOI222_X1 U10302 ( .A1(n8952), .A2(n8849), .B1(n8848), .B2(n5656), .C1(n8847), .C2(n8949), .ZN(n9034) );
  INV_X1 U10303 ( .A(n9034), .ZN(n8853) );
  OAI22_X1 U10304 ( .A1(n8851), .A2(n10023), .B1(n8850), .B2(n10021), .ZN(
        n8852) );
  OAI21_X1 U10305 ( .B1(n8853), .B2(n8852), .A(n8926), .ZN(n8855) );
  NAND2_X1 U10306 ( .A1(n10034), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8854) );
  OAI211_X1 U10307 ( .C1(n9039), .C2(n8959), .A(n8855), .B(n8854), .ZN(
        P2_U3209) );
  XOR2_X1 U10308 ( .A(n8857), .B(n8856), .Z(n9045) );
  INV_X1 U10309 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8862) );
  XNOR2_X1 U10310 ( .A(n8858), .B(n8857), .ZN(n8861) );
  AOI222_X1 U10311 ( .A1(n8952), .A2(n8861), .B1(n8860), .B2(n5656), .C1(n8859), .C2(n8949), .ZN(n9040) );
  MUX2_X1 U10312 ( .A(n8862), .B(n9040), .S(n8926), .Z(n8865) );
  AOI22_X1 U10313 ( .A1(n9042), .A2(n8956), .B1(n8955), .B2(n8863), .ZN(n8864)
         );
  OAI211_X1 U10314 ( .C1(n9045), .C2(n8959), .A(n8865), .B(n8864), .ZN(
        P2_U3210) );
  XOR2_X1 U10315 ( .A(n8870), .B(n8866), .Z(n8867) );
  OAI222_X1 U10316 ( .A1(n10030), .A2(n8868), .B1(n10028), .B2(n8893), .C1(
        n10026), .C2(n8867), .ZN(n8982) );
  AOI21_X1 U10317 ( .B1(n8955), .B2(n8869), .A(n8982), .ZN(n8875) );
  AOI22_X1 U10318 ( .A1(n9047), .A2(n8956), .B1(P2_REG2_REG_22__SCAN_IN), .B2(
        n10034), .ZN(n8874) );
  INV_X1 U10319 ( .A(n8870), .ZN(n8871) );
  XNOR2_X1 U10320 ( .A(n8872), .B(n8871), .ZN(n9049) );
  NAND2_X1 U10321 ( .A1(n9049), .A2(n8914), .ZN(n8873) );
  OAI211_X1 U10322 ( .C1(n8875), .C2(n10034), .A(n8874), .B(n8873), .ZN(
        P2_U3211) );
  XNOR2_X1 U10323 ( .A(n8876), .B(n8882), .ZN(n8879) );
  OAI22_X1 U10324 ( .A1(n8877), .A2(n10030), .B1(n8904), .B2(n10028), .ZN(
        n8878) );
  AOI21_X1 U10325 ( .B1(n8879), .B2(n8952), .A(n8878), .ZN(n8989) );
  NAND2_X1 U10326 ( .A1(n8881), .A2(n8880), .ZN(n8883) );
  XNOR2_X1 U10327 ( .A(n8883), .B(n5072), .ZN(n8987) );
  AOI22_X1 U10328 ( .A1(n8955), .A2(n8884), .B1(n10034), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n8885) );
  OAI21_X1 U10329 ( .B1(n9055), .B2(n8912), .A(n8885), .ZN(n8886) );
  AOI21_X1 U10330 ( .B1(n8987), .B2(n8914), .A(n8886), .ZN(n8887) );
  OAI21_X1 U10331 ( .B1(n8989), .B2(n10034), .A(n8887), .ZN(P2_U3212) );
  XOR2_X1 U10332 ( .A(n8889), .B(n8888), .Z(n9061) );
  NAND2_X1 U10333 ( .A1(n8890), .A2(n8889), .ZN(n8891) );
  NAND2_X1 U10334 ( .A1(n8892), .A2(n8891), .ZN(n8895) );
  OAI22_X1 U10335 ( .A1(n8893), .A2(n10030), .B1(n8925), .B2(n10028), .ZN(
        n8894) );
  AOI21_X1 U10336 ( .B1(n8895), .B2(n8952), .A(n8894), .ZN(n9057) );
  INV_X1 U10337 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8896) );
  MUX2_X1 U10338 ( .A(n9057), .B(n8896), .S(n10034), .Z(n8899) );
  AOI22_X1 U10339 ( .A1(n9058), .A2(n8956), .B1(n8955), .B2(n8897), .ZN(n8898)
         );
  OAI211_X1 U10340 ( .C1(n9061), .C2(n8959), .A(n8899), .B(n8898), .ZN(
        P2_U3213) );
  NAND2_X1 U10341 ( .A1(n8900), .A2(n8909), .ZN(n8901) );
  NAND3_X1 U10342 ( .A1(n8902), .A2(n8952), .A3(n8901), .ZN(n8907) );
  OAI22_X1 U10343 ( .A1(n8904), .A2(n10030), .B1(n8903), .B2(n10028), .ZN(
        n8905) );
  INV_X1 U10344 ( .A(n8905), .ZN(n8906) );
  NAND2_X1 U10345 ( .A1(n8907), .A2(n8906), .ZN(n9062) );
  AOI21_X1 U10346 ( .B1(n8955), .B2(n8908), .A(n9062), .ZN(n8917) );
  XNOR2_X1 U10347 ( .A(n8910), .B(n8909), .ZN(n9064) );
  INV_X1 U10348 ( .A(n9064), .ZN(n8915) );
  OAI22_X1 U10349 ( .A1(n9063), .A2(n8912), .B1(n8911), .B2(n8926), .ZN(n8913)
         );
  AOI21_X1 U10350 ( .B1(n8915), .B2(n8914), .A(n8913), .ZN(n8916) );
  OAI21_X1 U10351 ( .B1(n8917), .B2(n10034), .A(n8916), .ZN(P2_U3214) );
  NAND2_X1 U10352 ( .A1(n8918), .A2(n8921), .ZN(n8919) );
  INV_X1 U10353 ( .A(n8998), .ZN(n8934) );
  XNOR2_X1 U10354 ( .A(n8922), .B(n8921), .ZN(n8923) );
  OAI222_X1 U10355 ( .A1(n10030), .A2(n8925), .B1(n10028), .B2(n8924), .C1(
        n8923), .C2(n10026), .ZN(n8997) );
  NAND2_X1 U10356 ( .A1(n8997), .A2(n8926), .ZN(n8933) );
  INV_X1 U10357 ( .A(n8927), .ZN(n8928) );
  OAI22_X1 U10358 ( .A1(n8926), .A2(n8929), .B1(n8928), .B2(n10021), .ZN(n8930) );
  AOI21_X1 U10359 ( .B1(n8931), .B2(n8956), .A(n8930), .ZN(n8932) );
  OAI211_X1 U10360 ( .C1(n8934), .C2(n8959), .A(n8933), .B(n8932), .ZN(
        P2_U3215) );
  XNOR2_X1 U10361 ( .A(n8935), .B(n8936), .ZN(n9076) );
  XNOR2_X1 U10362 ( .A(n8937), .B(n8936), .ZN(n8940) );
  AOI222_X1 U10363 ( .A1(n8952), .A2(n8940), .B1(n8939), .B2(n8949), .C1(n8938), .C2(n5656), .ZN(n9071) );
  MUX2_X1 U10364 ( .A(n8941), .B(n9071), .S(n8926), .Z(n8944) );
  AOI22_X1 U10365 ( .A1(n9073), .A2(n8956), .B1(n8955), .B2(n8942), .ZN(n8943)
         );
  OAI211_X1 U10366 ( .C1(n9076), .C2(n8959), .A(n8944), .B(n8943), .ZN(
        P2_U3216) );
  XOR2_X1 U10367 ( .A(n8945), .B(n8946), .Z(n9084) );
  XOR2_X1 U10368 ( .A(n8947), .B(n8946), .Z(n8951) );
  AOI222_X1 U10369 ( .A1(n8952), .A2(n8951), .B1(n8950), .B2(n8949), .C1(n8948), .C2(n5656), .ZN(n9077) );
  MUX2_X1 U10370 ( .A(n8953), .B(n9077), .S(n8926), .Z(n8958) );
  AOI22_X1 U10371 ( .A1(n9080), .A2(n8956), .B1(n8955), .B2(n8954), .ZN(n8957)
         );
  OAI211_X1 U10372 ( .C1(n9084), .C2(n8959), .A(n8958), .B(n8957), .ZN(
        P2_U3217) );
  NAND2_X1 U10373 ( .A1(n9011), .A2(n10096), .ZN(n8962) );
  NAND2_X1 U10374 ( .A1(n10094), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8960) );
  OAI211_X1 U10375 ( .C1(n8961), .C2(n9001), .A(n8962), .B(n8960), .ZN(
        P2_U3490) );
  NAND2_X1 U10376 ( .A1(n10094), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8963) );
  OAI211_X1 U10377 ( .C1(n9016), .C2(n9001), .A(n8963), .B(n8962), .ZN(
        P2_U3489) );
  NAND2_X1 U10378 ( .A1(n8965), .A2(n10080), .ZN(n8966) );
  NAND2_X1 U10379 ( .A1(n8968), .A2(n8967), .ZN(n9017) );
  MUX2_X1 U10380 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9017), .S(n10096), .Z(
        P2_U3487) );
  MUX2_X1 U10381 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8969), .S(n10096), .Z(
        n8972) );
  OAI22_X1 U10382 ( .A1(n9027), .A2(n9009), .B1(n8970), .B2(n9001), .ZN(n8971)
         );
  OR2_X1 U10383 ( .A1(n8972), .A2(n8971), .ZN(P2_U3485) );
  INV_X1 U10384 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8973) );
  MUX2_X1 U10385 ( .A(n8973), .B(n9028), .S(n10096), .Z(n8975) );
  NAND2_X1 U10386 ( .A1(n9030), .A2(n9006), .ZN(n8974) );
  OAI211_X1 U10387 ( .C1(n9033), .C2(n9009), .A(n8975), .B(n8974), .ZN(
        P2_U3484) );
  MUX2_X1 U10388 ( .A(n8976), .B(n9034), .S(n10096), .Z(n8978) );
  NAND2_X1 U10389 ( .A1(n9036), .A2(n9006), .ZN(n8977) );
  OAI211_X1 U10390 ( .C1(n9009), .C2(n9039), .A(n8978), .B(n8977), .ZN(
        P2_U3483) );
  MUX2_X1 U10391 ( .A(n8979), .B(n9040), .S(n10096), .Z(n8981) );
  NAND2_X1 U10392 ( .A1(n9042), .A2(n9006), .ZN(n8980) );
  OAI211_X1 U10393 ( .C1(n9045), .C2(n9009), .A(n8981), .B(n8980), .ZN(
        P2_U3482) );
  INV_X1 U10394 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8983) );
  INV_X1 U10395 ( .A(n8982), .ZN(n9046) );
  MUX2_X1 U10396 ( .A(n8983), .B(n9046), .S(n10096), .Z(n8986) );
  AOI22_X1 U10397 ( .A1(n9049), .A2(n8984), .B1(n9006), .B2(n9047), .ZN(n8985)
         );
  NAND2_X1 U10398 ( .A1(n8986), .A2(n8985), .ZN(P2_U3481) );
  INV_X1 U10399 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8990) );
  NAND2_X1 U10400 ( .A1(n8987), .A2(n10075), .ZN(n8988) );
  AND2_X1 U10401 ( .A1(n8989), .A2(n8988), .ZN(n9053) );
  MUX2_X1 U10402 ( .A(n8990), .B(n9053), .S(n10096), .Z(n8991) );
  OAI21_X1 U10403 ( .B1(n9055), .B2(n9001), .A(n8991), .ZN(P2_U3480) );
  INV_X1 U10404 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8992) );
  MUX2_X1 U10405 ( .A(n8992), .B(n9057), .S(n10096), .Z(n8994) );
  NAND2_X1 U10406 ( .A1(n9058), .A2(n9006), .ZN(n8993) );
  OAI211_X1 U10407 ( .C1(n9009), .C2(n9061), .A(n8994), .B(n8993), .ZN(
        P2_U3479) );
  MUX2_X1 U10408 ( .A(n9062), .B(P2_REG1_REG_19__SCAN_IN), .S(n10094), .Z(
        n8996) );
  OAI22_X1 U10409 ( .A1(n9064), .A2(n9009), .B1(n9063), .B2(n9001), .ZN(n8995)
         );
  OR2_X1 U10410 ( .A1(n8996), .A2(n8995), .ZN(P2_U3478) );
  INV_X1 U10411 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8999) );
  AOI21_X1 U10412 ( .B1(n8998), .B2(n10075), .A(n8997), .ZN(n9067) );
  MUX2_X1 U10413 ( .A(n8999), .B(n9067), .S(n10096), .Z(n9000) );
  OAI21_X1 U10414 ( .B1(n5036), .B2(n9001), .A(n9000), .ZN(P2_U3477) );
  MUX2_X1 U10415 ( .A(n9002), .B(n9071), .S(n10096), .Z(n9004) );
  NAND2_X1 U10416 ( .A1(n9073), .A2(n9006), .ZN(n9003) );
  OAI211_X1 U10417 ( .C1(n9076), .C2(n9009), .A(n9004), .B(n9003), .ZN(
        P2_U3476) );
  MUX2_X1 U10418 ( .A(n9005), .B(n9077), .S(n10096), .Z(n9008) );
  NAND2_X1 U10419 ( .A1(n9080), .A2(n9006), .ZN(n9007) );
  OAI211_X1 U10420 ( .C1(n9084), .C2(n9009), .A(n9008), .B(n9007), .ZN(
        P2_U3475) );
  NAND2_X1 U10421 ( .A1(n9010), .A2(n9079), .ZN(n9012) );
  NAND2_X1 U10422 ( .A1(n10081), .A2(n9011), .ZN(n9014) );
  OAI211_X1 U10423 ( .C1(n10081), .C2(n9013), .A(n9012), .B(n9014), .ZN(
        P2_U3458) );
  NAND2_X1 U10424 ( .A1(n10082), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9015) );
  OAI211_X1 U10425 ( .C1(n9016), .C2(n9070), .A(n9015), .B(n9014), .ZN(
        P2_U3457) );
  MUX2_X1 U10426 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9017), .S(n10081), .Z(
        P2_U3455) );
  MUX2_X1 U10427 ( .A(n9019), .B(n9018), .S(n10081), .Z(n9020) );
  OAI21_X1 U10428 ( .B1(n9021), .B2(n9083), .A(n9020), .ZN(P2_U3454) );
  MUX2_X1 U10429 ( .A(n9023), .B(n9022), .S(n10081), .Z(n9026) );
  NAND2_X1 U10430 ( .A1(n9024), .A2(n9079), .ZN(n9025) );
  OAI211_X1 U10431 ( .C1(n9027), .C2(n9083), .A(n9026), .B(n9025), .ZN(
        P2_U3453) );
  MUX2_X1 U10432 ( .A(n9029), .B(n9028), .S(n10081), .Z(n9032) );
  NAND2_X1 U10433 ( .A1(n9030), .A2(n9079), .ZN(n9031) );
  OAI211_X1 U10434 ( .C1(n9033), .C2(n9083), .A(n9032), .B(n9031), .ZN(
        P2_U3452) );
  INV_X1 U10435 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9035) );
  MUX2_X1 U10436 ( .A(n9035), .B(n9034), .S(n10081), .Z(n9038) );
  NAND2_X1 U10437 ( .A1(n9036), .A2(n9079), .ZN(n9037) );
  OAI211_X1 U10438 ( .C1(n9039), .C2(n9083), .A(n9038), .B(n9037), .ZN(
        P2_U3451) );
  INV_X1 U10439 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9041) );
  MUX2_X1 U10440 ( .A(n9041), .B(n9040), .S(n10081), .Z(n9044) );
  NAND2_X1 U10441 ( .A1(n9042), .A2(n9079), .ZN(n9043) );
  OAI211_X1 U10442 ( .C1(n9045), .C2(n9083), .A(n9044), .B(n9043), .ZN(
        P2_U3450) );
  MUX2_X1 U10443 ( .A(n10158), .B(n9046), .S(n10081), .Z(n9051) );
  AOI22_X1 U10444 ( .A1(n9049), .A2(n9048), .B1(n9079), .B2(n9047), .ZN(n9050)
         );
  NAND2_X1 U10445 ( .A1(n9051), .A2(n9050), .ZN(P2_U3449) );
  INV_X1 U10446 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9052) );
  MUX2_X1 U10447 ( .A(n9053), .B(n9052), .S(n10082), .Z(n9054) );
  OAI21_X1 U10448 ( .B1(n9055), .B2(n9070), .A(n9054), .ZN(P2_U3448) );
  INV_X1 U10449 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9056) );
  MUX2_X1 U10450 ( .A(n9057), .B(n9056), .S(n10082), .Z(n9060) );
  NAND2_X1 U10451 ( .A1(n9058), .A2(n9079), .ZN(n9059) );
  OAI211_X1 U10452 ( .C1(n9061), .C2(n9083), .A(n9060), .B(n9059), .ZN(
        P2_U3447) );
  MUX2_X1 U10453 ( .A(n9062), .B(P2_REG0_REG_19__SCAN_IN), .S(n10082), .Z(
        n9066) );
  OAI22_X1 U10454 ( .A1(n9064), .A2(n9083), .B1(n9063), .B2(n9070), .ZN(n9065)
         );
  OR2_X1 U10455 ( .A1(n9066), .A2(n9065), .ZN(P2_U3446) );
  MUX2_X1 U10456 ( .A(n9068), .B(n9067), .S(n10081), .Z(n9069) );
  OAI21_X1 U10457 ( .B1(n5036), .B2(n9070), .A(n9069), .ZN(P2_U3444) );
  MUX2_X1 U10458 ( .A(n9072), .B(n9071), .S(n10081), .Z(n9075) );
  NAND2_X1 U10459 ( .A1(n9073), .A2(n9079), .ZN(n9074) );
  OAI211_X1 U10460 ( .C1(n9076), .C2(n9083), .A(n9075), .B(n9074), .ZN(
        P2_U3441) );
  INV_X1 U10461 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9078) );
  MUX2_X1 U10462 ( .A(n9078), .B(n9077), .S(n10081), .Z(n9082) );
  NAND2_X1 U10463 ( .A1(n9080), .A2(n9079), .ZN(n9081) );
  OAI211_X1 U10464 ( .C1(n9084), .C2(n9083), .A(n9082), .B(n9081), .ZN(
        P2_U3438) );
  INV_X1 U10465 ( .A(n9085), .ZN(n9783) );
  NOR4_X1 U10466 ( .A1(n9087), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n9086), .ZN(n9088) );
  AOI21_X1 U10467 ( .B1(n9100), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9088), .ZN(
        n9089) );
  OAI21_X1 U10468 ( .B1(n9783), .B2(n9103), .A(n9089), .ZN(P2_U3264) );
  AOI22_X1 U10469 ( .A1(n4607), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9100), .ZN(n9091) );
  OAI21_X1 U10470 ( .B1(n9092), .B2(n9103), .A(n9091), .ZN(P2_U3265) );
  INV_X1 U10471 ( .A(n9093), .ZN(n9786) );
  AOI22_X1 U10472 ( .A1(n9094), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9100), .ZN(n9095) );
  OAI21_X1 U10473 ( .B1(n9786), .B2(n9103), .A(n9095), .ZN(P2_U3266) );
  INV_X1 U10474 ( .A(n9096), .ZN(n9788) );
  AOI21_X1 U10475 ( .B1(n9100), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n9097), .ZN(
        n9098) );
  OAI21_X1 U10476 ( .B1(n9788), .B2(n9103), .A(n9098), .ZN(P2_U3267) );
  INV_X1 U10477 ( .A(n9099), .ZN(n9791) );
  NAND2_X1 U10478 ( .A1(n9100), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9101) );
  OAI211_X1 U10479 ( .C1(n9791), .C2(n9103), .A(n9102), .B(n9101), .ZN(
        P2_U3268) );
  AOI21_X1 U10480 ( .B1(n9106), .B2(n9105), .A(n4409), .ZN(n9113) );
  NAND2_X1 U10481 ( .A1(n9281), .A2(n9524), .ZN(n9108) );
  NAND2_X1 U10482 ( .A1(n9283), .A2(n9523), .ZN(n9107) );
  AND2_X1 U10483 ( .A1(n9108), .A2(n9107), .ZN(n9611) );
  NAND2_X1 U10484 ( .A1(n9267), .A2(n9616), .ZN(n9110) );
  OAI211_X1 U10485 ( .C1(n9611), .C2(n9265), .A(n9110), .B(n9109), .ZN(n9111)
         );
  AOI21_X1 U10486 ( .B1(n9770), .B2(n6649), .A(n9111), .ZN(n9112) );
  OAI21_X1 U10487 ( .B1(n9113), .B2(n9245), .A(n9112), .ZN(P1_U3215) );
  OAI21_X1 U10488 ( .B1(n9114), .B2(n9231), .A(n8450), .ZN(n9118) );
  NAND2_X1 U10489 ( .A1(n9462), .A2(n6649), .ZN(n9116) );
  OAI22_X1 U10490 ( .A1(n9172), .A2(n9490), .B1(n9491), .B2(n9488), .ZN(n9458)
         );
  AOI22_X1 U10491 ( .A1(n9458), .A2(n9254), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9115) );
  OAI211_X1 U10492 ( .C1(n9814), .C2(n9463), .A(n9116), .B(n9115), .ZN(n9117)
         );
  AOI21_X1 U10493 ( .B1(n9118), .B2(n9809), .A(n9117), .ZN(n9119) );
  INV_X1 U10494 ( .A(n9119), .ZN(P1_U3216) );
  XNOR2_X1 U10495 ( .A(n9120), .B(n9794), .ZN(n9123) );
  INV_X1 U10496 ( .A(n9121), .ZN(n9122) );
  NOR2_X1 U10497 ( .A1(n9123), .A2(n9122), .ZN(n9793) );
  AOI21_X1 U10498 ( .B1(n9123), .B2(n9122), .A(n9793), .ZN(n9130) );
  AOI22_X1 U10499 ( .A1(n9254), .A2(n9124), .B1(P1_REG3_REG_10__SCAN_IN), .B2(
        P1_U3086), .ZN(n9125) );
  OAI21_X1 U10500 ( .B1(n9814), .B2(n9126), .A(n9125), .ZN(n9127) );
  AOI21_X1 U10501 ( .B1(n9128), .B2(n6649), .A(n9127), .ZN(n9129) );
  OAI21_X1 U10502 ( .B1(n9130), .B2(n9245), .A(n9129), .ZN(P1_U3217) );
  XNOR2_X1 U10503 ( .A(n9131), .B(n9132), .ZN(n9240) );
  NOR2_X1 U10504 ( .A1(n9240), .A2(n9239), .ZN(n9238) );
  AOI21_X1 U10505 ( .B1(n9132), .B2(n9131), .A(n9238), .ZN(n9136) );
  XNOR2_X1 U10506 ( .A(n9134), .B(n9133), .ZN(n9135) );
  XNOR2_X1 U10507 ( .A(n9136), .B(n9135), .ZN(n9143) );
  NOR2_X1 U10508 ( .A1(n9803), .A2(n9137), .ZN(n9138) );
  AOI211_X1 U10509 ( .C1(n9802), .C2(n9525), .A(n9139), .B(n9138), .ZN(n9140)
         );
  OAI21_X1 U10510 ( .B1(n9814), .B2(n9529), .A(n9140), .ZN(n9141) );
  AOI21_X1 U10511 ( .B1(n9528), .B2(n6649), .A(n9141), .ZN(n9142) );
  OAI21_X1 U10512 ( .B1(n9143), .B2(n9245), .A(n9142), .ZN(P1_U3219) );
  OAI21_X1 U10513 ( .B1(n9146), .B2(n9145), .A(n9144), .ZN(n9147) );
  NAND2_X1 U10514 ( .A1(n9147), .A2(n9809), .ZN(n9152) );
  AOI22_X1 U10515 ( .A1(n9148), .A2(n6901), .B1(n9802), .B2(n9293), .ZN(n9151)
         );
  AOI22_X1 U10516 ( .A1(n6649), .A2(n4511), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n9149), .ZN(n9150) );
  NAND3_X1 U10517 ( .A1(n9152), .A2(n9151), .A3(n9150), .ZN(P1_U3222) );
  XOR2_X1 U10518 ( .A(n9154), .B(n9153), .Z(n9159) );
  AOI22_X1 U10519 ( .A1(n9276), .A2(n9802), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9156) );
  NAND2_X1 U10520 ( .A1(n9267), .A2(n9498), .ZN(n9155) );
  OAI211_X1 U10521 ( .C1(n9489), .C2(n9803), .A(n9156), .B(n9155), .ZN(n9157)
         );
  AOI21_X1 U10522 ( .B1(n9739), .B2(n6649), .A(n9157), .ZN(n9158) );
  OAI21_X1 U10523 ( .B1(n9159), .B2(n9245), .A(n9158), .ZN(P1_U3223) );
  OAI21_X1 U10524 ( .B1(n9162), .B2(n9161), .A(n9160), .ZN(n9163) );
  NAND2_X1 U10525 ( .A1(n9163), .A2(n9809), .ZN(n9168) );
  NAND2_X1 U10526 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n9838) );
  OAI21_X1 U10527 ( .B1(n9265), .B2(n9164), .A(n9838), .ZN(n9165) );
  AOI21_X1 U10528 ( .B1(n9267), .B2(n9166), .A(n9165), .ZN(n9167) );
  OAI211_X1 U10529 ( .C1(n9169), .C2(n9800), .A(n9168), .B(n9167), .ZN(
        P1_U3224) );
  AOI21_X1 U10530 ( .B1(n9171), .B2(n9170), .A(n4355), .ZN(n9179) );
  OAI22_X1 U10531 ( .A1(n9173), .A2(n9490), .B1(n9172), .B2(n9488), .ZN(n9425)
         );
  INV_X1 U10532 ( .A(n9430), .ZN(n9175) );
  OAI22_X1 U10533 ( .A1(n9175), .A2(n9814), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9174), .ZN(n9177) );
  NOR2_X1 U10534 ( .A1(n9722), .A2(n9800), .ZN(n9176) );
  AOI211_X1 U10535 ( .C1(n9254), .C2(n9425), .A(n9177), .B(n9176), .ZN(n9178)
         );
  OAI21_X1 U10536 ( .B1(n9179), .B2(n9245), .A(n9178), .ZN(P1_U3225) );
  INV_X1 U10537 ( .A(n9761), .ZN(n9577) );
  NAND2_X1 U10538 ( .A1(n9259), .A2(n9182), .ZN(n9183) );
  INV_X1 U10539 ( .A(n9187), .ZN(n9184) );
  NOR2_X1 U10540 ( .A1(n9185), .A2(n9184), .ZN(n9190) );
  NAND2_X1 U10541 ( .A1(n9259), .A2(n9258), .ZN(n9257) );
  NAND2_X1 U10542 ( .A1(n9257), .A2(n9180), .ZN(n9186) );
  AOI21_X1 U10543 ( .B1(n9188), .B2(n9187), .A(n9186), .ZN(n9189) );
  OAI21_X1 U10544 ( .B1(n9190), .B2(n9189), .A(n9809), .ZN(n9195) );
  NAND2_X1 U10545 ( .A1(n9281), .A2(n9523), .ZN(n9192) );
  NAND2_X1 U10546 ( .A1(n9279), .A2(n9524), .ZN(n9191) );
  AND2_X1 U10547 ( .A1(n9192), .A2(n9191), .ZN(n9572) );
  NAND2_X1 U10548 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9324) );
  OAI21_X1 U10549 ( .B1(n9265), .B2(n9572), .A(n9324), .ZN(n9193) );
  AOI21_X1 U10550 ( .B1(n9267), .B2(n9578), .A(n9193), .ZN(n9194) );
  OAI211_X1 U10551 ( .C1(n9577), .C2(n9800), .A(n9195), .B(n9194), .ZN(
        P1_U3226) );
  OAI21_X1 U10552 ( .B1(n9198), .B2(n9197), .A(n9196), .ZN(n9199) );
  NAND2_X1 U10553 ( .A1(n9199), .A2(n9809), .ZN(n9204) );
  OR2_X1 U10554 ( .A1(n9261), .A2(n9488), .ZN(n9201) );
  NAND2_X1 U10555 ( .A1(n9522), .A2(n9524), .ZN(n9200) );
  AND2_X1 U10556 ( .A1(n9201), .A2(n9200), .ZN(n9558) );
  NAND2_X1 U10557 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9854) );
  OAI21_X1 U10558 ( .B1(n9265), .B2(n9558), .A(n9854), .ZN(n9202) );
  AOI21_X1 U10559 ( .B1(n9267), .B2(n9562), .A(n9202), .ZN(n9203) );
  OAI211_X1 U10560 ( .C1(n9760), .C2(n9800), .A(n9204), .B(n9203), .ZN(
        P1_U3228) );
  XNOR2_X1 U10561 ( .A(n9206), .B(n9205), .ZN(n9207) );
  XNOR2_X1 U10562 ( .A(n9208), .B(n9207), .ZN(n9214) );
  NAND2_X1 U10563 ( .A1(n9277), .A2(n9524), .ZN(n9210) );
  NAND2_X1 U10564 ( .A1(n9278), .A2(n9523), .ZN(n9209) );
  NAND2_X1 U10565 ( .A1(n9210), .A2(n9209), .ZN(n9507) );
  AOI22_X1 U10566 ( .A1(n9507), .A2(n9254), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9211) );
  OAI21_X1 U10567 ( .B1(n9814), .B2(n9511), .A(n9211), .ZN(n9212) );
  AOI21_X1 U10568 ( .B1(n9744), .B2(n6649), .A(n9212), .ZN(n9213) );
  OAI21_X1 U10569 ( .B1(n9214), .B2(n9245), .A(n9213), .ZN(P1_U3233) );
  OAI21_X1 U10570 ( .B1(n9217), .B2(n9216), .A(n9215), .ZN(n9218) );
  NAND2_X1 U10571 ( .A1(n9218), .A2(n9809), .ZN(n9224) );
  OAI21_X1 U10572 ( .B1(n9265), .B2(n9220), .A(n9219), .ZN(n9221) );
  AOI21_X1 U10573 ( .B1(n9267), .B2(n9222), .A(n9221), .ZN(n9223) );
  OAI211_X1 U10574 ( .C1(n9225), .C2(n9800), .A(n9224), .B(n9223), .ZN(
        P1_U3234) );
  INV_X1 U10575 ( .A(n9226), .ZN(n9227) );
  NAND2_X1 U10576 ( .A1(n9227), .A2(n9230), .ZN(n9228) );
  AOI22_X1 U10577 ( .A1(n9231), .A2(n9230), .B1(n9229), .B2(n9228), .ZN(n9237)
         );
  NAND2_X1 U10578 ( .A1(n9275), .A2(n9524), .ZN(n9233) );
  NAND2_X1 U10579 ( .A1(n9277), .A2(n9523), .ZN(n9232) );
  NAND2_X1 U10580 ( .A1(n9233), .A2(n9232), .ZN(n9471) );
  AOI22_X1 U10581 ( .A1(n9471), .A2(n9254), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9234) );
  OAI21_X1 U10582 ( .B1(n9814), .B2(n9476), .A(n9234), .ZN(n9235) );
  AOI21_X1 U10583 ( .B1(n9734), .B2(n6649), .A(n9235), .ZN(n9236) );
  OAI21_X1 U10584 ( .B1(n9237), .B2(n9245), .A(n9236), .ZN(P1_U3235) );
  AOI21_X1 U10585 ( .B1(n9240), .B2(n9239), .A(n9238), .ZN(n9246) );
  NOR2_X1 U10586 ( .A1(n9814), .A2(n9545), .ZN(n9243) );
  AND2_X1 U10587 ( .A1(n9279), .A2(n9523), .ZN(n9241) );
  AOI21_X1 U10588 ( .B1(n9278), .B2(n9524), .A(n9241), .ZN(n9537) );
  NAND2_X1 U10589 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9342) );
  OAI21_X1 U10590 ( .B1(n9537), .B2(n9265), .A(n9342), .ZN(n9242) );
  AOI211_X1 U10591 ( .C1(n9751), .C2(n6649), .A(n9243), .B(n9242), .ZN(n9244)
         );
  OAI21_X1 U10592 ( .B1(n9246), .B2(n9245), .A(n9244), .ZN(P1_U3238) );
  OAI21_X1 U10593 ( .B1(n4355), .B2(n9248), .A(n9247), .ZN(n9249) );
  NAND3_X1 U10594 ( .A1(n4356), .A2(n9809), .A3(n9249), .ZN(n9256) );
  OAI22_X1 U10595 ( .A1(n9251), .A2(n9490), .B1(n9250), .B2(n9488), .ZN(n9410)
         );
  OAI22_X1 U10596 ( .A1(n9414), .A2(n9814), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9252), .ZN(n9253) );
  AOI21_X1 U10597 ( .B1(n9410), .B2(n9254), .A(n9253), .ZN(n9255) );
  OAI211_X1 U10598 ( .C1(n9413), .C2(n9800), .A(n9256), .B(n9255), .ZN(
        P1_U3240) );
  OAI21_X1 U10599 ( .B1(n9259), .B2(n9258), .A(n9257), .ZN(n9260) );
  NAND2_X1 U10600 ( .A1(n9260), .A2(n9809), .ZN(n9269) );
  OR2_X1 U10601 ( .A1(n9261), .A2(n9490), .ZN(n9263) );
  NAND2_X1 U10602 ( .A1(n9282), .A2(n9523), .ZN(n9262) );
  AND2_X1 U10603 ( .A1(n9263), .A2(n9262), .ZN(n9591) );
  OAI21_X1 U10604 ( .B1(n9265), .B2(n9591), .A(n9264), .ZN(n9266) );
  AOI21_X1 U10605 ( .B1(n9267), .B2(n9596), .A(n9266), .ZN(n9268) );
  OAI211_X1 U10606 ( .C1(n9599), .C2(n9800), .A(n9269), .B(n9268), .ZN(
        P1_U3241) );
  MUX2_X1 U10607 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9270), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10608 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9271), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10609 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9272), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10610 ( .A(n9395), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9294), .Z(
        P1_U3580) );
  MUX2_X1 U10611 ( .A(n9273), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9294), .Z(
        P1_U3579) );
  MUX2_X1 U10612 ( .A(n9274), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9294), .Z(
        P1_U3578) );
  MUX2_X1 U10613 ( .A(n9275), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9294), .Z(
        P1_U3577) );
  MUX2_X1 U10614 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9276), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10615 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9277), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10616 ( .A(n9525), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9294), .Z(
        P1_U3574) );
  MUX2_X1 U10617 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9278), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10618 ( .A(n9522), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9294), .Z(
        P1_U3572) );
  MUX2_X1 U10619 ( .A(n9279), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9294), .Z(
        P1_U3571) );
  MUX2_X1 U10620 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9280), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10621 ( .A(n9281), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9294), .Z(
        P1_U3569) );
  MUX2_X1 U10622 ( .A(n9282), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9294), .Z(
        P1_U3568) );
  MUX2_X1 U10623 ( .A(n9283), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9294), .Z(
        P1_U3567) );
  MUX2_X1 U10624 ( .A(n9284), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9294), .Z(
        P1_U3566) );
  MUX2_X1 U10625 ( .A(n9285), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9294), .Z(
        P1_U3565) );
  MUX2_X1 U10626 ( .A(n9286), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9294), .Z(
        P1_U3564) );
  MUX2_X1 U10627 ( .A(n9287), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9294), .Z(
        P1_U3563) );
  MUX2_X1 U10628 ( .A(n9288), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9294), .Z(
        P1_U3562) );
  MUX2_X1 U10629 ( .A(n9289), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9294), .Z(
        P1_U3560) );
  MUX2_X1 U10630 ( .A(n9290), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9294), .Z(
        P1_U3559) );
  MUX2_X1 U10631 ( .A(n9291), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9294), .Z(
        P1_U3558) );
  MUX2_X1 U10632 ( .A(n9292), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9294), .Z(
        P1_U3557) );
  MUX2_X1 U10633 ( .A(n9293), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9294), .Z(
        P1_U3556) );
  MUX2_X1 U10634 ( .A(n7140), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9294), .Z(
        P1_U3555) );
  INV_X1 U10635 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9295) );
  OAI22_X1 U10636 ( .A1(n9857), .A2(n9296), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9295), .ZN(n9297) );
  AOI21_X1 U10637 ( .B1(n9298), .B2(n9332), .A(n9297), .ZN(n9308) );
  MUX2_X1 U10638 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6773), .S(n9299), .Z(n9300)
         );
  OAI21_X1 U10639 ( .B1(n9816), .B2(n9819), .A(n9300), .ZN(n9301) );
  NAND3_X1 U10640 ( .A1(n9340), .A2(n9302), .A3(n9301), .ZN(n9307) );
  OAI211_X1 U10641 ( .C1(n9305), .C2(n9304), .A(n9853), .B(n9303), .ZN(n9306)
         );
  NAND3_X1 U10642 ( .A1(n9308), .A2(n9307), .A3(n9306), .ZN(P1_U3244) );
  AOI211_X1 U10643 ( .C1(n9311), .C2(n9310), .A(n9309), .B(n9849), .ZN(n9312)
         );
  INV_X1 U10644 ( .A(n9312), .ZN(n9320) );
  AOI22_X1 U10645 ( .A1(n9824), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(P1_U3086), .ZN(n9319) );
  NAND2_X1 U10646 ( .A1(n9332), .A2(n9313), .ZN(n9318) );
  OAI211_X1 U10647 ( .C1(n9316), .C2(n9315), .A(n9853), .B(n9314), .ZN(n9317)
         );
  NAND4_X1 U10648 ( .A1(n9320), .A2(n9319), .A3(n9318), .A4(n9317), .ZN(
        P1_U3246) );
  AOI21_X1 U10649 ( .B1(n9323), .B2(n9322), .A(n9321), .ZN(n9335) );
  INV_X1 U10650 ( .A(n9324), .ZN(n9330) );
  INV_X1 U10651 ( .A(n9325), .ZN(n9326) );
  AOI211_X1 U10652 ( .C1(n9328), .C2(n9327), .A(n9326), .B(n9343), .ZN(n9329)
         );
  AOI211_X1 U10653 ( .C1(n9824), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9330), .B(
        n9329), .ZN(n9334) );
  NAND2_X1 U10654 ( .A1(n9332), .A2(n9331), .ZN(n9333) );
  OAI211_X1 U10655 ( .C1(n9335), .C2(n9849), .A(n9334), .B(n9333), .ZN(
        P1_U3259) );
  INV_X1 U10656 ( .A(n9336), .ZN(n9341) );
  OAI21_X1 U10657 ( .B1(n9844), .B2(n9338), .A(n9337), .ZN(n9339) );
  NAND3_X1 U10658 ( .A1(n9341), .A2(n9340), .A3(n9339), .ZN(n9350) );
  INV_X1 U10659 ( .A(n9342), .ZN(n9348) );
  AOI211_X1 U10660 ( .C1(n9346), .C2(n9345), .A(n9344), .B(n9343), .ZN(n9347)
         );
  AOI211_X1 U10661 ( .C1(n9824), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9348), .B(
        n9347), .ZN(n9349) );
  OAI211_X1 U10662 ( .C1(n9847), .C2(n9351), .A(n9350), .B(n9349), .ZN(
        P1_U3261) );
  XOR2_X1 U10663 ( .A(n9359), .B(n9352), .Z(n9353) );
  NOR2_X1 U10664 ( .A1(n9353), .A2(n9595), .ZN(n9627) );
  NAND2_X1 U10665 ( .A1(n9627), .A2(n9858), .ZN(n9358) );
  NOR2_X1 U10666 ( .A1(n9355), .A2(n9354), .ZN(n9630) );
  INV_X1 U10667 ( .A(n9630), .ZN(n9356) );
  NOR2_X1 U10668 ( .A1(n9617), .A2(n9356), .ZN(n9363) );
  AOI21_X1 U10669 ( .B1(n9617), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9363), .ZN(
        n9357) );
  OAI211_X1 U10670 ( .C1(n9703), .C2(n9865), .A(n9358), .B(n9357), .ZN(
        P1_U3263) );
  AOI211_X1 U10671 ( .C1(n9361), .C2(n9360), .A(n9595), .B(n9359), .ZN(n9631)
         );
  NAND2_X1 U10672 ( .A1(n9631), .A2(n9858), .ZN(n9365) );
  AND2_X1 U10673 ( .A1(n9617), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9362) );
  NOR2_X1 U10674 ( .A1(n9363), .A2(n9362), .ZN(n9364) );
  OAI211_X1 U10675 ( .C1(n9707), .C2(n9865), .A(n9365), .B(n9364), .ZN(
        P1_U3264) );
  NAND2_X1 U10676 ( .A1(n9366), .A2(n9868), .ZN(n9374) );
  INV_X1 U10677 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9367) );
  OAI22_X1 U10678 ( .A1(n9368), .A2(n9544), .B1(n9367), .B2(n9623), .ZN(n9371)
         );
  NOR2_X1 U10679 ( .A1(n9369), .A2(n9621), .ZN(n9370) );
  AOI211_X1 U10680 ( .C1(n9618), .C2(n9372), .A(n9371), .B(n9370), .ZN(n9373)
         );
  OAI211_X1 U10681 ( .C1(n9375), .C2(n9617), .A(n9374), .B(n9373), .ZN(
        P1_U3356) );
  NAND2_X1 U10682 ( .A1(n9384), .A2(n9383), .ZN(n9635) );
  INV_X1 U10683 ( .A(n9709), .ZN(n9389) );
  NAND2_X1 U10684 ( .A1(n9634), .A2(n9858), .ZN(n9388) );
  AOI22_X1 U10685 ( .A1(n9386), .A2(n9861), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9617), .ZN(n9387) );
  OAI211_X1 U10686 ( .C1(n9389), .C2(n9865), .A(n9388), .B(n9387), .ZN(n9390)
         );
  AOI21_X1 U10687 ( .B1(n9623), .B2(n9635), .A(n9390), .ZN(n9391) );
  OAI21_X1 U10688 ( .B1(n9710), .B2(n9626), .A(n9391), .ZN(P1_U3265) );
  XNOR2_X1 U10689 ( .A(n9376), .B(n9393), .ZN(n9641) );
  INV_X1 U10690 ( .A(n9641), .ZN(n9406) );
  NAND2_X1 U10691 ( .A1(n9395), .A2(n9523), .ZN(n9396) );
  AOI211_X1 U10692 ( .C1(n9399), .C2(n9412), .A(n9595), .B(n9385), .ZN(n9640)
         );
  NAND2_X1 U10693 ( .A1(n9640), .A2(n9858), .ZN(n9403) );
  INV_X1 U10694 ( .A(n9400), .ZN(n9401) );
  AOI22_X1 U10695 ( .A1(n9401), .A2(n9861), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9617), .ZN(n9402) );
  OAI211_X1 U10696 ( .C1(n9713), .C2(n9865), .A(n9403), .B(n9402), .ZN(n9404)
         );
  AOI21_X1 U10697 ( .B1(n9639), .B2(n9623), .A(n9404), .ZN(n9405) );
  OAI21_X1 U10698 ( .B1(n9406), .B2(n9626), .A(n9405), .ZN(P1_U3266) );
  XNOR2_X1 U10699 ( .A(n9407), .B(n9408), .ZN(n9718) );
  XNOR2_X1 U10700 ( .A(n9409), .B(n9408), .ZN(n9411) );
  AOI21_X1 U10701 ( .B1(n9411), .B2(n9608), .A(n9410), .ZN(n9644) );
  INV_X1 U10702 ( .A(n9644), .ZN(n9419) );
  OAI211_X1 U10703 ( .C1(n9413), .C2(n9428), .A(n9613), .B(n9412), .ZN(n9643)
         );
  INV_X1 U10704 ( .A(n9414), .ZN(n9415) );
  AOI22_X1 U10705 ( .A1(n9415), .A2(n9861), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9617), .ZN(n9417) );
  NAND2_X1 U10706 ( .A1(n9716), .A2(n9618), .ZN(n9416) );
  OAI211_X1 U10707 ( .C1(n9643), .C2(n9621), .A(n9417), .B(n9416), .ZN(n9418)
         );
  AOI21_X1 U10708 ( .B1(n9419), .B2(n9623), .A(n9418), .ZN(n9420) );
  OAI21_X1 U10709 ( .B1(n9718), .B2(n9626), .A(n9420), .ZN(P1_U3267) );
  XOR2_X1 U10710 ( .A(n9423), .B(n9421), .Z(n9649) );
  INV_X1 U10711 ( .A(n9649), .ZN(n9435) );
  OAI211_X1 U10712 ( .C1(n9424), .C2(n9423), .A(n9422), .B(n9608), .ZN(n9427)
         );
  INV_X1 U10713 ( .A(n9425), .ZN(n9426) );
  NAND2_X1 U10714 ( .A1(n9427), .A2(n9426), .ZN(n9647) );
  OAI21_X1 U10715 ( .B1(n9722), .B2(n9443), .A(n9613), .ZN(n9429) );
  NOR2_X1 U10716 ( .A1(n9429), .A2(n9428), .ZN(n9648) );
  NAND2_X1 U10717 ( .A1(n9648), .A2(n9858), .ZN(n9432) );
  AOI22_X1 U10718 ( .A1(n9430), .A2(n9861), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9617), .ZN(n9431) );
  OAI211_X1 U10719 ( .C1(n9722), .C2(n9865), .A(n9432), .B(n9431), .ZN(n9433)
         );
  AOI21_X1 U10720 ( .B1(n9623), .B2(n9647), .A(n9433), .ZN(n9434) );
  OAI21_X1 U10721 ( .B1(n9435), .B2(n9626), .A(n9434), .ZN(P1_U3268) );
  XNOR2_X1 U10722 ( .A(n9436), .B(n9438), .ZN(n9727) );
  INV_X1 U10723 ( .A(n9437), .ZN(n9439) );
  AOI21_X1 U10724 ( .B1(n9439), .B2(n9438), .A(n9592), .ZN(n9442) );
  AOI21_X1 U10725 ( .B1(n9442), .B2(n9441), .A(n9440), .ZN(n9653) );
  INV_X1 U10726 ( .A(n9653), .ZN(n9451) );
  INV_X1 U10727 ( .A(n5088), .ZN(n9461) );
  INV_X1 U10728 ( .A(n9443), .ZN(n9444) );
  OAI211_X1 U10729 ( .C1(n9445), .C2(n9461), .A(n9444), .B(n9613), .ZN(n9652)
         );
  INV_X1 U10730 ( .A(n9446), .ZN(n9447) );
  AOI22_X1 U10731 ( .A1(n9447), .A2(n9861), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9617), .ZN(n9449) );
  NAND2_X1 U10732 ( .A1(n9725), .A2(n9618), .ZN(n9448) );
  OAI211_X1 U10733 ( .C1(n9652), .C2(n9621), .A(n9449), .B(n9448), .ZN(n9450)
         );
  AOI21_X1 U10734 ( .B1(n9451), .B2(n9623), .A(n9450), .ZN(n9452) );
  OAI21_X1 U10735 ( .B1(n9727), .B2(n9626), .A(n9452), .ZN(P1_U3269) );
  XOR2_X1 U10736 ( .A(n9456), .B(n9453), .Z(n9658) );
  INV_X1 U10737 ( .A(n9658), .ZN(n9469) );
  AND2_X1 U10738 ( .A1(n9472), .A2(n9454), .ZN(n9455) );
  XNOR2_X1 U10739 ( .A(n9456), .B(n9455), .ZN(n9457) );
  NAND2_X1 U10740 ( .A1(n9457), .A2(n9608), .ZN(n9460) );
  INV_X1 U10741 ( .A(n9458), .ZN(n9459) );
  NAND2_X1 U10742 ( .A1(n9460), .A2(n9459), .ZN(n9656) );
  AOI211_X1 U10743 ( .C1(n9462), .C2(n9478), .A(n9595), .B(n9461), .ZN(n9657)
         );
  NAND2_X1 U10744 ( .A1(n9657), .A2(n9858), .ZN(n9466) );
  INV_X1 U10745 ( .A(n9463), .ZN(n9464) );
  AOI22_X1 U10746 ( .A1(n9464), .A2(n9861), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9617), .ZN(n9465) );
  OAI211_X1 U10747 ( .C1(n9731), .C2(n9865), .A(n9466), .B(n9465), .ZN(n9467)
         );
  AOI21_X1 U10748 ( .B1(n9623), .B2(n9656), .A(n9467), .ZN(n9468) );
  OAI21_X1 U10749 ( .B1(n9469), .B2(n9626), .A(n9468), .ZN(P1_U3270) );
  AOI21_X1 U10750 ( .B1(n9474), .B2(n9470), .A(n9592), .ZN(n9473) );
  AOI21_X1 U10751 ( .B1(n9473), .B2(n9472), .A(n9471), .ZN(n9662) );
  XNOR2_X1 U10752 ( .A(n4395), .B(n9474), .ZN(n9736) );
  INV_X1 U10753 ( .A(n9736), .ZN(n9475) );
  NAND2_X1 U10754 ( .A1(n9475), .A2(n9868), .ZN(n9483) );
  INV_X1 U10755 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9477) );
  OAI22_X1 U10756 ( .A1(n9623), .A2(n9477), .B1(n9476), .B2(n9544), .ZN(n9481)
         );
  OAI211_X1 U10757 ( .C1(n9479), .C2(n9494), .A(n9613), .B(n9478), .ZN(n9661)
         );
  NOR2_X1 U10758 ( .A1(n9661), .A2(n9621), .ZN(n9480) );
  AOI211_X1 U10759 ( .C1(n9618), .C2(n9734), .A(n9481), .B(n9480), .ZN(n9482)
         );
  OAI211_X1 U10760 ( .C1(n9617), .C2(n9662), .A(n9483), .B(n9482), .ZN(
        P1_U3271) );
  XOR2_X1 U10761 ( .A(n9486), .B(n9484), .Z(n9741) );
  OR2_X1 U10762 ( .A1(n9506), .A2(n9505), .ZN(n9508) );
  AND2_X1 U10763 ( .A1(n9508), .A2(n9485), .ZN(n9487) );
  XNOR2_X1 U10764 ( .A(n9487), .B(n9486), .ZN(n9493) );
  OAI22_X1 U10765 ( .A1(n9491), .A2(n9490), .B1(n9489), .B2(n9488), .ZN(n9492)
         );
  AOI21_X1 U10766 ( .B1(n9493), .B2(n9608), .A(n9492), .ZN(n9666) );
  INV_X1 U10767 ( .A(n9666), .ZN(n9502) );
  INV_X1 U10768 ( .A(n9510), .ZN(n9496) );
  INV_X1 U10769 ( .A(n9494), .ZN(n9495) );
  OAI211_X1 U10770 ( .C1(n9497), .C2(n9496), .A(n9495), .B(n9613), .ZN(n9665)
         );
  AOI22_X1 U10771 ( .A1(n9617), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9498), .B2(
        n9861), .ZN(n9500) );
  NAND2_X1 U10772 ( .A1(n9739), .A2(n9618), .ZN(n9499) );
  OAI211_X1 U10773 ( .C1(n9665), .C2(n9621), .A(n9500), .B(n9499), .ZN(n9501)
         );
  AOI21_X1 U10774 ( .B1(n9502), .B2(n9623), .A(n9501), .ZN(n9503) );
  OAI21_X1 U10775 ( .B1(n9741), .B2(n9626), .A(n9503), .ZN(P1_U3272) );
  XNOR2_X1 U10776 ( .A(n9504), .B(n9505), .ZN(n9746) );
  AOI21_X1 U10777 ( .B1(n9506), .B2(n9505), .A(n9592), .ZN(n9509) );
  AOI21_X1 U10778 ( .B1(n9509), .B2(n9508), .A(n9507), .ZN(n9670) );
  INV_X1 U10779 ( .A(n9670), .ZN(n9516) );
  OAI211_X1 U10780 ( .C1(n4765), .C2(n4766), .A(n9510), .B(n9613), .ZN(n9669)
         );
  INV_X1 U10781 ( .A(n9511), .ZN(n9512) );
  AOI22_X1 U10782 ( .A1(n9617), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9512), .B2(
        n9861), .ZN(n9514) );
  NAND2_X1 U10783 ( .A1(n9744), .A2(n9618), .ZN(n9513) );
  OAI211_X1 U10784 ( .C1(n9669), .C2(n9621), .A(n9514), .B(n9513), .ZN(n9515)
         );
  AOI21_X1 U10785 ( .B1(n9516), .B2(n9623), .A(n9515), .ZN(n9517) );
  OAI21_X1 U10786 ( .B1(n9746), .B2(n9626), .A(n9517), .ZN(P1_U3273) );
  XNOR2_X1 U10787 ( .A(n9518), .B(n9520), .ZN(n9675) );
  INV_X1 U10788 ( .A(n9675), .ZN(n9535) );
  XNOR2_X1 U10789 ( .A(n9520), .B(n9519), .ZN(n9521) );
  NAND2_X1 U10790 ( .A1(n9521), .A2(n9608), .ZN(n9527) );
  AOI22_X1 U10791 ( .A1(n9525), .A2(n9524), .B1(n9523), .B2(n9522), .ZN(n9526)
         );
  NAND2_X1 U10792 ( .A1(n9527), .A2(n9526), .ZN(n9673) );
  AOI211_X1 U10793 ( .C1(n9528), .C2(n9547), .A(n9595), .B(n4766), .ZN(n9674)
         );
  NAND2_X1 U10794 ( .A1(n9674), .A2(n9858), .ZN(n9532) );
  INV_X1 U10795 ( .A(n9529), .ZN(n9530) );
  AOI22_X1 U10796 ( .A1(n9617), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9530), .B2(
        n9861), .ZN(n9531) );
  OAI211_X1 U10797 ( .C1(n9750), .C2(n9865), .A(n9532), .B(n9531), .ZN(n9533)
         );
  AOI21_X1 U10798 ( .B1(n9623), .B2(n9673), .A(n9533), .ZN(n9534) );
  OAI21_X1 U10799 ( .B1(n9535), .B2(n9626), .A(n9534), .ZN(P1_U3274) );
  XNOR2_X1 U10800 ( .A(n9536), .B(n9541), .ZN(n9539) );
  INV_X1 U10801 ( .A(n9537), .ZN(n9538) );
  AOI21_X1 U10802 ( .B1(n9539), .B2(n9608), .A(n9538), .ZN(n9679) );
  INV_X1 U10803 ( .A(n9540), .ZN(n9542) );
  XNOR2_X1 U10804 ( .A(n9542), .B(n9541), .ZN(n9755) );
  INV_X1 U10805 ( .A(n9755), .ZN(n9543) );
  NAND2_X1 U10806 ( .A1(n9543), .A2(n9868), .ZN(n9552) );
  OAI22_X1 U10807 ( .A1(n9623), .A2(n9546), .B1(n9545), .B2(n9544), .ZN(n9550)
         );
  OAI211_X1 U10808 ( .C1(n9548), .C2(n9560), .A(n9613), .B(n9547), .ZN(n9678)
         );
  NOR2_X1 U10809 ( .A1(n9678), .A2(n9621), .ZN(n9549) );
  AOI211_X1 U10810 ( .C1(n9618), .C2(n9751), .A(n9550), .B(n9549), .ZN(n9551)
         );
  OAI211_X1 U10811 ( .C1(n9617), .C2(n9679), .A(n9552), .B(n9551), .ZN(
        P1_U3275) );
  XNOR2_X1 U10812 ( .A(n9553), .B(n9554), .ZN(n9684) );
  INV_X1 U10813 ( .A(n9684), .ZN(n9567) );
  NAND2_X1 U10814 ( .A1(n9555), .A2(n9554), .ZN(n9556) );
  NAND3_X1 U10815 ( .A1(n9557), .A2(n9608), .A3(n9556), .ZN(n9559) );
  NAND2_X1 U10816 ( .A1(n9559), .A2(n9558), .ZN(n9682) );
  AOI211_X1 U10817 ( .C1(n9561), .C2(n9576), .A(n9595), .B(n9560), .ZN(n9683)
         );
  NAND2_X1 U10818 ( .A1(n9683), .A2(n9858), .ZN(n9564) );
  AOI22_X1 U10819 ( .A1(n9617), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9562), .B2(
        n9861), .ZN(n9563) );
  OAI211_X1 U10820 ( .C1(n9760), .C2(n9865), .A(n9564), .B(n9563), .ZN(n9565)
         );
  AOI21_X1 U10821 ( .B1(n9623), .B2(n9682), .A(n9565), .ZN(n9566) );
  OAI21_X1 U10822 ( .B1(n9567), .B2(n9626), .A(n9566), .ZN(P1_U3276) );
  XNOR2_X1 U10823 ( .A(n9568), .B(n9569), .ZN(n9765) );
  XNOR2_X1 U10824 ( .A(n9571), .B(n9570), .ZN(n9574) );
  INV_X1 U10825 ( .A(n9572), .ZN(n9573) );
  AOI21_X1 U10826 ( .B1(n9574), .B2(n9608), .A(n9573), .ZN(n9688) );
  INV_X1 U10827 ( .A(n9688), .ZN(n9582) );
  INV_X1 U10828 ( .A(n9575), .ZN(n9594) );
  OAI211_X1 U10829 ( .C1(n9577), .C2(n9594), .A(n9613), .B(n9576), .ZN(n9687)
         );
  AOI22_X1 U10830 ( .A1(n9617), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9578), .B2(
        n9861), .ZN(n9580) );
  NAND2_X1 U10831 ( .A1(n9761), .A2(n9618), .ZN(n9579) );
  OAI211_X1 U10832 ( .C1(n9687), .C2(n9621), .A(n9580), .B(n9579), .ZN(n9581)
         );
  AOI21_X1 U10833 ( .B1(n9582), .B2(n9623), .A(n9581), .ZN(n9583) );
  OAI21_X1 U10834 ( .B1(n9765), .B2(n9626), .A(n9583), .ZN(P1_U3277) );
  XOR2_X1 U10835 ( .A(n9585), .B(n9590), .Z(n9693) );
  INV_X1 U10836 ( .A(n9693), .ZN(n9602) );
  NAND2_X1 U10837 ( .A1(n9609), .A2(n9586), .ZN(n9589) );
  INV_X1 U10838 ( .A(n9587), .ZN(n9588) );
  AOI21_X1 U10839 ( .B1(n9590), .B2(n9589), .A(n9588), .ZN(n9593) );
  OAI21_X1 U10840 ( .B1(n9593), .B2(n9592), .A(n9591), .ZN(n9691) );
  AOI211_X1 U10841 ( .C1(n9766), .C2(n9614), .A(n9595), .B(n9594), .ZN(n9692)
         );
  NAND2_X1 U10842 ( .A1(n9692), .A2(n9858), .ZN(n9598) );
  AOI22_X1 U10843 ( .A1(n9617), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9596), .B2(
        n9861), .ZN(n9597) );
  OAI211_X1 U10844 ( .C1(n9599), .C2(n9865), .A(n9598), .B(n9597), .ZN(n9600)
         );
  AOI21_X1 U10845 ( .B1(n9691), .B2(n9623), .A(n9600), .ZN(n9601) );
  OAI21_X1 U10846 ( .B1(n9602), .B2(n9626), .A(n9601), .ZN(P1_U3278) );
  XOR2_X1 U10847 ( .A(n9603), .B(n9606), .Z(n9775) );
  NAND2_X1 U10848 ( .A1(n9605), .A2(n9604), .ZN(n9607) );
  NAND2_X1 U10849 ( .A1(n9607), .A2(n9606), .ZN(n9610) );
  NAND3_X1 U10850 ( .A1(n9610), .A2(n9609), .A3(n9608), .ZN(n9612) );
  AND2_X1 U10851 ( .A1(n9612), .A2(n9611), .ZN(n9697) );
  INV_X1 U10852 ( .A(n9697), .ZN(n9624) );
  OAI211_X1 U10853 ( .C1(n4420), .C2(n9615), .A(n9614), .B(n9613), .ZN(n9696)
         );
  AOI22_X1 U10854 ( .A1(n9617), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9616), .B2(
        n9861), .ZN(n9620) );
  NAND2_X1 U10855 ( .A1(n9770), .A2(n9618), .ZN(n9619) );
  OAI211_X1 U10856 ( .C1(n9696), .C2(n9621), .A(n9620), .B(n9619), .ZN(n9622)
         );
  AOI21_X1 U10857 ( .B1(n9624), .B2(n9623), .A(n9622), .ZN(n9625) );
  OAI21_X1 U10858 ( .B1(n9775), .B2(n9626), .A(n9625), .ZN(P1_U3279) );
  INV_X1 U10859 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9628) );
  NOR2_X1 U10860 ( .A1(n9627), .A2(n9630), .ZN(n9701) );
  MUX2_X1 U10861 ( .A(n9628), .B(n9701), .S(n9896), .Z(n9629) );
  OAI21_X1 U10862 ( .B1(n9703), .B2(n9686), .A(n9629), .ZN(P1_U3553) );
  INV_X1 U10863 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9632) );
  NOR2_X1 U10864 ( .A1(n9631), .A2(n9630), .ZN(n9704) );
  MUX2_X1 U10865 ( .A(n9632), .B(n9704), .S(n9896), .Z(n9633) );
  OAI21_X1 U10866 ( .B1(n9707), .B2(n9686), .A(n9633), .ZN(P1_U3552) );
  NOR2_X1 U10867 ( .A1(n9635), .A2(n9634), .ZN(n9708) );
  MUX2_X1 U10868 ( .A(n9636), .B(n9708), .S(n9896), .Z(n9638) );
  NAND2_X1 U10869 ( .A1(n9709), .A2(n9695), .ZN(n9637) );
  OAI211_X1 U10870 ( .C1(n9710), .C2(n9700), .A(n9638), .B(n9637), .ZN(
        P1_U3550) );
  NAND2_X1 U10871 ( .A1(n9644), .A2(n9643), .ZN(n9714) );
  MUX2_X1 U10872 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9714), .S(n9896), .Z(n9645) );
  AOI21_X1 U10873 ( .B1(n9695), .B2(n9716), .A(n9645), .ZN(n9646) );
  OAI21_X1 U10874 ( .B1(n9718), .B2(n9700), .A(n9646), .ZN(P1_U3548) );
  AOI211_X1 U10875 ( .C1(n9649), .C2(n9878), .A(n9648), .B(n9647), .ZN(n9719)
         );
  MUX2_X1 U10876 ( .A(n9650), .B(n9719), .S(n9896), .Z(n9651) );
  OAI21_X1 U10877 ( .B1(n9722), .B2(n9686), .A(n9651), .ZN(P1_U3547) );
  NAND2_X1 U10878 ( .A1(n9653), .A2(n9652), .ZN(n9723) );
  MUX2_X1 U10879 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9723), .S(n9896), .Z(n9654) );
  AOI21_X1 U10880 ( .B1(n9695), .B2(n9725), .A(n9654), .ZN(n9655) );
  OAI21_X1 U10881 ( .B1(n9727), .B2(n9700), .A(n9655), .ZN(P1_U3546) );
  AOI211_X1 U10882 ( .C1(n9658), .C2(n9878), .A(n9657), .B(n9656), .ZN(n9728)
         );
  MUX2_X1 U10883 ( .A(n9659), .B(n9728), .S(n9896), .Z(n9660) );
  OAI21_X1 U10884 ( .B1(n9731), .B2(n9686), .A(n9660), .ZN(P1_U3545) );
  NAND2_X1 U10885 ( .A1(n9662), .A2(n9661), .ZN(n9732) );
  MUX2_X1 U10886 ( .A(n9732), .B(P1_REG1_REG_22__SCAN_IN), .S(n9893), .Z(n9663) );
  AOI21_X1 U10887 ( .B1(n9695), .B2(n9734), .A(n9663), .ZN(n9664) );
  OAI21_X1 U10888 ( .B1(n9736), .B2(n9700), .A(n9664), .ZN(P1_U3544) );
  NAND2_X1 U10889 ( .A1(n9666), .A2(n9665), .ZN(n9737) );
  MUX2_X1 U10890 ( .A(n9737), .B(P1_REG1_REG_21__SCAN_IN), .S(n9893), .Z(n9667) );
  AOI21_X1 U10891 ( .B1(n9695), .B2(n9739), .A(n9667), .ZN(n9668) );
  OAI21_X1 U10892 ( .B1(n9741), .B2(n9700), .A(n9668), .ZN(P1_U3543) );
  NAND2_X1 U10893 ( .A1(n9670), .A2(n9669), .ZN(n9742) );
  MUX2_X1 U10894 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9742), .S(n9896), .Z(n9671) );
  AOI21_X1 U10895 ( .B1(n9695), .B2(n9744), .A(n9671), .ZN(n9672) );
  OAI21_X1 U10896 ( .B1(n9746), .B2(n9700), .A(n9672), .ZN(P1_U3542) );
  INV_X1 U10897 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9676) );
  AOI211_X1 U10898 ( .C1(n9675), .C2(n9878), .A(n9674), .B(n9673), .ZN(n9747)
         );
  MUX2_X1 U10899 ( .A(n9676), .B(n9747), .S(n9896), .Z(n9677) );
  OAI21_X1 U10900 ( .B1(n9750), .B2(n9686), .A(n9677), .ZN(P1_U3541) );
  AOI22_X1 U10901 ( .A1(n9751), .A2(n9695), .B1(P1_REG1_REG_18__SCAN_IN), .B2(
        n9893), .ZN(n9681) );
  NAND2_X1 U10902 ( .A1(n9679), .A2(n9678), .ZN(n9752) );
  NAND2_X1 U10903 ( .A1(n9752), .A2(n9896), .ZN(n9680) );
  OAI211_X1 U10904 ( .C1(n9755), .C2(n9700), .A(n9681), .B(n9680), .ZN(
        P1_U3540) );
  INV_X1 U10905 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10290) );
  AOI211_X1 U10906 ( .C1(n9684), .C2(n9878), .A(n9683), .B(n9682), .ZN(n9756)
         );
  MUX2_X1 U10907 ( .A(n10290), .B(n9756), .S(n9896), .Z(n9685) );
  OAI21_X1 U10908 ( .B1(n9760), .B2(n9686), .A(n9685), .ZN(P1_U3539) );
  AOI22_X1 U10909 ( .A1(n9761), .A2(n9695), .B1(P1_REG1_REG_16__SCAN_IN), .B2(
        n9893), .ZN(n9690) );
  NAND2_X1 U10910 ( .A1(n9688), .A2(n9687), .ZN(n9762) );
  NAND2_X1 U10911 ( .A1(n9762), .A2(n9896), .ZN(n9689) );
  OAI211_X1 U10912 ( .C1(n9765), .C2(n9700), .A(n9690), .B(n9689), .ZN(
        P1_U3538) );
  AOI211_X1 U10913 ( .C1(n9693), .C2(n9878), .A(n9692), .B(n9691), .ZN(n9768)
         );
  AOI22_X1 U10914 ( .A1(n9766), .A2(n9695), .B1(P1_REG1_REG_15__SCAN_IN), .B2(
        n9893), .ZN(n9694) );
  OAI21_X1 U10915 ( .B1(n9768), .B2(n9893), .A(n9694), .ZN(P1_U3537) );
  AOI22_X1 U10916 ( .A1(n9770), .A2(n9695), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n9893), .ZN(n9699) );
  NAND2_X1 U10917 ( .A1(n9697), .A2(n9696), .ZN(n9771) );
  NAND2_X1 U10918 ( .A1(n9771), .A2(n9896), .ZN(n9698) );
  OAI211_X1 U10919 ( .C1(n9775), .C2(n9700), .A(n9699), .B(n9698), .ZN(
        P1_U3536) );
  INV_X1 U10920 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10155) );
  MUX2_X1 U10921 ( .A(n10155), .B(n9701), .S(n9890), .Z(n9702) );
  OAI21_X1 U10922 ( .B1(n9703), .B2(n9759), .A(n9702), .ZN(P1_U3521) );
  INV_X1 U10923 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9705) );
  MUX2_X1 U10924 ( .A(n9705), .B(n9704), .S(n9890), .Z(n9706) );
  OAI21_X1 U10925 ( .B1(n9707), .B2(n9759), .A(n9706), .ZN(P1_U3520) );
  INV_X1 U10926 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9712) );
  MUX2_X1 U10927 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9714), .S(n9890), .Z(n9715) );
  AOI21_X1 U10928 ( .B1(n9769), .B2(n9716), .A(n9715), .ZN(n9717) );
  OAI21_X1 U10929 ( .B1(n9718), .B2(n9774), .A(n9717), .ZN(P1_U3516) );
  INV_X1 U10930 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9720) );
  MUX2_X1 U10931 ( .A(n9720), .B(n9719), .S(n9890), .Z(n9721) );
  OAI21_X1 U10932 ( .B1(n9722), .B2(n9759), .A(n9721), .ZN(P1_U3515) );
  MUX2_X1 U10933 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9723), .S(n9890), .Z(n9724) );
  AOI21_X1 U10934 ( .B1(n9769), .B2(n9725), .A(n9724), .ZN(n9726) );
  OAI21_X1 U10935 ( .B1(n9727), .B2(n9774), .A(n9726), .ZN(P1_U3514) );
  INV_X1 U10936 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9729) );
  MUX2_X1 U10937 ( .A(n9729), .B(n9728), .S(n9890), .Z(n9730) );
  OAI21_X1 U10938 ( .B1(n9731), .B2(n9759), .A(n9730), .ZN(P1_U3513) );
  MUX2_X1 U10939 ( .A(n9732), .B(P1_REG0_REG_22__SCAN_IN), .S(n9888), .Z(n9733) );
  AOI21_X1 U10940 ( .B1(n9769), .B2(n9734), .A(n9733), .ZN(n9735) );
  OAI21_X1 U10941 ( .B1(n9736), .B2(n9774), .A(n9735), .ZN(P1_U3512) );
  MUX2_X1 U10942 ( .A(n9737), .B(P1_REG0_REG_21__SCAN_IN), .S(n9888), .Z(n9738) );
  AOI21_X1 U10943 ( .B1(n9769), .B2(n9739), .A(n9738), .ZN(n9740) );
  OAI21_X1 U10944 ( .B1(n9741), .B2(n9774), .A(n9740), .ZN(P1_U3511) );
  MUX2_X1 U10945 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9742), .S(n9890), .Z(n9743) );
  AOI21_X1 U10946 ( .B1(n9769), .B2(n9744), .A(n9743), .ZN(n9745) );
  OAI21_X1 U10947 ( .B1(n9746), .B2(n9774), .A(n9745), .ZN(P1_U3510) );
  INV_X1 U10948 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9748) );
  MUX2_X1 U10949 ( .A(n9748), .B(n9747), .S(n9890), .Z(n9749) );
  OAI21_X1 U10950 ( .B1(n9750), .B2(n9759), .A(n9749), .ZN(P1_U3509) );
  AOI22_X1 U10951 ( .A1(n9751), .A2(n9769), .B1(P1_REG0_REG_18__SCAN_IN), .B2(
        n9888), .ZN(n9754) );
  NAND2_X1 U10952 ( .A1(n9752), .A2(n9890), .ZN(n9753) );
  OAI211_X1 U10953 ( .C1(n9755), .C2(n9774), .A(n9754), .B(n9753), .ZN(
        P1_U3507) );
  INV_X1 U10954 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9757) );
  MUX2_X1 U10955 ( .A(n9757), .B(n9756), .S(n9890), .Z(n9758) );
  OAI21_X1 U10956 ( .B1(n9760), .B2(n9759), .A(n9758), .ZN(P1_U3504) );
  AOI22_X1 U10957 ( .A1(n9761), .A2(n9769), .B1(P1_REG0_REG_16__SCAN_IN), .B2(
        n9888), .ZN(n9764) );
  NAND2_X1 U10958 ( .A1(n9762), .A2(n9890), .ZN(n9763) );
  OAI211_X1 U10959 ( .C1(n9765), .C2(n9774), .A(n9764), .B(n9763), .ZN(
        P1_U3501) );
  AOI22_X1 U10960 ( .A1(n9766), .A2(n9769), .B1(P1_REG0_REG_15__SCAN_IN), .B2(
        n9888), .ZN(n9767) );
  OAI21_X1 U10961 ( .B1(n9768), .B2(n9888), .A(n9767), .ZN(P1_U3498) );
  AOI22_X1 U10962 ( .A1(n9770), .A2(n9769), .B1(P1_REG0_REG_14__SCAN_IN), .B2(
        n9888), .ZN(n9773) );
  NAND2_X1 U10963 ( .A1(n9771), .A2(n9890), .ZN(n9772) );
  OAI211_X1 U10964 ( .C1(n9775), .C2(n9774), .A(n9773), .B(n9772), .ZN(
        P1_U3495) );
  MUX2_X1 U10965 ( .A(P1_D_REG_1__SCAN_IN), .B(n9776), .S(n9871), .Z(P1_U3440)
         );
  INV_X1 U10966 ( .A(n9777), .ZN(n9779) );
  NOR4_X1 U10967 ( .A1(n9779), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n6244), .ZN(n9780) );
  AOI21_X1 U10968 ( .B1(n9781), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9780), .ZN(
        n9782) );
  OAI21_X1 U10969 ( .B1(n9783), .B2(n4336), .A(n9782), .ZN(P1_U3324) );
  OAI222_X1 U10970 ( .A1(n4336), .A2(n9786), .B1(n9785), .B2(P1_U3086), .C1(
        n9784), .C2(n9789), .ZN(P1_U3326) );
  OAI222_X1 U10971 ( .A1(n4336), .A2(n9788), .B1(n4337), .B2(P1_U3086), .C1(
        n9787), .C2(n9789), .ZN(P1_U3327) );
  OAI222_X1 U10972 ( .A1(n4336), .A2(n9791), .B1(n9817), .B2(P1_U3086), .C1(
        n9790), .C2(n9789), .ZN(P1_U3328) );
  MUX2_X1 U10973 ( .A(n9792), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI21_X1 U10974 ( .B1(n9794), .B2(n9120), .A(n9793), .ZN(n9799) );
  OAI21_X1 U10975 ( .B1(n9797), .B2(n9796), .A(n9795), .ZN(n9798) );
  XNOR2_X1 U10976 ( .A(n9799), .B(n9798), .ZN(n9810) );
  NOR2_X1 U10977 ( .A1(n9801), .A2(n9800), .ZN(n9808) );
  INV_X1 U10978 ( .A(n9802), .ZN(n9806) );
  OAI22_X1 U10979 ( .A1(n9806), .A2(n9805), .B1(n9804), .B2(n9803), .ZN(n9807)
         );
  AOI211_X1 U10980 ( .C1(n9810), .C2(n9809), .A(n9808), .B(n9807), .ZN(n9812)
         );
  OAI211_X1 U10981 ( .C1(n9814), .C2(n9813), .A(n9812), .B(n9811), .ZN(
        P1_U3236) );
  XNOR2_X1 U10982 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10983 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10984 ( .A(n9815), .ZN(n9818) );
  NAND2_X1 U10985 ( .A1(n9817), .A2(n9816), .ZN(n9820) );
  NAND2_X1 U10986 ( .A1(n9818), .A2(n9820), .ZN(n9821) );
  MUX2_X1 U10987 ( .A(n9821), .B(n9820), .S(n9819), .Z(n9823) );
  NAND2_X1 U10988 ( .A1(n9823), .A2(n9822), .ZN(n9826) );
  AOI22_X1 U10989 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9824), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9825) );
  OAI21_X1 U10990 ( .B1(n9827), .B2(n9826), .A(n9825), .ZN(P1_U3243) );
  OAI21_X1 U10991 ( .B1(n9830), .B2(n9829), .A(n9828), .ZN(n9837) );
  AOI21_X1 U10992 ( .B1(n9833), .B2(n9832), .A(n9831), .ZN(n9835) );
  OAI22_X1 U10993 ( .A1(n9835), .A2(n9849), .B1(n9834), .B2(n9847), .ZN(n9836)
         );
  AOI21_X1 U10994 ( .B1(n9853), .B2(n9837), .A(n9836), .ZN(n9839) );
  OAI211_X1 U10995 ( .C1(n9857), .C2(n9840), .A(n9839), .B(n9838), .ZN(
        P1_U3255) );
  OAI21_X1 U10996 ( .B1(n9843), .B2(n9842), .A(n9841), .ZN(n9852) );
  AOI21_X1 U10997 ( .B1(n9846), .B2(n9845), .A(n9844), .ZN(n9850) );
  OAI22_X1 U10998 ( .A1(n9850), .A2(n9849), .B1(n9848), .B2(n9847), .ZN(n9851)
         );
  AOI21_X1 U10999 ( .B1(n9853), .B2(n9852), .A(n9851), .ZN(n9855) );
  OAI211_X1 U11000 ( .C1(n9857), .C2(n9856), .A(n9855), .B(n9854), .ZN(
        P1_U3260) );
  NAND2_X1 U11001 ( .A1(n9859), .A2(n9858), .ZN(n9863) );
  AOI22_X1 U11002 ( .A1(n9617), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9861), .B2(
        n9860), .ZN(n9862) );
  OAI211_X1 U11003 ( .C1(n9865), .C2(n9864), .A(n9863), .B(n9862), .ZN(n9866)
         );
  AOI21_X1 U11004 ( .B1(n9868), .B2(n9867), .A(n9866), .ZN(n9869) );
  OAI21_X1 U11005 ( .B1(n9617), .B2(n9870), .A(n9869), .ZN(P1_U3290) );
  AND2_X1 U11006 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9872), .ZN(P1_U3294) );
  INV_X1 U11007 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10262) );
  NOR2_X1 U11008 ( .A1(n9871), .A2(n10262), .ZN(P1_U3295) );
  AND2_X1 U11009 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9872), .ZN(P1_U3296) );
  AND2_X1 U11010 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9872), .ZN(P1_U3297) );
  AND2_X1 U11011 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9872), .ZN(P1_U3298) );
  AND2_X1 U11012 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9872), .ZN(P1_U3299) );
  AND2_X1 U11013 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9872), .ZN(P1_U3300) );
  INV_X1 U11014 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10245) );
  NOR2_X1 U11015 ( .A1(n9871), .A2(n10245), .ZN(P1_U3301) );
  AND2_X1 U11016 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9872), .ZN(P1_U3302) );
  AND2_X1 U11017 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9872), .ZN(P1_U3303) );
  AND2_X1 U11018 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9872), .ZN(P1_U3304) );
  AND2_X1 U11019 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9872), .ZN(P1_U3305) );
  AND2_X1 U11020 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9872), .ZN(P1_U3306) );
  AND2_X1 U11021 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9872), .ZN(P1_U3307) );
  AND2_X1 U11022 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9872), .ZN(P1_U3308) );
  AND2_X1 U11023 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9872), .ZN(P1_U3309) );
  AND2_X1 U11024 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9872), .ZN(P1_U3310) );
  AND2_X1 U11025 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9872), .ZN(P1_U3311) );
  AND2_X1 U11026 ( .A1(n9872), .A2(P1_D_REG_13__SCAN_IN), .ZN(P1_U3312) );
  AND2_X1 U11027 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9872), .ZN(P1_U3313) );
  AND2_X1 U11028 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9872), .ZN(P1_U3314) );
  AND2_X1 U11029 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9872), .ZN(P1_U3315) );
  AND2_X1 U11030 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9872), .ZN(P1_U3316) );
  AND2_X1 U11031 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9872), .ZN(P1_U3317) );
  AND2_X1 U11032 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9872), .ZN(P1_U3318) );
  AND2_X1 U11033 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9872), .ZN(P1_U3319) );
  AND2_X1 U11034 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9872), .ZN(P1_U3320) );
  AND2_X1 U11035 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9872), .ZN(P1_U3321) );
  AND2_X1 U11036 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9872), .ZN(P1_U3322) );
  AND2_X1 U11037 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9872), .ZN(P1_U3323) );
  OAI211_X1 U11038 ( .C1(n9875), .C2(n9881), .A(n9874), .B(n9873), .ZN(n9876)
         );
  AOI21_X1 U11039 ( .B1(n9878), .B2(n9877), .A(n9876), .ZN(n9892) );
  INV_X1 U11040 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9879) );
  AOI22_X1 U11041 ( .A1(n9890), .A2(n9892), .B1(n9879), .B2(n9888), .ZN(
        P1_U3471) );
  OAI21_X1 U11042 ( .B1(n9882), .B2(n9881), .A(n9880), .ZN(n9883) );
  AOI21_X1 U11043 ( .B1(n9885), .B2(n9884), .A(n9883), .ZN(n9886) );
  AND2_X1 U11044 ( .A1(n9887), .A2(n9886), .ZN(n9895) );
  INV_X1 U11045 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9889) );
  AOI22_X1 U11046 ( .A1(n9890), .A2(n9895), .B1(n9889), .B2(n9888), .ZN(
        P1_U3477) );
  AOI22_X1 U11047 ( .A1(n9896), .A2(n9892), .B1(n9891), .B2(n9893), .ZN(
        P1_U3528) );
  AOI22_X1 U11048 ( .A1(n9896), .A2(n9895), .B1(n9894), .B2(n9893), .ZN(
        P1_U3530) );
  OAI21_X1 U11049 ( .B1(n9899), .B2(n9898), .A(n9897), .ZN(n9901) );
  NOR2_X1 U11050 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10022), .ZN(n9900) );
  AOI21_X1 U11051 ( .B1(n10009), .B2(n9901), .A(n9900), .ZN(n9910) );
  NAND2_X1 U11052 ( .A1(n9962), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n9909) );
  NAND2_X1 U11053 ( .A1(n10003), .A2(n4602), .ZN(n9908) );
  OAI21_X1 U11054 ( .B1(n9904), .B2(n9903), .A(n9902), .ZN(n9905) );
  NAND2_X1 U11055 ( .A1(n9906), .A2(n9905), .ZN(n9907) );
  AND4_X1 U11056 ( .A1(n9910), .A2(n9909), .A3(n9908), .A4(n9907), .ZN(n9915)
         );
  XOR2_X1 U11057 ( .A(n9912), .B(n9911), .Z(n9913) );
  NAND2_X1 U11058 ( .A1(n9913), .A2(n9949), .ZN(n9914) );
  NAND2_X1 U11059 ( .A1(n9915), .A2(n9914), .ZN(P2_U3184) );
  INV_X1 U11060 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n9935) );
  AOI21_X1 U11061 ( .B1(n9918), .B2(n9917), .A(n9916), .ZN(n9927) );
  AOI21_X1 U11062 ( .B1(n9920), .B2(n5283), .A(n9919), .ZN(n9922) );
  OAI21_X1 U11063 ( .B1(n9980), .B2(n9922), .A(n9921), .ZN(n9923) );
  INV_X1 U11064 ( .A(n9923), .ZN(n9926) );
  NAND2_X1 U11065 ( .A1(n10003), .A2(n9924), .ZN(n9925) );
  OAI211_X1 U11066 ( .C1(n9927), .C2(n10005), .A(n9926), .B(n9925), .ZN(n9928)
         );
  INV_X1 U11067 ( .A(n9928), .ZN(n9934) );
  AOI21_X1 U11068 ( .B1(n9931), .B2(n9930), .A(n9929), .ZN(n9932) );
  OR2_X1 U11069 ( .A1(n9932), .A2(n10013), .ZN(n9933) );
  OAI211_X1 U11070 ( .C1(n9935), .C2(n10017), .A(n9934), .B(n9933), .ZN(
        P2_U3185) );
  INV_X1 U11071 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9953) );
  AOI21_X1 U11072 ( .B1(n10087), .B2(n9937), .A(n9936), .ZN(n9945) );
  AOI21_X1 U11073 ( .B1(n10003), .B2(n9939), .A(n9938), .ZN(n9944) );
  AOI21_X1 U11074 ( .B1(n7395), .B2(n9941), .A(n9940), .ZN(n9942) );
  OR2_X1 U11075 ( .A1(n9942), .A2(n9980), .ZN(n9943) );
  OAI211_X1 U11076 ( .C1(n9945), .C2(n10005), .A(n9944), .B(n9943), .ZN(n9946)
         );
  INV_X1 U11077 ( .A(n9946), .ZN(n9952) );
  XOR2_X1 U11078 ( .A(n9948), .B(n9947), .Z(n9950) );
  NAND2_X1 U11079 ( .A1(n9950), .A2(n9949), .ZN(n9951) );
  OAI211_X1 U11080 ( .C1(n9953), .C2(n10017), .A(n9952), .B(n9951), .ZN(
        P2_U3187) );
  INV_X1 U11081 ( .A(n9954), .ZN(n9955) );
  AOI21_X1 U11082 ( .B1(n9957), .B2(n9956), .A(n9955), .ZN(n9960) );
  OAI22_X1 U11083 ( .A1(n9960), .A2(n9980), .B1(n9959), .B2(n9958), .ZN(n9961)
         );
  AOI21_X1 U11084 ( .B1(n9962), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n9961), .ZN(
        n9975) );
  AOI21_X1 U11085 ( .B1(n9965), .B2(n9964), .A(n9963), .ZN(n9966) );
  OR2_X1 U11086 ( .A1(n9966), .A2(n10013), .ZN(n9973) );
  INV_X1 U11087 ( .A(n9967), .ZN(n9968) );
  AOI21_X1 U11088 ( .B1(n9970), .B2(n9969), .A(n9968), .ZN(n9971) );
  OR2_X1 U11089 ( .A1(n9971), .A2(n10005), .ZN(n9972) );
  NAND4_X1 U11090 ( .A1(n9975), .A2(n9974), .A3(n9973), .A4(n9972), .ZN(
        P2_U3188) );
  AOI21_X1 U11091 ( .B1(n7317), .B2(n9977), .A(n9976), .ZN(n9986) );
  AOI21_X1 U11092 ( .B1(n7376), .B2(n9979), .A(n9978), .ZN(n9981) );
  OR2_X1 U11093 ( .A1(n9981), .A2(n9980), .ZN(n9985) );
  AOI21_X1 U11094 ( .B1(n10003), .B2(n9983), .A(n9982), .ZN(n9984) );
  OAI211_X1 U11095 ( .C1(n9986), .C2(n10005), .A(n9985), .B(n9984), .ZN(n9987)
         );
  INV_X1 U11096 ( .A(n9987), .ZN(n9993) );
  AOI21_X1 U11097 ( .B1(n9990), .B2(n9989), .A(n9988), .ZN(n9991) );
  OR2_X1 U11098 ( .A1(n9991), .A2(n10013), .ZN(n9992) );
  OAI211_X1 U11099 ( .C1(n9994), .C2(n10017), .A(n9993), .B(n9992), .ZN(
        P2_U3189) );
  OAI21_X1 U11100 ( .B1(n4885), .B2(n4884), .A(n9996), .ZN(n10008) );
  INV_X1 U11101 ( .A(n9997), .ZN(n9998) );
  AOI21_X1 U11102 ( .B1(n10000), .B2(n9999), .A(n9998), .ZN(n10006) );
  AOI21_X1 U11103 ( .B1(n10003), .B2(n10002), .A(n10001), .ZN(n10004) );
  OAI21_X1 U11104 ( .B1(n10006), .B2(n10005), .A(n10004), .ZN(n10007) );
  AOI21_X1 U11105 ( .B1(n10009), .B2(n10008), .A(n10007), .ZN(n10016) );
  AOI21_X1 U11106 ( .B1(n10012), .B2(n10011), .A(n10010), .ZN(n10014) );
  OR2_X1 U11107 ( .A1(n10014), .A2(n10013), .ZN(n10015) );
  OAI211_X1 U11108 ( .C1(n10018), .C2(n10017), .A(n10016), .B(n10015), .ZN(
        P2_U3190) );
  OAI21_X1 U11109 ( .B1(n10020), .B2(n4724), .A(n10019), .ZN(n10038) );
  OAI22_X1 U11110 ( .A1(n10035), .A2(n10023), .B1(n10022), .B2(n10021), .ZN(
        n10031) );
  XNOR2_X1 U11111 ( .A(n10024), .B(n4724), .ZN(n10025) );
  OAI222_X1 U11112 ( .A1(n10030), .A2(n10029), .B1(n10028), .B2(n10027), .C1(
        n10026), .C2(n10025), .ZN(n10036) );
  AOI211_X1 U11113 ( .C1(n10032), .C2(n10038), .A(n10031), .B(n10036), .ZN(
        n10033) );
  AOI22_X1 U11114 ( .A1(n10034), .A2(n5267), .B1(n10033), .B2(n8926), .ZN(
        P2_U3231) );
  NOR2_X1 U11115 ( .A1(n10035), .A2(n10052), .ZN(n10037) );
  AOI211_X1 U11116 ( .C1(n10075), .C2(n10038), .A(n10037), .B(n10036), .ZN(
        n10084) );
  AOI22_X1 U11117 ( .A1(n10082), .A2(n5266), .B1(n10084), .B2(n10081), .ZN(
        P2_U3396) );
  OAI21_X1 U11118 ( .B1(n5315), .B2(n10052), .A(n10039), .ZN(n10040) );
  AOI21_X1 U11119 ( .B1(n10041), .B2(n10075), .A(n10040), .ZN(n10086) );
  AOI22_X1 U11120 ( .A1(n10082), .A2(n5300), .B1(n10086), .B2(n10081), .ZN(
        P2_U3402) );
  INV_X1 U11121 ( .A(n10042), .ZN(n10046) );
  OAI22_X1 U11122 ( .A1(n10044), .A2(n10068), .B1(n10043), .B2(n10052), .ZN(
        n10045) );
  NOR2_X1 U11123 ( .A1(n10046), .A2(n10045), .ZN(n10088) );
  AOI22_X1 U11124 ( .A1(n10082), .A2(n5318), .B1(n10088), .B2(n10081), .ZN(
        P2_U3405) );
  OAI22_X1 U11125 ( .A1(n10048), .A2(n10068), .B1(n10047), .B2(n10052), .ZN(
        n10049) );
  NOR2_X1 U11126 ( .A1(n10050), .A2(n10049), .ZN(n10089) );
  AOI22_X1 U11127 ( .A1(n10082), .A2(n5333), .B1(n10089), .B2(n10081), .ZN(
        P2_U3408) );
  INV_X1 U11128 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10058) );
  NOR2_X1 U11129 ( .A1(n10054), .A2(n10051), .ZN(n10056) );
  OAI22_X1 U11130 ( .A1(n10054), .A2(n10063), .B1(n10053), .B2(n10052), .ZN(
        n10055) );
  NOR3_X1 U11131 ( .A1(n10057), .A2(n10056), .A3(n10055), .ZN(n10090) );
  AOI22_X1 U11132 ( .A1(n10082), .A2(n10058), .B1(n10090), .B2(n10081), .ZN(
        P2_U3411) );
  NOR2_X1 U11133 ( .A1(n10059), .A2(n10063), .ZN(n10061) );
  AOI211_X1 U11134 ( .C1(n10080), .C2(n10062), .A(n10061), .B(n10060), .ZN(
        n10091) );
  AOI22_X1 U11135 ( .A1(n10082), .A2(n5388), .B1(n10091), .B2(n10081), .ZN(
        P2_U3417) );
  NOR2_X1 U11136 ( .A1(n10064), .A2(n10063), .ZN(n10066) );
  AOI211_X1 U11137 ( .C1(n10080), .C2(n10067), .A(n10066), .B(n10065), .ZN(
        n10092) );
  AOI22_X1 U11138 ( .A1(n10082), .A2(n5411), .B1(n10092), .B2(n10081), .ZN(
        P2_U3420) );
  INV_X1 U11139 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10073) );
  NOR2_X1 U11140 ( .A1(n10069), .A2(n10068), .ZN(n10071) );
  AOI211_X1 U11141 ( .C1(n10080), .C2(n10072), .A(n10071), .B(n10070), .ZN(
        n10093) );
  AOI22_X1 U11142 ( .A1(n10082), .A2(n10073), .B1(n10093), .B2(n10081), .ZN(
        P2_U3423) );
  AND3_X1 U11143 ( .A1(n10076), .A2(n10075), .A3(n10074), .ZN(n10078) );
  AOI211_X1 U11144 ( .C1(n10080), .C2(n10079), .A(n10078), .B(n10077), .ZN(
        n10095) );
  AOI22_X1 U11145 ( .A1(n10082), .A2(n5445), .B1(n10095), .B2(n10081), .ZN(
        P2_U3426) );
  AOI22_X1 U11146 ( .A1(n10096), .A2(n10084), .B1(n10083), .B2(n10094), .ZN(
        P2_U3461) );
  INV_X1 U11147 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10085) );
  AOI22_X1 U11148 ( .A1(n10096), .A2(n10086), .B1(n10085), .B2(n10094), .ZN(
        P2_U3463) );
  AOI22_X1 U11149 ( .A1(n10096), .A2(n10088), .B1(n10087), .B2(n10094), .ZN(
        P2_U3464) );
  AOI22_X1 U11150 ( .A1(n10096), .A2(n10089), .B1(n7311), .B2(n10094), .ZN(
        P2_U3465) );
  AOI22_X1 U11151 ( .A1(n10096), .A2(n10090), .B1(n7317), .B2(n10094), .ZN(
        P2_U3466) );
  AOI22_X1 U11152 ( .A1(n10096), .A2(n10091), .B1(n10121), .B2(n10094), .ZN(
        P2_U3468) );
  AOI22_X1 U11153 ( .A1(n10096), .A2(n10092), .B1(n7423), .B2(n10094), .ZN(
        P2_U3469) );
  AOI22_X1 U11154 ( .A1(n10096), .A2(n10093), .B1(n5425), .B2(n10094), .ZN(
        P2_U3470) );
  AOI22_X1 U11155 ( .A1(n10096), .A2(n10095), .B1(n5442), .B2(n10094), .ZN(
        P2_U3471) );
  NOR2_X1 U11156 ( .A1(n10098), .A2(n10097), .ZN(n10099) );
  XOR2_X1 U11157 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10099), .Z(ADD_1068_U5) );
  XOR2_X1 U11158 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11159 ( .A1(n10101), .A2(n10100), .ZN(n10102) );
  XOR2_X1 U11160 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n10102), .Z(ADD_1068_U55)
         );
  XNOR2_X1 U11161 ( .A(n10104), .B(n10103), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11162 ( .A(n10106), .B(n10105), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11163 ( .A(n10108), .B(n10107), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11164 ( .A(n10110), .B(n10109), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11165 ( .A(n10112), .B(n10111), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11166 ( .A(n10114), .B(n10113), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11167 ( .A(n10116), .B(n10115), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11168 ( .A(n10118), .B(n10117), .ZN(ADD_1068_U63) );
  NAND2_X1 U11169 ( .A1(n10119), .A2(P2_D_REG_4__SCAN_IN), .ZN(n10307) );
  AOI22_X1 U11170 ( .A1(n10122), .A2(keyinput67), .B1(n10121), .B2(keyinput96), 
        .ZN(n10120) );
  OAI221_X1 U11171 ( .B1(n10122), .B2(keyinput67), .C1(n10121), .C2(keyinput96), .A(n10120), .ZN(n10131) );
  INV_X1 U11172 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n10124) );
  AOI22_X1 U11173 ( .A1(n10124), .A2(keyinput73), .B1(keyinput107), .B2(n10271), .ZN(n10123) );
  OAI221_X1 U11174 ( .B1(n10124), .B2(keyinput73), .C1(n10271), .C2(
        keyinput107), .A(n10123), .ZN(n10130) );
  AOI22_X1 U11175 ( .A1(n10022), .A2(keyinput114), .B1(n10291), .B2(
        keyinput102), .ZN(n10125) );
  OAI221_X1 U11176 ( .B1(n10022), .B2(keyinput114), .C1(n10291), .C2(
        keyinput102), .A(n10125), .ZN(n10129) );
  INV_X1 U11177 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10127) );
  AOI22_X1 U11178 ( .A1(n10127), .A2(keyinput117), .B1(keyinput125), .B2(n9477), .ZN(n10126) );
  OAI221_X1 U11179 ( .B1(n10127), .B2(keyinput117), .C1(n9477), .C2(
        keyinput125), .A(n10126), .ZN(n10128) );
  NOR4_X1 U11180 ( .A1(n10131), .A2(n10130), .A3(n10129), .A4(n10128), .ZN(
        n10170) );
  AOI22_X1 U11181 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(keyinput108), .B1(
        P2_D_REG_21__SCAN_IN), .B2(keyinput88), .ZN(n10132) );
  OAI221_X1 U11182 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(keyinput108), .C1(
        P2_D_REG_21__SCAN_IN), .C2(keyinput88), .A(n10132), .ZN(n10135) );
  AOI22_X1 U11183 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(keyinput87), .B1(
        P2_REG2_REG_5__SCAN_IN), .B2(keyinput71), .ZN(n10133) );
  OAI221_X1 U11184 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(keyinput87), .C1(
        P2_REG2_REG_5__SCAN_IN), .C2(keyinput71), .A(n10133), .ZN(n10134) );
  NOR2_X1 U11185 ( .A1(n10135), .A2(n10134), .ZN(n10143) );
  INV_X1 U11186 ( .A(keyinput68), .ZN(n10136) );
  XNOR2_X1 U11187 ( .A(n10278), .B(n10136), .ZN(n10142) );
  XNOR2_X1 U11188 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput115), .ZN(n10141) );
  AOI22_X1 U11189 ( .A1(P2_D_REG_10__SCAN_IN), .A2(keyinput64), .B1(n10138), 
        .B2(keyinput103), .ZN(n10137) );
  OAI221_X1 U11190 ( .B1(P2_D_REG_10__SCAN_IN), .B2(keyinput64), .C1(n10138), 
        .C2(keyinput103), .A(n10137), .ZN(n10139) );
  INV_X1 U11191 ( .A(n10139), .ZN(n10140) );
  AND4_X1 U11192 ( .A1(n10143), .A2(n10142), .A3(n10141), .A4(n10140), .ZN(
        n10169) );
  AOI22_X1 U11193 ( .A1(n10145), .A2(keyinput124), .B1(n10255), .B2(keyinput90), .ZN(n10144) );
  OAI221_X1 U11194 ( .B1(n10145), .B2(keyinput124), .C1(n10255), .C2(
        keyinput90), .A(n10144), .ZN(n10153) );
  XNOR2_X1 U11195 ( .A(n10273), .B(keyinput123), .ZN(n10152) );
  INV_X1 U11196 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n10279) );
  XNOR2_X1 U11197 ( .A(keyinput85), .B(n10279), .ZN(n10151) );
  XNOR2_X1 U11198 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput76), .ZN(n10149) );
  XNOR2_X1 U11199 ( .A(P1_REG0_REG_24__SCAN_IN), .B(keyinput75), .ZN(n10148)
         );
  XNOR2_X1 U11200 ( .A(SI_29_), .B(keyinput78), .ZN(n10147) );
  XNOR2_X1 U11201 ( .A(P1_REG3_REG_4__SCAN_IN), .B(keyinput95), .ZN(n10146) );
  NAND4_X1 U11202 ( .A1(n10149), .A2(n10148), .A3(n10147), .A4(n10146), .ZN(
        n10150) );
  NOR4_X1 U11203 ( .A1(n10153), .A2(n10152), .A3(n10151), .A4(n10150), .ZN(
        n10168) );
  AOI22_X1 U11204 ( .A1(n10288), .A2(keyinput94), .B1(n10155), .B2(keyinput74), 
        .ZN(n10154) );
  OAI221_X1 U11205 ( .B1(n10288), .B2(keyinput94), .C1(n10155), .C2(keyinput74), .A(n10154), .ZN(n10166) );
  INV_X1 U11206 ( .A(SI_16_), .ZN(n10272) );
  AOI22_X1 U11207 ( .A1(n10272), .A2(keyinput120), .B1(keyinput86), .B2(n5245), 
        .ZN(n10156) );
  OAI221_X1 U11208 ( .B1(n10272), .B2(keyinput120), .C1(n5245), .C2(keyinput86), .A(n10156), .ZN(n10165) );
  AOI22_X1 U11209 ( .A1(n10159), .A2(keyinput110), .B1(n10158), .B2(keyinput80), .ZN(n10157) );
  OAI221_X1 U11210 ( .B1(n10159), .B2(keyinput110), .C1(n10158), .C2(
        keyinput80), .A(n10157), .ZN(n10164) );
  AOI22_X1 U11211 ( .A1(n10162), .A2(keyinput97), .B1(keyinput82), .B2(n10161), 
        .ZN(n10160) );
  OAI221_X1 U11212 ( .B1(n10162), .B2(keyinput97), .C1(n10161), .C2(keyinput82), .A(n10160), .ZN(n10163) );
  NOR4_X1 U11213 ( .A1(n10166), .A2(n10165), .A3(n10164), .A4(n10163), .ZN(
        n10167) );
  AND4_X1 U11214 ( .A1(n10170), .A2(n10169), .A3(n10168), .A4(n10167), .ZN(
        n10305) );
  OAI22_X1 U11215 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(keyinput104), .B1(
        keyinput83), .B2(P1_REG1_REG_3__SCAN_IN), .ZN(n10171) );
  AOI221_X1 U11216 ( .B1(P2_IR_REG_19__SCAN_IN), .B2(keyinput104), .C1(
        P1_REG1_REG_3__SCAN_IN), .C2(keyinput83), .A(n10171), .ZN(n10178) );
  OAI22_X1 U11217 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(keyinput84), .B1(
        keyinput101), .B2(P2_ADDR_REG_11__SCAN_IN), .ZN(n10172) );
  AOI221_X1 U11218 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(keyinput84), .C1(
        P2_ADDR_REG_11__SCAN_IN), .C2(keyinput101), .A(n10172), .ZN(n10177) );
  OAI22_X1 U11219 ( .A1(P2_D_REG_4__SCAN_IN), .A2(keyinput65), .B1(
        P2_REG1_REG_31__SCAN_IN), .B2(keyinput93), .ZN(n10173) );
  AOI221_X1 U11220 ( .B1(P2_D_REG_4__SCAN_IN), .B2(keyinput65), .C1(keyinput93), .C2(P2_REG1_REG_31__SCAN_IN), .A(n10173), .ZN(n10176) );
  OAI22_X1 U11221 ( .A1(P2_REG0_REG_28__SCAN_IN), .A2(keyinput122), .B1(
        P1_REG1_REG_29__SCAN_IN), .B2(keyinput127), .ZN(n10174) );
  AOI221_X1 U11222 ( .B1(P2_REG0_REG_28__SCAN_IN), .B2(keyinput122), .C1(
        keyinput127), .C2(P1_REG1_REG_29__SCAN_IN), .A(n10174), .ZN(n10175) );
  NAND4_X1 U11223 ( .A1(n10178), .A2(n10177), .A3(n10176), .A4(n10175), .ZN(
        n10206) );
  OAI22_X1 U11224 ( .A1(P2_D_REG_14__SCAN_IN), .A2(keyinput118), .B1(
        keyinput105), .B2(P2_D_REG_5__SCAN_IN), .ZN(n10179) );
  AOI221_X1 U11225 ( .B1(P2_D_REG_14__SCAN_IN), .B2(keyinput118), .C1(
        P2_D_REG_5__SCAN_IN), .C2(keyinput105), .A(n10179), .ZN(n10186) );
  OAI22_X1 U11226 ( .A1(SI_7_), .A2(keyinput92), .B1(P1_REG1_REG_17__SCAN_IN), 
        .B2(keyinput126), .ZN(n10180) );
  AOI221_X1 U11227 ( .B1(SI_7_), .B2(keyinput92), .C1(keyinput126), .C2(
        P1_REG1_REG_17__SCAN_IN), .A(n10180), .ZN(n10185) );
  OAI22_X1 U11228 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(keyinput116), .B1(
        P1_REG3_REG_14__SCAN_IN), .B2(keyinput69), .ZN(n10181) );
  AOI221_X1 U11229 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(keyinput116), .C1(
        keyinput69), .C2(P1_REG3_REG_14__SCAN_IN), .A(n10181), .ZN(n10184) );
  OAI22_X1 U11230 ( .A1(P1_D_REG_24__SCAN_IN), .A2(keyinput109), .B1(
        P2_ADDR_REG_14__SCAN_IN), .B2(keyinput106), .ZN(n10182) );
  AOI221_X1 U11231 ( .B1(P1_D_REG_24__SCAN_IN), .B2(keyinput109), .C1(
        keyinput106), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n10182), .ZN(n10183) );
  NAND4_X1 U11232 ( .A1(n10186), .A2(n10185), .A3(n10184), .A4(n10183), .ZN(
        n10205) );
  OAI22_X1 U11233 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(keyinput91), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(keyinput70), .ZN(n10187) );
  AOI221_X1 U11234 ( .B1(P2_IR_REG_30__SCAN_IN), .B2(keyinput91), .C1(
        keyinput70), .C2(P1_REG3_REG_0__SCAN_IN), .A(n10187), .ZN(n10194) );
  OAI22_X1 U11235 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(keyinput100), .B1(
        keyinput81), .B2(P1_D_REG_30__SCAN_IN), .ZN(n10188) );
  AOI221_X1 U11236 ( .B1(P1_DATAO_REG_15__SCAN_IN), .B2(keyinput100), .C1(
        P1_D_REG_30__SCAN_IN), .C2(keyinput81), .A(n10188), .ZN(n10193) );
  OAI22_X1 U11237 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(keyinput119), .B1(
        keyinput99), .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n10189) );
  AOI221_X1 U11238 ( .B1(P2_DATAO_REG_26__SCAN_IN), .B2(keyinput119), .C1(
        P1_DATAO_REG_18__SCAN_IN), .C2(keyinput99), .A(n10189), .ZN(n10192) );
  OAI22_X1 U11239 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput77), .B1(
        keyinput112), .B2(P2_REG2_REG_7__SCAN_IN), .ZN(n10190) );
  AOI221_X1 U11240 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput77), .C1(
        P2_REG2_REG_7__SCAN_IN), .C2(keyinput112), .A(n10190), .ZN(n10191) );
  NAND4_X1 U11241 ( .A1(n10194), .A2(n10193), .A3(n10192), .A4(n10191), .ZN(
        n10204) );
  OAI22_X1 U11242 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput72), .B1(
        keyinput98), .B2(P1_D_REG_13__SCAN_IN), .ZN(n10195) );
  AOI221_X1 U11243 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput72), .C1(
        P1_D_REG_13__SCAN_IN), .C2(keyinput98), .A(n10195), .ZN(n10202) );
  OAI22_X1 U11244 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(keyinput79), .B1(
        keyinput66), .B2(P1_REG2_REG_3__SCAN_IN), .ZN(n10196) );
  AOI221_X1 U11245 ( .B1(P2_IR_REG_28__SCAN_IN), .B2(keyinput79), .C1(
        P1_REG2_REG_3__SCAN_IN), .C2(keyinput66), .A(n10196), .ZN(n10201) );
  OAI22_X1 U11246 ( .A1(P2_D_REG_12__SCAN_IN), .A2(keyinput113), .B1(
        P1_REG0_REG_22__SCAN_IN), .B2(keyinput121), .ZN(n10197) );
  AOI221_X1 U11247 ( .B1(P2_D_REG_12__SCAN_IN), .B2(keyinput113), .C1(
        keyinput121), .C2(P1_REG0_REG_22__SCAN_IN), .A(n10197), .ZN(n10200) );
  OAI22_X1 U11248 ( .A1(SI_6_), .A2(keyinput89), .B1(P1_REG1_REG_15__SCAN_IN), 
        .B2(keyinput111), .ZN(n10198) );
  AOI221_X1 U11249 ( .B1(SI_6_), .B2(keyinput89), .C1(keyinput111), .C2(
        P1_REG1_REG_15__SCAN_IN), .A(n10198), .ZN(n10199) );
  NAND4_X1 U11250 ( .A1(n10202), .A2(n10201), .A3(n10200), .A4(n10199), .ZN(
        n10203) );
  NOR4_X1 U11251 ( .A1(n10206), .A2(n10205), .A3(n10204), .A4(n10203), .ZN(
        n10304) );
  AOI22_X1 U11252 ( .A1(P2_D_REG_10__SCAN_IN), .A2(keyinput0), .B1(
        P2_D_REG_14__SCAN_IN), .B2(keyinput54), .ZN(n10207) );
  OAI221_X1 U11253 ( .B1(P2_D_REG_10__SCAN_IN), .B2(keyinput0), .C1(
        P2_D_REG_14__SCAN_IN), .C2(keyinput54), .A(n10207), .ZN(n10214) );
  AOI22_X1 U11254 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(keyinput6), .B1(
        P2_REG3_REG_20__SCAN_IN), .B2(keyinput13), .ZN(n10208) );
  OAI221_X1 U11255 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(keyinput6), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput13), .A(n10208), .ZN(n10213) );
  AOI22_X1 U11256 ( .A1(P2_REG1_REG_31__SCAN_IN), .A2(keyinput29), .B1(
        P1_REG2_REG_22__SCAN_IN), .B2(keyinput61), .ZN(n10209) );
  OAI221_X1 U11257 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(keyinput29), .C1(
        P1_REG2_REG_22__SCAN_IN), .C2(keyinput61), .A(n10209), .ZN(n10212) );
  AOI22_X1 U11258 ( .A1(P2_REG2_REG_7__SCAN_IN), .A2(keyinput48), .B1(
        P2_REG0_REG_22__SCAN_IN), .B2(keyinput16), .ZN(n10210) );
  OAI221_X1 U11259 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(keyinput48), .C1(
        P2_REG0_REG_22__SCAN_IN), .C2(keyinput16), .A(n10210), .ZN(n10211) );
  NOR4_X1 U11260 ( .A1(n10214), .A2(n10213), .A3(n10212), .A4(n10211), .ZN(
        n10242) );
  AOI22_X1 U11261 ( .A1(P1_REG0_REG_31__SCAN_IN), .A2(keyinput10), .B1(
        P2_REG0_REG_28__SCAN_IN), .B2(keyinput58), .ZN(n10215) );
  OAI221_X1 U11262 ( .B1(P1_REG0_REG_31__SCAN_IN), .B2(keyinput10), .C1(
        P2_REG0_REG_28__SCAN_IN), .C2(keyinput58), .A(n10215), .ZN(n10222) );
  AOI22_X1 U11263 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(keyinput52), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(keyinput18), .ZN(n10216) );
  OAI221_X1 U11264 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(keyinput52), .C1(
        P1_DATAO_REG_14__SCAN_IN), .C2(keyinput18), .A(n10216), .ZN(n10221) );
  AOI22_X1 U11265 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(keyinput44), .B1(
        P1_REG3_REG_27__SCAN_IN), .B2(keyinput60), .ZN(n10217) );
  OAI221_X1 U11266 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(keyinput44), .C1(
        P1_REG3_REG_27__SCAN_IN), .C2(keyinput60), .A(n10217), .ZN(n10220) );
  AOI22_X1 U11267 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(keyinput3), .B1(
        P1_REG3_REG_14__SCAN_IN), .B2(keyinput5), .ZN(n10218) );
  OAI221_X1 U11268 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(keyinput3), .C1(
        P1_REG3_REG_14__SCAN_IN), .C2(keyinput5), .A(n10218), .ZN(n10219) );
  NOR4_X1 U11269 ( .A1(n10222), .A2(n10221), .A3(n10220), .A4(n10219), .ZN(
        n10241) );
  AOI22_X1 U11270 ( .A1(P1_REG0_REG_26__SCAN_IN), .A2(keyinput46), .B1(
        P1_IR_REG_28__SCAN_IN), .B2(keyinput51), .ZN(n10223) );
  OAI221_X1 U11271 ( .B1(P1_REG0_REG_26__SCAN_IN), .B2(keyinput46), .C1(
        P1_IR_REG_28__SCAN_IN), .C2(keyinput51), .A(n10223), .ZN(n10230) );
  AOI22_X1 U11272 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput8), .B1(
        P2_D_REG_12__SCAN_IN), .B2(keyinput49), .ZN(n10224) );
  OAI221_X1 U11273 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput8), .C1(
        P2_D_REG_12__SCAN_IN), .C2(keyinput49), .A(n10224), .ZN(n10229) );
  AOI22_X1 U11274 ( .A1(P2_REG0_REG_1__SCAN_IN), .A2(keyinput22), .B1(
        P2_IR_REG_30__SCAN_IN), .B2(keyinput27), .ZN(n10225) );
  OAI221_X1 U11275 ( .B1(P2_REG0_REG_1__SCAN_IN), .B2(keyinput22), .C1(
        P2_IR_REG_30__SCAN_IN), .C2(keyinput27), .A(n10225), .ZN(n10228) );
  AOI22_X1 U11276 ( .A1(P1_REG0_REG_22__SCAN_IN), .A2(keyinput57), .B1(SI_6_), 
        .B2(keyinput25), .ZN(n10226) );
  OAI221_X1 U11277 ( .B1(P1_REG0_REG_22__SCAN_IN), .B2(keyinput57), .C1(SI_6_), 
        .C2(keyinput25), .A(n10226), .ZN(n10227) );
  NOR4_X1 U11278 ( .A1(n10230), .A2(n10229), .A3(n10228), .A4(n10227), .ZN(
        n10240) );
  AOI22_X1 U11279 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(keyinput32), .B1(
        P2_REG1_REG_14__SCAN_IN), .B2(keyinput39), .ZN(n10231) );
  OAI221_X1 U11280 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(keyinput32), .C1(
        P2_REG1_REG_14__SCAN_IN), .C2(keyinput39), .A(n10231), .ZN(n10238) );
  AOI22_X1 U11281 ( .A1(P1_REG1_REG_29__SCAN_IN), .A2(keyinput63), .B1(
        P2_IR_REG_1__SCAN_IN), .B2(keyinput12), .ZN(n10232) );
  OAI221_X1 U11282 ( .B1(P1_REG1_REG_29__SCAN_IN), .B2(keyinput63), .C1(
        P2_IR_REG_1__SCAN_IN), .C2(keyinput12), .A(n10232), .ZN(n10237) );
  AOI22_X1 U11283 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(keyinput36), .B1(
        P2_D_REG_28__SCAN_IN), .B2(keyinput33), .ZN(n10233) );
  OAI221_X1 U11284 ( .B1(P1_DATAO_REG_15__SCAN_IN), .B2(keyinput36), .C1(
        P2_D_REG_28__SCAN_IN), .C2(keyinput33), .A(n10233), .ZN(n10236) );
  AOI22_X1 U11285 ( .A1(P1_REG1_REG_3__SCAN_IN), .A2(keyinput19), .B1(
        P1_D_REG_13__SCAN_IN), .B2(keyinput34), .ZN(n10234) );
  OAI221_X1 U11286 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(keyinput19), .C1(
        P1_D_REG_13__SCAN_IN), .C2(keyinput34), .A(n10234), .ZN(n10235) );
  NOR4_X1 U11287 ( .A1(n10238), .A2(n10237), .A3(n10236), .A4(n10235), .ZN(
        n10239) );
  NAND4_X1 U11288 ( .A1(n10242), .A2(n10241), .A3(n10240), .A4(n10239), .ZN(
        n10303) );
  AOI22_X1 U11289 ( .A1(n7314), .A2(keyinput20), .B1(n10244), .B2(keyinput35), 
        .ZN(n10243) );
  OAI221_X1 U11290 ( .B1(n7314), .B2(keyinput20), .C1(n10244), .C2(keyinput35), 
        .A(n10243), .ZN(n10249) );
  XNOR2_X1 U11291 ( .A(n10245), .B(keyinput45), .ZN(n10248) );
  XNOR2_X1 U11292 ( .A(n10246), .B(keyinput15), .ZN(n10247) );
  OR3_X1 U11293 ( .A1(n10249), .A2(n10248), .A3(n10247), .ZN(n10258) );
  AOI22_X1 U11294 ( .A1(n10252), .A2(keyinput37), .B1(n10251), .B2(keyinput24), 
        .ZN(n10250) );
  OAI221_X1 U11295 ( .B1(n10252), .B2(keyinput37), .C1(n10251), .C2(keyinput24), .A(n10250), .ZN(n10257) );
  INV_X1 U11296 ( .A(SI_29_), .ZN(n10254) );
  AOI22_X1 U11297 ( .A1(n10255), .A2(keyinput26), .B1(keyinput14), .B2(n10254), 
        .ZN(n10253) );
  OAI221_X1 U11298 ( .B1(n10255), .B2(keyinput26), .C1(n10254), .C2(keyinput14), .A(n10253), .ZN(n10256) );
  NOR3_X1 U11299 ( .A1(n10258), .A2(n10257), .A3(n10256), .ZN(n10301) );
  AOI22_X1 U11300 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(keyinput55), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput53), .ZN(n10259) );
  OAI221_X1 U11301 ( .B1(P2_DATAO_REG_26__SCAN_IN), .B2(keyinput55), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput53), .A(n10259), .ZN(n10267) );
  AOI22_X1 U11302 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(keyinput2), .B1(
        P1_REG0_REG_24__SCAN_IN), .B2(keyinput11), .ZN(n10260) );
  OAI221_X1 U11303 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(keyinput2), .C1(
        P1_REG0_REG_24__SCAN_IN), .C2(keyinput11), .A(n10260), .ZN(n10266) );
  AOI22_X1 U11304 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(keyinput9), .B1(n10262), 
        .B2(keyinput17), .ZN(n10261) );
  OAI221_X1 U11305 ( .B1(P2_IR_REG_29__SCAN_IN), .B2(keyinput9), .C1(n10262), 
        .C2(keyinput17), .A(n10261), .ZN(n10265) );
  AOI22_X1 U11306 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(keyinput23), .B1(
        P2_D_REG_4__SCAN_IN), .B2(keyinput1), .ZN(n10263) );
  OAI221_X1 U11307 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(keyinput23), .C1(
        P2_D_REG_4__SCAN_IN), .C2(keyinput1), .A(n10263), .ZN(n10264) );
  NOR4_X1 U11308 ( .A1(n10267), .A2(n10266), .A3(n10265), .A4(n10264), .ZN(
        n10300) );
  AOI22_X1 U11309 ( .A1(n7395), .A2(keyinput7), .B1(keyinput42), .B2(n10269), 
        .ZN(n10268) );
  OAI221_X1 U11310 ( .B1(n7395), .B2(keyinput7), .C1(n10269), .C2(keyinput42), 
        .A(n10268), .ZN(n10276) );
  AOI22_X1 U11311 ( .A1(n10272), .A2(keyinput56), .B1(n10271), .B2(keyinput43), 
        .ZN(n10270) );
  OAI221_X1 U11312 ( .B1(n10272), .B2(keyinput56), .C1(n10271), .C2(keyinput43), .A(n10270), .ZN(n10275) );
  XNOR2_X1 U11313 ( .A(n10273), .B(keyinput59), .ZN(n10274) );
  OR3_X1 U11314 ( .A1(n10276), .A2(n10275), .A3(n10274), .ZN(n10283) );
  AOI22_X1 U11315 ( .A1(n10279), .A2(keyinput21), .B1(keyinput4), .B2(n10278), 
        .ZN(n10277) );
  OAI221_X1 U11316 ( .B1(n10279), .B2(keyinput21), .C1(n10278), .C2(keyinput4), 
        .A(n10277), .ZN(n10282) );
  XNOR2_X1 U11317 ( .A(n10280), .B(keyinput41), .ZN(n10281) );
  NOR3_X1 U11318 ( .A1(n10283), .A2(n10282), .A3(n10281), .ZN(n10299) );
  INV_X1 U11319 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10285) );
  AOI22_X1 U11320 ( .A1(n10285), .A2(keyinput47), .B1(n10022), .B2(keyinput50), 
        .ZN(n10284) );
  OAI221_X1 U11321 ( .B1(n10285), .B2(keyinput47), .C1(n10022), .C2(keyinput50), .A(n10284), .ZN(n10297) );
  AOI22_X1 U11322 ( .A1(n10288), .A2(keyinput30), .B1(n10287), .B2(keyinput28), 
        .ZN(n10286) );
  OAI221_X1 U11323 ( .B1(n10288), .B2(keyinput30), .C1(n10287), .C2(keyinput28), .A(n10286), .ZN(n10296) );
  AOI22_X1 U11324 ( .A1(n10291), .A2(keyinput38), .B1(keyinput62), .B2(n10290), 
        .ZN(n10289) );
  OAI221_X1 U11325 ( .B1(n10291), .B2(keyinput38), .C1(n10290), .C2(keyinput62), .A(n10289), .ZN(n10295) );
  XNOR2_X1 U11326 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput40), .ZN(n10293) );
  XNOR2_X1 U11327 ( .A(P1_REG3_REG_4__SCAN_IN), .B(keyinput31), .ZN(n10292) );
  NAND2_X1 U11328 ( .A1(n10293), .A2(n10292), .ZN(n10294) );
  NOR4_X1 U11329 ( .A1(n10297), .A2(n10296), .A3(n10295), .A4(n10294), .ZN(
        n10298) );
  NAND4_X1 U11330 ( .A1(n10301), .A2(n10300), .A3(n10299), .A4(n10298), .ZN(
        n10302) );
  AOI211_X1 U11331 ( .C1(n10305), .C2(n10304), .A(n10303), .B(n10302), .ZN(
        n10306) );
  XNOR2_X1 U11332 ( .A(n10307), .B(n10306), .ZN(P2_U3261) );
  XNOR2_X1 U11333 ( .A(n10309), .B(n10308), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11334 ( .A(n10311), .B(n10310), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11335 ( .A(n10313), .B(n10312), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11336 ( .A(n10315), .B(n10314), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11337 ( .A(n10317), .B(n10316), .ZN(ADD_1068_U48) );
  XOR2_X1 U11338 ( .A(n10319), .B(n10318), .Z(ADD_1068_U54) );
  XOR2_X1 U11339 ( .A(n10321), .B(n10320), .Z(ADD_1068_U53) );
  XNOR2_X1 U11340 ( .A(n10323), .B(n10322), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4839 ( .A(n4527), .Z(n4329) );
  CLKBUF_X1 U4852 ( .A(n6114), .Z(n4333) );
  CLKBUF_X1 U4856 ( .A(n6114), .Z(n4332) );
  CLKBUF_X1 U4859 ( .A(n6617), .Z(n4337) );
endmodule

