

module b22_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P3_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, 
        P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN, 
        P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN, 
        P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN, 
        P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN, 
        P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN, 
        P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN, 
        P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN, 
        P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN, 
        P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN, 
        P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN,
         P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN,
         P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN,
         P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN,
         P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN,
         P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN,
         P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN,
         P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN,
         P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN,
         P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN,
         P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN,
         P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN,
         P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN,
         P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN,
         P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN,
         P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN,
         P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN,
         P3_ADDR_REG_3__SCAN_IN, P3_ADDR_REG_4__SCAN_IN,
         P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN,
         P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN,
         P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN,
         P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN,
         P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN,
         P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN,
         P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN,
         P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN,
         P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN,
         P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN,
         P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN,
         P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN,
         P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN,
         P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN,
         P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN,
         P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN,
         P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN,
         P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN,
         P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN,
         P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN,
         P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN,
         P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN,
         P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN,
         P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN,
         P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN,
         P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN,
         P3_REG0_REG_3__SCAN_IN, P3_REG0_REG_4__SCAN_IN,
         P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN,
         P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN,
         P3_REG0_REG_9__SCAN_IN, P3_REG0_REG_10__SCAN_IN,
         P3_REG0_REG_11__SCAN_IN, P3_REG0_REG_12__SCAN_IN,
         P3_REG0_REG_13__SCAN_IN, P3_REG0_REG_14__SCAN_IN,
         P3_REG0_REG_15__SCAN_IN, P3_REG0_REG_16__SCAN_IN,
         P3_REG0_REG_17__SCAN_IN, P3_REG0_REG_18__SCAN_IN,
         P3_REG0_REG_19__SCAN_IN, P3_REG0_REG_20__SCAN_IN,
         P3_REG0_REG_21__SCAN_IN, P3_REG0_REG_22__SCAN_IN,
         P3_REG0_REG_23__SCAN_IN, P3_REG0_REG_24__SCAN_IN,
         P3_REG0_REG_25__SCAN_IN, P3_REG0_REG_26__SCAN_IN,
         P3_REG0_REG_27__SCAN_IN, P3_REG0_REG_28__SCAN_IN,
         P3_REG0_REG_29__SCAN_IN, P3_REG0_REG_30__SCAN_IN,
         P3_REG0_REG_31__SCAN_IN, P3_REG1_REG_0__SCAN_IN,
         P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN,
         P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN,
         P3_REG1_REG_5__SCAN_IN, P3_REG1_REG_6__SCAN_IN,
         P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN,
         P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN,
         P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN,
         P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN,
         P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN,
         P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN,
         P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN,
         P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN,
         P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN,
         P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN,
         P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN,
         P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN,
         P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN,
         P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN,
         P3_REG2_REG_3__SCAN_IN, P3_REG2_REG_4__SCAN_IN,
         P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN,
         P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN,
         P3_REG2_REG_9__SCAN_IN, P3_REG2_REG_10__SCAN_IN,
         P3_REG2_REG_11__SCAN_IN, P3_REG2_REG_12__SCAN_IN,
         P3_REG2_REG_13__SCAN_IN, P3_REG2_REG_14__SCAN_IN,
         P3_REG2_REG_15__SCAN_IN, P3_REG2_REG_16__SCAN_IN,
         P3_REG2_REG_17__SCAN_IN, P3_REG2_REG_18__SCAN_IN,
         P3_REG2_REG_19__SCAN_IN, P3_REG2_REG_20__SCAN_IN,
         P3_REG2_REG_21__SCAN_IN, P3_REG2_REG_22__SCAN_IN,
         P3_REG2_REG_23__SCAN_IN, P3_REG2_REG_24__SCAN_IN,
         P3_REG2_REG_25__SCAN_IN, P3_REG2_REG_26__SCAN_IN,
         P3_REG2_REG_27__SCAN_IN, P3_REG2_REG_28__SCAN_IN,
         P3_REG2_REG_29__SCAN_IN, P3_REG2_REG_30__SCAN_IN,
         P3_REG2_REG_31__SCAN_IN, P3_ADDR_REG_19__SCAN_IN,
         P3_ADDR_REG_18__SCAN_IN, P3_ADDR_REG_17__SCAN_IN,
         P3_ADDR_REG_16__SCAN_IN, P3_ADDR_REG_15__SCAN_IN,
         P3_ADDR_REG_14__SCAN_IN, P3_ADDR_REG_13__SCAN_IN,
         P3_ADDR_REG_12__SCAN_IN, P3_ADDR_REG_11__SCAN_IN,
         P3_ADDR_REG_10__SCAN_IN;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165;

  AOI211_X1 U7278 ( .C1(n14918), .C2(n14917), .A(n16060), .B(n14916), .ZN(
        n14919) );
  AND2_X1 U7279 ( .A1(n14865), .A2(n7995), .ZN(n12541) );
  NOR2_X1 U7280 ( .A1(n14250), .A2(n7796), .ZN(n7795) );
  OR2_X1 U7281 ( .A1(n12973), .A2(n12974), .ZN(n12975) );
  OR2_X1 U7282 ( .A1(n11159), .A2(n13208), .ZN(n11185) );
  NAND2_X1 U7283 ( .A1(n11724), .A2(n11723), .ZN(n14526) );
  NAND2_X1 U7284 ( .A1(n10717), .A2(n10716), .ZN(n10793) );
  CLKBUF_X2 U7285 ( .A(n10225), .Z(n12519) );
  NAND2_X1 U7286 ( .A1(n10689), .A2(n10688), .ZN(n13190) );
  INV_X1 U7287 ( .A(n13059), .ZN(n14836) );
  NAND2_X2 U7288 ( .A1(n8968), .A2(n15165), .ZN(n10077) );
  CLKBUF_X2 U7289 ( .A(n8405), .Z(n8590) );
  AND2_X1 U7291 ( .A1(n9279), .A2(n15149), .ZN(n9340) );
  INV_X2 U7292 ( .A(n12239), .ZN(n13321) );
  MUX2_X1 U7293 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9070), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n9071) );
  INV_X2 U7294 ( .A(n7177), .ZN(n7180) );
  NAND2_X1 U7295 ( .A1(n9489), .A2(n9488), .ZN(n13408) );
  NOR2_X1 U7296 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n8940) );
  AND4_X1 U7297 ( .A1(n7879), .A2(n7878), .A3(n9650), .A4(n7880), .ZN(n7548)
         );
  AND2_X1 U7298 ( .A1(n7883), .A2(n9649), .ZN(n7549) );
  NOR2_X1 U7299 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n7881) );
  NOR2_X1 U7300 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n7334) );
  INV_X1 U7301 ( .A(n9956), .ZN(n9827) );
  NAND2_X1 U7302 ( .A1(n15874), .A2(n15912), .ZN(n12657) );
  NAND2_X1 U7303 ( .A1(n12596), .A2(n13670), .ZN(n10528) );
  INV_X1 U7304 ( .A(n7177), .ZN(n7179) );
  INV_X1 U7305 ( .A(n13411), .ZN(n8046) );
  INV_X1 U7306 ( .A(n9340), .ZN(n10239) );
  NAND2_X1 U7307 ( .A1(n12800), .A2(n12993), .ZN(n12808) );
  OR2_X1 U7308 ( .A1(n12885), .A2(n11454), .ZN(n11455) );
  OAI21_X1 U7309 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(n15514), .A(n15513), .ZN(
        n15525) );
  NAND2_X1 U7310 ( .A1(n8703), .A2(n13453), .ZN(n13455) );
  INV_X1 U7311 ( .A(n13656), .ZN(n13670) );
  INV_X1 U7312 ( .A(n8227), .ZN(n8226) );
  INV_X1 U7313 ( .A(n8605), .ZN(n12573) );
  INV_X1 U7314 ( .A(n13735), .ZN(n13771) );
  INV_X1 U7315 ( .A(n12762), .ZN(n12772) );
  INV_X1 U7316 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8221) );
  INV_X1 U7317 ( .A(n12339), .ZN(n13322) );
  CLKBUF_X2 U7318 ( .A(n10053), .Z(n13011) );
  NAND2_X1 U7319 ( .A1(n9291), .A2(n9290), .ZN(n9305) );
  INV_X1 U7320 ( .A(n12049), .ZN(n12008) );
  AOI21_X1 U7321 ( .B1(n13685), .B2(n13684), .A(n13683), .ZN(n13892) );
  NAND2_X1 U7322 ( .A1(n10006), .A2(n10005), .ZN(n13161) );
  OAI21_X1 U7323 ( .B1(n9310), .B2(n9285), .A(n9284), .ZN(n7942) );
  AND4_X1 U7324 ( .A1(n9309), .A2(n9308), .A3(n9307), .A4(n9306), .ZN(n10624)
         );
  AOI21_X1 U7325 ( .B1(n13055), .B2(n12163), .A(n12541), .ZN(n15039) );
  OR2_X1 U7326 ( .A1(n9282), .A2(n8947), .ZN(n9084) );
  INV_X1 U7328 ( .A(n10988), .ZN(n15874) );
  INV_X2 U7329 ( .A(n15899), .ZN(n13853) );
  OAI21_X1 U7330 ( .B1(n12418), .B2(n12374), .A(n12416), .ZN(n12422) );
  NAND2_X1 U7331 ( .A1(n15169), .A2(n12049), .ZN(n15075) );
  NAND2_X1 U7332 ( .A1(n13100), .A2(n13411), .ZN(n7177) );
  AND2_X2 U7333 ( .A1(n8958), .A2(n8957), .ZN(n15165) );
  OR2_X2 U7334 ( .A1(n13278), .A2(n13277), .ZN(n7240) );
  NAND2_X2 U7335 ( .A1(n13350), .A2(n13349), .ZN(n13368) );
  OR2_X2 U7336 ( .A1(n14940), .A2(n14939), .ZN(n7210) );
  AOI21_X2 U7337 ( .B1(n7717), .B2(n7715), .A(n7234), .ZN(n7714) );
  OR2_X2 U7338 ( .A1(n13150), .A2(n13149), .ZN(n8184) );
  OAI21_X2 U7339 ( .B1(n13472), .B2(n7849), .A(n7847), .ZN(n13440) );
  AOI21_X2 U7340 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n15550), .A(n15549), .ZN(
        n15554) );
  OR2_X2 U7341 ( .A1(n8987), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8989) );
  INV_X2 U7342 ( .A(n8987), .ZN(n8990) );
  NAND2_X2 U7343 ( .A1(n7621), .A2(n7620), .ZN(n8987) );
  INV_X2 U7344 ( .A(n12336), .ZN(n13325) );
  NAND2_X4 U7345 ( .A1(n9599), .A2(n14226), .ZN(n16107) );
  AND2_X2 U7346 ( .A1(n7665), .A2(n7664), .ZN(n13620) );
  OAI21_X2 U7347 ( .B1(n7524), .B2(n7274), .A(n7526), .ZN(n12973) );
  NOR4_X2 U7348 ( .A1(n7215), .A2(n7183), .A3(n7182), .A4(n13406), .ZN(n13414)
         );
  NAND2_X2 U7351 ( .A1(n12330), .A2(n12329), .ZN(n14250) );
  AOI21_X2 U7352 ( .B1(n10793), .B2(n10719), .A(n10718), .ZN(n10720) );
  NOR2_X2 U7353 ( .A1(n10063), .A2(n10062), .ZN(n10218) );
  XNOR2_X2 U7354 ( .A(n8292), .B(n8291), .ZN(n12193) );
  OAI21_X2 U7355 ( .B1(n10383), .B2(n10382), .A(n10381), .ZN(n10387) );
  AOI21_X2 U7356 ( .B1(n10220), .B2(n10219), .A(n10218), .ZN(n10383) );
  OAI21_X2 U7357 ( .B1(n14311), .B2(n7873), .A(n7871), .ZN(n14273) );
  AOI22_X2 U7358 ( .A1(n13708), .A2(n13710), .B1(n13971), .B2(n13725), .ZN(
        n13700) );
  OAI21_X2 U7359 ( .B1(n13721), .B2(n13722), .A(n12631), .ZN(n13708) );
  OAI22_X2 U7360 ( .A1(n9367), .A2(n9366), .B1(n9305), .B2(n9304), .ZN(n10044)
         );
  OAI21_X2 U7362 ( .B1(n7217), .B2(n7519), .A(n7520), .ZN(n12981) );
  XNOR2_X2 U7363 ( .A(n10773), .B(n15672), .ZN(n15662) );
  AOI21_X2 U7364 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n10772), .A(n10771), .ZN(
        n10773) );
  OAI22_X2 U7365 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n15527), .B1(n15526), .B2(
        n15525), .ZN(n15530) );
  AOI21_X2 U7366 ( .B1(n11382), .B2(n11381), .A(n11380), .ZN(n11684) );
  NAND2_X1 U7367 ( .A1(n11272), .A2(n11271), .ZN(n11382) );
  OR2_X2 U7368 ( .A1(n13700), .A2(n13701), .ZN(n7767) );
  OAI222_X1 U7369 ( .A1(n13083), .A2(n15289), .B1(P3_U3151), .B2(n8225), .C1(
        n13082), .C2(n12196), .ZN(P3_U3266) );
  BUF_X8 U7370 ( .A(n13007), .Z(n7178) );
  INV_X2 U7371 ( .A(n8990), .ZN(n13007) );
  OR2_X2 U7372 ( .A1(n8222), .A2(n8221), .ZN(n8224) );
  AOI22_X2 U7373 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n15532), .B1(n15531), .B2(
        n15530), .ZN(n15534) );
  OAI21_X2 U7374 ( .B1(n11684), .B2(n11683), .A(n11682), .ZN(n11706) );
  OAI21_X2 U7375 ( .B1(n11929), .B2(n11928), .A(n11927), .ZN(n11933) );
  AND2_X1 U7376 ( .A1(n7242), .A2(n7496), .ZN(n14542) );
  NAND2_X1 U7377 ( .A1(n8009), .A2(n14102), .ZN(n14106) );
  NAND2_X1 U7378 ( .A1(n7442), .A2(n12309), .ZN(n14259) );
  NAND2_X1 U7379 ( .A1(n12162), .A2(n12161), .ZN(n14863) );
  NAND2_X1 U7380 ( .A1(n14690), .A2(n14692), .ZN(n14613) );
  NAND2_X1 U7381 ( .A1(n7644), .A2(n15628), .ZN(n15638) );
  NAND2_X1 U7382 ( .A1(n12445), .A2(n12444), .ZN(n14648) );
  AOI21_X1 U7383 ( .B1(n12410), .B2(n10850), .A(n10860), .ZN(n11267) );
  NAND3_X1 U7384 ( .A1(n12401), .A2(n12402), .A3(n7559), .ZN(n12410) );
  OAI21_X1 U7385 ( .B1(n9997), .B2(n7558), .A(n7555), .ZN(n10328) );
  NAND2_X1 U7386 ( .A1(n8030), .A2(n8029), .ZN(n9997) );
  INV_X1 U7387 ( .A(n10624), .ZN(n14751) );
  NAND2_X1 U7388 ( .A1(n14196), .A2(n14416), .ZN(n9999) );
  INV_X4 U7389 ( .A(n12874), .ZN(n13015) );
  INV_X2 U7390 ( .A(n12868), .ZN(n12863) );
  INV_X2 U7391 ( .A(n12884), .ZN(n12874) );
  NAND2_X1 U7392 ( .A1(n9880), .A2(n9879), .ZN(n13127) );
  INV_X1 U7393 ( .A(n14198), .ZN(n9973) );
  INV_X2 U7394 ( .A(n7179), .ZN(n13351) );
  BUF_X4 U7395 ( .A(n7179), .Z(n13360) );
  INV_X4 U7398 ( .A(n8186), .ZN(n12526) );
  NAND2_X1 U7399 ( .A1(n9853), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9852) );
  CLKBUF_X2 U7400 ( .A(n8394), .Z(n8689) );
  INV_X1 U7401 ( .A(n12797), .ZN(n9279) );
  AND3_X1 U7402 ( .A1(n7951), .A2(n15144), .A3(n7950), .ZN(n9278) );
  BUF_X1 U7403 ( .A(n9598), .Z(n7182) );
  XNOR2_X1 U7404 ( .A(n9086), .B(P1_IR_REG_21__SCAN_IN), .ZN(n12800) );
  INV_X1 U7405 ( .A(n14218), .ZN(n14226) );
  CLKBUF_X1 U7406 ( .A(n14218), .Z(n7183) );
  AOI22_X1 U7407 ( .A1(n9286), .A2(n9077), .B1(n9076), .B2(n9075), .ZN(n9078)
         );
  NOR2_X4 U7408 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n8996) );
  AND2_X1 U7409 ( .A1(n14087), .A2(n14088), .ZN(n7337) );
  NAND2_X1 U7410 ( .A1(n14106), .A2(n7363), .ZN(n14169) );
  NAND2_X1 U7411 ( .A1(n14259), .A2(n14262), .ZN(n7797) );
  OAI21_X1 U7412 ( .B1(n12599), .B2(n8808), .A(n7766), .ZN(n13695) );
  NAND2_X1 U7413 ( .A1(n8013), .A2(n14117), .ZN(n8012) );
  AND2_X1 U7414 ( .A1(n7767), .A2(n12635), .ZN(n8808) );
  OR2_X1 U7415 ( .A1(n7993), .A2(n14863), .ZN(n7992) );
  NAND2_X1 U7416 ( .A1(n14283), .A2(n12363), .ZN(n7442) );
  AOI21_X1 U7417 ( .B1(n7795), .B2(n7793), .A(n7792), .ZN(n7791) );
  NAND2_X1 U7418 ( .A1(n7819), .A2(n7817), .ZN(n13097) );
  AOI21_X1 U7419 ( .B1(n7630), .B2(n7632), .A(n7206), .ZN(n7629) );
  NAND2_X1 U7420 ( .A1(n8015), .A2(n14030), .ZN(n8014) );
  NAND2_X1 U7421 ( .A1(n7443), .A2(n12308), .ZN(n14283) );
  XNOR2_X1 U7422 ( .A(n13010), .B(n13009), .ZN(n14581) );
  INV_X1 U7423 ( .A(n12330), .ZN(n7792) );
  NAND2_X1 U7424 ( .A1(n14691), .A2(n14693), .ZN(n14690) );
  INV_X1 U7425 ( .A(n14544), .ZN(n14076) );
  NAND2_X1 U7426 ( .A1(n12311), .A2(n12310), .ZN(n14463) );
  NAND2_X1 U7427 ( .A1(n7458), .A2(n12282), .ZN(n14319) );
  CLKBUF_X1 U7428 ( .A(n13763), .Z(n13801) );
  NOR2_X1 U7429 ( .A1(n14470), .A2(n14175), .ZN(n12362) );
  NAND2_X2 U7430 ( .A1(n7341), .A2(n12107), .ZN(n15051) );
  NAND2_X1 U7431 ( .A1(n8080), .A2(n7248), .ZN(n14700) );
  XNOR2_X1 U7432 ( .A(n12129), .B(n12180), .ZN(n14589) );
  NAND2_X1 U7433 ( .A1(n14351), .A2(n14350), .ZN(n7457) );
  XNOR2_X1 U7434 ( .A(n15638), .B(n7643), .ZN(n15640) );
  AOI21_X1 U7435 ( .B1(n12178), .B2(n12176), .A(n7356), .ZN(n12129) );
  NAND2_X1 U7436 ( .A1(n14648), .A2(n8077), .ZN(n8080) );
  NAND2_X1 U7437 ( .A1(n8007), .A2(n8006), .ZN(n12178) );
  AOI21_X1 U7438 ( .B1(n7196), .B2(n8019), .A(n7311), .ZN(n8018) );
  XNOR2_X1 U7439 ( .A(n15064), .B(n12085), .ZN(n14918) );
  OR2_X1 U7440 ( .A1(n11884), .A2(n11902), .ZN(n12154) );
  NAND2_X1 U7441 ( .A1(n7221), .A2(n7203), .ZN(n7815) );
  XNOR2_X1 U7442 ( .A(n12073), .B(n12072), .ZN(n14601) );
  NAND2_X1 U7443 ( .A1(n12061), .A2(n12060), .ZN(n15069) );
  NAND2_X1 U7444 ( .A1(n12273), .A2(n12272), .ZN(n14485) );
  NAND2_X1 U7445 ( .A1(n12285), .A2(n12284), .ZN(n14480) );
  XNOR2_X1 U7446 ( .A(n11979), .B(SI_24_), .ZN(n12073) );
  CLKBUF_X1 U7447 ( .A(n15387), .Z(n7362) );
  NAND2_X1 U7448 ( .A1(n8566), .A2(n8565), .ZN(n13472) );
  OAI21_X1 U7449 ( .B1(n11933), .B2(n8052), .A(n8050), .ZN(n12441) );
  NAND2_X1 U7450 ( .A1(n8841), .A2(n8114), .ZN(n13807) );
  NAND2_X1 U7451 ( .A1(n7684), .A2(n7683), .ZN(n14418) );
  INV_X1 U7452 ( .A(n14417), .ZN(n7684) );
  NAND2_X1 U7453 ( .A1(n12047), .A2(n11572), .ZN(n11750) );
  NAND2_X1 U7454 ( .A1(n15590), .A2(n7343), .ZN(n15600) );
  NAND2_X1 U7455 ( .A1(n7686), .A2(n7685), .ZN(n14417) );
  NOR2_X1 U7456 ( .A1(n15727), .A2(n8327), .ZN(n15726) );
  NAND2_X1 U7457 ( .A1(n11861), .A2(n12696), .ZN(n11860) );
  NAND2_X1 U7458 ( .A1(n8829), .A2(n7307), .ZN(n8124) );
  NAND2_X1 U7459 ( .A1(n11300), .A2(n11299), .ZN(n11477) );
  XNOR2_X1 U7460 ( .A(n11263), .B(n11262), .ZN(n12233) );
  NAND2_X1 U7461 ( .A1(n11629), .A2(n11628), .ZN(n15122) );
  NAND2_X1 U7462 ( .A1(n10693), .A2(n10692), .ZN(n13203) );
  NAND2_X1 U7463 ( .A1(n11072), .A2(n11071), .ZN(n11216) );
  XNOR2_X1 U7464 ( .A(n13629), .B(n15697), .ZN(n15704) );
  AND2_X1 U7465 ( .A1(n7898), .A2(n7897), .ZN(n13629) );
  CLKBUF_X1 U7466 ( .A(n9762), .Z(n7536) );
  NAND2_X1 U7467 ( .A1(n11000), .A2(n10999), .ZN(n12864) );
  AND2_X1 U7468 ( .A1(n10393), .A2(n10678), .ZN(n10479) );
  NAND2_X1 U7469 ( .A1(n10327), .A2(n10326), .ZN(n13170) );
  OR2_X1 U7470 ( .A1(n15565), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7652) );
  NAND2_X1 U7471 ( .A1(n9876), .A2(n8031), .ZN(n8030) );
  XNOR2_X1 U7472 ( .A(n11329), .B(n15685), .ZN(n15676) );
  XNOR2_X1 U7473 ( .A(n9440), .B(SI_9_), .ZN(n9439) );
  NOR2_X1 U7474 ( .A1(n7813), .A2(n10396), .ZN(n7811) );
  AND2_X2 U7475 ( .A1(n14430), .A2(n10515), .ZN(n14378) );
  AND2_X1 U7476 ( .A1(n7900), .A2(n7899), .ZN(n11329) );
  OAI21_X1 U7477 ( .B1(n15529), .B2(n15648), .A(n15645), .ZN(n15538) );
  INV_X2 U7478 ( .A(n8410), .ZN(n13084) );
  NAND2_X1 U7479 ( .A1(n15537), .A2(n15536), .ZN(n15547) );
  INV_X4 U7482 ( .A(n12523), .ZN(n7181) );
  OR2_X1 U7483 ( .A1(n15535), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n15536) );
  NAND2_X1 U7484 ( .A1(n16107), .A2(n9600), .ZN(n11374) );
  INV_X1 U7485 ( .A(n10524), .ZN(n8787) );
  NAND4_X1 U7486 ( .A1(n9606), .A2(n9605), .A3(n9604), .A4(n9603), .ZN(n14199)
         );
  AND4_X1 U7487 ( .A1(n9295), .A2(n9294), .A3(n9293), .A4(n9292), .ZN(n12809)
         );
  NAND2_X1 U7488 ( .A1(n8227), .A2(n8228), .ZN(n8556) );
  CLKBUF_X3 U7489 ( .A(n10051), .Z(n12089) );
  AND2_X1 U7490 ( .A1(n8750), .A2(n8304), .ZN(n9220) );
  INV_X1 U7491 ( .A(n12339), .ZN(n12345) );
  AND2_X2 U7492 ( .A1(n9278), .A2(n9279), .ZN(n12095) );
  AND2_X2 U7493 ( .A1(n12797), .A2(n15149), .ZN(n12014) );
  INV_X1 U7494 ( .A(n13317), .ZN(n7677) );
  AOI21_X1 U7495 ( .B1(n7615), .B2(n7617), .A(n7273), .ZN(n7612) );
  CLKBUF_X3 U7496 ( .A(n9620), .Z(n12239) );
  AND2_X1 U7497 ( .A1(n9580), .A2(n12174), .ZN(n8182) );
  OR2_X1 U7498 ( .A1(n8951), .A2(n8950), .ZN(n8958) );
  AND2_X1 U7499 ( .A1(n7658), .A2(n9806), .ZN(n9853) );
  INV_X1 U7500 ( .A(n9278), .ZN(n15149) );
  XNOR2_X1 U7501 ( .A(n7770), .B(n14018), .ZN(n8227) );
  NOR2_X1 U7502 ( .A1(n10506), .A2(n14226), .ZN(n13100) );
  NAND2_X1 U7503 ( .A1(n8963), .A2(n9067), .ZN(n15161) );
  CLKBUF_X3 U7504 ( .A(n8767), .Z(n13664) );
  OR2_X1 U7505 ( .A1(n15170), .A2(n12800), .ZN(n15832) );
  XNOR2_X1 U7506 ( .A(n8310), .B(n8309), .ZN(n12596) );
  XNOR2_X1 U7507 ( .A(n8293), .B(n8220), .ZN(n8767) );
  XNOR2_X1 U7508 ( .A(n8453), .B(P3_IR_REG_7__SCAN_IN), .ZN(n15672) );
  NAND2_X1 U7509 ( .A1(n7211), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8293) );
  NAND2_X1 U7510 ( .A1(n9283), .A2(n9282), .ZN(n12993) );
  NAND2_X1 U7511 ( .A1(n15144), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7436) );
  NAND2_X1 U7512 ( .A1(n8967), .A2(n8966), .ZN(n15159) );
  OR2_X1 U7513 ( .A1(n9274), .A2(n7952), .ZN(n7951) );
  XNOR2_X1 U7514 ( .A(n9475), .B(n9474), .ZN(n13411) );
  NAND2_X1 U7515 ( .A1(n9282), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9086) );
  XNOR2_X1 U7516 ( .A(n9564), .B(P2_IR_REG_21__SCAN_IN), .ZN(n9598) );
  NOR2_X1 U7517 ( .A1(n8298), .A2(n8118), .ZN(n8290) );
  OR2_X1 U7518 ( .A1(n9282), .A2(n8954), .ZN(n8959) );
  NAND2_X1 U7519 ( .A1(n9803), .A2(n9802), .ZN(n9938) );
  MUX2_X1 U7520 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9487), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n9489) );
  NAND2_X1 U7521 ( .A1(n7922), .A2(n7232), .ZN(n9282) );
  XNOR2_X1 U7522 ( .A(n9287), .B(P1_IR_REG_19__SCAN_IN), .ZN(n13059) );
  XNOR2_X1 U7523 ( .A(n9566), .B(P2_IR_REG_19__SCAN_IN), .ZN(n14218) );
  OR2_X1 U7524 ( .A1(n9476), .A2(n14582), .ZN(n9564) );
  NAND2_X2 U7525 ( .A1(n9540), .A2(P2_U3088), .ZN(n14593) );
  NAND2_X2 U7526 ( .A1(n7178), .A2(P1_U3086), .ZN(n15167) );
  NAND2_X1 U7527 ( .A1(n9540), .A2(P1_U3086), .ZN(n15157) );
  NAND2_X1 U7528 ( .A1(n9540), .A2(P3_U3151), .ZN(n13083) );
  INV_X1 U7529 ( .A(n7758), .ZN(n8308) );
  AND2_X1 U7530 ( .A1(n9561), .A2(n8173), .ZN(n9476) );
  AND2_X1 U7531 ( .A1(n7787), .A2(n7784), .ZN(n9484) );
  OR2_X1 U7532 ( .A1(n9561), .A2(n14582), .ZN(n9566) );
  NAND2_X1 U7533 ( .A1(n9801), .A2(n9800), .ZN(n9924) );
  NAND2_X2 U7534 ( .A1(n7892), .A2(n7891), .ZN(n9932) );
  AND3_X1 U7535 ( .A1(n8996), .A2(n8925), .A3(n7881), .ZN(n7547) );
  AND3_X1 U7536 ( .A1(n8049), .A2(n8048), .A3(n9050), .ZN(n8938) );
  AND4_X1 U7537 ( .A1(n8217), .A2(n8216), .A3(n8215), .A4(n8572), .ZN(n8218)
         );
  AND2_X1 U7538 ( .A1(n8996), .A2(n8926), .ZN(n9014) );
  AND2_X1 U7539 ( .A1(n8953), .A2(n8952), .ZN(n8962) );
  NOR2_X1 U7540 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), .ZN(
        n8210) );
  INV_X1 U7541 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n7435) );
  NOR2_X1 U7542 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n8049) );
  NOR2_X1 U7543 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n8048) );
  NOR2_X1 U7544 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n8212) );
  NOR2_X1 U7545 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8211) );
  INV_X4 U7546 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X4 U7547 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X2 U7548 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n8386) );
  NOR2_X1 U7549 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .ZN(
        n8217) );
  NOR2_X1 U7550 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n8216) );
  NOR2_X1 U7551 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), .ZN(
        n8215) );
  INV_X1 U7552 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8417) );
  INV_X1 U7553 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8572) );
  NOR2_X2 U7554 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n9650) );
  INV_X1 U7555 ( .A(n12523), .ZN(n12514) );
  XNOR2_X2 U7556 ( .A(n11352), .B(n11223), .ZN(n11350) );
  NAND2_X2 U7557 ( .A1(n11222), .A2(n11221), .ZN(n11352) );
  NOR2_X2 U7558 ( .A1(n10787), .A2(n13190), .ZN(n10788) );
  OAI21_X2 U7559 ( .B1(n11453), .B2(n7710), .A(n7708), .ZN(n11670) );
  AOI21_X2 U7560 ( .B1(n15604), .B2(n15603), .A(n15602), .ZN(n15611) );
  AOI21_X1 U7561 ( .B1(n15128), .B2(n16071), .A(n7949), .ZN(n7948) );
  OR4_X2 U7562 ( .A1(n14282), .A2(n13398), .A3(n14310), .A4(n13397), .ZN(
        n13399) );
  NOR2_X2 U7563 ( .A1(n10936), .A2(n10935), .ZN(n10938) );
  NOR2_X1 U7564 ( .A1(n15923), .A2(n15924), .ZN(n15922) );
  OAI22_X2 U7565 ( .A1(n10048), .A2(n10047), .B1(n10046), .B2(n10045), .ZN(
        n15923) );
  NOR2_X2 U7566 ( .A1(n11455), .A2(n16128), .ZN(n11638) );
  BUF_X1 U7567 ( .A(n14869), .Z(n7184) );
  INV_X4 U7570 ( .A(n13360), .ZN(n7188) );
  NAND2_X1 U7571 ( .A1(n9637), .A2(n9437), .ZN(n7627) );
  INV_X1 U7572 ( .A(n7626), .ZN(n7625) );
  INV_X1 U7573 ( .A(n9133), .ZN(n7617) );
  OR2_X1 U7574 ( .A1(n13432), .A2(n13811), .ZN(n13778) );
  INV_X1 U7575 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8219) );
  INV_X1 U7576 ( .A(n13392), .ZN(n7886) );
  NAND2_X1 U7577 ( .A1(n11785), .A2(n9540), .ZN(n13317) );
  NAND2_X1 U7578 ( .A1(n11459), .A2(n7709), .ZN(n11460) );
  AOI22_X2 U7579 ( .A1(n11393), .A2(n11394), .B1(n8463), .B2(n13572), .ZN(
        n11466) );
  AND2_X1 U7580 ( .A1(n8704), .A2(n8702), .ZN(n13453) );
  INV_X1 U7581 ( .A(n8590), .ZN(n8887) );
  XNOR2_X1 U7582 ( .A(n13153), .B(n14032), .ZN(n9998) );
  INV_X1 U7583 ( .A(n12014), .ZN(n12992) );
  XNOR2_X1 U7584 ( .A(n14871), .B(n14882), .ZN(n14862) );
  NAND2_X1 U7585 ( .A1(n12049), .A2(n7178), .ZN(n12994) );
  AND2_X1 U7586 ( .A1(n13226), .A2(n13225), .ZN(n8143) );
  NAND2_X1 U7587 ( .A1(n8144), .A2(n8145), .ZN(n8142) );
  INV_X1 U7588 ( .A(n13226), .ZN(n8144) );
  NAND2_X1 U7589 ( .A1(n8138), .A2(n8131), .ZN(n8136) );
  INV_X1 U7590 ( .A(n13241), .ZN(n8131) );
  NAND2_X1 U7591 ( .A1(n12954), .A2(n12951), .ZN(n7913) );
  AND2_X1 U7592 ( .A1(n12953), .A2(n7915), .ZN(n7914) );
  INV_X1 U7593 ( .A(n12951), .ZN(n7915) );
  AOI21_X1 U7594 ( .B1(n13278), .B2(n13277), .A(n13275), .ZN(n13276) );
  INV_X1 U7595 ( .A(n8258), .ZN(n7722) );
  NAND2_X1 U7596 ( .A1(n7743), .A2(n7742), .ZN(n12770) );
  NOR2_X1 U7597 ( .A1(n13722), .A2(n12767), .ZN(n7742) );
  NAND2_X1 U7598 ( .A1(n13312), .A2(n7198), .ZN(n8166) );
  NOR2_X1 U7599 ( .A1(n7633), .A2(n7543), .ZN(n7542) );
  NAND2_X1 U7600 ( .A1(n7985), .A2(n10886), .ZN(n7633) );
  INV_X1 U7601 ( .A(n7616), .ZN(n7615) );
  OAI21_X1 U7602 ( .B1(n9130), .B2(n7617), .A(n9173), .ZN(n7616) );
  INV_X1 U7603 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n15514) );
  OAI21_X1 U7604 ( .B1(n10184), .B2(n7584), .A(n7585), .ZN(n10766) );
  NAND2_X1 U7605 ( .A1(n10186), .A2(n7901), .ZN(n7585) );
  NAND2_X1 U7606 ( .A1(n7205), .A2(n7901), .ZN(n7584) );
  NAND2_X1 U7607 ( .A1(n10772), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7901) );
  NAND2_X1 U7608 ( .A1(n15796), .A2(n7329), .ZN(n7571) );
  NAND2_X1 U7609 ( .A1(n7573), .A2(n7329), .ZN(n7572) );
  AND2_X1 U7610 ( .A1(n7763), .A2(n8881), .ZN(n7762) );
  OR2_X1 U7611 ( .A1(n8909), .A2(n13681), .ZN(n12774) );
  AND2_X1 U7612 ( .A1(n8100), .A2(n8102), .ZN(n8895) );
  NOR2_X1 U7613 ( .A1(n12599), .A2(n8101), .ZN(n8100) );
  INV_X1 U7614 ( .A(n8103), .ZN(n8101) );
  OR2_X1 U7615 ( .A1(n13788), .A2(n13799), .ZN(n12748) );
  OR2_X1 U7616 ( .A1(n13514), .A2(n13824), .ZN(n12738) );
  INV_X1 U7617 ( .A(n8098), .ZN(n8097) );
  OAI21_X1 U7618 ( .B1(n8825), .B2(n8099), .A(n8827), .ZN(n8098) );
  OR2_X1 U7619 ( .A1(n8485), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8502) );
  NAND2_X1 U7620 ( .A1(n8278), .A2(n8277), .ZN(n8279) );
  INV_X1 U7621 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8214) );
  NOR2_X1 U7622 ( .A1(n8248), .A2(n7405), .ZN(n7404) );
  INV_X1 U7623 ( .A(n8246), .ZN(n7405) );
  NOR2_X1 U7624 ( .A1(n7200), .A2(n7270), .ZN(n7553) );
  NAND2_X1 U7625 ( .A1(n8164), .A2(n8166), .ZN(n8163) );
  NAND2_X1 U7626 ( .A1(n14358), .A2(n14357), .ZN(n12358) );
  OR2_X1 U7627 ( .A1(n14409), .A2(n14408), .ZN(n7805) );
  NAND2_X1 U7628 ( .A1(n7549), .A2(n7545), .ZN(n7882) );
  AND2_X1 U7629 ( .A1(n9650), .A2(n8925), .ZN(n7545) );
  NOR2_X1 U7630 ( .A1(n7706), .A2(n14966), .ZN(n7704) );
  OR2_X1 U7631 ( .A1(n15086), .A2(n14637), .ZN(n12035) );
  INV_X1 U7632 ( .A(n7961), .ZN(n7959) );
  NAND2_X1 U7633 ( .A1(n9416), .A2(n10936), .ZN(n12815) );
  INV_X1 U7634 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9066) );
  AND2_X1 U7635 ( .A1(n12105), .A2(n11986), .ZN(n8006) );
  XNOR2_X1 U7636 ( .A(n11088), .B(n15207), .ZN(n11086) );
  NAND2_X1 U7637 ( .A1(n7537), .A2(n7541), .ZN(n10024) );
  INV_X1 U7638 ( .A(n7543), .ZN(n7541) );
  AND2_X1 U7639 ( .A1(n10023), .A2(n9765), .ZN(n10021) );
  NAND2_X1 U7640 ( .A1(n9131), .A2(n7615), .ZN(n7613) );
  NAND2_X1 U7641 ( .A1(n8202), .A2(n8201), .ZN(n8692) );
  INV_X1 U7642 ( .A(n8674), .ZN(n8202) );
  AND2_X1 U7643 ( .A1(n8649), .A2(n8648), .ZN(n8655) );
  OR2_X1 U7644 ( .A1(n8647), .A2(n8646), .ZN(n8648) );
  CLKBUF_X1 U7645 ( .A(n8556), .Z(n8889) );
  AND2_X1 U7646 ( .A1(n8227), .A2(n8225), .ZN(n8438) );
  OR2_X1 U7647 ( .A1(n10769), .A2(n10768), .ZN(n7900) );
  NOR2_X1 U7648 ( .A1(n15676), .A2(n11319), .ZN(n15675) );
  NAND2_X1 U7649 ( .A1(n7588), .A2(n7587), .ZN(n7898) );
  INV_X1 U7650 ( .A(n11332), .ZN(n7587) );
  OR2_X1 U7651 ( .A1(n15694), .A2(n11863), .ZN(n7679) );
  OAI21_X1 U7652 ( .B1(n7574), .B2(n13641), .A(n7904), .ZN(n15820) );
  OR2_X1 U7653 ( .A1(n15820), .A2(n15819), .ZN(n7582) );
  NAND2_X1 U7654 ( .A1(n7581), .A2(n13643), .ZN(n13655) );
  NAND2_X1 U7655 ( .A1(n7582), .A2(n7904), .ZN(n7581) );
  NAND2_X1 U7656 ( .A1(n13094), .A2(n7408), .ZN(n7407) );
  AND2_X1 U7657 ( .A1(n8234), .A2(n8233), .ZN(n13678) );
  NAND2_X1 U7658 ( .A1(n8844), .A2(n8843), .ZN(n13782) );
  NAND2_X1 U7659 ( .A1(n13807), .A2(n8170), .ZN(n8844) );
  OR2_X1 U7660 ( .A1(n8345), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8485) );
  INV_X1 U7661 ( .A(n8689), .ZN(n12584) );
  INV_X1 U7662 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8223) );
  NAND2_X1 U7663 ( .A1(n8119), .A2(n8220), .ZN(n8118) );
  INV_X1 U7664 ( .A(n8121), .ZN(n8119) );
  INV_X1 U7665 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8291) );
  NAND2_X1 U7666 ( .A1(n8876), .A2(n8875), .ZN(n8883) );
  OAI21_X1 U7667 ( .B1(n8598), .B2(n8270), .A(n8271), .ZN(n8612) );
  OR2_X1 U7668 ( .A1(n8311), .A2(P3_IR_REG_19__SCAN_IN), .ZN(n8314) );
  NAND2_X1 U7669 ( .A1(n8254), .A2(n8253), .ZN(n8339) );
  XNOR2_X1 U7670 ( .A(n8340), .B(n8492), .ZN(n13628) );
  NAND2_X1 U7671 ( .A1(n7400), .A2(n7397), .ZN(n8465) );
  INV_X1 U7672 ( .A(n7398), .ZN(n7397) );
  OAI21_X1 U7673 ( .B1(n9137), .B2(P2_DATAO_REG_7__SCAN_IN), .A(n7399), .ZN(
        n7398) );
  OAI21_X1 U7674 ( .B1(n8375), .B2(n8239), .A(n8240), .ZN(n8416) );
  AND2_X1 U7675 ( .A1(n9018), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8239) );
  OAI211_X1 U7676 ( .C1(n16107), .C2(n15904), .A(n7566), .B(n7565), .ZN(n9607)
         );
  NAND2_X1 U7677 ( .A1(n7678), .A2(n13099), .ZN(n7565) );
  NAND2_X1 U7678 ( .A1(n16107), .A2(n7567), .ZN(n7566) );
  AND2_X1 U7679 ( .A1(n15904), .A2(n9600), .ZN(n7567) );
  OR2_X1 U7681 ( .A1(n9617), .A2(n9616), .ZN(n9618) );
  AND2_X1 U7682 ( .A1(n8033), .A2(n8034), .ZN(n8029) );
  INV_X1 U7683 ( .A(n9898), .ZN(n8033) );
  NAND2_X1 U7684 ( .A1(n7471), .A2(n7469), .ZN(n14311) );
  NAND2_X1 U7685 ( .A1(n7470), .A2(n12360), .ZN(n7469) );
  OR2_X1 U7686 ( .A1(n14358), .A2(n7472), .ZN(n7471) );
  INV_X1 U7687 ( .A(n7473), .ZN(n7470) );
  XNOR2_X1 U7688 ( .A(n14475), .B(n14104), .ZN(n14310) );
  AOI21_X1 U7689 ( .B1(n7194), .B2(n7479), .A(n7257), .ZN(n7478) );
  INV_X1 U7690 ( .A(n7884), .ZN(n7479) );
  INV_X1 U7691 ( .A(n7194), .ZN(n7480) );
  NAND2_X1 U7692 ( .A1(n7440), .A2(n11544), .ZN(n11733) );
  OR2_X1 U7693 ( .A1(n11542), .A2(n11541), .ZN(n7440) );
  NAND2_X2 U7694 ( .A1(n9960), .A2(n9959), .ZN(n13153) );
  NAND2_X1 U7695 ( .A1(n9975), .A2(n9974), .ZN(n10510) );
  INV_X1 U7696 ( .A(n10870), .ZN(n7675) );
  INV_X1 U7697 ( .A(n13329), .ZN(n14453) );
  INV_X1 U7698 ( .A(n9883), .ZN(n9957) );
  BUF_X1 U7699 ( .A(n7677), .Z(n7890) );
  INV_X2 U7700 ( .A(n11785), .ZN(n12234) );
  INV_X1 U7701 ( .A(n14483), .ZN(n16140) );
  NAND2_X1 U7702 ( .A1(n11415), .A2(n11414), .ZN(n12885) );
  INV_X1 U7703 ( .A(n12994), .ZN(n10051) );
  NAND2_X1 U7704 ( .A1(n7999), .A2(n7998), .ZN(n7997) );
  XNOR2_X1 U7705 ( .A(n14656), .B(n14664), .ZN(n13046) );
  NAND2_X1 U7706 ( .A1(n11622), .A2(n11621), .ZN(n11625) );
  NAND2_X1 U7707 ( .A1(n7963), .A2(n7438), .ZN(n7437) );
  NOR2_X1 U7708 ( .A1(n10923), .A2(n7439), .ZN(n7438) );
  INV_X1 U7709 ( .A(n10922), .ZN(n7439) );
  NAND2_X1 U7710 ( .A1(n10540), .A2(n9334), .ZN(n16058) );
  NAND2_X1 U7711 ( .A1(n13006), .A2(n13005), .ZN(n13010) );
  NAND2_X1 U7712 ( .A1(n7952), .A2(n9069), .ZN(n7950) );
  INV_X1 U7713 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8946) );
  NAND2_X1 U7714 ( .A1(n15626), .A2(n15627), .ZN(n7644) );
  OAI21_X1 U7715 ( .B1(n13455), .B2(n7822), .A(n7820), .ZN(n8723) );
  NAND2_X1 U7716 ( .A1(n7837), .A2(n7835), .ZN(n11868) );
  NOR2_X1 U7717 ( .A1(n7838), .A2(n7836), .ZN(n7835) );
  INV_X1 U7718 ( .A(n11869), .ZN(n7836) );
  NAND2_X1 U7719 ( .A1(n14169), .A2(n7237), .ZN(n14086) );
  INV_X1 U7720 ( .A(n8041), .ZN(n8037) );
  NAND2_X1 U7721 ( .A1(n14046), .A2(n14045), .ZN(n7335) );
  NAND2_X1 U7722 ( .A1(n7797), .A2(n7795), .ZN(n14246) );
  NAND2_X1 U7723 ( .A1(n12141), .A2(n12140), .ZN(n14857) );
  XOR2_X1 U7724 ( .A(n13058), .B(n12542), .Z(n15037) );
  NAND2_X1 U7725 ( .A1(n7991), .A2(n7994), .ZN(n7990) );
  NOR2_X1 U7726 ( .A1(n12994), .A2(n9615), .ZN(n7431) );
  AND2_X1 U7727 ( .A1(n7296), .A2(n7509), .ZN(n7508) );
  NAND2_X1 U7728 ( .A1(n12831), .A2(n12828), .ZN(n7509) );
  AND2_X1 U7729 ( .A1(n12830), .A2(n7511), .ZN(n7510) );
  INV_X1 U7730 ( .A(n12828), .ZN(n7511) );
  INV_X1 U7731 ( .A(n13162), .ZN(n7348) );
  NAND2_X1 U7732 ( .A1(n7347), .A2(n7346), .ZN(n13183) );
  INV_X1 U7733 ( .A(n13175), .ZN(n7346) );
  INV_X1 U7734 ( .A(n13176), .ZN(n7347) );
  NAND2_X1 U7735 ( .A1(n8127), .A2(n8126), .ZN(n8125) );
  INV_X1 U7736 ( .A(n13204), .ZN(n8126) );
  OAI211_X1 U7737 ( .C1(n12860), .C2(n7499), .A(n7498), .B(n12867), .ZN(n7504)
         );
  INV_X1 U7738 ( .A(n7502), .ZN(n7498) );
  INV_X1 U7739 ( .A(n7276), .ZN(n7499) );
  OAI21_X1 U7740 ( .B1(n12860), .B2(n7503), .A(n7500), .ZN(n7505) );
  NAND2_X1 U7741 ( .A1(n7276), .A2(n12866), .ZN(n7503) );
  AOI21_X1 U7742 ( .B1(n7502), .B2(n12866), .A(n7501), .ZN(n7500) );
  INV_X1 U7743 ( .A(n12865), .ZN(n7501) );
  NOR2_X1 U7744 ( .A1(n7202), .A2(n7267), .ZN(n7522) );
  NAND2_X1 U7745 ( .A1(n12886), .A2(n12888), .ZN(n7929) );
  AND2_X1 U7746 ( .A1(n8139), .A2(n13235), .ZN(n8140) );
  NAND2_X1 U7747 ( .A1(n8142), .A2(n8143), .ZN(n8139) );
  NAND2_X1 U7748 ( .A1(n7516), .A2(n12907), .ZN(n7515) );
  INV_X1 U7749 ( .A(n12908), .ZN(n7516) );
  INV_X1 U7750 ( .A(n8132), .ZN(n8137) );
  AND2_X1 U7751 ( .A1(n12921), .A2(n7514), .ZN(n7513) );
  NAND2_X1 U7752 ( .A1(n7517), .A2(n7515), .ZN(n7514) );
  AND2_X1 U7753 ( .A1(n12947), .A2(n12920), .ZN(n12921) );
  AND2_X1 U7754 ( .A1(n7518), .A2(n12908), .ZN(n7517) );
  AND2_X1 U7755 ( .A1(n12958), .A2(n7913), .ZN(n7528) );
  AND2_X1 U7756 ( .A1(n7911), .A2(n12957), .ZN(n7910) );
  NAND2_X1 U7757 ( .A1(n7914), .A2(n7913), .ZN(n7911) );
  INV_X1 U7758 ( .A(n13271), .ZN(n8155) );
  INV_X1 U7759 ( .A(n13287), .ZN(n8129) );
  INV_X1 U7760 ( .A(n13288), .ZN(n8130) );
  NAND2_X1 U7761 ( .A1(n7214), .A2(n13283), .ZN(n7490) );
  NAND2_X1 U7762 ( .A1(n12968), .A2(n12970), .ZN(n7526) );
  NAND2_X1 U7763 ( .A1(n8218), .A2(n7757), .ZN(n7756) );
  INV_X1 U7764 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7757) );
  INV_X1 U7765 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10436) );
  INV_X1 U7766 ( .A(n7727), .ZN(n7726) );
  OAI21_X1 U7767 ( .B1(n8520), .B2(n7728), .A(n8533), .ZN(n7727) );
  INV_X1 U7768 ( .A(n8262), .ZN(n7728) );
  INV_X1 U7769 ( .A(n8256), .ZN(n7396) );
  NOR2_X1 U7770 ( .A1(n7721), .A2(n7395), .ZN(n7394) );
  NOR2_X1 U7771 ( .A1(n8255), .A2(n7396), .ZN(n7395) );
  AOI21_X1 U7772 ( .B1(n7720), .B2(n7722), .A(n7316), .ZN(n7718) );
  INV_X1 U7773 ( .A(n12232), .ZN(n7804) );
  AND2_X1 U7774 ( .A1(n11220), .A2(n11260), .ZN(n11221) );
  INV_X1 U7775 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8939) );
  NAND2_X1 U7776 ( .A1(n10299), .A2(n15318), .ZN(n10433) );
  NAND2_X1 U7777 ( .A1(n9013), .A2(n7368), .ZN(n9033) );
  NAND2_X1 U7778 ( .A1(n9540), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7368) );
  NAND2_X1 U7779 ( .A1(n7178), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9013) );
  OAI21_X1 U7780 ( .B1(n15500), .B2(P1_ADDR_REG_2__SCAN_IN), .A(n15501), .ZN(
        n15502) );
  NAND2_X1 U7781 ( .A1(n12773), .A2(n12762), .ZN(n7744) );
  NAND2_X1 U7782 ( .A1(n7743), .A2(n7313), .ZN(n7741) );
  XNOR2_X1 U7783 ( .A(n10190), .B(n10174), .ZN(n10154) );
  AOI21_X1 U7784 ( .B1(P3_REG1_REG_14__SCAN_IN), .B2(n13634), .A(n15758), .ZN(
        n13635) );
  NOR2_X1 U7785 ( .A1(n8807), .A2(n7764), .ZN(n7763) );
  INV_X1 U7786 ( .A(n12635), .ZN(n7764) );
  OR2_X1 U7787 ( .A1(n13739), .A2(n13752), .ZN(n12763) );
  NOR2_X1 U7788 ( .A1(n7749), .A2(n13837), .ZN(n7748) );
  INV_X1 U7789 ( .A(n7751), .ZN(n7749) );
  NAND2_X1 U7790 ( .A1(n11959), .A2(n12709), .ZN(n15387) );
  INV_X1 U7791 ( .A(n8826), .ZN(n8099) );
  NAND2_X1 U7792 ( .A1(n12644), .A2(n12646), .ZN(n12604) );
  NAND2_X1 U7793 ( .A1(n13750), .A2(n7773), .ZN(n13743) );
  NOR2_X1 U7794 ( .A1(n13740), .A2(n7774), .ZN(n7773) );
  INV_X1 U7795 ( .A(n12758), .ZN(n7774) );
  NAND2_X1 U7796 ( .A1(n11077), .A2(n8115), .ZN(n11285) );
  NOR2_X1 U7797 ( .A1(n8116), .A2(n12668), .ZN(n8115) );
  INV_X1 U7798 ( .A(n8818), .ZN(n8116) );
  NAND2_X1 U7799 ( .A1(n11077), .A2(n8818), .ZN(n11283) );
  INV_X1 U7800 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8122) );
  NAND2_X1 U7801 ( .A1(n8299), .A2(n8301), .ZN(n8120) );
  OR2_X1 U7802 ( .A1(n8279), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8281) );
  INV_X1 U7803 ( .A(n7389), .ZN(n7388) );
  OAI21_X1 U7804 ( .B1(n8567), .B2(n7390), .A(n8268), .ZN(n7389) );
  INV_X1 U7805 ( .A(n8267), .ZN(n7390) );
  INV_X1 U7806 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n8269) );
  NOR2_X1 U7807 ( .A1(n8352), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n8493) );
  INV_X1 U7808 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8492) );
  INV_X1 U7809 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n8245) );
  INV_X1 U7810 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8123) );
  INV_X1 U7811 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8207) );
  OR4_X1 U7812 ( .A1(n14373), .A2(n14390), .A3(n14408), .A4(n13393), .ZN(
        n13394) );
  INV_X1 U7813 ( .A(n9887), .ZN(n12339) );
  OR2_X1 U7814 ( .A1(n14076), .A2(n14047), .ZN(n12330) );
  NOR2_X1 U7815 ( .A1(n13390), .A2(n7885), .ZN(n7884) );
  INV_X1 U7816 ( .A(n11720), .ZN(n7885) );
  INV_X1 U7817 ( .A(n11552), .ZN(n11550) );
  NOR2_X2 U7818 ( .A1(n11740), .A2(n14526), .ZN(n7686) );
  AND2_X1 U7819 ( .A1(n13380), .A2(n7487), .ZN(n7486) );
  NAND2_X1 U7820 ( .A1(n10969), .A2(n10557), .ZN(n7487) );
  NAND2_X1 U7821 ( .A1(n7805), .A2(n12232), .ZN(n14391) );
  NOR2_X1 U7822 ( .A1(n9486), .A2(n7785), .ZN(n7784) );
  NAND2_X1 U7823 ( .A1(n7786), .A2(n8996), .ZN(n7785) );
  OR2_X1 U7824 ( .A1(n9654), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n10305) );
  INV_X1 U7825 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8926) );
  INV_X1 U7826 ( .A(n12513), .ZN(n8063) );
  AND2_X1 U7827 ( .A1(n10049), .A2(n10050), .ZN(n7376) );
  INV_X1 U7828 ( .A(n12524), .ZN(n12518) );
  INV_X1 U7829 ( .A(n13058), .ZN(n8005) );
  NAND2_X1 U7830 ( .A1(n12555), .A2(n7603), .ZN(n7602) );
  INV_X1 U7831 ( .A(n7631), .ZN(n7630) );
  OAI21_X1 U7832 ( .B1(n14880), .B2(n7632), .A(n14862), .ZN(n7631) );
  INV_X1 U7833 ( .A(n12119), .ZN(n7632) );
  AND2_X1 U7834 ( .A1(n14918), .A2(n12159), .ZN(n7971) );
  NOR2_X1 U7835 ( .A1(n14918), .A2(n7639), .ZN(n7638) );
  INV_X1 U7836 ( .A(n12071), .ZN(n7639) );
  NOR2_X1 U7837 ( .A1(n12026), .A2(n12025), .ZN(n12024) );
  OAI21_X1 U7838 ( .B1(n7975), .B2(n7707), .A(n12157), .ZN(n7706) );
  INV_X1 U7839 ( .A(n12007), .ZN(n7956) );
  NAND2_X1 U7840 ( .A1(n7426), .A2(n7265), .ZN(n7423) );
  INV_X1 U7841 ( .A(n10281), .ZN(n7946) );
  INV_X1 U7842 ( .A(n12087), .ZN(n8008) );
  NAND2_X1 U7843 ( .A1(n8949), .A2(n8948), .ZN(n8970) );
  INV_X1 U7844 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8948) );
  NAND4_X1 U7845 ( .A1(n10892), .A2(n8943), .A3(n11094), .A4(n8942), .ZN(n8944) );
  INV_X1 U7846 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8943) );
  INV_X1 U7847 ( .A(n7542), .ZN(n7540) );
  NAND2_X1 U7848 ( .A1(n7542), .A2(n7539), .ZN(n7538) );
  NOR2_X1 U7849 ( .A1(n10295), .A2(n7989), .ZN(n7988) );
  INV_X1 U7850 ( .A(n10023), .ZN(n7989) );
  AOI21_X1 U7851 ( .B1(n9350), .B2(n9353), .A(n7534), .ZN(n7533) );
  INV_X1 U7852 ( .A(SI_9_), .ZN(n7534) );
  OAI211_X1 U7853 ( .C1(n7613), .C2(n9350), .A(n9353), .B(n7531), .ZN(n9440)
         );
  NAND2_X1 U7854 ( .A1(n9107), .A2(n9106), .ZN(n9131) );
  XNOR2_X1 U7855 ( .A(n9033), .B(n7966), .ZN(n9031) );
  INV_X1 U7856 ( .A(SI_3_), .ZN(n7966) );
  NAND3_X1 U7857 ( .A1(n8989), .A2(n8988), .A3(SI_0_), .ZN(n8992) );
  XNOR2_X1 U7858 ( .A(n15488), .B(n7344), .ZN(n15489) );
  OR2_X1 U7859 ( .A1(n15532), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n15531) );
  AOI21_X1 U7860 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n15700), .A(n15576), .ZN(
        n15583) );
  NOR2_X1 U7861 ( .A1(n15575), .A2(n15574), .ZN(n15576) );
  NOR2_X1 U7862 ( .A1(n15619), .A2(n15618), .ZN(n15629) );
  AND2_X1 U7863 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n15617), .ZN(n15618) );
  INV_X1 U7864 ( .A(n8582), .ZN(n7854) );
  NAND2_X1 U7865 ( .A1(n8200), .A2(n15253), .ZN(n8650) );
  OR2_X1 U7866 ( .A1(n8557), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8576) );
  NAND2_X1 U7867 ( .A1(n7806), .A2(n7807), .ZN(n13451) );
  AOI21_X1 U7868 ( .B1(n13480), .B2(n13559), .A(n7808), .ZN(n7807) );
  INV_X1 U7869 ( .A(n13481), .ZN(n7808) );
  NAND2_X1 U7870 ( .A1(n8414), .A2(n15874), .ZN(n7832) );
  NAND2_X1 U7871 ( .A1(n7207), .A2(n7815), .ZN(n13505) );
  NAND2_X1 U7872 ( .A1(n7856), .A2(n7310), .ZN(n7855) );
  INV_X1 U7873 ( .A(n13472), .ZN(n7856) );
  AND2_X1 U7874 ( .A1(n11206), .A2(n11203), .ZN(n7831) );
  NAND2_X1 U7875 ( .A1(n8196), .A2(n8195), .ZN(n8557) );
  INV_X1 U7876 ( .A(n8539), .ZN(n8196) );
  AND2_X1 U7877 ( .A1(n7739), .A2(n7738), .ZN(n12782) );
  NAND2_X1 U7878 ( .A1(n13675), .A2(n13556), .ZN(n7738) );
  NAND2_X1 U7879 ( .A1(n12588), .A2(n13555), .ZN(n7739) );
  NAND2_X1 U7880 ( .A1(n8750), .A2(n8749), .ZN(n8981) );
  AND2_X1 U7881 ( .A1(n8748), .A2(n8747), .ZN(n8749) );
  NAND2_X1 U7882 ( .A1(n9939), .A2(n7583), .ZN(n7896) );
  AND2_X1 U7883 ( .A1(n9834), .A2(n9790), .ZN(n7583) );
  NAND2_X1 U7884 ( .A1(n9791), .A2(n9872), .ZN(n9794) );
  NOR2_X1 U7885 ( .A1(n10194), .A2(n10193), .ZN(n10771) );
  NAND2_X1 U7886 ( .A1(n7586), .A2(n7205), .ZN(n7903) );
  OAI21_X1 U7887 ( .B1(n15662), .B2(n7660), .A(n7659), .ZN(n11308) );
  NAND2_X1 U7888 ( .A1(n7663), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7660) );
  INV_X1 U7889 ( .A(n10775), .ZN(n7663) );
  OR2_X1 U7890 ( .A1(n15662), .A2(n10761), .ZN(n7662) );
  NOR2_X1 U7891 ( .A1(n15659), .A2(n10767), .ZN(n10769) );
  NAND2_X1 U7892 ( .A1(n7352), .A2(n7351), .ZN(n15684) );
  INV_X1 U7893 ( .A(n15681), .ZN(n7351) );
  INV_X1 U7894 ( .A(n15682), .ZN(n7352) );
  OR2_X1 U7895 ( .A1(n15675), .A2(n11330), .ZN(n7588) );
  NOR2_X1 U7896 ( .A1(n15679), .A2(n11320), .ZN(n15678) );
  NAND2_X1 U7897 ( .A1(n7679), .A2(n7238), .ZN(n7358) );
  OR2_X1 U7898 ( .A1(n15714), .A2(n15715), .ZN(n15733) );
  NOR2_X1 U7899 ( .A1(n15719), .A2(n13631), .ZN(n13632) );
  OR2_X1 U7900 ( .A1(n15746), .A2(n7380), .ZN(n7379) );
  NOR2_X1 U7901 ( .A1(n15757), .A2(n13884), .ZN(n7380) );
  NAND2_X1 U7902 ( .A1(n7378), .A2(n7377), .ZN(n7665) );
  INV_X1 U7903 ( .A(n15785), .ZN(n7377) );
  INV_X1 U7904 ( .A(n15786), .ZN(n7378) );
  NOR2_X1 U7905 ( .A1(n8895), .A2(n7409), .ZN(n13677) );
  AND2_X1 U7906 ( .A1(n13898), .A2(n13678), .ZN(n7409) );
  NAND2_X1 U7907 ( .A1(n13677), .A2(n13685), .ZN(n13676) );
  NOR2_X1 U7908 ( .A1(n13685), .A2(n8880), .ZN(n7765) );
  NAND2_X1 U7909 ( .A1(n8881), .A2(n12777), .ZN(n13685) );
  NAND2_X1 U7910 ( .A1(n8102), .A2(n8103), .ZN(n8852) );
  AND2_X1 U7911 ( .A1(n12638), .A2(n13682), .ZN(n12599) );
  INV_X1 U7912 ( .A(n8692), .ZN(n8203) );
  OR2_X1 U7913 ( .A1(n8705), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8707) );
  NAND2_X1 U7914 ( .A1(n12632), .A2(n13725), .ZN(n8105) );
  INV_X1 U7915 ( .A(n13557), .ZN(n13712) );
  AND2_X1 U7916 ( .A1(n13743), .A2(n12763), .ZN(n13721) );
  AOI21_X1 U7917 ( .B1(n13763), .B2(n8801), .A(n7263), .ZN(n8806) );
  NAND2_X1 U7918 ( .A1(n8806), .A2(n7775), .ZN(n13750) );
  NOR2_X1 U7919 ( .A1(n12752), .A2(n7776), .ZN(n7775) );
  INV_X1 U7920 ( .A(n12753), .ZN(n7776) );
  OR2_X1 U7921 ( .A1(n13772), .A2(n13783), .ZN(n12753) );
  NOR2_X1 U7922 ( .A1(n13769), .A2(n8110), .ZN(n8109) );
  INV_X1 U7923 ( .A(n8845), .ZN(n8110) );
  NAND2_X1 U7924 ( .A1(n13782), .A2(n12615), .ZN(n8111) );
  AND2_X1 U7925 ( .A1(n12753), .A2(n12754), .ZN(n13769) );
  AND2_X1 U7926 ( .A1(n8842), .A2(n8840), .ZN(n8114) );
  INV_X1 U7927 ( .A(n13812), .ZN(n8842) );
  OR2_X1 U7928 ( .A1(n14003), .A2(n13564), .ZN(n12730) );
  AND2_X1 U7929 ( .A1(n12738), .A2(n12731), .ZN(n13812) );
  NAND2_X1 U7930 ( .A1(n13844), .A2(n8798), .ZN(n13827) );
  NAND2_X1 U7931 ( .A1(n13827), .A2(n13826), .ZN(n13825) );
  AOI21_X1 U7932 ( .B1(n12713), .B2(n7753), .A(n7752), .ZN(n7751) );
  INV_X1 U7933 ( .A(n12704), .ZN(n7753) );
  INV_X1 U7934 ( .A(n12713), .ZN(n7754) );
  INV_X1 U7935 ( .A(n13567), .ZN(n15393) );
  NAND2_X1 U7936 ( .A1(n11691), .A2(n8825), .ZN(n11695) );
  AND4_X1 U7937 ( .A1(n8479), .A2(n8478), .A3(n8477), .A4(n8476), .ZN(n12687)
         );
  NAND2_X1 U7938 ( .A1(n8189), .A2(n15338), .ZN(n8472) );
  INV_X1 U7939 ( .A(n8457), .ZN(n8189) );
  AND2_X1 U7940 ( .A1(n8854), .A2(n8853), .ZN(n13874) );
  AND2_X1 U7941 ( .A1(n8856), .A2(n12772), .ZN(n15876) );
  INV_X1 U7942 ( .A(n15873), .ZN(n15390) );
  INV_X1 U7943 ( .A(n15876), .ZN(n15392) );
  AND2_X1 U7944 ( .A1(n8812), .A2(n8811), .ZN(n15886) );
  NAND2_X1 U7945 ( .A1(n8886), .A2(n8885), .ZN(n8909) );
  NAND2_X1 U7946 ( .A1(n8295), .A2(n8294), .ZN(n8786) );
  OR2_X1 U7947 ( .A1(n8884), .A2(n15297), .ZN(n8294) );
  OR2_X1 U7948 ( .A1(n11828), .A2(n8689), .ZN(n8295) );
  NAND2_X1 U7949 ( .A1(n8587), .A2(n8586), .ZN(n13514) );
  NAND2_X1 U7950 ( .A1(n8307), .A2(n8306), .ZN(n8911) );
  NAND2_X1 U7951 ( .A1(n7730), .A2(n7729), .ZN(n12583) );
  AOI21_X1 U7952 ( .B1(n7731), .B2(n7733), .A(n7333), .ZN(n7729) );
  NAND2_X1 U7953 ( .A1(n8873), .A2(n8872), .ZN(n8876) );
  OAI21_X1 U7954 ( .B1(n8671), .B2(n14603), .A(n8281), .ZN(n8686) );
  INV_X1 U7955 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8301) );
  OAI21_X1 U7956 ( .B1(n8273), .B2(n7412), .A(n7410), .ZN(n8657) );
  INV_X1 U7957 ( .A(n7411), .ZN(n7410) );
  OAI21_X1 U7958 ( .B1(n7319), .B2(n7412), .A(n8276), .ZN(n7411) );
  NAND2_X1 U7959 ( .A1(n8273), .A2(n7319), .ZN(n8623) );
  NOR3_X1 U7960 ( .A1(n7189), .A2(P3_IR_REG_15__SCAN_IN), .A3(
        P3_IR_REG_18__SCAN_IN), .ZN(n7833) );
  XNOR2_X1 U7961 ( .A(n8264), .B(n10895), .ZN(n8552) );
  NAND2_X1 U7962 ( .A1(n8213), .A2(n8320), .ZN(n7810) );
  NAND2_X1 U7963 ( .A1(n8261), .A2(n8260), .ZN(n8521) );
  NAND2_X1 U7964 ( .A1(n7393), .A2(n8256), .ZN(n8497) );
  NAND2_X1 U7965 ( .A1(n8339), .A2(n8255), .ZN(n7393) );
  XNOR2_X1 U7966 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n8464) );
  INV_X1 U7967 ( .A(n7404), .ZN(n7403) );
  AOI21_X1 U7968 ( .B1(n7404), .B2(n8431), .A(n7402), .ZN(n7401) );
  INV_X1 U7969 ( .A(n8249), .ZN(n7402) );
  INV_X1 U7970 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8319) );
  AND2_X1 U7971 ( .A1(n8249), .A2(n8247), .ZN(n8366) );
  NAND2_X1 U7972 ( .A1(n8243), .A2(n8242), .ZN(n8432) );
  NAND2_X1 U7973 ( .A1(n8172), .A2(n8209), .ZN(n8433) );
  XNOR2_X1 U7974 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8236) );
  NAND2_X1 U7975 ( .A1(n7381), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8403) );
  INV_X1 U7976 ( .A(n10329), .ZN(n10334) );
  AND2_X1 U7977 ( .A1(n14177), .A2(n14416), .ZN(n8016) );
  OR2_X1 U7978 ( .A1(n10008), .A2(n10007), .ZN(n10345) );
  INV_X1 U7979 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10344) );
  OR2_X1 U7980 ( .A1(n10345), .A2(n10344), .ZN(n10453) );
  NAND2_X1 U7981 ( .A1(n8022), .A2(n8028), .ZN(n8021) );
  INV_X1 U7982 ( .A(n8025), .ZN(n8022) );
  AOI21_X1 U7983 ( .B1(n14062), .B2(n12383), .A(n8026), .ZN(n8025) );
  INV_X1 U7984 ( .A(n12388), .ZN(n8026) );
  AND2_X1 U7985 ( .A1(n14062), .A2(n8028), .ZN(n8023) );
  INV_X1 U7986 ( .A(n9996), .ZN(n7557) );
  OR2_X1 U7987 ( .A1(n11840), .A2(n11841), .ZN(n8043) );
  NAND2_X1 U7988 ( .A1(n7277), .A2(n8163), .ZN(n8162) );
  NOR2_X1 U7989 ( .A1(n13342), .A2(n8159), .ZN(n8158) );
  NAND2_X1 U7990 ( .A1(n7283), .A2(n8160), .ZN(n8159) );
  NAND2_X1 U7991 ( .A1(n8164), .A2(n8161), .ZN(n8160) );
  INV_X1 U7992 ( .A(n9622), .ZN(n12336) );
  NAND2_X1 U7993 ( .A1(n14290), .A2(n14294), .ZN(n7443) );
  AND2_X1 U7994 ( .A1(n13398), .A2(n12361), .ZN(n7874) );
  NAND2_X1 U7995 ( .A1(n14311), .A2(n14310), .ZN(n14309) );
  AND2_X1 U7996 ( .A1(n7875), .A2(n7474), .ZN(n7473) );
  NAND2_X1 U7997 ( .A1(n7877), .A2(n14350), .ZN(n7474) );
  NOR2_X1 U7998 ( .A1(n14324), .A2(n7876), .ZN(n7875) );
  INV_X1 U7999 ( .A(n12359), .ZN(n7876) );
  NAND2_X1 U8000 ( .A1(n12358), .A2(n7877), .ZN(n14334) );
  NAND2_X1 U8001 ( .A1(n7457), .A2(n7455), .ZN(n7458) );
  NOR2_X1 U8002 ( .A1(n12281), .A2(n7456), .ZN(n7455) );
  INV_X1 U8003 ( .A(n13396), .ZN(n14324) );
  AOI21_X1 U8004 ( .B1(n7866), .B2(n7868), .A(n7261), .ZN(n7865) );
  NAND2_X1 U8005 ( .A1(n14383), .A2(n14390), .ZN(n14385) );
  AOI21_X1 U8006 ( .B1(n7453), .B2(n7451), .A(n7260), .ZN(n7450) );
  INV_X1 U8007 ( .A(n7453), .ZN(n7452) );
  AOI21_X1 U8008 ( .B1(n7478), .B2(n7480), .A(n7801), .ZN(n7477) );
  NAND2_X1 U8009 ( .A1(n11721), .A2(n7884), .ZN(n11805) );
  OR2_X1 U8010 ( .A1(n11548), .A2(n13389), .ZN(n11721) );
  NOR2_X1 U8011 ( .A1(n13216), .A2(n14187), .ZN(n7862) );
  AOI21_X1 U8012 ( .B1(n13216), .B2(n7863), .A(n7861), .ZN(n7860) );
  NAND2_X1 U8013 ( .A1(n11183), .A2(n11711), .ZN(n7863) );
  NOR2_X1 U8014 ( .A1(n11183), .A2(n11711), .ZN(n7861) );
  XNOR2_X1 U8015 ( .A(n13216), .B(n14187), .ZN(n13386) );
  XNOR2_X1 U8016 ( .A(n14435), .B(n10857), .ZN(n13380) );
  OR2_X1 U8017 ( .A1(n10965), .A2(n10969), .ZN(n10963) );
  OAI21_X1 U8018 ( .B1(n10108), .B2(n10107), .A(n10109), .ZN(n10362) );
  NAND2_X1 U8019 ( .A1(n9972), .A2(n9971), .ZN(n10830) );
  INV_X1 U8020 ( .A(n14393), .ZN(n14413) );
  NAND2_X1 U8021 ( .A1(n13320), .A2(n13319), .ZN(n14232) );
  AOI21_X2 U8022 ( .B1(n12350), .B2(n14393), .A(n12349), .ZN(n14455) );
  XNOR2_X1 U8023 ( .A(n12343), .B(n13403), .ZN(n12350) );
  AOI22_X1 U8024 ( .A1(n14172), .A2(n14137), .B1(n14235), .B2(n14170), .ZN(
        n12348) );
  NAND2_X1 U8025 ( .A1(n14601), .A2(n7890), .ZN(n7535) );
  NAND2_X1 U8026 ( .A1(n12261), .A2(n12260), .ZN(n14361) );
  AND2_X1 U8027 ( .A1(n9545), .A2(n9544), .ZN(n9902) );
  NOR2_X1 U8028 ( .A1(n9573), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n9575) );
  NAND2_X1 U8029 ( .A1(n8929), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8934) );
  INV_X1 U8030 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8928) );
  INV_X1 U8031 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8927) );
  INV_X1 U8032 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n7381) );
  AND2_X1 U8033 ( .A1(n14606), .A2(n8062), .ZN(n8061) );
  OR2_X1 U8034 ( .A1(n14711), .A2(n8063), .ZN(n8062) );
  AND2_X1 U8035 ( .A1(n12475), .A2(n8074), .ZN(n8073) );
  AND2_X1 U8036 ( .A1(n14631), .A2(n14632), .ZN(n12475) );
  NAND2_X1 U8037 ( .A1(n12468), .A2(n8075), .ZN(n8074) );
  INV_X1 U8038 ( .A(n14622), .ZN(n8075) );
  INV_X1 U8039 ( .A(n12468), .ZN(n8076) );
  NAND2_X1 U8040 ( .A1(n11815), .A2(n11816), .ZN(n8084) );
  AND2_X1 U8041 ( .A1(n14673), .A2(n8069), .ZN(n8068) );
  OR2_X1 U8042 ( .A1(n14614), .A2(n8070), .ZN(n8069) );
  INV_X1 U8043 ( .A(n12492), .ZN(n8070) );
  NAND2_X1 U8044 ( .A1(n11418), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n11631) );
  NAND2_X1 U8045 ( .A1(n12443), .A2(n12442), .ZN(n8081) );
  OR2_X1 U8046 ( .A1(n12011), .A2(n14626), .ZN(n12026) );
  NOR2_X1 U8047 ( .A1(n11481), .A2(n8083), .ZN(n8082) );
  INV_X1 U8048 ( .A(n8086), .ZN(n8083) );
  AOI21_X1 U8049 ( .B1(n12432), .B2(n8051), .A(n7258), .ZN(n8050) );
  INV_X1 U8050 ( .A(n12432), .ZN(n8052) );
  NAND2_X1 U8051 ( .A1(n7369), .A2(n7935), .ZN(n13014) );
  OR2_X1 U8052 ( .A1(n13001), .A2(n7936), .ZN(n7935) );
  OR2_X1 U8053 ( .A1(n9766), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n10025) );
  NAND2_X1 U8054 ( .A1(n10077), .A2(n9064), .ZN(n9337) );
  INV_X1 U8055 ( .A(n15024), .ZN(n7599) );
  INV_X1 U8056 ( .A(n7997), .ZN(n7996) );
  OR2_X1 U8057 ( .A1(n15057), .A2(n14914), .ZN(n12102) );
  AND2_X1 U8058 ( .A1(n14894), .A2(n12160), .ZN(n7717) );
  NAND2_X1 U8059 ( .A1(n7210), .A2(n7971), .ZN(n14912) );
  OAI21_X1 U8060 ( .B1(n14959), .B2(n7419), .A(n7418), .ZN(n14930) );
  AOI21_X1 U8061 ( .B1(n7420), .B2(n7702), .A(n7259), .ZN(n7418) );
  INV_X1 U8062 ( .A(n7420), .ZN(n7419) );
  NAND2_X1 U8063 ( .A1(n14930), .A2(n14939), .ZN(n14929) );
  INV_X1 U8064 ( .A(n7972), .ZN(n7707) );
  INV_X1 U8065 ( .A(n7706), .ZN(n7705) );
  NOR2_X1 U8066 ( .A1(n12021), .A2(n7976), .ZN(n7975) );
  INV_X1 U8067 ( .A(n12156), .ZN(n7976) );
  NOR2_X1 U8068 ( .A1(n14974), .A2(n7973), .ZN(n7972) );
  INV_X1 U8069 ( .A(n7978), .ZN(n7973) );
  NAND2_X1 U8070 ( .A1(n15097), .A2(n15006), .ZN(n7978) );
  INV_X1 U8071 ( .A(n13047), .ZN(n14974) );
  OR2_X1 U8072 ( .A1(n11889), .A2(n11888), .ZN(n12011) );
  NAND2_X1 U8073 ( .A1(n12154), .A2(n12153), .ZN(n15002) );
  OR2_X1 U8074 ( .A1(n15009), .A2(n15010), .ZN(n15007) );
  AOI21_X1 U8075 ( .B1(n7962), .B2(n11669), .A(n7262), .ZN(n7961) );
  INV_X1 U8076 ( .A(n11624), .ZN(n7962) );
  NAND2_X1 U8077 ( .A1(n11460), .A2(n11428), .ZN(n11622) );
  AND2_X1 U8078 ( .A1(n13044), .A2(n11442), .ZN(n7711) );
  NAND2_X1 U8079 ( .A1(n11232), .A2(n11231), .ZN(n12875) );
  AOI21_X1 U8080 ( .B1(n7964), .B2(n7201), .A(n7256), .ZN(n11235) );
  OAI21_X1 U8081 ( .B1(n10905), .B2(n7696), .A(n7271), .ZN(n11040) );
  INV_X1 U8082 ( .A(n10995), .ZN(n7696) );
  NAND2_X1 U8083 ( .A1(n7695), .A2(n10995), .ZN(n7694) );
  NAND2_X1 U8084 ( .A1(n10920), .A2(n10919), .ZN(n7963) );
  NAND2_X1 U8085 ( .A1(n10905), .A2(n7698), .ZN(n10996) );
  INV_X1 U8086 ( .A(n7695), .ZN(n7698) );
  INV_X1 U8087 ( .A(n15003), .ZN(n14978) );
  AND2_X1 U8088 ( .A1(n10730), .A2(n10729), .ZN(n10735) );
  NAND2_X1 U8089 ( .A1(n10735), .A2(n13036), .ZN(n10905) );
  OR2_X1 U8090 ( .A1(n10469), .A2(n10468), .ZN(n10471) );
  NAND2_X1 U8091 ( .A1(n10479), .A2(n7595), .ZN(n10751) );
  NAND2_X1 U8092 ( .A1(n10672), .A2(n10281), .ZN(n10282) );
  NAND2_X1 U8093 ( .A1(n7417), .A2(n10276), .ZN(n10546) );
  OAI21_X1 U8094 ( .B1(n13028), .B2(n10933), .A(n9417), .ZN(n10250) );
  INV_X1 U8095 ( .A(n12869), .ZN(n16059) );
  INV_X1 U8096 ( .A(n16058), .ZN(n15948) );
  NAND2_X1 U8097 ( .A1(n7979), .A2(n12184), .ZN(n12189) );
  NAND2_X1 U8098 ( .A1(n12332), .A2(n12331), .ZN(n7979) );
  OR2_X1 U8099 ( .A1(n12189), .A2(n12188), .ZN(n13006) );
  INV_X1 U8100 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8950) );
  INV_X1 U8101 ( .A(n8959), .ZN(n8956) );
  OAI21_X1 U8102 ( .B1(n10024), .B2(n7984), .A(n7982), .ZN(n10887) );
  CLKBUF_X1 U8103 ( .A(n9007), .Z(n8995) );
  NAND2_X1 U8104 ( .A1(n7195), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7654) );
  INV_X1 U8105 ( .A(n15569), .ZN(n7653) );
  AOI22_X1 U8106 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n15594), .B1(n15593), 
        .B2(n15592), .ZN(n15597) );
  AND3_X1 U8107 ( .A1(n8456), .A2(n8455), .A3(n8454), .ZN(n11397) );
  AND4_X1 U8108 ( .A1(n8491), .A2(n8490), .A3(n8489), .A4(n8488), .ZN(n11961)
         );
  AND3_X1 U8109 ( .A1(n8343), .A2(n8342), .A3(n8341), .ZN(n13953) );
  NOR2_X1 U8110 ( .A1(n7812), .A2(n7811), .ZN(n10635) );
  OAI21_X1 U8111 ( .B1(n10396), .B2(n8411), .A(n7216), .ZN(n7812) );
  AND2_X1 U8112 ( .A1(n8618), .A2(n8617), .ZN(n13799) );
  OR2_X1 U8113 ( .A1(n12194), .A2(n8689), .ZN(n8879) );
  AOI21_X1 U8114 ( .B1(n7820), .B2(n7822), .A(n7818), .ZN(n7817) );
  INV_X1 U8115 ( .A(n8724), .ZN(n7818) );
  INV_X1 U8116 ( .A(n16005), .ZN(n12682) );
  NAND2_X1 U8117 ( .A1(n8625), .A2(n8624), .ZN(n13772) );
  OR2_X1 U8118 ( .A1(n8884), .A2(n15183), .ZN(n8624) );
  OR2_X1 U8119 ( .A1(n10632), .A2(n8689), .ZN(n8625) );
  AND4_X1 U8120 ( .A1(n8609), .A2(n8608), .A3(n8607), .A4(n8606), .ZN(n13811)
         );
  NAND2_X1 U8121 ( .A1(n8614), .A2(n8613), .ZN(n13788) );
  NAND2_X1 U8122 ( .A1(n8640), .A2(n8639), .ZN(n13757) );
  AND4_X1 U8123 ( .A1(n8337), .A2(n8336), .A3(n8335), .A4(n8334), .ZN(n11859)
         );
  AND2_X1 U8124 ( .A1(n8756), .A2(n9783), .ZN(n13527) );
  AND2_X1 U8125 ( .A1(n8759), .A2(n15892), .ZN(n13554) );
  NOR2_X1 U8126 ( .A1(n15748), .A2(n15747), .ZN(n15746) );
  XNOR2_X1 U8127 ( .A(n7379), .B(n16152), .ZN(n15766) );
  NOR2_X1 U8128 ( .A1(n15767), .A2(n15766), .ZN(n15765) );
  XNOR2_X1 U8129 ( .A(n13620), .B(n15816), .ZN(n15803) );
  NAND2_X1 U8130 ( .A1(n13655), .A2(n7579), .ZN(n7578) );
  NAND2_X1 U8131 ( .A1(n7580), .A2(n7582), .ZN(n7579) );
  NOR2_X1 U8132 ( .A1(n13644), .A2(n13643), .ZN(n7580) );
  NAND2_X1 U8133 ( .A1(n7577), .A2(n7576), .ZN(n7575) );
  NAND2_X1 U8134 ( .A1(n15817), .A2(n13647), .ZN(n7576) );
  INV_X1 U8135 ( .A(n13646), .ZN(n7577) );
  OR2_X1 U8136 ( .A1(n7674), .A2(n7671), .ZN(n7668) );
  AND2_X1 U8137 ( .A1(n13623), .A2(n13651), .ZN(n7674) );
  OAI211_X1 U8138 ( .C1(n15773), .C2(n13656), .A(n13659), .B(n13658), .ZN(
        n7909) );
  NAND2_X1 U8139 ( .A1(n7906), .A2(n10162), .ZN(n7905) );
  XNOR2_X1 U8140 ( .A(n13657), .B(n7907), .ZN(n7906) );
  INV_X1 U8141 ( .A(n13665), .ZN(n7907) );
  AND2_X1 U8142 ( .A1(n8515), .A2(n8514), .ZN(n11968) );
  AND3_X1 U8143 ( .A1(n8423), .A2(n8422), .A3(n8421), .ZN(n11030) );
  OR2_X1 U8144 ( .A1(n8394), .A2(n8984), .ZN(n8395) );
  INV_X1 U8145 ( .A(n8786), .ZN(n13898) );
  AND2_X1 U8146 ( .A1(n8291), .A2(n8223), .ZN(n7769) );
  AND2_X1 U8147 ( .A1(n14089), .A2(n8039), .ZN(n8038) );
  NOR2_X1 U8148 ( .A1(n8040), .A2(n14168), .ZN(n8039) );
  INV_X1 U8149 ( .A(n14085), .ZN(n8040) );
  INV_X1 U8150 ( .A(n14038), .ZN(n8010) );
  AND2_X1 U8151 ( .A1(n10003), .A2(n10002), .ZN(n10096) );
  NAND2_X1 U8152 ( .A1(n7562), .A2(n7563), .ZN(n7561) );
  NOR2_X1 U8153 ( .A1(n10030), .A2(n8032), .ZN(n8031) );
  INV_X1 U8154 ( .A(n9875), .ZN(n8032) );
  NAND2_X1 U8155 ( .A1(n8036), .A2(n8035), .ZN(n8034) );
  INV_X1 U8156 ( .A(n9881), .ZN(n8035) );
  INV_X1 U8157 ( .A(n9882), .ZN(n8036) );
  NAND2_X2 U8158 ( .A1(n9886), .A2(n9885), .ZN(n13145) );
  NAND2_X1 U8159 ( .A1(n12399), .A2(n7560), .ZN(n7559) );
  INV_X1 U8160 ( .A(n10847), .ZN(n7560) );
  NAND2_X1 U8161 ( .A1(n9887), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9623) );
  AND2_X1 U8162 ( .A1(n12334), .A2(n12333), .ZN(n13329) );
  INV_X1 U8163 ( .A(n14455), .ZN(n7889) );
  NAND2_X1 U8164 ( .A1(n11492), .A2(n11491), .ZN(n13224) );
  NAND2_X1 U8165 ( .A1(n14427), .A2(n10518), .ZN(n14366) );
  NAND2_X1 U8166 ( .A1(n12234), .A2(n9612), .ZN(n9613) );
  NAND2_X1 U8167 ( .A1(n7677), .A2(n7434), .ZN(n7676) );
  NAND2_X1 U8168 ( .A1(n13332), .A2(n13331), .ZN(n14233) );
  AND2_X2 U8169 ( .A1(n12323), .A2(n12322), .ZN(n14544) );
  AOI21_X1 U8170 ( .B1(n14457), .B2(n16140), .A(n8180), .ZN(n7496) );
  NAND2_X1 U8171 ( .A1(n9549), .A2(n9548), .ZN(n15408) );
  NAND2_X1 U8172 ( .A1(n8060), .A2(n12513), .ZN(n7367) );
  INV_X1 U8173 ( .A(n14606), .ZN(n7366) );
  NAND2_X1 U8174 ( .A1(n12368), .A2(n12089), .ZN(n11991) );
  NAND2_X1 U8175 ( .A1(n11411), .A2(n11410), .ZN(n16128) );
  NAND2_X1 U8176 ( .A1(n12131), .A2(n12130), .ZN(n15040) );
  NAND2_X1 U8177 ( .A1(n11649), .A2(n11648), .ZN(n14656) );
  NAND2_X2 U8178 ( .A1(n12075), .A2(n12074), .ZN(n15064) );
  NAND2_X1 U8179 ( .A1(n12005), .A2(n12004), .ZN(n15104) );
  NAND2_X1 U8180 ( .A1(n14594), .A2(n12089), .ZN(n7341) );
  AND2_X1 U8181 ( .A1(n15921), .A2(n15948), .ZN(n16129) );
  NAND2_X1 U8182 ( .A1(n8002), .A2(n8001), .ZN(n13072) );
  NAND2_X1 U8183 ( .A1(n12101), .A2(n12100), .ZN(n14881) );
  NAND2_X1 U8184 ( .A1(n12084), .A2(n12083), .ZN(n14900) );
  NAND2_X1 U8185 ( .A1(n12070), .A2(n12069), .ZN(n14951) );
  NAND2_X1 U8186 ( .A1(n12046), .A2(n12045), .ZN(n14981) );
  AND2_X1 U8187 ( .A1(n12134), .A2(n11995), .ZN(n14870) );
  NOR2_X1 U8188 ( .A1(n7360), .A2(n14860), .ZN(n7359) );
  OAI211_X1 U8189 ( .C1(n15037), .C2(n15933), .A(n15038), .B(n15036), .ZN(
        n15128) );
  AND2_X1 U8190 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n9077) );
  OR2_X1 U8191 ( .A1(n9086), .A2(n9082), .ZN(n9085) );
  NOR2_X1 U8192 ( .A1(n15569), .A2(n15568), .ZN(n15573) );
  NAND2_X1 U8193 ( .A1(n7651), .A2(n7650), .ZN(n15568) );
  NAND2_X1 U8194 ( .A1(n15566), .A2(n7652), .ZN(n7651) );
  XNOR2_X1 U8195 ( .A(n15578), .B(n15577), .ZN(n15579) );
  OAI21_X1 U8196 ( .B1(n15589), .B2(n15588), .A(P2_ADDR_REG_13__SCAN_IN), .ZN(
        n7343) );
  INV_X1 U8197 ( .A(n15639), .ZN(n7643) );
  NOR2_X1 U8198 ( .A1(n13129), .A2(n13128), .ZN(n13138) );
  NAND2_X1 U8199 ( .A1(n7507), .A2(n7937), .ZN(n12838) );
  OR2_X1 U8200 ( .A1(n7938), .A2(n12834), .ZN(n7937) );
  INV_X1 U8201 ( .A(n12833), .ZN(n7938) );
  NAND2_X1 U8202 ( .A1(n8146), .A2(n8148), .ZN(n13176) );
  NAND2_X1 U8203 ( .A1(n8149), .A2(n8150), .ZN(n8148) );
  OAI22_X1 U8204 ( .A1(n12846), .A2(n7940), .B1(n12847), .B2(n7939), .ZN(
        n12852) );
  INV_X1 U8205 ( .A(n12845), .ZN(n7939) );
  NOR2_X1 U8206 ( .A1(n12845), .A2(n12848), .ZN(n7940) );
  OR2_X1 U8207 ( .A1(n13186), .A2(n13187), .ZN(n8152) );
  INV_X1 U8208 ( .A(n13205), .ZN(n8127) );
  INV_X1 U8209 ( .A(n12859), .ZN(n7930) );
  OAI22_X1 U8210 ( .A1(n12871), .A2(n7934), .B1(n12872), .B2(n7933), .ZN(
        n12878) );
  INV_X1 U8211 ( .A(n12870), .ZN(n7933) );
  NOR2_X1 U8212 ( .A1(n12873), .A2(n12870), .ZN(n7934) );
  NAND2_X1 U8213 ( .A1(n7465), .A2(n7463), .ZN(n13220) );
  OAI22_X1 U8214 ( .A1(n12893), .A2(n7932), .B1(n12894), .B2(n7931), .ZN(
        n12898) );
  INV_X1 U8215 ( .A(n12892), .ZN(n7931) );
  NOR2_X1 U8216 ( .A1(n12895), .A2(n12892), .ZN(n7932) );
  AND2_X1 U8217 ( .A1(n8132), .A2(n13250), .ZN(n8134) );
  NAND2_X1 U8218 ( .A1(n13242), .A2(n13241), .ZN(n8132) );
  NAND2_X1 U8219 ( .A1(n7493), .A2(n7492), .ZN(n13237) );
  AND2_X1 U8220 ( .A1(n8142), .A2(n13236), .ZN(n7492) );
  INV_X1 U8221 ( .A(n12907), .ZN(n7518) );
  NAND2_X1 U8222 ( .A1(n12904), .A2(n12906), .ZN(n7928) );
  AND2_X1 U8223 ( .A1(n12930), .A2(n12919), .ZN(n12947) );
  NAND2_X1 U8224 ( .A1(n8128), .A2(n7247), .ZN(n13263) );
  OAI21_X1 U8225 ( .B1(n12952), .B2(n7914), .A(n7528), .ZN(n12959) );
  NAND2_X1 U8226 ( .A1(n8157), .A2(n8154), .ZN(n13278) );
  NAND2_X1 U8227 ( .A1(n8156), .A2(n8155), .ZN(n8154) );
  INV_X1 U8228 ( .A(n13272), .ZN(n8156) );
  NAND2_X1 U8229 ( .A1(n12969), .A2(n7527), .ZN(n7525) );
  NAND2_X1 U8230 ( .A1(n15848), .A2(n7222), .ZN(n13372) );
  AOI21_X1 U8231 ( .B1(n7197), .B2(n7491), .A(n7278), .ZN(n7489) );
  NOR2_X1 U8232 ( .A1(n7214), .A2(n13283), .ZN(n7491) );
  NAND2_X1 U8233 ( .A1(n12798), .A2(n12799), .ZN(n12801) );
  OR2_X1 U8234 ( .A1(n15170), .A2(n13059), .ZN(n12798) );
  INV_X1 U8235 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7619) );
  INV_X1 U8236 ( .A(n12771), .ZN(n7743) );
  INV_X1 U8237 ( .A(n13637), .ZN(n7573) );
  NAND2_X1 U8238 ( .A1(n10087), .A2(n8787), .ZN(n12644) );
  INV_X1 U8239 ( .A(n12391), .ZN(n8027) );
  INV_X1 U8240 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8925) );
  AND2_X1 U8241 ( .A1(n8926), .A2(n9483), .ZN(n7786) );
  OR2_X1 U8242 ( .A1(n9473), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n8935) );
  INV_X1 U8243 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7551) );
  NAND2_X1 U8244 ( .A1(n7921), .A2(n7920), .ZN(n12997) );
  INV_X1 U8245 ( .A(n12801), .ZN(n7921) );
  NAND2_X1 U8246 ( .A1(n12976), .A2(n12978), .ZN(n7520) );
  INV_X1 U8247 ( .A(n9760), .ZN(n7539) );
  INV_X1 U8248 ( .A(n7635), .ZN(n7634) );
  OAI21_X1 U8249 ( .B1(n7982), .B2(n7636), .A(n10888), .ZN(n7635) );
  INV_X1 U8250 ( .A(n10298), .ZN(n7986) );
  NAND2_X1 U8251 ( .A1(n10438), .A2(n10437), .ZN(n10888) );
  NAND2_X1 U8252 ( .A1(n10021), .A2(n7544), .ZN(n7543) );
  NAND2_X1 U8253 ( .A1(n9761), .A2(n9760), .ZN(n7544) );
  INV_X1 U8254 ( .A(n12618), .ZN(n7737) );
  NAND2_X1 U8255 ( .A1(n7896), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7895) );
  NAND2_X1 U8256 ( .A1(n11328), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7899) );
  NAND2_X1 U8257 ( .A1(n13628), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7897) );
  INV_X1 U8258 ( .A(n9254), .ZN(n7570) );
  NAND2_X1 U8259 ( .A1(n13622), .A2(n13651), .ZN(n7673) );
  NOR2_X1 U8260 ( .A1(n8104), .A2(n7255), .ZN(n8103) );
  NOR2_X1 U8261 ( .A1(n8851), .A2(n8105), .ZN(n8104) );
  OR2_X1 U8262 ( .A1(n13711), .A2(n7224), .ZN(n8102) );
  OR2_X1 U8263 ( .A1(n8786), .A2(n13678), .ZN(n12638) );
  INV_X1 U8264 ( .A(n11023), .ZN(n12659) );
  INV_X1 U8265 ( .A(n7732), .ZN(n7731) );
  OAI21_X1 U8266 ( .B1(n8875), .B2(n7733), .A(n12563), .ZN(n7732) );
  INV_X1 U8267 ( .A(n8882), .ZN(n7733) );
  INV_X1 U8268 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8220) );
  NAND2_X1 U8269 ( .A1(n7413), .A2(n8275), .ZN(n7412) );
  INV_X1 U8270 ( .A(n8637), .ZN(n7413) );
  INV_X1 U8271 ( .A(n8620), .ZN(n7414) );
  NAND2_X1 U8272 ( .A1(n7724), .A2(n7723), .ZN(n8264) );
  AOI21_X1 U8273 ( .B1(n7726), .B2(n7728), .A(n7317), .ZN(n7723) );
  NAND2_X1 U8274 ( .A1(n7392), .A2(n7243), .ZN(n8259) );
  NAND2_X1 U8275 ( .A1(n7394), .A2(n7396), .ZN(n7391) );
  OR2_X1 U8276 ( .A1(n8452), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8466) );
  INV_X1 U8277 ( .A(n8166), .ZN(n8165) );
  INV_X1 U8278 ( .A(n13316), .ZN(n8161) );
  INV_X1 U8279 ( .A(n13315), .ZN(n8164) );
  OR2_X1 U8280 ( .A1(n12324), .A2(n14081), .ZN(n12335) );
  NOR2_X1 U8281 ( .A1(n14470), .A2(n7690), .ZN(n7689) );
  NAND2_X1 U8282 ( .A1(n14551), .A2(n7691), .ZN(n7690) );
  NAND2_X1 U8283 ( .A1(n7877), .A2(n12360), .ZN(n7472) );
  INV_X1 U8284 ( .A(n12270), .ZN(n7456) );
  INV_X1 U8285 ( .A(n7867), .ZN(n7866) );
  OAI21_X1 U8286 ( .B1(n14390), .B2(n7868), .A(n14373), .ZN(n7867) );
  INV_X1 U8287 ( .A(n12356), .ZN(n7868) );
  OR2_X1 U8288 ( .A1(n7801), .A2(n7804), .ZN(n7800) );
  AND2_X1 U8289 ( .A1(n7454), .A2(n13392), .ZN(n7453) );
  NAND2_X1 U8290 ( .A1(n11790), .A2(n11791), .ZN(n7454) );
  INV_X1 U8291 ( .A(n11791), .ZN(n7451) );
  NAND2_X1 U8292 ( .A1(n13388), .A2(n7859), .ZN(n7858) );
  NAND2_X1 U8293 ( .A1(n7860), .A2(n7862), .ZN(n7859) );
  OR2_X1 U8294 ( .A1(n11145), .A2(n11144), .ZN(n11192) );
  NAND2_X1 U8295 ( .A1(n7783), .A2(n10562), .ZN(n7779) );
  NAND2_X1 U8296 ( .A1(n10559), .A2(n7782), .ZN(n7777) );
  INV_X1 U8297 ( .A(n10369), .ZN(n7782) );
  NAND2_X1 U8298 ( .A1(n13367), .A2(n9598), .ZN(n10506) );
  NAND2_X1 U8299 ( .A1(n7190), .A2(n13367), .ZN(n9772) );
  NAND2_X1 U8300 ( .A1(n10370), .A2(n10369), .ZN(n10560) );
  OAI21_X1 U8301 ( .B1(n8935), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8933) );
  OR2_X1 U8302 ( .A1(n9652), .A2(n14582), .ZN(n9135) );
  INV_X1 U8303 ( .A(n9014), .ZN(n9016) );
  OR2_X1 U8304 ( .A1(n9016), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n9059) );
  OAI22_X1 U8305 ( .A1(n10273), .A2(n12523), .B1(n10275), .B2(n12525), .ZN(
        n10043) );
  NOR2_X1 U8306 ( .A1(n10737), .A2(n10736), .ZN(n10911) );
  INV_X1 U8307 ( .A(n12525), .ZN(n10225) );
  INV_X1 U8308 ( .A(n11932), .ZN(n8051) );
  NOR2_X1 U8309 ( .A1(n14921), .A2(n15057), .ZN(n14884) );
  INV_X1 U8310 ( .A(n7971), .ZN(n7715) );
  AND2_X1 U8311 ( .A1(n13052), .A2(n7228), .ZN(n7420) );
  AND2_X1 U8312 ( .A1(n7610), .A2(n7609), .ZN(n7608) );
  NOR2_X1 U8313 ( .A1(n15086), .A2(n14995), .ZN(n7610) );
  NOR2_X1 U8314 ( .A1(n11651), .A2(n14656), .ZN(n7605) );
  NAND2_X1 U8315 ( .A1(n10923), .A2(n10904), .ZN(n7695) );
  NOR2_X1 U8316 ( .A1(n7944), .A2(n10258), .ZN(n7425) );
  INV_X1 U8317 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10067) );
  NAND2_X1 U8318 ( .A1(n11427), .A2(n11426), .ZN(n11459) );
  INV_X1 U8319 ( .A(n10751), .ZN(n7594) );
  NAND2_X1 U8320 ( .A1(n12181), .A2(n7980), .ZN(n12332) );
  NOR2_X1 U8321 ( .A1(n7321), .A2(n7981), .ZN(n7980) );
  INV_X1 U8322 ( .A(n12182), .ZN(n7981) );
  NAND2_X1 U8323 ( .A1(n11978), .A2(n12072), .ZN(n11981) );
  NAND2_X1 U8324 ( .A1(n11750), .A2(n11749), .ZN(n11974) );
  INV_X1 U8325 ( .A(n11351), .ZN(n8000) );
  INV_X1 U8326 ( .A(n7983), .ZN(n7982) );
  OAI21_X1 U8327 ( .B1(n7988), .B2(n7984), .A(n10433), .ZN(n7983) );
  OR2_X1 U8328 ( .A1(n9111), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n9138) );
  NAND2_X1 U8329 ( .A1(n15487), .A2(n7642), .ZN(n15499) );
  NAND2_X1 U8330 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n7344), .ZN(n7642) );
  OR2_X1 U8331 ( .A1(n15503), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n15504) );
  OAI21_X1 U8332 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(n15564), .A(n15563), .ZN(
        n15574) );
  INV_X1 U8333 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n9857) );
  AOI21_X1 U8334 ( .B1(n7852), .B2(n7851), .A(n7314), .ZN(n7850) );
  INV_X1 U8335 ( .A(n7310), .ZN(n7851) );
  NAND2_X1 U8336 ( .A1(n8199), .A2(n8198), .ZN(n8615) );
  INV_X1 U8337 ( .A(n8603), .ZN(n8199) );
  INV_X1 U8338 ( .A(n13526), .ZN(n7822) );
  AOI21_X1 U8339 ( .B1(n13526), .B2(n7821), .A(n8722), .ZN(n7820) );
  INV_X1 U8340 ( .A(n8704), .ZN(n7821) );
  OR2_X1 U8341 ( .A1(n8615), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8626) );
  INV_X1 U8342 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n15253) );
  OAI21_X1 U8343 ( .B1(n8519), .B2(n13566), .A(n8518), .ZN(n13537) );
  AND2_X1 U8344 ( .A1(n13452), .A2(n8684), .ZN(n13481) );
  INV_X1 U8345 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n15365) );
  INV_X1 U8346 ( .A(n7844), .ZN(n7841) );
  OR2_X1 U8347 ( .A1(n8480), .A2(n12687), .ZN(n7844) );
  NAND2_X1 U8348 ( .A1(n7843), .A2(n7845), .ZN(n7842) );
  INV_X1 U8349 ( .A(n11466), .ZN(n7843) );
  NAND2_X1 U8350 ( .A1(n8193), .A2(n8192), .ZN(n8504) );
  INV_X1 U8351 ( .A(n8502), .ZN(n8193) );
  NAND2_X1 U8352 ( .A1(n8194), .A2(n15272), .ZN(n8527) );
  INV_X1 U8353 ( .A(n8504), .ZN(n8194) );
  INV_X1 U8354 ( .A(SI_22_), .ZN(n15181) );
  OR2_X1 U8355 ( .A1(n8527), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8539) );
  NAND2_X1 U8356 ( .A1(n7735), .A2(n7734), .ZN(n12625) );
  INV_X1 U8357 ( .A(n12619), .ZN(n7734) );
  NOR2_X1 U8358 ( .A1(n7736), .A2(n12620), .ZN(n7735) );
  NAND2_X1 U8359 ( .A1(n12782), .A2(n7737), .ZN(n7736) );
  INV_X1 U8360 ( .A(n12625), .ZN(n12622) );
  AOI211_X1 U8361 ( .C1(n12778), .C2(n12777), .A(n12776), .B(n12775), .ZN(
        n12784) );
  NAND2_X1 U8362 ( .A1(n7744), .A2(n7740), .ZN(n12778) );
  AND2_X1 U8363 ( .A1(n12581), .A2(n12580), .ZN(n13555) );
  NAND2_X1 U8364 ( .A1(n9804), .A2(n9934), .ZN(n9933) );
  NAND2_X1 U8365 ( .A1(n7894), .A2(n9794), .ZN(n9856) );
  INV_X1 U8366 ( .A(n7895), .ZN(n7894) );
  AND2_X1 U8367 ( .A1(n10192), .A2(n10191), .ZN(n10194) );
  XNOR2_X1 U8368 ( .A(n10766), .B(n15672), .ZN(n15660) );
  OR2_X1 U8369 ( .A1(n10757), .A2(n10756), .ZN(n10759) );
  AND2_X1 U8370 ( .A1(n15684), .A2(n11324), .ZN(n11326) );
  INV_X1 U8371 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n15564) );
  NOR2_X1 U8372 ( .A1(n13611), .A2(n7680), .ZN(n13612) );
  AND2_X1 U8373 ( .A1(n13628), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7680) );
  NOR2_X1 U8374 ( .A1(n15721), .A2(n15720), .ZN(n15719) );
  AND2_X1 U8375 ( .A1(n15735), .A2(n13595), .ZN(n15753) );
  OR2_X1 U8376 ( .A1(n15790), .A2(n15789), .ZN(n15792) );
  NAND2_X1 U8377 ( .A1(n13639), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7664) );
  NAND2_X1 U8378 ( .A1(n7354), .A2(n7353), .ZN(n15809) );
  INV_X1 U8379 ( .A(n15813), .ZN(n7353) );
  INV_X1 U8380 ( .A(n15812), .ZN(n7354) );
  NAND2_X1 U8381 ( .A1(n7673), .A2(n7672), .ZN(n7671) );
  NOR2_X1 U8382 ( .A1(n15825), .A2(n7330), .ZN(n7670) );
  NAND2_X1 U8383 ( .A1(n7761), .A2(n7759), .ZN(n12587) );
  NAND2_X1 U8384 ( .A1(n7760), .A2(n8881), .ZN(n7759) );
  INV_X1 U8385 ( .A(n7765), .ZN(n7760) );
  OR2_X1 U8386 ( .A1(n13899), .A2(n13712), .ZN(n12635) );
  NAND2_X1 U8387 ( .A1(n12635), .A2(n12634), .ZN(n13701) );
  OR2_X1 U8388 ( .A1(n13711), .A2(n13710), .ZN(n8106) );
  NAND2_X1 U8389 ( .A1(n8112), .A2(n7415), .ZN(n13727) );
  NAND2_X1 U8390 ( .A1(n13722), .A2(n8113), .ZN(n8112) );
  INV_X1 U8391 ( .A(n8850), .ZN(n8113) );
  NAND2_X1 U8392 ( .A1(n13734), .A2(n8850), .ZN(n13723) );
  OR2_X1 U8393 ( .A1(n8849), .A2(n12760), .ZN(n13734) );
  OAI21_X1 U8394 ( .B1(n13782), .B2(n8108), .A(n8107), .ZN(n13749) );
  AOI21_X1 U8395 ( .B1(n8109), .B2(n13781), .A(n7264), .ZN(n8107) );
  INV_X1 U8396 ( .A(n8109), .ZN(n8108) );
  OR2_X1 U8397 ( .A1(n8804), .A2(n8803), .ZN(n13765) );
  AND3_X1 U8398 ( .A1(n8630), .A2(n8629), .A3(n8628), .ZN(n13783) );
  INV_X1 U8399 ( .A(n13800), .ZN(n13796) );
  NAND2_X1 U8400 ( .A1(n8197), .A2(n15356), .ZN(n8588) );
  OR2_X1 U8401 ( .A1(n8588), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8603) );
  AND4_X1 U8402 ( .A1(n8594), .A2(n8593), .A3(n8592), .A4(n8591), .ZN(n13824)
         );
  AND2_X1 U8403 ( .A1(n12722), .A2(n12726), .ZN(n13840) );
  AOI21_X1 U8404 ( .B1(n7748), .B2(n7754), .A(n7746), .ZN(n7745) );
  INV_X1 U8405 ( .A(n12718), .ZN(n7746) );
  INV_X1 U8406 ( .A(n13840), .ZN(n13845) );
  INV_X1 U8407 ( .A(SI_15_), .ZN(n10437) );
  NAND2_X1 U8408 ( .A1(n8096), .A2(n8095), .ZN(n11960) );
  AOI21_X1 U8409 ( .B1(n8097), .B2(n8099), .A(n7269), .ZN(n8095) );
  AND4_X1 U8410 ( .A1(n8331), .A2(n8330), .A3(n8329), .A4(n8328), .ZN(n13876)
         );
  AND2_X1 U8411 ( .A1(n12709), .A2(n12706), .ZN(n12609) );
  NAND2_X1 U8412 ( .A1(n11697), .A2(n12694), .ZN(n11861) );
  NAND2_X1 U8413 ( .A1(n8797), .A2(n7768), .ZN(n11697) );
  NOR2_X1 U8414 ( .A1(n8824), .A2(n12685), .ZN(n7768) );
  AND2_X1 U8415 ( .A1(n12694), .A2(n12695), .ZN(n12691) );
  AND3_X1 U8416 ( .A1(n8356), .A2(n8355), .A3(n8354), .ZN(n8822) );
  NAND2_X1 U8417 ( .A1(n8191), .A2(n8190), .ZN(n8345) );
  INV_X1 U8418 ( .A(n8474), .ZN(n8191) );
  INV_X1 U8419 ( .A(n8796), .ZN(n11580) );
  OR2_X1 U8420 ( .A1(n8472), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8474) );
  AOI21_X1 U8421 ( .B1(n11594), .B2(n11591), .A(n8820), .ZN(n11402) );
  AND2_X1 U8422 ( .A1(n8821), .A2(n8794), .ZN(n12603) );
  OR2_X1 U8423 ( .A1(n8441), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8457) );
  NAND2_X1 U8424 ( .A1(n8817), .A2(n7244), .ZN(n11077) );
  AND4_X1 U8425 ( .A1(n8361), .A2(n8360), .A3(n8359), .A4(n8358), .ZN(n11596)
         );
  INV_X1 U8426 ( .A(n10879), .ZN(n12600) );
  NAND2_X1 U8427 ( .A1(n15870), .A2(n8813), .ZN(n15877) );
  CLKBUF_X1 U8428 ( .A(n12604), .Z(n7361) );
  NAND2_X1 U8429 ( .A1(n10316), .A2(n10315), .ZN(n10317) );
  NAND2_X1 U8430 ( .A1(n8719), .A2(n8718), .ZN(n13899) );
  OR2_X1 U8431 ( .A1(n8884), .A2(n15301), .ZN(n8718) );
  OR2_X1 U8432 ( .A1(n11757), .A2(n8689), .ZN(n8719) );
  NAND2_X1 U8433 ( .A1(n8691), .A2(n8690), .ZN(n12632) );
  OR2_X1 U8434 ( .A1(n8884), .A2(n11982), .ZN(n8690) );
  OR2_X1 U8435 ( .A1(n11589), .A2(n8689), .ZN(n8691) );
  NAND2_X1 U8436 ( .A1(n8673), .A2(n8672), .ZN(n13479) );
  OR2_X1 U8437 ( .A1(n8884), .A2(n15201), .ZN(n8672) );
  NAND2_X1 U8438 ( .A1(n13750), .A2(n12758), .ZN(n13741) );
  AND2_X1 U8439 ( .A1(n15886), .A2(n16097), .ZN(n13944) );
  INV_X1 U8440 ( .A(n13944), .ZN(n13955) );
  INV_X1 U8441 ( .A(n16097), .ZN(n16082) );
  AND2_X1 U8442 ( .A1(n8855), .A2(n12772), .ZN(n15873) );
  INV_X1 U8443 ( .A(n16096), .ZN(n13954) );
  INV_X1 U8444 ( .A(n8751), .ZN(n8752) );
  NAND2_X1 U8445 ( .A1(n8717), .A2(n8285), .ZN(n8288) );
  NAND2_X1 U8446 ( .A1(n8288), .A2(n8287), .ZN(n8873) );
  NAND2_X1 U8447 ( .A1(n8688), .A2(n8283), .ZN(n8715) );
  NAND2_X1 U8448 ( .A1(n8715), .A2(n8714), .ZN(n8717) );
  AND2_X1 U8449 ( .A1(n8297), .A2(n7211), .ZN(n8750) );
  NAND2_X1 U8450 ( .A1(n8686), .A2(n8685), .ZN(n8688) );
  NAND2_X1 U8451 ( .A1(n8281), .A2(n8280), .ZN(n8671) );
  NAND2_X1 U8452 ( .A1(n7386), .A2(n7385), .ZN(n8598) );
  AOI21_X1 U8453 ( .B1(n7388), .B2(n7390), .A(n7328), .ZN(n7385) );
  NAND2_X1 U8454 ( .A1(n8568), .A2(n7388), .ZN(n7386) );
  NOR2_X1 U8455 ( .A1(n7189), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n7834) );
  NAND2_X1 U8456 ( .A1(n8308), .A2(n8535), .ZN(n8553) );
  XNOR2_X1 U8457 ( .A(n8259), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8318) );
  NAND2_X1 U8458 ( .A1(n8251), .A2(n8250), .ZN(n8351) );
  OR2_X1 U8459 ( .A1(n8466), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8352) );
  OAI21_X1 U8460 ( .B1(n8392), .B2(n7384), .A(n7382), .ZN(n8375) );
  INV_X1 U8461 ( .A(n8238), .ZN(n7384) );
  AOI21_X1 U8462 ( .B1(n7383), .B2(n8238), .A(n7218), .ZN(n7382) );
  AND2_X1 U8463 ( .A1(n10445), .A2(n10340), .ZN(n10341) );
  OR2_X1 U8464 ( .A1(n12312), .A2(n14050), .ZN(n12324) );
  AND2_X1 U8465 ( .A1(n11715), .A2(n11705), .ZN(n8044) );
  INV_X1 U8466 ( .A(n9711), .ZN(n9629) );
  INV_X1 U8467 ( .A(n8023), .ZN(n8019) );
  INV_X1 U8468 ( .A(n8044), .ZN(n7562) );
  NAND2_X1 U8469 ( .A1(n14055), .A2(n7225), .ZN(n8011) );
  INV_X1 U8470 ( .A(n8014), .ZN(n8013) );
  CLKBUF_X1 U8471 ( .A(n13102), .Z(n9774) );
  NAND2_X1 U8472 ( .A1(n12206), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n12274) );
  NAND2_X1 U8473 ( .A1(n10451), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n10696) );
  OR3_X1 U8474 ( .A1(n10696), .A2(n10695), .A3(n10694), .ZN(n10707) );
  INV_X1 U8475 ( .A(n8043), .ZN(n7564) );
  OR2_X1 U8476 ( .A1(n12239), .A2(n9587), .ZN(n9589) );
  OR2_X1 U8477 ( .A1(n9622), .A2(n9579), .ZN(n9582) );
  AOI21_X1 U8478 ( .B1(n14254), .B2(n12342), .A(n12328), .ZN(n14047) );
  INV_X1 U8479 ( .A(n12321), .ZN(n7796) );
  NAND2_X1 U8480 ( .A1(n7797), .A2(n12321), .ZN(n14244) );
  NAND2_X1 U8481 ( .A1(n7689), .A2(n7688), .ZN(n14274) );
  INV_X1 U8482 ( .A(n14326), .ZN(n7688) );
  NOR2_X1 U8483 ( .A1(n7692), .A2(n14326), .ZN(n14300) );
  OR2_X1 U8484 ( .A1(n14470), .A2(n14475), .ZN(n7692) );
  AOI21_X1 U8485 ( .B1(n7874), .B2(n7872), .A(n12362), .ZN(n7871) );
  INV_X1 U8486 ( .A(n7874), .ZN(n7873) );
  INV_X1 U8487 ( .A(n14310), .ZN(n7872) );
  OAI21_X1 U8488 ( .B1(n12296), .B2(n14310), .A(n7789), .ZN(n14290) );
  INV_X1 U8489 ( .A(n7790), .ZN(n7789) );
  OAI21_X1 U8490 ( .B1(n14310), .B2(n12295), .A(n12307), .ZN(n7790) );
  INV_X1 U8491 ( .A(n11795), .ZN(n11793) );
  OR3_X1 U8492 ( .A1(n12248), .A2(n14132), .A3(n12247), .ZN(n12262) );
  INV_X1 U8493 ( .A(n14577), .ZN(n7685) );
  INV_X1 U8494 ( .A(n7686), .ZN(n11806) );
  NAND2_X1 U8495 ( .A1(n11721), .A2(n11720), .ZN(n11725) );
  NAND2_X1 U8496 ( .A1(n11190), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n11497) );
  INV_X1 U8497 ( .A(n11192), .ZN(n11190) );
  OR2_X1 U8498 ( .A1(n11497), .A2(n11496), .ZN(n11552) );
  OAI21_X1 U8499 ( .B1(n11494), .B2(n11493), .A(n11495), .ZN(n11542) );
  INV_X1 U8500 ( .A(n14354), .ZN(n14137) );
  AOI21_X1 U8501 ( .B1(n7486), .B2(n7484), .A(n7230), .ZN(n7483) );
  INV_X1 U8502 ( .A(n7486), .ZN(n7485) );
  INV_X1 U8503 ( .A(n10557), .ZN(n7484) );
  NAND2_X1 U8504 ( .A1(n7373), .A2(n7372), .ZN(n10787) );
  INV_X1 U8505 ( .A(n10966), .ZN(n7373) );
  NAND2_X1 U8506 ( .A1(n7682), .A2(n7681), .ZN(n10966) );
  OAI21_X1 U8507 ( .B1(n10362), .B2(n10361), .A(n10363), .ZN(n10364) );
  NAND2_X1 U8508 ( .A1(n10364), .A2(n13378), .ZN(n10555) );
  NAND2_X1 U8509 ( .A1(n7371), .A2(n7370), .ZN(n10366) );
  INV_X1 U8510 ( .A(n13161), .ZN(n7370) );
  INV_X1 U8511 ( .A(n10110), .ZN(n7371) );
  NAND2_X1 U8512 ( .A1(n10514), .A2(n9967), .ZN(n10110) );
  NAND2_X1 U8513 ( .A1(n9966), .A2(n9965), .ZN(n10108) );
  NAND2_X1 U8514 ( .A1(n10867), .A2(n10868), .ZN(n9962) );
  AND2_X1 U8515 ( .A1(n16107), .A2(n16106), .ZN(n14483) );
  NAND2_X1 U8516 ( .A1(n12358), .A2(n12357), .ZN(n14336) );
  NAND2_X1 U8517 ( .A1(n7805), .A2(n7803), .ZN(n14394) );
  NAND2_X1 U8518 ( .A1(n9541), .A2(n7677), .ZN(n9543) );
  INV_X1 U8519 ( .A(n7788), .ZN(n7550) );
  INV_X1 U8520 ( .A(n7882), .ZN(n7552) );
  XNOR2_X1 U8521 ( .A(n8934), .B(P2_IR_REG_25__SCAN_IN), .ZN(n9546) );
  INV_X1 U8522 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n9562) );
  OR2_X1 U8523 ( .A1(n10305), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n10590) );
  AND2_X1 U8524 ( .A1(n9655), .A2(n10305), .ZN(n11137) );
  INV_X1 U8525 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10265) );
  OR2_X1 U8526 ( .A1(n11430), .A2(n11429), .ZN(n11432) );
  AOI21_X1 U8527 ( .B1(n8061), .B2(n8063), .A(n7252), .ZN(n8059) );
  OR2_X1 U8528 ( .A1(n10266), .A2(n10265), .ZN(n10481) );
  INV_X1 U8529 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10480) );
  INV_X1 U8530 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n11041) );
  NAND2_X1 U8531 ( .A1(n11121), .A2(n11122), .ZN(n8092) );
  NOR2_X1 U8532 ( .A1(n10821), .A2(n8091), .ZN(n8090) );
  INV_X1 U8533 ( .A(n10818), .ZN(n8091) );
  INV_X1 U8534 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10736) );
  OR2_X1 U8535 ( .A1(n10481), .A2(n10480), .ZN(n10737) );
  NAND2_X1 U8536 ( .A1(n9301), .A2(n9300), .ZN(n9363) );
  NAND2_X1 U8537 ( .A1(n9362), .A2(n9363), .ZN(n9361) );
  NAND2_X1 U8538 ( .A1(n14621), .A2(n14622), .ZN(n14680) );
  AOI21_X1 U8539 ( .B1(n8073), .B2(n8076), .A(n7254), .ZN(n8071) );
  NAND2_X1 U8540 ( .A1(n8088), .A2(n8087), .ZN(n8086) );
  INV_X1 U8541 ( .A(n11479), .ZN(n8087) );
  NAND2_X1 U8542 ( .A1(n14660), .A2(n14659), .ZN(n8079) );
  NOR2_X1 U8543 ( .A1(n12451), .A2(n8078), .ZN(n8077) );
  INV_X1 U8544 ( .A(n8081), .ZN(n8078) );
  XNOR2_X1 U8545 ( .A(n8003), .B(n13059), .ZN(n8002) );
  NAND2_X1 U8546 ( .A1(n13023), .A2(n8004), .ZN(n8003) );
  AND2_X1 U8547 ( .A1(n13057), .A2(n7226), .ZN(n8004) );
  INV_X1 U8548 ( .A(n13060), .ZN(n8001) );
  NOR2_X1 U8549 ( .A1(n15028), .A2(n7602), .ZN(n7601) );
  OR2_X1 U8550 ( .A1(n12540), .A2(n14862), .ZN(n7993) );
  INV_X1 U8551 ( .A(n7995), .ZN(n7991) );
  INV_X1 U8552 ( .A(n12540), .ZN(n7994) );
  INV_X1 U8553 ( .A(n7602), .ZN(n7600) );
  AND2_X1 U8554 ( .A1(n14861), .A2(n15955), .ZN(n7360) );
  OAI21_X1 U8555 ( .B1(n14879), .B2(n7632), .A(n7630), .ZN(n14855) );
  NAND2_X1 U8556 ( .A1(n14878), .A2(n12119), .ZN(n14856) );
  NAND2_X1 U8557 ( .A1(n14879), .A2(n14880), .ZN(n14878) );
  NAND2_X1 U8558 ( .A1(n14895), .A2(n12104), .ZN(n14879) );
  AND2_X1 U8559 ( .A1(n14915), .A2(n12086), .ZN(n14896) );
  NAND2_X1 U8560 ( .A1(n14896), .A2(n12103), .ZN(n14895) );
  NAND2_X1 U8561 ( .A1(n11992), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n12077) );
  INV_X1 U8562 ( .A(n12063), .ZN(n11992) );
  OR2_X1 U8563 ( .A1(n12077), .A2(n12076), .ZN(n12093) );
  NAND2_X1 U8564 ( .A1(n15013), .A2(n7606), .ZN(n14949) );
  NOR2_X1 U8565 ( .A1(n7611), .A2(n7607), .ZN(n7606) );
  INV_X1 U8566 ( .A(n7608), .ZN(n7607) );
  AOI21_X1 U8567 ( .B1(n7705), .B2(n7236), .A(n7701), .ZN(n7700) );
  NOR2_X1 U8568 ( .A1(n15082), .A2(n14981), .ZN(n7701) );
  NAND2_X1 U8569 ( .A1(n14948), .A2(n14947), .ZN(n14946) );
  NAND2_X1 U8570 ( .A1(n15013), .A2(n7610), .ZN(n14975) );
  OAI21_X1 U8571 ( .B1(n15009), .B2(n7954), .A(n7953), .ZN(n14972) );
  NAND2_X1 U8572 ( .A1(n7193), .A2(n7955), .ZN(n7954) );
  NAND2_X1 U8573 ( .A1(n7282), .A2(n7193), .ZN(n7953) );
  NAND2_X1 U8574 ( .A1(n15013), .A2(n15097), .ZN(n14990) );
  NAND2_X1 U8575 ( .A1(n7605), .A2(n7604), .ZN(n15014) );
  NAND2_X1 U8576 ( .A1(n11653), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n11889) );
  AOI21_X1 U8577 ( .B1(n7958), .B2(n13048), .A(n7235), .ZN(n7637) );
  NOR2_X1 U8578 ( .A1(n13046), .A2(n7959), .ZN(n7958) );
  INV_X1 U8579 ( .A(n7605), .ZN(n11887) );
  AOI21_X1 U8580 ( .B1(n7711), .B2(n7709), .A(n7233), .ZN(n7708) );
  INV_X1 U8581 ( .A(n7711), .ZN(n7710) );
  NAND2_X1 U8582 ( .A1(n11638), .A2(n14732), .ZN(n11651) );
  OR2_X1 U8583 ( .A1(n11247), .A2(n12875), .ZN(n11454) );
  NAND2_X1 U8584 ( .A1(n7592), .A2(n7591), .ZN(n11008) );
  INV_X1 U8585 ( .A(n10926), .ZN(n7592) );
  NAND2_X1 U8586 ( .A1(n7943), .A2(n7945), .ZN(n10744) );
  INV_X1 U8587 ( .A(n7423), .ZN(n7945) );
  OR2_X1 U8588 ( .A1(n10672), .A2(n7947), .ZN(n7943) );
  NAND2_X1 U8589 ( .A1(n10673), .A2(n13031), .ZN(n10672) );
  NOR2_X1 U8590 ( .A1(n10621), .A2(n15949), .ZN(n10677) );
  AND2_X1 U8591 ( .A1(n10682), .A2(n10677), .ZN(n10678) );
  INV_X1 U8592 ( .A(n15832), .ZN(n10540) );
  OR2_X1 U8593 ( .A1(n10620), .A2(n15918), .ZN(n10621) );
  XNOR2_X1 U8594 ( .A(n15918), .B(n14750), .ZN(n13027) );
  NAND2_X1 U8595 ( .A1(n10272), .A2(n12816), .ZN(n10619) );
  NAND2_X1 U8596 ( .A1(n12014), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n7433) );
  INV_X1 U8597 ( .A(n15854), .ZN(n10936) );
  OR2_X1 U8598 ( .A1(n10535), .A2(n10534), .ZN(n12167) );
  AND2_X1 U8599 ( .A1(n15041), .A2(n13059), .ZN(n10536) );
  INV_X1 U8600 ( .A(n15041), .ZN(n15952) );
  INV_X1 U8601 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9068) );
  BUF_X1 U8602 ( .A(n9275), .Z(n9273) );
  INV_X1 U8603 ( .A(n12179), .ZN(n7356) );
  NAND2_X1 U8604 ( .A1(n10442), .A2(n8945), .ZN(n9286) );
  XNOR2_X1 U8605 ( .A(n11989), .B(n11988), .ZN(n12368) );
  INV_X1 U8606 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9072) );
  NOR2_X1 U8607 ( .A1(n8944), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n7925) );
  INV_X1 U8608 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n11094) );
  XNOR2_X1 U8609 ( .A(n7970), .B(n11092), .ZN(n11880) );
  OAI21_X1 U8610 ( .B1(n11086), .B2(n11067), .A(n11089), .ZN(n7970) );
  NAND2_X1 U8611 ( .A1(n10024), .A2(n7988), .ZN(n7987) );
  XNOR2_X1 U8612 ( .A(n10296), .B(n10294), .ZN(n11412) );
  OAI21_X1 U8613 ( .B1(n7536), .B2(n9761), .A(n9760), .ZN(n10022) );
  OAI21_X1 U8614 ( .B1(n9439), .B2(n9438), .A(n9441), .ZN(n9638) );
  XNOR2_X1 U8615 ( .A(n9439), .B(n9437), .ZN(n10906) );
  NAND2_X1 U8616 ( .A1(n7613), .A2(n7612), .ZN(n9351) );
  NAND2_X1 U8617 ( .A1(n9130), .A2(n9131), .ZN(n7614) );
  XNOR2_X1 U8618 ( .A(n9131), .B(n9129), .ZN(n10261) );
  OR2_X1 U8619 ( .A1(n9089), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n9091) );
  INV_X1 U8620 ( .A(n9031), .ZN(n7965) );
  XNOR2_X1 U8621 ( .A(n15499), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n15500) );
  INV_X1 U8622 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n15532) );
  OAI21_X1 U8623 ( .B1(n15540), .B2(n15539), .A(n7266), .ZN(n7641) );
  NOR2_X1 U8624 ( .A1(n15548), .A2(n15547), .ZN(n15549) );
  OAI21_X1 U8625 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n15585), .A(n15584), .ZN(
        n15593) );
  OR2_X1 U8626 ( .A1(n15632), .A2(n15631), .ZN(n15634) );
  NAND2_X1 U8627 ( .A1(n13480), .A2(n8662), .ZN(n13426) );
  NAND2_X1 U8628 ( .A1(n8659), .A2(n8658), .ZN(n13739) );
  AND2_X1 U8629 ( .A1(n7837), .A2(n7839), .ZN(n11870) );
  AND4_X2 U8630 ( .A1(n8383), .A2(n8382), .A3(n8381), .A4(n8380), .ZN(n10636)
         );
  OR2_X1 U8631 ( .A1(n8556), .A2(n9825), .ZN(n8381) );
  AND4_X1 U8632 ( .A1(n8428), .A2(n8427), .A3(n8426), .A4(n8425), .ZN(n11113)
         );
  INV_X1 U8633 ( .A(n7850), .ZN(n7849) );
  AOI21_X1 U8634 ( .B1(n7850), .B2(n7853), .A(n7848), .ZN(n7847) );
  INV_X1 U8635 ( .A(n13433), .ZN(n7848) );
  NAND2_X1 U8636 ( .A1(n7846), .A2(n7850), .ZN(n13434) );
  NAND2_X1 U8637 ( .A1(n13472), .A2(n7852), .ZN(n7846) );
  AND4_X1 U8638 ( .A1(n8462), .A2(n8461), .A3(n8460), .A4(n8459), .ZN(n11469)
         );
  OR2_X1 U8639 ( .A1(n10166), .A2(n10167), .ZN(n7813) );
  AOI22_X1 U8640 ( .A1(n8973), .A2(n8972), .B1(n8501), .B2(n13568), .ZN(n11951) );
  AND2_X1 U8641 ( .A1(n8681), .A2(n8680), .ZN(n13738) );
  NAND2_X1 U8642 ( .A1(n8555), .A2(n8554), .ZN(n13847) );
  AND3_X1 U8643 ( .A1(n8437), .A2(n8436), .A3(n8435), .ZN(n11116) );
  NAND2_X1 U8644 ( .A1(n7842), .A2(n7844), .ZN(n11604) );
  AND4_X2 U8645 ( .A1(n8400), .A2(n8399), .A3(n8398), .A4(n8397), .ZN(n9769)
         );
  OR2_X1 U8646 ( .A1(n8556), .A2(n9818), .ZN(n8398) );
  NAND2_X1 U8647 ( .A1(n7815), .A2(n8655), .ZN(n13507) );
  AND2_X1 U8648 ( .A1(n7813), .A2(n8411), .ZN(n10395) );
  NAND2_X1 U8649 ( .A1(n7855), .A2(n8582), .ZN(n13516) );
  NAND2_X1 U8650 ( .A1(n7855), .A2(n7852), .ZN(n13517) );
  NAND2_X1 U8651 ( .A1(n7823), .A2(n7326), .ZN(n11204) );
  INV_X1 U8652 ( .A(n7824), .ZN(n7823) );
  OAI21_X1 U8653 ( .B1(n10633), .B2(n11110), .A(n11109), .ZN(n7824) );
  OAI21_X1 U8654 ( .B1(n7829), .B2(n7827), .A(n7825), .ZN(n11205) );
  AND2_X1 U8655 ( .A1(n7826), .A2(n7831), .ZN(n7825) );
  NAND2_X1 U8656 ( .A1(n11110), .A2(n11109), .ZN(n7826) );
  NAND2_X1 U8657 ( .A1(n13525), .A2(n13526), .ZN(n13524) );
  OR2_X1 U8658 ( .A1(n12597), .A2(n12595), .ZN(n12630) );
  INV_X1 U8659 ( .A(n13555), .ZN(n13960) );
  INV_X1 U8660 ( .A(n13678), .ZN(n13698) );
  NAND2_X1 U8661 ( .A1(n8713), .A2(n8712), .ZN(n13557) );
  NAND2_X1 U8662 ( .A1(n8699), .A2(n8698), .ZN(n13725) );
  INV_X1 U8663 ( .A(n13824), .ZN(n13563) );
  INV_X1 U8664 ( .A(n11961), .ZN(n13568) );
  INV_X1 U8665 ( .A(n11469), .ZN(n13572) );
  NAND4_X1 U8666 ( .A1(n8409), .A2(n8408), .A3(n8407), .A4(n8406), .ZN(n13578)
         );
  NAND2_X1 U8667 ( .A1(n9920), .A2(n15655), .ZN(n9947) );
  NAND2_X1 U8668 ( .A1(n7896), .A2(n9794), .ZN(n9854) );
  NAND2_X1 U8669 ( .A1(n9838), .A2(n9865), .ZN(n9867) );
  INV_X1 U8670 ( .A(n7903), .ZN(n10187) );
  INV_X1 U8671 ( .A(n7662), .ZN(n15661) );
  INV_X1 U8672 ( .A(n10774), .ZN(n7661) );
  INV_X1 U8673 ( .A(n7900), .ZN(n11327) );
  INV_X1 U8674 ( .A(n7588), .ZN(n11333) );
  INV_X1 U8675 ( .A(n7898), .ZN(n13627) );
  NOR2_X1 U8676 ( .A1(n15678), .A2(n11310), .ZN(n11313) );
  XNOR2_X1 U8677 ( .A(n13612), .B(n15697), .ZN(n15694) );
  INV_X1 U8678 ( .A(n7679), .ZN(n15693) );
  INV_X1 U8679 ( .A(n15709), .ZN(n7357) );
  INV_X1 U8680 ( .A(n7358), .ZN(n15710) );
  XNOR2_X1 U8681 ( .A(n13615), .B(n15739), .ZN(n15727) );
  INV_X1 U8682 ( .A(n7379), .ZN(n13617) );
  INV_X1 U8683 ( .A(n7665), .ZN(n15784) );
  NOR2_X1 U8684 ( .A1(n15777), .A2(n13637), .ZN(n15797) );
  INV_X1 U8685 ( .A(n7582), .ZN(n15818) );
  OAI21_X1 U8686 ( .B1(n8906), .B2(n13874), .A(n8905), .ZN(n12197) );
  NAND2_X1 U8687 ( .A1(n13676), .A2(n7407), .ZN(n8897) );
  AND2_X1 U8688 ( .A1(n7766), .A2(n7765), .ZN(n13683) );
  NAND2_X1 U8689 ( .A1(n8862), .A2(n8861), .ZN(n13691) );
  INV_X1 U8690 ( .A(n8860), .ZN(n8861) );
  OAI21_X1 U8691 ( .B1(n8859), .B2(n13874), .A(n8858), .ZN(n8860) );
  NAND2_X1 U8692 ( .A1(n8111), .A2(n8845), .ZN(n13768) );
  NAND2_X1 U8693 ( .A1(n8841), .A2(n8840), .ZN(n13809) );
  NAND2_X1 U8694 ( .A1(n13825), .A2(n12730), .ZN(n13813) );
  NAND2_X1 U8695 ( .A1(n7750), .A2(n7751), .ZN(n13855) );
  OR2_X1 U8696 ( .A1(n7362), .A2(n7754), .ZN(n7750) );
  NAND2_X1 U8697 ( .A1(n7362), .A2(n12704), .ZN(n13879) );
  NAND2_X1 U8698 ( .A1(n11695), .A2(n8826), .ZN(n11857) );
  INV_X1 U8699 ( .A(n13868), .ZN(n13887) );
  INV_X1 U8700 ( .A(n8822), .ZN(n16026) );
  AND3_X1 U8701 ( .A1(n8470), .A2(n8469), .A3(n8468), .ZN(n16005) );
  INV_X1 U8702 ( .A(n10528), .ZN(n15893) );
  NAND2_X1 U8703 ( .A1(n8758), .A2(n15893), .ZN(n15892) );
  INV_X1 U8704 ( .A(n15892), .ZN(n13829) );
  INV_X1 U8705 ( .A(n12588), .ZN(n13962) );
  NAND2_X1 U8706 ( .A1(n12586), .A2(n12585), .ZN(n16162) );
  INV_X1 U8707 ( .A(n8909), .ZN(n12199) );
  INV_X1 U8708 ( .A(n12632), .ZN(n13971) );
  INV_X1 U8709 ( .A(n13479), .ZN(n13975) );
  NAND2_X1 U8710 ( .A1(n8575), .A2(n8574), .ZN(n14003) );
  INV_X1 U8711 ( .A(n11030), .ZN(n11061) );
  INV_X1 U8712 ( .A(n8911), .ZN(n14017) );
  INV_X1 U8713 ( .A(n9116), .ZN(n14016) );
  NAND2_X1 U8714 ( .A1(n14021), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7770) );
  NAND2_X1 U8715 ( .A1(n8883), .A2(n8882), .ZN(n12564) );
  INV_X1 U8716 ( .A(n8750), .ZN(n11758) );
  XNOR2_X1 U8717 ( .A(n8302), .B(n8301), .ZN(n11590) );
  XNOR2_X1 U8718 ( .A(n8300), .B(n8299), .ZN(n11452) );
  NAND2_X1 U8719 ( .A1(n8623), .A2(n8275), .ZN(n8638) );
  XNOR2_X1 U8720 ( .A(n8738), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12792) );
  NAND2_X1 U8721 ( .A1(n8308), .A2(n8218), .ZN(n8737) );
  NAND2_X1 U8722 ( .A1(n8273), .A2(n8272), .ZN(n8621) );
  XNOR2_X1 U8723 ( .A(n8316), .B(n8315), .ZN(n12623) );
  INV_X1 U8724 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8315) );
  OAI21_X1 U8725 ( .B1(n8314), .B2(P3_IR_REG_20__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8316) );
  INV_X1 U8726 ( .A(SI_20_), .ZN(n11223) );
  NAND2_X1 U8727 ( .A1(n8314), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8310) );
  INV_X1 U8728 ( .A(SI_19_), .ZN(n15180) );
  NAND2_X1 U8729 ( .A1(n7387), .A2(n8267), .ZN(n8584) );
  NAND2_X1 U8730 ( .A1(n8568), .A2(n8567), .ZN(n7387) );
  INV_X1 U8731 ( .A(SI_18_), .ZN(n15184) );
  INV_X1 U8732 ( .A(SI_16_), .ZN(n15207) );
  NAND2_X1 U8733 ( .A1(n7725), .A2(n8262), .ZN(n8534) );
  NAND2_X1 U8734 ( .A1(n8521), .A2(n8520), .ZN(n7725) );
  NOR2_X1 U8735 ( .A1(n7810), .A2(n8433), .ZN(n8522) );
  INV_X1 U8736 ( .A(SI_14_), .ZN(n15318) );
  INV_X1 U8737 ( .A(SI_13_), .ZN(n15311) );
  XNOR2_X1 U8738 ( .A(n8513), .B(n8512), .ZN(n15711) );
  NAND2_X1 U8739 ( .A1(n7719), .A2(n8258), .ZN(n8510) );
  NAND2_X1 U8740 ( .A1(n8497), .A2(n8257), .ZN(n7719) );
  INV_X1 U8741 ( .A(SI_11_), .ZN(n15208) );
  INV_X1 U8742 ( .A(n11315), .ZN(n11328) );
  OAI21_X1 U8743 ( .B1(n8432), .B2(n7403), .A(n7401), .ZN(n8451) );
  OR2_X1 U8744 ( .A1(n8365), .A2(n8364), .ZN(n10772) );
  NAND2_X1 U8745 ( .A1(n7406), .A2(n8246), .ZN(n8367) );
  NAND2_X1 U8746 ( .A1(n8432), .A2(n8244), .ZN(n7406) );
  XNOR2_X1 U8747 ( .A(n8420), .B(P3_IR_REG_4__SCAN_IN), .ZN(n10151) );
  NOR2_X1 U8748 ( .A1(n8386), .A2(n8221), .ZN(n7687) );
  NAND2_X1 U8749 ( .A1(n8392), .A2(n8237), .ZN(n8385) );
  INV_X1 U8750 ( .A(n8236), .ZN(n8391) );
  INV_X1 U8751 ( .A(n8386), .ZN(n7891) );
  MUX2_X1 U8752 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7893), .S(
        P3_IR_REG_1__SCAN_IN), .Z(n7892) );
  NAND2_X1 U8753 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7893) );
  NAND2_X1 U8754 ( .A1(n11706), .A2(n8044), .ZN(n11839) );
  NAND2_X1 U8755 ( .A1(n14055), .A2(n8016), .ZN(n14054) );
  NAND2_X1 U8756 ( .A1(n8024), .A2(n14062), .ZN(n14127) );
  OR2_X1 U8757 ( .A1(n14145), .A2(n12383), .ZN(n8024) );
  NAND2_X1 U8758 ( .A1(n9997), .A2(n9996), .ZN(n10095) );
  NAND2_X1 U8759 ( .A1(n10095), .A2(n10096), .ZN(n10094) );
  NAND2_X1 U8760 ( .A1(n14054), .A2(n8014), .ZN(n14116) );
  NAND2_X1 U8761 ( .A1(n14145), .A2(n8023), .ZN(n8020) );
  NOR2_X1 U8762 ( .A1(n12392), .A2(n7336), .ZN(n14029) );
  NAND2_X1 U8763 ( .A1(n14178), .A2(n14416), .ZN(n7336) );
  AND2_X1 U8764 ( .A1(n11269), .A2(n11268), .ZN(n8042) );
  NAND2_X1 U8765 ( .A1(n12422), .A2(n7338), .ZN(n14147) );
  OR2_X1 U8766 ( .A1(n12375), .A2(n12376), .ZN(n7338) );
  AOI21_X1 U8767 ( .B1(n10096), .B2(n7557), .A(n7556), .ZN(n7555) );
  INV_X1 U8768 ( .A(n10003), .ZN(n7556) );
  AND2_X1 U8769 ( .A1(n14154), .A2(n14040), .ZN(n7363) );
  NAND2_X1 U8770 ( .A1(n9904), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14161) );
  AND2_X1 U8771 ( .A1(n9597), .A2(n9571), .ZN(n14165) );
  NAND2_X1 U8772 ( .A1(n11839), .A2(n8043), .ZN(n11923) );
  NAND2_X1 U8773 ( .A1(n11537), .A2(n11536), .ZN(n13230) );
  NOR2_X1 U8774 ( .A1(n13348), .A2(n13347), .ZN(n13349) );
  AND2_X1 U8775 ( .A1(n14233), .A2(n13353), .ZN(n13362) );
  OR2_X1 U8776 ( .A1(n9622), .A2(n9601), .ZN(n9605) );
  NAND2_X1 U8777 ( .A1(n14309), .A2(n12361), .ZN(n14293) );
  AND2_X1 U8778 ( .A1(n12296), .A2(n12295), .ZN(n14306) );
  NAND2_X1 U8779 ( .A1(n14334), .A2(n12359), .ZN(n14323) );
  OR2_X1 U8780 ( .A1(n14358), .A2(n7475), .ZN(n7468) );
  NAND2_X1 U8781 ( .A1(n7457), .A2(n12270), .ZN(n14341) );
  NAND2_X1 U8782 ( .A1(n14385), .A2(n12356), .ZN(n14374) );
  OAI21_X1 U8783 ( .B1(n11721), .B2(n7480), .A(n7478), .ZN(n14405) );
  NAND2_X1 U8784 ( .A1(n11805), .A2(n11804), .ZN(n12354) );
  OAI21_X1 U8785 ( .B1(n11184), .B2(n7862), .A(n7860), .ZN(n11545) );
  NAND2_X1 U8786 ( .A1(n11184), .A2(n11183), .ZN(n11510) );
  NAND2_X1 U8787 ( .A1(n10963), .A2(n10557), .ZN(n10686) );
  NAND2_X1 U8788 ( .A1(n7447), .A2(n9976), .ZN(n10113) );
  INV_X1 U8789 ( .A(n10869), .ZN(n10834) );
  INV_X1 U8790 ( .A(n14366), .ZN(n14434) );
  INV_X1 U8791 ( .A(n14303), .ZN(n14436) );
  INV_X1 U8792 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n7461) );
  NAND2_X1 U8793 ( .A1(n12246), .A2(n12245), .ZN(n14502) );
  AND2_X2 U8794 ( .A1(n10136), .A2(n9994), .ZN(n16142) );
  INV_X1 U8795 ( .A(n14232), .ZN(n14540) );
  NAND2_X1 U8796 ( .A1(n14461), .A2(n7246), .ZN(n14545) );
  INV_X2 U8797 ( .A(n14277), .ZN(n14551) );
  INV_X1 U8798 ( .A(n14502), .ZN(n14567) );
  INV_X1 U8799 ( .A(n13230), .ZN(n11837) );
  AND2_X1 U8800 ( .A1(n9902), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15409) );
  INV_X1 U8801 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n7869) );
  MUX2_X1 U8802 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9574), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n9576) );
  INV_X1 U8803 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8931) );
  INV_X1 U8804 ( .A(n9546), .ZN(n14599) );
  INV_X1 U8805 ( .A(n9547), .ZN(n14602) );
  INV_X1 U8806 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n9474) );
  INV_X1 U8807 ( .A(n7182), .ZN(n13405) );
  INV_X1 U8808 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10592) );
  INV_X1 U8809 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n11489) );
  INV_X1 U8810 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9851) );
  INV_X1 U8811 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9137) );
  INV_X1 U8812 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9110) );
  INV_X1 U8813 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9006) );
  NAND2_X1 U8814 ( .A1(n16121), .A2(n12432), .ZN(n16124) );
  NAND2_X1 U8815 ( .A1(n11295), .A2(n7364), .ZN(n11300) );
  NAND2_X1 U8816 ( .A1(n11294), .A2(n7365), .ZN(n7364) );
  INV_X1 U8817 ( .A(n11296), .ZN(n7365) );
  OAI21_X1 U8818 ( .B1(n8059), .B2(n8064), .A(n8055), .ZN(n8054) );
  NAND2_X1 U8819 ( .A1(n8059), .A2(n8056), .ZN(n8055) );
  NAND2_X1 U8820 ( .A1(n12530), .A2(n8057), .ZN(n8056) );
  INV_X1 U8821 ( .A(n8061), .ZN(n8057) );
  NAND2_X1 U8822 ( .A1(n8059), .A2(n12530), .ZN(n8058) );
  NAND2_X1 U8823 ( .A1(n10819), .A2(n10818), .ZN(n10820) );
  OAI21_X1 U8824 ( .B1(n14621), .B2(n8076), .A(n8073), .ZN(n14630) );
  NAND2_X1 U8825 ( .A1(n8085), .A2(n7229), .ZN(n11927) );
  AND2_X1 U8826 ( .A1(n8085), .A2(n8084), .ZN(n11820) );
  INV_X1 U8827 ( .A(n14899), .ZN(n14859) );
  AOI21_X1 U8828 ( .B1(n8068), .B2(n8070), .A(n7250), .ZN(n8066) );
  NAND2_X1 U8829 ( .A1(n14648), .A2(n8081), .ZN(n14662) );
  NAND2_X1 U8830 ( .A1(n8067), .A2(n12492), .ZN(n14672) );
  NAND2_X1 U8831 ( .A1(n14613), .A2(n14614), .ZN(n8067) );
  NAND2_X1 U8832 ( .A1(n8093), .A2(n8089), .ZN(n11295) );
  AND2_X1 U8833 ( .A1(n11127), .A2(n8092), .ZN(n8089) );
  AND2_X1 U8834 ( .A1(n8093), .A2(n8092), .ZN(n11128) );
  AND2_X1 U8835 ( .A1(n12023), .A2(n12022), .ZN(n14976) );
  NAND2_X1 U8836 ( .A1(n14680), .A2(n12468), .ZN(n14681) );
  AND2_X1 U8837 ( .A1(n12039), .A2(n12027), .ZN(n14982) );
  NAND2_X1 U8838 ( .A1(n11933), .A2(n11932), .ZN(n16121) );
  NAND2_X1 U8839 ( .A1(n11477), .A2(n8086), .ZN(n11480) );
  AOI21_X1 U8840 ( .B1(n10053), .B2(P2_DATAO_REG_2__SCAN_IN), .A(n7590), .ZN(
        n7589) );
  NOR2_X1 U8841 ( .A1(n12049), .A2(n14781), .ZN(n7590) );
  NAND2_X1 U8842 ( .A1(n8080), .A2(n8079), .ZN(n14702) );
  INV_X1 U8843 ( .A(n16123), .ZN(n14719) );
  INV_X1 U8844 ( .A(n16133), .ZN(n14728) );
  NAND2_X1 U8845 ( .A1(n12058), .A2(n12057), .ZN(n14961) );
  INV_X1 U8846 ( .A(n9416), .ZN(n14753) );
  AND2_X1 U8847 ( .A1(n10302), .A2(n10028), .ZN(n11413) );
  INV_X1 U8848 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7623) );
  NAND2_X1 U8849 ( .A1(n13013), .A2(n13012), .ZN(n15024) );
  INV_X1 U8850 ( .A(n15040), .ZN(n12555) );
  NAND2_X1 U8851 ( .A1(n14865), .A2(n7997), .ZN(n12163) );
  AOI21_X1 U8852 ( .B1(n12152), .B2(n15955), .A(n12151), .ZN(n15044) );
  NAND2_X1 U8853 ( .A1(n14912), .A2(n7717), .ZN(n14893) );
  NAND2_X1 U8854 ( .A1(n14929), .A2(n12071), .ZN(n14917) );
  AND2_X1 U8855 ( .A1(n7421), .A2(n7228), .ZN(n14945) );
  NAND2_X1 U8856 ( .A1(n14959), .A2(n14966), .ZN(n7421) );
  OAI21_X1 U8857 ( .B1(n7977), .B2(n7707), .A(n7705), .ZN(n14965) );
  INV_X1 U8858 ( .A(n14976), .ZN(n15086) );
  NAND2_X1 U8859 ( .A1(n7974), .A2(n7978), .ZN(n14973) );
  NAND2_X1 U8860 ( .A1(n7977), .A2(n7975), .ZN(n7974) );
  NAND2_X1 U8861 ( .A1(n7977), .A2(n12156), .ZN(n14989) );
  NAND2_X1 U8862 ( .A1(n15007), .A2(n12007), .ZN(n14988) );
  NAND2_X1 U8863 ( .A1(n7960), .A2(n7961), .ZN(n11901) );
  OR2_X1 U8864 ( .A1(n11625), .A2(n13048), .ZN(n7960) );
  INV_X1 U8865 ( .A(n15122), .ZN(n14732) );
  NAND2_X1 U8866 ( .A1(n11625), .A2(n11624), .ZN(n11650) );
  NAND2_X1 U8867 ( .A1(n7712), .A2(n11442), .ZN(n11443) );
  NAND2_X1 U8868 ( .A1(n11453), .A2(n13043), .ZN(n7712) );
  NAND2_X1 U8869 ( .A1(n11038), .A2(n11037), .ZN(n12869) );
  NAND2_X1 U8870 ( .A1(n7437), .A2(n11011), .ZN(n11013) );
  NAND2_X1 U8871 ( .A1(n10996), .A2(n10995), .ZN(n11001) );
  NAND2_X1 U8872 ( .A1(n7963), .A2(n10922), .ZN(n11010) );
  NOR2_X1 U8873 ( .A1(n7697), .A2(n7699), .ZN(n10910) );
  INV_X1 U8874 ( .A(n10904), .ZN(n7699) );
  INV_X1 U8875 ( .A(n10905), .ZN(n7697) );
  INV_X1 U8876 ( .A(n15977), .ZN(n16034) );
  NAND2_X1 U8877 ( .A1(n10471), .A2(n10470), .ZN(n10477) );
  NAND2_X1 U8878 ( .A1(n10282), .A2(n13032), .ZN(n10492) );
  INV_X1 U8879 ( .A(n14997), .ZN(n16035) );
  NAND2_X1 U8880 ( .A1(n7941), .A2(n10277), .ZN(n15956) );
  INV_X1 U8881 ( .A(n13029), .ZN(n10277) );
  NAND2_X1 U8882 ( .A1(n11899), .A2(n11009), .ZN(n14967) );
  INV_X1 U8883 ( .A(n16037), .ZN(n15016) );
  INV_X1 U8884 ( .A(n10755), .ZN(n16044) );
  AND2_X2 U8885 ( .A1(n10289), .A2(n10534), .ZN(n16067) );
  INV_X1 U8886 ( .A(n15049), .ZN(n7430) );
  OR2_X1 U8887 ( .A1(n15054), .A2(n15933), .ZN(n7345) );
  NAND2_X1 U8888 ( .A1(n13006), .A2(n12190), .ZN(n13318) );
  NOR2_X1 U8889 ( .A1(n8956), .A2(n8955), .ZN(n8957) );
  XNOR2_X1 U8890 ( .A(n12048), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15169) );
  INV_X1 U8891 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10895) );
  INV_X1 U8892 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10304) );
  INV_X1 U8893 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9768) );
  INV_X1 U8894 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9443) );
  INV_X1 U8895 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9360) );
  INV_X1 U8896 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9180) );
  INV_X1 U8897 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9114) );
  INV_X1 U8898 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9038) );
  INV_X1 U8899 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U8900 ( .A1(n7342), .A2(n15492), .ZN(n15494) );
  XNOR2_X1 U8901 ( .A(n15516), .B(n7647), .ZN(n15518) );
  INV_X1 U8902 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7647) );
  NOR2_X1 U8903 ( .A1(n15509), .A2(n15510), .ZN(n15517) );
  XNOR2_X1 U8904 ( .A(n15520), .B(n7645), .ZN(n15522) );
  INV_X1 U8905 ( .A(n15521), .ZN(n7645) );
  AND2_X1 U8906 ( .A1(n15542), .A2(n15541), .ZN(n15544) );
  AOI21_X1 U8907 ( .B1(n7654), .B2(n7649), .A(n7280), .ZN(n15571) );
  AND2_X1 U8908 ( .A1(n15558), .A2(n7650), .ZN(n7649) );
  INV_X1 U8909 ( .A(n7652), .ZN(n7648) );
  NOR2_X1 U8910 ( .A1(n15581), .A2(n15580), .ZN(n15589) );
  OAI21_X1 U8911 ( .B1(n15624), .B2(n15623), .A(n15622), .ZN(n15626) );
  OAI21_X1 U8912 ( .B1(n13898), .B2(n13554), .A(n8782), .ZN(n8783) );
  AOI21_X1 U8913 ( .B1(n7578), .B2(n10162), .A(n7575), .ZN(n13648) );
  NAND2_X1 U8914 ( .A1(n15802), .A2(n7331), .ZN(n7355) );
  NOR2_X1 U8915 ( .A1(n13669), .A2(n7909), .ZN(n7908) );
  OR2_X1 U8916 ( .A1(n7666), .A2(n15802), .ZN(n7669) );
  NAND2_X1 U8917 ( .A1(n9876), .A2(n9875), .ZN(n10031) );
  NAND2_X1 U8918 ( .A1(n8030), .A2(n8034), .ZN(n9899) );
  OAI211_X1 U8919 ( .C1(n14456), .C2(n14303), .A(n7888), .B(n7887), .ZN(
        P2_U3236) );
  AOI21_X1 U8920 ( .B1(n14452), .B2(n14438), .A(n12367), .ZN(n7887) );
  NAND2_X1 U8921 ( .A1(n7889), .A2(n14427), .ZN(n7888) );
  NAND2_X1 U8922 ( .A1(n14233), .A2(n14524), .ZN(n7339) );
  NAND2_X1 U8923 ( .A1(n14542), .A2(n16142), .ZN(n7530) );
  NAND2_X1 U8924 ( .A1(n7462), .A2(n7459), .ZN(P2_U3526) );
  AOI21_X1 U8925 ( .B1(n14463), .B2(n14524), .A(n7460), .ZN(n7459) );
  NAND2_X1 U8926 ( .A1(n14545), .A2(n16142), .ZN(n7462) );
  NOR2_X1 U8927 ( .A1(n16142), .A2(n7461), .ZN(n7460) );
  NAND2_X1 U8928 ( .A1(n14233), .A2(n14578), .ZN(n7340) );
  OAI21_X1 U8929 ( .B1(n14542), .B2(n16143), .A(n7494), .ZN(P2_U3495) );
  INV_X1 U8930 ( .A(n7495), .ZN(n7494) );
  OAI22_X1 U8931 ( .A1(n14544), .A2(n14566), .B1(n16146), .B2(n14543), .ZN(
        n7495) );
  XNOR2_X1 U8932 ( .A(n7367), .B(n7366), .ZN(n14612) );
  AND3_X1 U8933 ( .A1(n13074), .A2(n13073), .A3(n8179), .ZN(n13079) );
  OR2_X1 U8934 ( .A1(n16067), .A2(n7968), .ZN(n7967) );
  NAND2_X1 U8935 ( .A1(n15128), .A2(n16067), .ZN(n7969) );
  INV_X1 U8936 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7968) );
  NAND2_X1 U8937 ( .A1(n7429), .A2(n7427), .ZN(P1_U3555) );
  OR2_X1 U8938 ( .A1(n16067), .A2(n7428), .ZN(n7427) );
  NAND2_X1 U8939 ( .A1(n15130), .A2(n16067), .ZN(n7429) );
  INV_X1 U8940 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n7428) );
  INV_X1 U8941 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7622) );
  NOR2_X1 U8942 ( .A1(n15566), .A2(n15565), .ZN(n15567) );
  XNOR2_X1 U8943 ( .A(n15644), .B(n7656), .ZN(n7655) );
  NAND2_X1 U8944 ( .A1(n15641), .A2(n15642), .ZN(n7657) );
  XNOR2_X1 U8945 ( .A(n15643), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n7656) );
  OR2_X1 U8946 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .ZN(
        n7189) );
  NOR2_X1 U8947 ( .A1(n8046), .A2(n7182), .ZN(n7190) );
  NOR2_X1 U8948 ( .A1(n13631), .A2(n9254), .ZN(n7191) );
  INV_X1 U8949 ( .A(n8438), .ZN(n8605) );
  INV_X1 U8950 ( .A(n14966), .ZN(n7702) );
  INV_X1 U8951 ( .A(n13043), .ZN(n7709) );
  INV_X1 U8952 ( .A(n8896), .ZN(n7408) );
  AND2_X1 U8953 ( .A1(n7809), .A2(n13752), .ZN(n7192) );
  OR2_X1 U8954 ( .A1(n15097), .A2(n14979), .ZN(n7193) );
  AND2_X1 U8955 ( .A1(n7886), .A2(n11804), .ZN(n7194) );
  OR2_X1 U8956 ( .A1(n15557), .A2(n15556), .ZN(n7195) );
  NOR2_X1 U8957 ( .A1(n10434), .A2(n7986), .ZN(n7985) );
  INV_X1 U8958 ( .A(n11075), .ZN(n8117) );
  AND2_X1 U8959 ( .A1(n8021), .A2(n12389), .ZN(n7196) );
  AND2_X1 U8960 ( .A1(n7279), .A2(n7490), .ZN(n7197) );
  AND2_X1 U8961 ( .A1(n13309), .A2(n13308), .ZN(n7198) );
  INV_X1 U8962 ( .A(n12615), .ZN(n13781) );
  AND2_X1 U8963 ( .A1(n12763), .A2(n12764), .ZN(n12760) );
  AND3_X1 U8964 ( .A1(n12883), .A2(n7298), .A3(n12882), .ZN(n7199) );
  AND2_X1 U8965 ( .A1(n8018), .A2(n8017), .ZN(n7200) );
  OR2_X1 U8966 ( .A1(n12869), .A2(n11476), .ZN(n7201) );
  NOR2_X1 U8967 ( .A1(n11922), .A2(n7564), .ZN(n7563) );
  AND2_X1 U8968 ( .A1(n7929), .A2(n12889), .ZN(n7202) );
  AND2_X1 U8969 ( .A1(n8644), .A2(n8647), .ZN(n7203) );
  OR2_X1 U8970 ( .A1(n7923), .A2(n7924), .ZN(n7204) );
  NAND2_X1 U8971 ( .A1(n10185), .A2(n10189), .ZN(n7205) );
  AND2_X1 U8972 ( .A1(n14871), .A2(n7998), .ZN(n7206) );
  AND2_X1 U8973 ( .A1(n8655), .A2(n13771), .ZN(n7207) );
  INV_X1 U8974 ( .A(n14233), .ZN(n14536) );
  MUX2_X1 U8975 ( .A(n14899), .B(n15051), .S(n13015), .Z(n12969) );
  INV_X1 U8976 ( .A(n12969), .ZN(n12970) );
  INV_X1 U8977 ( .A(n8849), .ZN(n7416) );
  AND2_X1 U8978 ( .A1(n8482), .A2(n11693), .ZN(n7208) );
  NAND2_X1 U8979 ( .A1(n15565), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7650) );
  INV_X1 U8980 ( .A(n14178), .ZN(n14355) );
  AND2_X1 U8981 ( .A1(n13631), .A2(n9254), .ZN(n7209) );
  AOI21_X1 U8982 ( .B1(n7191), .B2(n15720), .A(n7209), .ZN(n7569) );
  INV_X1 U8983 ( .A(n12844), .ZN(n7595) );
  INV_X1 U8984 ( .A(n13177), .ZN(n7681) );
  NAND2_X1 U8985 ( .A1(n7594), .A2(n7593), .ZN(n10926) );
  INV_X1 U8986 ( .A(n9339), .ZN(n11659) );
  INV_X1 U8987 ( .A(n14262), .ZN(n7793) );
  INV_X1 U8988 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n14582) );
  OR2_X1 U8989 ( .A1(n8298), .A2(n8121), .ZN(n7211) );
  NAND2_X1 U8990 ( .A1(n15002), .A2(n12155), .ZN(n7977) );
  AND2_X1 U8991 ( .A1(n8011), .A2(n8012), .ZN(n7212) );
  AND2_X1 U8992 ( .A1(n15013), .A2(n7608), .ZN(n7213) );
  OR2_X1 U8993 ( .A1(n13515), .A2(n7854), .ZN(n7853) );
  INV_X1 U8994 ( .A(n13050), .ZN(n12021) );
  INV_X1 U8995 ( .A(n12530), .ZN(n8064) );
  AND2_X1 U8996 ( .A1(n13281), .A2(n13280), .ZN(n7214) );
  OR3_X2 U8997 ( .A1(n13404), .A2(n13403), .A3(n13402), .ZN(n7215) );
  NAND2_X1 U8998 ( .A1(n8413), .A2(n10636), .ZN(n7216) );
  AND2_X1 U8999 ( .A1(n12972), .A2(n12971), .ZN(n7217) );
  AND2_X1 U9000 ( .A1(n9000), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7218) );
  NOR2_X1 U9001 ( .A1(n11847), .A2(n11846), .ZN(n7219) );
  OR2_X1 U9002 ( .A1(n14326), .A2(n14475), .ZN(n7220) );
  AND2_X1 U9003 ( .A1(n8633), .A2(n8645), .ZN(n7221) );
  INV_X1 U9004 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n15488) );
  OR2_X1 U9005 ( .A1(n13094), .A2(n8896), .ZN(n8881) );
  AND3_X1 U9006 ( .A1(n13369), .A2(n13370), .A3(n7441), .ZN(n7222) );
  XNOR2_X1 U9007 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n8450) );
  AND2_X1 U9008 ( .A1(n7358), .A2(n7357), .ZN(n7223) );
  INV_X1 U9009 ( .A(n13032), .ZN(n7947) );
  INV_X1 U9010 ( .A(n15075), .ZN(n7611) );
  OR2_X1 U9011 ( .A1(n8851), .A2(n13710), .ZN(n7224) );
  AND2_X1 U9012 ( .A1(n14117), .A2(n8016), .ZN(n7225) );
  OAI21_X1 U9013 ( .B1(n15777), .B2(n7572), .A(n7571), .ZN(n13640) );
  INV_X1 U9014 ( .A(n13640), .ZN(n7574) );
  AND4_X1 U9015 ( .A1(n8005), .A2(n13056), .A3(n14862), .A4(n13055), .ZN(n7226) );
  NOR2_X1 U9016 ( .A1(n8181), .A2(n13835), .ZN(n7227) );
  OR2_X1 U9017 ( .A1(n15082), .A2(n12914), .ZN(n7228) );
  INV_X1 U9018 ( .A(n9615), .ZN(n7434) );
  AND2_X1 U9019 ( .A1(n11819), .A2(n8084), .ZN(n7229) );
  AND2_X1 U9020 ( .A1(n14435), .A2(n14191), .ZN(n7230) );
  AND2_X1 U9021 ( .A1(n8806), .A2(n12753), .ZN(n7231) );
  INV_X1 U9022 ( .A(n15028), .ZN(n14851) );
  OAI21_X1 U9023 ( .B1(n13318), .B2(n12994), .A(n12995), .ZN(n15028) );
  AND3_X1 U9024 ( .A1(n8938), .A2(n9036), .A3(n8946), .ZN(n7232) );
  NAND2_X1 U9025 ( .A1(n12538), .A2(n12537), .ZN(n15031) );
  INV_X1 U9026 ( .A(n15031), .ZN(n7603) );
  INV_X1 U9027 ( .A(n13038), .ZN(n11014) );
  AND2_X1 U9028 ( .A1(n16128), .A2(n14739), .ZN(n7233) );
  AND2_X1 U9029 ( .A1(n15057), .A2(n14881), .ZN(n7234) );
  AND2_X1 U9030 ( .A1(n14656), .A2(n14664), .ZN(n7235) );
  AND2_X1 U9031 ( .A1(n12010), .A2(n12009), .ZN(n15097) );
  AND2_X1 U9032 ( .A1(n7707), .A2(n7702), .ZN(n7236) );
  INV_X1 U9033 ( .A(n14463), .ZN(n7375) );
  NOR2_X1 U9034 ( .A1(n14045), .A2(n8037), .ZN(n7237) );
  INV_X1 U9035 ( .A(n15006), .ZN(n14979) );
  AND2_X1 U9036 ( .A1(n12020), .A2(n12019), .ZN(n15006) );
  OR2_X1 U9037 ( .A1(n15697), .A2(n13612), .ZN(n7238) );
  NOR2_X1 U9038 ( .A1(n15797), .A2(n15796), .ZN(n7239) );
  AND2_X1 U9039 ( .A1(n8111), .A2(n8109), .ZN(n7241) );
  AND2_X1 U9040 ( .A1(n14249), .A2(n14248), .ZN(n7242) );
  AND2_X1 U9041 ( .A1(n7391), .A2(n7718), .ZN(n7243) );
  AND2_X1 U9042 ( .A1(n8117), .A2(n8816), .ZN(n7244) );
  OR2_X1 U9043 ( .A1(n13220), .A2(n13219), .ZN(n7245) );
  INV_X1 U9044 ( .A(n10886), .ZN(n7636) );
  AND2_X1 U9045 ( .A1(n14462), .A2(n14460), .ZN(n7246) );
  INV_X1 U9046 ( .A(n10186), .ZN(n7902) );
  INV_X1 U9047 ( .A(n7721), .ZN(n7720) );
  OAI21_X1 U9048 ( .B1(n8257), .B2(n7722), .A(n8509), .ZN(n7721) );
  OR2_X1 U9049 ( .A1(n13255), .A2(n13256), .ZN(n7247) );
  AND2_X1 U9050 ( .A1(n12458), .A2(n8079), .ZN(n7248) );
  AND2_X1 U9051 ( .A1(n7974), .A2(n7972), .ZN(n7249) );
  AND2_X1 U9052 ( .A1(n12498), .A2(n12497), .ZN(n7250) );
  AND2_X1 U9053 ( .A1(n14309), .A2(n7874), .ZN(n7251) );
  INV_X1 U9054 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7344) );
  INV_X1 U9055 ( .A(n7904), .ZN(n13644) );
  NAND2_X1 U9056 ( .A1(n7574), .A2(n13641), .ZN(n7904) );
  AND2_X1 U9057 ( .A1(n12522), .A2(n12521), .ZN(n7252) );
  OR2_X1 U9058 ( .A1(n8754), .A2(P3_IR_REG_24__SCAN_IN), .ZN(n7253) );
  AND2_X1 U9059 ( .A1(n12478), .A2(n12477), .ZN(n7254) );
  NOR2_X1 U9060 ( .A1(n13704), .A2(n13712), .ZN(n7255) );
  AND2_X1 U9061 ( .A1(n12869), .A2(n11476), .ZN(n7256) );
  NOR2_X1 U9062 ( .A1(n14577), .A2(n14183), .ZN(n7257) );
  NOR2_X1 U9063 ( .A1(n12435), .A2(n12434), .ZN(n7258) );
  NOR2_X1 U9064 ( .A1(n15075), .A2(n14961), .ZN(n7259) );
  NOR2_X1 U9065 ( .A1(n14577), .A2(n12227), .ZN(n7260) );
  NOR2_X1 U9066 ( .A1(n14502), .A2(n14180), .ZN(n7261) );
  NOR2_X1 U9067 ( .A1(n15122), .A2(n16116), .ZN(n7262) );
  NOR2_X1 U9068 ( .A1(n8805), .A2(n13765), .ZN(n7263) );
  NOR2_X1 U9069 ( .A1(n13772), .A2(n13560), .ZN(n7264) );
  OR2_X1 U9070 ( .A1(n15991), .A2(n10491), .ZN(n7265) );
  OR2_X1 U9071 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n15538), .ZN(n7266) );
  AND2_X1 U9072 ( .A1(n7929), .A2(n12891), .ZN(n7267) );
  AND2_X1 U9073 ( .A1(n7468), .A2(n7473), .ZN(n7268) );
  AND2_X1 U9074 ( .A1(n13568), .A2(n8828), .ZN(n7269) );
  AND2_X1 U9075 ( .A1(n12390), .A2(n8027), .ZN(n7270) );
  AND2_X1 U9076 ( .A1(n11014), .A2(n7694), .ZN(n7271) );
  AND2_X1 U9077 ( .A1(n7210), .A2(n12159), .ZN(n7272) );
  AND2_X1 U9078 ( .A1(n9175), .A2(SI_7_), .ZN(n7273) );
  AND2_X1 U9079 ( .A1(n12962), .A2(n12961), .ZN(n7274) );
  AND2_X1 U9080 ( .A1(n7634), .A2(n7538), .ZN(n7275) );
  INV_X1 U9081 ( .A(n7985), .ZN(n7984) );
  NOR2_X1 U9082 ( .A1(n7930), .A2(n12861), .ZN(n7502) );
  OR2_X1 U9083 ( .A1(n12862), .A2(n12859), .ZN(n7276) );
  INV_X1 U9084 ( .A(n7829), .ZN(n7828) );
  NAND2_X1 U9085 ( .A1(n7832), .A2(n7830), .ZN(n7829) );
  INV_X1 U9086 ( .A(n13094), .ZN(n13966) );
  NAND2_X1 U9087 ( .A1(n8879), .A2(n8878), .ZN(n13094) );
  OR2_X1 U9088 ( .A1(n8165), .A2(n13316), .ZN(n7277) );
  AND2_X1 U9089 ( .A1(n8130), .A2(n8129), .ZN(n7278) );
  INV_X1 U9090 ( .A(n13242), .ZN(n8138) );
  INV_X1 U9091 ( .A(n7877), .ZN(n7475) );
  AND2_X1 U9092 ( .A1(n13395), .A2(n12357), .ZN(n7877) );
  NAND2_X1 U9093 ( .A1(n13287), .A2(n13288), .ZN(n7279) );
  OR2_X1 U9094 ( .A1(n7653), .A2(n7648), .ZN(n7280) );
  NAND2_X1 U9095 ( .A1(n7219), .A2(n7561), .ZN(n7281) );
  OR2_X1 U9096 ( .A1(n13050), .A2(n7956), .ZN(n7282) );
  OR2_X1 U9097 ( .A1(n13339), .A2(n13338), .ZN(n7283) );
  INV_X1 U9098 ( .A(n13000), .ZN(n7936) );
  AND2_X1 U9099 ( .A1(n12687), .A2(n12682), .ZN(n7284) );
  AND2_X1 U9100 ( .A1(n7401), .A2(n8450), .ZN(n7285) );
  AND2_X1 U9101 ( .A1(n8106), .A2(n8105), .ZN(n7286) );
  AND2_X1 U9102 ( .A1(n9072), .A2(n9066), .ZN(n7287) );
  INV_X1 U9103 ( .A(n13171), .ZN(n8150) );
  NOR2_X1 U9104 ( .A1(n11605), .A2(n7841), .ZN(n7840) );
  AND2_X1 U9105 ( .A1(n12731), .A2(n12730), .ZN(n7288) );
  AND2_X1 U9106 ( .A1(n8655), .A2(n7816), .ZN(n7289) );
  OR2_X1 U9107 ( .A1(n8754), .A2(n8120), .ZN(n7290) );
  AND2_X1 U9108 ( .A1(n11980), .A2(n8008), .ZN(n7291) );
  AND2_X1 U9109 ( .A1(n10476), .A2(n10470), .ZN(n7292) );
  AND2_X1 U9110 ( .A1(n7359), .A2(n14866), .ZN(n7293) );
  AND2_X1 U9111 ( .A1(n14912), .A2(n12160), .ZN(n7294) );
  AND2_X1 U9112 ( .A1(n8064), .A2(n8061), .ZN(n7295) );
  OR2_X1 U9113 ( .A1(n12833), .A2(n12835), .ZN(n7296) );
  INV_X1 U9114 ( .A(n12760), .ZN(n13740) );
  OR2_X1 U9115 ( .A1(n12906), .A2(n12904), .ZN(n7297) );
  OR2_X1 U9116 ( .A1(n12888), .A2(n12886), .ZN(n7298) );
  AND2_X1 U9117 ( .A1(n8926), .A2(n7551), .ZN(n7299) );
  INV_X1 U9118 ( .A(n10743), .ZN(n7944) );
  NAND2_X1 U9119 ( .A1(n7936), .A2(n13001), .ZN(n7300) );
  NAND2_X1 U9120 ( .A1(n13204), .A2(n13205), .ZN(n7301) );
  NAND2_X1 U9121 ( .A1(n13271), .A2(n13272), .ZN(n7302) );
  AND2_X1 U9122 ( .A1(n7287), .A2(n9068), .ZN(n7303) );
  NAND2_X1 U9123 ( .A1(n13256), .A2(n13255), .ZN(n7304) );
  OR2_X1 U9124 ( .A1(n13312), .A2(n7198), .ZN(n7305) );
  INV_X1 U9125 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7952) );
  NAND2_X1 U9126 ( .A1(n12977), .A2(n7521), .ZN(n7306) );
  INV_X1 U9127 ( .A(n14408), .ZN(n7801) );
  INV_X1 U9128 ( .A(n15010), .ZN(n7955) );
  NAND2_X1 U9129 ( .A1(n13567), .A2(n11968), .ZN(n7307) );
  INV_X1 U9130 ( .A(n13613), .ZN(n15697) );
  INV_X1 U9131 ( .A(n14475), .ZN(n7691) );
  AND2_X1 U9132 ( .A1(n11839), .A2(n7563), .ZN(n7308) );
  AND2_X1 U9133 ( .A1(n8020), .A2(n8021), .ZN(n7309) );
  OR2_X1 U9134 ( .A1(n13470), .A2(n13843), .ZN(n7310) );
  AND2_X1 U9135 ( .A1(n8670), .A2(n8669), .ZN(n13752) );
  NAND2_X1 U9136 ( .A1(n12001), .A2(n12000), .ZN(n14882) );
  INV_X1 U9137 ( .A(n14882), .ZN(n7998) );
  XOR2_X1 U9138 ( .A(n12390), .B(n12391), .Z(n7311) );
  NAND4_X1 U9139 ( .A1(n8941), .A2(n8940), .A3(n8939), .A4(n7334), .ZN(n10441)
         );
  INV_X1 U9140 ( .A(n14470), .ZN(n7693) );
  OR2_X1 U9141 ( .A1(n13966), .A2(n16159), .ZN(n7312) );
  INV_X1 U9142 ( .A(n11087), .ZN(n11067) );
  INV_X1 U9143 ( .A(n12714), .ZN(n7752) );
  AND2_X1 U9144 ( .A1(n13479), .A2(n13738), .ZN(n7313) );
  AND2_X1 U9145 ( .A1(n8595), .A2(n13563), .ZN(n7314) );
  INV_X1 U9146 ( .A(n13752), .ZN(n13559) );
  INV_X1 U9147 ( .A(n10442), .ZN(n7923) );
  AND2_X1 U9148 ( .A1(n7712), .A2(n7711), .ZN(n7315) );
  AND2_X1 U9149 ( .A1(n9768), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7316) );
  AND2_X1 U9150 ( .A1(n10436), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7317) );
  OR2_X1 U9151 ( .A1(n15720), .A2(n7570), .ZN(n7318) );
  INV_X1 U9152 ( .A(n16047), .ZN(n11899) );
  INV_X1 U9153 ( .A(n14115), .ZN(n14168) );
  NAND2_X1 U9154 ( .A1(n11883), .A2(n11882), .ZN(n14669) );
  INV_X1 U9155 ( .A(n14669), .ZN(n7604) );
  INV_X1 U9156 ( .A(n15082), .ZN(n7609) );
  INV_X1 U9157 ( .A(n14496), .ZN(n14524) );
  AND2_X2 U9158 ( .A1(n10136), .A2(n15408), .ZN(n16146) );
  NOR2_X1 U9159 ( .A1(n10366), .A2(n13170), .ZN(n7682) );
  AND2_X1 U9160 ( .A1(n7414), .A2(n8272), .ZN(n7319) );
  NAND2_X1 U9161 ( .A1(n12230), .A2(n12229), .ZN(n14511) );
  INV_X1 U9162 ( .A(n14511), .ZN(n7683) );
  AND2_X1 U9163 ( .A1(n7777), .A2(n10562), .ZN(n7781) );
  AND2_X1 U9164 ( .A1(n7828), .A2(n10633), .ZN(n7320) );
  NOR2_X1 U9165 ( .A1(n12180), .A2(n12179), .ZN(n7321) );
  INV_X1 U9166 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9477) );
  AND2_X1 U9167 ( .A1(n8817), .A2(n8816), .ZN(n7322) );
  AND2_X1 U9168 ( .A1(n8797), .A2(n11578), .ZN(n7323) );
  AND2_X1 U9169 ( .A1(n7842), .A2(n7840), .ZN(n7324) );
  AND2_X1 U9170 ( .A1(n7662), .A2(n7661), .ZN(n7325) );
  INV_X1 U9171 ( .A(n7853), .ZN(n7852) );
  OR2_X1 U9172 ( .A1(n7828), .A2(n11110), .ZN(n7326) );
  NAND2_X1 U9173 ( .A1(n8308), .A2(n7834), .ZN(n7327) );
  AND2_X1 U9174 ( .A1(n8269), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7328) );
  INV_X1 U9175 ( .A(n7839), .ZN(n7838) );
  AOI21_X1 U9176 ( .B1(n11467), .B2(n7840), .A(n7208), .ZN(n7839) );
  INV_X1 U9177 ( .A(n12849), .ZN(n7593) );
  INV_X1 U9178 ( .A(n14435), .ZN(n7372) );
  INV_X1 U9179 ( .A(n12858), .ZN(n7591) );
  INV_X1 U9180 ( .A(n12800), .ZN(n7920) );
  NAND2_X1 U9181 ( .A1(n13639), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7329) );
  NAND2_X1 U9182 ( .A1(n12641), .A2(n12792), .ZN(n12762) );
  INV_X1 U9183 ( .A(n13663), .ZN(n7672) );
  INV_X1 U9184 ( .A(n9772), .ZN(n14397) );
  INV_X1 U9185 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9478) );
  AND2_X1 U9186 ( .A1(n10150), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n10184) );
  NOR2_X1 U9187 ( .A1(n7673), .A2(n7672), .ZN(n7330) );
  AND2_X1 U9188 ( .A1(n7670), .A2(n7671), .ZN(n7331) );
  AND2_X1 U9189 ( .A1(n15977), .A2(n15856), .ZN(n15933) );
  AND2_X1 U9190 ( .A1(n7903), .A2(n7902), .ZN(n7332) );
  NAND2_X1 U9191 ( .A1(n8313), .A2(n8314), .ZN(n13656) );
  AND2_X1 U9192 ( .A1(n15148), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7333) );
  INV_X1 U9193 ( .A(n7717), .ZN(n7716) );
  OR2_X1 U9194 ( .A1(n8184), .A2(n13157), .ZN(n8185) );
  AND2_X1 U9195 ( .A1(n9773), .A2(n13101), .ZN(n13106) );
  NAND2_X1 U9196 ( .A1(n8135), .A2(n8134), .ZN(n13249) );
  NAND2_X1 U9197 ( .A1(n8141), .A2(n8140), .ZN(n13234) );
  OAI21_X1 U9198 ( .B1(n13303), .B2(n7482), .A(n8162), .ZN(n7481) );
  NAND3_X1 U9199 ( .A1(n7335), .A2(n14086), .A3(n14115), .ZN(n14053) );
  NOR2_X2 U9200 ( .A1(n14029), .A2(n14028), .ZN(n14031) );
  OAI21_X1 U9201 ( .B1(n14090), .B2(n14089), .A(n7337), .ZN(P2_U3192) );
  NAND2_X1 U9202 ( .A1(n7293), .A2(n7430), .ZN(n15130) );
  NAND2_X1 U9203 ( .A1(n14447), .A2(n7339), .ZN(P2_U3530) );
  NAND2_X1 U9204 ( .A1(n14535), .A2(n7340), .ZN(P2_U3498) );
  NAND2_X1 U9205 ( .A1(n7689), .A2(n7375), .ZN(n7374) );
  AOI22_X1 U9206 ( .A1(n12557), .A2(n12556), .B1(n14609), .B2(n15040), .ZN(
        n12558) );
  NAND2_X1 U9207 ( .A1(n7969), .A2(n7967), .ZN(P1_U3557) );
  NAND2_X1 U9208 ( .A1(n15651), .A2(n15650), .ZN(n7342) );
  XNOR2_X1 U9209 ( .A(n15489), .B(n15490), .ZN(n15491) );
  OAI21_X1 U9210 ( .B1(n15498), .B2(n15497), .A(n15496), .ZN(n15507) );
  NAND2_X1 U9211 ( .A1(n15517), .A2(n15518), .ZN(n7646) );
  INV_X1 U9212 ( .A(n7641), .ZN(n15541) );
  XNOR2_X1 U9213 ( .A(n15538), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15540) );
  NOR2_X1 U9214 ( .A1(n15546), .A2(n15545), .ZN(n15557) );
  XNOR2_X1 U9215 ( .A(n7657), .B(n7655), .ZN(SUB_1596_U4) );
  NAND3_X1 U9216 ( .A1(n7437), .A2(n13038), .A3(n11011), .ZN(n11034) );
  NAND3_X1 U9217 ( .A1(n15053), .A2(n15052), .A3(n7345), .ZN(n15131) );
  NAND2_X1 U9218 ( .A1(n12003), .A2(n12002), .ZN(n15009) );
  NAND2_X1 U9219 ( .A1(n11235), .A2(n11234), .ZN(n11427) );
  NAND2_X1 U9220 ( .A1(n7423), .A2(n10743), .ZN(n7422) );
  NAND2_X1 U9221 ( .A1(n7957), .A2(n7637), .ZN(n11903) );
  NAND2_X1 U9222 ( .A1(n14972), .A2(n14974), .ZN(n14971) );
  INV_X1 U9223 ( .A(n11233), .ZN(n7964) );
  AND3_X2 U9224 ( .A1(n7432), .A2(n9280), .A3(n7433), .ZN(n9416) );
  INV_X1 U9225 ( .A(n9275), .ZN(n7506) );
  NAND2_X1 U9226 ( .A1(n7506), .A2(n7952), .ZN(n15144) );
  INV_X1 U9227 ( .A(n7948), .ZN(P1_U3525) );
  NAND2_X1 U9228 ( .A1(n13307), .A2(n7305), .ZN(n7482) );
  NAND2_X1 U9229 ( .A1(n7349), .A2(n7348), .ZN(n13167) );
  NAND2_X1 U9230 ( .A1(n13164), .A2(n13163), .ZN(n7349) );
  NAND2_X1 U9231 ( .A1(n7481), .A2(n8158), .ZN(n13350) );
  OR2_X1 U9232 ( .A1(n13243), .A2(n8137), .ZN(n8133) );
  NAND2_X1 U9233 ( .A1(n7350), .A2(n8125), .ZN(n7467) );
  NAND3_X1 U9234 ( .A1(n13200), .A2(n13199), .A3(n7301), .ZN(n7350) );
  NOR2_X1 U9235 ( .A1(n9773), .A2(n13101), .ZN(n13102) );
  INV_X1 U9236 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7618) );
  OR4_X2 U9237 ( .A1(n13396), .A2(n13395), .A3(n14357), .A4(n13394), .ZN(
        n13397) );
  NAND4_X1 U9238 ( .A1(n7908), .A2(n7905), .A3(n7669), .A4(n7355), .ZN(
        P3_U3201) );
  OAI21_X1 U9239 ( .B1(n14259), .B2(n7794), .A(n7791), .ZN(n12343) );
  NOR2_X2 U9240 ( .A1(n15726), .A2(n13616), .ZN(n15748) );
  NAND2_X1 U9241 ( .A1(n10774), .A2(n7663), .ZN(n7659) );
  NAND2_X1 U9242 ( .A1(n7987), .A2(n10298), .ZN(n10435) );
  OR2_X2 U9243 ( .A1(n14863), .A2(n14862), .ZN(n14865) );
  NAND2_X1 U9244 ( .A1(n7703), .A2(n7700), .ZN(n14948) );
  AOI21_X1 U9245 ( .B1(n11400), .B2(n12680), .A(n7284), .ZN(n8796) );
  NAND2_X1 U9246 ( .A1(n8751), .A2(n8219), .ZN(n8298) );
  NAND2_X1 U9247 ( .A1(n13695), .A2(n13754), .ZN(n8862) );
  NAND2_X1 U9248 ( .A1(n9476), .A2(n8927), .ZN(n9473) );
  NAND2_X1 U9249 ( .A1(n10342), .A2(n10341), .ZN(n10446) );
  NAND2_X1 U9250 ( .A1(n14169), .A2(n8041), .ZN(n14046) );
  NAND2_X1 U9251 ( .A1(n9049), .A2(n9048), .ZN(n9104) );
  NAND2_X1 U9252 ( .A1(n7614), .A2(n9133), .ZN(n9174) );
  NAND2_X1 U9253 ( .A1(n14145), .A2(n8018), .ZN(n7554) );
  NAND2_X4 U9254 ( .A1(n10077), .A2(n12808), .ZN(n12523) );
  OAI21_X1 U9255 ( .B1(n10596), .B2(n10595), .A(n10594), .ZN(n10600) );
  INV_X1 U9256 ( .A(n7924), .ZN(n7922) );
  NAND2_X1 U9257 ( .A1(n7815), .A2(n13771), .ZN(n7814) );
  NAND2_X1 U9258 ( .A1(n13965), .A2(n7312), .ZN(P3_U3455) );
  NAND2_X1 U9259 ( .A1(n11957), .A2(n12609), .ZN(n11959) );
  NAND3_X1 U9260 ( .A1(n12986), .A2(n12985), .A3(n7300), .ZN(n7369) );
  NAND2_X1 U9261 ( .A1(n8007), .A2(n11986), .ZN(n12106) );
  NAND2_X1 U9262 ( .A1(n10869), .A2(n15944), .ZN(n10836) );
  AND2_X1 U9263 ( .A1(n7675), .A2(n7678), .ZN(n10869) );
  OR2_X2 U9264 ( .A1(n14375), .A2(n14361), .ZN(n14359) );
  OR2_X2 U9265 ( .A1(n13216), .A2(n11185), .ZN(n11506) );
  NOR2_X2 U9266 ( .A1(n14326), .A2(n7374), .ZN(n14264) );
  NOR2_X2 U9267 ( .A1(n15922), .A2(n7376), .ZN(n10063) );
  NAND2_X4 U9268 ( .A1(n15154), .A2(n15151), .ZN(n12049) );
  NAND2_X1 U9269 ( .A1(n7713), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9070) );
  NOR2_X1 U9270 ( .A1(n7882), .A2(n7788), .ZN(n7787) );
  NAND2_X1 U9271 ( .A1(n7554), .A2(n7553), .ZN(n14027) );
  INV_X1 U9272 ( .A(n10096), .ZN(n7558) );
  NOR2_X1 U9273 ( .A1(n11267), .A2(n8042), .ZN(n11272) );
  INV_X1 U9274 ( .A(n10328), .ZN(n10335) );
  AOI21_X2 U9275 ( .B1(n12399), .B2(n10846), .A(n10845), .ZN(n12401) );
  NOR2_X2 U9276 ( .A1(n14147), .A2(n14146), .ZN(n14145) );
  NAND3_X1 U9277 ( .A1(n7772), .A2(n12650), .A3(n12649), .ZN(n7771) );
  NAND2_X1 U9278 ( .A1(n8793), .A2(n12677), .ZN(n11400) );
  NAND2_X1 U9279 ( .A1(n7747), .A2(n7745), .ZN(n13846) );
  XNOR2_X2 U9280 ( .A(n12088), .B(n12087), .ZN(n14598) );
  XNOR2_X1 U9281 ( .A(n12366), .B(n13403), .ZN(n14456) );
  OR2_X1 U9282 ( .A1(n13414), .A2(n13413), .ZN(n13415) );
  NAND2_X1 U9283 ( .A1(n7926), .A2(n7925), .ZN(n7924) );
  XNOR2_X1 U9284 ( .A(n12441), .B(n12439), .ZN(n14722) );
  NAND2_X1 U9285 ( .A1(n8072), .A2(n8071), .ZN(n14691) );
  AOI21_X2 U9286 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n11328), .A(n11308), .ZN(
        n11309) );
  NAND2_X4 U9287 ( .A1(n10077), .A2(n10642), .ZN(n12525) );
  XNOR2_X1 U9288 ( .A(n9626), .B(n7381), .ZN(n14604) );
  INV_X1 U9289 ( .A(n8237), .ZN(n7383) );
  NAND2_X1 U9290 ( .A1(n8339), .A2(n7394), .ZN(n7392) );
  NAND2_X1 U9291 ( .A1(n8432), .A2(n7285), .ZN(n7400) );
  NAND3_X1 U9292 ( .A1(n7401), .A2(n7403), .A3(n8450), .ZN(n7399) );
  NAND3_X1 U9293 ( .A1(n7416), .A2(n13722), .A3(n13740), .ZN(n7415) );
  XNOR2_X2 U9294 ( .A(n13479), .B(n13738), .ZN(n13722) );
  NAND2_X1 U9295 ( .A1(n10619), .A2(n10274), .ZN(n7417) );
  NAND2_X1 U9296 ( .A1(n9423), .A2(n13026), .ZN(n10272) );
  NAND3_X1 U9297 ( .A1(n7422), .A2(n7424), .A3(n10746), .ZN(n10920) );
  NAND3_X1 U9298 ( .A1(n10673), .A2(n7425), .A3(n13032), .ZN(n7424) );
  NAND2_X1 U9299 ( .A1(n13032), .A2(n7946), .ZN(n7426) );
  NOR2_X4 U9300 ( .A1(n7942), .A2(n7431), .ZN(n15854) );
  AND2_X1 U9301 ( .A1(n9277), .A2(n9276), .ZN(n7432) );
  NAND2_X1 U9302 ( .A1(n15854), .A2(n14753), .ZN(n12813) );
  AND2_X2 U9303 ( .A1(n9278), .A2(n12797), .ZN(n9339) );
  XNOR2_X2 U9304 ( .A(n7436), .B(n7435), .ZN(n12797) );
  NAND2_X1 U9305 ( .A1(n11189), .A2(n11188), .ZN(n11494) );
  NAND2_X1 U9306 ( .A1(n9774), .A2(n7441), .ZN(n9970) );
  OAI22_X1 U9307 ( .A1(n7441), .A2(n10660), .B1(n13109), .B2(n14200), .ZN(
        n10868) );
  XNOR2_X1 U9308 ( .A(n10661), .B(n7441), .ZN(n10663) );
  XNOR2_X1 U9309 ( .A(n7441), .B(n10660), .ZN(n15862) );
  XNOR2_X2 U9310 ( .A(n13109), .B(n14200), .ZN(n7441) );
  NAND3_X1 U9311 ( .A1(n10510), .A2(n10112), .A3(n7448), .ZN(n7446) );
  NAND2_X1 U9312 ( .A1(n7444), .A2(n9976), .ZN(n7448) );
  INV_X1 U9313 ( .A(n13374), .ZN(n7444) );
  NAND3_X1 U9314 ( .A1(n7446), .A2(n7445), .A3(n10115), .ZN(n10367) );
  NAND3_X1 U9315 ( .A1(n7448), .A2(n10112), .A3(n7449), .ZN(n7445) );
  NAND2_X1 U9316 ( .A1(n10510), .A2(n13374), .ZN(n7447) );
  INV_X1 U9317 ( .A(n9976), .ZN(n7449) );
  OAI21_X1 U9318 ( .B1(n11789), .B2(n7452), .A(n7450), .ZN(n14409) );
  OAI21_X1 U9319 ( .B1(n11789), .B2(n11790), .A(n11791), .ZN(n12226) );
  NOR2_X2 U9320 ( .A1(n9578), .A2(n12174), .ZN(n9887) );
  NAND2_X1 U9321 ( .A1(n7464), .A2(n13213), .ZN(n7463) );
  INV_X1 U9322 ( .A(n7467), .ZN(n7464) );
  NAND2_X1 U9323 ( .A1(n7466), .A2(n13211), .ZN(n7465) );
  NAND2_X1 U9324 ( .A1(n7467), .A2(n13212), .ZN(n7466) );
  NAND2_X2 U9325 ( .A1(n9492), .A2(n13408), .ZN(n11785) );
  XNOR2_X2 U9326 ( .A(n9485), .B(n9572), .ZN(n9492) );
  NAND2_X1 U9327 ( .A1(n11721), .A2(n7478), .ZN(n7476) );
  NAND2_X1 U9328 ( .A1(n7476), .A2(n7477), .ZN(n14406) );
  OAI21_X1 U9329 ( .B1(n10965), .B2(n7485), .A(n7483), .ZN(n10784) );
  NAND2_X1 U9330 ( .A1(n13284), .A2(n7197), .ZN(n7488) );
  NAND2_X1 U9331 ( .A1(n7488), .A2(n7489), .ZN(n13295) );
  OR2_X1 U9332 ( .A1(n13227), .A2(n8143), .ZN(n7493) );
  NAND3_X1 U9333 ( .A1(n13252), .A2(n7304), .A3(n7497), .ZN(n8128) );
  NAND3_X1 U9334 ( .A1(n8133), .A2(n8136), .A3(n13251), .ZN(n7497) );
  NAND2_X1 U9335 ( .A1(n7505), .A2(n7504), .ZN(n12871) );
  NAND4_X1 U9336 ( .A1(n8945), .A2(n10442), .A3(n8094), .A4(n7303), .ZN(n9275)
         );
  OAI21_X1 U9337 ( .B1(n7510), .B2(n12829), .A(n7508), .ZN(n7507) );
  NAND2_X1 U9338 ( .A1(n7512), .A2(n7513), .ZN(n12950) );
  NAND2_X1 U9339 ( .A1(n12909), .A2(n7515), .ZN(n7512) );
  NAND2_X1 U9340 ( .A1(n12975), .A2(n7306), .ZN(n7519) );
  INV_X1 U9341 ( .A(n12976), .ZN(n7521) );
  OAI22_X1 U9342 ( .A1(n7199), .A2(n7522), .B1(n12890), .B2(n7523), .ZN(n12893) );
  INV_X1 U9343 ( .A(n12889), .ZN(n7523) );
  NAND2_X1 U9344 ( .A1(n12967), .A2(n7525), .ZN(n7524) );
  INV_X1 U9345 ( .A(n12968), .ZN(n7527) );
  NAND2_X1 U9346 ( .A1(n7530), .A2(n7529), .ZN(n14458) );
  OR2_X1 U9347 ( .A1(n16142), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n7529) );
  OR2_X1 U9348 ( .A1(n7612), .A2(n9350), .ZN(n7531) );
  NAND3_X1 U9349 ( .A1(n7613), .A2(n9353), .A3(n7612), .ZN(n7532) );
  NAND2_X1 U9350 ( .A1(n7532), .A2(n7533), .ZN(n9441) );
  NAND2_X2 U9351 ( .A1(n7535), .A2(n12297), .ZN(n14475) );
  NAND2_X1 U9352 ( .A1(n9762), .A2(n9760), .ZN(n7537) );
  OAI21_X2 U9353 ( .B1(n9439), .B2(n7627), .A(n7625), .ZN(n9762) );
  OAI21_X2 U9354 ( .B1(n9762), .B2(n7540), .A(n7275), .ZN(n11088) );
  NAND3_X1 U9355 ( .A1(n8012), .A2(n8010), .A3(n8011), .ZN(n8009) );
  XNOR2_X2 U9356 ( .A(n14031), .B(n14030), .ZN(n14055) );
  NAND4_X1 U9357 ( .A1(n7881), .A2(n7879), .A3(n7878), .A4(n7880), .ZN(n7788)
         );
  INV_X1 U9358 ( .A(n7546), .ZN(n9561) );
  NAND4_X1 U9359 ( .A1(n7548), .A2(n7549), .A3(n7547), .A4(n7299), .ZN(n7546)
         );
  NAND3_X1 U9360 ( .A1(n7552), .A2(n9014), .A3(n7550), .ZN(n8047) );
  XNOR2_X1 U9361 ( .A(n14027), .B(n14026), .ZN(n12392) );
  AND2_X2 U9362 ( .A1(n10446), .A2(n10445), .ZN(n12399) );
  AOI21_X2 U9363 ( .B1(n11714), .B2(n7563), .A(n7281), .ZN(n12418) );
  INV_X2 U9364 ( .A(n11374), .ZN(n14032) );
  NAND2_X1 U9365 ( .A1(n15721), .A2(n7191), .ZN(n7568) );
  OAI211_X1 U9366 ( .C1(n15721), .C2(n7318), .A(n7568), .B(n7569), .ZN(n15741)
         );
  NOR2_X1 U9367 ( .A1(n15741), .A2(n8325), .ZN(n15740) );
  NAND2_X1 U9368 ( .A1(n9939), .A2(n9790), .ZN(n9791) );
  INV_X1 U9369 ( .A(n10184), .ZN(n7586) );
  NOR2_X2 U9370 ( .A1(n10441), .A2(n8944), .ZN(n8945) );
  AND2_X2 U9371 ( .A1(n8938), .A2(n9036), .ZN(n10442) );
  NOR2_X2 U9373 ( .A1(n11008), .A2(n12864), .ZN(n11050) );
  AND2_X1 U9374 ( .A1(n7185), .A2(n7600), .ZN(n14850) );
  NAND2_X1 U9375 ( .A1(n7184), .A2(n12555), .ZN(n12543) );
  NAND2_X1 U9376 ( .A1(n7185), .A2(n7601), .ZN(n14849) );
  OAI211_X1 U9377 ( .C1(n7601), .C2(n7599), .A(n7598), .B(n7596), .ZN(n15023)
         );
  NAND2_X1 U9378 ( .A1(n7185), .A2(n7597), .ZN(n7596) );
  AND2_X1 U9379 ( .A1(n7601), .A2(n7599), .ZN(n7597) );
  OR2_X1 U9380 ( .A1(n7185), .A2(n7599), .ZN(n7598) );
  NAND4_X1 U9381 ( .A1(n7619), .A2(n7618), .A3(P2_ADDR_REG_19__SCAN_IN), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n7620) );
  NAND4_X1 U9382 ( .A1(n7624), .A2(n7623), .A3(P3_ADDR_REG_19__SCAN_IN), .A4(
        n15828), .ZN(n7621) );
  INV_X1 U9383 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7624) );
  OAI21_X1 U9384 ( .B1(n9441), .B2(n9636), .A(n9640), .ZN(n7626) );
  NAND2_X1 U9385 ( .A1(n14879), .A2(n7630), .ZN(n7628) );
  NAND2_X1 U9386 ( .A1(n7629), .A2(n7628), .ZN(n12557) );
  NAND2_X1 U9387 ( .A1(n14929), .A2(n7638), .ZN(n14915) );
  NAND2_X1 U9388 ( .A1(n7640), .A2(n15955), .ZN(n15038) );
  XNOR2_X1 U9389 ( .A(n12558), .B(n13058), .ZN(n7640) );
  NAND2_X1 U9390 ( .A1(n7646), .A2(n15519), .ZN(n15520) );
  NAND2_X1 U9391 ( .A1(n7654), .A2(n15558), .ZN(n15566) );
  NAND2_X1 U9392 ( .A1(n9852), .A2(n9806), .ZN(n9805) );
  NAND2_X1 U9393 ( .A1(n9933), .A2(n9872), .ZN(n9806) );
  OR2_X1 U9394 ( .A1(n9933), .A2(n9872), .ZN(n7658) );
  NOR2_X2 U9395 ( .A1(n7223), .A2(n13614), .ZN(n13615) );
  NOR2_X2 U9396 ( .A1(n15803), .A2(n15804), .ZN(n15802) );
  NAND3_X1 U9397 ( .A1(n7668), .A2(n7667), .A3(n7670), .ZN(n7666) );
  NAND2_X1 U9398 ( .A1(n7674), .A2(n13663), .ZN(n7667) );
  AOI21_X1 U9399 ( .B1(n13624), .B2(n13623), .A(n13622), .ZN(n13652) );
  INV_X2 U9400 ( .A(n15864), .ZN(n13109) );
  NAND2_X1 U9401 ( .A1(n15864), .A2(n13101), .ZN(n10870) );
  AND3_X2 U9402 ( .A1(n9613), .A2(n9614), .A3(n7676), .ZN(n15864) );
  INV_X2 U9403 ( .A(n15904), .ZN(n7678) );
  NOR2_X2 U9404 ( .A1(n14418), .A2(n14570), .ZN(n14400) );
  XNOR2_X2 U9405 ( .A(n7687), .B(P3_IR_REG_2__SCAN_IN), .ZN(n9956) );
  NAND2_X2 U9406 ( .A1(n9078), .A2(n7713), .ZN(n15154) );
  NAND2_X2 U9407 ( .A1(n9071), .A2(n9273), .ZN(n15151) );
  NAND2_X1 U9408 ( .A1(n7977), .A2(n7704), .ZN(n7703) );
  NAND3_X1 U9409 ( .A1(n8945), .A2(n10442), .A3(n8094), .ZN(n9067) );
  NAND4_X1 U9410 ( .A1(n8945), .A2(n10442), .A3(n8094), .A4(n7287), .ZN(n7713)
         );
  NAND2_X1 U9411 ( .A1(n10471), .A2(n7292), .ZN(n10730) );
  OAI21_X2 U9412 ( .B1(n7210), .B2(n7716), .A(n7714), .ZN(n14877) );
  NAND2_X1 U9413 ( .A1(n8521), .A2(n7726), .ZN(n7724) );
  NAND2_X1 U9414 ( .A1(n8876), .A2(n7731), .ZN(n7730) );
  NAND4_X1 U9415 ( .A1(n12770), .A2(n12769), .A3(n12772), .A4(n7741), .ZN(
        n7740) );
  NAND2_X1 U9416 ( .A1(n15387), .A2(n7748), .ZN(n7747) );
  NAND4_X2 U9417 ( .A1(n8320), .A2(n8213), .A3(n7755), .A4(n8209), .ZN(n7758)
         );
  AND2_X2 U9418 ( .A1(n8172), .A2(n8214), .ZN(n7755) );
  NOR2_X2 U9419 ( .A1(n7758), .A2(n7756), .ZN(n8751) );
  NAND2_X1 U9420 ( .A1(n7767), .A2(n7762), .ZN(n7761) );
  NAND2_X1 U9421 ( .A1(n7767), .A2(n7763), .ZN(n7766) );
  NAND2_X1 U9422 ( .A1(n13825), .A2(n7288), .ZN(n8799) );
  AND2_X1 U9423 ( .A1(n8290), .A2(n8291), .ZN(n8222) );
  NAND2_X1 U9424 ( .A1(n8290), .A2(n7769), .ZN(n14021) );
  OAI21_X1 U9425 ( .B1(n12604), .B2(n10420), .A(n12646), .ZN(n7772) );
  NAND2_X1 U9426 ( .A1(n7771), .A2(n12650), .ZN(n10876) );
  AND2_X1 U9427 ( .A1(n12649), .A2(n12650), .ZN(n15879) );
  OAI21_X1 U9428 ( .B1(n7361), .B2(n10420), .A(n12646), .ZN(n15871) );
  INV_X1 U9429 ( .A(n15879), .ZN(n15870) );
  NAND2_X1 U9430 ( .A1(n10370), .A2(n7781), .ZN(n7780) );
  INV_X1 U9431 ( .A(n10559), .ZN(n7783) );
  NAND2_X1 U9432 ( .A1(n7780), .A2(n7778), .ZN(n10565) );
  AND2_X1 U9433 ( .A1(n7779), .A2(n10563), .ZN(n7778) );
  OAI21_X1 U9434 ( .B1(n10370), .B2(n7783), .A(n7781), .ZN(n10970) );
  INV_X1 U9435 ( .A(n7795), .ZN(n7794) );
  NAND3_X1 U9436 ( .A1(n11153), .A2(n11152), .A3(n13384), .ZN(n11189) );
  OAI21_X2 U9437 ( .B1(n11733), .B2(n11732), .A(n11734), .ZN(n11789) );
  NAND2_X1 U9438 ( .A1(n7802), .A2(n7798), .ZN(n14370) );
  INV_X1 U9439 ( .A(n7799), .ZN(n7798) );
  OAI21_X1 U9440 ( .B1(n14390), .B2(n7800), .A(n12243), .ZN(n7799) );
  NAND2_X1 U9441 ( .A1(n14409), .A2(n7803), .ZN(n7802) );
  NOR2_X1 U9442 ( .A1(n14390), .A2(n7804), .ZN(n7803) );
  NAND2_X1 U9443 ( .A1(n10720), .A2(n13383), .ZN(n11153) );
  NOR3_X4 U9444 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .A3(
        P3_IR_REG_6__SCAN_IN), .ZN(n8213) );
  NAND2_X1 U9445 ( .A1(n10565), .A2(n10564), .ZN(n10567) );
  XNOR2_X2 U9446 ( .A(n13127), .B(n9973), .ZN(n13371) );
  INV_X1 U9447 ( .A(n8376), .ZN(n8209) );
  OR2_X2 U9448 ( .A1(n14485), .A2(n14359), .ZN(n14344) );
  NOR2_X2 U9449 ( .A1(n13224), .A2(n11506), .ZN(n11538) );
  OR2_X2 U9450 ( .A1(n15064), .A2(n14934), .ZN(n14921) );
  NOR2_X2 U9451 ( .A1(n14871), .A2(n14885), .ZN(n14869) );
  NOR2_X4 U9452 ( .A1(n15014), .A2(n15104), .ZN(n15013) );
  NAND2_X1 U9453 ( .A1(n8612), .A2(n8611), .ZN(n8273) );
  NAND2_X1 U9454 ( .A1(n8657), .A2(n8656), .ZN(n8278) );
  NAND2_X1 U9455 ( .A1(n8266), .A2(n8265), .ZN(n8568) );
  NOR2_X2 U9456 ( .A1(n15573), .A2(n15572), .ZN(n15578) );
  AOI21_X2 U9457 ( .B1(n15614), .B2(n15613), .A(n15612), .ZN(n15621) );
  OR2_X2 U9458 ( .A1(n13380), .A2(n10567), .ZN(n10717) );
  NAND2_X1 U9459 ( .A1(n13426), .A2(n13480), .ZN(n7806) );
  INV_X1 U9460 ( .A(n13426), .ZN(n7809) );
  NAND2_X1 U9461 ( .A1(n13451), .A2(n13452), .ZN(n8703) );
  AND3_X2 U9462 ( .A1(n8211), .A2(n8212), .A3(n8210), .ZN(n8320) );
  NOR2_X1 U9463 ( .A1(n10395), .A2(n10396), .ZN(n10394) );
  INV_X1 U9464 ( .A(n7813), .ZN(n10165) );
  NAND2_X1 U9465 ( .A1(n7814), .A2(n8655), .ZN(n8661) );
  NAND2_X1 U9466 ( .A1(n13505), .A2(n7289), .ZN(n8662) );
  INV_X1 U9467 ( .A(n8660), .ZN(n7816) );
  NAND2_X1 U9468 ( .A1(n13455), .A2(n7820), .ZN(n7819) );
  NAND2_X1 U9469 ( .A1(n13455), .A2(n8704), .ZN(n13525) );
  NAND2_X1 U9470 ( .A1(n10633), .A2(n11109), .ZN(n7827) );
  NAND2_X1 U9471 ( .A1(n10633), .A2(n7832), .ZN(n10987) );
  INV_X1 U9472 ( .A(n10986), .ZN(n7830) );
  NAND2_X1 U9473 ( .A1(n8308), .A2(n7833), .ZN(n8311) );
  NAND2_X1 U9474 ( .A1(n11466), .A2(n7840), .ZN(n7837) );
  INV_X1 U9475 ( .A(n11467), .ZN(n7845) );
  AOI21_X1 U9476 ( .B1(n11184), .B2(n7860), .A(n7858), .ZN(n7857) );
  INV_X1 U9477 ( .A(n7857), .ZN(n11547) );
  NAND2_X1 U9478 ( .A1(n14383), .A2(n7866), .ZN(n7864) );
  NAND2_X1 U9479 ( .A1(n7864), .A2(n7865), .ZN(n14358) );
  XNOR2_X2 U9480 ( .A(n7870), .B(n7869), .ZN(n12174) );
  NOR2_X1 U9481 ( .A1(n9575), .A2(n14582), .ZN(n7870) );
  NOR2_X2 U9482 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n9649) );
  NOR2_X2 U9483 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7878) );
  NOR2_X2 U9485 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n7880) );
  NOR2_X1 U9486 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n7883) );
  NAND2_X1 U9487 ( .A1(n9877), .A2(n7677), .ZN(n9880) );
  NAND2_X1 U9488 ( .A1(n10052), .A2(n7677), .ZN(n9886) );
  NAND2_X1 U9489 ( .A1(n10221), .A2(n7677), .ZN(n9960) );
  NAND2_X1 U9490 ( .A1(n10261), .A2(n7677), .ZN(n10006) );
  NAND2_X1 U9491 ( .A1(n10472), .A2(n7677), .ZN(n10327) );
  NAND2_X1 U9492 ( .A1(n10731), .A2(n7677), .ZN(n10449) );
  NAND2_X1 U9493 ( .A1(n10906), .A2(n7890), .ZN(n10553) );
  NAND2_X1 U9494 ( .A1(n10997), .A2(n7890), .ZN(n10689) );
  NAND2_X1 U9495 ( .A1(n11035), .A2(n7890), .ZN(n10693) );
  NAND2_X1 U9496 ( .A1(n11229), .A2(n7890), .ZN(n11139) );
  NAND2_X1 U9497 ( .A1(n11412), .A2(n7890), .ZN(n11182) );
  NAND2_X1 U9498 ( .A1(n11626), .A2(n7890), .ZN(n11537) );
  NAND2_X1 U9499 ( .A1(n11488), .A2(n7890), .ZN(n11492) );
  NAND2_X1 U9500 ( .A1(n11722), .A2(n7890), .ZN(n11724) );
  NAND2_X1 U9501 ( .A1(n11880), .A2(n7890), .ZN(n11788) );
  NAND2_X1 U9502 ( .A1(n12228), .A2(n7890), .ZN(n12230) );
  NAND2_X1 U9503 ( .A1(n12244), .A2(n7890), .ZN(n12246) );
  NAND2_X1 U9504 ( .A1(n12233), .A2(n7890), .ZN(n12236) );
  NAND2_X1 U9505 ( .A1(n12259), .A2(n7890), .ZN(n12261) );
  NAND2_X1 U9506 ( .A1(n12271), .A2(n7890), .ZN(n12273) );
  NAND2_X1 U9507 ( .A1(n12283), .A2(n7890), .ZN(n12285) );
  NAND2_X1 U9508 ( .A1(n14598), .A2(n7890), .ZN(n12217) );
  NAND2_X1 U9509 ( .A1(n14594), .A2(n7890), .ZN(n12205) );
  NAND2_X1 U9510 ( .A1(n12368), .A2(n7890), .ZN(n12311) );
  NAND2_X1 U9511 ( .A1(n14586), .A2(n7890), .ZN(n12334) );
  NAND2_X1 U9512 ( .A1(n14589), .A2(n7890), .ZN(n12323) );
  NAND2_X1 U9513 ( .A1(n14581), .A2(n7890), .ZN(n13332) );
  NAND2_X1 U9514 ( .A1(n7895), .A2(n9794), .ZN(n9792) );
  NAND2_X1 U9515 ( .A1(n7912), .A2(n7910), .ZN(n12956) );
  NAND2_X1 U9516 ( .A1(n12952), .A2(n7913), .ZN(n7912) );
  OAI211_X1 U9517 ( .C1(n7919), .C2(n7918), .A(n12812), .B(n7916), .ZN(n12819)
         );
  NAND2_X1 U9518 ( .A1(n7917), .A2(n12807), .ZN(n7916) );
  INV_X1 U9519 ( .A(n12804), .ZN(n7917) );
  INV_X1 U9520 ( .A(n12807), .ZN(n7918) );
  NAND2_X1 U9521 ( .A1(n12803), .A2(n12805), .ZN(n7919) );
  NAND2_X2 U9522 ( .A1(n12997), .A2(n12998), .ZN(n12884) );
  INV_X1 U9523 ( .A(n10441), .ZN(n7926) );
  NAND2_X1 U9524 ( .A1(n7927), .A2(n7928), .ZN(n12909) );
  NAND3_X1 U9525 ( .A1(n12903), .A2(n7297), .A3(n12902), .ZN(n7927) );
  NAND2_X1 U9526 ( .A1(n12898), .A2(n12899), .ZN(n12897) );
  NAND2_X1 U9527 ( .A1(n12878), .A2(n12879), .ZN(n12877) );
  INV_X1 U9528 ( .A(n13014), .ZN(n13022) );
  NAND2_X1 U9529 ( .A1(n12852), .A2(n12853), .ZN(n12851) );
  INV_X1 U9530 ( .A(n10546), .ZN(n7941) );
  AND2_X2 U9531 ( .A1(n12813), .A2(n12815), .ZN(n13028) );
  NOR2_X1 U9532 ( .A1(n16071), .A2(n12145), .ZN(n7949) );
  NAND2_X1 U9533 ( .A1(n11625), .A2(n7958), .ZN(n7957) );
  XNOR2_X1 U9534 ( .A(n9032), .B(n7965), .ZN(n9877) );
  NAND2_X1 U9535 ( .A1(n10024), .A2(n10023), .ZN(n10296) );
  NOR2_X1 U9536 ( .A1(n13055), .A2(n7996), .ZN(n7995) );
  NAND2_X1 U9537 ( .A1(n7992), .A2(n7990), .ZN(n12542) );
  INV_X1 U9538 ( .A(n14871), .ZN(n7999) );
  OAI21_X2 U9539 ( .B1(n11350), .B2(n8000), .A(n11354), .ZN(n11567) );
  NAND2_X1 U9540 ( .A1(n11981), .A2(n11980), .ZN(n12088) );
  NAND2_X1 U9541 ( .A1(n11981), .A2(n7291), .ZN(n8007) );
  OAI21_X2 U9542 ( .B1(n11974), .B2(n11973), .A(n11977), .ZN(n11979) );
  INV_X1 U9543 ( .A(n14031), .ZN(n8015) );
  OAI21_X1 U9544 ( .B1(n14145), .B2(n8017), .A(n8018), .ZN(n14092) );
  INV_X1 U9545 ( .A(n7196), .ZN(n8017) );
  INV_X1 U9546 ( .A(n14126), .ZN(n8028) );
  INV_X1 U9547 ( .A(n14086), .ZN(n14075) );
  NAND2_X1 U9548 ( .A1(n14086), .A2(n8038), .ZN(n14087) );
  OR2_X1 U9549 ( .A1(n14041), .A2(n14042), .ZN(n8041) );
  NAND2_X1 U9550 ( .A1(n9708), .A2(n9630), .ZN(n9631) );
  NAND2_X1 U9551 ( .A1(n8045), .A2(n9629), .ZN(n9708) );
  INV_X1 U9552 ( .A(n9710), .ZN(n8045) );
  NAND2_X1 U9553 ( .A1(n9618), .A2(n9630), .ZN(n9710) );
  NAND2_X1 U9554 ( .A1(n8047), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n11106) );
  OAI21_X1 U9555 ( .B1(n8047), .B2(n9486), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9487) );
  OR2_X1 U9556 ( .A1(n12049), .A2(n14758), .ZN(n9284) );
  NAND2_X1 U9557 ( .A1(n14710), .A2(n7295), .ZN(n8053) );
  NAND2_X1 U9558 ( .A1(n14710), .A2(n14711), .ZN(n8060) );
  OAI211_X1 U9559 ( .C1(n14710), .C2(n8058), .A(n8054), .B(n8053), .ZN(n12536)
         );
  NAND2_X1 U9560 ( .A1(n14613), .A2(n8068), .ZN(n8065) );
  NAND2_X1 U9561 ( .A1(n8065), .A2(n8066), .ZN(n14641) );
  NAND2_X1 U9562 ( .A1(n14621), .A2(n8073), .ZN(n8072) );
  NAND2_X1 U9563 ( .A1(n11477), .A2(n8082), .ZN(n8085) );
  INV_X1 U9564 ( .A(n8085), .ZN(n11814) );
  INV_X1 U9565 ( .A(n11478), .ZN(n8088) );
  NAND2_X1 U9566 ( .A1(n10819), .A2(n8090), .ZN(n8093) );
  INV_X1 U9567 ( .A(n8093), .ZN(n11120) );
  INV_X1 U9568 ( .A(n9074), .ZN(n8094) );
  NAND2_X1 U9569 ( .A1(n11691), .A2(n8097), .ZN(n8096) );
  INV_X1 U9570 ( .A(n8106), .ZN(n13709) );
  NAND3_X1 U9571 ( .A1(n8301), .A2(n8299), .A3(n8122), .ZN(n8121) );
  NAND3_X1 U9572 ( .A1(n9798), .A2(n8123), .A3(n8207), .ZN(n8376) );
  OAI21_X2 U9573 ( .B1(n15389), .B2(n8833), .A(n8839), .ZN(n13821) );
  NAND2_X2 U9574 ( .A1(n8124), .A2(n8830), .ZN(n15389) );
  INV_X1 U9575 ( .A(n13295), .ZN(n13296) );
  NAND2_X1 U9576 ( .A1(n13243), .A2(n8136), .ZN(n8135) );
  NAND2_X1 U9577 ( .A1(n13227), .A2(n8142), .ZN(n8141) );
  INV_X1 U9578 ( .A(n13225), .ZN(n8145) );
  INV_X1 U9579 ( .A(n13172), .ZN(n8149) );
  NAND3_X1 U9580 ( .A1(n13167), .A2(n13166), .A3(n8147), .ZN(n8146) );
  NAND2_X1 U9581 ( .A1(n13171), .A2(n13172), .ZN(n8147) );
  NAND3_X1 U9582 ( .A1(n13182), .A2(n13183), .A3(n8151), .ZN(n8153) );
  NAND2_X1 U9583 ( .A1(n13187), .A2(n13186), .ZN(n8151) );
  NAND2_X1 U9584 ( .A1(n8153), .A2(n8152), .ZN(n13195) );
  NAND3_X1 U9585 ( .A1(n13268), .A2(n13267), .A3(n7302), .ZN(n8157) );
  NAND2_X1 U9586 ( .A1(n11570), .A2(n11569), .ZN(n11748) );
  AOI21_X1 U9587 ( .B1(n13537), .B2(n8551), .A(n8174), .ZN(n13464) );
  NAND2_X1 U9588 ( .A1(n12597), .A2(n8178), .ZN(n12629) );
  XNOR2_X1 U9589 ( .A(n12332), .B(n12331), .ZN(n14586) );
  OR2_X1 U9590 ( .A1(n11748), .A2(SI_22_), .ZN(n11749) );
  XNOR2_X1 U9591 ( .A(n12557), .B(n13055), .ZN(n12152) );
  NAND2_X1 U9592 ( .A1(n11088), .A2(n11066), .ZN(n11072) );
  NAND2_X1 U9593 ( .A1(n11567), .A2(n11566), .ZN(n11570) );
  XNOR2_X1 U9594 ( .A(n11567), .B(n11565), .ZN(n12259) );
  OR2_X1 U9595 ( .A1(n8290), .A2(n8221), .ZN(n8292) );
  INV_X1 U9596 ( .A(n12095), .ZN(n12142) );
  NAND2_X1 U9597 ( .A1(n8226), .A2(n8228), .ZN(n8405) );
  CLKBUF_X1 U9598 ( .A(n10087), .Z(n15875) );
  NAND4_X2 U9599 ( .A1(n8183), .A2(n9625), .A3(n9624), .A4(n9623), .ZN(n9773)
         );
  OR2_X1 U9600 ( .A1(n12199), .A2(n16154), .ZN(n8167) );
  OR2_X1 U9601 ( .A1(n12199), .A2(n16159), .ZN(n8168) );
  OR2_X1 U9602 ( .A1(n13898), .A2(n16159), .ZN(n8169) );
  NAND2_X2 U9603 ( .A1(n10317), .A2(n15892), .ZN(n15899) );
  AND2_X1 U9604 ( .A1(n13800), .A2(n13795), .ZN(n8170) );
  AND2_X1 U9605 ( .A1(n10333), .A2(n10332), .ZN(n8171) );
  AND2_X2 U9606 ( .A1(n8417), .A2(n8208), .ZN(n8172) );
  AND2_X1 U9607 ( .A1(n9562), .A2(n9563), .ZN(n8173) );
  NOR2_X1 U9608 ( .A1(n8550), .A2(n13542), .ZN(n8174) );
  AND3_X1 U9609 ( .A1(n12628), .A2(n12627), .A3(n12626), .ZN(n8175) );
  OR2_X1 U9610 ( .A1(n12441), .A2(n12440), .ZN(n8176) );
  CLKBUF_X3 U9611 ( .A(n8390), .Z(n8884) );
  INV_X1 U9612 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n8195) );
  NOR2_X1 U9613 ( .A1(n12685), .A2(n11579), .ZN(n8177) );
  INV_X1 U9614 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n15585) );
  AND2_X1 U9615 ( .A1(n12624), .A2(n12641), .ZN(n8178) );
  AND2_X1 U9616 ( .A1(n13072), .A2(n13071), .ZN(n8179) );
  NOR3_X1 U9617 ( .A1(n14253), .A2(n14252), .A3(n14416), .ZN(n8180) );
  NAND2_X1 U9618 ( .A1(n13837), .A2(n13840), .ZN(n8181) );
  INV_X1 U9619 ( .A(n13037), .ZN(n10923) );
  OR2_X1 U9620 ( .A1(n9620), .A2(n9619), .ZN(n8183) );
  INV_X1 U9621 ( .A(n13034), .ZN(n10476) );
  AND2_X1 U9622 ( .A1(n9288), .A2(n12808), .ZN(n8186) );
  AND2_X1 U9623 ( .A1(n14198), .A2(n13351), .ZN(n13128) );
  NAND2_X1 U9624 ( .A1(n12825), .A2(n12824), .ZN(n12826) );
  INV_X1 U9625 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8208) );
  INV_X1 U9626 ( .A(n11256), .ZN(n11217) );
  INV_X1 U9627 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8942) );
  AND2_X1 U9628 ( .A1(n11070), .A2(n11090), .ZN(n11071) );
  INV_X1 U9629 ( .A(n8576), .ZN(n8197) );
  INV_X1 U9630 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n15356) );
  INV_X1 U9631 ( .A(n8857), .ZN(n8858) );
  NOR2_X1 U9632 ( .A1(n7227), .A2(n8838), .ZN(n8839) );
  INV_X1 U9633 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n8192) );
  AND2_X1 U9634 ( .A1(n13878), .A2(n12704), .ZN(n12703) );
  INV_X1 U9635 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10007) );
  INV_X1 U9636 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n9572) );
  OAI22_X1 U9637 ( .A1(n9416), .A2(n12525), .B1(n15854), .B2(n12523), .ZN(
        n9289) );
  INV_X1 U9638 ( .A(n11432), .ZN(n11418) );
  INV_X1 U9639 ( .A(n14961), .ZN(n12911) );
  INV_X1 U9640 ( .A(n11655), .ZN(n11653) );
  INV_X1 U9641 ( .A(n15051), .ZN(n12164) );
  INV_X1 U9642 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11752) );
  INV_X1 U9643 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9255) );
  INV_X1 U9644 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8190) );
  OR2_X1 U9645 ( .A1(n8663), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8674) );
  INV_X1 U9646 ( .A(n12623), .ZN(n12641) );
  OR2_X1 U9647 ( .A1(n8650), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8663) );
  INV_X1 U9648 ( .A(n8225), .ZN(n8228) );
  AND2_X1 U9649 ( .A1(n15711), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n13631) );
  INV_X1 U9650 ( .A(n13664), .ZN(n9817) );
  INV_X1 U9651 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n15272) );
  INV_X1 U9652 ( .A(n12703), .ZN(n15388) );
  INV_X1 U9653 ( .A(n12792), .ZN(n8742) );
  NOR2_X1 U9654 ( .A1(n8743), .A2(n10312), .ZN(n8866) );
  INV_X1 U9655 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10694) );
  OR2_X1 U9656 ( .A1(n12298), .A2(n14119), .ZN(n12300) );
  NAND2_X1 U9657 ( .A1(n12207), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n12298) );
  NAND2_X1 U9658 ( .A1(n11550), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n11728) );
  OR2_X1 U9659 ( .A1(n12274), .A2(n12394), .ZN(n12287) );
  AND2_X1 U9660 ( .A1(n9109), .A2(n9108), .ZN(n9652) );
  AND2_X1 U9661 ( .A1(n16119), .A2(n16120), .ZN(n12432) );
  INV_X1 U9662 ( .A(n10815), .ZN(n10816) );
  INV_X1 U9663 ( .A(n14651), .ZN(n12444) );
  NOR2_X1 U9664 ( .A1(n11042), .A2(n11041), .ZN(n11236) );
  OR2_X1 U9665 ( .A1(n12111), .A2(n11994), .ZN(n12134) );
  OR2_X1 U9666 ( .A1(n12093), .A2(n12092), .ZN(n12109) );
  INV_X1 U9667 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n11630) );
  INV_X1 U9668 ( .A(n14894), .ZN(n12103) );
  INV_X1 U9669 ( .A(n15097), .ZN(n14995) );
  NAND2_X1 U9670 ( .A1(n14884), .A2(n12164), .ZN(n14885) );
  INV_X1 U9671 ( .A(n14884), .ZN(n14897) );
  INV_X1 U9672 ( .A(n12993), .ZN(n13017) );
  NOR2_X1 U9673 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n8955) );
  NAND2_X1 U9674 ( .A1(n11353), .A2(SI_20_), .ZN(n11354) );
  OR2_X1 U9675 ( .A1(n10889), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n10891) );
  OR2_X1 U9676 ( .A1(n9374), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n9396) );
  INV_X1 U9677 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8937) );
  NOR2_X1 U9678 ( .A1(n15554), .A2(n15553), .ZN(n15555) );
  OAI21_X1 U9679 ( .B1(P3_ADDR_REG_15__SCAN_IN), .B2(n15609), .A(n15608), .ZN(
        n15616) );
  NAND2_X1 U9680 ( .A1(n8203), .A2(n15250), .ZN(n8705) );
  INV_X1 U9681 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8187) );
  INV_X1 U9682 ( .A(n13546), .ZN(n13519) );
  INV_X1 U9683 ( .A(n8889), .ZN(n8898) );
  OR2_X1 U9684 ( .A1(n13631), .A2(n13589), .ZN(n15720) );
  AND2_X1 U9685 ( .A1(n15711), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n13614) );
  OR2_X1 U9686 ( .A1(n8760), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n12198) );
  INV_X1 U9687 ( .A(n13564), .ZN(n13843) );
  AND2_X1 U9688 ( .A1(n12700), .A2(n12707), .ZN(n12696) );
  INV_X1 U9689 ( .A(n15886), .ZN(n13754) );
  AND2_X1 U9690 ( .A1(n9783), .A2(n13954), .ZN(n8758) );
  OR2_X1 U9691 ( .A1(n8884), .A2(n15293), .ZN(n8878) );
  OR2_X1 U9692 ( .A1(n8884), .A2(n15287), .ZN(n8658) );
  INV_X1 U9693 ( .A(n9782), .ZN(n8599) );
  INV_X1 U9694 ( .A(n11968), .ZN(n16078) );
  AND2_X1 U9695 ( .A1(n12670), .A2(n12671), .ZN(n12668) );
  NAND2_X1 U9696 ( .A1(n12623), .A2(n8742), .ZN(n16096) );
  OR2_X1 U9697 ( .A1(n10528), .A2(n12792), .ZN(n16097) );
  INV_X1 U9698 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n14018) );
  NAND2_X1 U9700 ( .A1(n8318), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8261) );
  AOI21_X1 U9701 ( .B1(n10335), .B2(n10334), .A(n8171), .ZN(n10342) );
  NAND2_X1 U9702 ( .A1(n11793), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n12248) );
  AOI22_X1 U9703 ( .A1(n9883), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n12234), .B2(
        n14204), .ZN(n9542) );
  AND2_X1 U9704 ( .A1(n13367), .A2(n14226), .ZN(n9571) );
  INV_X1 U9705 ( .A(n14082), .ZN(n14254) );
  OR2_X1 U9706 ( .A1(n11728), .A2(n11727), .ZN(n11795) );
  OR2_X1 U9707 ( .A1(n9491), .A2(n9490), .ZN(n9512) );
  AND2_X1 U9708 ( .A1(n9512), .A2(n14590), .ZN(n9494) );
  INV_X1 U9709 ( .A(n14175), .ZN(n14158) );
  INV_X1 U9710 ( .A(n13395), .ZN(n14340) );
  INV_X1 U9711 ( .A(n14180), .ZN(n14353) );
  OR2_X1 U9712 ( .A1(n9593), .A2(n9592), .ZN(n14356) );
  INV_X1 U9713 ( .A(n13398), .ZN(n14294) );
  INV_X1 U9714 ( .A(n9571), .ZN(n13407) );
  CLKBUF_X3 U9715 ( .A(n9772), .Z(n14416) );
  INV_X1 U9716 ( .A(n15905), .ZN(n16136) );
  XNOR2_X1 U9717 ( .A(n8936), .B(n9478), .ZN(n9544) );
  INV_X1 U9718 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n11429) );
  NAND2_X1 U9719 ( .A1(n10817), .A2(n10816), .ZN(n10818) );
  AND2_X1 U9720 ( .A1(n14682), .A2(n14679), .ZN(n12468) );
  OR2_X1 U9721 ( .A1(n12051), .A2(n12050), .ZN(n12063) );
  OR2_X1 U9722 ( .A1(n11002), .A2(n11482), .ZN(n11042) );
  OR2_X1 U9723 ( .A1(n9338), .A2(n13075), .ZN(n14725) );
  OR2_X1 U9724 ( .A1(n11631), .A2(n11630), .ZN(n11655) );
  INV_X1 U9725 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n15527) );
  INV_X1 U9726 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n15533) );
  INV_X1 U9727 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n11482) );
  INV_X1 U9728 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n14626) );
  AND2_X1 U9729 ( .A1(n15040), .A2(n14857), .ZN(n12540) );
  INV_X1 U9730 ( .A(n14881), .ZN(n14914) );
  OAI21_X1 U9731 ( .B1(n11670), .B2(n11669), .A(n11668), .ZN(n11877) );
  INV_X1 U9732 ( .A(n15990), .ZN(n16041) );
  INV_X1 U9733 ( .A(n13044), .ZN(n11444) );
  OR2_X1 U9734 ( .A1(n10538), .A2(n13059), .ZN(n15977) );
  INV_X1 U9735 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9082) );
  INV_X1 U9736 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n10892) );
  AND2_X1 U9737 ( .A1(n10888), .A2(n10440), .ZN(n10886) );
  OR2_X1 U9738 ( .A1(n8769), .A2(n8855), .ZN(n13548) );
  INV_X1 U9739 ( .A(n13554), .ZN(n13511) );
  NAND2_X1 U9740 ( .A1(n8779), .A2(n8778), .ZN(n13550) );
  AOI21_X1 U9741 ( .B1(n13686), .B2(n8887), .A(n8765), .ZN(n8896) );
  OR2_X1 U9742 ( .A1(n13614), .A2(n13588), .ZN(n15709) );
  INV_X1 U9743 ( .A(n15811), .ZN(n15775) );
  NAND2_X1 U9744 ( .A1(n9812), .A2(n13664), .ZN(n15822) );
  MUX2_X1 U9745 ( .A(n9812), .B(P3_U3897), .S(n12788), .Z(n15817) );
  INV_X1 U9746 ( .A(n13874), .ZN(n15881) );
  AND2_X1 U9747 ( .A1(n15899), .A2(n15898), .ZN(n13792) );
  AND2_X1 U9748 ( .A1(n15873), .A2(n8904), .ZN(n13959) );
  AND2_X1 U9749 ( .A1(n8981), .A2(n9116), .ZN(n9783) );
  AND2_X1 U9750 ( .A1(n8726), .A2(n8725), .ZN(n10312) );
  INV_X1 U9751 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8299) );
  INV_X1 U9752 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8309) );
  INV_X1 U9753 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8535) );
  OR3_X1 U9754 ( .A1(n14596), .A2(n14602), .A3(n14599), .ZN(n9545) );
  AND2_X1 U9755 ( .A1(n9597), .A2(n9596), .ZN(n14115) );
  AND2_X1 U9756 ( .A1(n9494), .A2(n9493), .ZN(n15477) );
  AND2_X1 U9757 ( .A1(n9494), .A2(n13408), .ZN(n15473) );
  INV_X1 U9758 ( .A(n12348), .ZN(n12349) );
  NAND2_X1 U9759 ( .A1(n15409), .A2(n9567), .ZN(n14430) );
  AND2_X1 U9760 ( .A1(n10516), .A2(n14226), .ZN(n14438) );
  NAND2_X1 U9761 ( .A1(n9977), .A2(n13358), .ZN(n14393) );
  AND2_X1 U9762 ( .A1(n7190), .A2(n13407), .ZN(n15905) );
  INV_X1 U9763 ( .A(n16106), .ZN(n16092) );
  NOR2_X1 U9764 ( .A1(n15173), .A2(n9993), .ZN(n10136) );
  NAND2_X1 U9765 ( .A1(n8930), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8932) );
  AND2_X1 U9766 ( .A1(n11097), .A2(n10983), .ZN(n11767) );
  AND2_X1 U9767 ( .A1(n10080), .A2(n10537), .ZN(n15921) );
  INV_X1 U9768 ( .A(n14725), .ZN(n15927) );
  OR2_X1 U9769 ( .A1(n13002), .A2(n15151), .ZN(n15003) );
  OR2_X1 U9770 ( .A1(n12168), .A2(n12142), .ZN(n12141) );
  AND2_X1 U9771 ( .A1(n12033), .A2(n12032), .ZN(n14637) );
  AND2_X1 U9772 ( .A1(n10130), .A2(n10129), .ZN(n10210) );
  INV_X1 U9773 ( .A(n14828), .ZN(n14787) );
  AND2_X1 U9774 ( .A1(n9125), .A2(n15154), .ZN(n14834) );
  INV_X1 U9775 ( .A(n14829), .ZN(n14833) );
  NAND2_X1 U9776 ( .A1(n12150), .A2(n12149), .ZN(n12151) );
  INV_X1 U9777 ( .A(n13052), .ZN(n14947) );
  INV_X1 U9778 ( .A(n15005), .ZN(n14980) );
  AND2_X1 U9779 ( .A1(n10537), .A2(n10536), .ZN(n16037) );
  AOI21_X1 U9780 ( .B1(n9432), .B2(n9330), .A(n9329), .ZN(n10534) );
  INV_X1 U9781 ( .A(n15955), .ZN(n16060) );
  INV_X1 U9782 ( .A(n15933), .ZN(n16064) );
  NAND2_X1 U9783 ( .A1(n12799), .A2(n9425), .ZN(n15955) );
  AND3_X1 U9784 ( .A1(n9435), .A2(n9434), .A3(n9433), .ZN(n10289) );
  AND2_X1 U9785 ( .A1(n9787), .A2(n9786), .ZN(n15771) );
  INV_X1 U9786 ( .A(n13527), .ZN(n13539) );
  INV_X1 U9787 ( .A(n13550), .ZN(n13531) );
  AND2_X1 U9788 ( .A1(n12581), .A2(n8894), .ZN(n13681) );
  INV_X1 U9789 ( .A(n13876), .ZN(n13566) );
  OR2_X1 U9790 ( .A1(n8981), .A2(n14016), .ZN(n13577) );
  AND4_X1 U9791 ( .A1(n15689), .A2(n15688), .A3(n15687), .A4(n15686), .ZN(
        n15691) );
  NAND2_X1 U9792 ( .A1(n9812), .A2(n9811), .ZN(n15825) );
  INV_X1 U9793 ( .A(n13792), .ZN(n15402) );
  NAND2_X1 U9794 ( .A1(n16101), .A2(n13954), .ZN(n16154) );
  AND2_X2 U9795 ( .A1(n10316), .A2(n8921), .ZN(n16101) );
  INV_X1 U9796 ( .A(n13514), .ZN(n13999) );
  NAND2_X1 U9797 ( .A1(n16104), .A2(n13954), .ZN(n16159) );
  AND2_X2 U9798 ( .A1(n8869), .A2(n9783), .ZN(n16104) );
  AND2_X1 U9799 ( .A1(n8775), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9116) );
  INV_X1 U9800 ( .A(SI_17_), .ZN(n15205) );
  INV_X1 U9801 ( .A(SI_12_), .ZN(n15319) );
  NOR2_X1 U9802 ( .A1(n9545), .A2(n11753), .ZN(n9491) );
  AND2_X1 U9803 ( .A1(n9568), .A2(n14430), .ZN(n14162) );
  NAND2_X1 U9804 ( .A1(n12320), .A2(n12319), .ZN(n14173) );
  OR2_X1 U9805 ( .A1(n15469), .A2(P2_U3088), .ZN(n15466) );
  INV_X1 U9806 ( .A(n14438), .ZN(n14420) );
  AND3_X1 U9807 ( .A1(n11738), .A2(n11737), .A3(n11736), .ZN(n14532) );
  INV_X1 U9808 ( .A(n16142), .ZN(n16141) );
  INV_X1 U9809 ( .A(n14361), .ZN(n14562) );
  INV_X1 U9810 ( .A(n16146), .ZN(n16143) );
  OR2_X1 U9811 ( .A1(n15406), .A2(n15176), .ZN(n15177) );
  INV_X1 U9812 ( .A(n15409), .ZN(n15406) );
  XNOR2_X1 U9813 ( .A(n8932), .B(n8931), .ZN(n14596) );
  INV_X1 U9814 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11264) );
  INV_X1 U9815 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9644) );
  INV_X1 U9816 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9018) );
  INV_X1 U9817 ( .A(n14842), .ZN(n14797) );
  NAND2_X1 U9818 ( .A1(n10081), .A2(P1_STATE_REG_SCAN_IN), .ZN(n16133) );
  OR2_X1 U9819 ( .A1(n9338), .A2(n9332), .ZN(n16123) );
  INV_X1 U9820 ( .A(n16129), .ZN(n14731) );
  NAND2_X1 U9821 ( .A1(n12117), .A2(n12116), .ZN(n14899) );
  OR2_X1 U9822 ( .A1(n9166), .A2(n14769), .ZN(n14828) );
  INV_X1 U9823 ( .A(n11899), .ZN(n15998) );
  AND2_X1 U9824 ( .A1(n12167), .A2(n15016), .ZN(n16047) );
  INV_X1 U9825 ( .A(n16067), .ZN(n16066) );
  INV_X1 U9826 ( .A(n16071), .ZN(n16068) );
  AND2_X2 U9827 ( .A1(n10290), .A2(n10289), .ZN(n16071) );
  NOR2_X1 U9828 ( .A1(n15165), .A2(n9097), .ZN(n9329) );
  INV_X1 U9829 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11096) );
  INV_X1 U9830 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9646) );
  INV_X1 U9831 ( .A(P2_RD_REG_SCAN_IN), .ZN(n15829) );
  INV_X2 U9832 ( .A(n13577), .ZN(P3_U3897) );
  OR4_X1 U9833 ( .A1(n8980), .A2(n8979), .A3(n8978), .A4(n8977), .ZN(P3_U3176)
         );
  AND2_X1 U9834 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9491), .ZN(P2_U3947) );
  INV_X1 U9835 ( .A(n14752), .ZN(P1_U4016) );
  INV_X2 U9836 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NAND2_X1 U9837 ( .A1(n9857), .A2(n15365), .ZN(n8439) );
  INV_X1 U9838 ( .A(n8439), .ZN(n8188) );
  NAND2_X1 U9839 ( .A1(n8188), .A2(n8187), .ZN(n8441) );
  INV_X1 U9840 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8198) );
  INV_X1 U9841 ( .A(n8626), .ZN(n8200) );
  INV_X1 U9842 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n8201) );
  INV_X1 U9843 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n15250) );
  INV_X1 U9844 ( .A(n8707), .ZN(n8205) );
  INV_X1 U9845 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8204) );
  NAND2_X1 U9846 ( .A1(n8205), .A2(n8204), .ZN(n8760) );
  NAND2_X1 U9847 ( .A1(n8707), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8206) );
  NAND2_X1 U9848 ( .A1(n8760), .A2(n8206), .ZN(n13692) );
  XNOR2_X2 U9849 ( .A(n8224), .B(n8223), .ZN(n8225) );
  NAND2_X1 U9850 ( .A1(n13692), .A2(n8887), .ZN(n8234) );
  NAND2_X4 U9851 ( .A1(n8226), .A2(n8225), .ZN(n12577) );
  INV_X1 U9852 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n8231) );
  NAND2_X1 U9853 ( .A1(n12573), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8230) );
  NAND2_X1 U9854 ( .A1(n8898), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8229) );
  OAI211_X1 U9855 ( .C1(n12577), .C2(n8231), .A(n8230), .B(n8229), .ZN(n8232)
         );
  INV_X1 U9856 ( .A(n8232), .ZN(n8233) );
  INV_X1 U9857 ( .A(n8403), .ZN(n8235) );
  NAND2_X1 U9858 ( .A1(n8236), .A2(n8235), .ZN(n8392) );
  NAND2_X1 U9859 ( .A1(n9006), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8237) );
  INV_X1 U9860 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9058) );
  NAND2_X1 U9861 ( .A1(n9058), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8238) );
  INV_X1 U9862 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9000) );
  NAND2_X1 U9863 ( .A1(n9094), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8240) );
  XNOR2_X1 U9864 ( .A(n9038), .B(P1_DATAO_REG_4__SCAN_IN), .ZN(n8415) );
  INV_X1 U9865 ( .A(n8415), .ZN(n8241) );
  NAND2_X1 U9866 ( .A1(n8416), .A2(n8241), .ZN(n8243) );
  NAND2_X1 U9867 ( .A1(n9038), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8242) );
  XNOR2_X1 U9868 ( .A(n8245), .B(P1_DATAO_REG_5__SCAN_IN), .ZN(n8431) );
  INV_X1 U9869 ( .A(n8431), .ZN(n8244) );
  NAND2_X1 U9870 ( .A1(n8245), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8246) );
  NAND2_X1 U9871 ( .A1(n9110), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8249) );
  NAND2_X1 U9872 ( .A1(n9114), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8247) );
  INV_X1 U9873 ( .A(n8366), .ZN(n8248) );
  NAND2_X1 U9874 ( .A1(n8465), .A2(n8464), .ZN(n8251) );
  NAND2_X1 U9875 ( .A1(n9180), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8250) );
  XNOR2_X1 U9876 ( .A(n9360), .B(P1_DATAO_REG_9__SCAN_IN), .ZN(n8350) );
  INV_X1 U9877 ( .A(n8350), .ZN(n8252) );
  NAND2_X1 U9878 ( .A1(n8351), .A2(n8252), .ZN(n8254) );
  NAND2_X1 U9879 ( .A1(n9360), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8253) );
  XNOR2_X1 U9880 ( .A(n9443), .B(P1_DATAO_REG_10__SCAN_IN), .ZN(n8338) );
  INV_X1 U9881 ( .A(n8338), .ZN(n8255) );
  NAND2_X1 U9882 ( .A1(n9443), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8256) );
  XNOR2_X1 U9883 ( .A(n9644), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n8496) );
  INV_X1 U9884 ( .A(n8496), .ZN(n8257) );
  NAND2_X1 U9885 ( .A1(n9646), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8258) );
  XNOR2_X1 U9886 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n8509) );
  INV_X1 U9887 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10029) );
  NAND2_X1 U9888 ( .A1(n8259), .A2(n10029), .ZN(n8260) );
  XNOR2_X1 U9889 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8520) );
  NAND2_X1 U9890 ( .A1(n10304), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8262) );
  XNOR2_X1 U9891 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n8533) );
  INV_X1 U9892 ( .A(n8552), .ZN(n8263) );
  NAND2_X1 U9893 ( .A1(n8263), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8266) );
  NAND2_X1 U9894 ( .A1(n8264), .A2(n10895), .ZN(n8265) );
  XNOR2_X1 U9895 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .ZN(n8567) );
  NAND2_X1 U9896 ( .A1(n11096), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8267) );
  XNOR2_X1 U9897 ( .A(n8269), .B(P1_DATAO_REG_18__SCAN_IN), .ZN(n8583) );
  INV_X1 U9898 ( .A(n8583), .ZN(n8268) );
  NOR2_X1 U9899 ( .A1(n11264), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8270) );
  NAND2_X1 U9900 ( .A1(n11264), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8271) );
  XNOR2_X1 U9901 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .ZN(n8611) );
  INV_X1 U9902 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11349) );
  NAND2_X1 U9903 ( .A1(n11349), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8272) );
  INV_X1 U9904 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11355) );
  NAND2_X1 U9905 ( .A1(n11355), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8275) );
  INV_X1 U9906 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11357) );
  NAND2_X1 U9907 ( .A1(n11357), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8274) );
  NAND2_X1 U9908 ( .A1(n8275), .A2(n8274), .ZN(n8620) );
  INV_X1 U9909 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n11571) );
  XNOR2_X1 U9910 ( .A(n11571), .B(P1_DATAO_REG_22__SCAN_IN), .ZN(n8637) );
  INV_X1 U9911 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11577) );
  NAND2_X1 U9912 ( .A1(n11577), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8276) );
  XNOR2_X1 U9913 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8656) );
  NAND2_X1 U9914 ( .A1(n11752), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8277) );
  NAND2_X1 U9915 ( .A1(n8279), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8280) );
  INV_X1 U9916 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n14603) );
  INV_X1 U9917 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n15163) );
  NAND2_X1 U9918 ( .A1(n15163), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8283) );
  INV_X1 U9919 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n14600) );
  NAND2_X1 U9920 ( .A1(n14600), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8282) );
  AND2_X1 U9921 ( .A1(n8283), .A2(n8282), .ZN(n8685) );
  INV_X1 U9922 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15158) );
  NAND2_X1 U9923 ( .A1(n15158), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8285) );
  INV_X1 U9924 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14595) );
  NAND2_X1 U9925 ( .A1(n14595), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8284) );
  AND2_X1 U9926 ( .A1(n8285), .A2(n8284), .ZN(n8714) );
  INV_X1 U9927 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15156) );
  NAND2_X1 U9928 ( .A1(n15156), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8872) );
  INV_X1 U9929 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n12369) );
  NAND2_X1 U9930 ( .A1(n12369), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8286) );
  AND2_X1 U9931 ( .A1(n8872), .A2(n8286), .ZN(n8287) );
  OR2_X1 U9932 ( .A1(n8288), .A2(n8287), .ZN(n8289) );
  NAND2_X1 U9933 ( .A1(n8873), .A2(n8289), .ZN(n11828) );
  NAND2_X4 U9934 ( .A1(n12193), .A2(n8767), .ZN(n9782) );
  NAND2_X1 U9935 ( .A1(n9782), .A2(n7178), .ZN(n8394) );
  NAND2_X1 U9936 ( .A1(n9782), .A2(n9540), .ZN(n8390) );
  INV_X1 U9937 ( .A(SI_27_), .ZN(n15297) );
  NAND2_X1 U9938 ( .A1(n7290), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8296) );
  MUX2_X1 U9939 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8296), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n8297) );
  NAND2_X1 U9940 ( .A1(n8754), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8300) );
  XNOR2_X1 U9941 ( .A(n11452), .B(P3_B_REG_SCAN_IN), .ZN(n8303) );
  NAND2_X1 U9942 ( .A1(n7253), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8302) );
  NAND2_X1 U9943 ( .A1(n8303), .A2(n11590), .ZN(n8304) );
  INV_X1 U9944 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8305) );
  NAND2_X1 U9945 ( .A1(n9220), .A2(n8305), .ZN(n8307) );
  NAND2_X1 U9946 ( .A1(n11758), .A2(n11452), .ZN(n8306) );
  NAND2_X1 U9947 ( .A1(n8311), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8312) );
  MUX2_X1 U9948 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8312), .S(
        P3_IR_REG_19__SCAN_IN), .Z(n8313) );
  MUX2_X1 U9949 ( .A(n12596), .B(n10528), .S(n12623), .Z(n8317) );
  NAND2_X2 U9950 ( .A1(n14017), .A2(n8317), .ZN(n8410) );
  INV_X4 U9951 ( .A(n13084), .ZN(n8720) );
  XNOR2_X1 U9952 ( .A(n8786), .B(n8720), .ZN(n13090) );
  NOR2_X1 U9953 ( .A1(n13090), .A2(n13698), .ZN(n13086) );
  AOI21_X1 U9954 ( .B1(n13698), .B2(n13090), .A(n13086), .ZN(n8724) );
  XNOR2_X1 U9955 ( .A(n8318), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n9253) );
  NAND2_X1 U9956 ( .A1(n9253), .A2(n12584), .ZN(n8324) );
  INV_X1 U9957 ( .A(n8884), .ZN(n8600) );
  NOR2_X1 U9958 ( .A1(n8433), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8362) );
  NAND2_X1 U9959 ( .A1(n8362), .A2(n8319), .ZN(n8452) );
  INV_X1 U9960 ( .A(n8320), .ZN(n8321) );
  OAI21_X1 U9961 ( .B1(n8452), .B2(n8321), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8322) );
  XNOR2_X1 U9962 ( .A(n8322), .B(P3_IR_REG_13__SCAN_IN), .ZN(n15739) );
  INV_X1 U9963 ( .A(n15739), .ZN(n9254) );
  AOI22_X1 U9964 ( .A1(n8600), .A2(n15311), .B1(n8599), .B2(n9254), .ZN(n8323)
         );
  NAND2_X1 U9965 ( .A1(n8324), .A2(n8323), .ZN(n16095) );
  XNOR2_X1 U9966 ( .A(n16095), .B(n8720), .ZN(n8517) );
  INV_X1 U9967 ( .A(n8517), .ZN(n8519) );
  NAND2_X1 U9968 ( .A1(n12573), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8331) );
  INV_X1 U9969 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n8325) );
  OR2_X1 U9970 ( .A1(n8889), .A2(n8325), .ZN(n8330) );
  NAND2_X1 U9971 ( .A1(n8504), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8326) );
  AND2_X1 U9972 ( .A1(n8527), .A2(n8326), .ZN(n15397) );
  OR2_X1 U9973 ( .A1(n8590), .A2(n15397), .ZN(n8329) );
  INV_X1 U9974 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n8327) );
  OR2_X1 U9975 ( .A1(n12577), .A2(n8327), .ZN(n8328) );
  NAND2_X1 U9976 ( .A1(n12573), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8337) );
  INV_X1 U9977 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n8332) );
  OR2_X1 U9978 ( .A1(n8889), .A2(n8332), .ZN(n8336) );
  NAND2_X1 U9979 ( .A1(n8345), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8333) );
  AND2_X1 U9980 ( .A1(n8485), .A2(n8333), .ZN(n11876) );
  OR2_X1 U9981 ( .A1(n8590), .A2(n11876), .ZN(n8335) );
  INV_X1 U9982 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11700) );
  OR2_X1 U9983 ( .A1(n12577), .A2(n11700), .ZN(n8334) );
  XNOR2_X1 U9984 ( .A(n8339), .B(n8338), .ZN(n9042) );
  OR2_X1 U9985 ( .A1(n8689), .A2(n9042), .ZN(n8343) );
  OR2_X1 U9986 ( .A1(n8884), .A2(SI_10_), .ZN(n8342) );
  OR2_X1 U9987 ( .A1(n8493), .A2(n8221), .ZN(n8340) );
  INV_X1 U9988 ( .A(n13628), .ZN(n13580) );
  OR2_X1 U9989 ( .A1(n9782), .A2(n13580), .ZN(n8341) );
  XNOR2_X1 U9990 ( .A(n13953), .B(n8720), .ZN(n8483) );
  INV_X1 U9991 ( .A(n8483), .ZN(n8484) );
  NAND2_X1 U9992 ( .A1(n12573), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8349) );
  INV_X1 U9993 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11319) );
  OR2_X1 U9994 ( .A1(n8889), .A2(n11319), .ZN(n8348) );
  NAND2_X1 U9995 ( .A1(n8474), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n8344) );
  AND2_X1 U9996 ( .A1(n8345), .A2(n8344), .ZN(n11608) );
  OR2_X1 U9997 ( .A1(n8590), .A2(n11608), .ZN(n8347) );
  INV_X1 U9998 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11320) );
  OR2_X1 U9999 ( .A1(n12577), .A2(n11320), .ZN(n8346) );
  NAND4_X1 U10000 ( .A1(n8349), .A2(n8348), .A3(n8347), .A4(n8346), .ZN(n13570) );
  INV_X1 U10001 ( .A(n13570), .ZN(n11693) );
  XNOR2_X1 U10002 ( .A(n8351), .B(n8350), .ZN(n9027) );
  OR2_X1 U10003 ( .A1(n8689), .A2(n9027), .ZN(n8356) );
  OR2_X1 U10004 ( .A1(n8884), .A2(SI_9_), .ZN(n8355) );
  NAND2_X1 U10005 ( .A1(n8352), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8353) );
  XNOR2_X1 U10006 ( .A(n8353), .B(P3_IR_REG_9__SCAN_IN), .ZN(n15685) );
  OR2_X1 U10007 ( .A1(n9782), .A2(n15685), .ZN(n8354) );
  XNOR2_X1 U10008 ( .A(n8822), .B(n8720), .ZN(n8481) );
  INV_X1 U10009 ( .A(n8481), .ZN(n8482) );
  NAND2_X1 U10010 ( .A1(n8438), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8361) );
  INV_X1 U10011 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10179) );
  OR2_X1 U10012 ( .A1(n12577), .A2(n10179), .ZN(n8360) );
  NAND2_X1 U10013 ( .A1(n8441), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8357) );
  AND2_X1 U10014 ( .A1(n8457), .A2(n8357), .ZN(n11290) );
  OR2_X1 U10015 ( .A1(n8590), .A2(n11290), .ZN(n8359) );
  INV_X1 U10016 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10178) );
  OR2_X1 U10017 ( .A1(n8556), .A2(n10178), .ZN(n8358) );
  NOR2_X1 U10018 ( .A1(n8362), .A2(n8221), .ZN(n8363) );
  MUX2_X1 U10019 ( .A(n8221), .B(n8363), .S(P3_IR_REG_6__SCAN_IN), .Z(n8365)
         );
  INV_X1 U10020 ( .A(n8452), .ZN(n8364) );
  INV_X1 U10021 ( .A(SI_6_), .ZN(n8982) );
  OR2_X1 U10022 ( .A1(n8884), .A2(n8982), .ZN(n8369) );
  XNOR2_X1 U10023 ( .A(n8367), .B(n8366), .ZN(n8983) );
  OR2_X1 U10024 ( .A1(n8689), .A2(n8983), .ZN(n8368) );
  OAI211_X1 U10025 ( .C1(n9782), .C2(n10772), .A(n8369), .B(n8368), .ZN(n11211) );
  XNOR2_X1 U10026 ( .A(n11211), .B(n8720), .ZN(n8447) );
  INV_X1 U10027 ( .A(n8447), .ZN(n8449) );
  NAND2_X1 U10028 ( .A1(n8438), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8373) );
  INV_X1 U10029 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n9833) );
  OR2_X1 U10030 ( .A1(n12577), .A2(n9833), .ZN(n8372) );
  INV_X1 U10031 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n9832) );
  OR2_X1 U10032 ( .A1(n8556), .A2(n9832), .ZN(n8371) );
  OR2_X1 U10033 ( .A1(n8590), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8370) );
  AND4_X2 U10034 ( .A1(n8373), .A2(n8372), .A3(n8371), .A4(n8370), .ZN(n10988)
         );
  OR2_X1 U10035 ( .A1(n8884), .A2(SI_3_), .ZN(n8379) );
  XNOR2_X1 U10036 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8374) );
  XNOR2_X1 U10037 ( .A(n8375), .B(n8374), .ZN(n9019) );
  OR2_X1 U10038 ( .A1(n8689), .A2(n9019), .ZN(n8378) );
  NAND2_X1 U10039 ( .A1(n8376), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8418) );
  XNOR2_X1 U10040 ( .A(n8418), .B(P3_IR_REG_3__SCAN_IN), .ZN(n9834) );
  OR2_X1 U10041 ( .A1(n9782), .A2(n9834), .ZN(n8377) );
  AND3_X2 U10042 ( .A1(n8379), .A2(n8378), .A3(n8377), .ZN(n10639) );
  XNOR2_X1 U10043 ( .A(n10639), .B(n8720), .ZN(n8414) );
  NAND2_X1 U10044 ( .A1(n8438), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8383) );
  INV_X1 U10045 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n9826) );
  OR2_X1 U10046 ( .A1(n12577), .A2(n9826), .ZN(n8382) );
  INV_X1 U10047 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9825) );
  INV_X1 U10048 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15891) );
  OR2_X1 U10049 ( .A1(n8405), .A2(n15891), .ZN(n8380) );
  OR2_X1 U10050 ( .A1(n8884), .A2(SI_2_), .ZN(n8389) );
  XNOR2_X1 U10051 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8384) );
  XNOR2_X1 U10052 ( .A(n8385), .B(n8384), .ZN(n9029) );
  OR2_X1 U10053 ( .A1(n8689), .A2(n9029), .ZN(n8388) );
  OR2_X1 U10054 ( .A1(n9782), .A2(n9827), .ZN(n8387) );
  AND3_X2 U10055 ( .A1(n8389), .A2(n8388), .A3(n8387), .ZN(n8788) );
  XNOR2_X1 U10056 ( .A(n8788), .B(n8410), .ZN(n8412) );
  INV_X1 U10057 ( .A(n8412), .ZN(n8413) );
  INV_X1 U10058 ( .A(SI_1_), .ZN(n8991) );
  OR2_X1 U10059 ( .A1(n8390), .A2(n8991), .ZN(n8396) );
  NAND2_X1 U10060 ( .A1(n8391), .A2(n8403), .ZN(n8393) );
  AND2_X1 U10061 ( .A1(n8393), .A2(n8392), .ZN(n8984) );
  OAI211_X1 U10062 ( .C1(n9782), .C2(n9932), .A(n8396), .B(n8395), .ZN(n10524)
         );
  XNOR2_X1 U10063 ( .A(n8787), .B(n8410), .ZN(n8401) );
  NAND2_X1 U10064 ( .A1(n8438), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8400) );
  INV_X1 U10065 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10527) );
  OR2_X1 U10066 ( .A1(n12577), .A2(n10527), .ZN(n8399) );
  INV_X1 U10067 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n9818) );
  INV_X1 U10068 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10168) );
  OR2_X1 U10069 ( .A1(n8405), .A2(n10168), .ZN(n8397) );
  NAND2_X1 U10070 ( .A1(n8401), .A2(n9769), .ZN(n8411) );
  OAI21_X1 U10071 ( .B1(n8401), .B2(n9769), .A(n8411), .ZN(n10166) );
  INV_X1 U10072 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9296) );
  NAND2_X1 U10073 ( .A1(n9296), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8402) );
  AND2_X1 U10074 ( .A1(n8403), .A2(n8402), .ZN(n8404) );
  NAND2_X1 U10075 ( .A1(n9540), .A2(SI_0_), .ZN(n9626) );
  OAI21_X1 U10076 ( .B1(n9540), .B2(n8404), .A(n9626), .ZN(n14025) );
  MUX2_X1 U10077 ( .A(P3_IR_REG_0__SCAN_IN), .B(n14025), .S(n9782), .Z(n10319)
         );
  NAND2_X1 U10078 ( .A1(n8438), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8409) );
  INV_X1 U10079 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n9823) );
  OR2_X1 U10080 ( .A1(n8556), .A2(n9823), .ZN(n8408) );
  INV_X1 U10081 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n9824) );
  OR2_X1 U10082 ( .A1(n12577), .A2(n9824), .ZN(n8407) );
  INV_X1 U10083 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n15658) );
  OR2_X1 U10084 ( .A1(n8405), .A2(n15658), .ZN(n8406) );
  NAND2_X1 U10085 ( .A1(n13578), .A2(n10319), .ZN(n10421) );
  OAI21_X1 U10086 ( .B1(n10319), .B2(n8410), .A(n10421), .ZN(n10167) );
  INV_X1 U10087 ( .A(n10636), .ZN(n13576) );
  XNOR2_X1 U10088 ( .A(n13576), .B(n8412), .ZN(n10396) );
  XNOR2_X1 U10089 ( .A(n8414), .B(n10988), .ZN(n10634) );
  NAND2_X1 U10090 ( .A1(n10635), .A2(n10634), .ZN(n10633) );
  OR2_X1 U10091 ( .A1(n8884), .A2(SI_4_), .ZN(n8423) );
  XNOR2_X1 U10092 ( .A(n8416), .B(n8415), .ZN(n9023) );
  OR2_X1 U10093 ( .A1(n8689), .A2(n9023), .ZN(n8422) );
  NAND2_X1 U10094 ( .A1(n8418), .A2(n8417), .ZN(n8419) );
  NAND2_X1 U10095 ( .A1(n8419), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8420) );
  OR2_X1 U10096 ( .A1(n9782), .A2(n10151), .ZN(n8421) );
  XNOR2_X1 U10097 ( .A(n11061), .B(n8410), .ZN(n8429) );
  NAND2_X1 U10098 ( .A1(n8438), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8428) );
  INV_X1 U10099 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11028) );
  OR2_X1 U10100 ( .A1(n12577), .A2(n11028), .ZN(n8427) );
  NAND2_X1 U10101 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8424) );
  AND2_X1 U10102 ( .A1(n8439), .A2(n8424), .ZN(n10991) );
  OR2_X1 U10103 ( .A1(n8590), .A2(n10991), .ZN(n8426) );
  INV_X1 U10104 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10147) );
  OR2_X1 U10105 ( .A1(n8556), .A2(n10147), .ZN(n8425) );
  NAND2_X1 U10106 ( .A1(n8429), .A2(n11113), .ZN(n8430) );
  OAI21_X1 U10107 ( .B1(n8429), .B2(n11113), .A(n8430), .ZN(n10986) );
  INV_X1 U10108 ( .A(n8430), .ZN(n11110) );
  OR2_X1 U10109 ( .A1(n8884), .A2(SI_5_), .ZN(n8437) );
  XNOR2_X1 U10110 ( .A(n8432), .B(n8431), .ZN(n9021) );
  OR2_X1 U10111 ( .A1(n8689), .A2(n9021), .ZN(n8436) );
  NAND2_X1 U10112 ( .A1(n8433), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8434) );
  XNOR2_X1 U10113 ( .A(n8434), .B(P3_IR_REG_5__SCAN_IN), .ZN(n10174) );
  OR2_X1 U10114 ( .A1(n9782), .A2(n10174), .ZN(n8435) );
  XNOR2_X1 U10115 ( .A(n11116), .B(n13084), .ZN(n8448) );
  NAND2_X1 U10116 ( .A1(n8438), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8446) );
  INV_X1 U10117 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n11280) );
  OR2_X1 U10118 ( .A1(n8889), .A2(n11280), .ZN(n8445) );
  NAND2_X1 U10119 ( .A1(n8439), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8440) );
  AND2_X1 U10120 ( .A1(n8441), .A2(n8440), .ZN(n11119) );
  OR2_X1 U10121 ( .A1(n8590), .A2(n11119), .ZN(n8444) );
  INV_X1 U10122 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n8442) );
  OR2_X1 U10123 ( .A1(n12577), .A2(n8442), .ZN(n8443) );
  NAND4_X1 U10124 ( .A1(n8446), .A2(n8445), .A3(n8444), .A4(n8443), .ZN(n13574) );
  XNOR2_X1 U10125 ( .A(n8448), .B(n13574), .ZN(n11109) );
  XNOR2_X1 U10126 ( .A(n11596), .B(n8447), .ZN(n11206) );
  INV_X1 U10127 ( .A(n13574), .ZN(n11208) );
  NAND2_X1 U10128 ( .A1(n8448), .A2(n11208), .ZN(n11203) );
  OAI21_X1 U10129 ( .B1(n11596), .B2(n8449), .A(n11205), .ZN(n11393) );
  OR2_X1 U10130 ( .A1(n8884), .A2(SI_7_), .ZN(n8456) );
  XNOR2_X1 U10131 ( .A(n8451), .B(n8450), .ZN(n9025) );
  OR2_X1 U10132 ( .A1(n8689), .A2(n9025), .ZN(n8455) );
  NAND2_X1 U10133 ( .A1(n8452), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8453) );
  OR2_X1 U10134 ( .A1(n9782), .A2(n15672), .ZN(n8454) );
  XNOR2_X1 U10135 ( .A(n11397), .B(n8720), .ZN(n8463) );
  NAND2_X1 U10136 ( .A1(n12573), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8462) );
  INV_X1 U10137 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n10760) );
  OR2_X1 U10138 ( .A1(n8889), .A2(n10760), .ZN(n8461) );
  NAND2_X1 U10139 ( .A1(n8457), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8458) );
  AND2_X1 U10140 ( .A1(n8472), .A2(n8458), .ZN(n11593) );
  OR2_X1 U10141 ( .A1(n8590), .A2(n11593), .ZN(n8460) );
  INV_X1 U10142 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10761) );
  OR2_X1 U10143 ( .A1(n12577), .A2(n10761), .ZN(n8459) );
  XNOR2_X1 U10144 ( .A(n8463), .B(n11469), .ZN(n11394) );
  XNOR2_X1 U10145 ( .A(n8465), .B(n8464), .ZN(n8985) );
  OR2_X1 U10146 ( .A1(n8689), .A2(n8985), .ZN(n8470) );
  INV_X1 U10147 ( .A(SI_8_), .ZN(n8986) );
  OR2_X1 U10148 ( .A1(n8884), .A2(n8986), .ZN(n8469) );
  NAND2_X1 U10149 ( .A1(n8466), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8467) );
  XNOR2_X1 U10150 ( .A(n8467), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11315) );
  OR2_X1 U10151 ( .A1(n9782), .A2(n11328), .ZN(n8468) );
  XNOR2_X1 U10152 ( .A(n16005), .B(n8720), .ZN(n8480) );
  NAND2_X1 U10153 ( .A1(n12573), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8479) );
  INV_X1 U10154 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n8471) );
  OR2_X1 U10155 ( .A1(n8556), .A2(n8471), .ZN(n8478) );
  NAND2_X1 U10156 ( .A1(n8472), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8473) );
  AND2_X1 U10157 ( .A1(n8474), .A2(n8473), .ZN(n11474) );
  OR2_X1 U10158 ( .A1(n8590), .A2(n11474), .ZN(n8477) );
  INV_X1 U10159 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n8475) );
  OR2_X1 U10160 ( .A1(n12577), .A2(n8475), .ZN(n8476) );
  XNOR2_X1 U10161 ( .A(n8480), .B(n12687), .ZN(n11467) );
  XNOR2_X1 U10162 ( .A(n8481), .B(n13570), .ZN(n11605) );
  XNOR2_X1 U10163 ( .A(n8483), .B(n11859), .ZN(n11869) );
  OAI21_X1 U10164 ( .B1(n11859), .B2(n8484), .A(n11868), .ZN(n8973) );
  NAND2_X1 U10165 ( .A1(n12573), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8491) );
  INV_X1 U10166 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11863) );
  OR2_X1 U10167 ( .A1(n12577), .A2(n11863), .ZN(n8490) );
  NAND2_X1 U10168 ( .A1(n8485), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8486) );
  AND2_X1 U10169 ( .A1(n8502), .A2(n8486), .ZN(n11862) );
  OR2_X1 U10170 ( .A1(n8590), .A2(n11862), .ZN(n8489) );
  INV_X1 U10171 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n8487) );
  OR2_X1 U10172 ( .A1(n8889), .A2(n8487), .ZN(n8488) );
  NAND2_X1 U10173 ( .A1(n8493), .A2(n8492), .ZN(n8511) );
  NAND2_X1 U10174 ( .A1(n8511), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8495) );
  INV_X1 U10175 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8494) );
  XNOR2_X1 U10176 ( .A(n8495), .B(n8494), .ZN(n13613) );
  XNOR2_X1 U10177 ( .A(n8497), .B(n8496), .ZN(n9118) );
  OR2_X1 U10178 ( .A1(n9118), .A2(n8689), .ZN(n8499) );
  OR2_X1 U10179 ( .A1(n8884), .A2(SI_11_), .ZN(n8498) );
  OAI211_X1 U10180 ( .C1(n15697), .C2(n9782), .A(n8499), .B(n8498), .ZN(n11947) );
  XNOR2_X1 U10181 ( .A(n11947), .B(n8720), .ZN(n8500) );
  XNOR2_X1 U10182 ( .A(n13568), .B(n8500), .ZN(n8972) );
  INV_X1 U10183 ( .A(n8500), .ZN(n8501) );
  NAND2_X1 U10184 ( .A1(n12573), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8508) );
  INV_X1 U10185 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n16083) );
  OR2_X1 U10186 ( .A1(n8556), .A2(n16083), .ZN(n8507) );
  NAND2_X1 U10187 ( .A1(n8502), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8503) );
  AND2_X1 U10188 ( .A1(n8504), .A2(n8503), .ZN(n11965) );
  OR2_X1 U10189 ( .A1(n8590), .A2(n11965), .ZN(n8506) );
  INV_X1 U10190 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11966) );
  OR2_X1 U10191 ( .A1(n12577), .A2(n11966), .ZN(n8505) );
  NAND4_X1 U10192 ( .A1(n8508), .A2(n8507), .A3(n8506), .A4(n8505), .ZN(n13567) );
  XNOR2_X1 U10193 ( .A(n8510), .B(n8509), .ZN(n9120) );
  NAND2_X1 U10194 ( .A1(n9120), .A2(n12584), .ZN(n8515) );
  OAI21_X1 U10195 ( .B1(n8511), .B2(P3_IR_REG_11__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8513) );
  INV_X1 U10196 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8512) );
  AOI22_X1 U10197 ( .A1(n8600), .A2(n15319), .B1(n8599), .B2(n15711), .ZN(
        n8514) );
  NAND2_X1 U10198 ( .A1(n13567), .A2(n16078), .ZN(n12706) );
  MUX2_X1 U10199 ( .A(n12706), .B(n7307), .S(n8720), .Z(n11949) );
  NAND2_X1 U10200 ( .A1(n11951), .A2(n11949), .ZN(n8516) );
  NAND2_X1 U10201 ( .A1(n15393), .A2(n11968), .ZN(n12709) );
  NAND2_X1 U10202 ( .A1(n15393), .A2(n16078), .ZN(n8830) );
  MUX2_X1 U10203 ( .A(n12709), .B(n8830), .S(n8720), .Z(n11948) );
  NAND2_X1 U10204 ( .A1(n8516), .A2(n11948), .ZN(n13499) );
  XNOR2_X1 U10205 ( .A(n8517), .B(n13566), .ZN(n13498) );
  NAND2_X1 U10206 ( .A1(n13499), .A2(n13498), .ZN(n8518) );
  XNOR2_X1 U10207 ( .A(n8521), .B(n8520), .ZN(n9272) );
  NAND2_X1 U10208 ( .A1(n9272), .A2(n12584), .ZN(n8526) );
  NOR2_X1 U10209 ( .A1(n8522), .A2(n8221), .ZN(n8523) );
  MUX2_X1 U10210 ( .A(n8221), .B(n8523), .S(P3_IR_REG_14__SCAN_IN), .Z(n8524)
         );
  OR2_X1 U10211 ( .A1(n8524), .A2(n8308), .ZN(n13634) );
  AOI22_X1 U10212 ( .A1(n8600), .A2(n15318), .B1(n8599), .B2(n13634), .ZN(
        n8525) );
  NAND2_X1 U10213 ( .A1(n8526), .A2(n8525), .ZN(n14014) );
  XNOR2_X1 U10214 ( .A(n14014), .B(n8720), .ZN(n8547) );
  NAND2_X1 U10215 ( .A1(n12573), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8532) );
  NAND2_X1 U10216 ( .A1(n8527), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8528) );
  AND2_X1 U10217 ( .A1(n8539), .A2(n8528), .ZN(n13883) );
  OR2_X1 U10218 ( .A1(n8590), .A2(n13883), .ZN(n8531) );
  INV_X1 U10219 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13884) );
  OR2_X1 U10220 ( .A1(n12577), .A2(n13884), .ZN(n8530) );
  INV_X1 U10221 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13951) );
  OR2_X1 U10222 ( .A1(n8556), .A2(n13951), .ZN(n8529) );
  NAND4_X1 U10223 ( .A1(n8532), .A2(n8531), .A3(n8530), .A4(n8529), .ZN(n13860) );
  XNOR2_X1 U10224 ( .A(n8547), .B(n13860), .ZN(n13536) );
  XNOR2_X1 U10225 ( .A(n8534), .B(n8533), .ZN(n16147) );
  NAND2_X1 U10226 ( .A1(n16147), .A2(n12584), .ZN(n8538) );
  OR2_X1 U10227 ( .A1(n8308), .A2(n8221), .ZN(n8536) );
  XNOR2_X1 U10228 ( .A(n8536), .B(n8535), .ZN(n16152) );
  AOI22_X1 U10229 ( .A1(n8600), .A2(n10437), .B1(n8599), .B2(n16152), .ZN(
        n8537) );
  NAND2_X1 U10230 ( .A1(n8538), .A2(n8537), .ZN(n13943) );
  XNOR2_X1 U10231 ( .A(n13943), .B(n8720), .ZN(n8548) );
  INV_X1 U10232 ( .A(n8548), .ZN(n8545) );
  NAND2_X1 U10233 ( .A1(n12573), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8544) );
  INV_X1 U10234 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n15778) );
  OR2_X1 U10235 ( .A1(n8889), .A2(n15778), .ZN(n8543) );
  NAND2_X1 U10236 ( .A1(n8539), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8540) );
  AND2_X1 U10237 ( .A1(n8557), .A2(n8540), .ZN(n13863) );
  OR2_X1 U10238 ( .A1(n8590), .A2(n13863), .ZN(n8542) );
  INV_X1 U10239 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n15767) );
  OR2_X1 U10240 ( .A1(n12577), .A2(n15767), .ZN(n8541) );
  NAND4_X1 U10241 ( .A1(n8544), .A2(n8543), .A3(n8542), .A4(n8541), .ZN(n13565) );
  NAND2_X1 U10242 ( .A1(n8545), .A2(n13565), .ZN(n8546) );
  AND2_X1 U10243 ( .A1(n13536), .A2(n8546), .ZN(n8551) );
  INV_X1 U10244 ( .A(n8546), .ZN(n8550) );
  INV_X1 U10245 ( .A(n13860), .ZN(n15391) );
  NAND2_X1 U10246 ( .A1(n8547), .A2(n15391), .ZN(n13538) );
  INV_X1 U10247 ( .A(n13565), .ZN(n13877) );
  XNOR2_X1 U10248 ( .A(n8548), .B(n13877), .ZN(n13540) );
  INV_X1 U10249 ( .A(n13540), .ZN(n8549) );
  AND2_X1 U10250 ( .A1(n13538), .A2(n8549), .ZN(n13542) );
  XNOR2_X1 U10251 ( .A(n8552), .B(P1_DATAO_REG_16__SCAN_IN), .ZN(n9873) );
  NAND2_X1 U10252 ( .A1(n9873), .A2(n12584), .ZN(n8555) );
  NAND2_X1 U10253 ( .A1(n8553), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8570) );
  INV_X1 U10254 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8569) );
  XNOR2_X1 U10255 ( .A(n8570), .B(n8569), .ZN(n13639) );
  INV_X1 U10256 ( .A(n13639), .ZN(n15795) );
  AOI22_X1 U10257 ( .A1(n8600), .A2(SI_16_), .B1(n8599), .B2(n15795), .ZN(
        n8554) );
  XNOR2_X1 U10258 ( .A(n13847), .B(n13084), .ZN(n13462) );
  NAND2_X1 U10259 ( .A1(n12573), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8562) );
  INV_X1 U10260 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13941) );
  OR2_X1 U10261 ( .A1(n8556), .A2(n13941), .ZN(n8561) );
  NAND2_X1 U10262 ( .A1(n8557), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8558) );
  AND2_X1 U10263 ( .A1(n8576), .A2(n8558), .ZN(n13848) );
  OR2_X1 U10264 ( .A1(n8590), .A2(n13848), .ZN(n8560) );
  INV_X1 U10265 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13849) );
  OR2_X1 U10266 ( .A1(n12577), .A2(n13849), .ZN(n8559) );
  NAND4_X1 U10267 ( .A1(n8562), .A2(n8561), .A3(n8560), .A4(n8559), .ZN(n13859) );
  INV_X1 U10268 ( .A(n13859), .ZN(n13823) );
  NAND2_X1 U10269 ( .A1(n13462), .A2(n13823), .ZN(n8563) );
  NAND2_X1 U10270 ( .A1(n13464), .A2(n8563), .ZN(n8566) );
  INV_X1 U10271 ( .A(n13462), .ZN(n8564) );
  NAND2_X1 U10272 ( .A1(n8564), .A2(n13859), .ZN(n8565) );
  XNOR2_X1 U10273 ( .A(n8568), .B(n8567), .ZN(n10039) );
  NAND2_X1 U10274 ( .A1(n10039), .A2(n12584), .ZN(n8575) );
  NAND2_X1 U10275 ( .A1(n8570), .A2(n8569), .ZN(n8571) );
  NAND2_X1 U10276 ( .A1(n8571), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8573) );
  XNOR2_X1 U10277 ( .A(n8573), .B(n8572), .ZN(n13641) );
  AOI22_X1 U10278 ( .A1(n8600), .A2(n15205), .B1(n8599), .B2(n13641), .ZN(
        n8574) );
  XNOR2_X1 U10279 ( .A(n14003), .B(n8720), .ZN(n13470) );
  NAND2_X1 U10280 ( .A1(n12573), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8581) );
  INV_X1 U10281 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n15804) );
  OR2_X1 U10282 ( .A1(n12577), .A2(n15804), .ZN(n8580) );
  NAND2_X1 U10283 ( .A1(n8576), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8577) );
  AND2_X1 U10284 ( .A1(n8588), .A2(n8577), .ZN(n13473) );
  OR2_X1 U10285 ( .A1(n8590), .A2(n13473), .ZN(n8579) );
  INV_X1 U10286 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n15819) );
  OR2_X1 U10287 ( .A1(n8889), .A2(n15819), .ZN(n8578) );
  NAND4_X1 U10288 ( .A1(n8581), .A2(n8580), .A3(n8579), .A4(n8578), .ZN(n13564) );
  NAND2_X1 U10289 ( .A1(n13470), .A2(n13843), .ZN(n8582) );
  XNOR2_X1 U10290 ( .A(n8584), .B(n8583), .ZN(n10323) );
  NAND2_X1 U10291 ( .A1(n10323), .A2(n12584), .ZN(n8587) );
  NAND2_X1 U10292 ( .A1(n7327), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8585) );
  XNOR2_X1 U10293 ( .A(n8585), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13647) );
  AOI22_X1 U10294 ( .A1(n8600), .A2(SI_18_), .B1(n8599), .B2(n13647), .ZN(
        n8586) );
  XNOR2_X1 U10295 ( .A(n13514), .B(n8720), .ZN(n8595) );
  NAND2_X1 U10296 ( .A1(n8898), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8594) );
  INV_X1 U10297 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13997) );
  OR2_X1 U10298 ( .A1(n8605), .A2(n13997), .ZN(n8593) );
  NAND2_X1 U10299 ( .A1(n8588), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8589) );
  AND2_X1 U10300 ( .A1(n8603), .A2(n8589), .ZN(n13814) );
  OR2_X1 U10301 ( .A1(n8590), .A2(n13814), .ZN(n8592) );
  INV_X1 U10302 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13815) );
  OR2_X1 U10303 ( .A1(n12577), .A2(n13815), .ZN(n8591) );
  XNOR2_X1 U10304 ( .A(n8595), .B(n13563), .ZN(n13515) );
  INV_X1 U10305 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11266) );
  AOI22_X1 U10306 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n11264), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n11266), .ZN(n8596) );
  INV_X1 U10307 ( .A(n8596), .ZN(n8597) );
  XNOR2_X1 U10308 ( .A(n8598), .B(n8597), .ZN(n10379) );
  NAND2_X1 U10309 ( .A1(n10379), .A2(n12584), .ZN(n8602) );
  AOI22_X1 U10310 ( .A1(n8600), .A2(SI_19_), .B1(n13670), .B2(n8599), .ZN(
        n8601) );
  NAND2_X1 U10311 ( .A1(n8602), .A2(n8601), .ZN(n13432) );
  XNOR2_X1 U10312 ( .A(n13432), .B(n8720), .ZN(n8610) );
  NAND2_X1 U10313 ( .A1(n8603), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8604) );
  NAND2_X1 U10314 ( .A1(n8615), .A2(n8604), .ZN(n13802) );
  NAND2_X1 U10315 ( .A1(n8887), .A2(n13802), .ZN(n8609) );
  INV_X1 U10316 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13993) );
  OR2_X1 U10317 ( .A1(n8605), .A2(n13993), .ZN(n8608) );
  INV_X1 U10318 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13930) );
  OR2_X1 U10319 ( .A1(n8889), .A2(n13930), .ZN(n8607) );
  INV_X1 U10320 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13653) );
  OR2_X1 U10321 ( .A1(n12577), .A2(n13653), .ZN(n8606) );
  XNOR2_X1 U10322 ( .A(n8610), .B(n13811), .ZN(n13433) );
  INV_X1 U10323 ( .A(n13811), .ZN(n13562) );
  NAND2_X1 U10324 ( .A1(n8610), .A2(n13562), .ZN(n13439) );
  XNOR2_X1 U10325 ( .A(n8612), .B(n8611), .ZN(n10606) );
  NAND2_X1 U10326 ( .A1(n10606), .A2(n12584), .ZN(n8614) );
  OR2_X1 U10327 ( .A1(n8884), .A2(n11223), .ZN(n8613) );
  XNOR2_X1 U10328 ( .A(n13788), .B(n13084), .ZN(n13490) );
  INV_X1 U10329 ( .A(n13490), .ZN(n8619) );
  NAND2_X1 U10330 ( .A1(n8615), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8616) );
  NAND2_X1 U10331 ( .A1(n8626), .A2(n8616), .ZN(n13789) );
  INV_X1 U10332 ( .A(n12577), .ZN(n8890) );
  AOI22_X1 U10333 ( .A1(n13789), .A2(n8887), .B1(n8890), .B2(
        P3_REG2_REG_20__SCAN_IN), .ZN(n8618) );
  AOI22_X1 U10334 ( .A1(n12573), .A2(P3_REG0_REG_20__SCAN_IN), .B1(n8898), 
        .B2(P3_REG1_REG_20__SCAN_IN), .ZN(n8617) );
  INV_X1 U10335 ( .A(n13799), .ZN(n13561) );
  NAND2_X1 U10336 ( .A1(n8619), .A2(n13561), .ZN(n13442) );
  NAND2_X1 U10337 ( .A1(n8621), .A2(n8620), .ZN(n8622) );
  NAND2_X1 U10338 ( .A1(n8623), .A2(n8622), .ZN(n10632) );
  INV_X1 U10339 ( .A(SI_21_), .ZN(n15183) );
  XNOR2_X1 U10340 ( .A(n13772), .B(n8720), .ZN(n8635) );
  NAND2_X1 U10341 ( .A1(n8626), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8627) );
  NAND2_X1 U10342 ( .A1(n8650), .A2(n8627), .ZN(n13773) );
  NAND2_X1 U10343 ( .A1(n13773), .A2(n8887), .ZN(n8630) );
  AOI22_X1 U10344 ( .A1(n12573), .A2(P3_REG0_REG_21__SCAN_IN), .B1(n8898), 
        .B2(P3_REG1_REG_21__SCAN_IN), .ZN(n8629) );
  NAND2_X1 U10345 ( .A1(n8890), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8628) );
  INV_X1 U10346 ( .A(n13783), .ZN(n13560) );
  NAND2_X1 U10347 ( .A1(n8635), .A2(n13560), .ZN(n8634) );
  AND2_X1 U10348 ( .A1(n13442), .A2(n8634), .ZN(n8631) );
  AND2_X1 U10349 ( .A1(n13439), .A2(n8631), .ZN(n8642) );
  NAND2_X1 U10350 ( .A1(n13440), .A2(n8642), .ZN(n8633) );
  INV_X1 U10351 ( .A(n8631), .ZN(n8632) );
  NAND2_X1 U10352 ( .A1(n13490), .A2(n13799), .ZN(n13441) );
  OR2_X1 U10353 ( .A1(n8632), .A2(n13441), .ZN(n8645) );
  INV_X1 U10354 ( .A(n8634), .ZN(n8636) );
  XNOR2_X1 U10355 ( .A(n8635), .B(n13783), .ZN(n13444) );
  OR2_X1 U10356 ( .A1(n8636), .A2(n13444), .ZN(n8644) );
  XNOR2_X1 U10357 ( .A(n8638), .B(n8637), .ZN(n10841) );
  NAND2_X1 U10358 ( .A1(n10841), .A2(n12584), .ZN(n8640) );
  OR2_X1 U10359 ( .A1(n8884), .A2(n15181), .ZN(n8639) );
  XNOR2_X1 U10360 ( .A(n13757), .B(n8720), .ZN(n8647) );
  INV_X1 U10361 ( .A(n8647), .ZN(n8641) );
  AND2_X1 U10362 ( .A1(n8642), .A2(n8641), .ZN(n8643) );
  NAND2_X1 U10363 ( .A1(n13440), .A2(n8643), .ZN(n8649) );
  AND2_X1 U10364 ( .A1(n8645), .A2(n8644), .ZN(n8646) );
  INV_X1 U10365 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n8654) );
  NAND2_X1 U10366 ( .A1(n8650), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U10367 ( .A1(n8663), .A2(n8651), .ZN(n13758) );
  NAND2_X1 U10368 ( .A1(n13758), .A2(n8887), .ZN(n8653) );
  AOI22_X1 U10369 ( .A1(n12573), .A2(P3_REG0_REG_22__SCAN_IN), .B1(n8898), 
        .B2(P3_REG1_REG_22__SCAN_IN), .ZN(n8652) );
  OAI211_X1 U10370 ( .C1(n12577), .C2(n8654), .A(n8653), .B(n8652), .ZN(n13735) );
  XNOR2_X1 U10371 ( .A(n8657), .B(n8656), .ZN(n11178) );
  NAND2_X1 U10372 ( .A1(n11178), .A2(n12584), .ZN(n8659) );
  INV_X1 U10373 ( .A(SI_23_), .ZN(n15287) );
  XOR2_X1 U10374 ( .A(n8720), .B(n13739), .Z(n8660) );
  NAND2_X1 U10375 ( .A1(n8661), .A2(n8660), .ZN(n13480) );
  NAND2_X1 U10376 ( .A1(n8663), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8664) );
  NAND2_X1 U10377 ( .A1(n8674), .A2(n8664), .ZN(n13744) );
  NAND2_X1 U10378 ( .A1(n13744), .A2(n8887), .ZN(n8670) );
  INV_X1 U10379 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n8667) );
  NAND2_X1 U10380 ( .A1(n8898), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8666) );
  NAND2_X1 U10381 ( .A1(n12573), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8665) );
  OAI211_X1 U10382 ( .C1(n8667), .C2(n12577), .A(n8666), .B(n8665), .ZN(n8668)
         );
  INV_X1 U10383 ( .A(n8668), .ZN(n8669) );
  XNOR2_X1 U10384 ( .A(n8671), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n11450) );
  NAND2_X1 U10385 ( .A1(n11450), .A2(n12584), .ZN(n8673) );
  INV_X1 U10386 ( .A(SI_24_), .ZN(n15201) );
  XNOR2_X1 U10387 ( .A(n13479), .B(n13084), .ZN(n8682) );
  NAND2_X1 U10388 ( .A1(n8674), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8675) );
  NAND2_X1 U10389 ( .A1(n8692), .A2(n8675), .ZN(n13729) );
  NAND2_X1 U10390 ( .A1(n13729), .A2(n8887), .ZN(n8681) );
  INV_X1 U10391 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n8678) );
  NAND2_X1 U10392 ( .A1(n8898), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8677) );
  NAND2_X1 U10393 ( .A1(n12573), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8676) );
  OAI211_X1 U10394 ( .C1(n8678), .C2(n12577), .A(n8677), .B(n8676), .ZN(n8679)
         );
  INV_X1 U10395 ( .A(n8679), .ZN(n8680) );
  NAND2_X1 U10396 ( .A1(n8682), .A2(n13738), .ZN(n13452) );
  INV_X1 U10397 ( .A(n8682), .ZN(n8683) );
  INV_X1 U10398 ( .A(n13738), .ZN(n13558) );
  NAND2_X1 U10399 ( .A1(n8683), .A2(n13558), .ZN(n8684) );
  OR2_X1 U10400 ( .A1(n8686), .A2(n8685), .ZN(n8687) );
  NAND2_X1 U10401 ( .A1(n8688), .A2(n8687), .ZN(n11589) );
  INV_X1 U10402 ( .A(SI_25_), .ZN(n11982) );
  XNOR2_X1 U10403 ( .A(n12632), .B(n13084), .ZN(n8700) );
  NAND2_X1 U10404 ( .A1(n8692), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8693) );
  NAND2_X1 U10405 ( .A1(n8705), .A2(n8693), .ZN(n13715) );
  NAND2_X1 U10406 ( .A1(n13715), .A2(n8887), .ZN(n8699) );
  INV_X1 U10407 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n8696) );
  NAND2_X1 U10408 ( .A1(n8898), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8695) );
  NAND2_X1 U10409 ( .A1(n12573), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8694) );
  OAI211_X1 U10410 ( .C1(n8696), .C2(n12577), .A(n8695), .B(n8694), .ZN(n8697)
         );
  INV_X1 U10411 ( .A(n8697), .ZN(n8698) );
  INV_X1 U10412 ( .A(n13725), .ZN(n13486) );
  NAND2_X1 U10413 ( .A1(n8700), .A2(n13486), .ZN(n8704) );
  INV_X1 U10414 ( .A(n8700), .ZN(n8701) );
  NAND2_X1 U10415 ( .A1(n8701), .A2(n13725), .ZN(n8702) );
  NAND2_X1 U10416 ( .A1(n8705), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8706) );
  NAND2_X1 U10417 ( .A1(n8707), .A2(n8706), .ZN(n13702) );
  NAND2_X1 U10418 ( .A1(n13702), .A2(n8887), .ZN(n8713) );
  INV_X1 U10419 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n8710) );
  NAND2_X1 U10420 ( .A1(n12573), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8709) );
  NAND2_X1 U10421 ( .A1(n8898), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8708) );
  OAI211_X1 U10422 ( .C1(n12577), .C2(n8710), .A(n8709), .B(n8708), .ZN(n8711)
         );
  INV_X1 U10423 ( .A(n8711), .ZN(n8712) );
  OR2_X1 U10424 ( .A1(n8715), .A2(n8714), .ZN(n8716) );
  NAND2_X1 U10425 ( .A1(n8717), .A2(n8716), .ZN(n11757) );
  INV_X1 U10426 ( .A(SI_26_), .ZN(n15301) );
  XNOR2_X1 U10427 ( .A(n13899), .B(n8720), .ZN(n8721) );
  NOR2_X1 U10428 ( .A1(n8721), .A2(n13557), .ZN(n8722) );
  AOI21_X1 U10429 ( .B1(n13557), .B2(n8721), .A(n8722), .ZN(n13526) );
  OAI21_X1 U10430 ( .B1(n8724), .B2(n8723), .A(n13097), .ZN(n8757) );
  INV_X1 U10431 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9117) );
  NAND2_X1 U10432 ( .A1(n9220), .A2(n9117), .ZN(n8726) );
  NAND2_X1 U10433 ( .A1(n11758), .A2(n11590), .ZN(n8725) );
  NOR2_X1 U10434 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .ZN(
        n8730) );
  NOR4_X1 U10435 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n8729) );
  NOR4_X1 U10436 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8728) );
  NOR4_X1 U10437 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8727) );
  NAND4_X1 U10438 ( .A1(n8730), .A2(n8729), .A3(n8728), .A4(n8727), .ZN(n8736)
         );
  NOR4_X1 U10439 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n8734) );
  NOR4_X1 U10440 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n8733) );
  NOR4_X1 U10441 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n8732) );
  NOR4_X1 U10442 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n8731) );
  NAND4_X1 U10443 ( .A1(n8734), .A2(n8733), .A3(n8732), .A4(n8731), .ZN(n8735)
         );
  OAI21_X1 U10444 ( .B1(n8736), .B2(n8735), .A(n9220), .ZN(n8912) );
  AND3_X1 U10445 ( .A1(n14017), .A2(n10312), .A3(n8912), .ZN(n8863) );
  NAND2_X1 U10446 ( .A1(n12623), .A2(n12596), .ZN(n8739) );
  NAND2_X1 U10447 ( .A1(n8737), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8738) );
  NAND2_X1 U10448 ( .A1(n8739), .A2(n8742), .ZN(n8917) );
  INV_X1 U10449 ( .A(n12596), .ZN(n12786) );
  OAI21_X1 U10450 ( .B1(n12786), .B2(n8742), .A(n13670), .ZN(n8740) );
  NAND2_X1 U10451 ( .A1(n8740), .A2(n12623), .ZN(n8741) );
  NAND2_X1 U10452 ( .A1(n8917), .A2(n8741), .ZN(n8865) );
  NAND3_X1 U10453 ( .A1(n8863), .A2(n8865), .A3(n16096), .ZN(n8746) );
  NAND2_X1 U10454 ( .A1(n8911), .A2(n8912), .ZN(n8743) );
  MUX2_X1 U10455 ( .A(n12792), .B(n12596), .S(n13656), .Z(n8744) );
  NAND2_X1 U10456 ( .A1(n8744), .A2(n12623), .ZN(n8916) );
  NOR2_X1 U10457 ( .A1(n8916), .A2(n12596), .ZN(n8864) );
  NAND2_X1 U10458 ( .A1(n8866), .A2(n8864), .ZN(n8745) );
  NAND2_X1 U10459 ( .A1(n8746), .A2(n8745), .ZN(n8756) );
  INV_X1 U10460 ( .A(n11590), .ZN(n8748) );
  INV_X1 U10461 ( .A(n11452), .ZN(n8747) );
  NAND2_X1 U10462 ( .A1(n8752), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8753) );
  MUX2_X1 U10463 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8753), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n8755) );
  NAND2_X1 U10464 ( .A1(n8755), .A2(n8754), .ZN(n8775) );
  NAND2_X1 U10465 ( .A1(n8757), .A2(n13527), .ZN(n8785) );
  NAND2_X1 U10466 ( .A1(n8863), .A2(n8758), .ZN(n8759) );
  NAND2_X1 U10467 ( .A1(n8760), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8761) );
  NAND2_X1 U10468 ( .A1(n12198), .A2(n8761), .ZN(n13686) );
  INV_X1 U10469 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n8764) );
  NAND2_X1 U10470 ( .A1(n12573), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8763) );
  NAND2_X1 U10471 ( .A1(n8898), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8762) );
  OAI211_X1 U10472 ( .C1(n8764), .C2(n12577), .A(n8763), .B(n8762), .ZN(n8765)
         );
  AND2_X1 U10473 ( .A1(n12596), .A2(n13656), .ZN(n8809) );
  INV_X1 U10474 ( .A(n8809), .ZN(n8766) );
  NOR2_X1 U10475 ( .A1(n8766), .A2(n12762), .ZN(n10086) );
  NAND2_X1 U10476 ( .A1(n9783), .A2(n10086), .ZN(n8776) );
  INV_X1 U10477 ( .A(n8776), .ZN(n12789) );
  NAND2_X1 U10478 ( .A1(n8866), .A2(n12789), .ZN(n8769) );
  INV_X1 U10479 ( .A(n8769), .ZN(n8768) );
  INV_X1 U10480 ( .A(n12193), .ZN(n12788) );
  NAND2_X1 U10481 ( .A1(n12788), .A2(n9817), .ZN(n9810) );
  NAND2_X1 U10482 ( .A1(n9782), .A2(n9810), .ZN(n8855) );
  AND2_X1 U10483 ( .A1(n8768), .A2(n8855), .ZN(n13546) );
  INV_X1 U10484 ( .A(n8865), .ZN(n8773) );
  INV_X1 U10485 ( .A(n8864), .ZN(n8770) );
  OR2_X1 U10486 ( .A1(n8866), .A2(n8770), .ZN(n8772) );
  OR2_X1 U10487 ( .A1(n12762), .A2(n8809), .ZN(n8915) );
  AND2_X1 U10488 ( .A1(n8915), .A2(n8981), .ZN(n8771) );
  OAI211_X1 U10489 ( .C1(n8863), .C2(n8773), .A(n8772), .B(n8771), .ZN(n8774)
         );
  NAND2_X1 U10490 ( .A1(n8774), .A2(P3_STATE_REG_SCAN_IN), .ZN(n8779) );
  INV_X1 U10491 ( .A(n8775), .ZN(n9780) );
  NAND2_X1 U10492 ( .A1(n9780), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12791) );
  OAI21_X1 U10493 ( .B1(n8866), .B2(n8776), .A(n12791), .ZN(n8777) );
  INV_X1 U10494 ( .A(n8777), .ZN(n8778) );
  AOI22_X1 U10495 ( .A1(n13692), .A2(n13550), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n8780) );
  OAI21_X1 U10496 ( .B1(n13712), .B2(n13548), .A(n8780), .ZN(n8781) );
  AOI21_X1 U10497 ( .B1(n7408), .B2(n13546), .A(n8781), .ZN(n8782) );
  INV_X1 U10498 ( .A(n8783), .ZN(n8784) );
  NAND2_X1 U10499 ( .A1(n8785), .A2(n8784), .ZN(P3_U3154) );
  INV_X1 U10500 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n8870) );
  NAND2_X1 U10501 ( .A1(n8786), .A2(n13678), .ZN(n13682) );
  INV_X1 U10502 ( .A(n9769), .ZN(n10087) );
  NAND2_X1 U10503 ( .A1(n9769), .A2(n10524), .ZN(n12646) );
  INV_X1 U10504 ( .A(n13578), .ZN(n10422) );
  NAND2_X1 U10505 ( .A1(n10422), .A2(n10319), .ZN(n10420) );
  NAND2_X1 U10506 ( .A1(n10636), .A2(n8788), .ZN(n12650) );
  INV_X1 U10507 ( .A(n8788), .ZN(n15872) );
  NAND2_X1 U10508 ( .A1(n13576), .A2(n15872), .ZN(n12649) );
  INV_X1 U10509 ( .A(n10639), .ZN(n15912) );
  NAND2_X1 U10510 ( .A1(n10988), .A2(n10639), .ZN(n12656) );
  NAND2_X1 U10511 ( .A1(n12657), .A2(n12656), .ZN(n10879) );
  NAND2_X1 U10512 ( .A1(n10876), .A2(n12600), .ZN(n8789) );
  NAND2_X1 U10513 ( .A1(n8789), .A2(n12656), .ZN(n11021) );
  NAND2_X1 U10514 ( .A1(n11113), .A2(n11030), .ZN(n12661) );
  INV_X1 U10515 ( .A(n11113), .ZN(n13575) );
  NAND2_X1 U10516 ( .A1(n13575), .A2(n11061), .ZN(n12662) );
  NAND2_X1 U10517 ( .A1(n12661), .A2(n12662), .ZN(n11023) );
  NAND2_X1 U10518 ( .A1(n11021), .A2(n12659), .ZN(n8790) );
  NAND2_X1 U10519 ( .A1(n8790), .A2(n12661), .ZN(n11076) );
  XNOR2_X1 U10520 ( .A(n13574), .B(n11116), .ZN(n11075) );
  NAND2_X1 U10521 ( .A1(n11076), .A2(n11075), .ZN(n8791) );
  NAND2_X1 U10522 ( .A1(n11208), .A2(n11116), .ZN(n12666) );
  NAND2_X1 U10523 ( .A1(n8791), .A2(n12666), .ZN(n11282) );
  NAND2_X1 U10524 ( .A1(n11596), .A2(n11211), .ZN(n12670) );
  INV_X1 U10525 ( .A(n11596), .ZN(n13573) );
  INV_X1 U10526 ( .A(n11211), .ZN(n15983) );
  NAND2_X1 U10527 ( .A1(n13573), .A2(n15983), .ZN(n12671) );
  NAND2_X1 U10528 ( .A1(n11282), .A2(n12668), .ZN(n8792) );
  NAND2_X1 U10529 ( .A1(n8792), .A2(n12670), .ZN(n11592) );
  NAND2_X1 U10530 ( .A1(n11469), .A2(n11397), .ZN(n12677) );
  INV_X1 U10531 ( .A(n11397), .ZN(n15999) );
  NAND2_X1 U10532 ( .A1(n13572), .A2(n15999), .ZN(n12678) );
  NAND2_X1 U10533 ( .A1(n12677), .A2(n12678), .ZN(n11591) );
  INV_X1 U10534 ( .A(n11591), .ZN(n12675) );
  NAND2_X1 U10535 ( .A1(n11592), .A2(n12675), .ZN(n8793) );
  NAND2_X1 U10536 ( .A1(n12687), .A2(n16005), .ZN(n8821) );
  INV_X1 U10537 ( .A(n12687), .ZN(n13571) );
  NAND2_X1 U10538 ( .A1(n13571), .A2(n12682), .ZN(n8794) );
  INV_X1 U10539 ( .A(n12603), .ZN(n12680) );
  NOR2_X1 U10540 ( .A1(n13570), .A2(n16026), .ZN(n11579) );
  INV_X1 U10541 ( .A(n11579), .ZN(n8795) );
  NAND2_X1 U10542 ( .A1(n8796), .A2(n8795), .ZN(n8797) );
  NAND2_X1 U10543 ( .A1(n13570), .A2(n16026), .ZN(n11578) );
  NAND2_X1 U10544 ( .A1(n11859), .A2(n13953), .ZN(n12694) );
  INV_X1 U10545 ( .A(n11859), .ZN(n13569) );
  INV_X1 U10546 ( .A(n13953), .ZN(n11701) );
  NAND2_X1 U10547 ( .A1(n13569), .A2(n11701), .ZN(n12695) );
  INV_X1 U10548 ( .A(n12691), .ZN(n8824) );
  INV_X1 U10549 ( .A(n11947), .ZN(n8828) );
  NAND2_X1 U10550 ( .A1(n11961), .A2(n8828), .ZN(n12700) );
  NAND2_X1 U10551 ( .A1(n13568), .A2(n11947), .ZN(n12707) );
  NAND2_X1 U10552 ( .A1(n11860), .A2(n12700), .ZN(n11957) );
  NAND2_X1 U10553 ( .A1(n16095), .A2(n13566), .ZN(n12704) );
  OR2_X1 U10554 ( .A1(n14014), .A2(n13860), .ZN(n8831) );
  OR2_X1 U10555 ( .A1(n16095), .A2(n13566), .ZN(n13878) );
  AND2_X1 U10556 ( .A1(n8831), .A2(n13878), .ZN(n12713) );
  NAND2_X1 U10557 ( .A1(n14014), .A2(n13860), .ZN(n12714) );
  OR2_X1 U10558 ( .A1(n13943), .A2(n13565), .ZN(n12718) );
  NAND2_X1 U10559 ( .A1(n13943), .A2(n13565), .ZN(n12719) );
  NAND2_X1 U10560 ( .A1(n12718), .A2(n12719), .ZN(n13837) );
  OR2_X1 U10561 ( .A1(n13847), .A2(n13859), .ZN(n12722) );
  NAND2_X1 U10562 ( .A1(n13847), .A2(n13859), .ZN(n12726) );
  NAND2_X1 U10563 ( .A1(n13846), .A2(n13845), .ZN(n13844) );
  NAND2_X1 U10564 ( .A1(n13847), .A2(n13823), .ZN(n8798) );
  NAND2_X1 U10565 ( .A1(n14003), .A2(n13564), .ZN(n12735) );
  NAND2_X1 U10566 ( .A1(n12730), .A2(n12735), .ZN(n13820) );
  INV_X1 U10567 ( .A(n13820), .ZN(n13826) );
  NAND2_X1 U10568 ( .A1(n13514), .A2(n13824), .ZN(n12731) );
  NAND2_X1 U10569 ( .A1(n8799), .A2(n12738), .ZN(n13763) );
  NAND2_X1 U10570 ( .A1(n13432), .A2(n13811), .ZN(n12745) );
  NAND2_X1 U10571 ( .A1(n13778), .A2(n12745), .ZN(n13800) );
  INV_X1 U10572 ( .A(n12748), .ZN(n8800) );
  NAND2_X1 U10573 ( .A1(n13788), .A2(n13799), .ZN(n12749) );
  NAND2_X1 U10574 ( .A1(n12748), .A2(n12749), .ZN(n12615) );
  OR2_X1 U10575 ( .A1(n8800), .A2(n13781), .ZN(n8802) );
  AND2_X1 U10576 ( .A1(n13796), .A2(n8802), .ZN(n13764) );
  NAND2_X1 U10577 ( .A1(n13772), .A2(n13783), .ZN(n12754) );
  AND2_X1 U10578 ( .A1(n13764), .A2(n13769), .ZN(n8801) );
  INV_X1 U10579 ( .A(n13769), .ZN(n8805) );
  INV_X1 U10580 ( .A(n8802), .ZN(n8804) );
  AND2_X1 U10581 ( .A1(n13778), .A2(n12748), .ZN(n8803) );
  OR2_X1 U10582 ( .A1(n13757), .A2(n13771), .ZN(n12757) );
  NAND2_X1 U10583 ( .A1(n13757), .A2(n13771), .ZN(n12758) );
  NAND2_X1 U10584 ( .A1(n12757), .A2(n12758), .ZN(n12752) );
  NAND2_X1 U10585 ( .A1(n13739), .A2(n13752), .ZN(n12764) );
  OR2_X1 U10586 ( .A1(n13479), .A2(n13738), .ZN(n12631) );
  XNOR2_X1 U10587 ( .A(n12632), .B(n13725), .ZN(n13710) );
  NAND2_X1 U10588 ( .A1(n13899), .A2(n13712), .ZN(n12634) );
  INV_X1 U10589 ( .A(n12599), .ZN(n8807) );
  AND2_X1 U10590 ( .A1(n16096), .A2(n8809), .ZN(n8810) );
  NAND2_X1 U10591 ( .A1(n8865), .A2(n8810), .ZN(n8812) );
  NAND3_X1 U10592 ( .A1(n12786), .A2(n12792), .A3(n13656), .ZN(n8811) );
  NAND2_X1 U10593 ( .A1(n12604), .A2(n10421), .ZN(n15880) );
  NAND2_X1 U10594 ( .A1(n9769), .A2(n8787), .ZN(n15878) );
  NAND2_X1 U10595 ( .A1(n15880), .A2(n15878), .ZN(n8813) );
  NAND2_X1 U10596 ( .A1(n10636), .A2(n15872), .ZN(n10877) );
  AND2_X1 U10597 ( .A1(n10879), .A2(n10877), .ZN(n8814) );
  NAND2_X1 U10598 ( .A1(n15877), .A2(n8814), .ZN(n10878) );
  NAND2_X1 U10599 ( .A1(n15874), .A2(n10639), .ZN(n8815) );
  NAND2_X1 U10600 ( .A1(n10878), .A2(n8815), .ZN(n11022) );
  NAND2_X1 U10601 ( .A1(n11022), .A2(n11023), .ZN(n8817) );
  NAND2_X1 U10602 ( .A1(n13575), .A2(n11030), .ZN(n8816) );
  INV_X1 U10603 ( .A(n11116), .ZN(n12665) );
  NAND2_X1 U10604 ( .A1(n11208), .A2(n12665), .ZN(n8818) );
  NAND2_X1 U10605 ( .A1(n13573), .A2(n11211), .ZN(n8819) );
  NAND2_X1 U10606 ( .A1(n11285), .A2(n8819), .ZN(n11594) );
  AND2_X1 U10607 ( .A1(n13572), .A2(n11397), .ZN(n8820) );
  NAND2_X1 U10608 ( .A1(n11402), .A2(n12603), .ZN(n11401) );
  NAND2_X1 U10609 ( .A1(n11401), .A2(n8821), .ZN(n11581) );
  NAND2_X1 U10610 ( .A1(n13570), .A2(n8822), .ZN(n8823) );
  NAND2_X1 U10611 ( .A1(n11581), .A2(n8823), .ZN(n11691) );
  NAND2_X1 U10612 ( .A1(n11693), .A2(n16026), .ZN(n11690) );
  AND2_X1 U10613 ( .A1(n8824), .A2(n11690), .ZN(n8825) );
  NAND2_X1 U10614 ( .A1(n13569), .A2(n13953), .ZN(n8826) );
  NAND2_X1 U10615 ( .A1(n11961), .A2(n11947), .ZN(n8827) );
  INV_X1 U10616 ( .A(n11960), .ZN(n8829) );
  AND2_X1 U10617 ( .A1(n16095), .A2(n13876), .ZN(n13869) );
  OR2_X1 U10618 ( .A1(n14014), .A2(n15391), .ZN(n8834) );
  INV_X1 U10619 ( .A(n8834), .ZN(n8832) );
  NAND2_X1 U10620 ( .A1(n8831), .A2(n12714), .ZN(n13872) );
  NOR2_X1 U10621 ( .A1(n8832), .A2(n13872), .ZN(n8836) );
  OR2_X1 U10622 ( .A1(n13869), .A2(n8836), .ZN(n13834) );
  OR2_X1 U10623 ( .A1(n13834), .A2(n8181), .ZN(n8833) );
  OR2_X1 U10624 ( .A1(n16095), .A2(n13876), .ZN(n13870) );
  AND2_X1 U10625 ( .A1(n13870), .A2(n8834), .ZN(n8835) );
  OR2_X1 U10626 ( .A1(n8836), .A2(n8835), .ZN(n13835) );
  OR2_X1 U10627 ( .A1(n13943), .A2(n13877), .ZN(n13838) );
  OR2_X1 U10628 ( .A1(n13845), .A2(n13838), .ZN(n8837) );
  NAND2_X1 U10629 ( .A1(n8837), .A2(n12726), .ZN(n8838) );
  NAND2_X1 U10630 ( .A1(n13821), .A2(n13820), .ZN(n8841) );
  OR2_X1 U10631 ( .A1(n14003), .A2(n13843), .ZN(n8840) );
  OR2_X1 U10632 ( .A1(n13514), .A2(n13563), .ZN(n13795) );
  NAND2_X1 U10633 ( .A1(n13432), .A2(n13562), .ZN(n8843) );
  NAND2_X1 U10634 ( .A1(n13788), .A2(n13561), .ZN(n8845) );
  NAND2_X1 U10635 ( .A1(n13757), .A2(n13735), .ZN(n8846) );
  NAND2_X1 U10636 ( .A1(n13749), .A2(n8846), .ZN(n8848) );
  OR2_X1 U10637 ( .A1(n13757), .A2(n13735), .ZN(n8847) );
  NAND2_X1 U10638 ( .A1(n8848), .A2(n8847), .ZN(n8849) );
  NAND2_X1 U10639 ( .A1(n13739), .A2(n13559), .ZN(n8850) );
  AOI21_X2 U10640 ( .B1(n13558), .B2(n13479), .A(n13727), .ZN(n13711) );
  NOR2_X1 U10641 ( .A1(n13899), .A2(n13557), .ZN(n8851) );
  INV_X1 U10642 ( .A(n13899), .ZN(n13704) );
  AOI21_X1 U10643 ( .B1(n12599), .B2(n8852), .A(n8895), .ZN(n8859) );
  NAND2_X1 U10644 ( .A1(n12641), .A2(n12786), .ZN(n8854) );
  NAND2_X1 U10645 ( .A1(n13670), .A2(n12792), .ZN(n8853) );
  INV_X1 U10646 ( .A(n8855), .ZN(n8856) );
  OAI22_X1 U10647 ( .A1(n8896), .A2(n15390), .B1(n13712), .B2(n15392), .ZN(
        n8857) );
  AOI21_X1 U10648 ( .B1(n16082), .B2(n13695), .A(n13691), .ZN(n13895) );
  OAI21_X1 U10649 ( .B1(n10086), .B2(n8864), .A(n8863), .ZN(n8868) );
  NAND2_X1 U10650 ( .A1(n8866), .A2(n8865), .ZN(n8867) );
  NAND2_X1 U10651 ( .A1(n8868), .A2(n8867), .ZN(n8869) );
  MUX2_X1 U10652 ( .A(n8870), .B(n13895), .S(n16104), .Z(n8871) );
  NAND2_X1 U10653 ( .A1(n8871), .A2(n8169), .ZN(P3_U3454) );
  INV_X1 U10654 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8908) );
  INV_X1 U10655 ( .A(n13682), .ZN(n8880) );
  INV_X1 U10656 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n15153) );
  NAND2_X1 U10657 ( .A1(n15153), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8882) );
  INV_X1 U10658 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n12125) );
  NAND2_X1 U10659 ( .A1(n12125), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8874) );
  AND2_X1 U10660 ( .A1(n8882), .A2(n8874), .ZN(n8875) );
  OR2_X1 U10661 ( .A1(n8876), .A2(n8875), .ZN(n8877) );
  NAND2_X1 U10662 ( .A1(n8883), .A2(n8877), .ZN(n12194) );
  INV_X1 U10663 ( .A(SI_28_), .ZN(n15293) );
  NAND2_X1 U10664 ( .A1(n13094), .A2(n8896), .ZN(n12777) );
  INV_X1 U10665 ( .A(n8881), .ZN(n12776) );
  INV_X1 U10666 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14587) );
  XNOR2_X1 U10667 ( .A(n14587), .B(P2_DATAO_REG_29__SCAN_IN), .ZN(n12562) );
  XNOR2_X1 U10668 ( .A(n12564), .B(n12562), .ZN(n12195) );
  NAND2_X1 U10669 ( .A1(n12195), .A2(n12584), .ZN(n8886) );
  INV_X1 U10670 ( .A(SI_29_), .ZN(n15289) );
  OR2_X1 U10671 ( .A1(n8884), .A2(n15289), .ZN(n8885) );
  INV_X1 U10672 ( .A(n12198), .ZN(n8888) );
  NAND2_X1 U10673 ( .A1(n8888), .A2(n8887), .ZN(n12581) );
  INV_X1 U10674 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8923) );
  NAND2_X1 U10675 ( .A1(n12573), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8892) );
  NAND2_X1 U10676 ( .A1(n8890), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8891) );
  OAI211_X1 U10677 ( .C1(n8923), .C2(n8889), .A(n8892), .B(n8891), .ZN(n8893)
         );
  INV_X1 U10678 ( .A(n8893), .ZN(n8894) );
  NAND2_X1 U10679 ( .A1(n8909), .A2(n13681), .ZN(n12591) );
  NAND2_X1 U10680 ( .A1(n12774), .A2(n12591), .ZN(n12618) );
  XNOR2_X1 U10681 ( .A(n12587), .B(n12618), .ZN(n12203) );
  NOR2_X1 U10682 ( .A1(n12203), .A2(n13944), .ZN(n8907) );
  XNOR2_X1 U10683 ( .A(n8897), .B(n12618), .ZN(n8906) );
  INV_X1 U10684 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n8901) );
  NAND2_X1 U10685 ( .A1(n8898), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8900) );
  NAND2_X1 U10686 ( .A1(n12573), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8899) );
  OAI211_X1 U10687 ( .C1(n8901), .C2(n12577), .A(n8900), .B(n8899), .ZN(n8902)
         );
  INV_X1 U10688 ( .A(n8902), .ZN(n8903) );
  NAND2_X1 U10689 ( .A1(n12581), .A2(n8903), .ZN(n13556) );
  NAND2_X1 U10690 ( .A1(n12788), .A2(P3_B_REG_SCAN_IN), .ZN(n8904) );
  AOI22_X1 U10691 ( .A1(n15876), .A2(n7408), .B1(n13556), .B2(n13959), .ZN(
        n8905) );
  NOR2_X1 U10692 ( .A1(n8907), .A2(n12197), .ZN(n8922) );
  MUX2_X1 U10693 ( .A(n8908), .B(n8922), .S(n16104), .Z(n8910) );
  NAND2_X1 U10694 ( .A1(n8910), .A2(n8168), .ZN(P3_U3456) );
  XNOR2_X1 U10695 ( .A(n10312), .B(n8911), .ZN(n8914) );
  AND2_X1 U10696 ( .A1(n8912), .A2(n9783), .ZN(n8913) );
  AND2_X1 U10697 ( .A1(n8914), .A2(n8913), .ZN(n10316) );
  AND2_X1 U10698 ( .A1(n8916), .A2(n12792), .ZN(n10310) );
  NAND2_X1 U10699 ( .A1(n10310), .A2(n8915), .ZN(n10309) );
  NAND2_X1 U10700 ( .A1(n10312), .A2(n10309), .ZN(n8920) );
  INV_X1 U10701 ( .A(n10312), .ZN(n8918) );
  NAND3_X1 U10702 ( .A1(n8918), .A2(n8917), .A3(n8916), .ZN(n8919) );
  AND2_X1 U10703 ( .A1(n8920), .A2(n8919), .ZN(n8921) );
  MUX2_X1 U10704 ( .A(n8923), .B(n8922), .S(n16101), .Z(n8924) );
  NAND2_X1 U10705 ( .A1(n8924), .A2(n8167), .ZN(P3_U3488) );
  INV_X2 U10706 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9563) );
  NAND2_X1 U10707 ( .A1(n8933), .A2(n8928), .ZN(n8929) );
  NAND2_X1 U10708 ( .A1(n8934), .A2(n9477), .ZN(n8930) );
  XNOR2_X1 U10709 ( .A(n8933), .B(P2_IR_REG_24__SCAN_IN), .ZN(n9547) );
  NAND2_X1 U10710 ( .A1(n8935), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8936) );
  INV_X1 U10711 ( .A(n9544), .ZN(n11753) );
  NOR2_X2 U10712 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9054) );
  AND2_X2 U10713 ( .A1(n9054), .A2(n8937), .ZN(n9036) );
  NOR2_X1 U10714 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n8941) );
  NOR2_X2 U10715 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n8953) );
  INV_X1 U10716 ( .A(n8953), .ZN(n8947) );
  INV_X1 U10717 ( .A(n9084), .ZN(n8949) );
  NAND2_X1 U10718 ( .A1(n8970), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8951) );
  NOR2_X1 U10719 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n8952) );
  INV_X1 U10720 ( .A(n8962), .ZN(n8954) );
  NAND2_X1 U10721 ( .A1(n8959), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8960) );
  MUX2_X1 U10722 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8960), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n8963) );
  NOR3_X1 U10723 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .A3(P1_IR_REG_25__SCAN_IN), .ZN(n8961) );
  NAND2_X1 U10724 ( .A1(n8962), .A2(n8961), .ZN(n9074) );
  NAND2_X1 U10725 ( .A1(n9067), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8964) );
  MUX2_X1 U10726 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8964), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n8967) );
  INV_X1 U10727 ( .A(n9067), .ZN(n8965) );
  NAND2_X1 U10728 ( .A1(n8965), .A2(n9072), .ZN(n8966) );
  NOR2_X1 U10729 ( .A1(n15161), .A2(n15159), .ZN(n8968) );
  NAND2_X1 U10730 ( .A1(n9084), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8969) );
  MUX2_X1 U10731 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8969), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n8971) );
  NAND2_X1 U10732 ( .A1(n8971), .A2(n8970), .ZN(n10076) );
  NAND2_X1 U10733 ( .A1(n10076), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9063) );
  OR2_X2 U10734 ( .A1(n10077), .A2(n9063), .ZN(n14752) );
  XNOR2_X1 U10735 ( .A(n8973), .B(n8972), .ZN(n8974) );
  NOR2_X1 U10736 ( .A1(n8974), .A2(n13539), .ZN(n8980) );
  NOR2_X1 U10737 ( .A1(n13554), .A2(n11947), .ZN(n8979) );
  INV_X1 U10738 ( .A(n11862), .ZN(n8975) );
  AND2_X1 U10739 ( .A1(n13550), .A2(n8975), .ZN(n8978) );
  INV_X1 U10740 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n15373) );
  OR2_X1 U10741 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15373), .ZN(n15698) );
  NAND2_X1 U10742 ( .A1(n13546), .A2(n13567), .ZN(n8976) );
  OAI211_X1 U10743 ( .C1(n11859), .C2(n13548), .A(n15698), .B(n8976), .ZN(
        n8977) );
  NOR2_X1 U10744 ( .A1(n9540), .A2(P3_STATE_REG_SCAN_IN), .ZN(n16149) );
  INV_X1 U10745 ( .A(n16149), .ZN(n13082) );
  OAI222_X1 U10746 ( .A1(P3_U3151), .A2(n10772), .B1(n13082), .B2(n8983), .C1(
        n8982), .C2(n13083), .ZN(P3_U3289) );
  OAI222_X1 U10747 ( .A1(n9932), .A2(P3_U3151), .B1(n13082), .B2(n8984), .C1(
        n8991), .C2(n13083), .ZN(P3_U3294) );
  OAI222_X1 U10748 ( .A1(P3_U3151), .A2(n11328), .B1(n13083), .B2(n8986), .C1(
        n13082), .C2(n8985), .ZN(P3_U3287) );
  NOR2_X1 U10749 ( .A1(n9540), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14591) );
  INV_X2 U10750 ( .A(n14591), .ZN(n14588) );
  NAND2_X1 U10751 ( .A1(n8987), .A2(n9296), .ZN(n8988) );
  XNOR2_X1 U10752 ( .A(n8992), .B(SI_1_), .ZN(n9001) );
  MUX2_X1 U10753 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n8990), .Z(n9002) );
  NAND2_X1 U10754 ( .A1(n9001), .A2(n9002), .ZN(n8994) );
  OR2_X1 U10755 ( .A1(n8992), .A2(n8991), .ZN(n8993) );
  NAND2_X1 U10756 ( .A1(n8994), .A2(n8993), .ZN(n9010) );
  XNOR2_X1 U10757 ( .A(n9010), .B(SI_2_), .ZN(n9007) );
  MUX2_X1 U10758 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n7178), .Z(n9008) );
  XNOR2_X1 U10759 ( .A(n8995), .B(n9008), .ZN(n9541) );
  INV_X1 U10760 ( .A(n9541), .ZN(n9057) );
  NOR2_X1 U10761 ( .A1(n8996), .A2(n14582), .ZN(n8997) );
  MUX2_X1 U10762 ( .A(n14582), .B(n8997), .S(P2_IR_REG_2__SCAN_IN), .Z(n8998)
         );
  NOR2_X1 U10763 ( .A1(n8998), .A2(n9014), .ZN(n14204) );
  INV_X1 U10764 ( .A(n14204), .ZN(n8999) );
  OAI222_X1 U10765 ( .A1(n14588), .A2(n9000), .B1(n14593), .B2(n9057), .C1(
        P2_U3088), .C2(n8999), .ZN(P2_U3325) );
  XNOR2_X1 U10766 ( .A(n9002), .B(n9001), .ZN(n9615) );
  NAND2_X1 U10767 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9003) );
  MUX2_X1 U10768 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9003), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n9005) );
  INV_X1 U10769 ( .A(n8996), .ZN(n9004) );
  NAND2_X1 U10770 ( .A1(n9005), .A2(n9004), .ZN(n9706) );
  OAI222_X1 U10771 ( .A1(n14588), .A2(n9006), .B1(n14593), .B2(n9615), .C1(
        n9706), .C2(P2_U3088), .ZN(P2_U3326) );
  INV_X1 U10772 ( .A(n9007), .ZN(n9009) );
  NAND2_X1 U10773 ( .A1(n9009), .A2(n9008), .ZN(n9012) );
  NAND2_X1 U10774 ( .A1(n9010), .A2(SI_2_), .ZN(n9011) );
  NAND2_X1 U10775 ( .A1(n9012), .A2(n9011), .ZN(n9032) );
  INV_X1 U10776 ( .A(n9877), .ZN(n10040) );
  NAND2_X1 U10777 ( .A1(n9016), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9015) );
  MUX2_X1 U10778 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9015), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n9017) );
  AND2_X1 U10779 ( .A1(n9017), .A2(n9059), .ZN(n9878) );
  INV_X1 U10780 ( .A(n9878), .ZN(n15410) );
  OAI222_X1 U10781 ( .A1(n14588), .A2(n9018), .B1(n14593), .B2(n10040), .C1(
        P2_U3088), .C2(n15410), .ZN(P2_U3324) );
  INV_X1 U10782 ( .A(n13083), .ZN(n16148) );
  AOI222_X1 U10783 ( .A1(n9019), .A2(n16149), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9834), .C1(SI_3_), .C2(n16148), .ZN(n9020) );
  INV_X1 U10784 ( .A(n9020), .ZN(P3_U3292) );
  AOI222_X1 U10785 ( .A1(n9021), .A2(n16149), .B1(SI_5_), .B2(n16148), .C1(
        n10174), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9022) );
  INV_X1 U10786 ( .A(n9022), .ZN(P3_U3290) );
  AOI222_X1 U10787 ( .A1(n9023), .A2(n16149), .B1(n10151), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_4_), .C2(n16148), .ZN(n9024) );
  INV_X1 U10788 ( .A(n9024), .ZN(P3_U3291) );
  AOI222_X1 U10789 ( .A1(n9025), .A2(n16149), .B1(n15672), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_7_), .C2(n16148), .ZN(n9026) );
  INV_X1 U10790 ( .A(n9026), .ZN(P3_U3288) );
  AOI222_X1 U10791 ( .A1(n9027), .A2(n16149), .B1(SI_9_), .B2(n16148), .C1(
        n15685), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9028) );
  INV_X1 U10792 ( .A(n9028), .ZN(P3_U3286) );
  INV_X1 U10793 ( .A(n9029), .ZN(n9030) );
  INV_X1 U10794 ( .A(SI_2_), .ZN(n15328) );
  OAI222_X1 U10795 ( .A1(n9956), .A2(P3_U3151), .B1(n13082), .B2(n9030), .C1(
        n15328), .C2(n13083), .ZN(P3_U3293) );
  NAND2_X1 U10796 ( .A1(n9032), .A2(n9031), .ZN(n9035) );
  NAND2_X1 U10797 ( .A1(n9033), .A2(SI_3_), .ZN(n9034) );
  NAND2_X1 U10798 ( .A1(n9035), .A2(n9034), .ZN(n9046) );
  MUX2_X1 U10799 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n7178), .Z(n9047) );
  XNOR2_X1 U10800 ( .A(n9047), .B(SI_4_), .ZN(n9044) );
  XNOR2_X1 U10801 ( .A(n9046), .B(n9044), .ZN(n10052) );
  INV_X1 U10802 ( .A(n10052), .ZN(n9040) );
  INV_X1 U10803 ( .A(n9036), .ZN(n9089) );
  NAND2_X1 U10804 ( .A1(n9091), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9037) );
  XNOR2_X1 U10805 ( .A(n9037), .B(P1_IR_REG_4__SCAN_IN), .ZN(n14808) );
  INV_X1 U10806 ( .A(n14808), .ZN(n14800) );
  OAI222_X1 U10807 ( .A1(n15157), .A2(n9038), .B1(n15167), .B2(n9040), .C1(
        P1_U3086), .C2(n14800), .ZN(P1_U3351) );
  INV_X1 U10808 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9041) );
  NAND2_X1 U10809 ( .A1(n9059), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9039) );
  XNOR2_X1 U10810 ( .A(n9039), .B(P2_IR_REG_4__SCAN_IN), .ZN(n9884) );
  INV_X1 U10811 ( .A(n9884), .ZN(n9694) );
  OAI222_X1 U10812 ( .A1(n14588), .A2(n9041), .B1(n14593), .B2(n9040), .C1(
        P2_U3088), .C2(n9694), .ZN(P2_U3323) );
  AOI222_X1 U10813 ( .A1(n9042), .A2(n16149), .B1(SI_10_), .B2(n16148), .C1(
        n13580), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9043) );
  INV_X1 U10814 ( .A(n9043), .ZN(P3_U3285) );
  INV_X1 U10815 ( .A(n9044), .ZN(n9045) );
  NAND2_X1 U10816 ( .A1(n9046), .A2(n9045), .ZN(n9049) );
  NAND2_X1 U10817 ( .A1(n9047), .A2(SI_4_), .ZN(n9048) );
  MUX2_X1 U10818 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n7178), .Z(n9105) );
  XNOR2_X1 U10819 ( .A(n9105), .B(SI_5_), .ZN(n9102) );
  XNOR2_X1 U10820 ( .A(n9104), .B(n9102), .ZN(n10221) );
  INV_X1 U10821 ( .A(n10221), .ZN(n9061) );
  INV_X1 U10822 ( .A(n9091), .ZN(n9051) );
  INV_X1 U10823 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9050) );
  NAND2_X1 U10824 ( .A1(n9051), .A2(n9050), .ZN(n9111) );
  NAND2_X1 U10825 ( .A1(n9111), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9052) );
  XNOR2_X1 U10826 ( .A(n9052), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10222) );
  INV_X1 U10827 ( .A(n15157), .ZN(n15164) );
  AOI22_X1 U10828 ( .A1(n10222), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n15164), .ZN(n9053) );
  OAI21_X1 U10829 ( .B1(n9061), .B2(n15167), .A(n9053), .ZN(P1_U3350) );
  INV_X1 U10830 ( .A(n9054), .ZN(n9100) );
  NAND2_X1 U10831 ( .A1(n9100), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9055) );
  MUX2_X1 U10832 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9055), .S(
        P1_IR_REG_2__SCAN_IN), .Z(n9056) );
  NAND2_X1 U10833 ( .A1(n9056), .A2(n9089), .ZN(n14781) );
  OAI222_X1 U10834 ( .A1(n15157), .A2(n9058), .B1(n15167), .B2(n9057), .C1(
        P1_U3086), .C2(n14781), .ZN(P1_U3353) );
  INV_X1 U10835 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9062) );
  NOR2_X1 U10836 ( .A1(n9059), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n9109) );
  OR2_X1 U10837 ( .A1(n9109), .A2(n14582), .ZN(n9060) );
  XNOR2_X1 U10838 ( .A(n9060), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9958) );
  INV_X1 U10839 ( .A(n9958), .ZN(n15421) );
  OAI222_X1 U10840 ( .A1(n14588), .A2(n9062), .B1(n14593), .B2(n9061), .C1(
        P2_U3088), .C2(n15421), .ZN(P2_U3322) );
  INV_X1 U10841 ( .A(n9063), .ZN(n9064) );
  INV_X1 U10842 ( .A(n10076), .ZN(n9065) );
  NAND2_X1 U10843 ( .A1(n9065), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13078) );
  NAND2_X1 U10844 ( .A1(n9337), .A2(n13078), .ZN(n9079) );
  INV_X1 U10845 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9069) );
  NAND2_X1 U10846 ( .A1(n9072), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n9073) );
  OR2_X1 U10847 ( .A1(n9074), .A2(n9073), .ZN(n9076) );
  XNOR2_X1 U10848 ( .A(P1_IR_REG_31__SCAN_IN), .B(P1_IR_REG_27__SCAN_IN), .ZN(
        n9075) );
  NAND2_X1 U10849 ( .A1(n9079), .A2(n12008), .ZN(n9088) );
  NAND2_X1 U10850 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n9080) );
  NAND2_X1 U10851 ( .A1(n9080), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9081) );
  OAI21_X1 U10852 ( .B1(n9082), .B2(P1_IR_REG_31__SCAN_IN), .A(n9081), .ZN(
        n9083) );
  NAND2_X1 U10854 ( .A1(n15170), .A2(n12800), .ZN(n13002) );
  OR2_X1 U10855 ( .A1(n9337), .A2(n13002), .ZN(n9087) );
  AND2_X1 U10856 ( .A1(n9088), .A2(n9087), .ZN(n14842) );
  NOR2_X1 U10857 ( .A1(n14797), .A2(P1_U4016), .ZN(P1_U3085) );
  NAND2_X1 U10858 ( .A1(n9089), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9090) );
  MUX2_X1 U10859 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9090), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n9092) );
  AND2_X1 U10860 ( .A1(n9092), .A2(n9091), .ZN(n14788) );
  INV_X1 U10861 ( .A(n14788), .ZN(n9093) );
  OAI222_X1 U10862 ( .A1(n15157), .A2(n9094), .B1(n15167), .B2(n10040), .C1(
        P1_U3086), .C2(n9093), .ZN(P1_U3352) );
  NAND2_X1 U10863 ( .A1(n15161), .A2(P1_B_REG_SCAN_IN), .ZN(n9095) );
  MUX2_X1 U10864 ( .A(n9095), .B(P1_B_REG_SCAN_IN), .S(n15165), .Z(n9096) );
  INV_X1 U10865 ( .A(n15159), .ZN(n9097) );
  NAND2_X1 U10866 ( .A1(n9096), .A2(n9097), .ZN(n9430) );
  INV_X1 U10867 ( .A(n9337), .ZN(n10537) );
  NAND2_X2 U10868 ( .A1(n9430), .A2(n10537), .ZN(n15172) );
  NAND2_X1 U10869 ( .A1(n15172), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9098) );
  OAI21_X1 U10870 ( .B1(n15172), .B2(n9329), .A(n9098), .ZN(P1_U3445) );
  NAND2_X1 U10871 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9099) );
  MUX2_X1 U10872 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9099), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n9101) );
  NAND2_X1 U10873 ( .A1(n9101), .A2(n9100), .ZN(n14758) );
  INV_X1 U10874 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9285) );
  OAI222_X1 U10875 ( .A1(n15167), .A2(n9615), .B1(n14758), .B2(P1_U3086), .C1(
        n9285), .C2(n15157), .ZN(P1_U3354) );
  INV_X1 U10876 ( .A(n9102), .ZN(n9103) );
  NAND2_X1 U10877 ( .A1(n9104), .A2(n9103), .ZN(n9107) );
  NAND2_X1 U10878 ( .A1(n9105), .A2(SI_5_), .ZN(n9106) );
  MUX2_X1 U10879 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n8987), .Z(n9132) );
  XNOR2_X1 U10880 ( .A(n9132), .B(SI_6_), .ZN(n9129) );
  INV_X1 U10881 ( .A(n10261), .ZN(n9113) );
  INV_X1 U10882 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9108) );
  XNOR2_X1 U10883 ( .A(n9135), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10004) );
  INV_X1 U10884 ( .A(n10004), .ZN(n9681) );
  OAI222_X1 U10885 ( .A1(n14588), .A2(n9110), .B1(n14593), .B2(n9113), .C1(
        P2_U3088), .C2(n9681), .ZN(P2_U3321) );
  NAND2_X1 U10886 ( .A1(n9138), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9112) );
  XNOR2_X1 U10887 ( .A(n9112), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10262) );
  INV_X1 U10888 ( .A(n10262), .ZN(n9204) );
  OAI222_X1 U10889 ( .A1(n15157), .A2(n9114), .B1(n15167), .B2(n9113), .C1(
        P1_U3086), .C2(n9204), .ZN(P1_U3349) );
  NAND2_X1 U10890 ( .A1(n10312), .A2(n9116), .ZN(n9115) );
  OAI21_X1 U10891 ( .B1(n9117), .B2(n9116), .A(n9115), .ZN(P3_U3377) );
  INV_X1 U10892 ( .A(n9118), .ZN(n9119) );
  OAI222_X1 U10893 ( .A1(P3_U3151), .A2(n13613), .B1(n13083), .B2(n15208), 
        .C1(n13082), .C2(n9119), .ZN(P3_U3284) );
  OAI222_X1 U10894 ( .A1(P3_U3151), .A2(n15711), .B1(n13083), .B2(n15319), 
        .C1(n13082), .C2(n9120), .ZN(P3_U3283) );
  NOR2_X1 U10895 ( .A1(n15154), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9121) );
  NOR2_X1 U10896 ( .A1(n15151), .A2(n9121), .ZN(n14772) );
  INV_X1 U10897 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n15836) );
  NAND2_X1 U10898 ( .A1(n15154), .A2(n15836), .ZN(n9122) );
  NAND2_X1 U10899 ( .A1(n14772), .A2(n9122), .ZN(n9123) );
  INV_X1 U10900 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14760) );
  MUX2_X1 U10901 ( .A(n14772), .B(n9123), .S(n14760), .Z(n9128) );
  INV_X1 U10902 ( .A(n13002), .ZN(n9335) );
  OAI21_X1 U10903 ( .B1(n9337), .B2(n9335), .A(n13078), .ZN(n9124) );
  NAND2_X1 U10904 ( .A1(n9124), .A2(n12049), .ZN(n9166) );
  AOI22_X1 U10905 ( .A1(n14797), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9127) );
  INV_X1 U10906 ( .A(n9166), .ZN(n9125) );
  NAND3_X1 U10907 ( .A1(n14834), .A2(P1_IR_REG_0__SCAN_IN), .A3(n15836), .ZN(
        n9126) );
  OAI211_X1 U10908 ( .C1(n9128), .C2(n9166), .A(n9127), .B(n9126), .ZN(
        P1_U3243) );
  INV_X1 U10909 ( .A(n9129), .ZN(n9130) );
  NAND2_X1 U10910 ( .A1(n9132), .A2(SI_6_), .ZN(n9133) );
  MUX2_X1 U10911 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n13007), .Z(n9175) );
  XNOR2_X1 U10912 ( .A(n9175), .B(SI_7_), .ZN(n9172) );
  XNOR2_X1 U10913 ( .A(n9174), .B(n9172), .ZN(n10472) );
  INV_X1 U10914 ( .A(n10472), .ZN(n9140) );
  INV_X1 U10915 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n9134) );
  NAND2_X1 U10916 ( .A1(n9135), .A2(n9134), .ZN(n9136) );
  NAND2_X1 U10917 ( .A1(n9136), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9176) );
  XNOR2_X1 U10918 ( .A(n9176), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10325) );
  INV_X1 U10919 ( .A(n10325), .ZN(n9725) );
  OAI222_X1 U10920 ( .A1(n14588), .A2(n9137), .B1(n14593), .B2(n9140), .C1(
        P2_U3088), .C2(n9725), .ZN(P2_U3320) );
  INV_X1 U10921 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9141) );
  OAI21_X1 U10922 ( .B1(n9138), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9139) );
  XNOR2_X1 U10923 ( .A(n9139), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10473) );
  INV_X1 U10924 ( .A(n10473), .ZN(n9219) );
  OAI222_X1 U10925 ( .A1(n15157), .A2(n9141), .B1(n15167), .B2(n9140), .C1(
        P1_U3086), .C2(n9219), .ZN(P1_U3348) );
  INV_X1 U10926 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9142) );
  MUX2_X1 U10927 ( .A(n9142), .B(P1_REG2_REG_2__SCAN_IN), .S(n14781), .Z(
        n14774) );
  XNOR2_X1 U10928 ( .A(n14758), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n14756) );
  AND2_X1 U10929 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14768) );
  NAND2_X1 U10930 ( .A1(n14756), .A2(n14768), .ZN(n14755) );
  INV_X1 U10931 ( .A(n14758), .ZN(n14757) );
  NAND2_X1 U10932 ( .A1(n14757), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9143) );
  NAND2_X1 U10933 ( .A1(n14755), .A2(n9143), .ZN(n14773) );
  NAND2_X1 U10934 ( .A1(n14774), .A2(n14773), .ZN(n14790) );
  INV_X1 U10935 ( .A(n14781), .ZN(n9311) );
  NAND2_X1 U10936 ( .A1(n9311), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14789) );
  NAND2_X1 U10937 ( .A1(n14790), .A2(n14789), .ZN(n9145) );
  INV_X1 U10938 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10627) );
  MUX2_X1 U10939 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10627), .S(n14788), .Z(
        n9144) );
  NAND2_X1 U10940 ( .A1(n9145), .A2(n9144), .ZN(n14812) );
  NAND2_X1 U10941 ( .A1(n14788), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n14811) );
  NAND2_X1 U10942 ( .A1(n14812), .A2(n14811), .ZN(n9147) );
  INV_X1 U10943 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n14809) );
  MUX2_X1 U10944 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n14809), .S(n14808), .Z(
        n9146) );
  NAND2_X1 U10945 ( .A1(n9147), .A2(n9146), .ZN(n14814) );
  NAND2_X1 U10946 ( .A1(n14808), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9185) );
  INV_X1 U10947 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9148) );
  MUX2_X1 U10948 ( .A(n9148), .B(P1_REG2_REG_5__SCAN_IN), .S(n10222), .Z(n9184) );
  AOI21_X1 U10949 ( .B1(n14814), .B2(n9185), .A(n9184), .ZN(n9187) );
  AOI21_X1 U10950 ( .B1(n10222), .B2(P1_REG2_REG_5__SCAN_IN), .A(n9187), .ZN(
        n9198) );
  INV_X1 U10951 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9149) );
  MUX2_X1 U10952 ( .A(n9149), .B(P1_REG2_REG_6__SCAN_IN), .S(n10262), .Z(n9197) );
  NOR2_X1 U10953 ( .A1(n9198), .A2(n9197), .ZN(n9196) );
  AOI21_X1 U10954 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n10262), .A(n9196), .ZN(
        n9213) );
  INV_X1 U10955 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9150) );
  MUX2_X1 U10956 ( .A(n9150), .B(P1_REG2_REG_7__SCAN_IN), .S(n10473), .Z(n9212) );
  NOR2_X1 U10957 ( .A1(n9213), .A2(n9212), .ZN(n9211) );
  NOR2_X1 U10958 ( .A1(n9219), .A2(n9150), .ZN(n9156) );
  INV_X1 U10959 ( .A(n9156), .ZN(n9154) );
  INV_X1 U10960 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9152) );
  NAND2_X1 U10961 ( .A1(n7923), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9151) );
  XNOR2_X1 U10962 ( .A(n9151), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10732) );
  MUX2_X1 U10963 ( .A(n9152), .B(P1_REG2_REG_8__SCAN_IN), .S(n10732), .Z(n9153) );
  NAND2_X1 U10964 ( .A1(n9154), .A2(n9153), .ZN(n9157) );
  MUX2_X1 U10965 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n9152), .S(n10732), .Z(n9155) );
  OAI21_X1 U10966 ( .B1(n9211), .B2(n9156), .A(n9155), .ZN(n9259) );
  OR3_X1 U10967 ( .A1(n9166), .A2(n15154), .A3(n15151), .ZN(n14829) );
  OAI211_X1 U10968 ( .C1(n9211), .C2(n9157), .A(n9259), .B(n14833), .ZN(n9171)
         );
  INV_X1 U10969 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n16018) );
  MUX2_X1 U10970 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n16018), .S(n10732), .Z(
        n9165) );
  INV_X1 U10971 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9158) );
  MUX2_X1 U10972 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9158), .S(n14788), .Z(
        n14786) );
  XNOR2_X1 U10973 ( .A(n14781), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n14776) );
  NAND2_X1 U10974 ( .A1(n14757), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9161) );
  INV_X1 U10975 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n15859) );
  NAND2_X1 U10976 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9159) );
  AOI21_X1 U10977 ( .B1(n14758), .B2(n15859), .A(n9159), .ZN(n9160) );
  NAND2_X1 U10978 ( .A1(n9161), .A2(n9160), .ZN(n14762) );
  NAND2_X1 U10979 ( .A1(n14762), .A2(n9161), .ZN(n14775) );
  NAND2_X1 U10980 ( .A1(n14776), .A2(n14775), .ZN(n9163) );
  NAND2_X1 U10981 ( .A1(n9311), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9162) );
  NAND2_X1 U10982 ( .A1(n9163), .A2(n9162), .ZN(n14785) );
  NAND2_X1 U10983 ( .A1(n14786), .A2(n14785), .ZN(n14805) );
  NAND2_X1 U10984 ( .A1(n14788), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n14804) );
  INV_X1 U10985 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n15960) );
  MUX2_X1 U10986 ( .A(n15960), .B(P1_REG1_REG_4__SCAN_IN), .S(n14808), .Z(
        n14803) );
  AOI21_X1 U10987 ( .B1(n14805), .B2(n14804), .A(n14803), .ZN(n14802) );
  AOI21_X1 U10988 ( .B1(n14808), .B2(P1_REG1_REG_4__SCAN_IN), .A(n14802), .ZN(
        n9182) );
  INV_X1 U10989 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n15980) );
  MUX2_X1 U10990 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n15980), .S(n10222), .Z(
        n9183) );
  NAND2_X1 U10991 ( .A1(n9182), .A2(n9183), .ZN(n9181) );
  OAI21_X1 U10992 ( .B1(n10222), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9181), .ZN(
        n9194) );
  INV_X1 U10993 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10288) );
  MUX2_X1 U10994 ( .A(n10288), .B(P1_REG1_REG_6__SCAN_IN), .S(n10262), .Z(
        n9193) );
  OR2_X1 U10995 ( .A1(n9194), .A2(n9193), .ZN(n9208) );
  NAND2_X1 U10996 ( .A1(n10262), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9207) );
  INV_X1 U10997 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10501) );
  MUX2_X1 U10998 ( .A(n10501), .B(P1_REG1_REG_7__SCAN_IN), .S(n10473), .Z(
        n9206) );
  AOI21_X1 U10999 ( .B1(n9208), .B2(n9207), .A(n9206), .ZN(n9205) );
  AOI21_X1 U11000 ( .B1(n10473), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9205), .ZN(
        n9164) );
  NAND2_X1 U11001 ( .A1(n9164), .A2(n9165), .ZN(n9265) );
  OAI21_X1 U11002 ( .B1(n9165), .B2(n9164), .A(n9265), .ZN(n9169) );
  INV_X1 U11003 ( .A(n15151), .ZN(n14769) );
  NAND2_X1 U11004 ( .A1(n14787), .A2(n10732), .ZN(n9167) );
  NAND2_X1 U11005 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n10822) );
  OAI211_X1 U11006 ( .C1(n14842), .C2(n15533), .A(n9167), .B(n10822), .ZN(
        n9168) );
  AOI21_X1 U11007 ( .B1(n9169), .B2(n14834), .A(n9168), .ZN(n9170) );
  NAND2_X1 U11008 ( .A1(n9171), .A2(n9170), .ZN(P1_U3251) );
  INV_X1 U11009 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9178) );
  INV_X1 U11010 ( .A(n9172), .ZN(n9173) );
  MUX2_X1 U11011 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n7178), .Z(n9352) );
  XNOR2_X1 U11012 ( .A(n9352), .B(SI_8_), .ZN(n9350) );
  XNOR2_X1 U11013 ( .A(n9351), .B(n9350), .ZN(n10731) );
  INV_X1 U11014 ( .A(n10731), .ZN(n9179) );
  INV_X1 U11015 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n9648) );
  NAND2_X1 U11016 ( .A1(n9176), .A2(n9648), .ZN(n9177) );
  NAND2_X1 U11017 ( .A1(n9177), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9355) );
  XNOR2_X1 U11018 ( .A(n9355), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10447) );
  INV_X1 U11019 ( .A(n10447), .ZN(n9738) );
  OAI222_X1 U11020 ( .A1(n14588), .A2(n9178), .B1(n14593), .B2(n9179), .C1(
        P2_U3088), .C2(n9738), .ZN(P2_U3319) );
  INV_X1 U11021 ( .A(n10732), .ZN(n9261) );
  OAI222_X1 U11022 ( .A1(n15157), .A2(n9180), .B1(n15167), .B2(n9179), .C1(
        P1_U3086), .C2(n9261), .ZN(P1_U3347) );
  OAI21_X1 U11023 ( .B1(n9183), .B2(n9182), .A(n9181), .ZN(n9191) );
  AND3_X1 U11024 ( .A1(n14814), .A2(n9185), .A3(n9184), .ZN(n9186) );
  NOR3_X1 U11025 ( .A1(n14829), .A2(n9187), .A3(n9186), .ZN(n9190) );
  NAND2_X1 U11026 ( .A1(n14787), .A2(n10222), .ZN(n9188) );
  NAND2_X1 U11027 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10244) );
  OAI211_X1 U11028 ( .C1(n14842), .C2(n15527), .A(n9188), .B(n10244), .ZN(
        n9189) );
  AOI211_X1 U11029 ( .C1(n14834), .C2(n9191), .A(n9190), .B(n9189), .ZN(n9192)
         );
  INV_X1 U11030 ( .A(n9192), .ZN(P1_U3248) );
  NAND2_X1 U11031 ( .A1(n9194), .A2(n9193), .ZN(n9195) );
  NAND3_X1 U11032 ( .A1(n14834), .A2(n9208), .A3(n9195), .ZN(n9203) );
  NAND2_X1 U11033 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n10388) );
  AOI211_X1 U11034 ( .C1(n9198), .C2(n9197), .A(n9196), .B(n14829), .ZN(n9199)
         );
  INV_X1 U11035 ( .A(n9199), .ZN(n9200) );
  NAND2_X1 U11036 ( .A1(n10388), .A2(n9200), .ZN(n9201) );
  AOI21_X1 U11037 ( .B1(n14797), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n9201), .ZN(
        n9202) );
  OAI211_X1 U11038 ( .C1(n14828), .C2(n9204), .A(n9203), .B(n9202), .ZN(
        P1_U3249) );
  INV_X1 U11039 ( .A(n9205), .ZN(n9210) );
  NAND3_X1 U11040 ( .A1(n9208), .A2(n9207), .A3(n9206), .ZN(n9209) );
  NAND3_X1 U11041 ( .A1(n14834), .A2(n9210), .A3(n9209), .ZN(n9218) );
  NAND2_X1 U11042 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n10601) );
  AOI211_X1 U11043 ( .C1(n9213), .C2(n9212), .A(n9211), .B(n14829), .ZN(n9214)
         );
  INV_X1 U11044 ( .A(n9214), .ZN(n9215) );
  NAND2_X1 U11045 ( .A1(n10601), .A2(n9215), .ZN(n9216) );
  AOI21_X1 U11046 ( .B1(n14797), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n9216), .ZN(
        n9217) );
  OAI211_X1 U11047 ( .C1(n14828), .C2(n9219), .A(n9218), .B(n9217), .ZN(
        P1_U3250) );
  NOR2_X1 U11048 ( .A1(n9220), .A2(n14016), .ZN(n9222) );
  INV_X1 U11049 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n9221) );
  NOR2_X1 U11050 ( .A1(n9250), .A2(n9221), .ZN(P3_U3260) );
  CLKBUF_X1 U11051 ( .A(n9222), .Z(n9250) );
  INV_X1 U11052 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9223) );
  NOR2_X1 U11053 ( .A1(n9250), .A2(n9223), .ZN(P3_U3259) );
  INV_X1 U11054 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n9224) );
  NOR2_X1 U11055 ( .A1(n9222), .A2(n9224), .ZN(P3_U3258) );
  INV_X1 U11056 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9225) );
  NOR2_X1 U11057 ( .A1(n9250), .A2(n9225), .ZN(P3_U3255) );
  INV_X1 U11058 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9226) );
  NOR2_X1 U11059 ( .A1(n9250), .A2(n9226), .ZN(P3_U3254) );
  INV_X1 U11060 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n9227) );
  NOR2_X1 U11061 ( .A1(n9250), .A2(n9227), .ZN(P3_U3253) );
  INV_X1 U11062 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9228) );
  NOR2_X1 U11063 ( .A1(n9250), .A2(n9228), .ZN(P3_U3257) );
  INV_X1 U11064 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n9229) );
  NOR2_X1 U11065 ( .A1(n9250), .A2(n9229), .ZN(P3_U3256) );
  INV_X1 U11066 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n9230) );
  NOR2_X1 U11067 ( .A1(n9250), .A2(n9230), .ZN(P3_U3250) );
  INV_X1 U11068 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9231) );
  NOR2_X1 U11069 ( .A1(n9250), .A2(n9231), .ZN(P3_U3263) );
  INV_X1 U11070 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n9232) );
  NOR2_X1 U11071 ( .A1(n9250), .A2(n9232), .ZN(P3_U3249) );
  INV_X1 U11072 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9233) );
  NOR2_X1 U11073 ( .A1(n9250), .A2(n9233), .ZN(P3_U3248) );
  INV_X1 U11074 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9234) );
  NOR2_X1 U11075 ( .A1(n9250), .A2(n9234), .ZN(P3_U3247) );
  INV_X1 U11076 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n9235) );
  NOR2_X1 U11077 ( .A1(n9250), .A2(n9235), .ZN(P3_U3246) );
  INV_X1 U11078 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n9236) );
  NOR2_X1 U11079 ( .A1(n9222), .A2(n9236), .ZN(P3_U3245) );
  INV_X1 U11080 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n9237) );
  NOR2_X1 U11081 ( .A1(n9222), .A2(n9237), .ZN(P3_U3234) );
  INV_X1 U11082 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n9238) );
  NOR2_X1 U11083 ( .A1(n9222), .A2(n9238), .ZN(P3_U3244) );
  INV_X1 U11084 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n9239) );
  NOR2_X1 U11085 ( .A1(n9222), .A2(n9239), .ZN(P3_U3243) );
  INV_X1 U11086 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n9240) );
  NOR2_X1 U11087 ( .A1(n9222), .A2(n9240), .ZN(P3_U3242) );
  INV_X1 U11088 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n9241) );
  NOR2_X1 U11089 ( .A1(n9222), .A2(n9241), .ZN(P3_U3241) );
  INV_X1 U11090 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9242) );
  NOR2_X1 U11091 ( .A1(n9250), .A2(n9242), .ZN(P3_U3252) );
  INV_X1 U11092 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9243) );
  NOR2_X1 U11093 ( .A1(n9222), .A2(n9243), .ZN(P3_U3262) );
  INV_X1 U11094 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9244) );
  NOR2_X1 U11095 ( .A1(n9250), .A2(n9244), .ZN(P3_U3261) );
  INV_X1 U11096 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9245) );
  NOR2_X1 U11097 ( .A1(n9222), .A2(n9245), .ZN(P3_U3237) );
  INV_X1 U11098 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n9246) );
  NOR2_X1 U11099 ( .A1(n9222), .A2(n9246), .ZN(P3_U3236) );
  INV_X1 U11100 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9247) );
  NOR2_X1 U11101 ( .A1(n9222), .A2(n9247), .ZN(P3_U3235) );
  INV_X1 U11102 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n9248) );
  NOR2_X1 U11103 ( .A1(n9250), .A2(n9248), .ZN(P3_U3238) );
  INV_X1 U11104 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n9249) );
  NOR2_X1 U11105 ( .A1(n9250), .A2(n9249), .ZN(P3_U3251) );
  INV_X1 U11106 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n9251) );
  NOR2_X1 U11107 ( .A1(n9250), .A2(n9251), .ZN(P3_U3239) );
  INV_X1 U11108 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n9252) );
  NOR2_X1 U11109 ( .A1(n9250), .A2(n9252), .ZN(P3_U3240) );
  OAI222_X1 U11110 ( .A1(P3_U3151), .A2(n9254), .B1(n13083), .B2(n15311), .C1(
        n13082), .C2(n9253), .ZN(P3_U3282) );
  NAND2_X1 U11111 ( .A1(n10732), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9258) );
  INV_X1 U11112 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9385) );
  NAND2_X1 U11113 ( .A1(n10442), .A2(n9255), .ZN(n9374) );
  NAND2_X1 U11114 ( .A1(n9374), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9256) );
  XNOR2_X1 U11115 ( .A(n9256), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10907) );
  MUX2_X1 U11116 ( .A(n9385), .B(P1_REG2_REG_9__SCAN_IN), .S(n10907), .Z(n9257) );
  AOI21_X1 U11117 ( .B1(n9259), .B2(n9258), .A(n9257), .ZN(n9393) );
  NAND3_X1 U11118 ( .A1(n9259), .A2(n9258), .A3(n9257), .ZN(n9260) );
  NAND2_X1 U11119 ( .A1(n9260), .A2(n14833), .ZN(n9271) );
  INV_X1 U11120 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n15551) );
  NAND2_X1 U11121 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n11129) );
  OAI21_X1 U11122 ( .B1(n14842), .B2(n15551), .A(n11129), .ZN(n9269) );
  NAND2_X1 U11123 ( .A1(n9261), .A2(n16018), .ZN(n9263) );
  INV_X1 U11124 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9262) );
  MUX2_X1 U11125 ( .A(n9262), .B(P1_REG1_REG_9__SCAN_IN), .S(n10907), .Z(n9264) );
  AOI21_X1 U11126 ( .B1(n9265), .B2(n9263), .A(n9264), .ZN(n9377) );
  INV_X1 U11127 ( .A(n9377), .ZN(n9267) );
  NAND3_X1 U11128 ( .A1(n9265), .A2(n9264), .A3(n9263), .ZN(n9266) );
  INV_X1 U11129 ( .A(n14834), .ZN(n10134) );
  AOI21_X1 U11130 ( .B1(n9267), .B2(n9266), .A(n10134), .ZN(n9268) );
  AOI211_X1 U11131 ( .C1(n14787), .C2(n10907), .A(n9269), .B(n9268), .ZN(n9270) );
  OAI21_X1 U11132 ( .B1(n9393), .B2(n9271), .A(n9270), .ZN(P1_U3252) );
  OAI222_X1 U11133 ( .A1(P3_U3151), .A2(n13634), .B1(n13083), .B2(n15318), 
        .C1(n13082), .C2(n9272), .ZN(P3_U3281) );
  NAND2_X1 U11134 ( .A1(n9273), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9274) );
  NAND2_X1 U11135 ( .A1(n9339), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9277) );
  NAND2_X1 U11136 ( .A1(n9340), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9276) );
  NAND2_X1 U11137 ( .A1(n12095), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n9280) );
  NAND2_X1 U11138 ( .A1(n7204), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9281) );
  MUX2_X1 U11139 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9281), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n9283) );
  INV_X1 U11140 ( .A(n12808), .ZN(n10642) );
  NAND2_X1 U11141 ( .A1(n12049), .A2(n9540), .ZN(n9310) );
  NAND2_X1 U11142 ( .A1(n9286), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9287) );
  NAND2_X1 U11143 ( .A1(n15170), .A2(n14836), .ZN(n9288) );
  XNOR2_X1 U11144 ( .A(n9289), .B(n12526), .ZN(n9304) );
  NOR2_X4 U11145 ( .A1(n15832), .A2(n13017), .ZN(n15041) );
  NAND2_X1 U11146 ( .A1(n15041), .A2(n14836), .ZN(n14952) );
  OR2_X1 U11147 ( .A1(n9416), .A2(n12524), .ZN(n9291) );
  NAND2_X1 U11148 ( .A1(n10225), .A2(n10936), .ZN(n9290) );
  NAND2_X1 U11149 ( .A1(n9339), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9295) );
  NAND2_X1 U11150 ( .A1(n12095), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9294) );
  NAND2_X1 U11151 ( .A1(n12014), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U11152 ( .A1(n9340), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9292) );
  OR2_X1 U11153 ( .A1(n12809), .A2(n12525), .ZN(n9301) );
  NAND3_X1 U11154 ( .A1(n7178), .A2(SI_0_), .A3(P2_DATAO_REG_0__SCAN_IN), .ZN(
        n9299) );
  INV_X1 U11155 ( .A(SI_0_), .ZN(n9297) );
  OAI21_X1 U11156 ( .B1(n9540), .B2(n9297), .A(n9296), .ZN(n9298) );
  AND2_X1 U11157 ( .A1(n9299), .A2(n9298), .ZN(n15171) );
  MUX2_X1 U11158 ( .A(P1_IR_REG_0__SCAN_IN), .B(n15171), .S(n12049), .Z(n10935) );
  INV_X1 U11159 ( .A(n10077), .ZN(n9302) );
  AOI22_X1 U11160 ( .A1(n12514), .A2(n10935), .B1(n9302), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n9300) );
  AOI22_X1 U11161 ( .A1(n10225), .A2(n10935), .B1(n9302), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n9303) );
  OAI21_X1 U11162 ( .B1(n12524), .B2(n12809), .A(n9303), .ZN(n9362) );
  OAI21_X1 U11163 ( .B1(n9363), .B2(n12526), .A(n9361), .ZN(n9366) );
  NAND2_X1 U11164 ( .A1(n12095), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9309) );
  NAND2_X1 U11165 ( .A1(n9339), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9308) );
  NAND2_X1 U11166 ( .A1(n9340), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9307) );
  NAND2_X1 U11167 ( .A1(n12014), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9306) );
  INV_X2 U11168 ( .A(n9310), .ZN(n10053) );
  NAND2_X1 U11169 ( .A1(n9541), .A2(n10051), .ZN(n9312) );
  INV_X2 U11170 ( .A(n12802), .ZN(n12805) );
  OAI22_X1 U11171 ( .A1(n10624), .A2(n12525), .B1(n12805), .B2(n12523), .ZN(
        n9313) );
  XNOR2_X1 U11172 ( .A(n9313), .B(n12526), .ZN(n10046) );
  OR2_X1 U11173 ( .A1(n10624), .A2(n12524), .ZN(n9315) );
  NAND2_X1 U11174 ( .A1(n10225), .A2(n12802), .ZN(n9314) );
  NAND2_X1 U11175 ( .A1(n9315), .A2(n9314), .ZN(n10045) );
  XNOR2_X1 U11176 ( .A(n10046), .B(n10045), .ZN(n10047) );
  XNOR2_X1 U11177 ( .A(n10044), .B(n10047), .ZN(n9349) );
  INV_X1 U11178 ( .A(n9430), .ZN(n9432) );
  NOR4_X1 U11179 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n9319) );
  NOR4_X1 U11180 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n9318) );
  NOR4_X1 U11181 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n9317) );
  NOR4_X1 U11182 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n9316) );
  AND4_X1 U11183 ( .A1(n9319), .A2(n9318), .A3(n9317), .A4(n9316), .ZN(n9325)
         );
  NOR2_X1 U11184 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n9323) );
  NOR4_X1 U11185 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n9322) );
  NOR4_X1 U11186 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n9321) );
  NOR4_X1 U11187 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n9320) );
  AND4_X1 U11188 ( .A1(n9323), .A2(n9322), .A3(n9321), .A4(n9320), .ZN(n9324)
         );
  NAND2_X1 U11189 ( .A1(n9325), .A2(n9324), .ZN(n9431) );
  INV_X1 U11190 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9326) );
  OR2_X1 U11191 ( .A1(n9431), .A2(n9326), .ZN(n9328) );
  NAND2_X1 U11192 ( .A1(n15161), .A2(n15159), .ZN(n15143) );
  INV_X1 U11193 ( .A(n15143), .ZN(n9327) );
  AOI21_X1 U11194 ( .B1(n9432), .B2(n9328), .A(n9327), .ZN(n10533) );
  INV_X1 U11195 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9330) );
  NAND2_X1 U11196 ( .A1(n10533), .A2(n10534), .ZN(n9338) );
  NAND2_X1 U11197 ( .A1(n12993), .A2(n14836), .ZN(n9334) );
  NAND2_X1 U11198 ( .A1(n16058), .A2(n13002), .ZN(n9331) );
  OR2_X1 U11199 ( .A1(n9337), .A2(n9331), .ZN(n9332) );
  INV_X1 U11200 ( .A(n10536), .ZN(n9333) );
  NAND2_X1 U11201 ( .A1(n9338), .A2(n9333), .ZN(n10080) );
  AND2_X1 U11202 ( .A1(n9335), .A2(n9334), .ZN(n9336) );
  INV_X1 U11203 ( .A(n9336), .ZN(n10078) );
  NAND2_X1 U11204 ( .A1(n15921), .A2(n10078), .ZN(n9371) );
  OR2_X1 U11205 ( .A1(n9337), .A2(n9336), .ZN(n13075) );
  OR2_X1 U11206 ( .A1(n9416), .A2(n15003), .ZN(n9346) );
  INV_X1 U11207 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10623) );
  NAND2_X1 U11208 ( .A1(n12095), .A2(n10623), .ZN(n9344) );
  NAND2_X1 U11209 ( .A1(n9339), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9343) );
  NAND2_X1 U11210 ( .A1(n12014), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9342) );
  NAND2_X1 U11211 ( .A1(n9340), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9341) );
  NAND4_X1 U11212 ( .A1(n9344), .A2(n9343), .A3(n9342), .A4(n9341), .ZN(n14750) );
  OR2_X1 U11213 ( .A1(n13002), .A2(n14769), .ZN(n15005) );
  NAND2_X1 U11214 ( .A1(n14750), .A2(n14980), .ZN(n9345) );
  NAND2_X1 U11215 ( .A1(n9346), .A2(n9345), .ZN(n10896) );
  AOI22_X1 U11216 ( .A1(n9371), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n15927), .B2(
        n10896), .ZN(n9348) );
  NAND2_X1 U11217 ( .A1(n16129), .A2(n12802), .ZN(n9347) );
  OAI211_X1 U11218 ( .C1(n9349), .C2(n16123), .A(n9348), .B(n9347), .ZN(
        P1_U3237) );
  INV_X1 U11219 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9358) );
  NAND2_X1 U11220 ( .A1(n9352), .A2(SI_8_), .ZN(n9353) );
  MUX2_X1 U11221 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n7178), .Z(n9437) );
  INV_X1 U11222 ( .A(n10906), .ZN(n9359) );
  INV_X1 U11223 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n9354) );
  NAND2_X1 U11224 ( .A1(n9355), .A2(n9354), .ZN(n9356) );
  NAND2_X1 U11225 ( .A1(n9356), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9445) );
  XNOR2_X1 U11226 ( .A(n9445), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10551) );
  INV_X1 U11227 ( .A(n10551), .ZN(n9357) );
  OAI222_X1 U11228 ( .A1(n14588), .A2(n9358), .B1(n14593), .B2(n9359), .C1(
        P2_U3088), .C2(n9357), .ZN(P2_U3318) );
  INV_X1 U11229 ( .A(n10907), .ZN(n9386) );
  OAI222_X1 U11230 ( .A1(n15157), .A2(n9360), .B1(n15167), .B2(n9359), .C1(
        P1_U3086), .C2(n9386), .ZN(P1_U3346) );
  INV_X1 U11231 ( .A(n10935), .ZN(n15839) );
  OAI21_X1 U11232 ( .B1(n9363), .B2(n9362), .A(n9361), .ZN(n14767) );
  OR2_X1 U11233 ( .A1(n9416), .A2(n15005), .ZN(n15830) );
  OAI22_X1 U11234 ( .A1(n16123), .A2(n14767), .B1(n14725), .B2(n15830), .ZN(
        n9364) );
  AOI21_X1 U11235 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n9371), .A(n9364), .ZN(
        n9365) );
  OAI21_X1 U11236 ( .B1(n14731), .B2(n15839), .A(n9365), .ZN(P1_U3232) );
  XNOR2_X1 U11237 ( .A(n9367), .B(n9366), .ZN(n9368) );
  NAND2_X1 U11238 ( .A1(n9368), .A2(n14719), .ZN(n9373) );
  OR2_X1 U11239 ( .A1(n12809), .A2(n15003), .ZN(n9370) );
  OR2_X1 U11240 ( .A1(n10624), .A2(n15005), .ZN(n9369) );
  NAND2_X1 U11241 ( .A1(n9370), .A2(n9369), .ZN(n10941) );
  AOI22_X1 U11242 ( .A1(n9371), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n15927), .B2(
        n10941), .ZN(n9372) );
  OAI211_X1 U11243 ( .C1(n14731), .C2(n15854), .A(n9373), .B(n9372), .ZN(
        P1_U3222) );
  NAND2_X1 U11244 ( .A1(n9396), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9375) );
  XNOR2_X1 U11245 ( .A(n9375), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10998) );
  INV_X1 U11246 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9376) );
  NAND2_X1 U11247 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11301)
         );
  OAI21_X1 U11248 ( .B1(n14842), .B2(n9376), .A(n11301), .ZN(n9384) );
  AOI21_X1 U11249 ( .B1(n9262), .B2(n9386), .A(n9377), .ZN(n9379) );
  INV_X1 U11250 ( .A(n9379), .ZN(n9382) );
  INV_X1 U11251 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n11174) );
  MUX2_X1 U11252 ( .A(n11174), .B(P1_REG1_REG_10__SCAN_IN), .S(n10998), .Z(
        n9381) );
  MUX2_X1 U11253 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n11174), .S(n10998), .Z(
        n9378) );
  NAND2_X1 U11254 ( .A1(n9379), .A2(n9378), .ZN(n9401) );
  INV_X1 U11255 ( .A(n9401), .ZN(n9380) );
  AOI211_X1 U11256 ( .C1(n9382), .C2(n9381), .A(n10134), .B(n9380), .ZN(n9383)
         );
  AOI211_X1 U11257 ( .C1(n14787), .C2(n10998), .A(n9384), .B(n9383), .ZN(n9395) );
  NOR2_X1 U11258 ( .A1(n9386), .A2(n9385), .ZN(n9391) );
  INV_X1 U11259 ( .A(n9391), .ZN(n9389) );
  INV_X1 U11260 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9387) );
  MUX2_X1 U11261 ( .A(n9387), .B(P1_REG2_REG_10__SCAN_IN), .S(n10998), .Z(
        n9388) );
  NAND2_X1 U11262 ( .A1(n9389), .A2(n9388), .ZN(n9392) );
  MUX2_X1 U11263 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n9387), .S(n10998), .Z(
        n9390) );
  OAI21_X1 U11264 ( .B1(n9393), .B2(n9391), .A(n9390), .ZN(n9409) );
  OAI211_X1 U11265 ( .C1(n9393), .C2(n9392), .A(n9409), .B(n14833), .ZN(n9394)
         );
  NAND2_X1 U11266 ( .A1(n9395), .A2(n9394), .ZN(P1_U3253) );
  INV_X1 U11267 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9400) );
  INV_X1 U11268 ( .A(n9396), .ZN(n9398) );
  INV_X1 U11269 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9397) );
  NAND2_X1 U11270 ( .A1(n9398), .A2(n9397), .ZN(n9766) );
  NAND2_X1 U11271 ( .A1(n9766), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9399) );
  XNOR2_X1 U11272 ( .A(n9399), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11036) );
  MUX2_X1 U11273 ( .A(n9400), .B(P1_REG1_REG_11__SCAN_IN), .S(n11036), .Z(
        n9403) );
  INV_X1 U11274 ( .A(n10998), .ZN(n9442) );
  OAI21_X1 U11275 ( .B1(n11174), .B2(n9442), .A(n9401), .ZN(n9402) );
  NOR2_X1 U11276 ( .A1(n9402), .A2(n9403), .ZN(n10119) );
  AOI21_X1 U11277 ( .B1(n9403), .B2(n9402), .A(n10119), .ZN(n9414) );
  NOR2_X1 U11278 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11482), .ZN(n9405) );
  INV_X1 U11279 ( .A(n11036), .ZN(n10120) );
  NOR2_X1 U11280 ( .A1(n14828), .A2(n10120), .ZN(n9404) );
  AOI211_X1 U11281 ( .C1(P1_ADDR_REG_11__SCAN_IN), .C2(n14797), .A(n9405), .B(
        n9404), .ZN(n9413) );
  NAND2_X1 U11282 ( .A1(n10998), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9408) );
  INV_X1 U11283 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9406) );
  MUX2_X1 U11284 ( .A(n9406), .B(P1_REG2_REG_11__SCAN_IN), .S(n11036), .Z(
        n9407) );
  AOI21_X1 U11285 ( .B1(n9409), .B2(n9408), .A(n9407), .ZN(n10127) );
  INV_X1 U11286 ( .A(n10127), .ZN(n9411) );
  NAND3_X1 U11287 ( .A1(n9409), .A2(n9408), .A3(n9407), .ZN(n9410) );
  NAND3_X1 U11288 ( .A1(n9411), .A2(n14833), .A3(n9410), .ZN(n9412) );
  OAI211_X1 U11289 ( .C1(n9414), .C2(n10134), .A(n9413), .B(n9412), .ZN(
        P1_U3254) );
  INV_X1 U11290 ( .A(n15170), .ZN(n9415) );
  OAI21_X1 U11291 ( .B1(n9415), .B2(n12808), .A(n12526), .ZN(n10538) );
  NOR2_X1 U11292 ( .A1(n12809), .A2(n15839), .ZN(n10933) );
  NAND2_X1 U11293 ( .A1(n9416), .A2(n15854), .ZN(n9417) );
  NAND2_X1 U11294 ( .A1(n10624), .A2(n12805), .ZN(n10251) );
  NAND2_X1 U11295 ( .A1(n14751), .A2(n12802), .ZN(n9418) );
  NAND2_X1 U11296 ( .A1(n10251), .A2(n9418), .ZN(n13026) );
  XNOR2_X1 U11297 ( .A(n10250), .B(n13026), .ZN(n10903) );
  INV_X1 U11298 ( .A(n10903), .ZN(n9429) );
  NOR2_X1 U11299 ( .A1(n15170), .A2(n14836), .ZN(n9419) );
  NAND2_X1 U11300 ( .A1(n9419), .A2(n12993), .ZN(n15856) );
  INV_X1 U11301 ( .A(n10938), .ZN(n9421) );
  NAND2_X1 U11302 ( .A1(n10938), .A2(n12805), .ZN(n10620) );
  INV_X1 U11303 ( .A(n10620), .ZN(n9420) );
  AOI211_X1 U11304 ( .C1(n12802), .C2(n9421), .A(n15952), .B(n9420), .ZN(
        n10897) );
  AOI211_X1 U11305 ( .C1(n15948), .C2(n12802), .A(n10896), .B(n10897), .ZN(
        n9427) );
  NAND2_X1 U11306 ( .A1(n12809), .A2(n10935), .ZN(n13025) );
  INV_X1 U11307 ( .A(n13025), .ZN(n12814) );
  NAND2_X1 U11308 ( .A1(n13028), .A2(n12814), .ZN(n9422) );
  NAND2_X1 U11309 ( .A1(n9422), .A2(n12815), .ZN(n9423) );
  OR2_X1 U11310 ( .A1(n9423), .A2(n13026), .ZN(n9424) );
  NAND2_X1 U11311 ( .A1(n10272), .A2(n9424), .ZN(n10901) );
  NAND2_X1 U11312 ( .A1(n15170), .A2(n13059), .ZN(n12799) );
  NAND2_X1 U11313 ( .A1(n12800), .A2(n13017), .ZN(n9425) );
  NAND2_X1 U11314 ( .A1(n10901), .A2(n15955), .ZN(n9426) );
  OAI211_X1 U11315 ( .C1(n10903), .C2(n15856), .A(n9427), .B(n9426), .ZN(n9428) );
  AOI21_X1 U11316 ( .B1(n16034), .B2(n9429), .A(n9428), .ZN(n15902) );
  OAI21_X1 U11317 ( .B1(n9430), .B2(P1_D_REG_1__SCAN_IN), .A(n15143), .ZN(
        n9435) );
  NOR2_X1 U11318 ( .A1(n13075), .A2(n10536), .ZN(n9434) );
  NAND2_X1 U11319 ( .A1(n9432), .A2(n9431), .ZN(n9433) );
  NAND2_X1 U11320 ( .A1(n16066), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9436) );
  OAI21_X1 U11321 ( .B1(n15902), .B2(n16066), .A(n9436), .ZN(P1_U3530) );
  INV_X1 U11322 ( .A(n9437), .ZN(n9438) );
  MUX2_X1 U11323 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n7178), .Z(n9639) );
  XNOR2_X1 U11324 ( .A(n9639), .B(SI_10_), .ZN(n9636) );
  XNOR2_X1 U11325 ( .A(n9638), .B(n9636), .ZN(n10997) );
  INV_X1 U11326 ( .A(n10997), .ZN(n9447) );
  OAI222_X1 U11327 ( .A1(n15157), .A2(n9443), .B1(n15167), .B2(n9447), .C1(
        P1_U3086), .C2(n9442), .ZN(P1_U3345) );
  INV_X1 U11328 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9448) );
  INV_X1 U11329 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9444) );
  NAND2_X1 U11330 ( .A1(n9445), .A2(n9444), .ZN(n9446) );
  NAND2_X1 U11331 ( .A1(n9446), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9523) );
  XNOR2_X1 U11332 ( .A(n9523), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10687) );
  INV_X1 U11333 ( .A(n10687), .ZN(n9751) );
  OAI222_X1 U11334 ( .A1(n14588), .A2(n9448), .B1(n14593), .B2(n9447), .C1(
        P2_U3088), .C2(n9751), .ZN(P2_U3317) );
  INV_X1 U11335 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9449) );
  MUX2_X1 U11336 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n9449), .S(n14204), .Z(
        n14203) );
  INV_X1 U11337 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9450) );
  MUX2_X1 U11338 ( .A(n9450), .B(P2_REG1_REG_1__SCAN_IN), .S(n9706), .Z(n9452)
         );
  AND2_X1 U11339 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9451) );
  NAND2_X1 U11340 ( .A1(n9452), .A2(n9451), .ZN(n9698) );
  INV_X1 U11341 ( .A(n9706), .ZN(n9612) );
  NAND2_X1 U11342 ( .A1(n9612), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9453) );
  NAND2_X1 U11343 ( .A1(n9698), .A2(n9453), .ZN(n14202) );
  NAND2_X1 U11344 ( .A1(n14203), .A2(n14202), .ZN(n14201) );
  NAND2_X1 U11345 ( .A1(n14204), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9454) );
  NAND2_X1 U11346 ( .A1(n14201), .A2(n9454), .ZN(n15417) );
  INV_X1 U11347 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9455) );
  MUX2_X1 U11348 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9455), .S(n9878), .Z(n15416) );
  NAND2_X1 U11349 ( .A1(n15417), .A2(n15416), .ZN(n15415) );
  NAND2_X1 U11350 ( .A1(n9878), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9683) );
  NAND2_X1 U11351 ( .A1(n15415), .A2(n9683), .ZN(n9458) );
  INV_X1 U11352 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9456) );
  MUX2_X1 U11353 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9456), .S(n9884), .Z(n9457)
         );
  NAND2_X1 U11354 ( .A1(n9458), .A2(n9457), .ZN(n9685) );
  NAND2_X1 U11355 ( .A1(n9884), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9459) );
  NAND2_X1 U11356 ( .A1(n9685), .A2(n9459), .ZN(n15428) );
  INV_X1 U11357 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9460) );
  MUX2_X1 U11358 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9460), .S(n9958), .Z(n15427) );
  NAND2_X1 U11359 ( .A1(n15428), .A2(n15427), .ZN(n15426) );
  NAND2_X1 U11360 ( .A1(n9958), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9670) );
  NAND2_X1 U11361 ( .A1(n15426), .A2(n9670), .ZN(n9463) );
  INV_X1 U11362 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9461) );
  MUX2_X1 U11363 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9461), .S(n10004), .Z(n9462) );
  NAND2_X1 U11364 ( .A1(n9463), .A2(n9462), .ZN(n9672) );
  NAND2_X1 U11365 ( .A1(n10004), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9464) );
  NAND2_X1 U11366 ( .A1(n9672), .A2(n9464), .ZN(n9717) );
  INV_X1 U11367 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9465) );
  MUX2_X1 U11368 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9465), .S(n10325), .Z(n9716) );
  NAND2_X1 U11369 ( .A1(n9717), .A2(n9716), .ZN(n9715) );
  NAND2_X1 U11370 ( .A1(n10325), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9466) );
  NAND2_X1 U11371 ( .A1(n9715), .A2(n9466), .ZN(n9733) );
  INV_X1 U11372 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9467) );
  MUX2_X1 U11373 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9467), .S(n10447), .Z(n9732) );
  NAND2_X1 U11374 ( .A1(n9733), .A2(n9732), .ZN(n9731) );
  NAND2_X1 U11375 ( .A1(n10447), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9468) );
  NAND2_X1 U11376 ( .A1(n9731), .A2(n9468), .ZN(n9472) );
  INV_X1 U11377 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9469) );
  MUX2_X1 U11378 ( .A(n9469), .B(P2_REG1_REG_9__SCAN_IN), .S(n10551), .Z(n9471) );
  OR2_X1 U11379 ( .A1(n9472), .A2(n9471), .ZN(n9530) );
  INV_X1 U11380 ( .A(n9530), .ZN(n9470) );
  AOI21_X1 U11381 ( .B1(n9472), .B2(n9471), .A(n9470), .ZN(n9518) );
  NAND2_X1 U11382 ( .A1(n9473), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9475) );
  NAND2_X1 U11383 ( .A1(n8046), .A2(n7182), .ZN(n9593) );
  INV_X1 U11384 ( .A(n9593), .ZN(n9595) );
  NOR2_X1 U11386 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n9481) );
  NOR2_X1 U11387 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .ZN(n9480) );
  NOR2_X1 U11388 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n9479) );
  NAND4_X1 U11389 ( .A1(n9482), .A2(n9481), .A3(n9480), .A4(n9479), .ZN(n9486)
         );
  INV_X1 U11390 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n9483) );
  INV_X1 U11391 ( .A(n9484), .ZN(n9488) );
  NAND2_X2 U11392 ( .A1(n9488), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9485) );
  AOI21_X1 U11393 ( .B1(n9595), .B2(n9544), .A(n12234), .ZN(n9490) );
  NOR2_X1 U11394 ( .A1(n9492), .A2(P2_U3088), .ZN(n14590) );
  INV_X1 U11395 ( .A(n15473), .ZN(n14230) );
  INV_X1 U11396 ( .A(n13408), .ZN(n9493) );
  INV_X1 U11397 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9602) );
  MUX2_X1 U11398 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n9602), .S(n14204), .Z(
        n14208) );
  INV_X1 U11399 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9577) );
  MUX2_X1 U11400 ( .A(n9577), .B(P2_REG2_REG_1__SCAN_IN), .S(n9706), .Z(n9496)
         );
  AND2_X1 U11401 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9495) );
  NAND2_X1 U11402 ( .A1(n9496), .A2(n9495), .ZN(n9703) );
  NAND2_X1 U11403 ( .A1(n9612), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9497) );
  NAND2_X1 U11404 ( .A1(n9703), .A2(n9497), .ZN(n14207) );
  NAND2_X1 U11405 ( .A1(n14208), .A2(n14207), .ZN(n14206) );
  NAND2_X1 U11406 ( .A1(n14204), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9498) );
  NAND2_X1 U11407 ( .A1(n14206), .A2(n9498), .ZN(n15414) );
  INV_X1 U11408 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9587) );
  MUX2_X1 U11409 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n9587), .S(n9878), .Z(n15413) );
  NAND2_X1 U11410 ( .A1(n15414), .A2(n15413), .ZN(n15412) );
  NAND2_X1 U11411 ( .A1(n9878), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9689) );
  NAND2_X1 U11412 ( .A1(n15412), .A2(n9689), .ZN(n9500) );
  INV_X1 U11413 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10513) );
  MUX2_X1 U11414 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10513), .S(n9884), .Z(n9499) );
  NAND2_X1 U11415 ( .A1(n9500), .A2(n9499), .ZN(n9691) );
  NAND2_X1 U11416 ( .A1(n9884), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9501) );
  NAND2_X1 U11417 ( .A1(n9691), .A2(n9501), .ZN(n15425) );
  INV_X1 U11418 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9909) );
  MUX2_X1 U11419 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n9909), .S(n9958), .Z(n15424) );
  NAND2_X1 U11420 ( .A1(n15425), .A2(n15424), .ZN(n15423) );
  NAND2_X1 U11421 ( .A1(n9958), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9676) );
  NAND2_X1 U11422 ( .A1(n15423), .A2(n9676), .ZN(n9503) );
  INV_X1 U11423 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n9982) );
  MUX2_X1 U11424 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n9982), .S(n10004), .Z(n9502) );
  NAND2_X1 U11425 ( .A1(n9503), .A2(n9502), .ZN(n9678) );
  NAND2_X1 U11426 ( .A1(n10004), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9504) );
  NAND2_X1 U11427 ( .A1(n9678), .A2(n9504), .ZN(n9719) );
  INV_X1 U11428 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10010) );
  MUX2_X1 U11429 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10010), .S(n10325), .Z(
        n9718) );
  NAND2_X1 U11430 ( .A1(n9719), .A2(n9718), .ZN(n9728) );
  NAND2_X1 U11431 ( .A1(n10325), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9727) );
  NAND2_X1 U11432 ( .A1(n9728), .A2(n9727), .ZN(n9506) );
  INV_X1 U11433 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10347) );
  MUX2_X1 U11434 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10347), .S(n10447), .Z(
        n9505) );
  NAND2_X1 U11435 ( .A1(n9506), .A2(n9505), .ZN(n9730) );
  NAND2_X1 U11436 ( .A1(n10447), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9507) );
  NAND2_X1 U11437 ( .A1(n9730), .A2(n9507), .ZN(n9509) );
  INV_X1 U11438 ( .A(n9509), .ZN(n9511) );
  INV_X1 U11439 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n14432) );
  MUX2_X1 U11440 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n14432), .S(n10551), .Z(
        n9510) );
  MUX2_X1 U11441 ( .A(n14432), .B(P2_REG2_REG_9__SCAN_IN), .S(n10551), .Z(
        n9508) );
  OR2_X1 U11442 ( .A1(n9509), .A2(n9508), .ZN(n9520) );
  OAI21_X1 U11443 ( .B1(n9511), .B2(n9510), .A(n9520), .ZN(n9516) );
  INV_X1 U11444 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n15559) );
  OR2_X1 U11445 ( .A1(n9512), .A2(P2_U3088), .ZN(n11766) );
  NAND2_X1 U11446 ( .A1(n9512), .A2(n9492), .ZN(n15469) );
  INV_X1 U11447 ( .A(n15466), .ZN(n14205) );
  NAND2_X1 U11448 ( .A1(n14205), .A2(n10551), .ZN(n9514) );
  NAND2_X1 U11449 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n9513) );
  OAI211_X1 U11450 ( .C1(n15559), .C2(n11766), .A(n9514), .B(n9513), .ZN(n9515) );
  AOI21_X1 U11451 ( .B1(n15477), .B2(n9516), .A(n9515), .ZN(n9517) );
  OAI21_X1 U11452 ( .B1(n9518), .B2(n14230), .A(n9517), .ZN(P2_U3223) );
  OR2_X1 U11453 ( .A1(n10551), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9519) );
  NAND2_X1 U11454 ( .A1(n9520), .A2(n9519), .ZN(n9743) );
  INV_X1 U11455 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10786) );
  MUX2_X1 U11456 ( .A(n10786), .B(P2_REG2_REG_10__SCAN_IN), .S(n10687), .Z(
        n9744) );
  OR2_X1 U11457 ( .A1(n9743), .A2(n9744), .ZN(n9745) );
  NAND2_X1 U11458 ( .A1(n10687), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9521) );
  NAND2_X1 U11459 ( .A1(n9745), .A2(n9521), .ZN(n9527) );
  INV_X1 U11460 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10698) );
  INV_X1 U11461 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n9522) );
  NAND2_X1 U11462 ( .A1(n9523), .A2(n9522), .ZN(n9524) );
  NAND2_X1 U11463 ( .A1(n9524), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9525) );
  XNOR2_X1 U11464 ( .A(n9525), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10691) );
  MUX2_X1 U11465 ( .A(n10698), .B(P2_REG2_REG_11__SCAN_IN), .S(n10691), .Z(
        n9526) );
  NOR2_X1 U11466 ( .A1(n9527), .A2(n9526), .ZN(n9656) );
  AOI21_X1 U11467 ( .B1(n9527), .B2(n9526), .A(n9656), .ZN(n9539) );
  INV_X1 U11468 ( .A(n15477), .ZN(n11778) );
  INV_X1 U11469 ( .A(n11766), .ZN(n15471) );
  AND2_X1 U11470 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n11275) );
  INV_X1 U11471 ( .A(n10691), .ZN(n9657) );
  NOR2_X1 U11472 ( .A1(n15466), .A2(n9657), .ZN(n9528) );
  AOI211_X1 U11473 ( .C1(n15471), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n11275), 
        .B(n9528), .ZN(n9538) );
  OR2_X1 U11474 ( .A1(n10551), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n9529) );
  NAND2_X1 U11475 ( .A1(n9530), .A2(n9529), .ZN(n9740) );
  INV_X1 U11476 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n16054) );
  MUX2_X1 U11477 ( .A(n16054), .B(P2_REG1_REG_10__SCAN_IN), .S(n10687), .Z(
        n9739) );
  OR2_X1 U11478 ( .A1(n9740), .A2(n9739), .ZN(n9741) );
  NAND2_X1 U11479 ( .A1(n10687), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9535) );
  NAND2_X1 U11480 ( .A1(n9741), .A2(n9535), .ZN(n9533) );
  INV_X1 U11481 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9531) );
  MUX2_X1 U11482 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9531), .S(n10691), .Z(
        n9532) );
  NAND2_X1 U11483 ( .A1(n9533), .A2(n9532), .ZN(n9660) );
  MUX2_X1 U11484 ( .A(n9531), .B(P2_REG1_REG_11__SCAN_IN), .S(n10691), .Z(
        n9534) );
  NAND3_X1 U11485 ( .A1(n9741), .A2(n9535), .A3(n9534), .ZN(n9536) );
  NAND3_X1 U11486 ( .A1(n9660), .A2(n15473), .A3(n9536), .ZN(n9537) );
  OAI211_X1 U11487 ( .C1(n9539), .C2(n11778), .A(n9538), .B(n9537), .ZN(
        P2_U3225) );
  AND2_X2 U11488 ( .A1(n11785), .A2(n7178), .ZN(n9883) );
  NAND2_X2 U11489 ( .A1(n9543), .A2(n9542), .ZN(n15904) );
  INV_X1 U11490 ( .A(P2_B_REG_SCAN_IN), .ZN(n13410) );
  AOI221_X1 U11491 ( .B1(n14602), .B2(n13410), .C1(n9547), .C2(
        P2_B_REG_SCAN_IN), .A(n9546), .ZN(n9550) );
  OR3_X1 U11492 ( .A1(n14596), .A2(P2_D_REG_0__SCAN_IN), .A3(n9550), .ZN(n9549) );
  NAND2_X1 U11493 ( .A1(n14596), .A2(n14602), .ZN(n9548) );
  NOR2_X1 U11494 ( .A1(n14596), .A2(n9550), .ZN(n15176) );
  INV_X1 U11495 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15175) );
  AOI22_X1 U11496 ( .A1(n15176), .A2(n15175), .B1(n14596), .B2(n14599), .ZN(
        n9990) );
  NOR4_X1 U11497 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n9554) );
  NOR4_X1 U11498 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n9553) );
  NOR4_X1 U11499 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n9552) );
  NOR4_X1 U11500 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9551) );
  NAND4_X1 U11501 ( .A1(n9554), .A2(n9553), .A3(n9552), .A4(n9551), .ZN(n9560)
         );
  NOR2_X1 U11502 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n9558) );
  NOR4_X1 U11503 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9557) );
  NOR4_X1 U11504 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n9556) );
  NOR4_X1 U11505 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n9555) );
  NAND4_X1 U11506 ( .A1(n9558), .A2(n9557), .A3(n9556), .A4(n9555), .ZN(n9559)
         );
  OAI21_X1 U11507 ( .B1(n9560), .B2(n9559), .A(n15176), .ZN(n9992) );
  NAND2_X1 U11508 ( .A1(n9990), .A2(n9992), .ZN(n10502) );
  NOR2_X1 U11509 ( .A1(n15408), .A2(n10502), .ZN(n9900) );
  AND2_X1 U11510 ( .A1(n15409), .A2(n9900), .ZN(n9597) );
  INV_X1 U11511 ( .A(n9597), .ZN(n9570) );
  AOI21_X1 U11512 ( .B1(n9566), .B2(n9562), .A(n14582), .ZN(n9565) );
  MUX2_X2 U11513 ( .A(n9565), .B(n9564), .S(n9563), .Z(n13367) );
  INV_X1 U11514 ( .A(n13367), .ZN(n13370) );
  NAND2_X1 U11515 ( .A1(n7190), .A2(n13370), .ZN(n10517) );
  OR2_X1 U11516 ( .A1(n9570), .A2(n10517), .ZN(n9568) );
  NAND2_X1 U11517 ( .A1(n14397), .A2(n7183), .ZN(n9991) );
  INV_X1 U11518 ( .A(n9991), .ZN(n9567) );
  NAND2_X1 U11519 ( .A1(n9595), .A2(n13407), .ZN(n10504) );
  INV_X1 U11520 ( .A(n10504), .ZN(n9569) );
  AOI21_X1 U11521 ( .B1(n9570), .B2(n14430), .A(n9569), .ZN(n9776) );
  INV_X1 U11522 ( .A(n9776), .ZN(n9594) );
  INV_X1 U11523 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10871) );
  NAND2_X1 U11524 ( .A1(n9484), .A2(n9572), .ZN(n9573) );
  NAND2_X1 U11525 ( .A1(n9573), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9574) );
  INV_X1 U11526 ( .A(n9575), .ZN(n14583) );
  NAND2_X2 U11527 ( .A1(n9576), .A2(n14583), .ZN(n9578) );
  NAND2_X1 U11528 ( .A1(n12174), .A2(n9578), .ZN(n9620) );
  OR2_X1 U11529 ( .A1(n9620), .A2(n9577), .ZN(n9584) );
  NAND2_X1 U11530 ( .A1(n9887), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9583) );
  INV_X1 U11531 ( .A(n9578), .ZN(n9580) );
  OR2_X2 U11532 ( .A1(n12174), .A2(n9580), .ZN(n9622) );
  INV_X1 U11533 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9579) );
  NAND2_X1 U11534 ( .A1(n8182), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9581) );
  NAND4_X2 U11535 ( .A1(n9584), .A2(n9583), .A3(n9582), .A4(n9581), .ZN(n14200) );
  INV_X1 U11536 ( .A(n14200), .ZN(n9968) );
  OR2_X1 U11537 ( .A1(n9593), .A2(n9492), .ZN(n14354) );
  INV_X1 U11538 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9585) );
  NAND2_X1 U11539 ( .A1(n8182), .A2(n9585), .ZN(n9591) );
  INV_X1 U11540 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9586) );
  OR2_X1 U11541 ( .A1(n9622), .A2(n9586), .ZN(n9590) );
  NAND2_X1 U11542 ( .A1(n9887), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9588) );
  NAND4_X1 U11543 ( .A1(n9591), .A2(n9590), .A3(n9589), .A4(n9588), .ZN(n14198) );
  INV_X1 U11544 ( .A(n9492), .ZN(n9592) );
  OAI22_X1 U11545 ( .A1(n9968), .A2(n14354), .B1(n9973), .B2(n14356), .ZN(
        n10865) );
  AOI22_X1 U11546 ( .A1(n9594), .A2(P2_REG3_REG_2__SCAN_IN), .B1(n14165), .B2(
        n10865), .ZN(n9635) );
  NOR2_X1 U11547 ( .A1(n15905), .A2(n9595), .ZN(n9596) );
  INV_X1 U11548 ( .A(n10506), .ZN(n13099) );
  NAND2_X1 U11549 ( .A1(n13099), .A2(n13411), .ZN(n13354) );
  OAI21_X1 U11550 ( .B1(n13099), .B2(n13411), .A(n13354), .ZN(n9599) );
  INV_X1 U11551 ( .A(n13099), .ZN(n9600) );
  NAND2_X1 U11552 ( .A1(n8182), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n9606) );
  INV_X1 U11553 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9601) );
  NAND2_X1 U11554 ( .A1(n9887), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9604) );
  OR2_X1 U11555 ( .A1(n9620), .A2(n9602), .ZN(n9603) );
  NAND2_X1 U11556 ( .A1(n14199), .A2(n9772), .ZN(n9608) );
  NAND2_X1 U11557 ( .A1(n9607), .A2(n9608), .ZN(n9875) );
  INV_X1 U11558 ( .A(n9607), .ZN(n9610) );
  INV_X1 U11559 ( .A(n9608), .ZN(n9609) );
  NAND2_X1 U11560 ( .A1(n9610), .A2(n9609), .ZN(n9611) );
  AND2_X1 U11561 ( .A1(n9875), .A2(n9611), .ZN(n9632) );
  NAND2_X1 U11562 ( .A1(n9883), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n9614) );
  XNOR2_X1 U11563 ( .A(n11374), .B(n15864), .ZN(n9617) );
  NAND2_X1 U11564 ( .A1(n14200), .A2(n9772), .ZN(n9616) );
  NAND2_X1 U11565 ( .A1(n9617), .A2(n9616), .ZN(n9630) );
  INV_X1 U11566 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9619) );
  NAND2_X1 U11567 ( .A1(n8182), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n9625) );
  INV_X1 U11568 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9621) );
  OR2_X1 U11569 ( .A1(n9622), .A2(n9621), .ZN(n9624) );
  INV_X1 U11570 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9754) );
  MUX2_X1 U11571 ( .A(n9754), .B(n14604), .S(n11785), .Z(n13101) );
  INV_X1 U11572 ( .A(n13101), .ZN(n10664) );
  AND2_X1 U11573 ( .A1(n9773), .A2(n10664), .ZN(n10660) );
  NAND2_X1 U11574 ( .A1(n10660), .A2(n9772), .ZN(n9628) );
  NAND2_X1 U11575 ( .A1(n14032), .A2(n13101), .ZN(n9627) );
  NAND2_X1 U11576 ( .A1(n9628), .A2(n9627), .ZN(n9711) );
  NAND2_X1 U11577 ( .A1(n9631), .A2(n9632), .ZN(n9876) );
  OAI21_X1 U11578 ( .B1(n9632), .B2(n9631), .A(n9876), .ZN(n9633) );
  NAND2_X1 U11579 ( .A1(n14115), .A2(n9633), .ZN(n9634) );
  OAI211_X1 U11580 ( .C1(n7678), .C2(n14162), .A(n9635), .B(n9634), .ZN(
        P2_U3209) );
  INV_X1 U11581 ( .A(n9636), .ZN(n9637) );
  NAND2_X1 U11582 ( .A1(n9639), .A2(SI_10_), .ZN(n9640) );
  MUX2_X1 U11583 ( .A(n9644), .B(n9646), .S(n7178), .Z(n9641) );
  NAND2_X1 U11584 ( .A1(n9641), .A2(n15208), .ZN(n9760) );
  INV_X1 U11585 ( .A(n9641), .ZN(n9642) );
  NAND2_X1 U11586 ( .A1(n9642), .A2(SI_11_), .ZN(n9643) );
  NAND2_X1 U11587 ( .A1(n9760), .A2(n9643), .ZN(n9761) );
  XNOR2_X1 U11588 ( .A(n7536), .B(n9761), .ZN(n11035) );
  INV_X1 U11589 ( .A(n11035), .ZN(n9645) );
  OAI222_X1 U11590 ( .A1(n14588), .A2(n9644), .B1(n14593), .B2(n9645), .C1(
        P2_U3088), .C2(n9657), .ZN(P2_U3316) );
  OAI222_X1 U11591 ( .A1(n15157), .A2(n9646), .B1(n15167), .B2(n9645), .C1(
        P1_U3086), .C2(n10120), .ZN(P1_U3344) );
  INV_X1 U11592 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n9647) );
  AND4_X1 U11593 ( .A1(n9650), .A2(n9649), .A3(n9648), .A4(n9647), .ZN(n9651)
         );
  NAND2_X1 U11594 ( .A1(n9652), .A2(n9651), .ZN(n9654) );
  NAND2_X1 U11595 ( .A1(n9654), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9653) );
  MUX2_X1 U11596 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9653), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n9655) );
  AOI21_X1 U11597 ( .B1(n9657), .B2(n10698), .A(n9656), .ZN(n10408) );
  XNOR2_X1 U11598 ( .A(n11137), .B(n10408), .ZN(n9658) );
  NOR2_X1 U11599 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n9658), .ZN(n10409) );
  AOI21_X1 U11600 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n9658), .A(n10409), .ZN(
        n9668) );
  NAND2_X1 U11601 ( .A1(n10691), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9659) );
  AND2_X1 U11602 ( .A1(n9660), .A2(n9659), .ZN(n9662) );
  INV_X1 U11603 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n16093) );
  MUX2_X1 U11604 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n16093), .S(n11137), .Z(
        n9661) );
  NAND2_X1 U11605 ( .A1(n9662), .A2(n9661), .ZN(n10402) );
  OAI21_X1 U11606 ( .B1(n9662), .B2(n9661), .A(n10402), .ZN(n9666) );
  INV_X1 U11607 ( .A(n11137), .ZN(n10404) );
  INV_X1 U11608 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n11386) );
  NOR2_X1 U11609 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11386), .ZN(n9663) );
  AOI21_X1 U11610 ( .B1(n15471), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n9663), .ZN(
        n9664) );
  OAI21_X1 U11611 ( .B1(n10404), .B2(n15466), .A(n9664), .ZN(n9665) );
  AOI21_X1 U11612 ( .B1(n9666), .B2(n15473), .A(n9665), .ZN(n9667) );
  OAI21_X1 U11613 ( .B1(n9668), .B2(n11778), .A(n9667), .ZN(P2_U3226) );
  NAND2_X1 U11614 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10017) );
  INV_X1 U11615 ( .A(n10017), .ZN(n9674) );
  MUX2_X1 U11616 ( .A(n9461), .B(P2_REG1_REG_6__SCAN_IN), .S(n10004), .Z(n9669) );
  NAND3_X1 U11617 ( .A1(n15426), .A2(n9670), .A3(n9669), .ZN(n9671) );
  AND3_X1 U11618 ( .A1(n15473), .A2(n9672), .A3(n9671), .ZN(n9673) );
  AOI211_X1 U11619 ( .C1(n15471), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n9674), .B(
        n9673), .ZN(n9680) );
  MUX2_X1 U11620 ( .A(n9982), .B(P2_REG2_REG_6__SCAN_IN), .S(n10004), .Z(n9675) );
  NAND3_X1 U11621 ( .A1(n15423), .A2(n9676), .A3(n9675), .ZN(n9677) );
  NAND3_X1 U11622 ( .A1(n15477), .A2(n9678), .A3(n9677), .ZN(n9679) );
  OAI211_X1 U11623 ( .C1(n15466), .C2(n9681), .A(n9680), .B(n9679), .ZN(
        P2_U3220) );
  NAND2_X1 U11624 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n9915) );
  INV_X1 U11625 ( .A(n9915), .ZN(n9687) );
  MUX2_X1 U11626 ( .A(n9456), .B(P2_REG1_REG_4__SCAN_IN), .S(n9884), .Z(n9682)
         );
  NAND3_X1 U11627 ( .A1(n15415), .A2(n9683), .A3(n9682), .ZN(n9684) );
  AND3_X1 U11628 ( .A1(n15473), .A2(n9685), .A3(n9684), .ZN(n9686) );
  AOI211_X1 U11629 ( .C1(n15471), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n9687), .B(
        n9686), .ZN(n9693) );
  MUX2_X1 U11630 ( .A(n10513), .B(P2_REG2_REG_4__SCAN_IN), .S(n9884), .Z(n9688) );
  NAND3_X1 U11631 ( .A1(n15412), .A2(n9689), .A3(n9688), .ZN(n9690) );
  NAND3_X1 U11632 ( .A1(n15477), .A2(n9691), .A3(n9690), .ZN(n9692) );
  OAI211_X1 U11633 ( .C1(n15466), .C2(n9694), .A(n9693), .B(n9692), .ZN(
        P2_U3218) );
  INV_X1 U11634 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9695) );
  NOR2_X1 U11635 ( .A1(n11766), .A2(n9695), .ZN(n9700) );
  INV_X1 U11636 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n15850) );
  MUX2_X1 U11637 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n9450), .S(n9706), .Z(n9696)
         );
  OAI21_X1 U11638 ( .B1(n15850), .B2(n9754), .A(n9696), .ZN(n9697) );
  AND3_X1 U11639 ( .A1(n15473), .A2(n9698), .A3(n9697), .ZN(n9699) );
  AOI211_X1 U11640 ( .C1(P2_REG3_REG_1__SCAN_IN), .C2(P2_U3088), .A(n9700), 
        .B(n9699), .ZN(n9705) );
  MUX2_X1 U11641 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n9577), .S(n9706), .Z(n9701)
         );
  OAI21_X1 U11642 ( .B1(n9619), .B2(n9754), .A(n9701), .ZN(n9702) );
  NAND3_X1 U11643 ( .A1(n15477), .A2(n9703), .A3(n9702), .ZN(n9704) );
  OAI211_X1 U11644 ( .C1(n15466), .C2(n9706), .A(n9705), .B(n9704), .ZN(
        P2_U3215) );
  INV_X1 U11645 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9707) );
  INV_X1 U11646 ( .A(n14165), .ZN(n14144) );
  INV_X1 U11647 ( .A(n14356), .ZN(n14139) );
  AOI22_X1 U11648 ( .A1(n14137), .A2(n9773), .B1(n14199), .B2(n14139), .ZN(
        n10662) );
  OAI22_X1 U11649 ( .A1(n9776), .A2(n9707), .B1(n14144), .B2(n10662), .ZN(
        n9714) );
  INV_X1 U11650 ( .A(n9708), .ZN(n9709) );
  AOI21_X1 U11651 ( .B1(n9711), .B2(n9710), .A(n9709), .ZN(n9712) );
  OAI22_X1 U11652 ( .A1(n14168), .A2(n9712), .B1(n14162), .B2(n15864), .ZN(
        n9713) );
  OR2_X1 U11653 ( .A1(n9714), .A2(n9713), .ZN(P2_U3194) );
  OAI211_X1 U11654 ( .C1(n9717), .C2(n9716), .A(n15473), .B(n9715), .ZN(n9721)
         );
  OAI211_X1 U11655 ( .C1(n9719), .C2(n9718), .A(n15477), .B(n9728), .ZN(n9720)
         );
  NAND2_X1 U11656 ( .A1(n9721), .A2(n9720), .ZN(n9723) );
  NAND2_X1 U11657 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n10356) );
  INV_X1 U11658 ( .A(n10356), .ZN(n9722) );
  AOI211_X1 U11659 ( .C1(n15471), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n9723), .B(
        n9722), .ZN(n9724) );
  OAI21_X1 U11660 ( .B1(n9725), .B2(n15466), .A(n9724), .ZN(P2_U3221) );
  MUX2_X1 U11661 ( .A(n10347), .B(P2_REG2_REG_8__SCAN_IN), .S(n10447), .Z(
        n9726) );
  NAND3_X1 U11662 ( .A1(n9728), .A2(n9727), .A3(n9726), .ZN(n9729) );
  NAND3_X1 U11663 ( .A1(n15477), .A2(n9730), .A3(n9729), .ZN(n9737) );
  NAND2_X1 U11664 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n10462) );
  OAI211_X1 U11665 ( .C1(n9733), .C2(n9732), .A(n15473), .B(n9731), .ZN(n9734)
         );
  NAND2_X1 U11666 ( .A1(n10462), .A2(n9734), .ZN(n9735) );
  AOI21_X1 U11667 ( .B1(n15471), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n9735), .ZN(
        n9736) );
  OAI211_X1 U11668 ( .C1(n15466), .C2(n9738), .A(n9737), .B(n9736), .ZN(
        P2_U3222) );
  AOI21_X1 U11669 ( .B1(n9740), .B2(n9739), .A(n14230), .ZN(n9742) );
  NAND2_X1 U11670 ( .A1(n9742), .A2(n9741), .ZN(n9750) );
  NAND2_X1 U11671 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n10853)
         );
  AOI21_X1 U11672 ( .B1(n9744), .B2(n9743), .A(n11778), .ZN(n9746) );
  NAND2_X1 U11673 ( .A1(n9746), .A2(n9745), .ZN(n9747) );
  NAND2_X1 U11674 ( .A1(n10853), .A2(n9747), .ZN(n9748) );
  AOI21_X1 U11675 ( .B1(n15471), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n9748), .ZN(
        n9749) );
  OAI211_X1 U11676 ( .C1(n15466), .C2(n9751), .A(n9750), .B(n9749), .ZN(
        P2_U3224) );
  INV_X1 U11677 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9759) );
  NAND2_X1 U11678 ( .A1(n15473), .A2(n15850), .ZN(n9753) );
  NAND2_X1 U11679 ( .A1(n15477), .A2(n9619), .ZN(n9752) );
  AND3_X1 U11680 ( .A1(n9753), .A2(n9752), .A3(n15466), .ZN(n9756) );
  AOI22_X1 U11681 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n15473), .B1(n15477), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n9755) );
  MUX2_X1 U11682 ( .A(n9756), .B(n9755), .S(n9754), .Z(n9758) );
  NAND2_X1 U11683 ( .A1(n15471), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n9757) );
  OAI211_X1 U11684 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n9759), .A(n9758), .B(
        n9757), .ZN(P2_U3214) );
  MUX2_X1 U11685 ( .A(n9851), .B(n9768), .S(n7178), .Z(n9763) );
  NAND2_X1 U11686 ( .A1(n9763), .A2(n15319), .ZN(n10023) );
  INV_X1 U11687 ( .A(n9763), .ZN(n9764) );
  NAND2_X1 U11688 ( .A1(n9764), .A2(SI_12_), .ZN(n9765) );
  XNOR2_X1 U11689 ( .A(n10022), .B(n10021), .ZN(n11229) );
  INV_X1 U11690 ( .A(n11229), .ZN(n9850) );
  NAND2_X1 U11691 ( .A1(n10025), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9767) );
  XNOR2_X1 U11692 ( .A(n9767), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11230) );
  INV_X1 U11693 ( .A(n11230), .ZN(n10204) );
  OAI222_X1 U11694 ( .A1(n15167), .A2(n9850), .B1(n10204), .B2(P1_U3086), .C1(
        n9768), .C2(n15157), .ZN(P1_U3343) );
  NOR2_X1 U11695 ( .A1(n13550), .A2(P3_U3151), .ZN(n10397) );
  INV_X1 U11696 ( .A(n10319), .ZN(n10104) );
  NAND2_X1 U11697 ( .A1(n13578), .A2(n10104), .ZN(n12643) );
  NAND2_X1 U11698 ( .A1(n10420), .A2(n12643), .ZN(n12602) );
  OAI22_X1 U11699 ( .A1(n13519), .A2(n9769), .B1(n10104), .B2(n13554), .ZN(
        n9770) );
  AOI21_X1 U11700 ( .B1(n13527), .B2(n12602), .A(n9770), .ZN(n9771) );
  OAI21_X1 U11701 ( .B1(n10397), .B2(n15658), .A(n9771), .ZN(P3_U3172) );
  NAND2_X1 U11702 ( .A1(n14115), .A2(n14416), .ZN(n14152) );
  INV_X1 U11703 ( .A(n14152), .ZN(n14063) );
  AOI21_X1 U11704 ( .B1(n10664), .B2(n14397), .A(n9774), .ZN(n9775) );
  NAND2_X1 U11705 ( .A1(n14200), .A2(n14139), .ZN(n10653) );
  OAI22_X1 U11706 ( .A1(n9775), .A2(n14168), .B1(n14144), .B2(n10653), .ZN(
        n9778) );
  OAI22_X1 U11707 ( .A1(n9776), .A2(n9759), .B1(n14162), .B2(n13101), .ZN(
        n9777) );
  AOI211_X1 U11708 ( .C1(n14063), .C2(n13106), .A(n9778), .B(n9777), .ZN(n9779) );
  INV_X1 U11709 ( .A(n9779), .ZN(P2_U3204) );
  OR2_X1 U11710 ( .A1(n12762), .A2(n9780), .ZN(n9781) );
  AND2_X1 U11711 ( .A1(n9782), .A2(n9781), .ZN(n9785) );
  INV_X1 U11712 ( .A(n9783), .ZN(n9784) );
  NAND2_X1 U11713 ( .A1(n9784), .A2(n12791), .ZN(n9786) );
  AND2_X1 U11714 ( .A1(n9785), .A2(n9786), .ZN(n9812) );
  INV_X1 U11715 ( .A(n15817), .ZN(n15773) );
  INV_X1 U11716 ( .A(n10151), .ZN(n9840) );
  INV_X1 U11717 ( .A(n9785), .ZN(n9787) );
  NOR2_X1 U11718 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15365), .ZN(n10990) );
  MUX2_X1 U11719 ( .A(n9825), .B(P3_REG1_REG_2__SCAN_IN), .S(n9827), .Z(n9941)
         );
  NOR2_X1 U11720 ( .A1(n9823), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9788) );
  NAND2_X1 U11721 ( .A1(n8386), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9789) );
  OAI21_X1 U11722 ( .B1(n9932), .B2(n9788), .A(n9789), .ZN(n9921) );
  OR2_X1 U11723 ( .A1(n9921), .A2(n9818), .ZN(n9923) );
  NAND2_X1 U11724 ( .A1(n9923), .A2(n9789), .ZN(n9940) );
  NAND2_X1 U11725 ( .A1(n9941), .A2(n9940), .ZN(n9939) );
  NAND2_X1 U11726 ( .A1(n9956), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9790) );
  INV_X1 U11727 ( .A(n9834), .ZN(n9872) );
  MUX2_X1 U11728 ( .A(n10147), .B(P3_REG1_REG_4__SCAN_IN), .S(n10151), .Z(
        n9793) );
  NAND2_X1 U11729 ( .A1(n9792), .A2(n9793), .ZN(n10149) );
  INV_X1 U11730 ( .A(n9793), .ZN(n9795) );
  NAND3_X1 U11731 ( .A1(n9856), .A2(n9795), .A3(n9794), .ZN(n9796) );
  AOI21_X1 U11732 ( .B1(n10149), .B2(n9796), .A(n15822), .ZN(n9797) );
  AOI211_X1 U11733 ( .C1(n15771), .C2(P3_ADDR_REG_4__SCAN_IN), .A(n10990), .B(
        n9797), .ZN(n9816) );
  NAND2_X1 U11734 ( .A1(n8386), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9802) );
  NAND2_X1 U11735 ( .A1(n9932), .A2(n9802), .ZN(n9801) );
  INV_X1 U11736 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n9798) );
  NAND2_X1 U11737 ( .A1(n9798), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9799) );
  OR2_X1 U11738 ( .A1(n9799), .A2(n8386), .ZN(n9800) );
  NAND2_X1 U11739 ( .A1(n9924), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n9803) );
  NAND2_X1 U11740 ( .A1(n9827), .A2(n9826), .ZN(n9937) );
  NAND2_X1 U11741 ( .A1(n9938), .A2(n9937), .ZN(n9804) );
  NAND2_X1 U11742 ( .A1(n9956), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9934) );
  MUX2_X1 U11743 ( .A(n11028), .B(P3_REG2_REG_4__SCAN_IN), .S(n10151), .Z(
        n9808) );
  NAND2_X1 U11744 ( .A1(n9805), .A2(n9808), .ZN(n10153) );
  INV_X1 U11745 ( .A(n10153), .ZN(n9814) );
  INV_X1 U11746 ( .A(n9852), .ZN(n9809) );
  INV_X1 U11747 ( .A(n9806), .ZN(n9807) );
  NOR3_X1 U11748 ( .A1(n9809), .A2(n9808), .A3(n9807), .ZN(n9813) );
  INV_X1 U11749 ( .A(n9810), .ZN(n9811) );
  INV_X1 U11750 ( .A(n15825), .ZN(n13625) );
  OAI21_X1 U11751 ( .B1(n9814), .B2(n9813), .A(n13625), .ZN(n9815) );
  OAI211_X1 U11752 ( .C1(n15773), .C2(n9840), .A(n9816), .B(n9815), .ZN(n9849)
         );
  MUX2_X1 U11753 ( .A(n10527), .B(n9818), .S(n8767), .Z(n9820) );
  INV_X1 U11754 ( .A(n9932), .ZN(n9819) );
  NAND2_X1 U11755 ( .A1(n9820), .A2(n9819), .ZN(n9948) );
  INV_X1 U11756 ( .A(n9820), .ZN(n9821) );
  NAND2_X1 U11757 ( .A1(n9821), .A2(n9932), .ZN(n9822) );
  AND2_X1 U11758 ( .A1(n9948), .A2(n9822), .ZN(n9920) );
  MUX2_X1 U11759 ( .A(n9824), .B(n9823), .S(n13664), .Z(n15652) );
  AND2_X1 U11760 ( .A1(n15652), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15655) );
  NAND2_X1 U11761 ( .A1(n9947), .A2(n9948), .ZN(n9831) );
  MUX2_X1 U11762 ( .A(n9826), .B(n9825), .S(n13664), .Z(n9828) );
  NAND2_X1 U11763 ( .A1(n9828), .A2(n9827), .ZN(n9864) );
  INV_X1 U11764 ( .A(n9828), .ZN(n9829) );
  NAND2_X1 U11765 ( .A1(n9829), .A2(n9956), .ZN(n9830) );
  AND2_X1 U11766 ( .A1(n9864), .A2(n9830), .ZN(n9949) );
  NAND2_X1 U11767 ( .A1(n9831), .A2(n9949), .ZN(n9863) );
  NAND2_X1 U11768 ( .A1(n9863), .A2(n9864), .ZN(n9838) );
  MUX2_X1 U11769 ( .A(n9833), .B(n9832), .S(n13664), .Z(n9835) );
  NAND2_X1 U11770 ( .A1(n9835), .A2(n9834), .ZN(n9846) );
  INV_X1 U11771 ( .A(n9835), .ZN(n9836) );
  NAND2_X1 U11772 ( .A1(n9836), .A2(n9872), .ZN(n9837) );
  AND2_X1 U11773 ( .A1(n9846), .A2(n9837), .ZN(n9865) );
  NAND2_X1 U11774 ( .A1(n9867), .A2(n9846), .ZN(n9843) );
  MUX2_X1 U11775 ( .A(n11028), .B(n10147), .S(n13664), .Z(n9839) );
  NAND2_X1 U11776 ( .A1(n9839), .A2(n10151), .ZN(n10142) );
  INV_X1 U11777 ( .A(n9839), .ZN(n9841) );
  NAND2_X1 U11778 ( .A1(n9841), .A2(n9840), .ZN(n9842) );
  AND2_X1 U11779 ( .A1(n10142), .A2(n9842), .ZN(n9844) );
  NAND2_X1 U11780 ( .A1(n9843), .A2(n9844), .ZN(n10143) );
  INV_X1 U11781 ( .A(n9844), .ZN(n9845) );
  NAND3_X1 U11782 ( .A1(n9867), .A2(n9846), .A3(n9845), .ZN(n9847) );
  NAND2_X1 U11783 ( .A1(P3_U3897), .A2(n12193), .ZN(n15811) );
  AOI21_X1 U11784 ( .B1(n10143), .B2(n9847), .A(n15811), .ZN(n9848) );
  OR2_X1 U11785 ( .A1(n9849), .A2(n9848), .ZN(P3_U3186) );
  OAI222_X1 U11786 ( .A1(n14588), .A2(n9851), .B1(n14593), .B2(n9850), .C1(
        n10404), .C2(P2_U3088), .ZN(P2_U3315) );
  OAI21_X1 U11787 ( .B1(n9853), .B2(P3_REG2_REG_3__SCAN_IN), .A(n9852), .ZN(
        n9862) );
  NAND2_X1 U11788 ( .A1(n9854), .A2(n9832), .ZN(n9855) );
  AOI21_X1 U11789 ( .B1(n9856), .B2(n9855), .A(n15822), .ZN(n9861) );
  INV_X1 U11790 ( .A(n15771), .ZN(n15808) );
  INV_X1 U11791 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n9859) );
  NOR2_X1 U11792 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9857), .ZN(n10638) );
  INV_X1 U11793 ( .A(n10638), .ZN(n9858) );
  OAI21_X1 U11794 ( .B1(n15808), .B2(n9859), .A(n9858), .ZN(n9860) );
  AOI211_X1 U11795 ( .C1(n13625), .C2(n9862), .A(n9861), .B(n9860), .ZN(n9871)
         );
  INV_X1 U11796 ( .A(n9863), .ZN(n9952) );
  INV_X1 U11797 ( .A(n9864), .ZN(n9866) );
  NOR3_X1 U11798 ( .A1(n9952), .A2(n9866), .A3(n9865), .ZN(n9869) );
  INV_X1 U11799 ( .A(n9867), .ZN(n9868) );
  OAI21_X1 U11800 ( .B1(n9869), .B2(n9868), .A(n15775), .ZN(n9870) );
  OAI211_X1 U11801 ( .C1(n15773), .C2(n9872), .A(n9871), .B(n9870), .ZN(
        P3_U3185) );
  INV_X1 U11802 ( .A(n9873), .ZN(n9874) );
  OAI222_X1 U11803 ( .A1(P3_U3151), .A2(n13639), .B1(n13083), .B2(n15207), 
        .C1(n13082), .C2(n9874), .ZN(P3_U3279) );
  AOI22_X1 U11804 ( .A1(n9883), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n12234), 
        .B2(n9878), .ZN(n9879) );
  XNOR2_X1 U11805 ( .A(n13127), .B(n14032), .ZN(n9882) );
  NAND2_X1 U11806 ( .A1(n14198), .A2(n9772), .ZN(n9881) );
  XNOR2_X1 U11807 ( .A(n9882), .B(n9881), .ZN(n10030) );
  INV_X2 U11808 ( .A(n9957), .ZN(n13330) );
  AOI22_X1 U11809 ( .A1(n13330), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n12234), 
        .B2(n9884), .ZN(n9885) );
  XNOR2_X1 U11810 ( .A(n13145), .B(n14032), .ZN(n9892) );
  NAND2_X1 U11811 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n9907) );
  OAI21_X1 U11812 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n9907), .ZN(n10519) );
  OR2_X1 U11813 ( .A1(n12314), .A2(n10519), .ZN(n9891) );
  NAND2_X1 U11814 ( .A1(n13321), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9890) );
  NAND2_X1 U11815 ( .A1(n12345), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9889) );
  NAND2_X1 U11816 ( .A1(n12336), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9888) );
  NAND4_X2 U11817 ( .A1(n9891), .A2(n9890), .A3(n9889), .A4(n9888), .ZN(n14197) );
  NAND2_X1 U11818 ( .A1(n14197), .A2(n9772), .ZN(n9893) );
  NAND2_X1 U11819 ( .A1(n9892), .A2(n9893), .ZN(n9996) );
  INV_X1 U11820 ( .A(n9892), .ZN(n9895) );
  INV_X1 U11821 ( .A(n9893), .ZN(n9894) );
  NAND2_X1 U11822 ( .A1(n9895), .A2(n9894), .ZN(n9896) );
  NAND2_X1 U11823 ( .A1(n9996), .A2(n9896), .ZN(n9898) );
  INV_X1 U11824 ( .A(n9997), .ZN(n9897) );
  AOI21_X1 U11825 ( .B1(n9899), .B2(n9898), .A(n9897), .ZN(n9919) );
  INV_X1 U11826 ( .A(n14162), .ZN(n14150) );
  INV_X1 U11827 ( .A(n9900), .ZN(n9901) );
  NAND2_X1 U11828 ( .A1(n9901), .A2(n9991), .ZN(n9903) );
  NAND3_X1 U11829 ( .A1(n9903), .A2(n9902), .A3(n10504), .ZN(n9904) );
  NAND2_X1 U11830 ( .A1(n12345), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9914) );
  INV_X1 U11831 ( .A(n9907), .ZN(n9905) );
  NAND2_X1 U11832 ( .A1(n9905), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9980) );
  INV_X1 U11833 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9906) );
  NAND2_X1 U11834 ( .A1(n9907), .A2(n9906), .ZN(n9908) );
  AND2_X1 U11835 ( .A1(n9980), .A2(n9908), .ZN(n10946) );
  NAND2_X1 U11836 ( .A1(n12342), .A2(n10946), .ZN(n9913) );
  OR2_X1 U11837 ( .A1(n12239), .A2(n9909), .ZN(n9912) );
  INV_X1 U11838 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9910) );
  OR2_X1 U11839 ( .A1(n9622), .A2(n9910), .ZN(n9911) );
  NAND4_X1 U11840 ( .A1(n9914), .A2(n9913), .A3(n9912), .A4(n9911), .ZN(n14196) );
  INV_X1 U11841 ( .A(n14196), .ZN(n10114) );
  OAI22_X1 U11842 ( .A1(n9973), .A2(n14354), .B1(n10114), .B2(n14356), .ZN(
        n10511) );
  NAND2_X1 U11843 ( .A1(n14165), .A2(n10511), .ZN(n9916) );
  OAI211_X1 U11844 ( .C1(n14161), .C2(n10519), .A(n9916), .B(n9915), .ZN(n9917) );
  AOI21_X1 U11845 ( .B1(n13145), .B2(n14150), .A(n9917), .ZN(n9918) );
  OAI21_X1 U11846 ( .B1(n9919), .B2(n14168), .A(n9918), .ZN(P2_U3202) );
  OAI21_X1 U11847 ( .B1(n9920), .B2(n15655), .A(n9947), .ZN(n9930) );
  NAND2_X1 U11848 ( .A1(n9921), .A2(n9818), .ZN(n9922) );
  AND2_X1 U11849 ( .A1(n9923), .A2(n9922), .ZN(n9928) );
  AOI22_X1 U11850 ( .A1(n15771), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n9927) );
  XNOR2_X1 U11851 ( .A(n9924), .B(P3_REG2_REG_1__SCAN_IN), .ZN(n9925) );
  NAND2_X1 U11852 ( .A1(n13625), .A2(n9925), .ZN(n9926) );
  OAI211_X1 U11853 ( .C1(n9928), .C2(n15822), .A(n9927), .B(n9926), .ZN(n9929)
         );
  AOI21_X1 U11854 ( .B1(n15775), .B2(n9930), .A(n9929), .ZN(n9931) );
  OAI21_X1 U11855 ( .B1(n9932), .B2(n15773), .A(n9931), .ZN(P3_U3183) );
  INV_X1 U11856 ( .A(n9938), .ZN(n9935) );
  OAI21_X1 U11857 ( .B1(n9935), .B2(n9934), .A(n9933), .ZN(n9936) );
  OAI21_X1 U11858 ( .B1(n9938), .B2(n9937), .A(n9936), .ZN(n9946) );
  INV_X1 U11859 ( .A(n15822), .ZN(n10162) );
  OAI21_X1 U11860 ( .B1(n9941), .B2(n9940), .A(n9939), .ZN(n9942) );
  AND2_X1 U11861 ( .A1(n10162), .A2(n9942), .ZN(n9945) );
  INV_X1 U11862 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n9943) );
  OAI22_X1 U11863 ( .A1(n15808), .A2(n9943), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15891), .ZN(n9944) );
  AOI211_X1 U11864 ( .C1(n13625), .C2(n9946), .A(n9945), .B(n9944), .ZN(n9955)
         );
  INV_X1 U11865 ( .A(n9947), .ZN(n9951) );
  INV_X1 U11866 ( .A(n9948), .ZN(n9950) );
  NOR3_X1 U11867 ( .A1(n9951), .A2(n9950), .A3(n9949), .ZN(n9953) );
  OAI21_X1 U11868 ( .B1(n9953), .B2(n9952), .A(n15775), .ZN(n9954) );
  OAI211_X1 U11869 ( .C1(n15773), .C2(n9956), .A(n9955), .B(n9954), .ZN(
        P3_U3184) );
  AOI22_X1 U11870 ( .A1(n13330), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n12234), 
        .B2(n9958), .ZN(n9959) );
  XNOR2_X1 U11871 ( .A(n13153), .B(n14196), .ZN(n13373) );
  XNOR2_X1 U11872 ( .A(n15904), .B(n14199), .ZN(n13369) );
  INV_X1 U11873 ( .A(n13369), .ZN(n10867) );
  INV_X1 U11874 ( .A(n14199), .ZN(n10032) );
  NAND2_X1 U11875 ( .A1(n7678), .A2(n10032), .ZN(n9961) );
  NAND2_X1 U11876 ( .A1(n9962), .A2(n9961), .ZN(n10833) );
  NAND2_X1 U11877 ( .A1(n10833), .A2(n13371), .ZN(n9964) );
  OR2_X1 U11878 ( .A1(n13127), .A2(n14198), .ZN(n9963) );
  NAND2_X1 U11879 ( .A1(n9964), .A2(n9963), .ZN(n10509) );
  XNOR2_X1 U11880 ( .A(n13145), .B(n14197), .ZN(n13374) );
  NAND2_X1 U11881 ( .A1(n10509), .A2(n7444), .ZN(n9966) );
  OR2_X1 U11882 ( .A1(n13145), .A2(n14197), .ZN(n9965) );
  XOR2_X1 U11883 ( .A(n13373), .B(n10108), .Z(n10952) );
  AND2_X1 U11884 ( .A1(n13367), .A2(n7183), .ZN(n13326) );
  NAND2_X1 U11885 ( .A1(n13326), .A2(n13411), .ZN(n16106) );
  INV_X1 U11886 ( .A(n13153), .ZN(n9967) );
  INV_X1 U11887 ( .A(n13127), .ZN(n15944) );
  NOR2_X2 U11888 ( .A1(n10836), .A2(n13145), .ZN(n10514) );
  OAI211_X1 U11889 ( .C1(n9967), .C2(n10514), .A(n14397), .B(n10110), .ZN(
        n10948) );
  OAI21_X1 U11890 ( .B1(n9967), .B2(n16136), .A(n10948), .ZN(n9989) );
  NAND2_X1 U11891 ( .A1(n9968), .A2(n13109), .ZN(n9969) );
  NAND2_X1 U11892 ( .A1(n9970), .A2(n9969), .ZN(n10864) );
  NAND2_X1 U11893 ( .A1(n10864), .A2(n13369), .ZN(n9972) );
  NAND2_X1 U11894 ( .A1(n10032), .A2(n15904), .ZN(n9971) );
  INV_X1 U11895 ( .A(n13371), .ZN(n10829) );
  NAND2_X1 U11896 ( .A1(n10830), .A2(n10829), .ZN(n9975) );
  NAND2_X1 U11897 ( .A1(n13127), .A2(n9973), .ZN(n9974) );
  INV_X1 U11898 ( .A(n14197), .ZN(n10033) );
  NAND2_X1 U11899 ( .A1(n13145), .A2(n10033), .ZN(n9976) );
  XOR2_X1 U11900 ( .A(n13373), .B(n10113), .Z(n9988) );
  OR2_X1 U11901 ( .A1(n13411), .A2(n14226), .ZN(n9977) );
  NAND2_X1 U11902 ( .A1(n13370), .A2(n7182), .ZN(n13358) );
  NAND2_X1 U11903 ( .A1(n12345), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9987) );
  INV_X1 U11904 ( .A(n9980), .ZN(n9978) );
  NAND2_X1 U11905 ( .A1(n9978), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10008) );
  INV_X1 U11906 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9979) );
  NAND2_X1 U11907 ( .A1(n9980), .A2(n9979), .ZN(n9981) );
  AND2_X1 U11908 ( .A1(n10008), .A2(n9981), .ZN(n10955) );
  NAND2_X1 U11909 ( .A1(n12342), .A2(n10955), .ZN(n9986) );
  OR2_X1 U11910 ( .A1(n12239), .A2(n9982), .ZN(n9985) );
  INV_X1 U11911 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9983) );
  OR2_X1 U11912 ( .A1(n13325), .A2(n9983), .ZN(n9984) );
  NAND4_X1 U11913 ( .A1(n9987), .A2(n9986), .A3(n9985), .A4(n9984), .ZN(n14195) );
  AOI22_X1 U11914 ( .A1(n14137), .A2(n14197), .B1(n14195), .B2(n14139), .ZN(
        n10099) );
  OAI21_X1 U11915 ( .B1(n9988), .B2(n14413), .A(n10099), .ZN(n10949) );
  AOI211_X1 U11916 ( .C1(n10952), .C2(n16140), .A(n9989), .B(n10949), .ZN(
        n10137) );
  OR2_X1 U11917 ( .A1(n9990), .A2(n15406), .ZN(n15173) );
  NAND3_X1 U11918 ( .A1(n9992), .A2(n9991), .A3(n10504), .ZN(n9993) );
  INV_X1 U11919 ( .A(n15408), .ZN(n9994) );
  NAND2_X1 U11920 ( .A1(n16141), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9995) );
  OAI21_X1 U11921 ( .B1(n10137), .B2(n16141), .A(n9995), .ZN(P2_U3504) );
  NAND2_X1 U11922 ( .A1(n9998), .A2(n9999), .ZN(n10003) );
  INV_X1 U11923 ( .A(n9998), .ZN(n10001) );
  INV_X1 U11924 ( .A(n9999), .ZN(n10000) );
  NAND2_X1 U11925 ( .A1(n10001), .A2(n10000), .ZN(n10002) );
  AOI22_X1 U11926 ( .A1(n13330), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n12234), 
        .B2(n10004), .ZN(n10005) );
  XNOR2_X1 U11927 ( .A(n13161), .B(n14032), .ZN(n10330) );
  NAND2_X1 U11928 ( .A1(n14195), .A2(n14416), .ZN(n10331) );
  XNOR2_X1 U11929 ( .A(n10330), .B(n10331), .ZN(n10329) );
  XNOR2_X1 U11930 ( .A(n10328), .B(n10329), .ZN(n10020) );
  NAND2_X1 U11931 ( .A1(n13322), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10015) );
  NAND2_X1 U11932 ( .A1(n10008), .A2(n10007), .ZN(n10009) );
  AND2_X1 U11933 ( .A1(n10345), .A2(n10009), .ZN(n10355) );
  NAND2_X1 U11934 ( .A1(n12342), .A2(n10355), .ZN(n10014) );
  OR2_X1 U11935 ( .A1(n12239), .A2(n10010), .ZN(n10013) );
  INV_X1 U11936 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10011) );
  OR2_X1 U11937 ( .A1(n13325), .A2(n10011), .ZN(n10012) );
  NAND4_X1 U11938 ( .A1(n10015), .A2(n10014), .A3(n10013), .A4(n10012), .ZN(
        n14194) );
  AOI22_X1 U11939 ( .A1(n14137), .A2(n14196), .B1(n14194), .B2(n14139), .ZN(
        n10116) );
  INV_X1 U11940 ( .A(n14161), .ZN(n14141) );
  NAND2_X1 U11941 ( .A1(n14141), .A2(n10955), .ZN(n10016) );
  OAI211_X1 U11942 ( .C1(n14144), .C2(n10116), .A(n10017), .B(n10016), .ZN(
        n10018) );
  AOI21_X1 U11943 ( .B1(n13161), .B2(n14150), .A(n10018), .ZN(n10019) );
  OAI21_X1 U11944 ( .B1(n10020), .B2(n14168), .A(n10019), .ZN(P2_U3211) );
  MUX2_X1 U11945 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7178), .Z(n10297) );
  XNOR2_X1 U11946 ( .A(n10297), .B(n15311), .ZN(n10294) );
  INV_X1 U11947 ( .A(n11412), .ZN(n10092) );
  OAI21_X1 U11948 ( .B1(n10025), .B2(P1_IR_REG_12__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10027) );
  INV_X1 U11949 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10026) );
  NAND2_X1 U11950 ( .A1(n10027), .A2(n10026), .ZN(n10302) );
  OR2_X1 U11951 ( .A1(n10027), .A2(n10026), .ZN(n10028) );
  INV_X1 U11952 ( .A(n11413), .ZN(n10612) );
  OAI222_X1 U11953 ( .A1(n15167), .A2(n10092), .B1(n10612), .B2(P1_U3086), 
        .C1(n10029), .C2(n15157), .ZN(P1_U3342) );
  XNOR2_X1 U11954 ( .A(n10031), .B(n10030), .ZN(n10038) );
  OAI22_X1 U11955 ( .A1(n10033), .A2(n14356), .B1(n10032), .B2(n14354), .ZN(
        n10831) );
  INV_X1 U11956 ( .A(n10831), .ZN(n10035) );
  AOI22_X1 U11957 ( .A1(n14141), .A2(n9585), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        P2_U3088), .ZN(n10034) );
  OAI21_X1 U11958 ( .B1(n14144), .B2(n10035), .A(n10034), .ZN(n10036) );
  AOI21_X1 U11959 ( .B1(n13127), .B2(n14150), .A(n10036), .ZN(n10037) );
  OAI21_X1 U11960 ( .B1(n10038), .B2(n14168), .A(n10037), .ZN(P2_U3190) );
  OAI222_X1 U11961 ( .A1(P3_U3151), .A2(n13641), .B1(n13083), .B2(n15205), 
        .C1(n13082), .C2(n10039), .ZN(P3_U3278) );
  NAND2_X1 U11962 ( .A1(n9877), .A2(n10051), .ZN(n10042) );
  AOI22_X1 U11963 ( .A1(n10053), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n12008), 
        .B2(n14788), .ZN(n10041) );
  NAND2_X1 U11964 ( .A1(n10042), .A2(n10041), .ZN(n15918) );
  INV_X1 U11965 ( .A(n15918), .ZN(n10273) );
  INV_X1 U11966 ( .A(n14750), .ZN(n10275) );
  OAI22_X1 U11967 ( .A1(n10273), .A2(n12525), .B1(n10275), .B2(n12524), .ZN(
        n10050) );
  XNOR2_X1 U11968 ( .A(n10043), .B(n12526), .ZN(n10049) );
  INV_X1 U11969 ( .A(n10044), .ZN(n10048) );
  XNOR2_X1 U11970 ( .A(n10049), .B(n10050), .ZN(n15924) );
  NAND2_X1 U11971 ( .A1(n10052), .A2(n12089), .ZN(n10055) );
  AOI22_X1 U11972 ( .A1(n13011), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n12008), 
        .B2(n14808), .ZN(n10054) );
  NAND2_X1 U11973 ( .A1(n10055), .A2(n10054), .ZN(n15949) );
  NAND2_X1 U11974 ( .A1(n9339), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10061) );
  INV_X1 U11975 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n10056) );
  NAND2_X1 U11976 ( .A1(n10623), .A2(n10056), .ZN(n10057) );
  NAND2_X1 U11977 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n10068) );
  AND2_X1 U11978 ( .A1(n10057), .A2(n10068), .ZN(n10543) );
  NAND2_X1 U11979 ( .A1(n12095), .A2(n10543), .ZN(n10060) );
  NAND2_X1 U11980 ( .A1(n12988), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10059) );
  NAND2_X1 U11981 ( .A1(n12014), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n10058) );
  NAND4_X1 U11982 ( .A1(n10061), .A2(n10060), .A3(n10059), .A4(n10058), .ZN(
        n14749) );
  AOI22_X1 U11983 ( .A1(n15949), .A2(n12519), .B1(n12518), .B2(n14749), .ZN(
        n10062) );
  NAND2_X1 U11984 ( .A1(n10063), .A2(n10062), .ZN(n10220) );
  INV_X1 U11985 ( .A(n10220), .ZN(n10064) );
  NOR2_X1 U11986 ( .A1(n10218), .A2(n10064), .ZN(n10066) );
  AOI22_X1 U11987 ( .A1(n15949), .A2(n7181), .B1(n12519), .B2(n14749), .ZN(
        n10065) );
  XOR2_X1 U11988 ( .A(n12526), .B(n10065), .Z(n10219) );
  XNOR2_X1 U11989 ( .A(n10066), .B(n10219), .ZN(n10085) );
  NAND2_X1 U11990 ( .A1(n12987), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n10073) );
  NOR2_X1 U11991 ( .A1(n10068), .A2(n10067), .ZN(n10235) );
  INV_X1 U11992 ( .A(n10235), .ZN(n10237) );
  NAND2_X1 U11993 ( .A1(n10068), .A2(n10067), .ZN(n10069) );
  AND2_X1 U11994 ( .A1(n10237), .A2(n10069), .ZN(n10680) );
  NAND2_X1 U11995 ( .A1(n12095), .A2(n10680), .ZN(n10072) );
  NAND2_X1 U11996 ( .A1(n12988), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10071) );
  NAND2_X1 U11997 ( .A1(n12014), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n10070) );
  NAND4_X1 U11998 ( .A1(n10073), .A2(n10072), .A3(n10071), .A4(n10070), .ZN(
        n14748) );
  NAND2_X1 U11999 ( .A1(n14748), .A2(n14980), .ZN(n10075) );
  NAND2_X1 U12000 ( .A1(n14750), .A2(n14978), .ZN(n10074) );
  AND2_X1 U12001 ( .A1(n10075), .A2(n10074), .ZN(n15951) );
  AND3_X1 U12002 ( .A1(n10078), .A2(n10077), .A3(n10076), .ZN(n10079) );
  NAND2_X1 U12003 ( .A1(n10080), .A2(n10079), .ZN(n10081) );
  NAND2_X1 U12004 ( .A1(n14728), .A2(n10543), .ZN(n10082) );
  NAND2_X1 U12005 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14798) );
  OAI211_X1 U12006 ( .C1(n15951), .C2(n14725), .A(n10082), .B(n14798), .ZN(
        n10083) );
  AOI21_X1 U12007 ( .B1(n16129), .B2(n15949), .A(n10083), .ZN(n10084) );
  OAI21_X1 U12008 ( .B1(n10085), .B2(n16123), .A(n10084), .ZN(P1_U3230) );
  NOR2_X1 U12009 ( .A1(n10086), .A2(n13954), .ZN(n10088) );
  AOI22_X1 U12010 ( .A1(n12602), .A2(n10088), .B1(n15873), .B2(n15875), .ZN(
        n10322) );
  INV_X1 U12011 ( .A(n16101), .ZN(n16155) );
  OAI22_X1 U12012 ( .A1(n16154), .A2(n10104), .B1(n16101), .B2(n9823), .ZN(
        n10089) );
  INV_X1 U12013 ( .A(n10089), .ZN(n10090) );
  OAI21_X1 U12014 ( .B1(n10322), .B2(n16155), .A(n10090), .ZN(P3_U3459) );
  INV_X1 U12015 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10093) );
  NAND2_X1 U12016 ( .A1(n10305), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10091) );
  XNOR2_X1 U12017 ( .A(n10091), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11180) );
  INV_X1 U12018 ( .A(n11180), .ZN(n15468) );
  OAI222_X1 U12019 ( .A1(n14588), .A2(n10093), .B1(n14593), .B2(n10092), .C1(
        n15468), .C2(P2_U3088), .ZN(P2_U3314) );
  OAI21_X1 U12020 ( .B1(n10096), .B2(n10095), .A(n10094), .ZN(n10101) );
  NAND2_X1 U12021 ( .A1(n14150), .A2(n13153), .ZN(n10098) );
  AOI22_X1 U12022 ( .A1(n14141), .A2(n10946), .B1(P2_REG3_REG_5__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10097) );
  OAI211_X1 U12023 ( .C1(n10099), .C2(n14144), .A(n10098), .B(n10097), .ZN(
        n10100) );
  AOI21_X1 U12024 ( .B1(n10101), .B2(n14115), .A(n10100), .ZN(n10102) );
  INV_X1 U12025 ( .A(n10102), .ZN(P2_U3199) );
  INV_X1 U12026 ( .A(n16104), .ZN(n16160) );
  INV_X1 U12027 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10103) );
  OAI22_X1 U12028 ( .A1(n16159), .A2(n10104), .B1(n16104), .B2(n10103), .ZN(
        n10105) );
  INV_X1 U12029 ( .A(n10105), .ZN(n10106) );
  OAI21_X1 U12030 ( .B1(n10322), .B2(n16160), .A(n10106), .ZN(P3_U3390) );
  NOR2_X1 U12031 ( .A1(n13153), .A2(n14196), .ZN(n10107) );
  NAND2_X1 U12032 ( .A1(n13153), .A2(n14196), .ZN(n10109) );
  OR2_X1 U12033 ( .A1(n13161), .A2(n14195), .ZN(n10363) );
  NAND2_X1 U12034 ( .A1(n13161), .A2(n14195), .ZN(n10360) );
  NAND2_X1 U12035 ( .A1(n10363), .A2(n10360), .ZN(n13376) );
  XNOR2_X1 U12036 ( .A(n10362), .B(n13376), .ZN(n10961) );
  AOI21_X1 U12037 ( .B1(n10110), .B2(n13161), .A(n14416), .ZN(n10111) );
  AND2_X1 U12038 ( .A1(n10111), .A2(n10366), .ZN(n10954) );
  OR2_X1 U12039 ( .A1(n13153), .A2(n10114), .ZN(n10112) );
  NAND2_X1 U12040 ( .A1(n13153), .A2(n10114), .ZN(n10115) );
  XOR2_X1 U12041 ( .A(n10367), .B(n13376), .Z(n10117) );
  OAI21_X1 U12042 ( .B1(n10117), .B2(n14413), .A(n10116), .ZN(n10958) );
  AOI211_X1 U12043 ( .C1(n16140), .C2(n10961), .A(n10954), .B(n10958), .ZN(
        n10141) );
  NAND2_X1 U12044 ( .A1(n16142), .A2(n15905), .ZN(n14496) );
  AOI22_X1 U12045 ( .A1(n14524), .A2(n13161), .B1(n16141), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n10118) );
  OAI21_X1 U12046 ( .B1(n10141), .B2(n16141), .A(n10118), .ZN(P2_U3505) );
  AOI21_X1 U12047 ( .B1(n9400), .B2(n10120), .A(n10119), .ZN(n10203) );
  XOR2_X1 U12048 ( .A(n11230), .B(n10203), .Z(n10122) );
  INV_X1 U12049 ( .A(n10122), .ZN(n10124) );
  INV_X1 U12050 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10121) );
  NAND2_X1 U12051 ( .A1(n10122), .A2(n10121), .ZN(n10208) );
  INV_X1 U12052 ( .A(n10208), .ZN(n10123) );
  AOI21_X1 U12053 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n10124), .A(n10123), 
        .ZN(n10135) );
  INV_X1 U12054 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10125) );
  NAND2_X1 U12055 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n11821)
         );
  OAI21_X1 U12056 ( .B1(n14842), .B2(n10125), .A(n11821), .ZN(n10126) );
  AOI21_X1 U12057 ( .B1(n11230), .B2(n14787), .A(n10126), .ZN(n10133) );
  AOI21_X1 U12058 ( .B1(n11036), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10127), 
        .ZN(n10130) );
  INV_X1 U12059 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10128) );
  MUX2_X1 U12060 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n10128), .S(n11230), .Z(
        n10129) );
  NOR2_X1 U12061 ( .A1(n10130), .A2(n10129), .ZN(n10131) );
  OAI21_X1 U12062 ( .B1(n10131), .B2(n10210), .A(n14833), .ZN(n10132) );
  OAI211_X1 U12063 ( .C1(n10135), .C2(n10134), .A(n10133), .B(n10132), .ZN(
        P1_U3255) );
  OR2_X1 U12064 ( .A1(n10137), .A2(n16143), .ZN(n10138) );
  OAI21_X1 U12065 ( .B1(n16146), .B2(n9910), .A(n10138), .ZN(P2_U3445) );
  NAND2_X1 U12066 ( .A1(n16146), .A2(n15905), .ZN(n14566) );
  INV_X1 U12067 ( .A(n14566), .ZN(n14578) );
  NOR2_X1 U12068 ( .A1(n16146), .A2(n9983), .ZN(n10139) );
  AOI21_X1 U12069 ( .B1(n14578), .B2(n13161), .A(n10139), .ZN(n10140) );
  OAI21_X1 U12070 ( .B1(n10141), .B2(n16143), .A(n10140), .ZN(P2_U3448) );
  NAND2_X1 U12071 ( .A1(n10143), .A2(n10142), .ZN(n10145) );
  MUX2_X1 U12072 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n13664), .Z(n10173) );
  XNOR2_X1 U12073 ( .A(n10173), .B(n10174), .ZN(n10144) );
  NAND2_X1 U12074 ( .A1(n10145), .A2(n10144), .ZN(n10177) );
  OAI21_X1 U12075 ( .B1(n10145), .B2(n10144), .A(n10177), .ZN(n10146) );
  NAND2_X1 U12076 ( .A1(n10146), .A2(n15775), .ZN(n10164) );
  OR2_X1 U12077 ( .A1(n10151), .A2(n10147), .ZN(n10148) );
  NAND2_X1 U12078 ( .A1(n10149), .A2(n10148), .ZN(n10185) );
  XNOR2_X1 U12079 ( .A(n10185), .B(n10174), .ZN(n10150) );
  OAI21_X1 U12080 ( .B1(n10150), .B2(P3_REG1_REG_5__SCAN_IN), .A(n7586), .ZN(
        n10161) );
  OR2_X1 U12081 ( .A1(n10151), .A2(n11028), .ZN(n10152) );
  NAND2_X1 U12082 ( .A1(n10153), .A2(n10152), .ZN(n10190) );
  NAND2_X1 U12083 ( .A1(n10154), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n10192) );
  OAI21_X1 U12084 ( .B1(n10154), .B2(P3_REG2_REG_5__SCAN_IN), .A(n10192), .ZN(
        n10155) );
  INV_X1 U12085 ( .A(n10155), .ZN(n10158) );
  AND2_X1 U12086 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n11115) );
  INV_X1 U12087 ( .A(n11115), .ZN(n10157) );
  NAND2_X1 U12088 ( .A1(n15771), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n10156) );
  OAI211_X1 U12089 ( .C1(n15825), .C2(n10158), .A(n10157), .B(n10156), .ZN(
        n10160) );
  INV_X1 U12090 ( .A(n10174), .ZN(n10189) );
  NOR2_X1 U12091 ( .A1(n15773), .A2(n10189), .ZN(n10159) );
  AOI211_X1 U12092 ( .C1(n10162), .C2(n10161), .A(n10160), .B(n10159), .ZN(
        n10163) );
  NAND2_X1 U12093 ( .A1(n10164), .A2(n10163), .ZN(P3_U3187) );
  AOI21_X1 U12094 ( .B1(n10167), .B2(n10166), .A(n10165), .ZN(n10172) );
  INV_X1 U12095 ( .A(n13548), .ZN(n13529) );
  OAI22_X1 U12096 ( .A1(n13519), .A2(n10636), .B1(n8787), .B2(n13554), .ZN(
        n10170) );
  NOR2_X1 U12097 ( .A1(n10397), .A2(n10168), .ZN(n10169) );
  AOI211_X1 U12098 ( .C1(n13529), .C2(n13578), .A(n10170), .B(n10169), .ZN(
        n10171) );
  OAI21_X1 U12099 ( .B1(n10172), .B2(n13539), .A(n10171), .ZN(P3_U3162) );
  INV_X1 U12100 ( .A(n10173), .ZN(n10175) );
  NAND2_X1 U12101 ( .A1(n10175), .A2(n10174), .ZN(n10176) );
  NAND2_X1 U12102 ( .A1(n10177), .A2(n10176), .ZN(n10757) );
  MUX2_X1 U12103 ( .A(n10179), .B(n10178), .S(n13664), .Z(n10180) );
  INV_X1 U12104 ( .A(n10772), .ZN(n10200) );
  AND2_X1 U12105 ( .A1(n10180), .A2(n10200), .ZN(n10756) );
  INV_X1 U12106 ( .A(n10756), .ZN(n10182) );
  INV_X1 U12107 ( .A(n10180), .ZN(n10181) );
  NAND2_X1 U12108 ( .A1(n10181), .A2(n10772), .ZN(n10758) );
  NAND2_X1 U12109 ( .A1(n10182), .A2(n10758), .ZN(n10183) );
  XNOR2_X1 U12110 ( .A(n10757), .B(n10183), .ZN(n10202) );
  AOI22_X1 U12111 ( .A1(n10200), .A2(P3_REG1_REG_6__SCAN_IN), .B1(n10178), 
        .B2(n10772), .ZN(n10186) );
  AOI21_X1 U12112 ( .B1(n10187), .B2(n10186), .A(n7332), .ZN(n10188) );
  NOR2_X1 U12113 ( .A1(n15822), .A2(n10188), .ZN(n10199) );
  NAND2_X1 U12114 ( .A1(n10190), .A2(n10189), .ZN(n10191) );
  AOI22_X1 U12115 ( .A1(n10200), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n10179), 
        .B2(n10772), .ZN(n10193) );
  AOI21_X1 U12116 ( .B1(n10194), .B2(n10193), .A(n10771), .ZN(n10197) );
  INV_X1 U12117 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n15275) );
  NOR2_X1 U12118 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15275), .ZN(n11210) );
  INV_X1 U12119 ( .A(n11210), .ZN(n10196) );
  NAND2_X1 U12120 ( .A1(n15771), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n10195) );
  OAI211_X1 U12121 ( .C1(n15825), .C2(n10197), .A(n10196), .B(n10195), .ZN(
        n10198) );
  AOI211_X1 U12122 ( .C1(n15817), .C2(n10200), .A(n10199), .B(n10198), .ZN(
        n10201) );
  OAI21_X1 U12123 ( .B1(n10202), .B2(n15811), .A(n10201), .ZN(P3_U3188) );
  INV_X1 U12124 ( .A(n10203), .ZN(n10205) );
  NAND2_X1 U12125 ( .A1(n10205), .A2(n10204), .ZN(n10206) );
  INV_X1 U12126 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10611) );
  XNOR2_X1 U12127 ( .A(n11413), .B(n10611), .ZN(n10207) );
  AOI21_X1 U12128 ( .B1(n10208), .B2(n10206), .A(n10207), .ZN(n10217) );
  NAND3_X1 U12129 ( .A1(n10208), .A2(n10207), .A3(n10206), .ZN(n10610) );
  NAND2_X1 U12130 ( .A1(n10610), .A2(n14834), .ZN(n10216) );
  INV_X1 U12131 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n15594) );
  NAND2_X1 U12132 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n11934)
         );
  OAI21_X1 U12133 ( .B1(n14842), .B2(n15594), .A(n11934), .ZN(n10214) );
  XNOR2_X1 U12134 ( .A(n11413), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n10212) );
  NOR2_X1 U12135 ( .A1(n11230), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10209) );
  OR2_X1 U12136 ( .A1(n10210), .A2(n10209), .ZN(n10211) );
  NOR3_X1 U12137 ( .A1(n10210), .A2(n10209), .A3(n10212), .ZN(n10608) );
  AOI211_X1 U12138 ( .C1(n10212), .C2(n10211), .A(n14829), .B(n10608), .ZN(
        n10213) );
  AOI211_X1 U12139 ( .C1(n14787), .C2(n11413), .A(n10214), .B(n10213), .ZN(
        n10215) );
  OAI21_X1 U12140 ( .B1(n10217), .B2(n10216), .A(n10215), .ZN(P1_U3256) );
  NAND2_X1 U12141 ( .A1(n10221), .A2(n12089), .ZN(n10224) );
  AOI22_X1 U12142 ( .A1(n13011), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n12008), 
        .B2(n10222), .ZN(n10223) );
  NAND2_X1 U12143 ( .A1(n10224), .A2(n10223), .ZN(n12832) );
  NAND2_X1 U12144 ( .A1(n12832), .A2(n7181), .ZN(n10227) );
  NAND2_X1 U12145 ( .A1(n14748), .A2(n12519), .ZN(n10226) );
  NAND2_X1 U12146 ( .A1(n10227), .A2(n10226), .ZN(n10228) );
  XNOR2_X1 U12147 ( .A(n10228), .B(n12526), .ZN(n10232) );
  NAND2_X1 U12148 ( .A1(n12832), .A2(n12519), .ZN(n10230) );
  NAND2_X1 U12149 ( .A1(n12518), .A2(n14748), .ZN(n10229) );
  NAND2_X1 U12150 ( .A1(n10230), .A2(n10229), .ZN(n10231) );
  NOR2_X1 U12151 ( .A1(n10232), .A2(n10231), .ZN(n10382) );
  INV_X1 U12152 ( .A(n10382), .ZN(n10233) );
  NAND2_X1 U12153 ( .A1(n10232), .A2(n10231), .ZN(n10381) );
  NAND2_X1 U12154 ( .A1(n10233), .A2(n10381), .ZN(n10234) );
  XNOR2_X1 U12155 ( .A(n10383), .B(n10234), .ZN(n10248) );
  AND2_X1 U12156 ( .A1(n12832), .A2(n15948), .ZN(n15973) );
  INV_X2 U12157 ( .A(n11659), .ZN(n12987) );
  NAND2_X1 U12158 ( .A1(n12987), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10243) );
  NAND2_X1 U12159 ( .A1(n10235), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10266) );
  INV_X1 U12160 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n10236) );
  NAND2_X1 U12161 ( .A1(n10237), .A2(n10236), .ZN(n10238) );
  AND2_X1 U12162 ( .A1(n10266), .A2(n10238), .ZN(n15989) );
  NAND2_X1 U12163 ( .A1(n12095), .A2(n15989), .ZN(n10242) );
  INV_X2 U12164 ( .A(n10239), .ZN(n12988) );
  NAND2_X1 U12165 ( .A1(n12988), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10241) );
  NAND2_X1 U12166 ( .A1(n12014), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n10240) );
  NAND4_X1 U12167 ( .A1(n10243), .A2(n10242), .A3(n10241), .A4(n10240), .ZN(
        n14747) );
  AOI22_X1 U12168 ( .A1(n14978), .A2(n14749), .B1(n14747), .B2(n14980), .ZN(
        n10674) );
  NAND2_X1 U12169 ( .A1(n14728), .A2(n10680), .ZN(n10245) );
  OAI211_X1 U12170 ( .C1(n10674), .C2(n14725), .A(n10245), .B(n10244), .ZN(
        n10246) );
  AOI21_X1 U12171 ( .B1(n15921), .B2(n15973), .A(n10246), .ZN(n10247) );
  OAI21_X1 U12172 ( .B1(n10248), .B2(n16123), .A(n10247), .ZN(P1_U3227) );
  INV_X1 U12173 ( .A(n13026), .ZN(n10249) );
  NAND2_X1 U12174 ( .A1(n10250), .A2(n10249), .ZN(n10252) );
  NAND2_X1 U12175 ( .A1(n10252), .A2(n10251), .ZN(n10618) );
  INV_X1 U12176 ( .A(n13027), .ZN(n10253) );
  NAND2_X1 U12177 ( .A1(n10618), .A2(n10253), .ZN(n10255) );
  NAND2_X1 U12178 ( .A1(n10273), .A2(n10275), .ZN(n10254) );
  NAND2_X1 U12179 ( .A1(n10255), .A2(n10254), .ZN(n10539) );
  INV_X1 U12180 ( .A(n14749), .ZN(n10278) );
  XNOR2_X1 U12181 ( .A(n15949), .B(n10278), .ZN(n13029) );
  NAND2_X1 U12182 ( .A1(n10539), .A2(n13029), .ZN(n10257) );
  OR2_X1 U12183 ( .A1(n15949), .A2(n14749), .ZN(n10256) );
  NAND2_X1 U12184 ( .A1(n10257), .A2(n10256), .ZN(n10671) );
  XNOR2_X1 U12185 ( .A(n12832), .B(n14748), .ZN(n13031) );
  INV_X1 U12186 ( .A(n13031), .ZN(n10258) );
  NAND2_X1 U12187 ( .A1(n10671), .A2(n10258), .ZN(n10260) );
  OR2_X1 U12188 ( .A1(n12832), .A2(n14748), .ZN(n10259) );
  NAND2_X1 U12189 ( .A1(n10260), .A2(n10259), .ZN(n10469) );
  NAND2_X1 U12190 ( .A1(n10261), .A2(n12089), .ZN(n10264) );
  AOI22_X1 U12191 ( .A1(n13011), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n12008), 
        .B2(n10262), .ZN(n10263) );
  NAND2_X1 U12192 ( .A1(n10264), .A2(n10263), .ZN(n15991) );
  XNOR2_X1 U12193 ( .A(n15991), .B(n14747), .ZN(n13032) );
  XNOR2_X1 U12194 ( .A(n10469), .B(n13032), .ZN(n15992) );
  NAND2_X1 U12195 ( .A1(n12987), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10271) );
  NAND2_X1 U12196 ( .A1(n10266), .A2(n10265), .ZN(n10267) );
  AND2_X1 U12197 ( .A1(n10481), .A2(n10267), .ZN(n10644) );
  NAND2_X1 U12198 ( .A1(n12095), .A2(n10644), .ZN(n10270) );
  NAND2_X1 U12199 ( .A1(n12988), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10269) );
  NAND2_X1 U12200 ( .A1(n12014), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n10268) );
  NAND4_X1 U12201 ( .A1(n10271), .A2(n10270), .A3(n10269), .A4(n10268), .ZN(
        n14746) );
  AOI22_X1 U12202 ( .A1(n14978), .A2(n14748), .B1(n14746), .B2(n14980), .ZN(
        n10389) );
  NAND2_X1 U12203 ( .A1(n10624), .A2(n12802), .ZN(n12816) );
  NAND2_X1 U12204 ( .A1(n10273), .A2(n14750), .ZN(n10274) );
  NAND2_X1 U12205 ( .A1(n10275), .A2(n15918), .ZN(n10276) );
  OR2_X1 U12206 ( .A1(n10278), .A2(n15949), .ZN(n10279) );
  NAND2_X1 U12207 ( .A1(n15956), .A2(n10279), .ZN(n10673) );
  INV_X1 U12208 ( .A(n14748), .ZN(n10280) );
  OR2_X1 U12209 ( .A1(n12832), .A2(n10280), .ZN(n10281) );
  OAI211_X1 U12210 ( .C1(n10282), .C2(n13032), .A(n10492), .B(n15955), .ZN(
        n10283) );
  OAI211_X1 U12211 ( .C1(n15992), .C2(n15977), .A(n10389), .B(n10283), .ZN(
        n10284) );
  INV_X1 U12212 ( .A(n10284), .ZN(n15997) );
  INV_X1 U12213 ( .A(n12832), .ZN(n10682) );
  INV_X1 U12214 ( .A(n10678), .ZN(n10285) );
  INV_X1 U12215 ( .A(n15991), .ZN(n10393) );
  AOI211_X1 U12216 ( .C1(n15991), .C2(n10285), .A(n15952), .B(n10479), .ZN(
        n15993) );
  AOI21_X1 U12217 ( .B1(n15948), .B2(n15991), .A(n15993), .ZN(n10286) );
  OAI211_X1 U12218 ( .C1(n15856), .C2(n15992), .A(n15997), .B(n10286), .ZN(
        n10291) );
  NAND2_X1 U12219 ( .A1(n10291), .A2(n16067), .ZN(n10287) );
  OAI21_X1 U12220 ( .B1(n16067), .B2(n10288), .A(n10287), .ZN(P1_U3534) );
  INV_X1 U12221 ( .A(n10534), .ZN(n10290) );
  INV_X1 U12222 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10293) );
  NAND2_X1 U12223 ( .A1(n10291), .A2(n16071), .ZN(n10292) );
  OAI21_X1 U12224 ( .B1(n16071), .B2(n10293), .A(n10292), .ZN(P1_U3477) );
  INV_X1 U12225 ( .A(n10294), .ZN(n10295) );
  NAND2_X1 U12226 ( .A1(n10297), .A2(SI_13_), .ZN(n10298) );
  MUX2_X1 U12227 ( .A(n11489), .B(n10304), .S(n7178), .Z(n10299) );
  INV_X1 U12228 ( .A(n10299), .ZN(n10300) );
  NAND2_X1 U12229 ( .A1(n10300), .A2(SI_14_), .ZN(n10301) );
  NAND2_X1 U12230 ( .A1(n10433), .A2(n10301), .ZN(n10434) );
  XNOR2_X1 U12231 ( .A(n10435), .B(n10434), .ZN(n11488) );
  INV_X1 U12232 ( .A(n11488), .ZN(n10308) );
  NAND2_X1 U12233 ( .A1(n10302), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10303) );
  XNOR2_X1 U12234 ( .A(n10303), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11409) );
  INV_X1 U12235 ( .A(n11409), .ZN(n10800) );
  OAI222_X1 U12236 ( .A1(n15157), .A2(n10304), .B1(n15167), .B2(n10308), .C1(
        P1_U3086), .C2(n10800), .ZN(P1_U3341) );
  NAND2_X1 U12237 ( .A1(n10590), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10307) );
  INV_X1 U12238 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n10306) );
  XNOR2_X1 U12239 ( .A(n10307), .B(n10306), .ZN(n11769) );
  OAI222_X1 U12240 ( .A1(n14588), .A2(n11489), .B1(n14593), .B2(n10308), .C1(
        P2_U3088), .C2(n11769), .ZN(P2_U3313) );
  INV_X1 U12241 ( .A(n10309), .ZN(n10313) );
  NAND2_X1 U12242 ( .A1(n10312), .A2(n10310), .ZN(n10311) );
  OAI21_X1 U12243 ( .B1(n10313), .B2(n10312), .A(n10311), .ZN(n10314) );
  INV_X1 U12244 ( .A(n10314), .ZN(n10315) );
  INV_X1 U12245 ( .A(n10317), .ZN(n10318) );
  NOR2_X1 U12246 ( .A1(n16096), .A2(n15893), .ZN(n10525) );
  NAND2_X2 U12247 ( .A1(n10318), .A2(n10525), .ZN(n13882) );
  INV_X1 U12248 ( .A(n13882), .ZN(n15399) );
  AOI22_X1 U12249 ( .A1(n15399), .A2(n10319), .B1(n13829), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n10321) );
  NAND2_X1 U12250 ( .A1(n13853), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10320) );
  OAI211_X1 U12251 ( .C1(n10322), .C2(n13853), .A(n10321), .B(n10320), .ZN(
        P3_U3233) );
  INV_X1 U12252 ( .A(n13647), .ZN(n13661) );
  INV_X1 U12253 ( .A(n10323), .ZN(n10324) );
  OAI222_X1 U12254 ( .A1(P3_U3151), .A2(n13661), .B1(n13083), .B2(n15184), 
        .C1(n13082), .C2(n10324), .ZN(P3_U3277) );
  AOI22_X1 U12255 ( .A1(n13330), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n10325), 
        .B2(n12234), .ZN(n10326) );
  INV_X1 U12256 ( .A(n13170), .ZN(n10584) );
  INV_X1 U12257 ( .A(n10330), .ZN(n10333) );
  INV_X1 U12258 ( .A(n10331), .ZN(n10332) );
  XNOR2_X1 U12259 ( .A(n13170), .B(n14032), .ZN(n10336) );
  NAND2_X1 U12260 ( .A1(n14194), .A2(n14416), .ZN(n10337) );
  NAND2_X1 U12261 ( .A1(n10336), .A2(n10337), .ZN(n10445) );
  INV_X1 U12262 ( .A(n10336), .ZN(n10339) );
  INV_X1 U12263 ( .A(n10337), .ZN(n10338) );
  NAND2_X1 U12264 ( .A1(n10339), .A2(n10338), .ZN(n10340) );
  OAI21_X1 U12265 ( .B1(n10342), .B2(n10341), .A(n10446), .ZN(n10343) );
  NAND2_X1 U12266 ( .A1(n10343), .A2(n14115), .ZN(n10359) );
  NAND2_X1 U12267 ( .A1(n14195), .A2(n14137), .ZN(n10354) );
  NAND2_X1 U12268 ( .A1(n13322), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10352) );
  NAND2_X1 U12269 ( .A1(n10345), .A2(n10344), .ZN(n10346) );
  NAND2_X1 U12270 ( .A1(n10453), .A2(n10346), .ZN(n10464) );
  INV_X1 U12271 ( .A(n10464), .ZN(n10967) );
  NAND2_X1 U12272 ( .A1(n12342), .A2(n10967), .ZN(n10351) );
  OR2_X1 U12273 ( .A1(n12239), .A2(n10347), .ZN(n10350) );
  INV_X1 U12274 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10348) );
  OR2_X1 U12275 ( .A1(n13325), .A2(n10348), .ZN(n10349) );
  NAND4_X1 U12276 ( .A1(n10352), .A2(n10351), .A3(n10350), .A4(n10349), .ZN(
        n14193) );
  NAND2_X1 U12277 ( .A1(n14193), .A2(n14139), .ZN(n10353) );
  NAND2_X1 U12278 ( .A1(n10354), .A2(n10353), .ZN(n10371) );
  INV_X1 U12279 ( .A(n10355), .ZN(n10583) );
  OAI21_X1 U12280 ( .B1(n14161), .B2(n10583), .A(n10356), .ZN(n10357) );
  AOI21_X1 U12281 ( .B1(n14165), .B2(n10371), .A(n10357), .ZN(n10358) );
  OAI211_X1 U12282 ( .C1(n10584), .C2(n14162), .A(n10359), .B(n10358), .ZN(
        P2_U3185) );
  INV_X1 U12283 ( .A(n10360), .ZN(n10361) );
  INV_X1 U12284 ( .A(n14194), .ZN(n10561) );
  XNOR2_X1 U12285 ( .A(n13170), .B(n10561), .ZN(n13378) );
  OR2_X1 U12286 ( .A1(n10364), .A2(n13378), .ZN(n10365) );
  NAND2_X1 U12287 ( .A1(n10555), .A2(n10365), .ZN(n10580) );
  AOI211_X1 U12288 ( .C1(n13170), .C2(n10366), .A(n14416), .B(n7682), .ZN(
        n10586) );
  NAND2_X1 U12289 ( .A1(n10367), .A2(n13376), .ZN(n10370) );
  INV_X1 U12290 ( .A(n14195), .ZN(n10368) );
  NAND2_X1 U12291 ( .A1(n13161), .A2(n10368), .ZN(n10369) );
  XNOR2_X1 U12292 ( .A(n10560), .B(n13378), .ZN(n10374) );
  INV_X1 U12293 ( .A(n16107), .ZN(n15907) );
  NAND2_X1 U12294 ( .A1(n10580), .A2(n15907), .ZN(n10373) );
  INV_X1 U12295 ( .A(n10371), .ZN(n10372) );
  OAI211_X1 U12296 ( .C1(n14413), .C2(n10374), .A(n10373), .B(n10372), .ZN(
        n10581) );
  AOI211_X1 U12297 ( .C1(n16092), .C2(n10580), .A(n10586), .B(n10581), .ZN(
        n10378) );
  OAI22_X1 U12298 ( .A1(n14566), .A2(n10584), .B1(n16146), .B2(n10011), .ZN(
        n10375) );
  INV_X1 U12299 ( .A(n10375), .ZN(n10376) );
  OAI21_X1 U12300 ( .B1(n10378), .B2(n16143), .A(n10376), .ZN(P2_U3451) );
  AOI22_X1 U12301 ( .A1(n14524), .A2(n13170), .B1(n16141), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n10377) );
  OAI21_X1 U12302 ( .B1(n10378), .B2(n16141), .A(n10377), .ZN(P2_U3506) );
  INV_X1 U12303 ( .A(n10379), .ZN(n10380) );
  OAI222_X1 U12304 ( .A1(P3_U3151), .A2(n13656), .B1(n13082), .B2(n10380), 
        .C1(n15180), .C2(n13083), .ZN(P3_U3276) );
  INV_X1 U12305 ( .A(n14747), .ZN(n10491) );
  OAI22_X1 U12306 ( .A1(n10393), .A2(n12523), .B1(n10491), .B2(n12525), .ZN(
        n10384) );
  XNOR2_X1 U12307 ( .A(n10384), .B(n12526), .ZN(n10593) );
  AND2_X1 U12308 ( .A1(n12518), .A2(n14747), .ZN(n10385) );
  AOI21_X1 U12309 ( .B1(n15991), .B2(n12519), .A(n10385), .ZN(n10596) );
  XNOR2_X1 U12310 ( .A(n10593), .B(n10596), .ZN(n10386) );
  OAI211_X1 U12311 ( .C1(n10387), .C2(n10386), .A(n10594), .B(n14719), .ZN(
        n10392) );
  OAI21_X1 U12312 ( .B1(n14725), .B2(n10389), .A(n10388), .ZN(n10390) );
  AOI21_X1 U12313 ( .B1(n14728), .B2(n15989), .A(n10390), .ZN(n10391) );
  OAI211_X1 U12314 ( .C1(n10393), .C2(n14731), .A(n10392), .B(n10391), .ZN(
        P1_U3239) );
  AOI21_X1 U12315 ( .B1(n10396), .B2(n10395), .A(n10394), .ZN(n10401) );
  OAI22_X1 U12316 ( .A1(n13519), .A2(n10988), .B1(n13554), .B2(n15872), .ZN(
        n10399) );
  NOR2_X1 U12317 ( .A1(n10397), .A2(n15891), .ZN(n10398) );
  AOI211_X1 U12318 ( .C1(n13529), .C2(n15875), .A(n10399), .B(n10398), .ZN(
        n10400) );
  OAI21_X1 U12319 ( .B1(n10401), .B2(n13539), .A(n10400), .ZN(P3_U3177) );
  INV_X1 U12320 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n16113) );
  MUX2_X1 U12321 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n16113), .S(n11180), .Z(
        n15474) );
  INV_X1 U12322 ( .A(n10402), .ZN(n10403) );
  AOI21_X1 U12323 ( .B1(n16093), .B2(n10404), .A(n10403), .ZN(n15475) );
  NAND2_X1 U12324 ( .A1(n15474), .A2(n15475), .ZN(n15472) );
  OAI21_X1 U12325 ( .B1(n15468), .B2(n16113), .A(n15472), .ZN(n10407) );
  INV_X1 U12326 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10405) );
  MUX2_X1 U12327 ( .A(n10405), .B(P2_REG1_REG_14__SCAN_IN), .S(n11769), .Z(
        n10406) );
  NAND2_X1 U12328 ( .A1(n10406), .A2(n10407), .ZN(n11759) );
  OAI211_X1 U12329 ( .C1(n10407), .C2(n10406), .A(n15473), .B(n11759), .ZN(
        n10419) );
  NAND2_X1 U12330 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n11707)
         );
  NAND2_X1 U12331 ( .A1(n11180), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10413) );
  NOR2_X1 U12332 ( .A1(n11137), .A2(n10408), .ZN(n10410) );
  NOR2_X1 U12333 ( .A1(n10410), .A2(n10409), .ZN(n15479) );
  INV_X1 U12334 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10411) );
  MUX2_X1 U12335 ( .A(n10411), .B(P2_REG2_REG_13__SCAN_IN), .S(n11180), .Z(
        n10412) );
  INV_X1 U12336 ( .A(n10412), .ZN(n15478) );
  NAND2_X1 U12337 ( .A1(n15479), .A2(n15478), .ZN(n15476) );
  NAND2_X1 U12338 ( .A1(n10413), .A2(n15476), .ZN(n10415) );
  INV_X1 U12339 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11505) );
  MUX2_X1 U12340 ( .A(n11505), .B(P2_REG2_REG_14__SCAN_IN), .S(n11769), .Z(
        n10414) );
  NAND2_X1 U12341 ( .A1(n10414), .A2(n10415), .ZN(n11768) );
  OAI211_X1 U12342 ( .C1(n10415), .C2(n10414), .A(n15477), .B(n11768), .ZN(
        n10416) );
  NAND2_X1 U12343 ( .A1(n11707), .A2(n10416), .ZN(n10417) );
  AOI21_X1 U12344 ( .B1(n15471), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n10417), 
        .ZN(n10418) );
  OAI211_X1 U12345 ( .C1(n15466), .C2(n11769), .A(n10419), .B(n10418), .ZN(
        P2_U3228) );
  XOR2_X1 U12346 ( .A(n10420), .B(n7361), .Z(n10426) );
  INV_X1 U12347 ( .A(n10426), .ZN(n10529) );
  OAI21_X1 U12348 ( .B1(n10421), .B2(n7361), .A(n15880), .ZN(n10424) );
  OAI22_X1 U12349 ( .A1(n10422), .A2(n15392), .B1(n10636), .B2(n15390), .ZN(
        n10423) );
  AOI21_X1 U12350 ( .B1(n10424), .B2(n15881), .A(n10423), .ZN(n10425) );
  OAI21_X1 U12351 ( .B1(n10426), .B2(n15886), .A(n10425), .ZN(n10523) );
  AOI21_X1 U12352 ( .B1(n16082), .B2(n10529), .A(n10523), .ZN(n10432) );
  OAI22_X1 U12353 ( .A1(n16154), .A2(n8787), .B1(n16101), .B2(n9818), .ZN(
        n10427) );
  INV_X1 U12354 ( .A(n10427), .ZN(n10428) );
  OAI21_X1 U12355 ( .B1(n10432), .B2(n16155), .A(n10428), .ZN(P3_U3460) );
  INV_X1 U12356 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n10429) );
  OAI22_X1 U12357 ( .A1(n16159), .A2(n8787), .B1(n16104), .B2(n10429), .ZN(
        n10430) );
  INV_X1 U12358 ( .A(n10430), .ZN(n10431) );
  OAI21_X1 U12359 ( .B1(n10432), .B2(n16160), .A(n10431), .ZN(P3_U3393) );
  MUX2_X1 U12360 ( .A(n10592), .B(n10436), .S(n7178), .Z(n10438) );
  INV_X1 U12361 ( .A(n10438), .ZN(n10439) );
  NAND2_X1 U12362 ( .A1(n10439), .A2(SI_15_), .ZN(n10440) );
  XNOR2_X1 U12363 ( .A(n10887), .B(n10886), .ZN(n11626) );
  INV_X1 U12364 ( .A(n11626), .ZN(n10591) );
  NAND2_X1 U12365 ( .A1(n10442), .A2(n7926), .ZN(n10889) );
  NAND2_X1 U12366 ( .A1(n10889), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10443) );
  XNOR2_X1 U12367 ( .A(n10443), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11627) );
  AOI22_X1 U12368 ( .A1(n11627), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n15164), .ZN(n10444) );
  OAI21_X1 U12369 ( .B1(n10591), .B2(n15167), .A(n10444), .ZN(P1_U3340) );
  AOI22_X1 U12370 ( .A1(n10447), .A2(n12234), .B1(n13330), .B2(
        P1_DATAO_REG_8__SCAN_IN), .ZN(n10448) );
  NAND2_X1 U12371 ( .A1(n10449), .A2(n10448), .ZN(n13177) );
  XNOR2_X1 U12372 ( .A(n13177), .B(n14032), .ZN(n10844) );
  NAND2_X1 U12373 ( .A1(n14193), .A2(n14416), .ZN(n10847) );
  NOR2_X1 U12374 ( .A1(n10844), .A2(n10847), .ZN(n10845) );
  AOI21_X1 U12375 ( .B1(n10844), .B2(n10847), .A(n10845), .ZN(n10450) );
  XNOR2_X1 U12376 ( .A(n12399), .B(n10450), .ZN(n10467) );
  NAND2_X1 U12377 ( .A1(n14194), .A2(n14137), .ZN(n10461) );
  NAND2_X1 U12378 ( .A1(n13322), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n10459) );
  INV_X1 U12379 ( .A(n10453), .ZN(n10451) );
  INV_X1 U12380 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10452) );
  NAND2_X1 U12381 ( .A1(n10453), .A2(n10452), .ZN(n10454) );
  AND2_X1 U12382 ( .A1(n10696), .A2(n10454), .ZN(n14429) );
  NAND2_X1 U12383 ( .A1(n12342), .A2(n14429), .ZN(n10458) );
  OR2_X1 U12384 ( .A1(n12239), .A2(n14432), .ZN(n10457) );
  INV_X1 U12385 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10455) );
  OR2_X1 U12386 ( .A1(n13325), .A2(n10455), .ZN(n10456) );
  NAND4_X1 U12387 ( .A1(n10459), .A2(n10458), .A3(n10457), .A4(n10456), .ZN(
        n14191) );
  NAND2_X1 U12388 ( .A1(n14191), .A2(n14139), .ZN(n10460) );
  NAND2_X1 U12389 ( .A1(n10461), .A2(n10460), .ZN(n10972) );
  NAND2_X1 U12390 ( .A1(n14165), .A2(n10972), .ZN(n10463) );
  OAI211_X1 U12391 ( .C1(n14161), .C2(n10464), .A(n10463), .B(n10462), .ZN(
        n10465) );
  AOI21_X1 U12392 ( .B1(n13177), .B2(n14150), .A(n10465), .ZN(n10466) );
  OAI21_X1 U12393 ( .B1(n10467), .B2(n14168), .A(n10466), .ZN(P2_U3193) );
  INV_X1 U12394 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10498) );
  INV_X1 U12395 ( .A(n15856), .ZN(n16017) );
  NOR2_X1 U12396 ( .A1(n15991), .A2(n14747), .ZN(n10468) );
  NAND2_X1 U12397 ( .A1(n15991), .A2(n14747), .ZN(n10470) );
  NAND2_X1 U12398 ( .A1(n10472), .A2(n12089), .ZN(n10475) );
  AOI22_X1 U12399 ( .A1(n13011), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n12008), 
        .B2(n10473), .ZN(n10474) );
  NAND2_X1 U12400 ( .A1(n10475), .A2(n10474), .ZN(n12844) );
  XNOR2_X1 U12401 ( .A(n12844), .B(n14746), .ZN(n13034) );
  NAND2_X1 U12402 ( .A1(n10477), .A2(n13034), .ZN(n10478) );
  NAND2_X1 U12403 ( .A1(n10730), .A2(n10478), .ZN(n10650) );
  OAI211_X1 U12404 ( .C1(n10479), .C2(n7595), .A(n15041), .B(n10751), .ZN(
        n10646) );
  OAI21_X1 U12405 ( .B1(n7595), .B2(n16058), .A(n10646), .ZN(n10496) );
  NAND2_X1 U12406 ( .A1(n12987), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10487) );
  NAND2_X1 U12407 ( .A1(n10481), .A2(n10480), .ZN(n10482) );
  NAND2_X1 U12408 ( .A1(n10737), .A2(n10482), .ZN(n10825) );
  INV_X1 U12409 ( .A(n10825), .ZN(n10483) );
  NAND2_X1 U12410 ( .A1(n12095), .A2(n10483), .ZN(n10486) );
  NAND2_X1 U12411 ( .A1(n12988), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10485) );
  NAND2_X1 U12412 ( .A1(n12014), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10484) );
  NAND4_X1 U12413 ( .A1(n10487), .A2(n10486), .A3(n10485), .A4(n10484), .ZN(
        n14745) );
  NAND2_X1 U12414 ( .A1(n14745), .A2(n14980), .ZN(n10489) );
  NAND2_X1 U12415 ( .A1(n14747), .A2(n14978), .ZN(n10488) );
  NAND2_X1 U12416 ( .A1(n10489), .A2(n10488), .ZN(n10490) );
  AOI21_X1 U12417 ( .B1(n10650), .B2(n16034), .A(n10490), .ZN(n10495) );
  XNOR2_X1 U12418 ( .A(n10744), .B(n10476), .ZN(n10493) );
  NAND2_X1 U12419 ( .A1(n10493), .A2(n15955), .ZN(n10494) );
  NAND2_X1 U12420 ( .A1(n10495), .A2(n10494), .ZN(n10647) );
  AOI211_X1 U12421 ( .C1(n16017), .C2(n10650), .A(n10496), .B(n10647), .ZN(
        n10499) );
  OR2_X1 U12422 ( .A1(n10499), .A2(n16068), .ZN(n10497) );
  OAI21_X1 U12423 ( .B1(n16071), .B2(n10498), .A(n10497), .ZN(P1_U3480) );
  OR2_X1 U12424 ( .A1(n10499), .A2(n16066), .ZN(n10500) );
  OAI21_X1 U12425 ( .B1(n16067), .B2(n10501), .A(n10500), .ZN(P1_U3535) );
  INV_X1 U12426 ( .A(n10502), .ZN(n10503) );
  AND3_X1 U12427 ( .A1(n15408), .A2(n10504), .A3(n10503), .ZN(n10505) );
  NAND2_X1 U12428 ( .A1(n15409), .A2(n10505), .ZN(n10515) );
  INV_X2 U12429 ( .A(n14378), .ZN(n14427) );
  INV_X1 U12430 ( .A(n13100), .ZN(n10507) );
  NAND2_X1 U12431 ( .A1(n16107), .A2(n10507), .ZN(n10508) );
  NAND2_X1 U12432 ( .A1(n14427), .A2(n10508), .ZN(n14303) );
  XNOR2_X1 U12433 ( .A(n10509), .B(n13374), .ZN(n15967) );
  XNOR2_X1 U12434 ( .A(n10510), .B(n13374), .ZN(n10512) );
  AOI21_X1 U12435 ( .B1(n10512), .B2(n14393), .A(n10511), .ZN(n15964) );
  MUX2_X1 U12436 ( .A(n10513), .B(n15964), .S(n14427), .Z(n10522) );
  AOI211_X1 U12437 ( .C1(n13145), .C2(n10836), .A(n14416), .B(n10514), .ZN(
        n15963) );
  INV_X1 U12438 ( .A(n10515), .ZN(n10516) );
  INV_X1 U12439 ( .A(n10517), .ZN(n10518) );
  INV_X1 U12440 ( .A(n13145), .ZN(n15966) );
  OAI22_X1 U12441 ( .A1(n14366), .A2(n15966), .B1(n10519), .B2(n14430), .ZN(
        n10520) );
  AOI21_X1 U12442 ( .B1(n15963), .B2(n14438), .A(n10520), .ZN(n10521) );
  OAI211_X1 U12443 ( .C1(n14303), .C2(n15967), .A(n10522), .B(n10521), .ZN(
        P2_U3261) );
  AOI21_X1 U12444 ( .B1(n10525), .B2(n10524), .A(n10523), .ZN(n10526) );
  MUX2_X1 U12445 ( .A(n10527), .B(n10526), .S(n15899), .Z(n10531) );
  OR2_X1 U12446 ( .A1(n10528), .A2(n12623), .ZN(n11698) );
  INV_X1 U12447 ( .A(n11698), .ZN(n15898) );
  AOI22_X1 U12448 ( .A1(n10529), .A2(n13792), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n13829), .ZN(n10530) );
  NAND2_X1 U12449 ( .A1(n10531), .A2(n10530), .ZN(P3_U3232) );
  INV_X1 U12450 ( .A(n13075), .ZN(n10532) );
  NAND2_X1 U12451 ( .A1(n10533), .A2(n10532), .ZN(n10535) );
  INV_X1 U12452 ( .A(n10538), .ZN(n11009) );
  XNOR2_X1 U12453 ( .A(n10539), .B(n13029), .ZN(n15959) );
  INV_X1 U12454 ( .A(n15959), .ZN(n10550) );
  NAND2_X1 U12455 ( .A1(n10540), .A2(n13017), .ZN(n10541) );
  NOR2_X2 U12456 ( .A1(n15998), .A2(n10541), .ZN(n15990) );
  AND2_X1 U12457 ( .A1(n10621), .A2(n15949), .ZN(n10542) );
  OR2_X1 U12458 ( .A1(n10542), .A2(n10677), .ZN(n15953) );
  NAND2_X1 U12459 ( .A1(n16037), .A2(n10543), .ZN(n10544) );
  OAI211_X1 U12460 ( .C1(n15953), .C2(n14952), .A(n15951), .B(n10544), .ZN(
        n10545) );
  MUX2_X1 U12461 ( .A(n10545), .B(P1_REG2_REG_4__SCAN_IN), .S(n15998), .Z(
        n10548) );
  NOR2_X1 U12462 ( .A1(n16047), .A2(n16060), .ZN(n14910) );
  NAND2_X1 U12463 ( .A1(n10546), .A2(n13029), .ZN(n15954) );
  AND3_X1 U12464 ( .A1(n15956), .A2(n14910), .A3(n15954), .ZN(n10547) );
  AOI211_X1 U12465 ( .C1(n15990), .C2(n15949), .A(n10548), .B(n10547), .ZN(
        n10549) );
  OAI21_X1 U12466 ( .B1(n14967), .B2(n10550), .A(n10549), .ZN(P1_U3289) );
  AOI22_X1 U12467 ( .A1(n10551), .A2(n12234), .B1(n13330), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n10552) );
  NAND2_X2 U12468 ( .A1(n10553), .A2(n10552), .ZN(n14435) );
  INV_X1 U12469 ( .A(n14191), .ZN(n10857) );
  OR2_X1 U12470 ( .A1(n13170), .A2(n14194), .ZN(n10554) );
  NAND2_X1 U12471 ( .A1(n10555), .A2(n10554), .ZN(n10965) );
  NAND2_X1 U12472 ( .A1(n13177), .A2(n14193), .ZN(n10557) );
  OR2_X1 U12473 ( .A1(n13177), .A2(n14193), .ZN(n10556) );
  AND2_X1 U12474 ( .A1(n10557), .A2(n10556), .ZN(n13379) );
  INV_X1 U12475 ( .A(n13379), .ZN(n10969) );
  XOR2_X1 U12476 ( .A(n13380), .B(n10686), .Z(n14437) );
  AOI21_X1 U12477 ( .B1(n14435), .B2(n10966), .A(n14416), .ZN(n10558) );
  AND2_X1 U12478 ( .A1(n10558), .A2(n10787), .ZN(n14439) );
  OR2_X1 U12479 ( .A1(n13170), .A2(n10561), .ZN(n10559) );
  NAND2_X1 U12480 ( .A1(n13170), .A2(n10561), .ZN(n10562) );
  INV_X1 U12481 ( .A(n14193), .ZN(n13179) );
  OR2_X1 U12482 ( .A1(n13177), .A2(n13179), .ZN(n10563) );
  NAND2_X1 U12483 ( .A1(n13177), .A2(n13179), .ZN(n10564) );
  INV_X1 U12484 ( .A(n10717), .ZN(n10566) );
  AOI211_X1 U12485 ( .C1(n13380), .C2(n10567), .A(n14413), .B(n10566), .ZN(
        n10575) );
  NAND2_X1 U12486 ( .A1(n13322), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10572) );
  XNOR2_X1 U12487 ( .A(n10696), .B(P2_REG3_REG_10__SCAN_IN), .ZN(n10851) );
  NAND2_X1 U12488 ( .A1(n12342), .A2(n10851), .ZN(n10571) );
  OR2_X1 U12489 ( .A1(n12239), .A2(n10786), .ZN(n10570) );
  INV_X1 U12490 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10568) );
  OR2_X1 U12491 ( .A1(n13325), .A2(n10568), .ZN(n10569) );
  NAND4_X1 U12492 ( .A1(n10572), .A2(n10571), .A3(n10570), .A4(n10569), .ZN(
        n14190) );
  NAND2_X1 U12493 ( .A1(n14190), .A2(n14139), .ZN(n10574) );
  NAND2_X1 U12494 ( .A1(n14193), .A2(n14137), .ZN(n10573) );
  NAND2_X1 U12495 ( .A1(n10574), .A2(n10573), .ZN(n12403) );
  OR2_X1 U12496 ( .A1(n10575), .A2(n12403), .ZN(n14428) );
  AOI211_X1 U12497 ( .C1(n16140), .C2(n14437), .A(n14439), .B(n14428), .ZN(
        n10579) );
  AOI22_X1 U12498 ( .A1(n14435), .A2(n14524), .B1(n16141), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n10576) );
  OAI21_X1 U12499 ( .B1(n10579), .B2(n16141), .A(n10576), .ZN(P2_U3508) );
  OAI22_X1 U12500 ( .A1(n7372), .A2(n14566), .B1(n16146), .B2(n10455), .ZN(
        n10577) );
  INV_X1 U12501 ( .A(n10577), .ZN(n10578) );
  OAI21_X1 U12502 ( .B1(n10579), .B2(n16143), .A(n10578), .ZN(P2_U3457) );
  INV_X1 U12503 ( .A(n10580), .ZN(n10589) );
  NAND2_X1 U12504 ( .A1(n14427), .A2(n13100), .ZN(n14425) );
  MUX2_X1 U12505 ( .A(n10581), .B(P2_REG2_REG_7__SCAN_IN), .S(n14378), .Z(
        n10582) );
  INV_X1 U12506 ( .A(n10582), .ZN(n10588) );
  OAI22_X1 U12507 ( .A1(n10584), .A2(n14366), .B1(n14430), .B2(n10583), .ZN(
        n10585) );
  AOI21_X1 U12508 ( .B1(n10586), .B2(n14438), .A(n10585), .ZN(n10587) );
  OAI211_X1 U12509 ( .C1(n10589), .C2(n14425), .A(n10588), .B(n10587), .ZN(
        P2_U3258) );
  OAI21_X1 U12510 ( .B1(n10590), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n10979) );
  XNOR2_X1 U12511 ( .A(n10979), .B(P2_IR_REG_15__SCAN_IN), .ZN(n11770) );
  INV_X1 U12512 ( .A(n11770), .ZN(n15442) );
  OAI222_X1 U12513 ( .A1(n14588), .A2(n10592), .B1(n14593), .B2(n10591), .C1(
        n15442), .C2(P2_U3088), .ZN(P2_U3312) );
  INV_X1 U12514 ( .A(n10593), .ZN(n10595) );
  AND2_X1 U12515 ( .A1(n12518), .A2(n14746), .ZN(n10597) );
  AOI21_X1 U12516 ( .B1(n12844), .B2(n12519), .A(n10597), .ZN(n10815) );
  AOI22_X1 U12517 ( .A1(n12844), .A2(n7181), .B1(n12519), .B2(n14746), .ZN(
        n10598) );
  XNOR2_X1 U12518 ( .A(n10598), .B(n12526), .ZN(n10814) );
  XOR2_X1 U12519 ( .A(n10815), .B(n10814), .Z(n10599) );
  OAI211_X1 U12520 ( .C1(n10600), .C2(n10599), .A(n10819), .B(n14719), .ZN(
        n10605) );
  INV_X1 U12521 ( .A(n14745), .ZN(n10921) );
  NAND2_X1 U12522 ( .A1(n15927), .A2(n14980), .ZN(n16115) );
  NOR2_X1 U12523 ( .A1(n14725), .A2(n15003), .ZN(n14713) );
  NAND2_X1 U12524 ( .A1(n14713), .A2(n14747), .ZN(n10602) );
  OAI211_X1 U12525 ( .C1(n10921), .C2(n16115), .A(n10602), .B(n10601), .ZN(
        n10603) );
  AOI21_X1 U12526 ( .B1(n10644), .B2(n14728), .A(n10603), .ZN(n10604) );
  OAI211_X1 U12527 ( .C1(n7595), .C2(n14731), .A(n10605), .B(n10604), .ZN(
        P1_U3213) );
  INV_X1 U12528 ( .A(n10606), .ZN(n10607) );
  OAI222_X1 U12529 ( .A1(P3_U3151), .A2(n12596), .B1(n13082), .B2(n10607), 
        .C1(n11223), .C2(n13083), .ZN(P3_U3275) );
  AOI21_X1 U12530 ( .B1(n11413), .B2(P1_REG2_REG_13__SCAN_IN), .A(n10608), 
        .ZN(n10802) );
  XNOR2_X1 U12531 ( .A(n11409), .B(P1_REG2_REG_14__SCAN_IN), .ZN(n10801) );
  XNOR2_X1 U12532 ( .A(n10802), .B(n10801), .ZN(n10617) );
  AOI22_X1 U12533 ( .A1(n14787), .A2(n11409), .B1(n14797), .B2(
        P1_ADDR_REG_14__SCAN_IN), .ZN(n10616) );
  NAND2_X1 U12534 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n16130)
         );
  INV_X1 U12535 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10609) );
  XNOR2_X1 U12536 ( .A(n11409), .B(n10609), .ZN(n10804) );
  OAI21_X1 U12537 ( .B1(n10612), .B2(n10611), .A(n10610), .ZN(n10805) );
  XOR2_X1 U12538 ( .A(n10804), .B(n10805), .Z(n10613) );
  NAND2_X1 U12539 ( .A1(n10613), .A2(n14834), .ZN(n10614) );
  AND2_X1 U12540 ( .A1(n16130), .A2(n10614), .ZN(n10615) );
  OAI211_X1 U12541 ( .C1(n10617), .C2(n14829), .A(n10616), .B(n10615), .ZN(
        P1_U3257) );
  XNOR2_X1 U12542 ( .A(n10618), .B(n13027), .ZN(n15934) );
  XNOR2_X1 U12543 ( .A(n10619), .B(n13027), .ZN(n15937) );
  AOI21_X1 U12544 ( .B1(n10620), .B2(n15918), .A(n15952), .ZN(n10622) );
  NAND2_X1 U12545 ( .A1(n10622), .A2(n10621), .ZN(n15931) );
  INV_X1 U12546 ( .A(n12167), .ZN(n12550) );
  NAND2_X1 U12547 ( .A1(n12550), .A2(n14836), .ZN(n14997) );
  AOI22_X1 U12548 ( .A1(n15990), .A2(n15918), .B1(n16037), .B2(n10623), .ZN(
        n10629) );
  OR2_X1 U12549 ( .A1(n10624), .A2(n15003), .ZN(n10626) );
  NAND2_X1 U12550 ( .A1(n14749), .A2(n14980), .ZN(n10625) );
  NAND2_X1 U12551 ( .A1(n10626), .A2(n10625), .ZN(n15926) );
  INV_X1 U12552 ( .A(n15926), .ZN(n15932) );
  MUX2_X1 U12553 ( .A(n15932), .B(n10627), .S(n15998), .Z(n10628) );
  OAI211_X1 U12554 ( .C1(n15931), .C2(n14997), .A(n10629), .B(n10628), .ZN(
        n10630) );
  AOI21_X1 U12555 ( .B1(n14910), .B2(n15937), .A(n10630), .ZN(n10631) );
  OAI21_X1 U12556 ( .B1(n14967), .B2(n15934), .A(n10631), .ZN(P1_U3290) );
  OAI222_X1 U12557 ( .A1(n13082), .A2(n10632), .B1(n13083), .B2(n15183), .C1(
        P3_U3151), .C2(n12623), .ZN(P3_U3274) );
  OAI211_X1 U12558 ( .C1(n10635), .C2(n10634), .A(n10633), .B(n13527), .ZN(
        n10641) );
  OAI22_X1 U12559 ( .A1(n13519), .A2(n11113), .B1(n10636), .B2(n13548), .ZN(
        n10637) );
  AOI211_X1 U12560 ( .C1(n10639), .C2(n13511), .A(n10638), .B(n10637), .ZN(
        n10640) );
  OAI211_X1 U12561 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n13531), .A(n10641), .B(
        n10640), .ZN(P3_U3158) );
  NAND2_X1 U12562 ( .A1(n10642), .A2(n13059), .ZN(n13004) );
  INV_X1 U12563 ( .A(n13004), .ZN(n10643) );
  NAND2_X1 U12564 ( .A1(n11899), .A2(n10643), .ZN(n10755) );
  AOI22_X1 U12565 ( .A1(n15990), .A2(n12844), .B1(n10644), .B2(n16037), .ZN(
        n10645) );
  OAI21_X1 U12566 ( .B1(n10646), .B2(n14997), .A(n10645), .ZN(n10649) );
  MUX2_X1 U12567 ( .A(n10647), .B(P1_REG2_REG_7__SCAN_IN), .S(n16047), .Z(
        n10648) );
  AOI211_X1 U12568 ( .C1(n16044), .C2(n10650), .A(n10649), .B(n10648), .ZN(
        n10651) );
  INV_X1 U12569 ( .A(n10651), .ZN(P1_U3286) );
  NAND2_X1 U12570 ( .A1(n10664), .A2(n7190), .ZN(n15846) );
  INV_X1 U12571 ( .A(n9774), .ZN(n10661) );
  INV_X1 U12572 ( .A(n13106), .ZN(n10652) );
  AND2_X1 U12573 ( .A1(n10661), .A2(n10652), .ZN(n15848) );
  AOI21_X1 U12574 ( .B1(n14413), .B2(n16107), .A(n15848), .ZN(n10655) );
  INV_X1 U12575 ( .A(n10653), .ZN(n10654) );
  NOR2_X1 U12576 ( .A1(n10655), .A2(n10654), .ZN(n15847) );
  OAI21_X1 U12577 ( .B1(n13326), .B2(n15846), .A(n15847), .ZN(n10656) );
  INV_X1 U12578 ( .A(n14430), .ZN(n14376) );
  AOI22_X1 U12579 ( .A1(n10656), .A2(n14427), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n14376), .ZN(n10659) );
  INV_X1 U12580 ( .A(n14425), .ZN(n11746) );
  INV_X1 U12581 ( .A(n15848), .ZN(n10657) );
  NAND2_X1 U12582 ( .A1(n11746), .A2(n10657), .ZN(n10658) );
  OAI211_X1 U12583 ( .C1(n9619), .C2(n14427), .A(n10659), .B(n10658), .ZN(
        P2_U3265) );
  OAI21_X1 U12584 ( .B1(n10663), .B2(n14413), .A(n10662), .ZN(n15867) );
  MUX2_X1 U12585 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n15867), .S(n14427), .Z(
        n10668) );
  NAND2_X1 U12586 ( .A1(n10664), .A2(n13109), .ZN(n10665) );
  AND3_X1 U12587 ( .A1(n10870), .A2(n14397), .A3(n10665), .ZN(n15865) );
  AOI22_X1 U12588 ( .A1(n14438), .A2(n15865), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n14376), .ZN(n10666) );
  OAI21_X1 U12589 ( .B1(n15864), .B2(n14366), .A(n10666), .ZN(n10667) );
  AOI211_X1 U12590 ( .C1(n15862), .C2(n14436), .A(n10668), .B(n10667), .ZN(
        n10669) );
  INV_X1 U12591 ( .A(n10669), .ZN(P2_U3264) );
  NAND2_X1 U12592 ( .A1(n11899), .A2(n16034), .ZN(n10670) );
  NAND2_X1 U12593 ( .A1(n10755), .A2(n10670), .ZN(n12172) );
  INV_X1 U12594 ( .A(n12172), .ZN(n11254) );
  XNOR2_X1 U12595 ( .A(n10671), .B(n13031), .ZN(n15976) );
  OAI211_X1 U12596 ( .C1(n10673), .C2(n13031), .A(n10672), .B(n15955), .ZN(
        n10675) );
  NAND2_X1 U12597 ( .A1(n10675), .A2(n10674), .ZN(n15974) );
  INV_X1 U12598 ( .A(n15974), .ZN(n10676) );
  MUX2_X1 U12599 ( .A(n9148), .B(n10676), .S(n11899), .Z(n10685) );
  INV_X1 U12600 ( .A(n10677), .ZN(n10679) );
  AOI211_X1 U12601 ( .C1(n12832), .C2(n10679), .A(n15952), .B(n10678), .ZN(
        n15972) );
  INV_X1 U12602 ( .A(n10680), .ZN(n10681) );
  OAI22_X1 U12603 ( .A1(n16041), .A2(n10682), .B1(n10681), .B2(n15016), .ZN(
        n10683) );
  AOI21_X1 U12604 ( .B1(n16035), .B2(n15972), .A(n10683), .ZN(n10684) );
  OAI211_X1 U12605 ( .C1(n11254), .C2(n15976), .A(n10685), .B(n10684), .ZN(
        P1_U3288) );
  AOI22_X1 U12606 ( .A1(n10687), .A2(n12234), .B1(n13330), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n10688) );
  AND2_X1 U12607 ( .A1(n13190), .A2(n14190), .ZN(n10690) );
  OAI22_X1 U12608 ( .A1(n10784), .A2(n10690), .B1(n14190), .B2(n13190), .ZN(
        n10704) );
  AOI22_X1 U12609 ( .A1(n10691), .A2(n12234), .B1(n13330), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n10692) );
  NAND2_X1 U12610 ( .A1(n13322), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10703) );
  INV_X1 U12611 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10695) );
  OAI21_X1 U12612 ( .B1(n10696), .B2(n10695), .A(n10694), .ZN(n10697) );
  AND2_X1 U12613 ( .A1(n10697), .A2(n10707), .ZN(n11276) );
  NAND2_X1 U12614 ( .A1(n12342), .A2(n11276), .ZN(n10702) );
  OR2_X1 U12615 ( .A1(n12239), .A2(n10698), .ZN(n10701) );
  INV_X1 U12616 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10699) );
  OR2_X1 U12617 ( .A1(n13325), .A2(n10699), .ZN(n10700) );
  NAND4_X1 U12618 ( .A1(n10703), .A2(n10702), .A3(n10701), .A4(n10700), .ZN(
        n14189) );
  XNOR2_X1 U12619 ( .A(n13203), .B(n14189), .ZN(n13383) );
  OR2_X1 U12620 ( .A1(n10704), .A2(n13383), .ZN(n11136) );
  NAND2_X1 U12621 ( .A1(n10704), .A2(n13383), .ZN(n10705) );
  NAND2_X1 U12622 ( .A1(n11136), .A2(n10705), .ZN(n10723) );
  NAND2_X1 U12623 ( .A1(n13322), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10713) );
  INV_X1 U12624 ( .A(n10707), .ZN(n10706) );
  NAND2_X1 U12625 ( .A1(n10706), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n11145) );
  NAND2_X1 U12626 ( .A1(n10707), .A2(n11386), .ZN(n10708) );
  AND2_X1 U12627 ( .A1(n11145), .A2(n10708), .ZN(n11157) );
  NAND2_X1 U12628 ( .A1(n12342), .A2(n11157), .ZN(n10712) );
  INV_X1 U12629 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11158) );
  OR2_X1 U12630 ( .A1(n12239), .A2(n11158), .ZN(n10711) );
  INV_X1 U12631 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10709) );
  OR2_X1 U12632 ( .A1(n13325), .A2(n10709), .ZN(n10710) );
  NAND4_X1 U12633 ( .A1(n10713), .A2(n10712), .A3(n10711), .A4(n10710), .ZN(
        n14188) );
  NAND2_X1 U12634 ( .A1(n14188), .A2(n14139), .ZN(n10715) );
  NAND2_X1 U12635 ( .A1(n14190), .A2(n14137), .ZN(n10714) );
  AND2_X1 U12636 ( .A1(n10715), .A2(n10714), .ZN(n11273) );
  OR2_X1 U12637 ( .A1(n14435), .A2(n10857), .ZN(n10716) );
  INV_X1 U12638 ( .A(n14190), .ZN(n10783) );
  NAND2_X1 U12639 ( .A1(n13190), .A2(n10783), .ZN(n10719) );
  NOR2_X1 U12640 ( .A1(n13190), .A2(n10783), .ZN(n10718) );
  OAI21_X1 U12641 ( .B1(n10720), .B2(n13383), .A(n11153), .ZN(n10721) );
  NAND2_X1 U12642 ( .A1(n10721), .A2(n14393), .ZN(n10722) );
  OAI211_X1 U12643 ( .C1(n10723), .C2(n16107), .A(n11273), .B(n10722), .ZN(
        n16074) );
  INV_X1 U12644 ( .A(n16074), .ZN(n10728) );
  INV_X1 U12645 ( .A(n10723), .ZN(n16076) );
  INV_X1 U12646 ( .A(n13203), .ZN(n16073) );
  NAND2_X1 U12647 ( .A1(n16073), .A2(n10788), .ZN(n11159) );
  OAI211_X1 U12648 ( .C1(n16073), .C2(n10788), .A(n14397), .B(n11159), .ZN(
        n16072) );
  AOI22_X1 U12649 ( .A1(n14378), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11276), 
        .B2(n14376), .ZN(n10725) );
  NAND2_X1 U12650 ( .A1(n13203), .A2(n14434), .ZN(n10724) );
  OAI211_X1 U12651 ( .C1(n16072), .C2(n14420), .A(n10725), .B(n10724), .ZN(
        n10726) );
  AOI21_X1 U12652 ( .B1(n16076), .B2(n11746), .A(n10726), .ZN(n10727) );
  OAI21_X1 U12653 ( .B1(n10728), .B2(n14378), .A(n10727), .ZN(P2_U3254) );
  OR2_X1 U12654 ( .A1(n12844), .A2(n14746), .ZN(n10729) );
  NAND2_X1 U12655 ( .A1(n10731), .A2(n12089), .ZN(n10734) );
  AOI22_X1 U12656 ( .A1(n13011), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n12008), 
        .B2(n10732), .ZN(n10733) );
  NAND2_X1 U12657 ( .A1(n10734), .A2(n10733), .ZN(n12849) );
  XNOR2_X1 U12658 ( .A(n12849), .B(n10921), .ZN(n13036) );
  OAI21_X1 U12659 ( .B1(n10735), .B2(n13036), .A(n10905), .ZN(n16011) );
  NAND2_X1 U12660 ( .A1(n12987), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n10742) );
  INV_X1 U12661 ( .A(n10911), .ZN(n10913) );
  NAND2_X1 U12662 ( .A1(n10737), .A2(n10736), .ZN(n10738) );
  AND2_X1 U12663 ( .A1(n10913), .A2(n10738), .ZN(n16038) );
  NAND2_X1 U12664 ( .A1(n12095), .A2(n16038), .ZN(n10741) );
  NAND2_X1 U12665 ( .A1(n12988), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10740) );
  NAND2_X1 U12666 ( .A1(n12014), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10739) );
  NAND4_X1 U12667 ( .A1(n10742), .A2(n10741), .A3(n10740), .A4(n10739), .ZN(
        n14744) );
  AOI22_X1 U12668 ( .A1(n14978), .A2(n14746), .B1(n14744), .B2(n14980), .ZN(
        n10749) );
  INV_X1 U12669 ( .A(n14746), .ZN(n10745) );
  NAND2_X1 U12670 ( .A1(n12844), .A2(n10745), .ZN(n10743) );
  OR2_X1 U12671 ( .A1(n12844), .A2(n10745), .ZN(n10746) );
  XNOR2_X1 U12672 ( .A(n10920), .B(n13036), .ZN(n10747) );
  NAND2_X1 U12673 ( .A1(n10747), .A2(n15955), .ZN(n10748) );
  OAI211_X1 U12674 ( .C1(n16011), .C2(n15977), .A(n10749), .B(n10748), .ZN(
        n16014) );
  MUX2_X1 U12675 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n16014), .S(n11899), .Z(
        n10750) );
  INV_X1 U12676 ( .A(n10750), .ZN(n10754) );
  AOI211_X1 U12677 ( .C1(n12849), .C2(n10751), .A(n15952), .B(n7592), .ZN(
        n16012) );
  OAI22_X1 U12678 ( .A1(n16041), .A2(n7593), .B1(n15016), .B2(n10825), .ZN(
        n10752) );
  AOI21_X1 U12679 ( .B1(n16012), .B2(n16035), .A(n10752), .ZN(n10753) );
  OAI211_X1 U12680 ( .C1(n16011), .C2(n10755), .A(n10754), .B(n10753), .ZN(
        P1_U3285) );
  NAND2_X1 U12681 ( .A1(n10759), .A2(n10758), .ZN(n15668) );
  MUX2_X1 U12682 ( .A(n10761), .B(n10760), .S(n13664), .Z(n10762) );
  XNOR2_X1 U12683 ( .A(n10762), .B(n15672), .ZN(n15667) );
  OR2_X1 U12684 ( .A1(n15668), .A2(n15667), .ZN(n15670) );
  NAND2_X1 U12685 ( .A1(n10762), .A2(n15672), .ZN(n10763) );
  NAND2_X1 U12686 ( .A1(n15670), .A2(n10763), .ZN(n10765) );
  MUX2_X1 U12687 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n13664), .Z(n11314) );
  XNOR2_X1 U12688 ( .A(n11314), .B(n11315), .ZN(n10764) );
  NAND2_X1 U12689 ( .A1(n10765), .A2(n10764), .ZN(n11318) );
  OAI21_X1 U12690 ( .B1(n10765), .B2(n10764), .A(n11318), .ZN(n10781) );
  NOR2_X1 U12691 ( .A1(n15672), .A2(n10766), .ZN(n10767) );
  NOR2_X1 U12692 ( .A1(n10760), .A2(n15660), .ZN(n15659) );
  AOI22_X1 U12693 ( .A1(n11315), .A2(P3_REG1_REG_8__SCAN_IN), .B1(n8471), .B2(
        n11328), .ZN(n10768) );
  AOI21_X1 U12694 ( .B1(n10769), .B2(n10768), .A(n11327), .ZN(n10770) );
  NOR2_X1 U12695 ( .A1(n10770), .A2(n15822), .ZN(n10780) );
  NOR2_X1 U12696 ( .A1(n15672), .A2(n10773), .ZN(n10774) );
  AOI22_X1 U12697 ( .A1(n11315), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n8475), .B2(
        n11328), .ZN(n10775) );
  AOI21_X1 U12698 ( .B1(n7325), .B2(n10775), .A(n11308), .ZN(n10776) );
  OR2_X1 U12699 ( .A1(n10776), .A2(n15825), .ZN(n10778) );
  AND2_X1 U12700 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n11471) );
  AOI21_X1 U12701 ( .B1(n15771), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11471), .ZN(
        n10777) );
  OAI211_X1 U12702 ( .C1(n15773), .C2(n11328), .A(n10778), .B(n10777), .ZN(
        n10779) );
  AOI211_X1 U12703 ( .C1(n10781), .C2(n15775), .A(n10780), .B(n10779), .ZN(
        n10782) );
  INV_X1 U12704 ( .A(n10782), .ZN(P3_U3190) );
  XNOR2_X1 U12705 ( .A(n13190), .B(n10783), .ZN(n13382) );
  XNOR2_X1 U12706 ( .A(n10784), .B(n13382), .ZN(n16048) );
  INV_X1 U12707 ( .A(n10851), .ZN(n10785) );
  OAI22_X1 U12708 ( .A1(n14427), .A2(n10786), .B1(n10785), .B2(n14430), .ZN(
        n10792) );
  INV_X1 U12709 ( .A(n13190), .ZN(n16050) );
  INV_X1 U12710 ( .A(n10787), .ZN(n10790) );
  INV_X1 U12711 ( .A(n10788), .ZN(n10789) );
  OAI211_X1 U12712 ( .C1(n16050), .C2(n10790), .A(n10789), .B(n14397), .ZN(
        n16049) );
  NOR2_X1 U12713 ( .A1(n16049), .A2(n14420), .ZN(n10791) );
  AOI211_X1 U12714 ( .C1(n14434), .C2(n13190), .A(n10792), .B(n10791), .ZN(
        n10798) );
  XNOR2_X1 U12715 ( .A(n10793), .B(n13382), .ZN(n10795) );
  INV_X1 U12716 ( .A(n14189), .ZN(n11388) );
  OAI22_X1 U12717 ( .A1(n10857), .A2(n14354), .B1(n11388), .B2(n14356), .ZN(
        n10794) );
  AOI21_X1 U12718 ( .B1(n10795), .B2(n14393), .A(n10794), .ZN(n10796) );
  OAI21_X1 U12719 ( .B1(n16048), .B2(n16107), .A(n10796), .ZN(n16051) );
  NAND2_X1 U12720 ( .A1(n16051), .A2(n14427), .ZN(n10797) );
  OAI211_X1 U12721 ( .C1(n16048), .C2(n14425), .A(n10798), .B(n10797), .ZN(
        P2_U3255) );
  INV_X1 U12722 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10799) );
  OAI22_X1 U12723 ( .A1(n10802), .A2(n10801), .B1(n10800), .B2(n10799), .ZN(
        n11358) );
  XNOR2_X1 U12724 ( .A(n11358), .B(n11627), .ZN(n10803) );
  NOR2_X1 U12725 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n10803), .ZN(n11359) );
  AOI21_X1 U12726 ( .B1(n10803), .B2(P1_REG2_REG_15__SCAN_IN), .A(n11359), 
        .ZN(n10812) );
  AOI22_X1 U12727 ( .A1(n10805), .A2(n10804), .B1(n11409), .B2(
        P1_REG1_REG_14__SCAN_IN), .ZN(n11366) );
  XOR2_X1 U12728 ( .A(n11627), .B(n11366), .Z(n10806) );
  AND2_X1 U12729 ( .A1(n10806), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n10807) );
  NOR2_X1 U12730 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n10806), .ZN(n11364) );
  OAI21_X1 U12731 ( .B1(n10807), .B2(n11364), .A(n14834), .ZN(n10811) );
  INV_X1 U12732 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n14723) );
  NOR2_X1 U12733 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14723), .ZN(n10809) );
  INV_X1 U12734 ( .A(n11627), .ZN(n11365) );
  NOR2_X1 U12735 ( .A1(n14828), .A2(n11365), .ZN(n10808) );
  AOI211_X1 U12736 ( .C1(P1_ADDR_REG_15__SCAN_IN), .C2(n14797), .A(n10809), 
        .B(n10808), .ZN(n10810) );
  OAI211_X1 U12737 ( .C1(n10812), .C2(n14829), .A(n10811), .B(n10810), .ZN(
        P1_U3258) );
  AOI22_X1 U12738 ( .A1(n12849), .A2(n12514), .B1(n12519), .B2(n14745), .ZN(
        n10813) );
  XNOR2_X1 U12739 ( .A(n10813), .B(n12526), .ZN(n11121) );
  AOI22_X1 U12740 ( .A1(n12849), .A2(n12519), .B1(n12518), .B2(n14745), .ZN(
        n11122) );
  XNOR2_X1 U12741 ( .A(n11121), .B(n11122), .ZN(n10821) );
  INV_X1 U12742 ( .A(n10814), .ZN(n10817) );
  AOI21_X1 U12743 ( .B1(n10821), .B2(n10820), .A(n11120), .ZN(n10828) );
  INV_X1 U12744 ( .A(n14744), .ZN(n11015) );
  OAI21_X1 U12745 ( .B1(n16115), .B2(n11015), .A(n10822), .ZN(n10823) );
  AOI21_X1 U12746 ( .B1(n14713), .B2(n14746), .A(n10823), .ZN(n10824) );
  OAI21_X1 U12747 ( .B1(n10825), .B2(n16133), .A(n10824), .ZN(n10826) );
  AOI21_X1 U12748 ( .B1(n16129), .B2(n12849), .A(n10826), .ZN(n10827) );
  OAI21_X1 U12749 ( .B1(n10828), .B2(n16123), .A(n10827), .ZN(P1_U3221) );
  XNOR2_X1 U12750 ( .A(n10830), .B(n10829), .ZN(n10832) );
  AOI21_X1 U12751 ( .B1(n10832), .B2(n14393), .A(n10831), .ZN(n15943) );
  XNOR2_X1 U12752 ( .A(n10833), .B(n13371), .ZN(n15940) );
  AOI21_X1 U12753 ( .B1(n13127), .B2(n10834), .A(n14416), .ZN(n10835) );
  NAND2_X1 U12754 ( .A1(n10836), .A2(n10835), .ZN(n15942) );
  OAI22_X1 U12755 ( .A1(n14427), .A2(n9587), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n14430), .ZN(n10837) );
  AOI21_X1 U12756 ( .B1(n14434), .B2(n13127), .A(n10837), .ZN(n10838) );
  OAI21_X1 U12757 ( .B1(n14420), .B2(n15942), .A(n10838), .ZN(n10839) );
  AOI21_X1 U12758 ( .B1(n15940), .B2(n14436), .A(n10839), .ZN(n10840) );
  OAI21_X1 U12759 ( .B1(n14378), .B2(n15943), .A(n10840), .ZN(P2_U3262) );
  INV_X1 U12760 ( .A(n10841), .ZN(n10843) );
  OAI22_X1 U12761 ( .A1(n12792), .A2(P3_U3151), .B1(SI_22_), .B2(n13083), .ZN(
        n10842) );
  AOI21_X1 U12762 ( .B1(n10843), .B2(n16149), .A(n10842), .ZN(P3_U3273) );
  INV_X1 U12763 ( .A(n10844), .ZN(n10846) );
  XNOR2_X1 U12764 ( .A(n14435), .B(n14043), .ZN(n10848) );
  NAND2_X1 U12765 ( .A1(n14191), .A2(n14416), .ZN(n10849) );
  XNOR2_X1 U12766 ( .A(n10848), .B(n10849), .ZN(n12402) );
  INV_X1 U12767 ( .A(n10848), .ZN(n10858) );
  NAND2_X1 U12768 ( .A1(n10858), .A2(n10849), .ZN(n10850) );
  XNOR2_X1 U12769 ( .A(n13190), .B(n14032), .ZN(n11269) );
  NAND2_X1 U12770 ( .A1(n14190), .A2(n14416), .ZN(n11268) );
  XNOR2_X1 U12771 ( .A(n11269), .B(n11268), .ZN(n10860) );
  INV_X1 U12772 ( .A(n11267), .ZN(n10863) );
  NAND2_X1 U12773 ( .A1(n14165), .A2(n14137), .ZN(n14096) );
  NOR2_X1 U12774 ( .A1(n14096), .A2(n10857), .ZN(n10856) );
  NOR2_X1 U12775 ( .A1(n14144), .A2(n14356), .ZN(n14099) );
  INV_X1 U12776 ( .A(n14099), .ZN(n10854) );
  NAND2_X1 U12777 ( .A1(n14141), .A2(n10851), .ZN(n10852) );
  OAI211_X1 U12778 ( .C1(n10854), .C2(n11388), .A(n10853), .B(n10852), .ZN(
        n10855) );
  AOI211_X1 U12779 ( .C1(n13190), .C2(n14150), .A(n10856), .B(n10855), .ZN(
        n10862) );
  OAI22_X1 U12780 ( .A1(n10858), .A2(n14168), .B1(n10857), .B2(n14152), .ZN(
        n10859) );
  NAND3_X1 U12781 ( .A1(n12410), .A2(n10860), .A3(n10859), .ZN(n10861) );
  OAI211_X1 U12782 ( .C1(n10863), .C2(n14168), .A(n10862), .B(n10861), .ZN(
        P2_U3189) );
  XNOR2_X1 U12783 ( .A(n10864), .B(n13369), .ZN(n10866) );
  AOI21_X1 U12784 ( .B1(n10866), .B2(n14393), .A(n10865), .ZN(n15909) );
  XNOR2_X1 U12785 ( .A(n10868), .B(n10867), .ZN(n15906) );
  AOI211_X1 U12786 ( .C1(n15904), .C2(n10870), .A(n14416), .B(n10869), .ZN(
        n15903) );
  OAI22_X1 U12787 ( .A1(n14427), .A2(n9602), .B1(n10871), .B2(n14430), .ZN(
        n10872) );
  AOI21_X1 U12788 ( .B1(n14438), .B2(n15903), .A(n10872), .ZN(n10873) );
  OAI21_X1 U12789 ( .B1(n7678), .B2(n14366), .A(n10873), .ZN(n10874) );
  AOI21_X1 U12790 ( .B1(n15906), .B2(n14436), .A(n10874), .ZN(n10875) );
  OAI21_X1 U12791 ( .B1(n14378), .B2(n15909), .A(n10875), .ZN(P2_U3263) );
  XOR2_X1 U12792 ( .A(n10876), .B(n12600), .Z(n15913) );
  AOI22_X1 U12793 ( .A1(n15876), .A2(n13576), .B1(n13575), .B2(n15873), .ZN(
        n10882) );
  AND2_X1 U12794 ( .A1(n15877), .A2(n10877), .ZN(n10880) );
  OAI211_X1 U12795 ( .C1(n10880), .C2(n10879), .A(n15881), .B(n10878), .ZN(
        n10881) );
  OAI211_X1 U12796 ( .C1(n15913), .C2(n15886), .A(n10882), .B(n10881), .ZN(
        n15915) );
  NAND2_X1 U12797 ( .A1(n15915), .A2(n15899), .ZN(n10885) );
  OAI22_X1 U12798 ( .A1(n13882), .A2(n15912), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n15892), .ZN(n10883) );
  AOI21_X1 U12799 ( .B1(n13853), .B2(P3_REG2_REG_3__SCAN_IN), .A(n10883), .ZN(
        n10884) );
  OAI211_X1 U12800 ( .C1(n15913), .C2(n15402), .A(n10885), .B(n10884), .ZN(
        P3_U3230) );
  MUX2_X1 U12801 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n7178), .Z(n11087) );
  XNOR2_X1 U12802 ( .A(n11086), .B(n11087), .ZN(n11722) );
  INV_X1 U12803 ( .A(n11722), .ZN(n10984) );
  NAND2_X1 U12804 ( .A1(n10891), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10890) );
  MUX2_X1 U12805 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10890), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n10894) );
  INV_X1 U12806 ( .A(n10891), .ZN(n10893) );
  NAND2_X1 U12807 ( .A1(n10893), .A2(n10892), .ZN(n11093) );
  NAND2_X1 U12808 ( .A1(n10894), .A2(n11093), .ZN(n11646) );
  OAI222_X1 U12809 ( .A1(n15167), .A2(n10984), .B1(n11646), .B2(P1_U3086), 
        .C1(n10895), .C2(n15157), .ZN(P1_U3339) );
  MUX2_X1 U12810 ( .A(n10896), .B(P1_REG2_REG_2__SCAN_IN), .S(n16047), .Z(
        n10900) );
  AOI22_X1 U12811 ( .A1(n16035), .A2(n10897), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n16037), .ZN(n10898) );
  OAI21_X1 U12812 ( .B1(n16041), .B2(n12805), .A(n10898), .ZN(n10899) );
  AOI211_X1 U12813 ( .C1(n14910), .C2(n10901), .A(n10900), .B(n10899), .ZN(
        n10902) );
  OAI21_X1 U12814 ( .B1(n11254), .B2(n10903), .A(n10902), .ZN(P1_U3291) );
  NAND2_X1 U12815 ( .A1(n12849), .A2(n14745), .ZN(n10904) );
  NAND2_X1 U12816 ( .A1(n10906), .A2(n12089), .ZN(n10909) );
  AOI22_X1 U12817 ( .A1(n13011), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n12008), 
        .B2(n10907), .ZN(n10908) );
  NAND2_X2 U12818 ( .A1(n10909), .A2(n10908), .ZN(n12858) );
  XNOR2_X1 U12819 ( .A(n12858), .B(n14744), .ZN(n13037) );
  OAI21_X1 U12820 ( .B1(n10910), .B2(n10923), .A(n10996), .ZN(n16043) );
  INV_X1 U12821 ( .A(n16043), .ZN(n10928) );
  NAND2_X1 U12822 ( .A1(n12987), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10918) );
  NAND2_X1 U12823 ( .A1(n10911), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11002) );
  INV_X1 U12824 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10912) );
  NAND2_X1 U12825 ( .A1(n10913), .A2(n10912), .ZN(n10914) );
  AND2_X1 U12826 ( .A1(n11002), .A2(n10914), .ZN(n11304) );
  NAND2_X1 U12827 ( .A1(n12095), .A2(n11304), .ZN(n10917) );
  NAND2_X1 U12828 ( .A1(n12988), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10916) );
  NAND2_X1 U12829 ( .A1(n12014), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n10915) );
  NAND4_X1 U12830 ( .A1(n10918), .A2(n10917), .A3(n10916), .A4(n10915), .ZN(
        n14743) );
  INV_X1 U12831 ( .A(n13036), .ZN(n10919) );
  OR2_X1 U12832 ( .A1(n12849), .A2(n10921), .ZN(n10922) );
  XNOR2_X1 U12833 ( .A(n11010), .B(n10923), .ZN(n10924) );
  AOI222_X1 U12834 ( .A1(n14745), .A2(n14978), .B1(n14743), .B2(n14980), .C1(
        n15955), .C2(n10924), .ZN(n16032) );
  INV_X1 U12835 ( .A(n11008), .ZN(n10925) );
  AOI211_X1 U12836 ( .C1(n12858), .C2(n10926), .A(n15952), .B(n10925), .ZN(
        n16036) );
  AOI21_X1 U12837 ( .B1(n15948), .B2(n12858), .A(n16036), .ZN(n10927) );
  OAI211_X1 U12838 ( .C1(n15933), .C2(n10928), .A(n16032), .B(n10927), .ZN(
        n10930) );
  NAND2_X1 U12839 ( .A1(n10930), .A2(n16067), .ZN(n10929) );
  OAI21_X1 U12840 ( .B1(n16067), .B2(n9262), .A(n10929), .ZN(P1_U3537) );
  INV_X1 U12841 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10932) );
  NAND2_X1 U12842 ( .A1(n10930), .A2(n16071), .ZN(n10931) );
  OAI21_X1 U12843 ( .B1(n16071), .B2(n10932), .A(n10931), .ZN(P1_U3486) );
  INV_X1 U12844 ( .A(n10933), .ZN(n10934) );
  XNOR2_X1 U12845 ( .A(n10934), .B(n13028), .ZN(n15855) );
  NAND2_X1 U12846 ( .A1(n10936), .A2(n10935), .ZN(n10937) );
  NAND2_X1 U12847 ( .A1(n10937), .A2(n15041), .ZN(n10939) );
  OR2_X1 U12848 ( .A1(n10939), .A2(n10938), .ZN(n15852) );
  INV_X1 U12849 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10940) );
  OAI22_X1 U12850 ( .A1(n14997), .A2(n15852), .B1(n10940), .B2(n15016), .ZN(
        n10944) );
  XNOR2_X1 U12851 ( .A(n13028), .B(n12814), .ZN(n10942) );
  AOI21_X1 U12852 ( .B1(n10942), .B2(n15955), .A(n10941), .ZN(n15853) );
  OAI22_X1 U12853 ( .A1(n16041), .A2(n15854), .B1(n16047), .B2(n15853), .ZN(
        n10943) );
  AOI211_X1 U12854 ( .C1(P1_REG2_REG_1__SCAN_IN), .C2(n15998), .A(n10944), .B(
        n10943), .ZN(n10945) );
  OAI21_X1 U12855 ( .B1(n11254), .B2(n15855), .A(n10945), .ZN(P1_U3292) );
  AOI22_X1 U12856 ( .A1(n14434), .A2(n13153), .B1(n14376), .B2(n10946), .ZN(
        n10947) );
  OAI21_X1 U12857 ( .B1(n14420), .B2(n10948), .A(n10947), .ZN(n10951) );
  MUX2_X1 U12858 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10949), .S(n14427), .Z(
        n10950) );
  AOI211_X1 U12859 ( .C1(n14436), .C2(n10952), .A(n10951), .B(n10950), .ZN(
        n10953) );
  INV_X1 U12860 ( .A(n10953), .ZN(P2_U3260) );
  INV_X1 U12861 ( .A(n10954), .ZN(n10957) );
  AOI22_X1 U12862 ( .A1(n14434), .A2(n13161), .B1(n10955), .B2(n14376), .ZN(
        n10956) );
  OAI21_X1 U12863 ( .B1(n10957), .B2(n14420), .A(n10956), .ZN(n10960) );
  MUX2_X1 U12864 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10958), .S(n14427), .Z(
        n10959) );
  AOI211_X1 U12865 ( .C1(n14436), .C2(n10961), .A(n10960), .B(n10959), .ZN(
        n10962) );
  INV_X1 U12866 ( .A(n10962), .ZN(P2_U3259) );
  INV_X1 U12867 ( .A(n10963), .ZN(n10964) );
  AOI21_X1 U12868 ( .B1(n10969), .B2(n10965), .A(n10964), .ZN(n16024) );
  OAI211_X1 U12869 ( .C1(n7681), .C2(n7682), .A(n14397), .B(n10966), .ZN(
        n16021) );
  AOI22_X1 U12870 ( .A1(n13177), .A2(n14434), .B1(n10967), .B2(n14376), .ZN(
        n10968) );
  OAI21_X1 U12871 ( .B1(n16021), .B2(n14420), .A(n10968), .ZN(n10976) );
  XNOR2_X1 U12872 ( .A(n10970), .B(n10969), .ZN(n10971) );
  NAND2_X1 U12873 ( .A1(n10971), .A2(n14393), .ZN(n10974) );
  INV_X1 U12874 ( .A(n10972), .ZN(n10973) );
  NAND2_X1 U12875 ( .A1(n10974), .A2(n10973), .ZN(n16023) );
  MUX2_X1 U12876 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n16023), .S(n14427), .Z(
        n10975) );
  AOI211_X1 U12877 ( .C1(n14436), .C2(n16024), .A(n10976), .B(n10975), .ZN(
        n10977) );
  INV_X1 U12878 ( .A(n10977), .ZN(P2_U3257) );
  INV_X1 U12879 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10985) );
  INV_X1 U12880 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n10978) );
  NAND2_X1 U12881 ( .A1(n10979), .A2(n10978), .ZN(n10980) );
  NAND2_X1 U12882 ( .A1(n10980), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10982) );
  INV_X1 U12883 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n10981) );
  NAND2_X1 U12884 ( .A1(n10982), .A2(n10981), .ZN(n11097) );
  OR2_X1 U12885 ( .A1(n10982), .A2(n10981), .ZN(n10983) );
  INV_X1 U12886 ( .A(n11767), .ZN(n15454) );
  OAI222_X1 U12887 ( .A1(n14588), .A2(n10985), .B1(n14593), .B2(n10984), .C1(
        n15454), .C2(P2_U3088), .ZN(P2_U3311) );
  AOI21_X1 U12888 ( .B1(n10987), .B2(n10986), .A(n7320), .ZN(n10994) );
  OAI22_X1 U12889 ( .A1(n13519), .A2(n11208), .B1(n10988), .B2(n13548), .ZN(
        n10989) );
  AOI211_X1 U12890 ( .C1(n11030), .C2(n13511), .A(n10990), .B(n10989), .ZN(
        n10993) );
  INV_X1 U12891 ( .A(n10991), .ZN(n11029) );
  NAND2_X1 U12892 ( .A1(n13550), .A2(n11029), .ZN(n10992) );
  OAI211_X1 U12893 ( .C1(n10994), .C2(n13539), .A(n10993), .B(n10992), .ZN(
        P3_U3170) );
  OR2_X1 U12894 ( .A1(n12858), .A2(n14744), .ZN(n10995) );
  NAND2_X1 U12895 ( .A1(n10997), .A2(n12089), .ZN(n11000) );
  AOI22_X1 U12896 ( .A1(n13011), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n12008), 
        .B2(n10998), .ZN(n10999) );
  XNOR2_X1 U12897 ( .A(n12864), .B(n14743), .ZN(n13038) );
  OAI21_X1 U12898 ( .B1(n11001), .B2(n11014), .A(n11040), .ZN(n11165) );
  NAND2_X1 U12899 ( .A1(n9339), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n11007) );
  NAND2_X1 U12900 ( .A1(n11002), .A2(n11482), .ZN(n11003) );
  AND2_X1 U12901 ( .A1(n11042), .A2(n11003), .ZN(n11485) );
  NAND2_X1 U12902 ( .A1(n12095), .A2(n11485), .ZN(n11006) );
  NAND2_X1 U12903 ( .A1(n12014), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n11005) );
  NAND2_X1 U12904 ( .A1(n12988), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11004) );
  NAND4_X1 U12905 ( .A1(n11007), .A2(n11006), .A3(n11005), .A4(n11004), .ZN(
        n14742) );
  INV_X1 U12906 ( .A(n14742), .ZN(n11476) );
  NOR2_X1 U12907 ( .A1(n11476), .A2(n15005), .ZN(n11167) );
  AOI211_X1 U12908 ( .C1(n12864), .C2(n11008), .A(n15952), .B(n11050), .ZN(
        n11169) );
  AOI211_X1 U12909 ( .C1(n11165), .C2(n11009), .A(n11167), .B(n11169), .ZN(
        n11020) );
  NAND2_X1 U12910 ( .A1(n12858), .A2(n11015), .ZN(n11011) );
  INV_X1 U12911 ( .A(n11034), .ZN(n11012) );
  AOI211_X1 U12912 ( .C1(n11014), .C2(n11013), .A(n16060), .B(n11012), .ZN(
        n11170) );
  NOR2_X1 U12913 ( .A1(n11015), .A2(n15003), .ZN(n11166) );
  OAI21_X1 U12914 ( .B1(n11170), .B2(n11166), .A(n11899), .ZN(n11019) );
  INV_X1 U12915 ( .A(n12864), .ZN(n11307) );
  AOI22_X1 U12916 ( .A1(n16047), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n11304), 
        .B2(n16037), .ZN(n11016) );
  OAI21_X1 U12917 ( .B1(n11307), .B2(n16041), .A(n11016), .ZN(n11017) );
  AOI21_X1 U12918 ( .B1(n11165), .B2(n16044), .A(n11017), .ZN(n11018) );
  OAI211_X1 U12919 ( .C1(n11020), .C2(n14997), .A(n11019), .B(n11018), .ZN(
        P1_U3283) );
  XNOR2_X1 U12920 ( .A(n11021), .B(n12659), .ZN(n11027) );
  INV_X1 U12921 ( .A(n11027), .ZN(n11057) );
  XNOR2_X1 U12922 ( .A(n11022), .B(n11023), .ZN(n11025) );
  AOI22_X1 U12923 ( .A1(n15874), .A2(n15876), .B1(n15873), .B2(n13574), .ZN(
        n11024) );
  OAI21_X1 U12924 ( .B1(n11025), .B2(n13874), .A(n11024), .ZN(n11026) );
  AOI21_X1 U12925 ( .B1(n11027), .B2(n13754), .A(n11026), .ZN(n11056) );
  MUX2_X1 U12926 ( .A(n11028), .B(n11056), .S(n15899), .Z(n11032) );
  AOI22_X1 U12927 ( .A1(n15399), .A2(n11030), .B1(n13829), .B2(n11029), .ZN(
        n11031) );
  OAI211_X1 U12928 ( .C1(n11057), .C2(n15402), .A(n11032), .B(n11031), .ZN(
        P3_U3229) );
  INV_X1 U12929 ( .A(n14743), .ZN(n11131) );
  OR2_X1 U12930 ( .A1(n12864), .A2(n11131), .ZN(n11033) );
  NAND2_X1 U12931 ( .A1(n11034), .A2(n11033), .ZN(n11233) );
  NAND2_X1 U12932 ( .A1(n11035), .A2(n12089), .ZN(n11038) );
  AOI22_X1 U12933 ( .A1(n13011), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n12008), 
        .B2(n11036), .ZN(n11037) );
  OR2_X1 U12934 ( .A1(n12869), .A2(n14742), .ZN(n11227) );
  NAND2_X1 U12935 ( .A1(n12869), .A2(n14742), .ZN(n11225) );
  NAND2_X1 U12936 ( .A1(n11227), .A2(n11225), .ZN(n13040) );
  XNOR2_X1 U12937 ( .A(n11233), .B(n13040), .ZN(n16061) );
  INV_X1 U12938 ( .A(n14910), .ZN(n15001) );
  OR2_X1 U12939 ( .A1(n12864), .A2(n14743), .ZN(n11039) );
  NAND2_X1 U12940 ( .A1(n11040), .A2(n11039), .ZN(n11226) );
  XOR2_X1 U12941 ( .A(n13040), .B(n11226), .Z(n16065) );
  INV_X1 U12942 ( .A(n14967), .ZN(n14999) );
  NAND2_X1 U12943 ( .A1(n16065), .A2(n14999), .ZN(n11054) );
  NAND2_X1 U12944 ( .A1(n12987), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11047) );
  INV_X1 U12945 ( .A(n11236), .ZN(n11238) );
  NAND2_X1 U12946 ( .A1(n11042), .A2(n11041), .ZN(n11043) );
  AND2_X1 U12947 ( .A1(n11238), .A2(n11043), .ZN(n11824) );
  NAND2_X1 U12948 ( .A1(n12095), .A2(n11824), .ZN(n11046) );
  NAND2_X1 U12949 ( .A1(n12988), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11045) );
  NAND2_X1 U12950 ( .A1(n12014), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n11044) );
  NAND4_X1 U12951 ( .A1(n11047), .A2(n11046), .A3(n11045), .A4(n11044), .ZN(
        n14741) );
  AOI22_X1 U12952 ( .A1(n14978), .A2(n14743), .B1(n14741), .B2(n14980), .ZN(
        n16056) );
  INV_X1 U12953 ( .A(n16056), .ZN(n11048) );
  AOI22_X1 U12954 ( .A1(n11899), .A2(n11048), .B1(n11485), .B2(n16037), .ZN(
        n11049) );
  OAI21_X1 U12955 ( .B1(n9406), .B2(n11899), .A(n11049), .ZN(n11052) );
  NAND2_X1 U12956 ( .A1(n16059), .A2(n11050), .ZN(n11247) );
  OAI211_X1 U12957 ( .C1(n16059), .C2(n11050), .A(n15041), .B(n11247), .ZN(
        n16057) );
  NOR2_X1 U12958 ( .A1(n16057), .A2(n14997), .ZN(n11051) );
  AOI211_X1 U12959 ( .C1(n15990), .C2(n12869), .A(n11052), .B(n11051), .ZN(
        n11053) );
  OAI211_X1 U12960 ( .C1(n16061), .C2(n15001), .A(n11054), .B(n11053), .ZN(
        P1_U3282) );
  NAND2_X1 U12961 ( .A1(n13577), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n11055) );
  OAI21_X1 U12962 ( .B1(n13681), .B2(n13577), .A(n11055), .ZN(P3_U3520) );
  OAI21_X1 U12963 ( .B1(n16097), .B2(n11057), .A(n11056), .ZN(n11063) );
  INV_X1 U12964 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n11058) );
  OAI22_X1 U12965 ( .A1(n16159), .A2(n11061), .B1(n16104), .B2(n11058), .ZN(
        n11059) );
  AOI21_X1 U12966 ( .B1(n11063), .B2(n16104), .A(n11059), .ZN(n11060) );
  INV_X1 U12967 ( .A(n11060), .ZN(P3_U3402) );
  OAI22_X1 U12968 ( .A1(n16154), .A2(n11061), .B1(n16101), .B2(n10147), .ZN(
        n11062) );
  AOI21_X1 U12969 ( .B1(n11063), .B2(n16101), .A(n11062), .ZN(n11064) );
  INV_X1 U12970 ( .A(n11064), .ZN(P3_U3463) );
  MUX2_X1 U12971 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n7178), .Z(n11068) );
  NAND2_X1 U12972 ( .A1(n11068), .A2(SI_17_), .ZN(n11091) );
  OAI21_X1 U12973 ( .B1(n11067), .B2(n15207), .A(n11091), .ZN(n11065) );
  INV_X1 U12974 ( .A(n11065), .ZN(n11066) );
  NAND3_X1 U12975 ( .A1(n11091), .A2(n15207), .A3(n11067), .ZN(n11070) );
  INV_X1 U12976 ( .A(n11068), .ZN(n11069) );
  NAND2_X1 U12977 ( .A1(n11069), .A2(n15205), .ZN(n11090) );
  XNOR2_X1 U12978 ( .A(n11216), .B(n15184), .ZN(n11255) );
  MUX2_X1 U12979 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7178), .Z(n11256) );
  XNOR2_X1 U12980 ( .A(n11255), .B(n11256), .ZN(n12228) );
  INV_X1 U12981 ( .A(n12228), .ZN(n11107) );
  OAI21_X1 U12982 ( .B1(n11093), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n11073) );
  XNOR2_X1 U12983 ( .A(n11073), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14824) );
  AOI22_X1 U12984 ( .A1(n14824), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n15164), .ZN(n11074) );
  OAI21_X1 U12985 ( .B1(n11107), .B2(n15167), .A(n11074), .ZN(P1_U3337) );
  XNOR2_X1 U12986 ( .A(n11076), .B(n8117), .ZN(n11081) );
  OAI21_X1 U12987 ( .B1(n7322), .B2(n8117), .A(n11077), .ZN(n11079) );
  OAI22_X1 U12988 ( .A1(n11113), .A2(n15392), .B1(n11596), .B2(n15390), .ZN(
        n11078) );
  AOI21_X1 U12989 ( .B1(n11079), .B2(n15881), .A(n11078), .ZN(n11080) );
  OAI21_X1 U12990 ( .B1(n15886), .B2(n11081), .A(n11080), .ZN(n11101) );
  INV_X1 U12991 ( .A(n11101), .ZN(n11085) );
  INV_X1 U12992 ( .A(n11081), .ZN(n11102) );
  NOR2_X1 U12993 ( .A1(n15899), .A2(n8442), .ZN(n11083) );
  OAI22_X1 U12994 ( .A1(n13882), .A2(n12665), .B1(n11119), .B2(n15892), .ZN(
        n11082) );
  AOI211_X1 U12995 ( .C1(n11102), .C2(n13792), .A(n11083), .B(n11082), .ZN(
        n11084) );
  OAI21_X1 U12996 ( .B1(n11085), .B2(n13853), .A(n11084), .ZN(P3_U3228) );
  OR2_X1 U12997 ( .A1(n11088), .A2(n15207), .ZN(n11089) );
  NAND2_X1 U12998 ( .A1(n11091), .A2(n11090), .ZN(n11092) );
  INV_X1 U12999 ( .A(n11880), .ZN(n11100) );
  NAND2_X1 U13000 ( .A1(n11093), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n11095) );
  XNOR2_X1 U13001 ( .A(n11095), .B(n11094), .ZN(n11910) );
  OAI222_X1 U13002 ( .A1(n15157), .A2(n11096), .B1(n15167), .B2(n11100), .C1(
        P1_U3086), .C2(n11910), .ZN(P1_U3338) );
  INV_X1 U13003 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11784) );
  NAND2_X1 U13004 ( .A1(n11097), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n11099) );
  INV_X1 U13005 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n11098) );
  XNOR2_X1 U13006 ( .A(n11099), .B(n11098), .ZN(n15467) );
  OAI222_X1 U13007 ( .A1(n14588), .A2(n11784), .B1(n14593), .B2(n11100), .C1(
        P2_U3088), .C2(n15467), .ZN(P2_U3310) );
  AOI21_X1 U13008 ( .B1(n16082), .B2(n11102), .A(n11101), .ZN(n11279) );
  INV_X1 U13009 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n11103) );
  OAI22_X1 U13010 ( .A1(n16159), .A2(n12665), .B1(n16104), .B2(n11103), .ZN(
        n11104) );
  INV_X1 U13011 ( .A(n11104), .ZN(n11105) );
  OAI21_X1 U13012 ( .B1(n11279), .B2(n16160), .A(n11105), .ZN(P3_U3405) );
  INV_X1 U13013 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11108) );
  XNOR2_X1 U13014 ( .A(n11106), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14214) );
  INV_X1 U13015 ( .A(n14214), .ZN(n11764) );
  OAI222_X1 U13016 ( .A1(n14588), .A2(n11108), .B1(n14593), .B2(n11107), .C1(
        n11764), .C2(P2_U3088), .ZN(P2_U3309) );
  INV_X1 U13017 ( .A(n11204), .ZN(n11112) );
  NOR3_X1 U13018 ( .A1(n7320), .A2(n11110), .A3(n11109), .ZN(n11111) );
  OAI21_X1 U13019 ( .B1(n11112), .B2(n11111), .A(n13527), .ZN(n11118) );
  OAI22_X1 U13020 ( .A1(n13519), .A2(n11596), .B1(n11113), .B2(n13548), .ZN(
        n11114) );
  AOI211_X1 U13021 ( .C1(n11116), .C2(n13511), .A(n11115), .B(n11114), .ZN(
        n11117) );
  OAI211_X1 U13022 ( .C1(n11119), .C2(n13531), .A(n11118), .B(n11117), .ZN(
        P3_U3167) );
  NAND2_X1 U13023 ( .A1(n12858), .A2(n7181), .ZN(n11124) );
  NAND2_X1 U13024 ( .A1(n14744), .A2(n12519), .ZN(n11123) );
  NAND2_X1 U13025 ( .A1(n11124), .A2(n11123), .ZN(n11125) );
  XNOR2_X1 U13026 ( .A(n11125), .B(n12526), .ZN(n11294) );
  AND2_X1 U13027 ( .A1(n12518), .A2(n14744), .ZN(n11126) );
  AOI21_X1 U13028 ( .B1(n12858), .B2(n12519), .A(n11126), .ZN(n11296) );
  XNOR2_X1 U13029 ( .A(n11294), .B(n11296), .ZN(n11127) );
  OAI211_X1 U13030 ( .C1(n11128), .C2(n11127), .A(n11295), .B(n14719), .ZN(
        n11134) );
  NAND2_X1 U13031 ( .A1(n14713), .A2(n14745), .ZN(n11130) );
  OAI211_X1 U13032 ( .C1(n11131), .C2(n16115), .A(n11130), .B(n11129), .ZN(
        n11132) );
  AOI21_X1 U13033 ( .B1(n16038), .B2(n14728), .A(n11132), .ZN(n11133) );
  OAI211_X1 U13034 ( .C1(n7591), .C2(n14731), .A(n11134), .B(n11133), .ZN(
        P1_U3231) );
  NAND2_X1 U13035 ( .A1(n13203), .A2(n14189), .ZN(n11135) );
  NAND2_X1 U13036 ( .A1(n11136), .A2(n11135), .ZN(n11142) );
  AOI22_X1 U13037 ( .A1(n13330), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n12234), 
        .B2(n11137), .ZN(n11138) );
  NAND2_X2 U13038 ( .A1(n11139), .A2(n11138), .ZN(n13208) );
  NAND2_X1 U13039 ( .A1(n13208), .A2(n14188), .ZN(n11183) );
  OR2_X1 U13040 ( .A1(n13208), .A2(n14188), .ZN(n11140) );
  NAND2_X1 U13041 ( .A1(n11183), .A2(n11140), .ZN(n13384) );
  INV_X1 U13042 ( .A(n13384), .ZN(n11141) );
  NAND2_X1 U13043 ( .A1(n11142), .A2(n11141), .ZN(n11184) );
  OR2_X1 U13044 ( .A1(n11142), .A2(n11141), .ZN(n11143) );
  NAND2_X1 U13045 ( .A1(n11184), .A2(n11143), .ZN(n16086) );
  NAND2_X1 U13046 ( .A1(n13322), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11151) );
  INV_X1 U13047 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11144) );
  NAND2_X1 U13048 ( .A1(n11145), .A2(n11144), .ZN(n11146) );
  AND2_X1 U13049 ( .A1(n11192), .A2(n11146), .ZN(n11673) );
  NAND2_X1 U13050 ( .A1(n12342), .A2(n11673), .ZN(n11150) );
  OR2_X1 U13051 ( .A1(n12239), .A2(n10411), .ZN(n11149) );
  INV_X1 U13052 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11147) );
  OR2_X1 U13053 ( .A1(n13325), .A2(n11147), .ZN(n11148) );
  NAND4_X1 U13054 ( .A1(n11151), .A2(n11150), .A3(n11149), .A4(n11148), .ZN(
        n14187) );
  AOI22_X1 U13055 ( .A1(n14137), .A2(n14189), .B1(n14187), .B2(n14139), .ZN(
        n11156) );
  NAND2_X1 U13056 ( .A1(n13203), .A2(n11388), .ZN(n11152) );
  AND2_X1 U13057 ( .A1(n11153), .A2(n11152), .ZN(n11154) );
  OAI211_X1 U13058 ( .C1(n11154), .C2(n13384), .A(n11189), .B(n14393), .ZN(
        n11155) );
  OAI211_X1 U13059 ( .C1(n16086), .C2(n16107), .A(n11156), .B(n11155), .ZN(
        n16089) );
  NAND2_X1 U13060 ( .A1(n16089), .A2(n14427), .ZN(n11164) );
  INV_X1 U13061 ( .A(n11157), .ZN(n11387) );
  OAI22_X1 U13062 ( .A1(n14427), .A2(n11158), .B1(n11387), .B2(n14430), .ZN(
        n11162) );
  INV_X1 U13063 ( .A(n11159), .ZN(n11160) );
  INV_X1 U13064 ( .A(n13208), .ZN(n16088) );
  OAI211_X1 U13065 ( .C1(n11160), .C2(n16088), .A(n14397), .B(n11185), .ZN(
        n16087) );
  NOR2_X1 U13066 ( .A1(n16087), .A2(n14420), .ZN(n11161) );
  AOI211_X1 U13067 ( .C1(n14434), .C2(n13208), .A(n11162), .B(n11161), .ZN(
        n11163) );
  OAI211_X1 U13068 ( .C1(n16086), .C2(n14425), .A(n11164), .B(n11163), .ZN(
        P2_U3253) );
  INV_X1 U13069 ( .A(n11165), .ZN(n11172) );
  NOR2_X1 U13070 ( .A1(n11167), .A2(n11166), .ZN(n11302) );
  OAI21_X1 U13071 ( .B1(n11307), .B2(n16058), .A(n11302), .ZN(n11168) );
  NOR3_X1 U13072 ( .A1(n11170), .A2(n11169), .A3(n11168), .ZN(n11171) );
  OAI21_X1 U13073 ( .B1(n15933), .B2(n11172), .A(n11171), .ZN(n11175) );
  NAND2_X1 U13074 ( .A1(n11175), .A2(n16067), .ZN(n11173) );
  OAI21_X1 U13075 ( .B1(n16067), .B2(n11174), .A(n11173), .ZN(P1_U3538) );
  INV_X1 U13076 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n11177) );
  NAND2_X1 U13077 ( .A1(n11175), .A2(n16071), .ZN(n11176) );
  OAI21_X1 U13078 ( .B1(n16071), .B2(n11177), .A(n11176), .ZN(P1_U3489) );
  NAND2_X1 U13079 ( .A1(n11178), .A2(n16149), .ZN(n11179) );
  OAI211_X1 U13080 ( .C1(n15287), .C2(n13083), .A(n11179), .B(n12791), .ZN(
        P3_U3272) );
  AOI22_X1 U13081 ( .A1(n13330), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n11180), 
        .B2(n12234), .ZN(n11181) );
  NAND2_X2 U13082 ( .A1(n11182), .A2(n11181), .ZN(n13216) );
  XOR2_X1 U13083 ( .A(n13386), .B(n11510), .Z(n16105) );
  INV_X1 U13084 ( .A(n11506), .ZN(n11507) );
  AOI211_X1 U13085 ( .C1(n13216), .C2(n11185), .A(n14416), .B(n11507), .ZN(
        n16111) );
  INV_X1 U13086 ( .A(n13216), .ZN(n16108) );
  AOI22_X1 U13087 ( .A1(n14378), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11673), 
        .B2(n14376), .ZN(n11186) );
  OAI21_X1 U13088 ( .B1(n16108), .B2(n14366), .A(n11186), .ZN(n11187) );
  AOI21_X1 U13089 ( .B1(n16111), .B2(n14438), .A(n11187), .ZN(n11202) );
  INV_X1 U13090 ( .A(n14188), .ZN(n13210) );
  OR2_X1 U13091 ( .A1(n13208), .A2(n13210), .ZN(n11188) );
  XNOR2_X1 U13092 ( .A(n13386), .B(n11494), .ZN(n11200) );
  INV_X1 U13093 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n11191) );
  NAND2_X1 U13094 ( .A1(n11192), .A2(n11191), .ZN(n11193) );
  AND2_X1 U13095 ( .A1(n11497), .A2(n11193), .ZN(n11504) );
  NAND2_X1 U13096 ( .A1(n11504), .A2(n12342), .ZN(n11197) );
  NAND2_X1 U13097 ( .A1(n12345), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n11196) );
  NAND2_X1 U13098 ( .A1(n12336), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n11195) );
  OR2_X1 U13099 ( .A1(n12239), .A2(n11505), .ZN(n11194) );
  NAND4_X1 U13100 ( .A1(n11197), .A2(n11196), .A3(n11195), .A4(n11194), .ZN(
        n14186) );
  NAND2_X1 U13101 ( .A1(n14186), .A2(n14139), .ZN(n11199) );
  NAND2_X1 U13102 ( .A1(n14188), .A2(n14137), .ZN(n11198) );
  AND2_X1 U13103 ( .A1(n11199), .A2(n11198), .ZN(n11675) );
  OAI21_X1 U13104 ( .B1(n11200), .B2(n14413), .A(n11675), .ZN(n16109) );
  NAND2_X1 U13105 ( .A1(n16109), .A2(n14427), .ZN(n11201) );
  OAI211_X1 U13106 ( .C1(n16105), .C2(n14303), .A(n11202), .B(n11201), .ZN(
        P2_U3252) );
  AND2_X1 U13107 ( .A1(n11204), .A2(n11203), .ZN(n11207) );
  OAI211_X1 U13108 ( .C1(n11207), .C2(n11206), .A(n13527), .B(n11205), .ZN(
        n11213) );
  OAI22_X1 U13109 ( .A1(n13519), .A2(n11469), .B1(n11208), .B2(n13548), .ZN(
        n11209) );
  AOI211_X1 U13110 ( .C1(n11211), .C2(n13511), .A(n11210), .B(n11209), .ZN(
        n11212) );
  OAI211_X1 U13111 ( .C1(n11290), .C2(n13531), .A(n11213), .B(n11212), .ZN(
        P3_U3179) );
  MUX2_X1 U13112 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n7178), .Z(n11218) );
  NAND2_X1 U13113 ( .A1(n11218), .A2(SI_19_), .ZN(n11261) );
  OAI21_X1 U13114 ( .B1(n11217), .B2(n15184), .A(n11261), .ZN(n11214) );
  INV_X1 U13115 ( .A(n11214), .ZN(n11215) );
  NAND2_X1 U13116 ( .A1(n11216), .A2(n11215), .ZN(n11222) );
  NAND3_X1 U13117 ( .A1(n11261), .A2(n15184), .A3(n11217), .ZN(n11220) );
  INV_X1 U13118 ( .A(n11218), .ZN(n11219) );
  NAND2_X1 U13119 ( .A1(n11219), .A2(n15180), .ZN(n11260) );
  MUX2_X1 U13120 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n7178), .Z(n11351) );
  XNOR2_X1 U13121 ( .A(n11350), .B(n11351), .ZN(n12244) );
  INV_X1 U13122 ( .A(n12244), .ZN(n11348) );
  INV_X1 U13123 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11224) );
  OAI222_X1 U13124 ( .A1(n15167), .A2(n11348), .B1(P1_U3086), .B2(n12993), 
        .C1(n11224), .C2(n15157), .ZN(P1_U3335) );
  NAND2_X1 U13125 ( .A1(n11226), .A2(n11225), .ZN(n11228) );
  NAND2_X1 U13126 ( .A1(n11228), .A2(n11227), .ZN(n11439) );
  NAND2_X1 U13127 ( .A1(n11229), .A2(n12089), .ZN(n11232) );
  AOI22_X1 U13128 ( .A1(n13011), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n12008), 
        .B2(n11230), .ZN(n11231) );
  INV_X1 U13129 ( .A(n14741), .ZN(n11425) );
  XNOR2_X1 U13130 ( .A(n12875), .B(n11425), .ZN(n13042) );
  XNOR2_X1 U13131 ( .A(n11439), .B(n13042), .ZN(n11344) );
  INV_X1 U13132 ( .A(n11344), .ZN(n11253) );
  INV_X1 U13133 ( .A(n13042), .ZN(n11234) );
  OAI211_X1 U13134 ( .C1(n11235), .C2(n11234), .A(n11427), .B(n15955), .ZN(
        n11246) );
  NAND2_X1 U13135 ( .A1(n12987), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11243) );
  NAND2_X1 U13136 ( .A1(n11236), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n11430) );
  INV_X1 U13137 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n11237) );
  NAND2_X1 U13138 ( .A1(n11238), .A2(n11237), .ZN(n11239) );
  AND2_X1 U13139 ( .A1(n11430), .A2(n11239), .ZN(n11937) );
  NAND2_X1 U13140 ( .A1(n12095), .A2(n11937), .ZN(n11242) );
  NAND2_X1 U13141 ( .A1(n12988), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11241) );
  NAND2_X1 U13142 ( .A1(n12014), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n11240) );
  NAND4_X1 U13143 ( .A1(n11243), .A2(n11242), .A3(n11241), .A4(n11240), .ZN(
        n14740) );
  NAND2_X1 U13144 ( .A1(n14740), .A2(n14980), .ZN(n11245) );
  NAND2_X1 U13145 ( .A1(n14742), .A2(n14978), .ZN(n11244) );
  AND2_X1 U13146 ( .A1(n11245), .A2(n11244), .ZN(n11822) );
  NAND2_X1 U13147 ( .A1(n11246), .A2(n11822), .ZN(n11342) );
  NAND2_X1 U13148 ( .A1(n11247), .A2(n12875), .ZN(n11248) );
  NAND3_X1 U13149 ( .A1(n11454), .A2(n15041), .A3(n11248), .ZN(n11341) );
  AOI22_X1 U13150 ( .A1(n16047), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n11824), 
        .B2(n16037), .ZN(n11250) );
  NAND2_X1 U13151 ( .A1(n12875), .A2(n15990), .ZN(n11249) );
  OAI211_X1 U13152 ( .C1(n11341), .C2(n14997), .A(n11250), .B(n11249), .ZN(
        n11251) );
  AOI21_X1 U13153 ( .B1(n11342), .B2(n11899), .A(n11251), .ZN(n11252) );
  OAI21_X1 U13154 ( .B1(n11254), .B2(n11253), .A(n11252), .ZN(P1_U3281) );
  INV_X1 U13155 ( .A(n11255), .ZN(n11257) );
  NAND2_X1 U13156 ( .A1(n11257), .A2(n11256), .ZN(n11259) );
  OR2_X1 U13157 ( .A1(n11216), .A2(n15184), .ZN(n11258) );
  NAND2_X1 U13158 ( .A1(n11259), .A2(n11258), .ZN(n11263) );
  NAND2_X1 U13159 ( .A1(n11261), .A2(n11260), .ZN(n11262) );
  INV_X1 U13160 ( .A(n12233), .ZN(n11265) );
  OAI222_X1 U13161 ( .A1(n14588), .A2(n11264), .B1(n14593), .B2(n11265), .C1(
        P2_U3088), .C2(n14226), .ZN(P2_U3308) );
  OAI222_X1 U13162 ( .A1(n15157), .A2(n11266), .B1(n15167), .B2(n11265), .C1(
        n14836), .C2(P1_U3086), .ZN(P1_U3336) );
  XNOR2_X1 U13163 ( .A(n13203), .B(n14032), .ZN(n11373) );
  NAND2_X1 U13164 ( .A1(n14189), .A2(n14416), .ZN(n11270) );
  NOR2_X1 U13165 ( .A1(n11373), .A2(n11270), .ZN(n11379) );
  AOI21_X1 U13166 ( .B1(n11373), .B2(n11270), .A(n11379), .ZN(n11271) );
  OAI211_X1 U13167 ( .C1(n11272), .C2(n11271), .A(n11382), .B(n14115), .ZN(
        n11278) );
  NOR2_X1 U13168 ( .A1(n14144), .A2(n11273), .ZN(n11274) );
  AOI211_X1 U13169 ( .C1(n14141), .C2(n11276), .A(n11275), .B(n11274), .ZN(
        n11277) );
  OAI211_X1 U13170 ( .C1(n16073), .C2(n14162), .A(n11278), .B(n11277), .ZN(
        P2_U3208) );
  MUX2_X1 U13171 ( .A(n11280), .B(n11279), .S(n16101), .Z(n11281) );
  OAI21_X1 U13172 ( .B1(n16154), .B2(n12665), .A(n11281), .ZN(P3_U3464) );
  XNOR2_X1 U13173 ( .A(n11282), .B(n12668), .ZN(n15986) );
  NAND2_X1 U13174 ( .A1(n15986), .A2(n13754), .ZN(n11288) );
  NAND2_X1 U13175 ( .A1(n11283), .A2(n12668), .ZN(n11284) );
  NAND3_X1 U13176 ( .A1(n11285), .A2(n15881), .A3(n11284), .ZN(n11287) );
  AOI22_X1 U13177 ( .A1(n13572), .A2(n15873), .B1(n15876), .B2(n13574), .ZN(
        n11286) );
  NAND3_X1 U13178 ( .A1(n11288), .A2(n11287), .A3(n11286), .ZN(n15984) );
  MUX2_X1 U13179 ( .A(n15984), .B(P3_REG2_REG_6__SCAN_IN), .S(n13853), .Z(
        n11289) );
  INV_X1 U13180 ( .A(n11289), .ZN(n11293) );
  OAI22_X1 U13181 ( .A1(n13882), .A2(n15983), .B1(n11290), .B2(n15892), .ZN(
        n11291) );
  AOI21_X1 U13182 ( .B1(n15986), .B2(n13792), .A(n11291), .ZN(n11292) );
  NAND2_X1 U13183 ( .A1(n11293), .A2(n11292), .ZN(P3_U3227) );
  AND2_X1 U13184 ( .A1(n12518), .A2(n14743), .ZN(n11297) );
  AOI21_X1 U13185 ( .B1(n12864), .B2(n12519), .A(n11297), .ZN(n11479) );
  AOI22_X1 U13186 ( .A1(n12864), .A2(n12514), .B1(n12519), .B2(n14743), .ZN(
        n11298) );
  XNOR2_X1 U13187 ( .A(n11298), .B(n12526), .ZN(n11478) );
  XOR2_X1 U13188 ( .A(n11479), .B(n11478), .Z(n11299) );
  OAI211_X1 U13189 ( .C1(n11300), .C2(n11299), .A(n11477), .B(n14719), .ZN(
        n11306) );
  OAI21_X1 U13190 ( .B1(n14725), .B2(n11302), .A(n11301), .ZN(n11303) );
  AOI21_X1 U13191 ( .B1(n14728), .B2(n11304), .A(n11303), .ZN(n11305) );
  OAI211_X1 U13192 ( .C1(n11307), .C2(n14731), .A(n11306), .B(n11305), .ZN(
        P1_U3217) );
  NOR2_X1 U13193 ( .A1(n15685), .A2(n11309), .ZN(n11310) );
  XNOR2_X1 U13194 ( .A(n11309), .B(n15685), .ZN(n15679) );
  NAND2_X1 U13195 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n13628), .ZN(n11311) );
  OAI21_X1 U13196 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n13628), .A(n11311), 
        .ZN(n11312) );
  NOR2_X1 U13197 ( .A1(n11313), .A2(n11312), .ZN(n13611) );
  AOI21_X1 U13198 ( .B1(n11313), .B2(n11312), .A(n13611), .ZN(n11340) );
  INV_X1 U13199 ( .A(n11314), .ZN(n11316) );
  NAND2_X1 U13200 ( .A1(n11316), .A2(n11315), .ZN(n11317) );
  NAND2_X1 U13201 ( .A1(n11318), .A2(n11317), .ZN(n15682) );
  MUX2_X1 U13202 ( .A(n11320), .B(n11319), .S(n13664), .Z(n11321) );
  XNOR2_X1 U13203 ( .A(n11321), .B(n15685), .ZN(n15681) );
  INV_X1 U13204 ( .A(n11321), .ZN(n11323) );
  INV_X1 U13205 ( .A(n15685), .ZN(n11322) );
  NAND2_X1 U13206 ( .A1(n11323), .A2(n11322), .ZN(n11324) );
  MUX2_X1 U13207 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n13664), .Z(n13579) );
  XNOR2_X1 U13208 ( .A(n13579), .B(n13580), .ZN(n11325) );
  NAND2_X1 U13209 ( .A1(n11326), .A2(n11325), .ZN(n13583) );
  OAI21_X1 U13210 ( .B1(n11326), .B2(n11325), .A(n13583), .ZN(n11336) );
  NOR2_X1 U13211 ( .A1(n15685), .A2(n11329), .ZN(n11330) );
  NAND2_X1 U13212 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n13628), .ZN(n11331) );
  OAI21_X1 U13213 ( .B1(n13628), .B2(P3_REG1_REG_10__SCAN_IN), .A(n11331), 
        .ZN(n11332) );
  AOI21_X1 U13214 ( .B1(n11333), .B2(n11332), .A(n13627), .ZN(n11334) );
  NOR2_X1 U13215 ( .A1(n11334), .A2(n15822), .ZN(n11335) );
  AOI21_X1 U13216 ( .B1(n15775), .B2(n11336), .A(n11335), .ZN(n11339) );
  INV_X1 U13217 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n15347) );
  OR2_X1 U13218 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15347), .ZN(n11872) );
  OAI21_X1 U13219 ( .B1(n15808), .B2(n15564), .A(n11872), .ZN(n11337) );
  AOI21_X1 U13220 ( .B1(n13580), .B2(n15817), .A(n11337), .ZN(n11338) );
  OAI211_X1 U13221 ( .C1(n11340), .C2(n15825), .A(n11339), .B(n11338), .ZN(
        P3_U3192) );
  INV_X1 U13222 ( .A(n12875), .ZN(n11827) );
  OAI21_X1 U13223 ( .B1(n11827), .B2(n16058), .A(n11341), .ZN(n11343) );
  AOI211_X1 U13224 ( .C1(n11344), .C2(n16064), .A(n11343), .B(n11342), .ZN(
        n11347) );
  NAND2_X1 U13225 ( .A1(n16066), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11345) );
  OAI21_X1 U13226 ( .B1(n11347), .B2(n16066), .A(n11345), .ZN(P1_U3540) );
  NAND2_X1 U13227 ( .A1(n16068), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n11346) );
  OAI21_X1 U13228 ( .B1(n11347), .B2(n16068), .A(n11346), .ZN(P1_U3495) );
  OAI222_X1 U13229 ( .A1(n14588), .A2(n11349), .B1(P2_U3088), .B2(n13367), 
        .C1(n11348), .C2(n14593), .ZN(P2_U3307) );
  INV_X1 U13230 ( .A(n11352), .ZN(n11353) );
  MUX2_X1 U13231 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n7178), .Z(n11568) );
  XNOR2_X1 U13232 ( .A(n11568), .B(SI_21_), .ZN(n11565) );
  INV_X1 U13233 ( .A(n12259), .ZN(n11356) );
  OAI222_X1 U13234 ( .A1(n15157), .A2(n11355), .B1(n15167), .B2(n11356), .C1(
        n7920), .C2(P1_U3086), .ZN(P1_U3334) );
  OAI222_X1 U13235 ( .A1(n14588), .A2(n11357), .B1(n14593), .B2(n11356), .C1(
        P2_U3088), .C2(n13405), .ZN(P2_U3306) );
  INV_X1 U13236 ( .A(n11358), .ZN(n11360) );
  AOI21_X1 U13237 ( .B1(n11360), .B2(n11365), .A(n11359), .ZN(n11363) );
  INV_X1 U13238 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11361) );
  NOR2_X1 U13239 ( .A1(n11646), .A2(n11361), .ZN(n11522) );
  AOI21_X1 U13240 ( .B1(n11361), .B2(n11646), .A(n11522), .ZN(n11362) );
  NAND2_X1 U13241 ( .A1(n11362), .A2(n11363), .ZN(n11523) );
  OAI211_X1 U13242 ( .C1(n11363), .C2(n11362), .A(n14833), .B(n11523), .ZN(
        n11372) );
  NAND2_X1 U13243 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14653)
         );
  AOI21_X1 U13244 ( .B1(n11366), .B2(n11365), .A(n11364), .ZN(n11368) );
  XNOR2_X1 U13245 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n11646), .ZN(n11367) );
  NAND2_X1 U13246 ( .A1(n11367), .A2(n11368), .ZN(n11528) );
  OAI211_X1 U13247 ( .C1(n11368), .C2(n11367), .A(n14834), .B(n11528), .ZN(
        n11369) );
  NAND2_X1 U13248 ( .A1(n14653), .A2(n11369), .ZN(n11370) );
  AOI21_X1 U13249 ( .B1(n14797), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11370), 
        .ZN(n11371) );
  OAI211_X1 U13250 ( .C1(n14828), .C2(n11646), .A(n11372), .B(n11371), .ZN(
        P1_U3259) );
  NOR3_X1 U13251 ( .A1(n11373), .A2(n11388), .A3(n14152), .ZN(n11385) );
  XNOR2_X1 U13252 ( .A(n13208), .B(n14043), .ZN(n11676) );
  AND2_X1 U13253 ( .A1(n14188), .A2(n14416), .ZN(n11375) );
  NAND2_X1 U13254 ( .A1(n11676), .A2(n11375), .ZN(n11681) );
  INV_X1 U13255 ( .A(n11676), .ZN(n11377) );
  INV_X1 U13256 ( .A(n11375), .ZN(n11376) );
  NAND2_X1 U13257 ( .A1(n11377), .A2(n11376), .ZN(n11378) );
  NAND2_X1 U13258 ( .A1(n11681), .A2(n11378), .ZN(n11380) );
  AOI21_X1 U13259 ( .B1(n11382), .B2(n11380), .A(n14168), .ZN(n11384) );
  INV_X1 U13260 ( .A(n11379), .ZN(n11381) );
  INV_X1 U13261 ( .A(n11684), .ZN(n11383) );
  OAI21_X1 U13262 ( .B1(n11385), .B2(n11384), .A(n11383), .ZN(n11392) );
  OAI22_X1 U13263 ( .A1(n14161), .A2(n11387), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11386), .ZN(n11390) );
  NOR2_X1 U13264 ( .A1(n14096), .A2(n11388), .ZN(n11389) );
  AOI211_X1 U13265 ( .C1(n14099), .C2(n14187), .A(n11390), .B(n11389), .ZN(
        n11391) );
  OAI211_X1 U13266 ( .C1(n16088), .C2(n14162), .A(n11392), .B(n11391), .ZN(
        P2_U3196) );
  XOR2_X1 U13267 ( .A(n11394), .B(n11393), .Z(n11395) );
  NAND2_X1 U13268 ( .A1(n11395), .A2(n13527), .ZN(n11399) );
  INV_X1 U13269 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n15338) );
  NOR2_X1 U13270 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15338), .ZN(n15666) );
  OAI22_X1 U13271 ( .A1(n13519), .A2(n12687), .B1(n11596), .B2(n13548), .ZN(
        n11396) );
  AOI211_X1 U13272 ( .C1(n11397), .C2(n13511), .A(n15666), .B(n11396), .ZN(
        n11398) );
  OAI211_X1 U13273 ( .C1(n11593), .C2(n13531), .A(n11399), .B(n11398), .ZN(
        P3_U3153) );
  XNOR2_X1 U13274 ( .A(n11400), .B(n12603), .ZN(n16006) );
  OAI21_X1 U13275 ( .B1(n12603), .B2(n11402), .A(n11401), .ZN(n11404) );
  OAI22_X1 U13276 ( .A1(n11693), .A2(n15390), .B1(n11469), .B2(n15392), .ZN(
        n11403) );
  AOI21_X1 U13277 ( .B1(n11404), .B2(n15881), .A(n11403), .ZN(n11405) );
  OAI21_X1 U13278 ( .B1(n15886), .B2(n16006), .A(n11405), .ZN(n16008) );
  NAND2_X1 U13279 ( .A1(n16008), .A2(n15899), .ZN(n11408) );
  OAI22_X1 U13280 ( .A1(n13882), .A2(n16005), .B1(n11474), .B2(n15892), .ZN(
        n11406) );
  AOI21_X1 U13281 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n13853), .A(n11406), .ZN(
        n11407) );
  OAI211_X1 U13282 ( .C1(n16006), .C2(n15402), .A(n11408), .B(n11407), .ZN(
        P3_U3225) );
  NAND2_X1 U13283 ( .A1(n11488), .A2(n12089), .ZN(n11411) );
  AOI22_X1 U13284 ( .A1(n11409), .A2(n12008), .B1(n13011), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n11410) );
  NAND2_X1 U13285 ( .A1(n11412), .A2(n12089), .ZN(n11415) );
  AOI22_X1 U13286 ( .A1(n13011), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n11413), 
        .B2(n12008), .ZN(n11414) );
  AOI211_X1 U13287 ( .C1(n16128), .C2(n11455), .A(n15952), .B(n11638), .ZN(
        n11424) );
  INV_X1 U13288 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n11422) );
  NAND2_X1 U13289 ( .A1(n12987), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n11417) );
  NAND2_X1 U13290 ( .A1(n12988), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n11416) );
  AND2_X1 U13291 ( .A1(n11417), .A2(n11416), .ZN(n11421) );
  NAND2_X1 U13292 ( .A1(n11432), .A2(n14723), .ZN(n11419) );
  NAND2_X1 U13293 ( .A1(n11631), .A2(n11419), .ZN(n11641) );
  OR2_X1 U13294 ( .A1(n11641), .A2(n12142), .ZN(n11420) );
  OAI211_X1 U13295 ( .C1(n12992), .C2(n11422), .A(n11421), .B(n11420), .ZN(
        n14738) );
  INV_X1 U13296 ( .A(n14738), .ZN(n16116) );
  INV_X1 U13297 ( .A(n14740), .ZN(n16117) );
  OAI22_X1 U13298 ( .A1(n16116), .A2(n15005), .B1(n16117), .B2(n15003), .ZN(
        n11423) );
  NOR2_X1 U13299 ( .A1(n11424), .A2(n11423), .ZN(n11613) );
  INV_X1 U13300 ( .A(n11613), .ZN(n11438) );
  OR2_X1 U13301 ( .A1(n12875), .A2(n11425), .ZN(n11426) );
  XNOR2_X1 U13302 ( .A(n12885), .B(n16117), .ZN(n13043) );
  OR2_X1 U13303 ( .A1(n12885), .A2(n16117), .ZN(n11428) );
  NAND2_X1 U13304 ( .A1(n11430), .A2(n11429), .ZN(n11431) );
  NAND2_X1 U13305 ( .A1(n11432), .A2(n11431), .ZN(n16132) );
  INV_X1 U13306 ( .A(n16132), .ZN(n11445) );
  NAND2_X1 U13307 ( .A1(n11445), .A2(n12095), .ZN(n11436) );
  NAND2_X1 U13308 ( .A1(n12987), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11435) );
  NAND2_X1 U13309 ( .A1(n12014), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n11434) );
  NAND2_X1 U13310 ( .A1(n12988), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11433) );
  NAND4_X1 U13311 ( .A1(n11436), .A2(n11435), .A3(n11434), .A4(n11433), .ZN(
        n14739) );
  INV_X1 U13312 ( .A(n14739), .ZN(n11623) );
  XNOR2_X1 U13313 ( .A(n16128), .B(n11623), .ZN(n13044) );
  XNOR2_X1 U13314 ( .A(n11622), .B(n11444), .ZN(n11437) );
  NOR2_X1 U13315 ( .A1(n11437), .A2(n16060), .ZN(n11615) );
  AOI21_X1 U13316 ( .B1(n14836), .B2(n11438), .A(n11615), .ZN(n11449) );
  NAND2_X1 U13317 ( .A1(n11439), .A2(n13042), .ZN(n11441) );
  OR2_X1 U13318 ( .A1(n12875), .A2(n14741), .ZN(n11440) );
  NAND2_X1 U13319 ( .A1(n11441), .A2(n11440), .ZN(n11453) );
  OR2_X1 U13320 ( .A1(n12885), .A2(n14740), .ZN(n11442) );
  AOI21_X1 U13321 ( .B1(n11444), .B2(n11443), .A(n7315), .ZN(n11617) );
  INV_X1 U13322 ( .A(n16128), .ZN(n11614) );
  AOI22_X1 U13323 ( .A1(n16047), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n11445), 
        .B2(n16037), .ZN(n11446) );
  OAI21_X1 U13324 ( .B1(n11614), .B2(n16041), .A(n11446), .ZN(n11447) );
  AOI21_X1 U13325 ( .B1(n11617), .B2(n14999), .A(n11447), .ZN(n11448) );
  OAI21_X1 U13326 ( .B1(n11449), .B2(n15998), .A(n11448), .ZN(P1_U3279) );
  INV_X1 U13327 ( .A(n11450), .ZN(n11451) );
  OAI222_X1 U13328 ( .A1(P3_U3151), .A2(n11452), .B1(n13083), .B2(n15201), 
        .C1(n13082), .C2(n11451), .ZN(P3_U3271) );
  XNOR2_X1 U13329 ( .A(n11453), .B(n13043), .ZN(n11518) );
  INV_X1 U13330 ( .A(n11518), .ZN(n11465) );
  INV_X1 U13331 ( .A(n12885), .ZN(n11940) );
  INV_X1 U13332 ( .A(n11454), .ZN(n11456) );
  OAI211_X1 U13333 ( .C1(n11940), .C2(n11456), .A(n15041), .B(n11455), .ZN(
        n11513) );
  AOI22_X1 U13334 ( .A1(n14980), .A2(n14739), .B1(n14741), .B2(n14978), .ZN(
        n11935) );
  NAND2_X1 U13335 ( .A1(n16037), .A2(n11937), .ZN(n11457) );
  OAI211_X1 U13336 ( .C1(n11513), .C2(n13059), .A(n11935), .B(n11457), .ZN(
        n11463) );
  INV_X1 U13337 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11458) );
  OAI22_X1 U13338 ( .A1(n11940), .A2(n16041), .B1(n11458), .B2(n11899), .ZN(
        n11462) );
  NOR2_X1 U13339 ( .A1(n11459), .A2(n7709), .ZN(n11515) );
  INV_X1 U13340 ( .A(n11460), .ZN(n11514) );
  NOR3_X1 U13341 ( .A1(n11515), .A2(n11514), .A3(n15001), .ZN(n11461) );
  AOI211_X1 U13342 ( .C1(n11899), .C2(n11463), .A(n11462), .B(n11461), .ZN(
        n11464) );
  OAI21_X1 U13343 ( .B1(n14967), .B2(n11465), .A(n11464), .ZN(P1_U3280) );
  XOR2_X1 U13344 ( .A(n11467), .B(n11466), .Z(n11468) );
  NAND2_X1 U13345 ( .A1(n11468), .A2(n13527), .ZN(n11473) );
  OAI22_X1 U13346 ( .A1(n13519), .A2(n11693), .B1(n11469), .B2(n13548), .ZN(
        n11470) );
  AOI211_X1 U13347 ( .C1(n12682), .C2(n13511), .A(n11471), .B(n11470), .ZN(
        n11472) );
  OAI211_X1 U13348 ( .C1(n11474), .C2(n13531), .A(n11473), .B(n11472), .ZN(
        P3_U3161) );
  OAI22_X1 U13349 ( .A1(n16059), .A2(n12523), .B1(n11476), .B2(n12525), .ZN(
        n11475) );
  XNOR2_X1 U13350 ( .A(n11475), .B(n12526), .ZN(n11813) );
  OAI22_X1 U13351 ( .A1(n16059), .A2(n12525), .B1(n11476), .B2(n12524), .ZN(
        n11812) );
  XNOR2_X1 U13352 ( .A(n11813), .B(n11812), .ZN(n11481) );
  AOI21_X1 U13353 ( .B1(n11481), .B2(n11480), .A(n11814), .ZN(n11487) );
  OAI22_X1 U13354 ( .A1(n14725), .A2(n16056), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11482), .ZN(n11484) );
  NOR2_X1 U13355 ( .A1(n16059), .A2(n14731), .ZN(n11483) );
  AOI211_X1 U13356 ( .C1(n14728), .C2(n11485), .A(n11484), .B(n11483), .ZN(
        n11486) );
  OAI21_X1 U13357 ( .B1(n11487), .B2(n16123), .A(n11486), .ZN(P1_U3236) );
  OAI22_X1 U13358 ( .A1(n11769), .A2(n11785), .B1(n9957), .B2(n11489), .ZN(
        n11490) );
  INV_X1 U13359 ( .A(n11490), .ZN(n11491) );
  INV_X1 U13360 ( .A(n14186), .ZN(n11543) );
  XNOR2_X1 U13361 ( .A(n13224), .B(n11543), .ZN(n13388) );
  INV_X1 U13362 ( .A(n14187), .ZN(n11711) );
  NOR2_X1 U13363 ( .A1(n13216), .A2(n11711), .ZN(n11493) );
  NAND2_X1 U13364 ( .A1(n13216), .A2(n11711), .ZN(n11495) );
  XOR2_X1 U13365 ( .A(n13388), .B(n11542), .Z(n11503) );
  INV_X1 U13366 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n11496) );
  NAND2_X1 U13367 ( .A1(n11497), .A2(n11496), .ZN(n11498) );
  NAND2_X1 U13368 ( .A1(n11552), .A2(n11498), .ZN(n11918) );
  NAND2_X1 U13369 ( .A1(n13322), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n11500) );
  INV_X1 U13370 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n11560) );
  OR2_X1 U13371 ( .A1(n12239), .A2(n11560), .ZN(n11499) );
  AND2_X1 U13372 ( .A1(n11500), .A2(n11499), .ZN(n11502) );
  NAND2_X1 U13373 ( .A1(n12336), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n11501) );
  OAI211_X1 U13374 ( .C1(n11918), .C2(n12314), .A(n11502), .B(n11501), .ZN(
        n14185) );
  AOI222_X1 U13375 ( .A1(n14393), .A2(n11503), .B1(n14185), .B2(n14139), .C1(
        n14187), .C2(n14137), .ZN(n16135) );
  INV_X1 U13376 ( .A(n11504), .ZN(n11708) );
  OAI22_X1 U13377 ( .A1(n14427), .A2(n11505), .B1(n11708), .B2(n14430), .ZN(
        n11509) );
  INV_X1 U13378 ( .A(n13224), .ZN(n16137) );
  INV_X1 U13379 ( .A(n11538), .ZN(n11540) );
  OAI211_X1 U13380 ( .C1(n16137), .C2(n11507), .A(n11540), .B(n14397), .ZN(
        n16134) );
  NOR2_X1 U13381 ( .A1(n16134), .A2(n14420), .ZN(n11508) );
  AOI211_X1 U13382 ( .C1(n14434), .C2(n13224), .A(n11509), .B(n11508), .ZN(
        n11512) );
  XOR2_X1 U13383 ( .A(n13388), .B(n11545), .Z(n16139) );
  NAND2_X1 U13384 ( .A1(n16139), .A2(n14436), .ZN(n11511) );
  OAI211_X1 U13385 ( .C1(n16135), .C2(n14378), .A(n11512), .B(n11511), .ZN(
        P2_U3251) );
  OAI211_X1 U13386 ( .C1(n11940), .C2(n16058), .A(n11513), .B(n11935), .ZN(
        n11517) );
  NOR3_X1 U13387 ( .A1(n11515), .A2(n11514), .A3(n16060), .ZN(n11516) );
  AOI211_X1 U13388 ( .C1(n11518), .C2(n16064), .A(n11517), .B(n11516), .ZN(
        n11521) );
  NAND2_X1 U13389 ( .A1(n16068), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n11519) );
  OAI21_X1 U13390 ( .B1(n11521), .B2(n16068), .A(n11519), .ZN(P1_U3498) );
  NAND2_X1 U13391 ( .A1(n16066), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11520) );
  OAI21_X1 U13392 ( .B1(n11521), .B2(n16066), .A(n11520), .ZN(P1_U3541) );
  INV_X1 U13393 ( .A(n11522), .ZN(n11524) );
  NAND2_X1 U13394 ( .A1(n11524), .A2(n11523), .ZN(n11527) );
  INV_X1 U13395 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n11907) );
  NOR2_X1 U13396 ( .A1(n11910), .A2(n11907), .ZN(n11525) );
  AOI21_X1 U13397 ( .B1(n11907), .B2(n11910), .A(n11525), .ZN(n11526) );
  NAND2_X1 U13398 ( .A1(n11526), .A2(n11527), .ZN(n11906) );
  OAI211_X1 U13399 ( .C1(n11527), .C2(n11526), .A(n14833), .B(n11906), .ZN(
        n11535) );
  NAND2_X1 U13400 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14663)
         );
  XNOR2_X1 U13401 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n11910), .ZN(n11531) );
  INV_X1 U13402 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n11529) );
  OAI21_X1 U13403 ( .B1(n11646), .B2(n11529), .A(n11528), .ZN(n11530) );
  NAND2_X1 U13404 ( .A1(n11531), .A2(n11530), .ZN(n11909) );
  OAI211_X1 U13405 ( .C1(n11531), .C2(n11530), .A(n11909), .B(n14834), .ZN(
        n11532) );
  NAND2_X1 U13406 ( .A1(n14663), .A2(n11532), .ZN(n11533) );
  AOI21_X1 U13407 ( .B1(n14797), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n11533), 
        .ZN(n11534) );
  OAI211_X1 U13408 ( .C1(n14828), .C2(n11910), .A(n11535), .B(n11534), .ZN(
        P1_U3260) );
  AOI22_X1 U13409 ( .A1(n11770), .A2(n12234), .B1(n13330), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n11536) );
  NAND2_X1 U13410 ( .A1(n11837), .A2(n11538), .ZN(n11740) );
  INV_X1 U13411 ( .A(n11740), .ZN(n11539) );
  AOI211_X1 U13412 ( .C1(n13230), .C2(n11540), .A(n14416), .B(n11539), .ZN(
        n11830) );
  AND2_X1 U13413 ( .A1(n13224), .A2(n11543), .ZN(n11541) );
  OR2_X1 U13414 ( .A1(n13224), .A2(n11543), .ZN(n11544) );
  XNOR2_X1 U13415 ( .A(n13230), .B(n14185), .ZN(n13389) );
  XNOR2_X1 U13416 ( .A(n11733), .B(n13389), .ZN(n11559) );
  NAND2_X1 U13417 ( .A1(n13224), .A2(n14186), .ZN(n11546) );
  NAND2_X1 U13418 ( .A1(n11547), .A2(n11546), .ZN(n11548) );
  NAND2_X1 U13419 ( .A1(n11548), .A2(n13389), .ZN(n11549) );
  NAND2_X1 U13420 ( .A1(n11721), .A2(n11549), .ZN(n11831) );
  NAND2_X1 U13421 ( .A1(n11831), .A2(n15907), .ZN(n11558) );
  INV_X1 U13422 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n11556) );
  INV_X1 U13423 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n11551) );
  NAND2_X1 U13424 ( .A1(n11552), .A2(n11551), .ZN(n11553) );
  NAND2_X1 U13425 ( .A1(n11728), .A2(n11553), .ZN(n11848) );
  OR2_X1 U13426 ( .A1(n11848), .A2(n12314), .ZN(n11555) );
  AOI22_X1 U13427 ( .A1(n13321), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n13322), 
        .B2(P2_REG1_REG_16__SCAN_IN), .ZN(n11554) );
  OAI211_X1 U13428 ( .C1(n13325), .C2(n11556), .A(n11555), .B(n11554), .ZN(
        n14184) );
  AND2_X1 U13429 ( .A1(n14186), .A2(n14137), .ZN(n11557) );
  AOI21_X1 U13430 ( .B1(n14184), .B2(n14139), .A(n11557), .ZN(n11921) );
  OAI211_X1 U13431 ( .C1(n14413), .C2(n11559), .A(n11558), .B(n11921), .ZN(
        n11829) );
  AOI21_X1 U13432 ( .B1(n11830), .B2(n14226), .A(n11829), .ZN(n11564) );
  NOR2_X1 U13433 ( .A1(n11837), .A2(n14366), .ZN(n11562) );
  OAI22_X1 U13434 ( .A1(n14427), .A2(n11560), .B1(n11918), .B2(n14430), .ZN(
        n11561) );
  AOI211_X1 U13435 ( .C1(n11831), .C2(n11746), .A(n11562), .B(n11561), .ZN(
        n11563) );
  OAI21_X1 U13436 ( .B1(n11564), .B2(n14378), .A(n11563), .ZN(P2_U3250) );
  INV_X1 U13437 ( .A(n11565), .ZN(n11566) );
  NAND2_X1 U13438 ( .A1(n11568), .A2(SI_21_), .ZN(n11569) );
  XNOR2_X2 U13439 ( .A(n11748), .B(n15181), .ZN(n12047) );
  MUX2_X1 U13440 ( .A(n11577), .B(n11571), .S(n7178), .Z(n11572) );
  INV_X1 U13441 ( .A(n12047), .ZN(n11574) );
  INV_X1 U13442 ( .A(n11572), .ZN(n11573) );
  NAND2_X1 U13443 ( .A1(n11574), .A2(n11573), .ZN(n11575) );
  NAND2_X1 U13444 ( .A1(n11750), .A2(n11575), .ZN(n12271) );
  INV_X1 U13445 ( .A(n12271), .ZN(n11576) );
  OAI222_X1 U13446 ( .A1(n14588), .A2(n11577), .B1(n14593), .B2(n11576), .C1(
        n13411), .C2(P2_U3088), .ZN(P2_U3305) );
  INV_X1 U13447 ( .A(n11578), .ZN(n12685) );
  XNOR2_X1 U13448 ( .A(n11580), .B(n8177), .ZN(n11583) );
  INV_X1 U13449 ( .A(n11583), .ZN(n16027) );
  XNOR2_X1 U13450 ( .A(n11581), .B(n8177), .ZN(n11585) );
  OAI22_X1 U13451 ( .A1(n12687), .A2(n15392), .B1(n11859), .B2(n15390), .ZN(
        n11582) );
  AOI21_X1 U13452 ( .B1(n11583), .B2(n13754), .A(n11582), .ZN(n11584) );
  OAI21_X1 U13453 ( .B1(n11585), .B2(n13874), .A(n11584), .ZN(n16029) );
  NAND2_X1 U13454 ( .A1(n16029), .A2(n15899), .ZN(n11588) );
  OAI22_X1 U13455 ( .A1(n13882), .A2(n16026), .B1(n11608), .B2(n15892), .ZN(
        n11586) );
  AOI21_X1 U13456 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n13853), .A(n11586), .ZN(
        n11587) );
  OAI211_X1 U13457 ( .C1(n16027), .C2(n15402), .A(n11588), .B(n11587), .ZN(
        P3_U3224) );
  OAI222_X1 U13458 ( .A1(P3_U3151), .A2(n11590), .B1(n13083), .B2(n11982), 
        .C1(n13082), .C2(n11589), .ZN(P3_U3270) );
  XNOR2_X1 U13459 ( .A(n11592), .B(n11591), .ZN(n16000) );
  INV_X1 U13460 ( .A(n16000), .ZN(n11602) );
  OAI22_X1 U13461 ( .A1(n13882), .A2(n15999), .B1(n11593), .B2(n15892), .ZN(
        n11601) );
  XNOR2_X1 U13462 ( .A(n11594), .B(n12675), .ZN(n11595) );
  NAND2_X1 U13463 ( .A1(n11595), .A2(n15881), .ZN(n11599) );
  OAI22_X1 U13464 ( .A1(n11596), .A2(n15392), .B1(n12687), .B2(n15390), .ZN(
        n11597) );
  INV_X1 U13465 ( .A(n11597), .ZN(n11598) );
  OAI211_X1 U13466 ( .C1(n15886), .C2(n16000), .A(n11599), .B(n11598), .ZN(
        n16002) );
  MUX2_X1 U13467 ( .A(n16002), .B(P3_REG2_REG_7__SCAN_IN), .S(n13853), .Z(
        n11600) );
  AOI211_X1 U13468 ( .C1(n11602), .C2(n13792), .A(n11601), .B(n11600), .ZN(
        n11603) );
  INV_X1 U13469 ( .A(n11603), .ZN(P3_U3226) );
  AOI21_X1 U13470 ( .B1(n11605), .B2(n11604), .A(n7324), .ZN(n11612) );
  NAND2_X1 U13471 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n15690) );
  INV_X1 U13472 ( .A(n15690), .ZN(n11607) );
  OAI22_X1 U13473 ( .A1(n13519), .A2(n11859), .B1(n13554), .B2(n16026), .ZN(
        n11606) );
  AOI211_X1 U13474 ( .C1(n13529), .C2(n13571), .A(n11607), .B(n11606), .ZN(
        n11611) );
  INV_X1 U13475 ( .A(n11608), .ZN(n11609) );
  NAND2_X1 U13476 ( .A1(n13550), .A2(n11609), .ZN(n11610) );
  OAI211_X1 U13477 ( .C1(n11612), .C2(n13539), .A(n11611), .B(n11610), .ZN(
        P3_U3171) );
  OAI21_X1 U13478 ( .B1(n11614), .B2(n16058), .A(n11613), .ZN(n11616) );
  AOI211_X1 U13479 ( .C1(n11617), .C2(n16064), .A(n11616), .B(n11615), .ZN(
        n11620) );
  NAND2_X1 U13480 ( .A1(n16068), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n11618) );
  OAI21_X1 U13481 ( .B1(n11620), .B2(n16068), .A(n11618), .ZN(P1_U3501) );
  NAND2_X1 U13482 ( .A1(n16066), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11619) );
  OAI21_X1 U13483 ( .B1(n11620), .B2(n16066), .A(n11619), .ZN(P1_U3542) );
  NAND2_X1 U13484 ( .A1(n16128), .A2(n11623), .ZN(n11621) );
  OR2_X1 U13485 ( .A1(n16128), .A2(n11623), .ZN(n11624) );
  NAND2_X1 U13486 ( .A1(n11626), .A2(n12089), .ZN(n11629) );
  AOI22_X1 U13487 ( .A1(n13011), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n12008), 
        .B2(n11627), .ZN(n11628) );
  XNOR2_X1 U13488 ( .A(n15122), .B(n16116), .ZN(n13048) );
  XNOR2_X1 U13489 ( .A(n11650), .B(n13048), .ZN(n11637) );
  NAND2_X1 U13490 ( .A1(n11631), .A2(n11630), .ZN(n11632) );
  NAND2_X1 U13491 ( .A1(n11655), .A2(n11632), .ZN(n14652) );
  AOI22_X1 U13492 ( .A1(n12987), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n12014), 
        .B2(P1_REG0_REG_16__SCAN_IN), .ZN(n11634) );
  NAND2_X1 U13493 ( .A1(n12988), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11633) );
  OAI211_X1 U13494 ( .C1(n14652), .C2(n12142), .A(n11634), .B(n11633), .ZN(
        n14737) );
  AND2_X1 U13495 ( .A1(n14739), .A2(n14978), .ZN(n11635) );
  AOI21_X1 U13496 ( .B1(n14737), .B2(n14980), .A(n11635), .ZN(n14724) );
  INV_X1 U13497 ( .A(n14724), .ZN(n11636) );
  AOI21_X1 U13498 ( .B1(n11637), .B2(n15955), .A(n11636), .ZN(n15124) );
  INV_X1 U13499 ( .A(n11638), .ZN(n11640) );
  INV_X1 U13500 ( .A(n11651), .ZN(n11639) );
  AOI211_X1 U13501 ( .C1(n15122), .C2(n11640), .A(n15952), .B(n11639), .ZN(
        n15121) );
  INV_X1 U13502 ( .A(n11641), .ZN(n14727) );
  AOI22_X1 U13503 ( .A1(n16047), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n14727), 
        .B2(n16037), .ZN(n11642) );
  OAI21_X1 U13504 ( .B1(n14732), .B2(n16041), .A(n11642), .ZN(n11644) );
  XNOR2_X1 U13505 ( .A(n11670), .B(n13048), .ZN(n15125) );
  NOR2_X1 U13506 ( .A1(n15125), .A2(n14967), .ZN(n11643) );
  AOI211_X1 U13507 ( .C1(n15121), .C2(n16035), .A(n11644), .B(n11643), .ZN(
        n11645) );
  OAI21_X1 U13508 ( .B1(n15998), .B2(n15124), .A(n11645), .ZN(P1_U3278) );
  NAND2_X1 U13509 ( .A1(n11722), .A2(n12089), .ZN(n11649) );
  INV_X1 U13510 ( .A(n11646), .ZN(n11647) );
  AOI22_X1 U13511 ( .A1(n13011), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n12008), 
        .B2(n11647), .ZN(n11648) );
  INV_X1 U13512 ( .A(n14737), .ZN(n14664) );
  INV_X1 U13513 ( .A(n13048), .ZN(n11669) );
  XOR2_X1 U13514 ( .A(n13046), .B(n11901), .Z(n15120) );
  AOI21_X1 U13515 ( .B1(n14656), .B2(n11651), .A(n15952), .ZN(n11652) );
  NAND2_X1 U13516 ( .A1(n11652), .A2(n11887), .ZN(n15115) );
  INV_X1 U13517 ( .A(n15115), .ZN(n11667) );
  INV_X1 U13518 ( .A(n14656), .ZN(n15116) );
  INV_X1 U13519 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n11654) );
  NAND2_X1 U13520 ( .A1(n11655), .A2(n11654), .ZN(n11656) );
  NAND2_X1 U13521 ( .A1(n11889), .A2(n11656), .ZN(n14667) );
  OR2_X1 U13522 ( .A1(n14667), .A2(n12142), .ZN(n11662) );
  INV_X1 U13523 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n11911) );
  NAND2_X1 U13524 ( .A1(n12988), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11658) );
  NAND2_X1 U13525 ( .A1(n12014), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n11657) );
  OAI211_X1 U13526 ( .C1(n11659), .C2(n11911), .A(n11658), .B(n11657), .ZN(
        n11660) );
  INV_X1 U13527 ( .A(n11660), .ZN(n11661) );
  NAND2_X1 U13528 ( .A1(n11662), .A2(n11661), .ZN(n14736) );
  AND2_X1 U13529 ( .A1(n14738), .A2(n14978), .ZN(n11663) );
  AOI21_X1 U13530 ( .B1(n14736), .B2(n14980), .A(n11663), .ZN(n15114) );
  OAI22_X1 U13531 ( .A1(n16047), .A2(n15114), .B1(n14652), .B2(n15016), .ZN(
        n11664) );
  AOI21_X1 U13532 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n15998), .A(n11664), 
        .ZN(n11665) );
  OAI21_X1 U13533 ( .B1(n15116), .B2(n16041), .A(n11665), .ZN(n11666) );
  AOI21_X1 U13534 ( .B1(n11667), .B2(n16035), .A(n11666), .ZN(n11672) );
  OR2_X1 U13535 ( .A1(n15122), .A2(n14738), .ZN(n11668) );
  XNOR2_X1 U13536 ( .A(n11877), .B(n13046), .ZN(n15118) );
  NAND2_X1 U13537 ( .A1(n15118), .A2(n14999), .ZN(n11671) );
  OAI211_X1 U13538 ( .C1(n15120), .C2(n15001), .A(n11672), .B(n11671), .ZN(
        P1_U3277) );
  AOI22_X1 U13539 ( .A1(n14141), .A2(n11673), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11674) );
  OAI21_X1 U13540 ( .B1(n14144), .B2(n11675), .A(n11674), .ZN(n11688) );
  NAND3_X1 U13541 ( .A1(n11676), .A2(n14063), .A3(n14188), .ZN(n11686) );
  XNOR2_X1 U13542 ( .A(n13216), .B(n14043), .ZN(n11677) );
  AND2_X1 U13543 ( .A1(n14187), .A2(n14416), .ZN(n11678) );
  NAND2_X1 U13544 ( .A1(n11677), .A2(n11678), .ZN(n11705) );
  INV_X1 U13545 ( .A(n11677), .ZN(n11712) );
  INV_X1 U13546 ( .A(n11678), .ZN(n11679) );
  NAND2_X1 U13547 ( .A1(n11712), .A2(n11679), .ZN(n11680) );
  AND2_X1 U13548 ( .A1(n11705), .A2(n11680), .ZN(n11682) );
  OAI21_X1 U13549 ( .B1(n11684), .B2(n11682), .A(n14115), .ZN(n11685) );
  INV_X1 U13550 ( .A(n11681), .ZN(n11683) );
  INV_X1 U13551 ( .A(n11706), .ZN(n11714) );
  AOI21_X1 U13552 ( .B1(n11686), .B2(n11685), .A(n11714), .ZN(n11687) );
  AOI211_X1 U13553 ( .C1(n13216), .C2(n14150), .A(n11688), .B(n11687), .ZN(
        n11689) );
  INV_X1 U13554 ( .A(n11689), .ZN(P2_U3206) );
  NAND2_X1 U13555 ( .A1(n11691), .A2(n11690), .ZN(n11692) );
  AOI21_X1 U13556 ( .B1(n11692), .B2(n12691), .A(n13874), .ZN(n11696) );
  OAI22_X1 U13557 ( .A1(n11693), .A2(n15392), .B1(n11961), .B2(n15390), .ZN(
        n11694) );
  AOI21_X1 U13558 ( .B1(n11696), .B2(n11695), .A(n11694), .ZN(n13958) );
  OAI21_X1 U13559 ( .B1(n7323), .B2(n12691), .A(n11697), .ZN(n13956) );
  NAND2_X1 U13560 ( .A1(n15886), .A2(n11698), .ZN(n11699) );
  NAND2_X1 U13561 ( .A1(n15899), .A2(n11699), .ZN(n13868) );
  NOR2_X1 U13562 ( .A1(n15899), .A2(n11700), .ZN(n11703) );
  OAI22_X1 U13563 ( .A1(n13882), .A2(n11701), .B1(n11876), .B2(n15892), .ZN(
        n11702) );
  AOI211_X1 U13564 ( .C1(n13956), .C2(n13887), .A(n11703), .B(n11702), .ZN(
        n11704) );
  OAI21_X1 U13565 ( .B1(n13958), .B2(n13853), .A(n11704), .ZN(P3_U3223) );
  XNOR2_X1 U13566 ( .A(n13224), .B(n14043), .ZN(n11840) );
  NAND2_X1 U13567 ( .A1(n14186), .A2(n14416), .ZN(n11838) );
  XNOR2_X1 U13568 ( .A(n11840), .B(n11838), .ZN(n11715) );
  OAI21_X1 U13569 ( .B1(n14161), .B2(n11708), .A(n11707), .ZN(n11709) );
  AOI21_X1 U13570 ( .B1(n14099), .B2(n14185), .A(n11709), .ZN(n11710) );
  OAI21_X1 U13571 ( .B1(n11711), .B2(n14096), .A(n11710), .ZN(n11718) );
  NOR3_X1 U13572 ( .A1(n11712), .A2(n11711), .A3(n14152), .ZN(n11713) );
  AOI21_X1 U13573 ( .B1(n11714), .B2(n14115), .A(n11713), .ZN(n11716) );
  NOR2_X1 U13574 ( .A1(n11716), .A2(n11715), .ZN(n11717) );
  AOI211_X1 U13575 ( .C1(n13224), .C2(n14150), .A(n11718), .B(n11717), .ZN(
        n11719) );
  OAI21_X1 U13576 ( .B1(n14168), .B2(n11839), .A(n11719), .ZN(P2_U3187) );
  OR2_X1 U13577 ( .A1(n13230), .A2(n14185), .ZN(n11720) );
  AOI22_X1 U13578 ( .A1(n11767), .A2(n12234), .B1(n13330), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n11723) );
  XNOR2_X1 U13579 ( .A(n14526), .B(n14184), .ZN(n13390) );
  NAND2_X1 U13580 ( .A1(n11725), .A2(n13390), .ZN(n11726) );
  NAND2_X1 U13581 ( .A1(n11805), .A2(n11726), .ZN(n11739) );
  OR2_X1 U13582 ( .A1(n11739), .A2(n16107), .ZN(n11738) );
  INV_X1 U13583 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n11727) );
  NAND2_X1 U13584 ( .A1(n11728), .A2(n11727), .ZN(n11729) );
  NAND2_X1 U13585 ( .A1(n11795), .A2(n11729), .ZN(n12411) );
  AOI22_X1 U13586 ( .A1(n13321), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13322), 
        .B2(P2_REG1_REG_17__SCAN_IN), .ZN(n11731) );
  NAND2_X1 U13587 ( .A1(n12336), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n11730) );
  OAI211_X1 U13588 ( .C1(n12411), .C2(n12314), .A(n11731), .B(n11730), .ZN(
        n14183) );
  AOI22_X1 U13589 ( .A1(n14183), .A2(n14139), .B1(n14137), .B2(n14185), .ZN(
        n11737) );
  INV_X1 U13590 ( .A(n14185), .ZN(n11851) );
  NOR2_X1 U13591 ( .A1(n13230), .A2(n11851), .ZN(n11732) );
  NAND2_X1 U13592 ( .A1(n13230), .A2(n11851), .ZN(n11734) );
  XNOR2_X1 U13593 ( .A(n13390), .B(n11789), .ZN(n11735) );
  NAND2_X1 U13594 ( .A1(n11735), .A2(n14393), .ZN(n11736) );
  INV_X1 U13595 ( .A(n11739), .ZN(n14530) );
  AOI21_X1 U13596 ( .B1(n14526), .B2(n11740), .A(n14416), .ZN(n11741) );
  NAND2_X1 U13597 ( .A1(n11741), .A2(n11806), .ZN(n14528) );
  INV_X1 U13598 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11742) );
  OAI22_X1 U13599 ( .A1(n14427), .A2(n11742), .B1(n11848), .B2(n14430), .ZN(
        n11743) );
  AOI21_X1 U13600 ( .B1(n14526), .B2(n14434), .A(n11743), .ZN(n11744) );
  OAI21_X1 U13601 ( .B1(n14528), .B2(n14420), .A(n11744), .ZN(n11745) );
  AOI21_X1 U13602 ( .B1(n14530), .B2(n11746), .A(n11745), .ZN(n11747) );
  OAI21_X1 U13603 ( .B1(n14532), .B2(n14378), .A(n11747), .ZN(P2_U3249) );
  INV_X1 U13604 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11751) );
  MUX2_X1 U13605 ( .A(n11752), .B(n11751), .S(n7178), .Z(n11975) );
  XNOR2_X1 U13606 ( .A(n11975), .B(SI_23_), .ZN(n11972) );
  XNOR2_X1 U13607 ( .A(n11974), .B(n11972), .ZN(n12283) );
  INV_X1 U13608 ( .A(n12283), .ZN(n11756) );
  NAND2_X1 U13609 ( .A1(n11753), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13406) );
  INV_X1 U13610 ( .A(n13406), .ZN(n13412) );
  AOI21_X1 U13611 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n14591), .A(n13412), 
        .ZN(n11754) );
  OAI21_X1 U13612 ( .B1(n11756), .B2(n14593), .A(n11754), .ZN(P2_U3304) );
  NAND2_X1 U13613 ( .A1(n15164), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11755) );
  OAI211_X1 U13614 ( .C1(n11756), .C2(n15167), .A(n13078), .B(n11755), .ZN(
        P1_U3332) );
  OAI222_X1 U13615 ( .A1(P3_U3151), .A2(n11758), .B1(n13083), .B2(n15301), 
        .C1(n13082), .C2(n11757), .ZN(P3_U3269) );
  INV_X1 U13616 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n11763) );
  XNOR2_X1 U13617 ( .A(n15467), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15463) );
  INV_X1 U13618 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n11762) );
  XNOR2_X1 U13619 ( .A(n15454), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n15450) );
  OAI21_X1 U13620 ( .B1(n10405), .B2(n11769), .A(n11759), .ZN(n11760) );
  NAND2_X1 U13621 ( .A1(n11770), .A2(n11760), .ZN(n11761) );
  XNOR2_X1 U13622 ( .A(n15442), .B(n11760), .ZN(n15439) );
  NAND2_X1 U13623 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n15439), .ZN(n15438) );
  NAND2_X1 U13624 ( .A1(n11761), .A2(n15438), .ZN(n15451) );
  NAND2_X1 U13625 ( .A1(n15450), .A2(n15451), .ZN(n15449) );
  OAI21_X1 U13626 ( .B1(n15454), .B2(n11762), .A(n15449), .ZN(n15462) );
  NAND2_X1 U13627 ( .A1(n15463), .A2(n15462), .ZN(n15461) );
  OAI21_X1 U13628 ( .B1(n15467), .B2(n11763), .A(n15461), .ZN(n14213) );
  XNOR2_X1 U13629 ( .A(n14213), .B(n11764), .ZN(n14215) );
  XNOR2_X1 U13630 ( .A(n14215), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n11783) );
  INV_X1 U13631 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n11765) );
  NAND2_X1 U13632 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14143)
         );
  OAI21_X1 U13633 ( .B1(n11766), .B2(n11765), .A(n14143), .ZN(n11781) );
  INV_X1 U13634 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n11774) );
  MUX2_X1 U13635 ( .A(n11774), .B(P2_REG2_REG_17__SCAN_IN), .S(n15467), .Z(
        n15456) );
  NAND2_X1 U13636 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n11767), .ZN(n11773) );
  MUX2_X1 U13637 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n11742), .S(n11767), .Z(
        n15444) );
  OAI21_X1 U13638 ( .B1(n11505), .B2(n11769), .A(n11768), .ZN(n11771) );
  NAND2_X1 U13639 ( .A1(n11770), .A2(n11771), .ZN(n11772) );
  XNOR2_X1 U13640 ( .A(n15442), .B(n11771), .ZN(n15434) );
  NAND2_X1 U13641 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n15434), .ZN(n15433) );
  NAND2_X1 U13642 ( .A1(n11772), .A2(n15433), .ZN(n15445) );
  NAND2_X1 U13643 ( .A1(n15444), .A2(n15445), .ZN(n15443) );
  NAND2_X1 U13644 ( .A1(n11773), .A2(n15443), .ZN(n15457) );
  NAND2_X1 U13645 ( .A1(n15456), .A2(n15457), .ZN(n15455) );
  OAI21_X1 U13646 ( .B1(n15467), .B2(n11774), .A(n15455), .ZN(n11775) );
  NOR2_X1 U13647 ( .A1(n11775), .A2(n14214), .ZN(n14220) );
  AOI21_X1 U13648 ( .B1(n14214), .B2(n11775), .A(n14220), .ZN(n11776) );
  INV_X1 U13649 ( .A(n11776), .ZN(n11777) );
  NOR2_X1 U13650 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n11777), .ZN(n14219) );
  AOI21_X1 U13651 ( .B1(n11777), .B2(P2_REG2_REG_18__SCAN_IN), .A(n14219), 
        .ZN(n11779) );
  NOR2_X1 U13652 ( .A1(n11779), .A2(n11778), .ZN(n11780) );
  AOI211_X1 U13653 ( .C1(n14205), .C2(n14214), .A(n11781), .B(n11780), .ZN(
        n11782) );
  OAI21_X1 U13654 ( .B1(n11783), .B2(n14230), .A(n11782), .ZN(P2_U3232) );
  OAI22_X1 U13655 ( .A1(n15467), .A2(n11785), .B1(n9957), .B2(n11784), .ZN(
        n11786) );
  INV_X1 U13656 ( .A(n11786), .ZN(n11787) );
  NAND2_X2 U13657 ( .A1(n11788), .A2(n11787), .ZN(n14577) );
  XNOR2_X1 U13658 ( .A(n14577), .B(n14183), .ZN(n13392) );
  INV_X1 U13659 ( .A(n14184), .ZN(n12414) );
  AND2_X1 U13660 ( .A1(n14526), .A2(n12414), .ZN(n11790) );
  OR2_X1 U13661 ( .A1(n14526), .A2(n12414), .ZN(n11791) );
  XNOR2_X1 U13662 ( .A(n13392), .B(n12226), .ZN(n11792) );
  OR2_X1 U13663 ( .A1(n11792), .A2(n14413), .ZN(n11803) );
  INV_X1 U13664 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n11794) );
  NAND2_X1 U13665 ( .A1(n11795), .A2(n11794), .ZN(n11796) );
  NAND2_X1 U13666 ( .A1(n12248), .A2(n11796), .ZN(n14414) );
  OR2_X1 U13667 ( .A1(n14414), .A2(n12314), .ZN(n11801) );
  INV_X1 U13668 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n14573) );
  NAND2_X1 U13669 ( .A1(n13322), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n11798) );
  NAND2_X1 U13670 ( .A1(n13321), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n11797) );
  OAI211_X1 U13671 ( .C1(n13325), .C2(n14573), .A(n11798), .B(n11797), .ZN(
        n11799) );
  INV_X1 U13672 ( .A(n11799), .ZN(n11800) );
  NAND2_X1 U13673 ( .A1(n11801), .A2(n11800), .ZN(n14182) );
  AOI22_X1 U13674 ( .A1(n14182), .A2(n14139), .B1(n14137), .B2(n14184), .ZN(
        n11802) );
  AND2_X1 U13675 ( .A1(n11803), .A2(n11802), .ZN(n14521) );
  NAND2_X1 U13676 ( .A1(n14526), .A2(n14184), .ZN(n11804) );
  XNOR2_X1 U13677 ( .A(n12354), .B(n13392), .ZN(n14519) );
  NAND2_X1 U13678 ( .A1(n14577), .A2(n11806), .ZN(n11807) );
  NAND3_X1 U13679 ( .A1(n14417), .A2(n14397), .A3(n11807), .ZN(n14520) );
  OAI22_X1 U13680 ( .A1(n14427), .A2(n11774), .B1(n12411), .B2(n14430), .ZN(
        n11808) );
  AOI21_X1 U13681 ( .B1(n14577), .B2(n14434), .A(n11808), .ZN(n11809) );
  OAI21_X1 U13682 ( .B1(n14520), .B2(n14420), .A(n11809), .ZN(n11810) );
  AOI21_X1 U13683 ( .B1(n14519), .B2(n14436), .A(n11810), .ZN(n11811) );
  OAI21_X1 U13684 ( .B1(n14378), .B2(n14521), .A(n11811), .ZN(P2_U3248) );
  INV_X1 U13685 ( .A(n11812), .ZN(n11816) );
  INV_X1 U13686 ( .A(n11813), .ZN(n11815) );
  AND2_X1 U13687 ( .A1(n12518), .A2(n14741), .ZN(n11817) );
  AOI21_X1 U13688 ( .B1(n12875), .B2(n12519), .A(n11817), .ZN(n11929) );
  AOI22_X1 U13689 ( .A1(n12875), .A2(n7181), .B1(n12519), .B2(n14741), .ZN(
        n11818) );
  XNOR2_X1 U13690 ( .A(n11818), .B(n12526), .ZN(n11928) );
  XOR2_X1 U13691 ( .A(n11929), .B(n11928), .Z(n11819) );
  OAI211_X1 U13692 ( .C1(n11820), .C2(n11819), .A(n11927), .B(n14719), .ZN(
        n11826) );
  OAI21_X1 U13693 ( .B1(n14725), .B2(n11822), .A(n11821), .ZN(n11823) );
  AOI21_X1 U13694 ( .B1(n14728), .B2(n11824), .A(n11823), .ZN(n11825) );
  OAI211_X1 U13695 ( .C1(n11827), .C2(n14731), .A(n11826), .B(n11825), .ZN(
        P1_U3224) );
  OAI222_X1 U13696 ( .A1(n13082), .A2(n11828), .B1(n13083), .B2(n15297), .C1(
        P3_U3151), .C2(n13664), .ZN(P3_U3268) );
  INV_X1 U13697 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n11832) );
  AOI211_X1 U13698 ( .C1(n16092), .C2(n11831), .A(n11830), .B(n11829), .ZN(
        n11834) );
  MUX2_X1 U13699 ( .A(n11832), .B(n11834), .S(n16142), .Z(n11833) );
  OAI21_X1 U13700 ( .B1(n11837), .B2(n14496), .A(n11833), .ZN(P2_U3514) );
  INV_X1 U13701 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n11835) );
  MUX2_X1 U13702 ( .A(n11835), .B(n11834), .S(n16146), .Z(n11836) );
  OAI21_X1 U13703 ( .B1(n11837), .B2(n14566), .A(n11836), .ZN(P2_U3475) );
  INV_X1 U13704 ( .A(n11838), .ZN(n11841) );
  XNOR2_X1 U13705 ( .A(n13230), .B(n14043), .ZN(n11843) );
  AND2_X1 U13706 ( .A1(n14185), .A2(n14416), .ZN(n11842) );
  NAND2_X1 U13707 ( .A1(n11843), .A2(n11842), .ZN(n11845) );
  OAI21_X1 U13708 ( .B1(n11843), .B2(n11842), .A(n11845), .ZN(n11922) );
  NOR2_X1 U13709 ( .A1(n14152), .A2(n11851), .ZN(n11844) );
  AOI22_X1 U13710 ( .A1(n7308), .A2(n14115), .B1(n11844), .B2(n11843), .ZN(
        n11856) );
  XNOR2_X1 U13711 ( .A(n14526), .B(n14032), .ZN(n12370) );
  NAND2_X1 U13712 ( .A1(n14184), .A2(n14416), .ZN(n12371) );
  XNOR2_X1 U13713 ( .A(n12370), .B(n12371), .ZN(n11847) );
  INV_X1 U13714 ( .A(n11847), .ZN(n11855) );
  INV_X1 U13715 ( .A(n11845), .ZN(n11846) );
  NAND2_X1 U13716 ( .A1(n12418), .A2(n14115), .ZN(n11854) );
  NAND2_X1 U13717 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n15447)
         );
  OAI21_X1 U13718 ( .B1(n14161), .B2(n11848), .A(n15447), .ZN(n11849) );
  AOI21_X1 U13719 ( .B1(n14099), .B2(n14183), .A(n11849), .ZN(n11850) );
  OAI21_X1 U13720 ( .B1(n11851), .B2(n14096), .A(n11850), .ZN(n11852) );
  AOI21_X1 U13721 ( .B1(n14526), .B2(n14150), .A(n11852), .ZN(n11853) );
  OAI211_X1 U13722 ( .C1(n11856), .C2(n11855), .A(n11854), .B(n11853), .ZN(
        P2_U3198) );
  XOR2_X1 U13723 ( .A(n12696), .B(n11857), .Z(n11858) );
  OAI222_X1 U13724 ( .A1(n15390), .A2(n15393), .B1(n15392), .B2(n11859), .C1(
        n11858), .C2(n13874), .ZN(n11941) );
  INV_X1 U13725 ( .A(n11941), .ZN(n11867) );
  OAI21_X1 U13726 ( .B1(n11861), .B2(n12696), .A(n11860), .ZN(n11942) );
  NOR2_X1 U13727 ( .A1(n13882), .A2(n11947), .ZN(n11865) );
  OAI22_X1 U13728 ( .A1(n15899), .A2(n11863), .B1(n11862), .B2(n15892), .ZN(
        n11864) );
  AOI211_X1 U13729 ( .C1(n11942), .C2(n13887), .A(n11865), .B(n11864), .ZN(
        n11866) );
  OAI21_X1 U13730 ( .B1(n11867), .B2(n13853), .A(n11866), .ZN(P3_U3222) );
  OAI211_X1 U13731 ( .C1(n11870), .C2(n11869), .A(n11868), .B(n13527), .ZN(
        n11875) );
  NAND2_X1 U13732 ( .A1(n13529), .A2(n13570), .ZN(n11871) );
  OAI211_X1 U13733 ( .C1(n13519), .C2(n11961), .A(n11872), .B(n11871), .ZN(
        n11873) );
  AOI21_X1 U13734 ( .B1(n13953), .B2(n13511), .A(n11873), .ZN(n11874) );
  OAI211_X1 U13735 ( .C1(n11876), .C2(n13531), .A(n11875), .B(n11874), .ZN(
        P3_U3157) );
  NAND2_X1 U13736 ( .A1(n11877), .A2(n13046), .ZN(n11879) );
  OR2_X1 U13737 ( .A1(n14656), .A2(n14737), .ZN(n11878) );
  NAND2_X1 U13738 ( .A1(n11879), .A2(n11878), .ZN(n11884) );
  INV_X1 U13739 ( .A(n11884), .ZN(n11885) );
  NAND2_X1 U13740 ( .A1(n11880), .A2(n12089), .ZN(n11883) );
  INV_X1 U13741 ( .A(n11910), .ZN(n11881) );
  AOI22_X1 U13742 ( .A1(n10053), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n12008), 
        .B2(n11881), .ZN(n11882) );
  INV_X1 U13743 ( .A(n14736), .ZN(n15004) );
  XNOR2_X1 U13744 ( .A(n14669), .B(n15004), .ZN(n13049) );
  INV_X1 U13745 ( .A(n13049), .ZN(n11902) );
  OAI21_X1 U13746 ( .B1(n11885), .B2(n13049), .A(n12154), .ZN(n15113) );
  INV_X1 U13747 ( .A(n15014), .ZN(n11886) );
  AOI211_X1 U13748 ( .C1(n14669), .C2(n11887), .A(n15952), .B(n11886), .ZN(
        n15109) );
  NAND2_X1 U13749 ( .A1(n15109), .A2(n14836), .ZN(n11897) );
  INV_X1 U13750 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n11888) );
  NAND2_X1 U13751 ( .A1(n11889), .A2(n11888), .ZN(n11890) );
  NAND2_X1 U13752 ( .A1(n12011), .A2(n11890), .ZN(n15017) );
  OR2_X1 U13753 ( .A1(n15017), .A2(n12142), .ZN(n11895) );
  INV_X1 U13754 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n15018) );
  NAND2_X1 U13755 ( .A1(n12987), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n11892) );
  NAND2_X1 U13756 ( .A1(n12014), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n11891) );
  OAI211_X1 U13757 ( .C1(n15018), .C2(n10239), .A(n11892), .B(n11891), .ZN(
        n11893) );
  INV_X1 U13758 ( .A(n11893), .ZN(n11894) );
  NAND2_X1 U13759 ( .A1(n11895), .A2(n11894), .ZN(n14735) );
  AND2_X1 U13760 ( .A1(n14737), .A2(n14978), .ZN(n11896) );
  AOI21_X1 U13761 ( .B1(n14735), .B2(n14980), .A(n11896), .ZN(n15108) );
  OAI211_X1 U13762 ( .C1(n15016), .C2(n14667), .A(n11897), .B(n15108), .ZN(
        n11900) );
  OAI22_X1 U13763 ( .A1(n7604), .A2(n16041), .B1(n11907), .B2(n11899), .ZN(
        n11898) );
  AOI21_X1 U13764 ( .B1(n11900), .B2(n11899), .A(n11898), .ZN(n11905) );
  NAND2_X1 U13765 ( .A1(n11903), .A2(n11902), .ZN(n12003) );
  OAI21_X1 U13766 ( .B1(n11903), .B2(n11902), .A(n12003), .ZN(n15111) );
  NAND2_X1 U13767 ( .A1(n15111), .A2(n14910), .ZN(n11904) );
  OAI211_X1 U13768 ( .C1(n15113), .C2(n14967), .A(n11905), .B(n11904), .ZN(
        P1_U3276) );
  INV_X1 U13769 ( .A(n14824), .ZN(n11917) );
  OAI21_X1 U13770 ( .B1(n11907), .B2(n11910), .A(n11906), .ZN(n14823) );
  XOR2_X1 U13771 ( .A(n14823), .B(n14824), .Z(n11908) );
  NAND2_X1 U13772 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n11908), .ZN(n14826) );
  OAI211_X1 U13773 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n11908), .A(n14833), 
        .B(n14826), .ZN(n11916) );
  NAND2_X1 U13774 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14704)
         );
  OAI21_X1 U13775 ( .B1(n11911), .B2(n11910), .A(n11909), .ZN(n14819) );
  XNOR2_X1 U13776 ( .A(n14819), .B(n11917), .ZN(n11912) );
  NAND2_X1 U13777 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n11912), .ZN(n14821) );
  OAI211_X1 U13778 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n11912), .A(n14834), 
        .B(n14821), .ZN(n11913) );
  NAND2_X1 U13779 ( .A1(n14704), .A2(n11913), .ZN(n11914) );
  AOI21_X1 U13780 ( .B1(n14797), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n11914), 
        .ZN(n11915) );
  OAI211_X1 U13781 ( .C1(n14828), .C2(n11917), .A(n11916), .B(n11915), .ZN(
        P1_U3261) );
  NAND2_X1 U13782 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n15436)
         );
  INV_X1 U13783 ( .A(n11918), .ZN(n11919) );
  NAND2_X1 U13784 ( .A1(n14141), .A2(n11919), .ZN(n11920) );
  OAI211_X1 U13785 ( .C1(n14144), .C2(n11921), .A(n15436), .B(n11920), .ZN(
        n11925) );
  AOI211_X1 U13786 ( .C1(n11923), .C2(n11922), .A(n14168), .B(n7308), .ZN(
        n11924) );
  AOI211_X1 U13787 ( .C1(n13230), .C2(n14150), .A(n11925), .B(n11924), .ZN(
        n11926) );
  INV_X1 U13788 ( .A(n11926), .ZN(P2_U3213) );
  AND2_X1 U13789 ( .A1(n12518), .A2(n14740), .ZN(n11930) );
  AOI21_X1 U13790 ( .B1(n12885), .B2(n12519), .A(n11930), .ZN(n12429) );
  AOI22_X1 U13791 ( .A1(n12885), .A2(n12514), .B1(n12519), .B2(n14740), .ZN(
        n11931) );
  XNOR2_X1 U13792 ( .A(n11931), .B(n12526), .ZN(n12428) );
  XOR2_X1 U13793 ( .A(n12429), .B(n12428), .Z(n11932) );
  OAI211_X1 U13794 ( .C1(n11933), .C2(n11932), .A(n16121), .B(n14719), .ZN(
        n11939) );
  OAI21_X1 U13795 ( .B1(n14725), .B2(n11935), .A(n11934), .ZN(n11936) );
  AOI21_X1 U13796 ( .B1(n14728), .B2(n11937), .A(n11936), .ZN(n11938) );
  OAI211_X1 U13797 ( .C1(n11940), .C2(n14731), .A(n11939), .B(n11938), .ZN(
        P1_U3234) );
  INV_X1 U13798 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n11943) );
  AOI21_X1 U13799 ( .B1(n13955), .B2(n11942), .A(n11941), .ZN(n11945) );
  MUX2_X1 U13800 ( .A(n11943), .B(n11945), .S(n16104), .Z(n11944) );
  OAI21_X1 U13801 ( .B1(n16159), .B2(n11947), .A(n11944), .ZN(P3_U3423) );
  MUX2_X1 U13802 ( .A(n8487), .B(n11945), .S(n16101), .Z(n11946) );
  OAI21_X1 U13803 ( .B1(n16154), .B2(n11947), .A(n11946), .ZN(P3_U3470) );
  NAND2_X1 U13804 ( .A1(n11949), .A2(n11948), .ZN(n11950) );
  XNOR2_X1 U13805 ( .A(n11951), .B(n11950), .ZN(n11956) );
  NAND2_X1 U13806 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(P3_U3151), .ZN(n15712)
         );
  OAI21_X1 U13807 ( .B1(n13519), .B2(n13876), .A(n15712), .ZN(n11953) );
  NOR2_X1 U13808 ( .A1(n13531), .A2(n11965), .ZN(n11952) );
  AOI211_X1 U13809 ( .C1(n13529), .C2(n13568), .A(n11953), .B(n11952), .ZN(
        n11955) );
  NAND2_X1 U13810 ( .A1(n13511), .A2(n11968), .ZN(n11954) );
  OAI211_X1 U13811 ( .C1(n11956), .C2(n13539), .A(n11955), .B(n11954), .ZN(
        P3_U3164) );
  OR2_X1 U13812 ( .A1(n11957), .A2(n12609), .ZN(n11958) );
  NAND2_X1 U13813 ( .A1(n11959), .A2(n11958), .ZN(n16081) );
  INV_X1 U13814 ( .A(n16081), .ZN(n11971) );
  XOR2_X1 U13815 ( .A(n12609), .B(n11960), .Z(n11964) );
  OAI22_X1 U13816 ( .A1(n11961), .A2(n15392), .B1(n13876), .B2(n15390), .ZN(
        n11962) );
  AOI21_X1 U13817 ( .B1(n16081), .B2(n13754), .A(n11962), .ZN(n11963) );
  OAI21_X1 U13818 ( .B1(n11964), .B2(n13874), .A(n11963), .ZN(n16079) );
  NAND2_X1 U13819 ( .A1(n16079), .A2(n15899), .ZN(n11970) );
  OAI22_X1 U13820 ( .A1(n15899), .A2(n11966), .B1(n11965), .B2(n15892), .ZN(
        n11967) );
  AOI21_X1 U13821 ( .B1(n11968), .B2(n15399), .A(n11967), .ZN(n11969) );
  OAI211_X1 U13822 ( .C1(n11971), .C2(n15402), .A(n11970), .B(n11969), .ZN(
        P3_U3221) );
  INV_X1 U13823 ( .A(n11972), .ZN(n11973) );
  INV_X1 U13824 ( .A(n11975), .ZN(n11976) );
  NAND2_X1 U13825 ( .A1(n11976), .A2(SI_23_), .ZN(n11977) );
  INV_X1 U13826 ( .A(n12073), .ZN(n11978) );
  MUX2_X1 U13827 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n7178), .Z(n12072) );
  NAND2_X1 U13828 ( .A1(n11979), .A2(SI_24_), .ZN(n11980) );
  MUX2_X1 U13829 ( .A(n14600), .B(n15163), .S(n7178), .Z(n11983) );
  NAND2_X1 U13830 ( .A1(n11983), .A2(n11982), .ZN(n11986) );
  INV_X1 U13831 ( .A(n11983), .ZN(n11984) );
  NAND2_X1 U13832 ( .A1(n11984), .A2(SI_25_), .ZN(n11985) );
  NAND2_X1 U13833 ( .A1(n11986), .A2(n11985), .ZN(n12087) );
  MUX2_X1 U13834 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n7178), .Z(n11987) );
  XNOR2_X1 U13835 ( .A(n11987), .B(n15301), .ZN(n12105) );
  NAND2_X1 U13836 ( .A1(n11987), .A2(SI_26_), .ZN(n12121) );
  NAND2_X1 U13837 ( .A1(n12178), .A2(n12121), .ZN(n11989) );
  MUX2_X1 U13838 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n7178), .Z(n12120) );
  XNOR2_X1 U13839 ( .A(n12120), .B(n15297), .ZN(n12123) );
  INV_X1 U13840 ( .A(n12123), .ZN(n11988) );
  NAND2_X1 U13841 ( .A1(n13011), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n11990) );
  NAND2_X2 U13842 ( .A1(n11991), .A2(n11990), .ZN(n14871) );
  INV_X1 U13843 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n12025) );
  NAND2_X1 U13844 ( .A1(n12024), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n12051) );
  INV_X1 U13845 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n12050) );
  INV_X1 U13846 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n12076) );
  INV_X1 U13847 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n12092) );
  INV_X1 U13848 ( .A(n12109), .ZN(n11993) );
  NAND2_X1 U13849 ( .A1(n11993), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n12111) );
  INV_X1 U13850 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n11994) );
  NAND2_X1 U13851 ( .A1(n12111), .A2(n11994), .ZN(n11995) );
  NAND2_X1 U13852 ( .A1(n14870), .A2(n12095), .ZN(n12001) );
  INV_X1 U13853 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n11998) );
  NAND2_X1 U13854 ( .A1(n12987), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n11997) );
  NAND2_X1 U13855 ( .A1(n12988), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n11996) );
  OAI211_X1 U13856 ( .C1(n11998), .C2(n12992), .A(n11997), .B(n11996), .ZN(
        n11999) );
  INV_X1 U13857 ( .A(n11999), .ZN(n12000) );
  NAND2_X1 U13858 ( .A1(n14669), .A2(n15004), .ZN(n12002) );
  NAND2_X1 U13859 ( .A1(n12228), .A2(n12089), .ZN(n12005) );
  AOI22_X1 U13860 ( .A1(n13011), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n12008), 
        .B2(n14824), .ZN(n12004) );
  INV_X1 U13861 ( .A(n14735), .ZN(n12006) );
  XNOR2_X1 U13862 ( .A(n15104), .B(n12006), .ZN(n15010) );
  OR2_X1 U13863 ( .A1(n15104), .A2(n12006), .ZN(n12007) );
  NAND2_X1 U13864 ( .A1(n12233), .A2(n12089), .ZN(n12010) );
  AOI22_X1 U13865 ( .A1(n10053), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n13059), 
        .B2(n12008), .ZN(n12009) );
  NAND2_X1 U13866 ( .A1(n12011), .A2(n14626), .ZN(n12012) );
  NAND2_X1 U13867 ( .A1(n12026), .A2(n12012), .ZN(n14993) );
  INV_X1 U13868 ( .A(n14993), .ZN(n12013) );
  NAND2_X1 U13869 ( .A1(n12013), .A2(n12095), .ZN(n12020) );
  INV_X1 U13870 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n12017) );
  NAND2_X1 U13871 ( .A1(n12987), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n12016) );
  NAND2_X1 U13872 ( .A1(n12014), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n12015) );
  OAI211_X1 U13873 ( .C1(n10239), .C2(n12017), .A(n12016), .B(n12015), .ZN(
        n12018) );
  INV_X1 U13874 ( .A(n12018), .ZN(n12019) );
  XNOR2_X1 U13875 ( .A(n14995), .B(n15006), .ZN(n13050) );
  NAND2_X1 U13876 ( .A1(n12244), .A2(n12089), .ZN(n12023) );
  NAND2_X1 U13877 ( .A1(n13011), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n12022) );
  INV_X1 U13878 ( .A(n12024), .ZN(n12039) );
  NAND2_X1 U13879 ( .A1(n12026), .A2(n12025), .ZN(n12027) );
  NAND2_X1 U13880 ( .A1(n14982), .A2(n12095), .ZN(n12033) );
  INV_X1 U13881 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n12030) );
  NAND2_X1 U13882 ( .A1(n12987), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n12029) );
  NAND2_X1 U13883 ( .A1(n12988), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n12028) );
  OAI211_X1 U13884 ( .C1(n12992), .C2(n12030), .A(n12029), .B(n12028), .ZN(
        n12031) );
  INV_X1 U13885 ( .A(n12031), .ZN(n12032) );
  NAND2_X1 U13886 ( .A1(n15086), .A2(n14637), .ZN(n12034) );
  NAND2_X1 U13887 ( .A1(n12035), .A2(n12034), .ZN(n13047) );
  NAND2_X1 U13888 ( .A1(n14971), .A2(n12035), .ZN(n14959) );
  NAND2_X1 U13889 ( .A1(n12259), .A2(n12089), .ZN(n12037) );
  NAND2_X1 U13890 ( .A1(n13011), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n12036) );
  NAND2_X2 U13891 ( .A1(n12037), .A2(n12036), .ZN(n15082) );
  INV_X1 U13892 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n12038) );
  NAND2_X1 U13893 ( .A1(n12039), .A2(n12038), .ZN(n12040) );
  NAND2_X1 U13894 ( .A1(n12051), .A2(n12040), .ZN(n14635) );
  OR2_X1 U13895 ( .A1(n14635), .A2(n12142), .ZN(n12046) );
  INV_X1 U13896 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n12043) );
  NAND2_X1 U13897 ( .A1(n12987), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n12042) );
  NAND2_X1 U13898 ( .A1(n12988), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n12041) );
  OAI211_X1 U13899 ( .C1(n12043), .C2(n12992), .A(n12042), .B(n12041), .ZN(
        n12044) );
  INV_X1 U13900 ( .A(n12044), .ZN(n12045) );
  XNOR2_X1 U13901 ( .A(n15082), .B(n14981), .ZN(n14966) );
  INV_X1 U13902 ( .A(n14981), .ZN(n12914) );
  NAND2_X1 U13903 ( .A1(n12047), .A2(n7178), .ZN(n12048) );
  NAND2_X1 U13904 ( .A1(n12051), .A2(n12050), .ZN(n12052) );
  AND2_X1 U13905 ( .A1(n12063), .A2(n12052), .ZN(n14954) );
  NAND2_X1 U13906 ( .A1(n14954), .A2(n12095), .ZN(n12058) );
  INV_X1 U13907 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n12055) );
  NAND2_X1 U13908 ( .A1(n9339), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n12054) );
  NAND2_X1 U13909 ( .A1(n12988), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n12053) );
  OAI211_X1 U13910 ( .C1(n12055), .C2(n12992), .A(n12054), .B(n12053), .ZN(
        n12056) );
  INV_X1 U13911 ( .A(n12056), .ZN(n12057) );
  NAND2_X1 U13912 ( .A1(n15075), .A2(n12911), .ZN(n12158) );
  OR2_X1 U13913 ( .A1(n15075), .A2(n12911), .ZN(n12059) );
  NAND2_X1 U13914 ( .A1(n12158), .A2(n12059), .ZN(n13052) );
  NAND2_X1 U13915 ( .A1(n12283), .A2(n12089), .ZN(n12061) );
  NAND2_X1 U13916 ( .A1(n13011), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12060) );
  INV_X1 U13917 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n12062) );
  NAND2_X1 U13918 ( .A1(n12063), .A2(n12062), .ZN(n12064) );
  NAND2_X1 U13919 ( .A1(n12077), .A2(n12064), .ZN(n14616) );
  OR2_X1 U13920 ( .A1(n14616), .A2(n12142), .ZN(n12070) );
  INV_X1 U13921 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n12067) );
  NAND2_X1 U13922 ( .A1(n12987), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n12066) );
  NAND2_X1 U13923 ( .A1(n12988), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n12065) );
  OAI211_X1 U13924 ( .C1(n12067), .C2(n12992), .A(n12066), .B(n12065), .ZN(
        n12068) );
  INV_X1 U13925 ( .A(n12068), .ZN(n12069) );
  XNOR2_X1 U13926 ( .A(n15069), .B(n14951), .ZN(n14939) );
  INV_X1 U13927 ( .A(n14951), .ZN(n14913) );
  NAND2_X1 U13928 ( .A1(n15069), .A2(n14913), .ZN(n12071) );
  NAND2_X1 U13929 ( .A1(n14601), .A2(n12089), .ZN(n12075) );
  NAND2_X1 U13930 ( .A1(n10053), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12074) );
  NAND2_X1 U13931 ( .A1(n12077), .A2(n12076), .ZN(n12078) );
  AND2_X1 U13932 ( .A1(n12093), .A2(n12078), .ZN(n14923) );
  NAND2_X1 U13933 ( .A1(n14923), .A2(n12095), .ZN(n12084) );
  INV_X1 U13934 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n12081) );
  NAND2_X1 U13935 ( .A1(n9339), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n12080) );
  NAND2_X1 U13936 ( .A1(n12988), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n12079) );
  OAI211_X1 U13937 ( .C1(n12081), .C2(n12992), .A(n12080), .B(n12079), .ZN(
        n12082) );
  INV_X1 U13938 ( .A(n12082), .ZN(n12083) );
  INV_X1 U13939 ( .A(n14900), .ZN(n12085) );
  OR2_X1 U13940 ( .A1(n15064), .A2(n12085), .ZN(n12086) );
  NAND2_X1 U13941 ( .A1(n14598), .A2(n12089), .ZN(n12091) );
  NAND2_X1 U13942 ( .A1(n13011), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12090) );
  NAND2_X2 U13943 ( .A1(n12091), .A2(n12090), .ZN(n15057) );
  NAND2_X1 U13944 ( .A1(n12093), .A2(n12092), .ZN(n12094) );
  AND2_X1 U13945 ( .A1(n12109), .A2(n12094), .ZN(n14903) );
  NAND2_X1 U13946 ( .A1(n14903), .A2(n12095), .ZN(n12101) );
  INV_X1 U13947 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n12098) );
  NAND2_X1 U13948 ( .A1(n12987), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n12097) );
  NAND2_X1 U13949 ( .A1(n12988), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n12096) );
  OAI211_X1 U13950 ( .C1(n12992), .C2(n12098), .A(n12097), .B(n12096), .ZN(
        n12099) );
  INV_X1 U13951 ( .A(n12099), .ZN(n12100) );
  NAND2_X1 U13952 ( .A1(n15057), .A2(n14914), .ZN(n12104) );
  NAND2_X1 U13953 ( .A1(n12104), .A2(n12102), .ZN(n14894) );
  XNOR2_X1 U13954 ( .A(n12106), .B(n12105), .ZN(n14594) );
  NAND2_X1 U13955 ( .A1(n10053), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n12107) );
  INV_X1 U13956 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n12108) );
  NAND2_X1 U13957 ( .A1(n12109), .A2(n12108), .ZN(n12110) );
  NAND2_X1 U13958 ( .A1(n12111), .A2(n12110), .ZN(n14712) );
  OR2_X1 U13959 ( .A1(n14712), .A2(n12142), .ZN(n12117) );
  INV_X1 U13960 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n12114) );
  NAND2_X1 U13961 ( .A1(n12987), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n12113) );
  NAND2_X1 U13962 ( .A1(n12988), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n12112) );
  OAI211_X1 U13963 ( .C1(n12992), .C2(n12114), .A(n12113), .B(n12112), .ZN(
        n12115) );
  INV_X1 U13964 ( .A(n12115), .ZN(n12116) );
  NAND2_X1 U13965 ( .A1(n15051), .A2(n14859), .ZN(n12119) );
  OR2_X1 U13966 ( .A1(n15051), .A2(n14859), .ZN(n12118) );
  NAND2_X1 U13967 ( .A1(n12119), .A2(n12118), .ZN(n14876) );
  INV_X1 U13968 ( .A(n14876), .ZN(n14880) );
  NAND2_X1 U13969 ( .A1(n12120), .A2(SI_27_), .ZN(n12122) );
  AND2_X1 U13970 ( .A1(n12121), .A2(n12122), .ZN(n12176) );
  INV_X1 U13971 ( .A(n12122), .ZN(n12124) );
  OR2_X1 U13972 ( .A1(n12124), .A2(n12123), .ZN(n12179) );
  MUX2_X1 U13973 ( .A(n12125), .B(n15153), .S(n7178), .Z(n12126) );
  NAND2_X1 U13974 ( .A1(n12126), .A2(n15293), .ZN(n12182) );
  INV_X1 U13975 ( .A(n12126), .ZN(n12127) );
  NAND2_X1 U13976 ( .A1(n12127), .A2(SI_28_), .ZN(n12128) );
  NAND2_X1 U13977 ( .A1(n12182), .A2(n12128), .ZN(n12180) );
  NAND2_X1 U13978 ( .A1(n14589), .A2(n12089), .ZN(n12131) );
  NAND2_X1 U13979 ( .A1(n10053), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12130) );
  INV_X1 U13980 ( .A(n12134), .ZN(n12132) );
  NAND2_X1 U13981 ( .A1(n12132), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n12553) );
  INV_X1 U13982 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n12133) );
  NAND2_X1 U13983 ( .A1(n12134), .A2(n12133), .ZN(n12135) );
  NAND2_X1 U13984 ( .A1(n12553), .A2(n12135), .ZN(n12168) );
  INV_X1 U13985 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n12138) );
  NAND2_X1 U13986 ( .A1(n9339), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n12137) );
  NAND2_X1 U13987 ( .A1(n12988), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n12136) );
  OAI211_X1 U13988 ( .C1(n12138), .C2(n12992), .A(n12137), .B(n12136), .ZN(
        n12139) );
  INV_X1 U13989 ( .A(n12139), .ZN(n12140) );
  XNOR2_X1 U13990 ( .A(n15040), .B(n14857), .ZN(n13055) );
  OR2_X1 U13991 ( .A1(n12553), .A2(n12142), .ZN(n12148) );
  INV_X1 U13992 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n12145) );
  NAND2_X1 U13993 ( .A1(n12987), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n12144) );
  NAND2_X1 U13994 ( .A1(n12988), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n12143) );
  OAI211_X1 U13995 ( .C1(n12145), .C2(n12992), .A(n12144), .B(n12143), .ZN(
        n12146) );
  INV_X1 U13996 ( .A(n12146), .ZN(n12147) );
  NAND2_X1 U13997 ( .A1(n12148), .A2(n12147), .ZN(n14734) );
  NAND2_X1 U13998 ( .A1(n14734), .A2(n14980), .ZN(n12150) );
  NAND2_X1 U13999 ( .A1(n14882), .A2(n14978), .ZN(n12149) );
  NAND2_X1 U14000 ( .A1(n14669), .A2(n14736), .ZN(n12153) );
  OR2_X1 U14001 ( .A1(n15104), .A2(n14735), .ZN(n12155) );
  NAND2_X1 U14002 ( .A1(n15104), .A2(n14735), .ZN(n12156) );
  OR2_X1 U14003 ( .A1(n14976), .A2(n14637), .ZN(n12157) );
  NAND2_X1 U14004 ( .A1(n14946), .A2(n12158), .ZN(n14940) );
  NAND2_X1 U14005 ( .A1(n15069), .A2(n14951), .ZN(n12159) );
  OR2_X1 U14006 ( .A1(n15064), .A2(n14900), .ZN(n12160) );
  NAND2_X1 U14007 ( .A1(n14877), .A2(n14876), .ZN(n12162) );
  NAND2_X1 U14008 ( .A1(n15051), .A2(n14899), .ZN(n12161) );
  OR2_X1 U14009 ( .A1(n15069), .A2(n14949), .ZN(n14934) );
  INV_X1 U14010 ( .A(n7185), .ZN(n12166) );
  INV_X1 U14011 ( .A(n12543), .ZN(n12165) );
  AOI21_X1 U14012 ( .B1(n15040), .B2(n12166), .A(n12165), .ZN(n15042) );
  NOR2_X1 U14013 ( .A1(n12167), .A2(n14952), .ZN(n14843) );
  NAND2_X1 U14014 ( .A1(n15042), .A2(n14843), .ZN(n12170) );
  INV_X1 U14015 ( .A(n12168), .ZN(n12531) );
  AOI22_X1 U14016 ( .A1(n12531), .A2(n16037), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n15998), .ZN(n12169) );
  OAI211_X1 U14017 ( .C1(n12555), .C2(n16041), .A(n12170), .B(n12169), .ZN(
        n12171) );
  AOI21_X1 U14018 ( .B1(n15039), .B2(n12172), .A(n12171), .ZN(n12173) );
  OAI21_X1 U14019 ( .B1(n15044), .B2(n15998), .A(n12173), .ZN(P1_U3265) );
  INV_X1 U14020 ( .A(n12174), .ZN(n12192) );
  INV_X1 U14021 ( .A(n12180), .ZN(n12175) );
  AND2_X1 U14022 ( .A1(n12176), .A2(n12175), .ZN(n12177) );
  NAND2_X1 U14023 ( .A1(n12178), .A2(n12177), .ZN(n12181) );
  INV_X1 U14024 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15148) );
  MUX2_X1 U14025 ( .A(n14587), .B(n15148), .S(n7178), .Z(n12183) );
  XNOR2_X1 U14026 ( .A(n12183), .B(SI_29_), .ZN(n12331) );
  NAND2_X1 U14027 ( .A1(n12183), .A2(n15289), .ZN(n12184) );
  MUX2_X1 U14028 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n7178), .Z(n12185) );
  NAND2_X1 U14029 ( .A1(n12185), .A2(SI_30_), .ZN(n13005) );
  INV_X1 U14030 ( .A(n12185), .ZN(n12186) );
  INV_X1 U14031 ( .A(SI_30_), .ZN(n15290) );
  NAND2_X1 U14032 ( .A1(n12186), .A2(n15290), .ZN(n12187) );
  NAND2_X1 U14033 ( .A1(n13005), .A2(n12187), .ZN(n12188) );
  NAND2_X1 U14034 ( .A1(n12189), .A2(n12188), .ZN(n12190) );
  INV_X1 U14035 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12191) );
  OAI222_X1 U14036 ( .A1(n12192), .A2(P2_U3088), .B1(n14593), .B2(n13318), 
        .C1(n12191), .C2(n14588), .ZN(P2_U3297) );
  OAI222_X1 U14037 ( .A1(n13082), .A2(n12194), .B1(n13083), .B2(n15293), .C1(
        P3_U3151), .C2(n12193), .ZN(P3_U3267) );
  INV_X1 U14038 ( .A(n12195), .ZN(n12196) );
  NAND2_X1 U14039 ( .A1(n12197), .A2(n15899), .ZN(n12202) );
  NOR2_X1 U14040 ( .A1(n12198), .A2(n15892), .ZN(n13671) );
  NOR2_X1 U14041 ( .A1(n12199), .A2(n13882), .ZN(n12200) );
  AOI211_X1 U14042 ( .C1(n13853), .C2(P3_REG2_REG_29__SCAN_IN), .A(n13671), 
        .B(n12200), .ZN(n12201) );
  OAI211_X1 U14043 ( .C1(n12203), .C2(n13868), .A(n12202), .B(n12201), .ZN(
        P3_U3204) );
  NAND2_X1 U14044 ( .A1(n13330), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n12204) );
  NAND2_X2 U14045 ( .A1(n12205), .A2(n12204), .ZN(n14277) );
  INV_X1 U14046 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n14132) );
  INV_X1 U14047 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n12247) );
  INV_X1 U14048 ( .A(n12262), .ZN(n12206) );
  INV_X1 U14049 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n12394) );
  INV_X1 U14050 ( .A(n12287), .ZN(n12207) );
  INV_X1 U14051 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n14119) );
  INV_X1 U14052 ( .A(n12300), .ZN(n12208) );
  NAND2_X1 U14053 ( .A1(n12208), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n12219) );
  INV_X1 U14054 ( .A(n12219), .ZN(n12209) );
  NAND2_X1 U14055 ( .A1(n12209), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n12312) );
  INV_X1 U14056 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n14160) );
  NAND2_X1 U14057 ( .A1(n12219), .A2(n14160), .ZN(n12210) );
  NAND2_X1 U14058 ( .A1(n12312), .A2(n12210), .ZN(n14278) );
  OR2_X1 U14059 ( .A1(n14278), .A2(n12314), .ZN(n12215) );
  INV_X1 U14060 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n14549) );
  NAND2_X1 U14061 ( .A1(n13321), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n12212) );
  NAND2_X1 U14062 ( .A1(n13322), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n12211) );
  OAI211_X1 U14063 ( .C1(n14549), .C2(n13325), .A(n12212), .B(n12211), .ZN(
        n12213) );
  INV_X1 U14064 ( .A(n12213), .ZN(n12214) );
  NAND2_X1 U14065 ( .A1(n12215), .A2(n12214), .ZN(n14174) );
  INV_X1 U14066 ( .A(n14174), .ZN(n13311) );
  XNOR2_X1 U14067 ( .A(n14277), .B(n13311), .ZN(n14282) );
  INV_X1 U14068 ( .A(n14282), .ZN(n12363) );
  NAND2_X1 U14069 ( .A1(n13330), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12216) );
  NAND2_X2 U14070 ( .A1(n12217), .A2(n12216), .ZN(n14470) );
  INV_X1 U14071 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n14111) );
  NAND2_X1 U14072 ( .A1(n12300), .A2(n14111), .ZN(n12218) );
  NAND2_X1 U14073 ( .A1(n12219), .A2(n12218), .ZN(n14296) );
  OR2_X1 U14074 ( .A1(n14296), .A2(n12314), .ZN(n12225) );
  INV_X1 U14075 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n12222) );
  NAND2_X1 U14076 ( .A1(n13321), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n12221) );
  NAND2_X1 U14077 ( .A1(n12345), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n12220) );
  OAI211_X1 U14078 ( .C1(n12222), .C2(n13325), .A(n12221), .B(n12220), .ZN(
        n12223) );
  INV_X1 U14079 ( .A(n12223), .ZN(n12224) );
  NAND2_X1 U14080 ( .A1(n12225), .A2(n12224), .ZN(n14175) );
  XNOR2_X1 U14081 ( .A(n14470), .B(n14158), .ZN(n13398) );
  INV_X1 U14082 ( .A(n14183), .ZN(n12227) );
  AOI22_X1 U14083 ( .A1(n13330), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n12234), 
        .B2(n14214), .ZN(n12229) );
  INV_X1 U14084 ( .A(n14182), .ZN(n12231) );
  XNOR2_X1 U14085 ( .A(n14511), .B(n12231), .ZN(n14408) );
  NAND2_X1 U14086 ( .A1(n14511), .A2(n12231), .ZN(n12232) );
  AOI22_X1 U14087 ( .A1(n9883), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7183), 
        .B2(n12234), .ZN(n12235) );
  NAND2_X2 U14088 ( .A1(n12236), .A2(n12235), .ZN(n14570) );
  XNOR2_X1 U14089 ( .A(n12248), .B(P2_REG3_REG_19__SCAN_IN), .ZN(n14386) );
  NAND2_X1 U14090 ( .A1(n14386), .A2(n12342), .ZN(n12242) );
  INV_X1 U14091 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n14388) );
  NAND2_X1 U14092 ( .A1(n12336), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n12238) );
  NAND2_X1 U14093 ( .A1(n13322), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n12237) );
  OAI211_X1 U14094 ( .C1(n12239), .C2(n14388), .A(n12238), .B(n12237), .ZN(
        n12240) );
  INV_X1 U14095 ( .A(n12240), .ZN(n12241) );
  NAND2_X1 U14096 ( .A1(n12242), .A2(n12241), .ZN(n14181) );
  INV_X1 U14097 ( .A(n14181), .ZN(n14124) );
  XNOR2_X1 U14098 ( .A(n14570), .B(n14124), .ZN(n14390) );
  OR2_X1 U14099 ( .A1(n14570), .A2(n14124), .ZN(n12243) );
  NAND2_X1 U14100 ( .A1(n9883), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n12245) );
  OAI21_X1 U14101 ( .B1(n12248), .B2(n12247), .A(n14132), .ZN(n12249) );
  AND2_X1 U14102 ( .A1(n12249), .A2(n12262), .ZN(n14377) );
  NAND2_X1 U14103 ( .A1(n14377), .A2(n12342), .ZN(n12255) );
  INV_X1 U14104 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n12252) );
  NAND2_X1 U14105 ( .A1(n13322), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n12251) );
  NAND2_X1 U14106 ( .A1(n13321), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n12250) );
  OAI211_X1 U14107 ( .C1(n12252), .C2(n13325), .A(n12251), .B(n12250), .ZN(
        n12253) );
  INV_X1 U14108 ( .A(n12253), .ZN(n12254) );
  NAND2_X1 U14109 ( .A1(n12255), .A2(n12254), .ZN(n14180) );
  NAND2_X1 U14110 ( .A1(n14502), .A2(n14353), .ZN(n12256) );
  NAND2_X1 U14111 ( .A1(n14370), .A2(n12256), .ZN(n12258) );
  OR2_X1 U14112 ( .A1(n14502), .A2(n14353), .ZN(n12257) );
  NAND2_X1 U14113 ( .A1(n12258), .A2(n12257), .ZN(n14351) );
  NAND2_X1 U14114 ( .A1(n9883), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n12260) );
  INV_X1 U14115 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n14095) );
  NAND2_X1 U14116 ( .A1(n12262), .A2(n14095), .ZN(n12263) );
  NAND2_X1 U14117 ( .A1(n12274), .A2(n12263), .ZN(n14362) );
  OR2_X1 U14118 ( .A1(n14362), .A2(n12314), .ZN(n12268) );
  INV_X1 U14119 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n14560) );
  NAND2_X1 U14120 ( .A1(n12345), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n12265) );
  NAND2_X1 U14121 ( .A1(n13321), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n12264) );
  OAI211_X1 U14122 ( .C1(n14560), .C2(n13325), .A(n12265), .B(n12264), .ZN(
        n12266) );
  INV_X1 U14123 ( .A(n12266), .ZN(n12267) );
  NAND2_X1 U14124 ( .A1(n12268), .A2(n12267), .ZN(n14179) );
  INV_X1 U14125 ( .A(n14179), .ZN(n12269) );
  XNOR2_X1 U14126 ( .A(n14361), .B(n12269), .ZN(n14357) );
  INV_X1 U14127 ( .A(n14357), .ZN(n14350) );
  OR2_X1 U14128 ( .A1(n14361), .A2(n12269), .ZN(n12270) );
  NAND2_X1 U14129 ( .A1(n9883), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n12272) );
  NAND2_X1 U14130 ( .A1(n12274), .A2(n12394), .ZN(n12275) );
  NAND2_X1 U14131 ( .A1(n12287), .A2(n12275), .ZN(n14337) );
  OR2_X1 U14132 ( .A1(n14337), .A2(n12314), .ZN(n12280) );
  INV_X1 U14133 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n14556) );
  NAND2_X1 U14134 ( .A1(n12345), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n12277) );
  NAND2_X1 U14135 ( .A1(n13321), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n12276) );
  OAI211_X1 U14136 ( .C1(n13325), .C2(n14556), .A(n12277), .B(n12276), .ZN(
        n12278) );
  INV_X1 U14137 ( .A(n12278), .ZN(n12279) );
  NAND2_X1 U14138 ( .A1(n12280), .A2(n12279), .ZN(n14178) );
  NOR2_X1 U14139 ( .A1(n14485), .A2(n14355), .ZN(n12281) );
  NAND2_X1 U14140 ( .A1(n14485), .A2(n14355), .ZN(n12282) );
  NAND2_X1 U14141 ( .A1(n9883), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n12284) );
  INV_X1 U14142 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n12286) );
  NAND2_X1 U14143 ( .A1(n12287), .A2(n12286), .ZN(n12288) );
  NAND2_X1 U14144 ( .A1(n12298), .A2(n12288), .ZN(n14056) );
  OR2_X1 U14145 ( .A1(n14056), .A2(n12314), .ZN(n12294) );
  INV_X1 U14146 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n12291) );
  NAND2_X1 U14147 ( .A1(n13322), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n12290) );
  NAND2_X1 U14148 ( .A1(n13321), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n12289) );
  OAI211_X1 U14149 ( .C1(n12291), .C2(n13325), .A(n12290), .B(n12289), .ZN(
        n12292) );
  INV_X1 U14150 ( .A(n12292), .ZN(n12293) );
  NAND2_X1 U14151 ( .A1(n12294), .A2(n12293), .ZN(n14177) );
  INV_X1 U14152 ( .A(n14177), .ZN(n14118) );
  XNOR2_X1 U14153 ( .A(n14480), .B(n14118), .ZN(n13396) );
  NAND2_X1 U14154 ( .A1(n14319), .A2(n14324), .ZN(n12296) );
  NAND2_X1 U14155 ( .A1(n14480), .A2(n14118), .ZN(n12295) );
  NAND2_X1 U14156 ( .A1(n13330), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n12297) );
  NAND2_X1 U14157 ( .A1(n12298), .A2(n14119), .ZN(n12299) );
  AND2_X1 U14158 ( .A1(n12300), .A2(n12299), .ZN(n14313) );
  NAND2_X1 U14159 ( .A1(n14313), .A2(n12342), .ZN(n12306) );
  INV_X1 U14160 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n12303) );
  NAND2_X1 U14161 ( .A1(n13322), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n12302) );
  NAND2_X1 U14162 ( .A1(n13321), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n12301) );
  OAI211_X1 U14163 ( .C1(n12303), .C2(n13325), .A(n12302), .B(n12301), .ZN(
        n12304) );
  INV_X1 U14164 ( .A(n12304), .ZN(n12305) );
  NAND2_X1 U14165 ( .A1(n12306), .A2(n12305), .ZN(n14176) );
  INV_X1 U14166 ( .A(n14176), .ZN(n14104) );
  NAND2_X1 U14167 ( .A1(n14475), .A2(n14104), .ZN(n12307) );
  NAND2_X1 U14168 ( .A1(n14470), .A2(n14158), .ZN(n12308) );
  NAND2_X1 U14169 ( .A1(n14277), .A2(n13311), .ZN(n12309) );
  NAND2_X1 U14170 ( .A1(n13330), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12310) );
  INV_X1 U14171 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n14050) );
  NAND2_X1 U14172 ( .A1(n12312), .A2(n14050), .ZN(n12313) );
  NAND2_X1 U14173 ( .A1(n12324), .A2(n12313), .ZN(n14267) );
  OR2_X1 U14174 ( .A1(n14267), .A2(n12314), .ZN(n12320) );
  INV_X1 U14175 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n12317) );
  NAND2_X1 U14176 ( .A1(n13321), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n12316) );
  NAND2_X1 U14177 ( .A1(n12345), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n12315) );
  OAI211_X1 U14178 ( .C1(n12317), .C2(n13325), .A(n12316), .B(n12315), .ZN(
        n12318) );
  INV_X1 U14179 ( .A(n12318), .ZN(n12319) );
  XNOR2_X1 U14180 ( .A(n14463), .B(n14173), .ZN(n14262) );
  INV_X1 U14181 ( .A(n14173), .ZN(n14159) );
  NAND2_X1 U14182 ( .A1(n14463), .A2(n14159), .ZN(n12321) );
  NAND2_X1 U14183 ( .A1(n9883), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12322) );
  INV_X1 U14184 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n14081) );
  NAND2_X1 U14185 ( .A1(n12324), .A2(n14081), .ZN(n12325) );
  NAND2_X1 U14186 ( .A1(n12335), .A2(n12325), .ZN(n14082) );
  INV_X1 U14187 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n14543) );
  NAND2_X1 U14188 ( .A1(n13321), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n12327) );
  NAND2_X1 U14189 ( .A1(n13322), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n12326) );
  OAI211_X1 U14190 ( .C1(n14543), .C2(n13325), .A(n12327), .B(n12326), .ZN(
        n12328) );
  NAND2_X1 U14191 ( .A1(n14076), .A2(n14047), .ZN(n12329) );
  NAND2_X1 U14192 ( .A1(n9883), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12333) );
  INV_X1 U14193 ( .A(n12335), .ZN(n12352) );
  INV_X1 U14194 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n12340) );
  NAND2_X1 U14195 ( .A1(n13321), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n12338) );
  NAND2_X1 U14196 ( .A1(n12336), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n12337) );
  OAI211_X1 U14197 ( .C1(n12340), .C2(n12339), .A(n12338), .B(n12337), .ZN(
        n12341) );
  AOI21_X1 U14198 ( .B1(n12352), .B2(n12342), .A(n12341), .ZN(n14078) );
  XNOR2_X1 U14199 ( .A(n14453), .B(n14078), .ZN(n13403) );
  INV_X1 U14200 ( .A(n14047), .ZN(n14172) );
  NOR2_X1 U14201 ( .A1(n13408), .A2(n13410), .ZN(n12344) );
  NOR2_X1 U14202 ( .A1(n14356), .A2(n12344), .ZN(n14235) );
  INV_X1 U14203 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n14538) );
  NAND2_X1 U14204 ( .A1(n13321), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n12347) );
  NAND2_X1 U14205 ( .A1(n12345), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n12346) );
  OAI211_X1 U14206 ( .C1(n13325), .C2(n14538), .A(n12347), .B(n12346), .ZN(
        n14170) );
  NAND2_X1 U14207 ( .A1(n14400), .A2(n14567), .ZN(n14375) );
  OR2_X2 U14208 ( .A1(n14344), .A2(n14480), .ZN(n14326) );
  AND2_X2 U14209 ( .A1(n14544), .A2(n14264), .ZN(n14253) );
  INV_X1 U14210 ( .A(n14253), .ZN(n12351) );
  AND2_X2 U14211 ( .A1(n13329), .A2(n14253), .ZN(n14240) );
  AOI211_X1 U14212 ( .C1(n14453), .C2(n12351), .A(n14416), .B(n14240), .ZN(
        n14452) );
  AOI22_X1 U14213 ( .A1(n12352), .A2(n14376), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14378), .ZN(n12353) );
  OAI21_X1 U14214 ( .B1(n13329), .B2(n14366), .A(n12353), .ZN(n12367) );
  OR2_X1 U14215 ( .A1(n14511), .A2(n14182), .ZN(n12355) );
  NAND2_X1 U14216 ( .A1(n14406), .A2(n12355), .ZN(n14383) );
  OR2_X1 U14217 ( .A1(n14570), .A2(n14181), .ZN(n12356) );
  XNOR2_X1 U14218 ( .A(n14502), .B(n14353), .ZN(n14373) );
  OR2_X1 U14219 ( .A1(n14361), .A2(n14179), .ZN(n12357) );
  XNOR2_X1 U14220 ( .A(n14485), .B(n14355), .ZN(n13395) );
  NAND2_X1 U14221 ( .A1(n14485), .A2(n14178), .ZN(n12359) );
  OR2_X1 U14222 ( .A1(n14480), .A2(n14177), .ZN(n12360) );
  NAND2_X1 U14223 ( .A1(n14475), .A2(n14176), .ZN(n12361) );
  OAI22_X1 U14224 ( .A1(n14273), .A2(n12363), .B1(n13311), .B2(n14551), .ZN(
        n14263) );
  AND2_X1 U14225 ( .A1(n14463), .A2(n14173), .ZN(n12364) );
  AOI21_X1 U14226 ( .B1(n14263), .B2(n7793), .A(n12364), .ZN(n14251) );
  INV_X1 U14227 ( .A(n14250), .ZN(n12365) );
  OAI22_X1 U14228 ( .A1(n14251), .A2(n12365), .B1(n14047), .B2(n14544), .ZN(
        n12366) );
  INV_X1 U14229 ( .A(n12368), .ZN(n15155) );
  OAI222_X1 U14230 ( .A1(n14588), .A2(n12369), .B1(n14593), .B2(n15155), .C1(
        P2_U3088), .C2(n13408), .ZN(P2_U3300) );
  XNOR2_X1 U14231 ( .A(n14361), .B(n14043), .ZN(n12390) );
  NAND2_X1 U14232 ( .A1(n14179), .A2(n14416), .ZN(n12391) );
  NAND2_X1 U14233 ( .A1(n14183), .A2(n14416), .ZN(n12373) );
  INV_X1 U14234 ( .A(n12373), .ZN(n12376) );
  XNOR2_X1 U14235 ( .A(n14577), .B(n14043), .ZN(n12375) );
  INV_X1 U14236 ( .A(n12370), .ZN(n12415) );
  INV_X1 U14237 ( .A(n12371), .ZN(n12372) );
  NOR2_X1 U14238 ( .A1(n12415), .A2(n12372), .ZN(n12374) );
  XNOR2_X1 U14239 ( .A(n12375), .B(n12373), .ZN(n12416) );
  XNOR2_X1 U14240 ( .A(n14511), .B(n14043), .ZN(n14064) );
  AND2_X1 U14241 ( .A1(n14182), .A2(n14416), .ZN(n12377) );
  NAND2_X1 U14242 ( .A1(n14064), .A2(n12377), .ZN(n12378) );
  OAI21_X1 U14243 ( .B1(n14064), .B2(n12377), .A(n12378), .ZN(n14146) );
  INV_X1 U14244 ( .A(n12378), .ZN(n12383) );
  XNOR2_X1 U14245 ( .A(n14570), .B(n14043), .ZN(n12379) );
  AND2_X1 U14246 ( .A1(n14181), .A2(n14416), .ZN(n12380) );
  NAND2_X1 U14247 ( .A1(n12379), .A2(n12380), .ZN(n12388) );
  INV_X1 U14248 ( .A(n12379), .ZN(n14125) );
  INV_X1 U14249 ( .A(n12380), .ZN(n12381) );
  NAND2_X1 U14250 ( .A1(n14125), .A2(n12381), .ZN(n12382) );
  AND2_X1 U14251 ( .A1(n12388), .A2(n12382), .ZN(n14062) );
  XNOR2_X1 U14252 ( .A(n14502), .B(n14043), .ZN(n12384) );
  AND2_X1 U14253 ( .A1(n14180), .A2(n14416), .ZN(n12385) );
  NAND2_X1 U14254 ( .A1(n12384), .A2(n12385), .ZN(n12389) );
  INV_X1 U14255 ( .A(n12384), .ZN(n14091) );
  INV_X1 U14256 ( .A(n12385), .ZN(n12386) );
  NAND2_X1 U14257 ( .A1(n14091), .A2(n12386), .ZN(n12387) );
  NAND2_X1 U14258 ( .A1(n12389), .A2(n12387), .ZN(n14126) );
  XNOR2_X1 U14259 ( .A(n14485), .B(n14043), .ZN(n14026) );
  INV_X1 U14260 ( .A(n12392), .ZN(n12393) );
  AOI22_X1 U14261 ( .A1(n12393), .A2(n14115), .B1(n14063), .B2(n14178), .ZN(
        n12398) );
  AOI22_X1 U14262 ( .A1(n14177), .A2(n14139), .B1(n14137), .B2(n14179), .ZN(
        n14342) );
  NOR2_X1 U14263 ( .A1(n14342), .A2(n14144), .ZN(n12396) );
  OAI22_X1 U14264 ( .A1(n14337), .A2(n14161), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12394), .ZN(n12395) );
  AOI211_X1 U14265 ( .C1(n14485), .C2(n14150), .A(n12396), .B(n12395), .ZN(
        n12397) );
  OAI21_X1 U14266 ( .B1(n14029), .B2(n12398), .A(n12397), .ZN(P2_U3207) );
  NAND3_X1 U14267 ( .A1(n12399), .A2(n14063), .A3(n14193), .ZN(n12400) );
  OAI21_X1 U14268 ( .B1(n12401), .B2(n14168), .A(n12400), .ZN(n12408) );
  INV_X1 U14269 ( .A(n12402), .ZN(n12407) );
  AOI22_X1 U14270 ( .A1(n14141), .A2(n14429), .B1(P2_REG3_REG_9__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12405) );
  NAND2_X1 U14271 ( .A1(n14165), .A2(n12403), .ZN(n12404) );
  OAI211_X1 U14272 ( .C1(n7372), .C2(n14162), .A(n12405), .B(n12404), .ZN(
        n12406) );
  AOI21_X1 U14273 ( .B1(n12408), .B2(n12407), .A(n12406), .ZN(n12409) );
  OAI21_X1 U14274 ( .B1(n14168), .B2(n12410), .A(n12409), .ZN(P2_U3203) );
  NAND2_X1 U14275 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3088), .ZN(n15459)
         );
  OAI21_X1 U14276 ( .B1(n14161), .B2(n12411), .A(n15459), .ZN(n12412) );
  AOI21_X1 U14277 ( .B1(n14099), .B2(n14182), .A(n12412), .ZN(n12413) );
  OAI21_X1 U14278 ( .B1(n12414), .B2(n14096), .A(n12413), .ZN(n12420) );
  AOI22_X1 U14279 ( .A1(n12415), .A2(n14115), .B1(n14063), .B2(n14184), .ZN(
        n12417) );
  NOR3_X1 U14280 ( .A1(n12418), .A2(n12417), .A3(n12416), .ZN(n12419) );
  AOI211_X1 U14281 ( .C1(n14577), .C2(n14150), .A(n12420), .B(n12419), .ZN(
        n12421) );
  OAI21_X1 U14282 ( .B1(n14168), .B2(n12422), .A(n12421), .ZN(P2_U3200) );
  AOI22_X1 U14283 ( .A1(n14656), .A2(n12519), .B1(n12518), .B2(n14737), .ZN(
        n12442) );
  AOI22_X1 U14284 ( .A1(n14656), .A2(n7181), .B1(n12519), .B2(n14737), .ZN(
        n12423) );
  XNOR2_X1 U14285 ( .A(n12423), .B(n12526), .ZN(n12443) );
  NAND2_X1 U14286 ( .A1(n16128), .A2(n7181), .ZN(n12425) );
  NAND2_X1 U14287 ( .A1(n14739), .A2(n12519), .ZN(n12424) );
  NAND2_X1 U14288 ( .A1(n12425), .A2(n12424), .ZN(n12426) );
  XNOR2_X1 U14289 ( .A(n12426), .B(n12526), .ZN(n12435) );
  AND2_X1 U14290 ( .A1(n12518), .A2(n14739), .ZN(n12427) );
  AOI21_X1 U14291 ( .B1(n16128), .B2(n12519), .A(n12427), .ZN(n12433) );
  XNOR2_X1 U14292 ( .A(n12435), .B(n12433), .ZN(n16119) );
  INV_X1 U14293 ( .A(n12428), .ZN(n12431) );
  INV_X1 U14294 ( .A(n12429), .ZN(n12430) );
  NAND2_X1 U14295 ( .A1(n12431), .A2(n12430), .ZN(n16120) );
  INV_X1 U14296 ( .A(n12433), .ZN(n12434) );
  NAND2_X1 U14297 ( .A1(n15122), .A2(n12514), .ZN(n12437) );
  NAND2_X1 U14298 ( .A1(n14738), .A2(n12519), .ZN(n12436) );
  NAND2_X1 U14299 ( .A1(n12437), .A2(n12436), .ZN(n12438) );
  XNOR2_X1 U14300 ( .A(n12438), .B(n12526), .ZN(n12439) );
  OAI22_X1 U14301 ( .A1(n14732), .A2(n12525), .B1(n16116), .B2(n12524), .ZN(
        n14721) );
  NAND2_X1 U14302 ( .A1(n14722), .A2(n14721), .ZN(n14720) );
  INV_X1 U14303 ( .A(n12439), .ZN(n12440) );
  NAND2_X1 U14304 ( .A1(n14720), .A2(n8176), .ZN(n14650) );
  INV_X1 U14305 ( .A(n14650), .ZN(n12445) );
  XNOR2_X1 U14306 ( .A(n12443), .B(n12442), .ZN(n14651) );
  NAND2_X1 U14307 ( .A1(n14669), .A2(n7181), .ZN(n12447) );
  NAND2_X1 U14308 ( .A1(n14736), .A2(n12519), .ZN(n12446) );
  NAND2_X1 U14309 ( .A1(n12447), .A2(n12446), .ZN(n12448) );
  XNOR2_X1 U14310 ( .A(n12448), .B(n12526), .ZN(n14660) );
  NAND2_X1 U14311 ( .A1(n14669), .A2(n12519), .ZN(n12450) );
  NAND2_X1 U14312 ( .A1(n14736), .A2(n12518), .ZN(n12449) );
  NAND2_X1 U14313 ( .A1(n12450), .A2(n12449), .ZN(n14659) );
  NOR2_X1 U14314 ( .A1(n14660), .A2(n14659), .ZN(n12451) );
  NAND2_X1 U14315 ( .A1(n15104), .A2(n7181), .ZN(n12453) );
  NAND2_X1 U14316 ( .A1(n14735), .A2(n12519), .ZN(n12452) );
  NAND2_X1 U14317 ( .A1(n12453), .A2(n12452), .ZN(n12454) );
  XNOR2_X1 U14318 ( .A(n12454), .B(n8186), .ZN(n12457) );
  AND2_X1 U14319 ( .A1(n14735), .A2(n12518), .ZN(n12455) );
  AOI21_X1 U14320 ( .B1(n15104), .B2(n12519), .A(n12455), .ZN(n12456) );
  NAND2_X1 U14321 ( .A1(n12457), .A2(n12456), .ZN(n12459) );
  OAI21_X1 U14322 ( .B1(n12457), .B2(n12456), .A(n12459), .ZN(n14703) );
  INV_X1 U14323 ( .A(n14703), .ZN(n12458) );
  NAND2_X2 U14324 ( .A1(n14700), .A2(n12459), .ZN(n14621) );
  OR2_X1 U14325 ( .A1(n15097), .A2(n12525), .ZN(n12461) );
  NAND2_X1 U14326 ( .A1(n14979), .A2(n12518), .ZN(n12460) );
  NAND2_X1 U14327 ( .A1(n12461), .A2(n12460), .ZN(n12465) );
  OAI22_X1 U14328 ( .A1(n15097), .A2(n12523), .B1(n15006), .B2(n12525), .ZN(
        n12462) );
  XNOR2_X1 U14329 ( .A(n12462), .B(n12526), .ZN(n12464) );
  XOR2_X1 U14330 ( .A(n12465), .B(n12464), .Z(n14622) );
  OAI22_X1 U14331 ( .A1(n14976), .A2(n12525), .B1(n14637), .B2(n12524), .ZN(
        n12473) );
  OAI22_X1 U14332 ( .A1(n14976), .A2(n12523), .B1(n14637), .B2(n12525), .ZN(
        n12463) );
  XNOR2_X1 U14333 ( .A(n12463), .B(n12526), .ZN(n12474) );
  XOR2_X1 U14334 ( .A(n12473), .B(n12474), .Z(n14682) );
  INV_X1 U14335 ( .A(n12464), .ZN(n12467) );
  INV_X1 U14336 ( .A(n12465), .ZN(n12466) );
  NAND2_X1 U14337 ( .A1(n12467), .A2(n12466), .ZN(n14679) );
  NAND2_X1 U14338 ( .A1(n15082), .A2(n7181), .ZN(n12470) );
  NAND2_X1 U14339 ( .A1(n14981), .A2(n12519), .ZN(n12469) );
  NAND2_X1 U14340 ( .A1(n12470), .A2(n12469), .ZN(n12471) );
  XNOR2_X1 U14341 ( .A(n12471), .B(n12526), .ZN(n12476) );
  AND2_X1 U14342 ( .A1(n14981), .A2(n12518), .ZN(n12472) );
  AOI21_X1 U14343 ( .B1(n15082), .B2(n12519), .A(n12472), .ZN(n12477) );
  XNOR2_X1 U14344 ( .A(n12476), .B(n12477), .ZN(n14631) );
  NAND2_X1 U14345 ( .A1(n12474), .A2(n12473), .ZN(n14632) );
  INV_X1 U14346 ( .A(n12476), .ZN(n12478) );
  OAI22_X1 U14347 ( .A1(n15075), .A2(n12523), .B1(n12911), .B2(n12525), .ZN(
        n12479) );
  XNOR2_X1 U14348 ( .A(n12479), .B(n12526), .ZN(n12482) );
  OR2_X1 U14349 ( .A1(n15075), .A2(n12525), .ZN(n12481) );
  NAND2_X1 U14350 ( .A1(n14961), .A2(n12518), .ZN(n12480) );
  NAND2_X1 U14351 ( .A1(n12481), .A2(n12480), .ZN(n12483) );
  NAND2_X1 U14352 ( .A1(n12482), .A2(n12483), .ZN(n14693) );
  INV_X1 U14353 ( .A(n12482), .ZN(n12485) );
  INV_X1 U14354 ( .A(n12483), .ZN(n12484) );
  NAND2_X1 U14355 ( .A1(n12485), .A2(n12484), .ZN(n14692) );
  NAND2_X1 U14356 ( .A1(n15069), .A2(n12514), .ZN(n12487) );
  NAND2_X1 U14357 ( .A1(n14951), .A2(n12519), .ZN(n12486) );
  NAND2_X1 U14358 ( .A1(n12487), .A2(n12486), .ZN(n12488) );
  XNOR2_X1 U14359 ( .A(n12488), .B(n12526), .ZN(n12489) );
  AOI22_X1 U14360 ( .A1(n15069), .A2(n12519), .B1(n12518), .B2(n14951), .ZN(
        n12490) );
  XNOR2_X1 U14361 ( .A(n12489), .B(n12490), .ZN(n14614) );
  INV_X1 U14362 ( .A(n12489), .ZN(n12491) );
  NAND2_X1 U14363 ( .A1(n12491), .A2(n12490), .ZN(n12492) );
  NAND2_X1 U14364 ( .A1(n15064), .A2(n12514), .ZN(n12494) );
  NAND2_X1 U14365 ( .A1(n14900), .A2(n12519), .ZN(n12493) );
  NAND2_X1 U14366 ( .A1(n12494), .A2(n12493), .ZN(n12495) );
  XNOR2_X1 U14367 ( .A(n12495), .B(n12526), .ZN(n12496) );
  AOI22_X1 U14368 ( .A1(n15064), .A2(n12519), .B1(n12518), .B2(n14900), .ZN(
        n12497) );
  XNOR2_X1 U14369 ( .A(n12496), .B(n12497), .ZN(n14673) );
  INV_X1 U14370 ( .A(n12496), .ZN(n12498) );
  NAND2_X1 U14371 ( .A1(n15057), .A2(n12514), .ZN(n12500) );
  NAND2_X1 U14372 ( .A1(n14881), .A2(n12519), .ZN(n12499) );
  NAND2_X1 U14373 ( .A1(n12500), .A2(n12499), .ZN(n12501) );
  XNOR2_X1 U14374 ( .A(n12501), .B(n12526), .ZN(n12502) );
  AOI22_X1 U14375 ( .A1(n15057), .A2(n12519), .B1(n12518), .B2(n14881), .ZN(
        n12503) );
  XNOR2_X1 U14376 ( .A(n12502), .B(n12503), .ZN(n14642) );
  NAND2_X1 U14377 ( .A1(n14641), .A2(n14642), .ZN(n12506) );
  INV_X1 U14378 ( .A(n12502), .ZN(n12504) );
  NAND2_X1 U14379 ( .A1(n12504), .A2(n12503), .ZN(n12505) );
  NAND2_X1 U14380 ( .A1(n12506), .A2(n12505), .ZN(n14710) );
  NAND2_X1 U14381 ( .A1(n15051), .A2(n7181), .ZN(n12508) );
  NAND2_X1 U14382 ( .A1(n14899), .A2(n12519), .ZN(n12507) );
  NAND2_X1 U14383 ( .A1(n12508), .A2(n12507), .ZN(n12509) );
  XNOR2_X1 U14384 ( .A(n12509), .B(n12526), .ZN(n12510) );
  AOI22_X1 U14385 ( .A1(n15051), .A2(n12519), .B1(n12518), .B2(n14899), .ZN(
        n12511) );
  XNOR2_X1 U14386 ( .A(n12510), .B(n12511), .ZN(n14711) );
  INV_X1 U14387 ( .A(n12510), .ZN(n12512) );
  NAND2_X1 U14388 ( .A1(n12512), .A2(n12511), .ZN(n12513) );
  NAND2_X1 U14389 ( .A1(n14871), .A2(n7181), .ZN(n12516) );
  NAND2_X1 U14390 ( .A1(n14882), .A2(n12519), .ZN(n12515) );
  NAND2_X1 U14391 ( .A1(n12516), .A2(n12515), .ZN(n12517) );
  XNOR2_X1 U14392 ( .A(n12517), .B(n12526), .ZN(n12520) );
  AOI22_X1 U14393 ( .A1(n14871), .A2(n12519), .B1(n12518), .B2(n14882), .ZN(
        n12521) );
  XNOR2_X1 U14394 ( .A(n12520), .B(n12521), .ZN(n14606) );
  INV_X1 U14395 ( .A(n12520), .ZN(n12522) );
  INV_X1 U14396 ( .A(n14857), .ZN(n14609) );
  OAI22_X1 U14397 ( .A1(n12555), .A2(n12523), .B1(n14609), .B2(n12525), .ZN(
        n12529) );
  OAI22_X1 U14398 ( .A1(n12555), .A2(n12525), .B1(n14609), .B2(n12524), .ZN(
        n12527) );
  XNOR2_X1 U14399 ( .A(n12527), .B(n12526), .ZN(n12528) );
  XOR2_X1 U14400 ( .A(n12529), .B(n12528), .Z(n12530) );
  INV_X1 U14401 ( .A(n14734), .ZN(n12539) );
  AOI22_X1 U14402 ( .A1(n12531), .A2(n14728), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12533) );
  NAND2_X1 U14403 ( .A1(n14882), .A2(n14713), .ZN(n12532) );
  OAI211_X1 U14404 ( .C1(n12539), .C2(n16115), .A(n12533), .B(n12532), .ZN(
        n12534) );
  AOI21_X1 U14405 ( .B1(n15040), .B2(n16129), .A(n12534), .ZN(n12535) );
  OAI21_X1 U14406 ( .B1(n12536), .B2(n16123), .A(n12535), .ZN(P1_U3220) );
  NAND2_X1 U14407 ( .A1(n14586), .A2(n12089), .ZN(n12538) );
  NAND2_X1 U14408 ( .A1(n10053), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12537) );
  XNOR2_X1 U14409 ( .A(n15031), .B(n12539), .ZN(n13058) );
  AOI21_X1 U14410 ( .B1(n15031), .B2(n12543), .A(n14850), .ZN(n15035) );
  NAND2_X1 U14411 ( .A1(n15031), .A2(n15990), .ZN(n12552) );
  INV_X1 U14412 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n12546) );
  NAND2_X1 U14413 ( .A1(n12987), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n12545) );
  NAND2_X1 U14414 ( .A1(n12988), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n12544) );
  OAI211_X1 U14415 ( .C1(n12992), .C2(n12546), .A(n12545), .B(n12544), .ZN(
        n14733) );
  INV_X1 U14416 ( .A(P1_B_REG_SCAN_IN), .ZN(n12547) );
  NOR2_X1 U14417 ( .A1(n15154), .A2(n12547), .ZN(n12548) );
  NOR2_X1 U14418 ( .A1(n15005), .A2(n12548), .ZN(n14844) );
  NAND2_X1 U14419 ( .A1(n14733), .A2(n14844), .ZN(n15032) );
  INV_X1 U14420 ( .A(n15032), .ZN(n12549) );
  AOI22_X1 U14421 ( .A1(n16047), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n12550), 
        .B2(n12549), .ZN(n12551) );
  OAI211_X1 U14422 ( .C1(n15016), .C2(n12553), .A(n12552), .B(n12551), .ZN(
        n12554) );
  AOI21_X1 U14423 ( .B1(n15035), .B2(n14843), .A(n12554), .ZN(n12561) );
  NAND2_X1 U14424 ( .A1(n12555), .A2(n14857), .ZN(n12556) );
  NAND2_X1 U14425 ( .A1(n14857), .A2(n14978), .ZN(n15033) );
  AOI21_X1 U14426 ( .B1(n15038), .B2(n15033), .A(n15998), .ZN(n12559) );
  INV_X1 U14427 ( .A(n12559), .ZN(n12560) );
  OAI211_X1 U14428 ( .C1(n15037), .C2(n14967), .A(n12561), .B(n12560), .ZN(
        P1_U3356) );
  INV_X1 U14429 ( .A(n12562), .ZN(n12563) );
  INV_X1 U14430 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12796) );
  XNOR2_X1 U14431 ( .A(n12796), .B(P1_DATAO_REG_30__SCAN_IN), .ZN(n12582) );
  INV_X1 U14432 ( .A(n12582), .ZN(n12565) );
  NAND2_X1 U14433 ( .A1(n12583), .A2(n12565), .ZN(n12567) );
  NAND2_X1 U14434 ( .A1(n12796), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12566) );
  NAND2_X1 U14435 ( .A1(n12567), .A2(n12566), .ZN(n12570) );
  INV_X1 U14436 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n12568) );
  XNOR2_X1 U14437 ( .A(n12568), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n12569) );
  XNOR2_X1 U14438 ( .A(n12570), .B(n12569), .ZN(n14023) );
  NAND2_X1 U14439 ( .A1(n14023), .A2(n12584), .ZN(n12572) );
  INV_X1 U14440 ( .A(SI_31_), .ZN(n14019) );
  OR2_X1 U14441 ( .A1(n8390), .A2(n14019), .ZN(n12571) );
  NAND2_X1 U14442 ( .A1(n12572), .A2(n12571), .ZN(n12588) );
  INV_X1 U14443 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12578) );
  NAND2_X1 U14444 ( .A1(n12573), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12576) );
  INV_X1 U14445 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12574) );
  OR2_X1 U14446 ( .A1(n8889), .A2(n12574), .ZN(n12575) );
  OAI211_X1 U14447 ( .C1(n12578), .C2(n12577), .A(n12576), .B(n12575), .ZN(
        n12579) );
  INV_X1 U14448 ( .A(n12579), .ZN(n12580) );
  XNOR2_X1 U14449 ( .A(n12583), .B(n12582), .ZN(n13080) );
  NAND2_X1 U14450 ( .A1(n13080), .A2(n12584), .ZN(n12586) );
  OR2_X1 U14451 ( .A1(n8390), .A2(n15290), .ZN(n12585) );
  INV_X1 U14452 ( .A(n16162), .ZN(n13675) );
  AOI22_X1 U14453 ( .A1(n12587), .A2(n12774), .B1(n13555), .B2(n16162), .ZN(
        n12593) );
  OR2_X1 U14454 ( .A1(n12588), .A2(n13555), .ZN(n12780) );
  INV_X1 U14455 ( .A(n13556), .ZN(n12589) );
  NAND2_X1 U14456 ( .A1(n16162), .A2(n12589), .ZN(n12590) );
  NAND2_X1 U14457 ( .A1(n12780), .A2(n12590), .ZN(n12619) );
  INV_X1 U14458 ( .A(n12591), .ZN(n12592) );
  NOR2_X1 U14459 ( .A1(n12619), .A2(n12592), .ZN(n12779) );
  NAND2_X1 U14460 ( .A1(n12593), .A2(n12779), .ZN(n12594) );
  OAI21_X1 U14461 ( .B1(n13962), .B2(n12782), .A(n12594), .ZN(n12597) );
  NOR2_X1 U14462 ( .A1(n12596), .A2(n13656), .ZN(n12621) );
  NAND2_X1 U14463 ( .A1(n12621), .A2(n12641), .ZN(n12595) );
  NOR2_X1 U14464 ( .A1(n12596), .A2(n13670), .ZN(n12624) );
  INV_X1 U14465 ( .A(n13710), .ZN(n13707) );
  NOR2_X1 U14466 ( .A1(n13701), .A2(n13707), .ZN(n12598) );
  NAND2_X1 U14467 ( .A1(n12599), .A2(n12598), .ZN(n12771) );
  NAND4_X1 U14468 ( .A1(n12659), .A2(n12675), .A3(n12600), .A4(n12668), .ZN(
        n12601) );
  OR2_X1 U14469 ( .A1(n12601), .A2(n8117), .ZN(n12608) );
  NOR2_X1 U14470 ( .A1(n12603), .A2(n12602), .ZN(n12606) );
  NOR2_X1 U14471 ( .A1(n7361), .A2(n15870), .ZN(n12605) );
  NAND4_X1 U14472 ( .A1(n12606), .A2(n12605), .A3(n12691), .A4(n8177), .ZN(
        n12607) );
  NOR2_X1 U14473 ( .A1(n12608), .A2(n12607), .ZN(n12610) );
  NAND4_X1 U14474 ( .A1(n12610), .A2(n12696), .A3(n12609), .A4(n12703), .ZN(
        n12611) );
  OR4_X1 U14475 ( .A1(n13840), .A2(n13837), .A3(n13872), .A4(n12611), .ZN(
        n12612) );
  NOR2_X1 U14476 ( .A1(n13820), .A2(n12612), .ZN(n12613) );
  NAND4_X1 U14477 ( .A1(n13769), .A2(n13796), .A3(n13812), .A4(n12613), .ZN(
        n12614) );
  OR3_X1 U14478 ( .A1(n12752), .A2(n12615), .A3(n12614), .ZN(n12616) );
  OR3_X1 U14479 ( .A1(n13722), .A2(n13740), .A3(n12616), .ZN(n12617) );
  OR3_X1 U14480 ( .A1(n12771), .A2(n13685), .A3(n12617), .ZN(n12620) );
  NAND3_X1 U14481 ( .A1(n12622), .A2(n12621), .A3(n12623), .ZN(n12628) );
  NAND3_X1 U14482 ( .A1(n12625), .A2(n12624), .A3(n12623), .ZN(n12627) );
  INV_X1 U14483 ( .A(n12791), .ZN(n12626) );
  NAND3_X1 U14484 ( .A1(n12630), .A2(n12629), .A3(n8175), .ZN(n12795) );
  INV_X1 U14485 ( .A(n12631), .ZN(n12640) );
  NAND2_X1 U14486 ( .A1(n12632), .A2(n13486), .ZN(n12633) );
  NAND2_X1 U14487 ( .A1(n12634), .A2(n12633), .ZN(n12636) );
  NAND2_X1 U14488 ( .A1(n12636), .A2(n12635), .ZN(n12637) );
  NAND2_X1 U14489 ( .A1(n13682), .A2(n12637), .ZN(n12639) );
  NAND2_X1 U14490 ( .A1(n12639), .A2(n12638), .ZN(n12769) );
  OAI21_X1 U14491 ( .B1(n12771), .B2(n12640), .A(n12769), .ZN(n12768) );
  AND3_X1 U14492 ( .A1(n12644), .A2(n12643), .A3(n12641), .ZN(n12642) );
  NOR2_X1 U14493 ( .A1(n15871), .A2(n12642), .ZN(n12648) );
  NAND2_X1 U14494 ( .A1(n12644), .A2(n12643), .ZN(n12645) );
  NAND2_X1 U14495 ( .A1(n12646), .A2(n12645), .ZN(n12647) );
  MUX2_X1 U14496 ( .A(n12648), .B(n12647), .S(n12772), .Z(n12655) );
  NAND2_X1 U14497 ( .A1(n12657), .A2(n12649), .ZN(n12652) );
  NAND2_X1 U14498 ( .A1(n12656), .A2(n12650), .ZN(n12651) );
  MUX2_X1 U14499 ( .A(n12652), .B(n12651), .S(n12762), .Z(n12653) );
  INV_X1 U14500 ( .A(n12653), .ZN(n12654) );
  OAI21_X1 U14501 ( .B1(n12655), .B2(n15870), .A(n12654), .ZN(n12660) );
  MUX2_X1 U14502 ( .A(n12657), .B(n12656), .S(n12772), .Z(n12658) );
  NAND3_X1 U14503 ( .A1(n12660), .A2(n12659), .A3(n12658), .ZN(n12664) );
  MUX2_X1 U14504 ( .A(n12662), .B(n12661), .S(n12762), .Z(n12663) );
  AOI21_X1 U14505 ( .B1(n12664), .B2(n12663), .A(n8117), .ZN(n12674) );
  NAND2_X1 U14506 ( .A1(n13574), .A2(n12665), .ZN(n12667) );
  MUX2_X1 U14507 ( .A(n12667), .B(n12666), .S(n12762), .Z(n12669) );
  NAND2_X1 U14508 ( .A1(n12669), .A2(n12668), .ZN(n12673) );
  MUX2_X1 U14509 ( .A(n12671), .B(n12670), .S(n12772), .Z(n12672) );
  OAI21_X1 U14510 ( .B1(n12674), .B2(n12673), .A(n12672), .ZN(n12676) );
  NAND2_X1 U14511 ( .A1(n12676), .A2(n12675), .ZN(n12681) );
  MUX2_X1 U14512 ( .A(n12678), .B(n12677), .S(n12772), .Z(n12679) );
  NAND3_X1 U14513 ( .A1(n12681), .A2(n12680), .A3(n12679), .ZN(n12684) );
  NAND3_X1 U14514 ( .A1(n12687), .A2(n12682), .A3(n12762), .ZN(n12683) );
  NAND3_X1 U14515 ( .A1(n12684), .A2(n8177), .A3(n12683), .ZN(n12690) );
  NAND2_X1 U14516 ( .A1(n12685), .A2(n12762), .ZN(n12689) );
  NAND2_X1 U14517 ( .A1(n16005), .A2(n12772), .ZN(n12686) );
  NOR2_X1 U14518 ( .A1(n12687), .A2(n12686), .ZN(n12688) );
  AOI21_X1 U14519 ( .B1(n12690), .B2(n12689), .A(n12688), .ZN(n12693) );
  NOR3_X1 U14520 ( .A1(n13570), .A2(n16026), .A3(n12762), .ZN(n12692) );
  OAI21_X1 U14521 ( .B1(n12693), .B2(n12692), .A(n12691), .ZN(n12699) );
  MUX2_X1 U14522 ( .A(n12695), .B(n12694), .S(n12772), .Z(n12697) );
  AND2_X1 U14523 ( .A1(n12697), .A2(n12696), .ZN(n12698) );
  NAND2_X1 U14524 ( .A1(n12699), .A2(n12698), .ZN(n12708) );
  AND2_X1 U14525 ( .A1(n12709), .A2(n12700), .ZN(n12702) );
  NAND2_X1 U14526 ( .A1(n12706), .A2(n12762), .ZN(n12701) );
  AOI21_X1 U14527 ( .B1(n12708), .B2(n12702), .A(n12701), .ZN(n12705) );
  OAI22_X1 U14528 ( .A1(n12705), .A2(n15388), .B1(n12772), .B2(n12704), .ZN(
        n12712) );
  INV_X1 U14529 ( .A(n13872), .ZN(n13880) );
  NAND3_X1 U14530 ( .A1(n12708), .A2(n12707), .A3(n12706), .ZN(n12710) );
  NAND3_X1 U14531 ( .A1(n12710), .A2(n12772), .A3(n12709), .ZN(n12711) );
  NAND3_X1 U14532 ( .A1(n12712), .A2(n13880), .A3(n12711), .ZN(n12717) );
  INV_X1 U14533 ( .A(n13837), .ZN(n13856) );
  OR2_X1 U14534 ( .A1(n12713), .A2(n7752), .ZN(n12715) );
  MUX2_X1 U14535 ( .A(n12715), .B(n12714), .S(n12762), .Z(n12716) );
  NAND3_X1 U14536 ( .A1(n12717), .A2(n13856), .A3(n12716), .ZN(n12721) );
  MUX2_X1 U14537 ( .A(n12719), .B(n12718), .S(n12762), .Z(n12720) );
  NAND2_X1 U14538 ( .A1(n12721), .A2(n12720), .ZN(n12727) );
  INV_X1 U14539 ( .A(n12722), .ZN(n12724) );
  MUX2_X1 U14540 ( .A(n13859), .B(n13847), .S(n12762), .Z(n12723) );
  AOI21_X1 U14541 ( .B1(n12727), .B2(n12724), .A(n12723), .ZN(n12729) );
  NAND2_X1 U14542 ( .A1(n13514), .A2(n13563), .ZN(n12725) );
  AND2_X1 U14543 ( .A1(n13795), .A2(n12725), .ZN(n12734) );
  NOR2_X1 U14544 ( .A1(n12727), .A2(n12726), .ZN(n12728) );
  OR4_X1 U14545 ( .A1(n12729), .A2(n12734), .A3(n12728), .A4(n13820), .ZN(
        n12744) );
  NAND2_X1 U14546 ( .A1(n12731), .A2(n12730), .ZN(n12732) );
  NAND2_X1 U14547 ( .A1(n12732), .A2(n12738), .ZN(n12733) );
  NAND2_X1 U14548 ( .A1(n12745), .A2(n12733), .ZN(n12741) );
  INV_X1 U14549 ( .A(n12734), .ZN(n12737) );
  INV_X1 U14550 ( .A(n12735), .ZN(n12736) );
  NAND2_X1 U14551 ( .A1(n12737), .A2(n12736), .ZN(n12739) );
  NAND3_X1 U14552 ( .A1(n13778), .A2(n12739), .A3(n12738), .ZN(n12740) );
  MUX2_X1 U14553 ( .A(n12741), .B(n12740), .S(n12772), .Z(n12742) );
  INV_X1 U14554 ( .A(n12742), .ZN(n12743) );
  NAND2_X1 U14555 ( .A1(n12744), .A2(n12743), .ZN(n12747) );
  MUX2_X1 U14556 ( .A(n12745), .B(n13778), .S(n12762), .Z(n12746) );
  NAND3_X1 U14557 ( .A1(n12747), .A2(n13781), .A3(n12746), .ZN(n12751) );
  MUX2_X1 U14558 ( .A(n12749), .B(n12748), .S(n12772), .Z(n12750) );
  NAND3_X1 U14559 ( .A1(n12751), .A2(n13769), .A3(n12750), .ZN(n12756) );
  INV_X1 U14560 ( .A(n12752), .ZN(n13751) );
  MUX2_X1 U14561 ( .A(n12754), .B(n12753), .S(n12762), .Z(n12755) );
  NAND3_X1 U14562 ( .A1(n12756), .A2(n13751), .A3(n12755), .ZN(n12761) );
  MUX2_X1 U14563 ( .A(n12758), .B(n12757), .S(n12772), .Z(n12759) );
  NAND3_X1 U14564 ( .A1(n12761), .A2(n12760), .A3(n12759), .ZN(n12766) );
  MUX2_X1 U14565 ( .A(n12764), .B(n12763), .S(n12762), .Z(n12765) );
  AND2_X1 U14566 ( .A1(n12766), .A2(n12765), .ZN(n12767) );
  NAND2_X1 U14567 ( .A1(n12768), .A2(n12770), .ZN(n12773) );
  INV_X1 U14568 ( .A(n12774), .ZN(n12775) );
  INV_X1 U14569 ( .A(n12779), .ZN(n12783) );
  INV_X1 U14570 ( .A(n12780), .ZN(n12781) );
  OAI22_X1 U14571 ( .A1(n12784), .A2(n12783), .B1(n12782), .B2(n12781), .ZN(
        n12785) );
  XNOR2_X1 U14572 ( .A(n12785), .B(n13670), .ZN(n12787) );
  NOR2_X1 U14573 ( .A1(n12787), .A2(n12786), .ZN(n12794) );
  NAND3_X1 U14574 ( .A1(n12789), .A2(n12788), .A3(n13664), .ZN(n12790) );
  OAI211_X1 U14575 ( .C1(n12792), .C2(n12791), .A(n12790), .B(P3_B_REG_SCAN_IN), .ZN(n12793) );
  OAI21_X1 U14576 ( .B1(n12795), .B2(n12794), .A(n12793), .ZN(P3_U3296) );
  OAI222_X1 U14577 ( .A1(n15167), .A2(n13318), .B1(n12797), .B2(P1_U3086), 
        .C1(n12796), .C2(n15157), .ZN(P1_U3325) );
  NAND2_X1 U14578 ( .A1(n12801), .A2(n13017), .ZN(n12998) );
  OAI21_X1 U14579 ( .B1(n14751), .B2(n13015), .A(n12802), .ZN(n12804) );
  NAND2_X1 U14580 ( .A1(n14751), .A2(n13015), .ZN(n12803) );
  NAND2_X1 U14581 ( .A1(n14751), .A2(n12805), .ZN(n12806) );
  NAND3_X1 U14582 ( .A1(n12813), .A2(n12868), .A3(n12806), .ZN(n12807) );
  NAND2_X1 U14583 ( .A1(n13025), .A2(n12808), .ZN(n12810) );
  INV_X1 U14584 ( .A(n12809), .ZN(n14754) );
  NAND2_X1 U14585 ( .A1(n14754), .A2(n15839), .ZN(n13024) );
  NAND2_X1 U14586 ( .A1(n12810), .A2(n13024), .ZN(n12811) );
  NAND3_X1 U14587 ( .A1(n12811), .A2(n12816), .A3(n12815), .ZN(n12812) );
  NAND2_X1 U14588 ( .A1(n12814), .A2(n12813), .ZN(n12817) );
  NAND4_X1 U14589 ( .A1(n12817), .A2(n12863), .A3(n12816), .A4(n12815), .ZN(
        n12818) );
  NAND2_X1 U14590 ( .A1(n12819), .A2(n12818), .ZN(n12822) );
  MUX2_X1 U14591 ( .A(n15918), .B(n14750), .S(n12863), .Z(n12823) );
  NAND2_X1 U14592 ( .A1(n12822), .A2(n12823), .ZN(n12821) );
  MUX2_X1 U14593 ( .A(n14750), .B(n15918), .S(n12863), .Z(n12820) );
  NAND2_X1 U14594 ( .A1(n12821), .A2(n12820), .ZN(n12827) );
  INV_X1 U14595 ( .A(n12822), .ZN(n12825) );
  INV_X1 U14596 ( .A(n12823), .ZN(n12824) );
  NAND2_X1 U14597 ( .A1(n12827), .A2(n12826), .ZN(n12829) );
  MUX2_X1 U14598 ( .A(n14749), .B(n15949), .S(n12863), .Z(n12830) );
  MUX2_X1 U14599 ( .A(n14749), .B(n15949), .S(n12868), .Z(n12828) );
  INV_X1 U14600 ( .A(n12830), .ZN(n12831) );
  MUX2_X1 U14601 ( .A(n14748), .B(n12832), .S(n12868), .Z(n12834) );
  MUX2_X1 U14602 ( .A(n14748), .B(n12832), .S(n12863), .Z(n12833) );
  INV_X1 U14603 ( .A(n12834), .ZN(n12835) );
  MUX2_X1 U14604 ( .A(n14747), .B(n15991), .S(n12863), .Z(n12839) );
  NAND2_X1 U14605 ( .A1(n12838), .A2(n12839), .ZN(n12837) );
  MUX2_X1 U14606 ( .A(n14747), .B(n15991), .S(n12868), .Z(n12836) );
  NAND2_X1 U14607 ( .A1(n12837), .A2(n12836), .ZN(n12843) );
  INV_X1 U14608 ( .A(n12838), .ZN(n12841) );
  INV_X1 U14609 ( .A(n12839), .ZN(n12840) );
  NAND2_X1 U14610 ( .A1(n12841), .A2(n12840), .ZN(n12842) );
  NAND2_X1 U14611 ( .A1(n12843), .A2(n12842), .ZN(n12846) );
  MUX2_X1 U14612 ( .A(n14746), .B(n12844), .S(n12868), .Z(n12847) );
  MUX2_X1 U14613 ( .A(n14746), .B(n12844), .S(n12863), .Z(n12845) );
  INV_X1 U14614 ( .A(n12847), .ZN(n12848) );
  MUX2_X1 U14615 ( .A(n14745), .B(n12849), .S(n12863), .Z(n12853) );
  MUX2_X1 U14616 ( .A(n14745), .B(n12849), .S(n12874), .Z(n12850) );
  NAND2_X1 U14617 ( .A1(n12851), .A2(n12850), .ZN(n12857) );
  INV_X1 U14618 ( .A(n12852), .ZN(n12855) );
  INV_X1 U14619 ( .A(n12853), .ZN(n12854) );
  NAND2_X1 U14620 ( .A1(n12855), .A2(n12854), .ZN(n12856) );
  NAND2_X1 U14621 ( .A1(n12857), .A2(n12856), .ZN(n12860) );
  MUX2_X1 U14622 ( .A(n14744), .B(n12858), .S(n12868), .Z(n12861) );
  MUX2_X1 U14623 ( .A(n14744), .B(n12858), .S(n12863), .Z(n12859) );
  INV_X1 U14624 ( .A(n12861), .ZN(n12862) );
  MUX2_X1 U14625 ( .A(n14743), .B(n12864), .S(n12863), .Z(n12866) );
  MUX2_X1 U14626 ( .A(n14743), .B(n12864), .S(n12874), .Z(n12865) );
  INV_X1 U14627 ( .A(n12866), .ZN(n12867) );
  MUX2_X1 U14628 ( .A(n14742), .B(n12869), .S(n12874), .Z(n12872) );
  MUX2_X1 U14629 ( .A(n14742), .B(n12869), .S(n13015), .Z(n12870) );
  INV_X1 U14630 ( .A(n12872), .ZN(n12873) );
  MUX2_X1 U14631 ( .A(n14741), .B(n12875), .S(n12884), .Z(n12879) );
  MUX2_X1 U14632 ( .A(n14741), .B(n12875), .S(n12874), .Z(n12876) );
  NAND2_X1 U14633 ( .A1(n12877), .A2(n12876), .ZN(n12883) );
  INV_X1 U14634 ( .A(n12878), .ZN(n12881) );
  INV_X1 U14635 ( .A(n12879), .ZN(n12880) );
  NAND2_X1 U14636 ( .A1(n12881), .A2(n12880), .ZN(n12882) );
  MUX2_X1 U14637 ( .A(n14740), .B(n12885), .S(n12868), .Z(n12887) );
  MUX2_X1 U14638 ( .A(n14740), .B(n12885), .S(n12863), .Z(n12886) );
  INV_X1 U14639 ( .A(n12887), .ZN(n12888) );
  MUX2_X1 U14640 ( .A(n14739), .B(n16128), .S(n12884), .Z(n12890) );
  MUX2_X1 U14641 ( .A(n14739), .B(n16128), .S(n12874), .Z(n12889) );
  INV_X1 U14642 ( .A(n12890), .ZN(n12891) );
  MUX2_X1 U14643 ( .A(n14738), .B(n15122), .S(n12874), .Z(n12894) );
  MUX2_X1 U14644 ( .A(n14738), .B(n15122), .S(n12884), .Z(n12892) );
  INV_X1 U14645 ( .A(n12894), .ZN(n12895) );
  MUX2_X1 U14646 ( .A(n14737), .B(n14656), .S(n12884), .Z(n12899) );
  MUX2_X1 U14647 ( .A(n14737), .B(n14656), .S(n12868), .Z(n12896) );
  NAND2_X1 U14648 ( .A1(n12897), .A2(n12896), .ZN(n12903) );
  INV_X1 U14649 ( .A(n12898), .ZN(n12901) );
  INV_X1 U14650 ( .A(n12899), .ZN(n12900) );
  NAND2_X1 U14651 ( .A1(n12901), .A2(n12900), .ZN(n12902) );
  MUX2_X1 U14652 ( .A(n14736), .B(n14669), .S(n12874), .Z(n12905) );
  MUX2_X1 U14653 ( .A(n14736), .B(n14669), .S(n12884), .Z(n12904) );
  INV_X1 U14654 ( .A(n12905), .ZN(n12906) );
  MUX2_X1 U14655 ( .A(n14735), .B(n15104), .S(n13015), .Z(n12908) );
  MUX2_X1 U14656 ( .A(n14735), .B(n15104), .S(n12874), .Z(n12907) );
  MUX2_X1 U14657 ( .A(n14981), .B(n15082), .S(n12868), .Z(n12937) );
  NOR2_X1 U14658 ( .A1(n14981), .A2(n13015), .ZN(n12931) );
  AOI21_X1 U14659 ( .B1(n12937), .B2(n14961), .A(n12931), .ZN(n12910) );
  OR2_X1 U14660 ( .A1(n15075), .A2(n12910), .ZN(n12918) );
  NAND2_X1 U14661 ( .A1(n12937), .A2(n12911), .ZN(n12912) );
  OR2_X1 U14662 ( .A1(n15082), .A2(n12874), .ZN(n12922) );
  NAND2_X1 U14663 ( .A1(n12912), .A2(n12922), .ZN(n12913) );
  NAND2_X1 U14664 ( .A1(n15075), .A2(n12913), .ZN(n12917) );
  NAND2_X1 U14665 ( .A1(n14961), .A2(n13015), .ZN(n12923) );
  OR2_X1 U14666 ( .A1(n15082), .A2(n12923), .ZN(n12916) );
  NOR2_X1 U14667 ( .A1(n14961), .A2(n13015), .ZN(n12932) );
  NAND2_X1 U14668 ( .A1(n12932), .A2(n12914), .ZN(n12915) );
  AND2_X1 U14669 ( .A1(n12916), .A2(n12915), .ZN(n12935) );
  NAND3_X1 U14670 ( .A1(n12918), .A2(n12917), .A3(n12935), .ZN(n12930) );
  MUX2_X1 U14671 ( .A(n14637), .B(n14976), .S(n12868), .Z(n12927) );
  INV_X1 U14672 ( .A(n14637), .ZN(n14962) );
  MUX2_X1 U14673 ( .A(n14962), .B(n15086), .S(n12884), .Z(n12926) );
  NAND2_X1 U14674 ( .A1(n12927), .A2(n12926), .ZN(n12919) );
  MUX2_X1 U14675 ( .A(n15006), .B(n15097), .S(n12868), .Z(n12943) );
  MUX2_X1 U14676 ( .A(n14979), .B(n14995), .S(n12884), .Z(n12944) );
  NAND2_X1 U14677 ( .A1(n12943), .A2(n12944), .ZN(n12920) );
  INV_X1 U14678 ( .A(n12922), .ZN(n12925) );
  INV_X1 U14679 ( .A(n12923), .ZN(n12924) );
  AOI21_X1 U14680 ( .B1(n12937), .B2(n12925), .A(n12924), .ZN(n12941) );
  INV_X1 U14681 ( .A(n12926), .ZN(n12929) );
  INV_X1 U14682 ( .A(n12927), .ZN(n12928) );
  NAND3_X1 U14683 ( .A1(n12930), .A2(n12929), .A3(n12928), .ZN(n12940) );
  NAND2_X1 U14684 ( .A1(n12937), .A2(n12931), .ZN(n12934) );
  INV_X1 U14685 ( .A(n12932), .ZN(n12933) );
  NAND2_X1 U14686 ( .A1(n12934), .A2(n12933), .ZN(n12938) );
  INV_X1 U14687 ( .A(n12935), .ZN(n12936) );
  AOI22_X1 U14688 ( .A1(n7611), .A2(n12938), .B1(n12937), .B2(n12936), .ZN(
        n12939) );
  OAI211_X1 U14689 ( .C1(n7611), .C2(n12941), .A(n12940), .B(n12939), .ZN(
        n12942) );
  INV_X1 U14690 ( .A(n12942), .ZN(n12949) );
  INV_X1 U14691 ( .A(n12943), .ZN(n12946) );
  INV_X1 U14692 ( .A(n12944), .ZN(n12945) );
  NAND3_X1 U14693 ( .A1(n12947), .A2(n12946), .A3(n12945), .ZN(n12948) );
  NAND3_X1 U14694 ( .A1(n12950), .A2(n12949), .A3(n12948), .ZN(n12952) );
  MUX2_X1 U14695 ( .A(n14951), .B(n15069), .S(n12868), .Z(n12953) );
  MUX2_X1 U14696 ( .A(n14951), .B(n15069), .S(n12884), .Z(n12951) );
  INV_X1 U14697 ( .A(n12953), .ZN(n12954) );
  MUX2_X1 U14698 ( .A(n14900), .B(n15064), .S(n12884), .Z(n12957) );
  MUX2_X1 U14699 ( .A(n14900), .B(n15064), .S(n12868), .Z(n12955) );
  NAND2_X1 U14700 ( .A1(n12956), .A2(n12955), .ZN(n12960) );
  INV_X1 U14701 ( .A(n12957), .ZN(n12958) );
  NAND2_X1 U14702 ( .A1(n12960), .A2(n12959), .ZN(n12963) );
  MUX2_X1 U14703 ( .A(n14881), .B(n15057), .S(n12874), .Z(n12964) );
  NAND2_X1 U14704 ( .A1(n12963), .A2(n12964), .ZN(n12962) );
  MUX2_X1 U14705 ( .A(n14881), .B(n15057), .S(n12884), .Z(n12961) );
  INV_X1 U14706 ( .A(n12963), .ZN(n12966) );
  INV_X1 U14707 ( .A(n12964), .ZN(n12965) );
  NAND2_X1 U14708 ( .A1(n12966), .A2(n12965), .ZN(n12967) );
  MUX2_X1 U14709 ( .A(n14899), .B(n15051), .S(n12868), .Z(n12968) );
  MUX2_X1 U14710 ( .A(n14882), .B(n14871), .S(n12868), .Z(n12974) );
  NAND2_X1 U14711 ( .A1(n12973), .A2(n12974), .ZN(n12972) );
  MUX2_X1 U14712 ( .A(n14882), .B(n14871), .S(n13015), .Z(n12971) );
  MUX2_X1 U14713 ( .A(n14857), .B(n15040), .S(n13015), .Z(n12977) );
  MUX2_X1 U14714 ( .A(n15040), .B(n14857), .S(n13015), .Z(n12976) );
  INV_X1 U14715 ( .A(n12977), .ZN(n12978) );
  MUX2_X1 U14716 ( .A(n14734), .B(n15031), .S(n12868), .Z(n12982) );
  NAND2_X1 U14717 ( .A1(n12981), .A2(n12982), .ZN(n12980) );
  MUX2_X1 U14718 ( .A(n14734), .B(n15031), .S(n13015), .Z(n12979) );
  NAND2_X1 U14719 ( .A1(n12980), .A2(n12979), .ZN(n12986) );
  INV_X1 U14720 ( .A(n12981), .ZN(n12984) );
  INV_X1 U14721 ( .A(n12982), .ZN(n12983) );
  NAND2_X1 U14722 ( .A1(n12984), .A2(n12983), .ZN(n12985) );
  INV_X1 U14723 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n12991) );
  NAND2_X1 U14724 ( .A1(n12987), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n12990) );
  NAND2_X1 U14725 ( .A1(n12988), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n12989) );
  OAI211_X1 U14726 ( .C1(n12992), .C2(n12991), .A(n12990), .B(n12989), .ZN(
        n14845) );
  OAI21_X1 U14727 ( .B1(n14845), .B2(n12993), .A(n14733), .ZN(n12996) );
  NAND2_X1 U14728 ( .A1(n13011), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12995) );
  MUX2_X1 U14729 ( .A(n12996), .B(n14851), .S(n12884), .Z(n13000) );
  INV_X1 U14730 ( .A(n14845), .ZN(n13016) );
  OAI21_X1 U14731 ( .B1(n13016), .B2(n12998), .A(n12997), .ZN(n12999) );
  AOI22_X1 U14732 ( .A1(n15028), .A2(n12868), .B1(n14733), .B2(n12999), .ZN(
        n13001) );
  OAI21_X1 U14733 ( .B1(n15170), .B2(n13017), .A(n13002), .ZN(n13003) );
  AND2_X1 U14734 ( .A1(n13004), .A2(n13003), .ZN(n13068) );
  MUX2_X1 U14735 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7178), .Z(n13008) );
  XNOR2_X1 U14736 ( .A(n13008), .B(SI_31_), .ZN(n13009) );
  NAND2_X1 U14737 ( .A1(n14581), .A2(n12089), .ZN(n13013) );
  NAND2_X1 U14738 ( .A1(n13011), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n13012) );
  XNOR2_X1 U14739 ( .A(n15024), .B(n14845), .ZN(n13023) );
  NAND3_X1 U14740 ( .A1(n13014), .A2(n13068), .A3(n13023), .ZN(n13074) );
  NAND2_X1 U14741 ( .A1(n13016), .A2(n13015), .ZN(n13067) );
  INV_X1 U14742 ( .A(n13067), .ZN(n13020) );
  INV_X1 U14743 ( .A(n13068), .ZN(n13018) );
  NAND2_X1 U14744 ( .A1(n7920), .A2(n13017), .ZN(n13060) );
  NAND2_X1 U14745 ( .A1(n13018), .A2(n13060), .ZN(n13065) );
  NAND2_X1 U14746 ( .A1(n14845), .A2(n12874), .ZN(n13064) );
  NOR2_X1 U14747 ( .A1(n15024), .A2(n13064), .ZN(n13019) );
  AOI211_X1 U14748 ( .C1(n13020), .C2(n15024), .A(n13065), .B(n13019), .ZN(
        n13021) );
  NAND2_X1 U14749 ( .A1(n13022), .A2(n13021), .ZN(n13073) );
  XNOR2_X1 U14750 ( .A(n15028), .B(n14733), .ZN(n13057) );
  AND2_X1 U14751 ( .A1(n13025), .A2(n13024), .ZN(n15833) );
  NAND4_X1 U14752 ( .A1(n15833), .A2(n13028), .A3(n13027), .A4(n13026), .ZN(
        n13030) );
  NOR2_X1 U14753 ( .A1(n13030), .A2(n13029), .ZN(n13033) );
  NAND4_X1 U14754 ( .A1(n13034), .A2(n13033), .A3(n13032), .A4(n13031), .ZN(
        n13035) );
  NOR2_X1 U14755 ( .A1(n13036), .A2(n13035), .ZN(n13039) );
  NAND4_X1 U14756 ( .A1(n13040), .A2(n13039), .A3(n13038), .A4(n13037), .ZN(
        n13041) );
  OR4_X1 U14757 ( .A1(n13044), .A2(n13043), .A3(n13042), .A4(n13041), .ZN(
        n13045) );
  OR4_X1 U14758 ( .A1(n13048), .A2(n13047), .A3(n13046), .A4(n13045), .ZN(
        n13051) );
  NOR4_X1 U14759 ( .A1(n13051), .A2(n13050), .A3(n15010), .A4(n13049), .ZN(
        n13053) );
  NAND4_X1 U14760 ( .A1(n13053), .A2(n14939), .A3(n13052), .A4(n14966), .ZN(
        n13054) );
  NOR4_X1 U14761 ( .A1(n14876), .A2(n14918), .A3(n14894), .A4(n13054), .ZN(
        n13056) );
  INV_X1 U14762 ( .A(n13065), .ZN(n13061) );
  NAND2_X1 U14763 ( .A1(n14845), .A2(n13061), .ZN(n13062) );
  NAND2_X1 U14764 ( .A1(n13064), .A2(n13062), .ZN(n13063) );
  OAI21_X1 U14765 ( .B1(n13064), .B2(n13068), .A(n13063), .ZN(n13070) );
  OAI21_X1 U14766 ( .B1(n14845), .B2(n13065), .A(n13067), .ZN(n13066) );
  OAI21_X1 U14767 ( .B1(n13068), .B2(n13067), .A(n13066), .ZN(n13069) );
  MUX2_X1 U14768 ( .A(n13070), .B(n13069), .S(n15024), .Z(n13071) );
  NOR3_X1 U14769 ( .A1(n13075), .A2(n15154), .A3(n15003), .ZN(n13077) );
  OAI21_X1 U14770 ( .B1(n13078), .B2(n15170), .A(P1_B_REG_SCAN_IN), .ZN(n13076) );
  OAI22_X1 U14771 ( .A1(n13079), .A2(n13078), .B1(n13077), .B2(n13076), .ZN(
        P1_U3242) );
  INV_X1 U14772 ( .A(n13080), .ZN(n13081) );
  OAI222_X1 U14773 ( .A1(n8227), .A2(P3_U3151), .B1(n13083), .B2(n15290), .C1(
        n13082), .C2(n13081), .ZN(P3_U3265) );
  XNOR2_X1 U14774 ( .A(n13685), .B(n13084), .ZN(n13091) );
  INV_X1 U14775 ( .A(n13091), .ZN(n13085) );
  NAND2_X1 U14776 ( .A1(n13085), .A2(n13527), .ZN(n13098) );
  INV_X1 U14777 ( .A(n13086), .ZN(n13087) );
  NAND4_X1 U14778 ( .A1(n13097), .A2(n13527), .A3(n13091), .A4(n13087), .ZN(
        n13096) );
  AOI22_X1 U14779 ( .A1(n13686), .A2(n13550), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13089) );
  NAND2_X1 U14780 ( .A1(n13698), .A2(n13529), .ZN(n13088) );
  OAI211_X1 U14781 ( .C1(n13681), .C2(n13519), .A(n13089), .B(n13088), .ZN(
        n13093) );
  NOR4_X1 U14782 ( .A1(n13091), .A2(n13539), .A3(n13698), .A4(n13090), .ZN(
        n13092) );
  AOI211_X1 U14783 ( .C1(n13094), .C2(n13511), .A(n13093), .B(n13092), .ZN(
        n13095) );
  OAI211_X1 U14784 ( .C1(n13098), .C2(n13097), .A(n13096), .B(n13095), .ZN(
        P3_U3160) );
  OAI21_X1 U14785 ( .B1(n8046), .B2(n14226), .A(n13099), .ZN(n13105) );
  NAND3_X1 U14786 ( .A1(n9773), .A2(n7180), .A3(n13101), .ZN(n13104) );
  NAND2_X1 U14787 ( .A1(n13102), .A2(n13351), .ZN(n13103) );
  OAI211_X1 U14788 ( .C1(n13106), .C2(n13105), .A(n13104), .B(n13103), .ZN(
        n13114) );
  NAND2_X1 U14789 ( .A1(n13351), .A2(n13109), .ZN(n13108) );
  NAND2_X1 U14790 ( .A1(n7180), .A2(n14200), .ZN(n13107) );
  NAND2_X1 U14791 ( .A1(n13108), .A2(n13107), .ZN(n13115) );
  NAND2_X1 U14792 ( .A1(n13114), .A2(n13115), .ZN(n13113) );
  NAND2_X1 U14793 ( .A1(n14200), .A2(n13351), .ZN(n13111) );
  NAND2_X1 U14794 ( .A1(n7180), .A2(n13109), .ZN(n13110) );
  NAND2_X1 U14795 ( .A1(n13111), .A2(n13110), .ZN(n13112) );
  NAND2_X1 U14796 ( .A1(n13113), .A2(n13112), .ZN(n13124) );
  INV_X1 U14797 ( .A(n13114), .ZN(n13117) );
  INV_X1 U14798 ( .A(n13115), .ZN(n13116) );
  NAND2_X1 U14799 ( .A1(n13117), .A2(n13116), .ZN(n13123) );
  NAND2_X1 U14800 ( .A1(n14199), .A2(n7180), .ZN(n13119) );
  NAND2_X1 U14801 ( .A1(n15904), .A2(n13351), .ZN(n13118) );
  AND2_X1 U14802 ( .A1(n13119), .A2(n13118), .ZN(n13131) );
  NAND2_X1 U14803 ( .A1(n15904), .A2(n7180), .ZN(n13121) );
  NAND2_X1 U14804 ( .A1(n14199), .A2(n13351), .ZN(n13120) );
  NAND2_X1 U14805 ( .A1(n13121), .A2(n13120), .ZN(n13130) );
  NAND2_X1 U14806 ( .A1(n13131), .A2(n13130), .ZN(n13122) );
  NAND3_X1 U14807 ( .A1(n13124), .A2(n13123), .A3(n13122), .ZN(n13136) );
  NAND2_X1 U14808 ( .A1(n14198), .A2(n7180), .ZN(n13126) );
  NAND2_X1 U14809 ( .A1(n13127), .A2(n13351), .ZN(n13125) );
  NAND2_X1 U14810 ( .A1(n13126), .A2(n13125), .ZN(n13137) );
  AND2_X1 U14811 ( .A1(n13127), .A2(n13360), .ZN(n13129) );
  NAND2_X1 U14812 ( .A1(n13137), .A2(n13138), .ZN(n13135) );
  INV_X1 U14813 ( .A(n13130), .ZN(n13133) );
  INV_X1 U14814 ( .A(n13131), .ZN(n13132) );
  NAND2_X1 U14815 ( .A1(n13133), .A2(n13132), .ZN(n13134) );
  NAND3_X1 U14816 ( .A1(n13136), .A2(n13135), .A3(n13134), .ZN(n13142) );
  INV_X1 U14817 ( .A(n13137), .ZN(n13140) );
  INV_X1 U14818 ( .A(n13138), .ZN(n13139) );
  NAND2_X1 U14819 ( .A1(n13140), .A2(n13139), .ZN(n13141) );
  NAND2_X1 U14820 ( .A1(n13142), .A2(n13141), .ZN(n13148) );
  NAND2_X1 U14821 ( .A1(n13145), .A2(n13360), .ZN(n13144) );
  NAND2_X1 U14822 ( .A1(n14197), .A2(n13351), .ZN(n13143) );
  NAND2_X1 U14823 ( .A1(n13144), .A2(n13143), .ZN(n13147) );
  AOI22_X1 U14824 ( .A1(n13145), .A2(n13351), .B1(n13360), .B2(n14197), .ZN(
        n13146) );
  AOI21_X1 U14825 ( .B1(n13148), .B2(n13147), .A(n13146), .ZN(n13150) );
  NOR2_X1 U14826 ( .A1(n13148), .A2(n13147), .ZN(n13149) );
  NAND2_X1 U14827 ( .A1(n13153), .A2(n7188), .ZN(n13152) );
  NAND2_X1 U14828 ( .A1(n14196), .A2(n13360), .ZN(n13151) );
  NAND2_X1 U14829 ( .A1(n13152), .A2(n13151), .ZN(n13157) );
  NAND2_X1 U14830 ( .A1(n8184), .A2(n13157), .ZN(n13156) );
  AOI22_X1 U14831 ( .A1(n13153), .A2(n7180), .B1(n14196), .B2(n7188), .ZN(
        n13154) );
  INV_X1 U14832 ( .A(n13154), .ZN(n13155) );
  NAND2_X1 U14833 ( .A1(n13156), .A2(n13155), .ZN(n13158) );
  NAND2_X1 U14834 ( .A1(n13158), .A2(n8185), .ZN(n13164) );
  NAND2_X1 U14835 ( .A1(n13161), .A2(n13360), .ZN(n13160) );
  NAND2_X1 U14836 ( .A1(n14195), .A2(n7188), .ZN(n13159) );
  NAND2_X1 U14837 ( .A1(n13160), .A2(n13159), .ZN(n13163) );
  AOI22_X1 U14838 ( .A1(n13161), .A2(n7188), .B1(n13360), .B2(n14195), .ZN(
        n13162) );
  NOR2_X1 U14839 ( .A1(n13164), .A2(n13163), .ZN(n13165) );
  INV_X1 U14840 ( .A(n13165), .ZN(n13166) );
  NAND2_X1 U14841 ( .A1(n13170), .A2(n7188), .ZN(n13169) );
  NAND2_X1 U14842 ( .A1(n14194), .A2(n13360), .ZN(n13168) );
  NAND2_X1 U14843 ( .A1(n13169), .A2(n13168), .ZN(n13172) );
  AOI22_X1 U14844 ( .A1(n13170), .A2(n13360), .B1(n14194), .B2(n7188), .ZN(
        n13171) );
  NAND2_X1 U14845 ( .A1(n13177), .A2(n13360), .ZN(n13174) );
  NAND2_X1 U14846 ( .A1(n14193), .A2(n7188), .ZN(n13173) );
  NAND2_X1 U14847 ( .A1(n13174), .A2(n13173), .ZN(n13175) );
  NAND2_X1 U14848 ( .A1(n13176), .A2(n13175), .ZN(n13181) );
  NAND2_X1 U14849 ( .A1(n13177), .A2(n7188), .ZN(n13178) );
  OAI21_X1 U14850 ( .B1(n13179), .B2(n13351), .A(n13178), .ZN(n13180) );
  NAND2_X1 U14851 ( .A1(n13181), .A2(n13180), .ZN(n13182) );
  NAND2_X1 U14852 ( .A1(n14435), .A2(n7188), .ZN(n13185) );
  NAND2_X1 U14853 ( .A1(n14191), .A2(n13360), .ZN(n13184) );
  NAND2_X1 U14854 ( .A1(n13185), .A2(n13184), .ZN(n13187) );
  AOI22_X1 U14855 ( .A1(n14435), .A2(n13360), .B1(n14191), .B2(n7188), .ZN(
        n13186) );
  NAND2_X1 U14856 ( .A1(n13190), .A2(n13360), .ZN(n13189) );
  NAND2_X1 U14857 ( .A1(n14190), .A2(n7188), .ZN(n13188) );
  NAND2_X1 U14858 ( .A1(n13189), .A2(n13188), .ZN(n13196) );
  NAND2_X1 U14859 ( .A1(n13195), .A2(n13196), .ZN(n13194) );
  NAND2_X1 U14860 ( .A1(n13190), .A2(n7188), .ZN(n13192) );
  NAND2_X1 U14861 ( .A1(n14190), .A2(n13360), .ZN(n13191) );
  NAND2_X1 U14862 ( .A1(n13192), .A2(n13191), .ZN(n13193) );
  NAND2_X1 U14863 ( .A1(n13194), .A2(n13193), .ZN(n13200) );
  INV_X1 U14864 ( .A(n13195), .ZN(n13198) );
  INV_X1 U14865 ( .A(n13196), .ZN(n13197) );
  NAND2_X1 U14866 ( .A1(n13198), .A2(n13197), .ZN(n13199) );
  NAND2_X1 U14867 ( .A1(n13203), .A2(n7188), .ZN(n13202) );
  NAND2_X1 U14868 ( .A1(n14189), .A2(n13360), .ZN(n13201) );
  NAND2_X1 U14869 ( .A1(n13202), .A2(n13201), .ZN(n13205) );
  AOI22_X1 U14870 ( .A1(n13203), .A2(n13360), .B1(n14189), .B2(n7188), .ZN(
        n13204) );
  NAND2_X1 U14871 ( .A1(n13208), .A2(n13360), .ZN(n13207) );
  NAND2_X1 U14872 ( .A1(n14188), .A2(n7188), .ZN(n13206) );
  NAND2_X1 U14873 ( .A1(n13207), .A2(n13206), .ZN(n13212) );
  NAND2_X1 U14874 ( .A1(n13208), .A2(n7188), .ZN(n13209) );
  OAI21_X1 U14875 ( .B1(n13210), .B2(n13351), .A(n13209), .ZN(n13211) );
  INV_X1 U14876 ( .A(n13212), .ZN(n13213) );
  NAND2_X1 U14877 ( .A1(n13216), .A2(n7188), .ZN(n13215) );
  NAND2_X1 U14878 ( .A1(n14187), .A2(n7180), .ZN(n13214) );
  NAND2_X1 U14879 ( .A1(n13215), .A2(n13214), .ZN(n13219) );
  AOI22_X1 U14880 ( .A1(n13216), .A2(n13360), .B1(n14187), .B2(n7188), .ZN(
        n13217) );
  AOI21_X1 U14881 ( .B1(n13220), .B2(n13219), .A(n13217), .ZN(n13218) );
  INV_X1 U14882 ( .A(n13218), .ZN(n13221) );
  NAND2_X1 U14883 ( .A1(n13221), .A2(n7245), .ZN(n13227) );
  NAND2_X1 U14884 ( .A1(n13224), .A2(n13360), .ZN(n13223) );
  NAND2_X1 U14885 ( .A1(n14186), .A2(n7188), .ZN(n13222) );
  NAND2_X1 U14886 ( .A1(n13223), .A2(n13222), .ZN(n13226) );
  AOI22_X1 U14887 ( .A1(n13224), .A2(n7188), .B1(n7180), .B2(n14186), .ZN(
        n13225) );
  NAND2_X1 U14888 ( .A1(n13230), .A2(n7188), .ZN(n13229) );
  NAND2_X1 U14889 ( .A1(n14185), .A2(n7180), .ZN(n13228) );
  NAND2_X1 U14890 ( .A1(n13229), .A2(n13228), .ZN(n13235) );
  NAND2_X1 U14891 ( .A1(n13230), .A2(n13360), .ZN(n13232) );
  NAND2_X1 U14892 ( .A1(n14185), .A2(n7188), .ZN(n13231) );
  NAND2_X1 U14893 ( .A1(n13232), .A2(n13231), .ZN(n13233) );
  NAND2_X1 U14894 ( .A1(n13234), .A2(n13233), .ZN(n13238) );
  INV_X1 U14895 ( .A(n13235), .ZN(n13236) );
  NAND2_X1 U14896 ( .A1(n13238), .A2(n13237), .ZN(n13243) );
  NAND2_X1 U14897 ( .A1(n14526), .A2(n13360), .ZN(n13240) );
  NAND2_X1 U14898 ( .A1(n14184), .A2(n7188), .ZN(n13239) );
  NAND2_X1 U14899 ( .A1(n13240), .A2(n13239), .ZN(n13242) );
  AOI22_X1 U14900 ( .A1(n14526), .A2(n7188), .B1(n7180), .B2(n14184), .ZN(
        n13241) );
  NAND2_X1 U14901 ( .A1(n14577), .A2(n7188), .ZN(n13245) );
  NAND2_X1 U14902 ( .A1(n14183), .A2(n13360), .ZN(n13244) );
  NAND2_X1 U14903 ( .A1(n13245), .A2(n13244), .ZN(n13250) );
  NAND2_X1 U14904 ( .A1(n14577), .A2(n13360), .ZN(n13247) );
  NAND2_X1 U14905 ( .A1(n14183), .A2(n7188), .ZN(n13246) );
  NAND2_X1 U14906 ( .A1(n13247), .A2(n13246), .ZN(n13248) );
  NAND2_X1 U14907 ( .A1(n13249), .A2(n13248), .ZN(n13252) );
  INV_X1 U14908 ( .A(n13250), .ZN(n13251) );
  NAND2_X1 U14909 ( .A1(n14511), .A2(n13360), .ZN(n13254) );
  NAND2_X1 U14910 ( .A1(n14182), .A2(n7188), .ZN(n13253) );
  NAND2_X1 U14911 ( .A1(n13254), .A2(n13253), .ZN(n13256) );
  AOI22_X1 U14912 ( .A1(n14511), .A2(n7188), .B1(n13360), .B2(n14182), .ZN(
        n13255) );
  NAND2_X1 U14913 ( .A1(n14570), .A2(n7188), .ZN(n13258) );
  NAND2_X1 U14914 ( .A1(n14181), .A2(n13360), .ZN(n13257) );
  NAND2_X1 U14915 ( .A1(n13258), .A2(n13257), .ZN(n13264) );
  NAND2_X1 U14916 ( .A1(n13263), .A2(n13264), .ZN(n13262) );
  NAND2_X1 U14917 ( .A1(n14570), .A2(n13360), .ZN(n13260) );
  NAND2_X1 U14918 ( .A1(n14181), .A2(n7188), .ZN(n13259) );
  NAND2_X1 U14919 ( .A1(n13260), .A2(n13259), .ZN(n13261) );
  NAND2_X1 U14920 ( .A1(n13262), .A2(n13261), .ZN(n13268) );
  INV_X1 U14921 ( .A(n13263), .ZN(n13266) );
  INV_X1 U14922 ( .A(n13264), .ZN(n13265) );
  NAND2_X1 U14923 ( .A1(n13266), .A2(n13265), .ZN(n13267) );
  NAND2_X1 U14924 ( .A1(n14502), .A2(n13360), .ZN(n13270) );
  NAND2_X1 U14925 ( .A1(n14180), .A2(n7188), .ZN(n13269) );
  NAND2_X1 U14926 ( .A1(n13270), .A2(n13269), .ZN(n13272) );
  AOI22_X1 U14927 ( .A1(n14502), .A2(n7188), .B1(n13360), .B2(n14180), .ZN(
        n13271) );
  NAND2_X1 U14928 ( .A1(n14361), .A2(n7188), .ZN(n13274) );
  NAND2_X1 U14929 ( .A1(n14179), .A2(n13360), .ZN(n13273) );
  NAND2_X1 U14930 ( .A1(n13274), .A2(n13273), .ZN(n13277) );
  AOI22_X1 U14931 ( .A1(n14361), .A2(n7180), .B1(n14179), .B2(n7188), .ZN(
        n13275) );
  INV_X1 U14932 ( .A(n13276), .ZN(n13279) );
  NAND2_X1 U14933 ( .A1(n13279), .A2(n7240), .ZN(n13284) );
  NAND2_X1 U14934 ( .A1(n14485), .A2(n13360), .ZN(n13281) );
  NAND2_X1 U14935 ( .A1(n14178), .A2(n7188), .ZN(n13280) );
  NAND2_X1 U14936 ( .A1(n14485), .A2(n7188), .ZN(n13282) );
  OAI21_X1 U14937 ( .B1(n14355), .B2(n13351), .A(n13282), .ZN(n13283) );
  NAND2_X1 U14938 ( .A1(n14480), .A2(n7188), .ZN(n13286) );
  NAND2_X1 U14939 ( .A1(n14177), .A2(n13360), .ZN(n13285) );
  NAND2_X1 U14940 ( .A1(n13286), .A2(n13285), .ZN(n13288) );
  AOI22_X1 U14941 ( .A1(n14480), .A2(n7180), .B1(n14177), .B2(n7188), .ZN(
        n13287) );
  NAND2_X1 U14942 ( .A1(n14475), .A2(n7180), .ZN(n13290) );
  NAND2_X1 U14943 ( .A1(n14176), .A2(n7188), .ZN(n13289) );
  NAND2_X1 U14944 ( .A1(n13290), .A2(n13289), .ZN(n13294) );
  NAND2_X1 U14945 ( .A1(n13295), .A2(n13294), .ZN(n13293) );
  NAND2_X1 U14946 ( .A1(n14475), .A2(n7188), .ZN(n13291) );
  OAI21_X1 U14947 ( .B1(n14104), .B2(n13351), .A(n13291), .ZN(n13292) );
  NAND2_X1 U14948 ( .A1(n13293), .A2(n13292), .ZN(n13299) );
  INV_X1 U14949 ( .A(n13294), .ZN(n13297) );
  NAND2_X1 U14950 ( .A1(n13297), .A2(n13296), .ZN(n13298) );
  NAND2_X1 U14951 ( .A1(n13299), .A2(n13298), .ZN(n13305) );
  NAND2_X1 U14952 ( .A1(n14470), .A2(n7188), .ZN(n13301) );
  NAND2_X1 U14953 ( .A1(n14175), .A2(n13360), .ZN(n13300) );
  NAND2_X1 U14954 ( .A1(n13301), .A2(n13300), .ZN(n13304) );
  AOI22_X1 U14955 ( .A1(n14470), .A2(n7180), .B1(n14175), .B2(n7188), .ZN(
        n13302) );
  AOI21_X1 U14956 ( .B1(n13305), .B2(n13304), .A(n13302), .ZN(n13303) );
  NOR2_X1 U14957 ( .A1(n13305), .A2(n13304), .ZN(n13306) );
  INV_X1 U14958 ( .A(n13306), .ZN(n13307) );
  NAND2_X1 U14959 ( .A1(n14277), .A2(n13360), .ZN(n13309) );
  NAND2_X1 U14960 ( .A1(n14174), .A2(n7188), .ZN(n13308) );
  NAND2_X1 U14961 ( .A1(n14277), .A2(n7188), .ZN(n13310) );
  OAI21_X1 U14962 ( .B1(n13311), .B2(n13351), .A(n13310), .ZN(n13312) );
  NAND2_X1 U14963 ( .A1(n14463), .A2(n7188), .ZN(n13314) );
  NAND2_X1 U14964 ( .A1(n14173), .A2(n13360), .ZN(n13313) );
  NAND2_X1 U14965 ( .A1(n13314), .A2(n13313), .ZN(n13316) );
  AOI22_X1 U14966 ( .A1(n14076), .A2(n7180), .B1(n14172), .B2(n7188), .ZN(
        n13339) );
  OAI22_X1 U14967 ( .A1(n14544), .A2(n13360), .B1(n14047), .B2(n13351), .ZN(
        n13338) );
  AOI22_X1 U14968 ( .A1(n14463), .A2(n7180), .B1(n14173), .B2(n7188), .ZN(
        n13315) );
  OR2_X1 U14969 ( .A1(n13318), .A2(n13317), .ZN(n13320) );
  NAND2_X1 U14970 ( .A1(n13330), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13319) );
  INV_X1 U14971 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n14534) );
  NAND2_X1 U14972 ( .A1(n13321), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n13324) );
  NAND2_X1 U14973 ( .A1(n13322), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n13323) );
  OAI211_X1 U14974 ( .C1(n13325), .C2(n14534), .A(n13324), .B(n13323), .ZN(
        n14236) );
  NAND2_X1 U14975 ( .A1(n14236), .A2(n7188), .ZN(n13352) );
  NAND2_X1 U14976 ( .A1(n13326), .A2(n8046), .ZN(n13357) );
  NAND4_X1 U14977 ( .A1(n13352), .A2(n7182), .A3(n13357), .A4(n13407), .ZN(
        n13327) );
  AOI22_X1 U14978 ( .A1(n14232), .A2(n7180), .B1(n14170), .B2(n13327), .ZN(
        n13328) );
  INV_X1 U14979 ( .A(n13328), .ZN(n13346) );
  AOI22_X1 U14980 ( .A1(n14232), .A2(n7188), .B1(n7180), .B2(n14170), .ZN(
        n13345) );
  INV_X1 U14981 ( .A(n14078), .ZN(n14171) );
  AOI22_X1 U14982 ( .A1(n14453), .A2(n7188), .B1(n7180), .B2(n14171), .ZN(
        n13336) );
  OAI22_X1 U14983 ( .A1(n13329), .A2(n13351), .B1(n14078), .B2(n13360), .ZN(
        n13337) );
  AOI22_X1 U14984 ( .A1(n13346), .A2(n13345), .B1(n13336), .B2(n13337), .ZN(
        n13335) );
  NAND2_X1 U14985 ( .A1(n13330), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n13331) );
  INV_X1 U14986 ( .A(n14236), .ZN(n13333) );
  OR2_X1 U14987 ( .A1(n14233), .A2(n13333), .ZN(n13359) );
  NAND2_X1 U14988 ( .A1(n14233), .A2(n13333), .ZN(n13334) );
  NAND2_X1 U14989 ( .A1(n13359), .A2(n13334), .ZN(n13404) );
  NOR2_X1 U14990 ( .A1(n13335), .A2(n13404), .ZN(n13342) );
  INV_X1 U14991 ( .A(n13404), .ZN(n13344) );
  INV_X1 U14992 ( .A(n13336), .ZN(n13341) );
  INV_X1 U14993 ( .A(n13337), .ZN(n13340) );
  AOI22_X1 U14994 ( .A1(n13341), .A2(n13340), .B1(n13339), .B2(n13338), .ZN(
        n13343) );
  AOI21_X1 U14995 ( .B1(n13344), .B2(n13343), .A(n13342), .ZN(n13348) );
  NOR2_X1 U14996 ( .A1(n13346), .A2(n13345), .ZN(n13347) );
  INV_X1 U14997 ( .A(n13368), .ZN(n13356) );
  AND2_X1 U14998 ( .A1(n13352), .A2(n13351), .ZN(n13353) );
  OAI211_X1 U14999 ( .C1(n7183), .C2(n13405), .A(n13354), .B(n13407), .ZN(
        n13355) );
  NOR3_X1 U15000 ( .A1(n13356), .A2(n13362), .A3(n13355), .ZN(n13420) );
  OAI21_X1 U15001 ( .B1(n13358), .B2(n14226), .A(n13357), .ZN(n13365) );
  INV_X1 U15002 ( .A(n13359), .ZN(n13361) );
  AOI21_X1 U15003 ( .B1(n13361), .B2(n13360), .A(n13406), .ZN(n13364) );
  INV_X1 U15004 ( .A(n13362), .ZN(n13366) );
  OR2_X1 U15005 ( .A1(n13366), .A2(n13365), .ZN(n13363) );
  OAI211_X1 U15006 ( .C1(n13368), .C2(n13365), .A(n13364), .B(n13363), .ZN(
        n13419) );
  NAND3_X1 U15007 ( .A1(n13368), .A2(n13367), .A3(n13366), .ZN(n13417) );
  XNOR2_X1 U15008 ( .A(n14232), .B(n14170), .ZN(n13401) );
  NOR2_X1 U15009 ( .A1(n13372), .A2(n13371), .ZN(n13375) );
  NAND4_X1 U15010 ( .A1(n13376), .A2(n13375), .A3(n13374), .A4(n13373), .ZN(
        n13377) );
  OR4_X1 U15011 ( .A1(n13380), .A2(n13379), .A3(n13378), .A4(n13377), .ZN(
        n13381) );
  NOR2_X1 U15012 ( .A1(n13382), .A2(n13381), .ZN(n13385) );
  NAND4_X1 U15013 ( .A1(n13386), .A2(n13385), .A3(n13384), .A4(n13383), .ZN(
        n13387) );
  NOR2_X1 U15014 ( .A1(n13388), .A2(n13387), .ZN(n13391) );
  NAND4_X1 U15015 ( .A1(n13391), .A2(n13392), .A3(n13390), .A4(n13389), .ZN(
        n13393) );
  NOR2_X1 U15016 ( .A1(n14250), .A2(n13399), .ZN(n13400) );
  NAND3_X1 U15017 ( .A1(n13401), .A2(n13400), .A3(n14262), .ZN(n13402) );
  AND4_X1 U15018 ( .A1(n7215), .A2(n7183), .A3(n13412), .A4(n13405), .ZN(
        n13416) );
  NOR4_X1 U15019 ( .A1(n15406), .A2(n13408), .A3(n14354), .A4(n13407), .ZN(
        n13409) );
  AOI211_X1 U15020 ( .C1(n13412), .C2(n13411), .A(n13410), .B(n13409), .ZN(
        n13413) );
  AOI21_X1 U15021 ( .B1(n13417), .B2(n13416), .A(n13415), .ZN(n13418) );
  OAI21_X1 U15022 ( .B1(n13420), .B2(n13419), .A(n13418), .ZN(P2_U3328) );
  XNOR2_X1 U15023 ( .A(n13537), .B(n13536), .ZN(n13421) );
  NAND2_X1 U15024 ( .A1(n13421), .A2(n13527), .ZN(n13425) );
  NAND2_X1 U15025 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(P3_U3151), .ZN(n15749)
         );
  OAI21_X1 U15026 ( .B1(n13519), .B2(n13877), .A(n15749), .ZN(n13423) );
  NOR2_X1 U15027 ( .A1(n13531), .A2(n13883), .ZN(n13422) );
  AOI211_X1 U15028 ( .C1(n13529), .C2(n13566), .A(n13423), .B(n13422), .ZN(
        n13424) );
  OAI211_X1 U15029 ( .C1(n13554), .C2(n14014), .A(n13425), .B(n13424), .ZN(
        P3_U3155) );
  AOI21_X1 U15030 ( .B1(n13559), .B2(n13426), .A(n7192), .ZN(n13431) );
  AOI22_X1 U15031 ( .A1(n13735), .A2(n13529), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13428) );
  NAND2_X1 U15032 ( .A1(n13744), .A2(n13550), .ZN(n13427) );
  OAI211_X1 U15033 ( .C1(n13738), .C2(n13519), .A(n13428), .B(n13427), .ZN(
        n13429) );
  AOI21_X1 U15034 ( .B1(n13739), .B2(n13511), .A(n13429), .ZN(n13430) );
  OAI21_X1 U15035 ( .B1(n13431), .B2(n13539), .A(n13430), .ZN(P3_U3156) );
  INV_X1 U15036 ( .A(n13432), .ZN(n13995) );
  OAI211_X1 U15037 ( .C1(n13434), .C2(n13433), .A(n13440), .B(n13527), .ZN(
        n13438) );
  NAND2_X1 U15038 ( .A1(n13563), .A2(n13529), .ZN(n13435) );
  NAND2_X1 U15039 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13658)
         );
  OAI211_X1 U15040 ( .C1(n13799), .C2(n13519), .A(n13435), .B(n13658), .ZN(
        n13436) );
  AOI21_X1 U15041 ( .B1(n13802), .B2(n13550), .A(n13436), .ZN(n13437) );
  OAI211_X1 U15042 ( .C1(n13995), .C2(n13554), .A(n13438), .B(n13437), .ZN(
        P3_U3159) );
  NAND2_X1 U15043 ( .A1(n13440), .A2(n13439), .ZN(n13492) );
  NAND2_X1 U15044 ( .A1(n13492), .A2(n13441), .ZN(n13443) );
  NAND2_X1 U15045 ( .A1(n13443), .A2(n13442), .ZN(n13445) );
  XNOR2_X1 U15046 ( .A(n13445), .B(n13444), .ZN(n13450) );
  OAI22_X1 U15047 ( .A1(n13799), .A2(n13548), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15253), .ZN(n13447) );
  NOR2_X1 U15048 ( .A1(n13771), .A2(n13519), .ZN(n13446) );
  AOI211_X1 U15049 ( .C1(n13773), .C2(n13550), .A(n13447), .B(n13446), .ZN(
        n13449) );
  NAND2_X1 U15050 ( .A1(n13772), .A2(n13511), .ZN(n13448) );
  OAI211_X1 U15051 ( .C1(n13450), .C2(n13539), .A(n13449), .B(n13448), .ZN(
        P3_U3163) );
  INV_X1 U15052 ( .A(n13451), .ZN(n13483) );
  INV_X1 U15053 ( .A(n13452), .ZN(n13454) );
  NOR3_X1 U15054 ( .A1(n13483), .A2(n13454), .A3(n13453), .ZN(n13457) );
  INV_X1 U15055 ( .A(n13455), .ZN(n13456) );
  OAI21_X1 U15056 ( .B1(n13457), .B2(n13456), .A(n13527), .ZN(n13461) );
  OAI22_X1 U15057 ( .A1(n13738), .A2(n13548), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15250), .ZN(n13459) );
  NOR2_X1 U15058 ( .A1(n13712), .A2(n13519), .ZN(n13458) );
  AOI211_X1 U15059 ( .C1(n13715), .C2(n13550), .A(n13459), .B(n13458), .ZN(
        n13460) );
  OAI211_X1 U15060 ( .C1(n13971), .C2(n13554), .A(n13461), .B(n13460), .ZN(
        P3_U3165) );
  XNOR2_X1 U15061 ( .A(n13462), .B(n13859), .ZN(n13463) );
  XNOR2_X1 U15062 ( .A(n13464), .B(n13463), .ZN(n13469) );
  NAND2_X1 U15063 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n15787)
         );
  OAI21_X1 U15064 ( .B1(n13519), .B2(n13843), .A(n15787), .ZN(n13465) );
  AOI21_X1 U15065 ( .B1(n13529), .B2(n13565), .A(n13465), .ZN(n13466) );
  OAI21_X1 U15066 ( .B1(n13848), .B2(n13531), .A(n13466), .ZN(n13467) );
  AOI21_X1 U15067 ( .B1(n13847), .B2(n13511), .A(n13467), .ZN(n13468) );
  OAI21_X1 U15068 ( .B1(n13469), .B2(n13539), .A(n13468), .ZN(P3_U3166) );
  XNOR2_X1 U15069 ( .A(n13470), .B(n13564), .ZN(n13471) );
  XNOR2_X1 U15070 ( .A(n13472), .B(n13471), .ZN(n13478) );
  INV_X1 U15071 ( .A(n13473), .ZN(n13828) );
  NOR2_X1 U15072 ( .A1(n15356), .A2(P3_STATE_REG_SCAN_IN), .ZN(n15805) );
  AOI21_X1 U15073 ( .B1(n13563), .B2(n13546), .A(n15805), .ZN(n13474) );
  OAI21_X1 U15074 ( .B1(n13823), .B2(n13548), .A(n13474), .ZN(n13476) );
  NOR2_X1 U15075 ( .A1(n14003), .A2(n13554), .ZN(n13475) );
  AOI211_X1 U15076 ( .C1(n13828), .C2(n13550), .A(n13476), .B(n13475), .ZN(
        n13477) );
  OAI21_X1 U15077 ( .B1(n13478), .B2(n13539), .A(n13477), .ZN(P3_U3168) );
  INV_X1 U15078 ( .A(n13480), .ZN(n13482) );
  NOR3_X1 U15079 ( .A1(n7192), .A2(n13482), .A3(n13481), .ZN(n13484) );
  OAI21_X1 U15080 ( .B1(n13484), .B2(n13483), .A(n13527), .ZN(n13489) );
  AOI22_X1 U15081 ( .A1(n13559), .A2(n13529), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13485) );
  OAI21_X1 U15082 ( .B1(n13486), .B2(n13519), .A(n13485), .ZN(n13487) );
  AOI21_X1 U15083 ( .B1(n13729), .B2(n13550), .A(n13487), .ZN(n13488) );
  OAI211_X1 U15084 ( .C1(n13975), .C2(n13554), .A(n13489), .B(n13488), .ZN(
        P3_U3169) );
  XNOR2_X1 U15085 ( .A(n13490), .B(n13561), .ZN(n13491) );
  XNOR2_X1 U15086 ( .A(n13492), .B(n13491), .ZN(n13497) );
  AOI22_X1 U15087 ( .A1(n13560), .A2(n13546), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13494) );
  NAND2_X1 U15088 ( .A1(n13550), .A2(n13789), .ZN(n13493) );
  OAI211_X1 U15089 ( .C1(n13811), .C2(n13548), .A(n13494), .B(n13493), .ZN(
        n13495) );
  AOI21_X1 U15090 ( .B1(n13788), .B2(n13511), .A(n13495), .ZN(n13496) );
  OAI21_X1 U15091 ( .B1(n13497), .B2(n13539), .A(n13496), .ZN(P3_U3173) );
  XOR2_X1 U15092 ( .A(n13499), .B(n13498), .Z(n13504) );
  INV_X1 U15093 ( .A(n16095), .ZN(n15400) );
  NOR2_X1 U15094 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15272), .ZN(n15728) );
  NOR2_X1 U15095 ( .A1(n15393), .A2(n13548), .ZN(n13500) );
  AOI211_X1 U15096 ( .C1(n13546), .C2(n13860), .A(n15728), .B(n13500), .ZN(
        n13501) );
  OAI21_X1 U15097 ( .B1(n15397), .B2(n13531), .A(n13501), .ZN(n13502) );
  AOI21_X1 U15098 ( .B1(n15400), .B2(n13511), .A(n13502), .ZN(n13503) );
  OAI21_X1 U15099 ( .B1(n13504), .B2(n13539), .A(n13503), .ZN(P3_U3174) );
  INV_X1 U15100 ( .A(n13505), .ZN(n13506) );
  AOI21_X1 U15101 ( .B1(n13735), .B2(n13507), .A(n13506), .ZN(n13513) );
  AOI22_X1 U15102 ( .A1(n13560), .A2(n13529), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13509) );
  NAND2_X1 U15103 ( .A1(n13550), .A2(n13758), .ZN(n13508) );
  OAI211_X1 U15104 ( .C1(n13752), .C2(n13519), .A(n13509), .B(n13508), .ZN(
        n13510) );
  AOI21_X1 U15105 ( .B1(n13757), .B2(n13511), .A(n13510), .ZN(n13512) );
  OAI21_X1 U15106 ( .B1(n13513), .B2(n13539), .A(n13512), .ZN(P3_U3175) );
  AOI21_X1 U15107 ( .B1(n13516), .B2(n13515), .A(n13539), .ZN(n13518) );
  NAND2_X1 U15108 ( .A1(n13518), .A2(n13517), .ZN(n13523) );
  NAND2_X1 U15109 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13645)
         );
  OAI21_X1 U15110 ( .B1(n13519), .B2(n13811), .A(n13645), .ZN(n13521) );
  NOR2_X1 U15111 ( .A1(n13531), .A2(n13814), .ZN(n13520) );
  AOI211_X1 U15112 ( .C1(n13529), .C2(n13564), .A(n13521), .B(n13520), .ZN(
        n13522) );
  OAI211_X1 U15113 ( .C1(n13999), .C2(n13554), .A(n13523), .B(n13522), .ZN(
        P3_U3178) );
  OAI21_X1 U15114 ( .B1(n13526), .B2(n13525), .A(n13524), .ZN(n13528) );
  NAND2_X1 U15115 ( .A1(n13528), .A2(n13527), .ZN(n13535) );
  INV_X1 U15116 ( .A(n13702), .ZN(n13532) );
  AOI22_X1 U15117 ( .A1(n13725), .A2(n13529), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13530) );
  OAI21_X1 U15118 ( .B1(n13532), .B2(n13531), .A(n13530), .ZN(n13533) );
  AOI21_X1 U15119 ( .B1(n13698), .B2(n13546), .A(n13533), .ZN(n13534) );
  OAI211_X1 U15120 ( .C1(n13704), .C2(n13554), .A(n13535), .B(n13534), .ZN(
        P3_U3180) );
  NAND2_X1 U15121 ( .A1(n13537), .A2(n13536), .ZN(n13543) );
  NAND2_X1 U15122 ( .A1(n13543), .A2(n13538), .ZN(n13541) );
  AOI21_X1 U15123 ( .B1(n13541), .B2(n13540), .A(n13539), .ZN(n13545) );
  NAND2_X1 U15124 ( .A1(n13543), .A2(n13542), .ZN(n13544) );
  NAND2_X1 U15125 ( .A1(n13545), .A2(n13544), .ZN(n13553) );
  INV_X1 U15126 ( .A(n13863), .ZN(n13551) );
  NOR2_X1 U15127 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8195), .ZN(n15770) );
  AOI21_X1 U15128 ( .B1(n13546), .B2(n13859), .A(n15770), .ZN(n13547) );
  OAI21_X1 U15129 ( .B1(n15391), .B2(n13548), .A(n13547), .ZN(n13549) );
  AOI21_X1 U15130 ( .B1(n13551), .B2(n13550), .A(n13549), .ZN(n13552) );
  OAI211_X1 U15131 ( .C1(n13554), .C2(n13943), .A(n13553), .B(n13552), .ZN(
        P3_U3181) );
  MUX2_X1 U15132 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n13960), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U15133 ( .A(n13556), .B(P3_DATAO_REG_30__SCAN_IN), .S(n13577), .Z(
        P3_U3521) );
  MUX2_X1 U15134 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n7408), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U15135 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n13698), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15136 ( .A(n13557), .B(P3_DATAO_REG_26__SCAN_IN), .S(n13577), .Z(
        P3_U3517) );
  MUX2_X1 U15137 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n13725), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U15138 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n13558), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U15139 ( .A(n13559), .B(P3_DATAO_REG_23__SCAN_IN), .S(n13577), .Z(
        P3_U3514) );
  MUX2_X1 U15140 ( .A(n13735), .B(P3_DATAO_REG_22__SCAN_IN), .S(n13577), .Z(
        P3_U3513) );
  MUX2_X1 U15141 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n13560), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U15142 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13561), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15143 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n13562), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U15144 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13563), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15145 ( .A(n13564), .B(P3_DATAO_REG_17__SCAN_IN), .S(n13577), .Z(
        P3_U3508) );
  MUX2_X1 U15146 ( .A(n13859), .B(P3_DATAO_REG_16__SCAN_IN), .S(n13577), .Z(
        P3_U3507) );
  MUX2_X1 U15147 ( .A(n13565), .B(P3_DATAO_REG_15__SCAN_IN), .S(n13577), .Z(
        P3_U3506) );
  MUX2_X1 U15148 ( .A(n13860), .B(P3_DATAO_REG_14__SCAN_IN), .S(n13577), .Z(
        P3_U3505) );
  MUX2_X1 U15149 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n13566), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U15150 ( .A(n13567), .B(P3_DATAO_REG_12__SCAN_IN), .S(n13577), .Z(
        P3_U3503) );
  MUX2_X1 U15151 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n13568), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U15152 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n13569), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15153 ( .A(n13570), .B(P3_DATAO_REG_9__SCAN_IN), .S(n13577), .Z(
        P3_U3500) );
  MUX2_X1 U15154 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n13571), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U15155 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n13572), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U15156 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n13573), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15157 ( .A(n13574), .B(P3_DATAO_REG_5__SCAN_IN), .S(n13577), .Z(
        P3_U3496) );
  MUX2_X1 U15158 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n13575), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U15159 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n15874), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15160 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n13576), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15161 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n15875), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15162 ( .A(n13578), .B(P3_DATAO_REG_0__SCAN_IN), .S(n13577), .Z(
        P3_U3491) );
  INV_X1 U15163 ( .A(n13579), .ZN(n13581) );
  NAND2_X1 U15164 ( .A1(n13581), .A2(n13580), .ZN(n13582) );
  NAND2_X1 U15165 ( .A1(n13583), .A2(n13582), .ZN(n15696) );
  MUX2_X1 U15166 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13664), .Z(n13584) );
  XNOR2_X1 U15167 ( .A(n13584), .B(n15697), .ZN(n15695) );
  NAND2_X1 U15168 ( .A1(n15696), .A2(n15695), .ZN(n13587) );
  INV_X1 U15169 ( .A(n13584), .ZN(n13585) );
  NAND2_X1 U15170 ( .A1(n13585), .A2(n15697), .ZN(n13586) );
  NAND2_X1 U15171 ( .A1(n13587), .A2(n13586), .ZN(n15714) );
  NOR2_X1 U15172 ( .A1(n15711), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n13588) );
  NOR2_X1 U15173 ( .A1(n15711), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n13589) );
  MUX2_X1 U15174 ( .A(n15709), .B(n15720), .S(n13664), .Z(n15715) );
  MUX2_X1 U15175 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13664), .Z(n13593) );
  XNOR2_X1 U15176 ( .A(n13593), .B(n15739), .ZN(n15731) );
  INV_X1 U15177 ( .A(n13614), .ZN(n13591) );
  INV_X1 U15178 ( .A(n13631), .ZN(n13590) );
  MUX2_X1 U15179 ( .A(n13591), .B(n13590), .S(n13664), .Z(n15732) );
  AND2_X1 U15180 ( .A1(n15731), .A2(n15732), .ZN(n13592) );
  NAND2_X1 U15181 ( .A1(n15733), .A2(n13592), .ZN(n15735) );
  INV_X1 U15182 ( .A(n13593), .ZN(n13594) );
  NAND2_X1 U15183 ( .A1(n13594), .A2(n15739), .ZN(n13595) );
  MUX2_X1 U15184 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n13664), .Z(n13596) );
  INV_X1 U15185 ( .A(n13634), .ZN(n15757) );
  XNOR2_X1 U15186 ( .A(n13596), .B(n15757), .ZN(n15752) );
  NAND2_X1 U15187 ( .A1(n15753), .A2(n15752), .ZN(n15751) );
  NAND2_X1 U15188 ( .A1(n13596), .A2(n13634), .ZN(n13597) );
  NAND2_X1 U15189 ( .A1(n15751), .A2(n13597), .ZN(n13598) );
  INV_X1 U15190 ( .A(n16152), .ZN(n13636) );
  XNOR2_X1 U15191 ( .A(n13598), .B(n13636), .ZN(n15768) );
  MUX2_X1 U15192 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n13664), .Z(n15769) );
  NAND2_X1 U15193 ( .A1(n15768), .A2(n15769), .ZN(n13600) );
  NAND2_X1 U15194 ( .A1(n13598), .A2(n16152), .ZN(n13599) );
  NAND2_X1 U15195 ( .A1(n13600), .A2(n13599), .ZN(n15790) );
  MUX2_X1 U15196 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n13664), .Z(n13601) );
  XNOR2_X1 U15197 ( .A(n13601), .B(n13639), .ZN(n15789) );
  INV_X1 U15198 ( .A(n13601), .ZN(n13602) );
  NAND2_X1 U15199 ( .A1(n13602), .A2(n15795), .ZN(n13603) );
  NAND2_X1 U15200 ( .A1(n15792), .A2(n13603), .ZN(n15812) );
  MUX2_X1 U15201 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13664), .Z(n13604) );
  NAND2_X1 U15202 ( .A1(n13604), .A2(n13641), .ZN(n13607) );
  INV_X1 U15203 ( .A(n13604), .ZN(n13605) );
  INV_X1 U15204 ( .A(n13641), .ZN(n15816) );
  NAND2_X1 U15205 ( .A1(n13605), .A2(n15816), .ZN(n13606) );
  NAND2_X1 U15206 ( .A1(n13607), .A2(n13606), .ZN(n15813) );
  NAND2_X1 U15207 ( .A1(n15809), .A2(n13607), .ZN(n13662) );
  XNOR2_X1 U15208 ( .A(n13662), .B(n13647), .ZN(n13609) );
  INV_X1 U15209 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13934) );
  MUX2_X1 U15210 ( .A(n13815), .B(n13934), .S(n13664), .Z(n13608) );
  NAND2_X1 U15211 ( .A1(n13609), .A2(n13608), .ZN(n13660) );
  OAI21_X1 U15212 ( .B1(n13609), .B2(n13608), .A(n13660), .ZN(n13610) );
  INV_X1 U15213 ( .A(n13610), .ZN(n13650) );
  NOR2_X1 U15214 ( .A1(n15739), .A2(n13615), .ZN(n13616) );
  AOI22_X1 U15215 ( .A1(P3_REG2_REG_14__SCAN_IN), .A2(n15757), .B1(n13634), 
        .B2(n13884), .ZN(n15747) );
  NOR2_X1 U15216 ( .A1(n13636), .A2(n13617), .ZN(n13618) );
  NOR2_X1 U15217 ( .A1(n13618), .A2(n15765), .ZN(n15786) );
  NAND2_X1 U15218 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n13639), .ZN(n13619) );
  OAI21_X1 U15219 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n13639), .A(n13619), 
        .ZN(n15785) );
  INV_X1 U15220 ( .A(n15802), .ZN(n13624) );
  OR2_X1 U15221 ( .A1(n13620), .A2(n15816), .ZN(n13623) );
  NAND2_X1 U15222 ( .A1(n13661), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n13651) );
  NAND2_X1 U15223 ( .A1(n13647), .A2(n13815), .ZN(n13621) );
  NAND2_X1 U15224 ( .A1(n13651), .A2(n13621), .ZN(n13622) );
  AND3_X1 U15225 ( .A1(n13624), .A2(n13623), .A3(n13622), .ZN(n13626) );
  OAI21_X1 U15226 ( .B1(n13652), .B2(n13626), .A(n13625), .ZN(n13649) );
  NOR2_X1 U15227 ( .A1(n15697), .A2(n13629), .ZN(n13630) );
  NOR2_X1 U15228 ( .A1(n8487), .A2(n15704), .ZN(n15703) );
  NOR2_X1 U15229 ( .A1(n13630), .A2(n15703), .ZN(n15721) );
  NOR2_X1 U15230 ( .A1(n15739), .A2(n13632), .ZN(n13633) );
  NOR2_X1 U15231 ( .A1(n13633), .A2(n15740), .ZN(n15760) );
  XNOR2_X1 U15232 ( .A(n13634), .B(P3_REG1_REG_14__SCAN_IN), .ZN(n15759) );
  NOR2_X1 U15233 ( .A1(n15760), .A2(n15759), .ZN(n15758) );
  NOR2_X1 U15234 ( .A1(n13636), .A2(n13635), .ZN(n13637) );
  XNOR2_X1 U15235 ( .A(n13636), .B(n13635), .ZN(n15779) );
  NOR2_X1 U15236 ( .A1(n15778), .A2(n15779), .ZN(n15777) );
  NAND2_X1 U15237 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n13639), .ZN(n13638) );
  OAI21_X1 U15238 ( .B1(n13639), .B2(P3_REG1_REG_16__SCAN_IN), .A(n13638), 
        .ZN(n15796) );
  NAND2_X1 U15239 ( .A1(n13661), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n13654) );
  NAND2_X1 U15240 ( .A1(n13647), .A2(n13934), .ZN(n13642) );
  AND2_X1 U15241 ( .A1(n13654), .A2(n13642), .ZN(n13643) );
  INV_X1 U15242 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15637) );
  OAI21_X1 U15243 ( .B1(n15808), .B2(n15637), .A(n13645), .ZN(n13646) );
  OAI211_X1 U15244 ( .C1(n13650), .C2(n15811), .A(n13649), .B(n13648), .ZN(
        P3_U3200) );
  XNOR2_X1 U15245 ( .A(n13656), .B(n13653), .ZN(n13663) );
  NAND2_X1 U15246 ( .A1(n13655), .A2(n13654), .ZN(n13657) );
  XNOR2_X1 U15247 ( .A(n13656), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13665) );
  NAND2_X1 U15248 ( .A1(n15771), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n13659) );
  OAI21_X1 U15249 ( .B1(n13662), .B2(n13661), .A(n13660), .ZN(n13667) );
  MUX2_X1 U15250 ( .A(n7672), .B(n13665), .S(n13664), .Z(n13666) );
  XNOR2_X1 U15251 ( .A(n13667), .B(n13666), .ZN(n13668) );
  NOR2_X1 U15252 ( .A1(n13668), .A2(n15811), .ZN(n13669) );
  AOI211_X1 U15253 ( .C1(n13960), .C2(n13959), .A(n13853), .B(n13671), .ZN(
        n13674) );
  NOR2_X1 U15254 ( .A1(n15899), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n13672) );
  OAI22_X1 U15255 ( .A1(n13962), .A2(n13882), .B1(n13674), .B2(n13672), .ZN(
        P3_U3202) );
  NOR2_X1 U15256 ( .A1(n15899), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n13673) );
  OAI22_X1 U15257 ( .A1(n13675), .A2(n13882), .B1(n13674), .B2(n13673), .ZN(
        P3_U3203) );
  OAI211_X1 U15258 ( .C1(n13677), .C2(n13685), .A(n13676), .B(n15881), .ZN(
        n13680) );
  OR2_X1 U15259 ( .A1(n13678), .A2(n15392), .ZN(n13679) );
  OAI211_X1 U15260 ( .C1(n13681), .C2(n15390), .A(n13680), .B(n13679), .ZN(
        n13891) );
  INV_X1 U15261 ( .A(n13891), .ZN(n13690) );
  NAND2_X1 U15262 ( .A1(n7766), .A2(n13682), .ZN(n13684) );
  AOI22_X1 U15263 ( .A1(n13686), .A2(n13829), .B1(n13853), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n13687) );
  OAI21_X1 U15264 ( .B1(n13966), .B2(n13882), .A(n13687), .ZN(n13688) );
  AOI21_X1 U15265 ( .B1(n13892), .B2(n13887), .A(n13688), .ZN(n13689) );
  OAI21_X1 U15266 ( .B1(n13690), .B2(n13853), .A(n13689), .ZN(P3_U3205) );
  INV_X1 U15267 ( .A(n13691), .ZN(n13697) );
  AOI22_X1 U15268 ( .A1(n13692), .A2(n13829), .B1(n13853), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13693) );
  OAI21_X1 U15269 ( .B1(n13898), .B2(n13882), .A(n13693), .ZN(n13694) );
  AOI21_X1 U15270 ( .B1(n13695), .B2(n13792), .A(n13694), .ZN(n13696) );
  OAI21_X1 U15271 ( .B1(n13697), .B2(n13853), .A(n13696), .ZN(P3_U3206) );
  XNOR2_X1 U15272 ( .A(n7286), .B(n13701), .ZN(n13699) );
  AOI222_X1 U15273 ( .A1(n15881), .A2(n13699), .B1(n13698), .B2(n15873), .C1(
        n13725), .C2(n15876), .ZN(n13902) );
  XOR2_X1 U15274 ( .A(n13701), .B(n13700), .Z(n13900) );
  AOI22_X1 U15275 ( .A1(n13702), .A2(n13829), .B1(n13853), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13703) );
  OAI21_X1 U15276 ( .B1(n13704), .B2(n13882), .A(n13703), .ZN(n13705) );
  AOI21_X1 U15277 ( .B1(n13900), .B2(n13887), .A(n13705), .ZN(n13706) );
  OAI21_X1 U15278 ( .B1(n13902), .B2(n13853), .A(n13706), .ZN(P3_U3207) );
  XNOR2_X1 U15279 ( .A(n13708), .B(n13707), .ZN(n13904) );
  INV_X1 U15280 ( .A(n13904), .ZN(n13719) );
  AOI211_X1 U15281 ( .C1(n13711), .C2(n13710), .A(n13874), .B(n13709), .ZN(
        n13714) );
  OAI22_X1 U15282 ( .A1(n13712), .A2(n15390), .B1(n13738), .B2(n15392), .ZN(
        n13713) );
  OR2_X1 U15283 ( .A1(n13714), .A2(n13713), .ZN(n13903) );
  AOI22_X1 U15284 ( .A1(n13715), .A2(n13829), .B1(n13853), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n13716) );
  OAI21_X1 U15285 ( .B1(n13971), .B2(n13882), .A(n13716), .ZN(n13717) );
  AOI21_X1 U15286 ( .B1(n13903), .B2(n15899), .A(n13717), .ZN(n13718) );
  OAI21_X1 U15287 ( .B1(n13868), .B2(n13719), .A(n13718), .ZN(P3_U3208) );
  INV_X1 U15288 ( .A(n13722), .ZN(n13720) );
  XNOR2_X1 U15289 ( .A(n13721), .B(n13720), .ZN(n13907) );
  INV_X1 U15290 ( .A(n13907), .ZN(n13733) );
  OAI21_X1 U15291 ( .B1(n13723), .B2(n13722), .A(n15881), .ZN(n13728) );
  NOR2_X1 U15292 ( .A1(n13752), .A2(n15392), .ZN(n13724) );
  AOI21_X1 U15293 ( .B1(n13725), .B2(n15873), .A(n13724), .ZN(n13726) );
  OAI21_X1 U15294 ( .B1(n13728), .B2(n13727), .A(n13726), .ZN(n13909) );
  AOI22_X1 U15295 ( .A1(n13729), .A2(n13829), .B1(n13853), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n13730) );
  OAI21_X1 U15296 ( .B1(n13975), .B2(n13882), .A(n13730), .ZN(n13731) );
  AOI21_X1 U15297 ( .B1(n13909), .B2(n15899), .A(n13731), .ZN(n13732) );
  OAI21_X1 U15298 ( .B1(n13868), .B2(n13733), .A(n13732), .ZN(P3_U3209) );
  OAI211_X1 U15299 ( .C1(n7416), .C2(n13740), .A(n15881), .B(n13734), .ZN(
        n13737) );
  NAND2_X1 U15300 ( .A1(n13735), .A2(n15876), .ZN(n13736) );
  OAI211_X1 U15301 ( .C1(n13738), .C2(n15390), .A(n13737), .B(n13736), .ZN(
        n13912) );
  INV_X1 U15302 ( .A(n13739), .ZN(n13979) );
  NAND2_X1 U15303 ( .A1(n13741), .A2(n13740), .ZN(n13742) );
  AND2_X1 U15304 ( .A1(n13743), .A2(n13742), .ZN(n13913) );
  NAND2_X1 U15305 ( .A1(n13913), .A2(n13887), .ZN(n13746) );
  AOI22_X1 U15306 ( .A1(n13744), .A2(n13829), .B1(n13853), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n13745) );
  OAI211_X1 U15307 ( .C1(n13979), .C2(n13882), .A(n13746), .B(n13745), .ZN(
        n13747) );
  AOI21_X1 U15308 ( .B1(n13912), .B2(n15899), .A(n13747), .ZN(n13748) );
  INV_X1 U15309 ( .A(n13748), .ZN(P3_U3210) );
  XNOR2_X1 U15310 ( .A(n13749), .B(n13751), .ZN(n13756) );
  OAI21_X1 U15311 ( .B1(n7231), .B2(n13751), .A(n13750), .ZN(n13917) );
  OAI22_X1 U15312 ( .A1(n13752), .A2(n15390), .B1(n13783), .B2(n15392), .ZN(
        n13753) );
  AOI21_X1 U15313 ( .B1(n13917), .B2(n13754), .A(n13753), .ZN(n13755) );
  OAI21_X1 U15314 ( .B1(n13756), .B2(n13874), .A(n13755), .ZN(n13916) );
  INV_X1 U15315 ( .A(n13916), .ZN(n13762) );
  INV_X1 U15316 ( .A(n13757), .ZN(n13983) );
  AOI22_X1 U15317 ( .A1(n13853), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n13758), 
        .B2(n13829), .ZN(n13759) );
  OAI21_X1 U15318 ( .B1(n13983), .B2(n13882), .A(n13759), .ZN(n13760) );
  AOI21_X1 U15319 ( .B1(n13917), .B2(n13792), .A(n13760), .ZN(n13761) );
  OAI21_X1 U15320 ( .B1(n13762), .B2(n13853), .A(n13761), .ZN(P3_U3211) );
  NAND2_X1 U15321 ( .A1(n13801), .A2(n13764), .ZN(n13766) );
  NAND2_X1 U15322 ( .A1(n13766), .A2(n13765), .ZN(n13767) );
  XOR2_X1 U15323 ( .A(n13769), .B(n13767), .Z(n13921) );
  INV_X1 U15324 ( .A(n13921), .ZN(n13777) );
  AOI21_X1 U15325 ( .B1(n13769), .B2(n13768), .A(n7241), .ZN(n13770) );
  OAI222_X1 U15326 ( .A1(n15390), .A2(n13771), .B1(n15392), .B2(n13799), .C1(
        n13874), .C2(n13770), .ZN(n13920) );
  INV_X1 U15327 ( .A(n13772), .ZN(n13987) );
  AOI22_X1 U15328 ( .A1(n13853), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n13829), 
        .B2(n13773), .ZN(n13774) );
  OAI21_X1 U15329 ( .B1(n13987), .B2(n13882), .A(n13774), .ZN(n13775) );
  AOI21_X1 U15330 ( .B1(n13920), .B2(n15899), .A(n13775), .ZN(n13776) );
  OAI21_X1 U15331 ( .B1(n13777), .B2(n13868), .A(n13776), .ZN(P3_U3212) );
  NAND2_X1 U15332 ( .A1(n13801), .A2(n13796), .ZN(n13779) );
  NAND2_X1 U15333 ( .A1(n13779), .A2(n13778), .ZN(n13780) );
  XNOR2_X1 U15334 ( .A(n13780), .B(n13781), .ZN(n13787) );
  XNOR2_X1 U15335 ( .A(n13782), .B(n13781), .ZN(n13785) );
  OAI22_X1 U15336 ( .A1(n13783), .A2(n15390), .B1(n13811), .B2(n15392), .ZN(
        n13784) );
  AOI21_X1 U15337 ( .B1(n13785), .B2(n15881), .A(n13784), .ZN(n13786) );
  OAI21_X1 U15338 ( .B1(n15886), .B2(n13787), .A(n13786), .ZN(n13924) );
  INV_X1 U15339 ( .A(n13924), .ZN(n13794) );
  INV_X1 U15340 ( .A(n13787), .ZN(n13925) );
  INV_X1 U15341 ( .A(n13788), .ZN(n13991) );
  AOI22_X1 U15342 ( .A1(n13853), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n13829), 
        .B2(n13789), .ZN(n13790) );
  OAI21_X1 U15343 ( .B1(n13991), .B2(n13882), .A(n13790), .ZN(n13791) );
  AOI21_X1 U15344 ( .B1(n13925), .B2(n13792), .A(n13791), .ZN(n13793) );
  OAI21_X1 U15345 ( .B1(n13794), .B2(n13853), .A(n13793), .ZN(P3_U3213) );
  NAND2_X1 U15346 ( .A1(n13807), .A2(n13795), .ZN(n13797) );
  XNOR2_X1 U15347 ( .A(n13797), .B(n13796), .ZN(n13798) );
  OAI222_X1 U15348 ( .A1(n15390), .A2(n13799), .B1(n15392), .B2(n13824), .C1(
        n13874), .C2(n13798), .ZN(n13928) );
  INV_X1 U15349 ( .A(n13928), .ZN(n13806) );
  XNOR2_X1 U15350 ( .A(n13801), .B(n13800), .ZN(n13929) );
  AOI22_X1 U15351 ( .A1(n13853), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n13829), 
        .B2(n13802), .ZN(n13803) );
  OAI21_X1 U15352 ( .B1(n13995), .B2(n13882), .A(n13803), .ZN(n13804) );
  AOI21_X1 U15353 ( .B1(n13929), .B2(n13887), .A(n13804), .ZN(n13805) );
  OAI21_X1 U15354 ( .B1(n13806), .B2(n13853), .A(n13805), .ZN(P3_U3214) );
  INV_X1 U15355 ( .A(n13807), .ZN(n13808) );
  AOI21_X1 U15356 ( .B1(n13812), .B2(n13809), .A(n13808), .ZN(n13810) );
  OAI222_X1 U15357 ( .A1(n15390), .A2(n13811), .B1(n15392), .B2(n13843), .C1(
        n13874), .C2(n13810), .ZN(n13932) );
  INV_X1 U15358 ( .A(n13932), .ZN(n13819) );
  XNOR2_X1 U15359 ( .A(n13813), .B(n13812), .ZN(n13933) );
  NOR2_X1 U15360 ( .A1(n13999), .A2(n13882), .ZN(n13817) );
  OAI22_X1 U15361 ( .A1(n15899), .A2(n13815), .B1(n13814), .B2(n15892), .ZN(
        n13816) );
  AOI211_X1 U15362 ( .C1(n13933), .C2(n13887), .A(n13817), .B(n13816), .ZN(
        n13818) );
  OAI21_X1 U15363 ( .B1(n13819), .B2(n13853), .A(n13818), .ZN(P3_U3215) );
  XNOR2_X1 U15364 ( .A(n13821), .B(n13820), .ZN(n13822) );
  OAI222_X1 U15365 ( .A1(n15390), .A2(n13824), .B1(n15392), .B2(n13823), .C1(
        n13822), .C2(n13874), .ZN(n13936) );
  INV_X1 U15366 ( .A(n13936), .ZN(n13833) );
  OAI21_X1 U15367 ( .B1(n13827), .B2(n13826), .A(n13825), .ZN(n13937) );
  AOI22_X1 U15368 ( .A1(n13853), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n13829), 
        .B2(n13828), .ZN(n13830) );
  OAI21_X1 U15369 ( .B1(n14003), .B2(n13882), .A(n13830), .ZN(n13831) );
  AOI21_X1 U15370 ( .B1(n13937), .B2(n13887), .A(n13831), .ZN(n13832) );
  OAI21_X1 U15371 ( .B1(n13833), .B2(n13853), .A(n13832), .ZN(P3_U3216) );
  OR2_X1 U15372 ( .A1(n15389), .A2(n13834), .ZN(n13836) );
  NAND2_X1 U15373 ( .A1(n13836), .A2(n13835), .ZN(n13857) );
  NAND2_X1 U15374 ( .A1(n13857), .A2(n13837), .ZN(n13839) );
  NAND2_X1 U15375 ( .A1(n13839), .A2(n13838), .ZN(n13841) );
  XNOR2_X1 U15376 ( .A(n13841), .B(n13840), .ZN(n13842) );
  OAI222_X1 U15377 ( .A1(n15390), .A2(n13843), .B1(n15392), .B2(n13877), .C1(
        n13874), .C2(n13842), .ZN(n13939) );
  INV_X1 U15378 ( .A(n13939), .ZN(n13854) );
  OAI21_X1 U15379 ( .B1(n13846), .B2(n13845), .A(n13844), .ZN(n13940) );
  INV_X1 U15380 ( .A(n13847), .ZN(n14007) );
  NOR2_X1 U15381 ( .A1(n14007), .A2(n13882), .ZN(n13851) );
  OAI22_X1 U15382 ( .A1(n15899), .A2(n13849), .B1(n13848), .B2(n15892), .ZN(
        n13850) );
  AOI211_X1 U15383 ( .C1(n13940), .C2(n13887), .A(n13851), .B(n13850), .ZN(
        n13852) );
  OAI21_X1 U15384 ( .B1(n13854), .B2(n13853), .A(n13852), .ZN(P3_U3217) );
  XNOR2_X1 U15385 ( .A(n13855), .B(n13856), .ZN(n13945) );
  XNOR2_X1 U15386 ( .A(n13857), .B(n13856), .ZN(n13858) );
  NAND2_X1 U15387 ( .A1(n13858), .A2(n15881), .ZN(n13862) );
  AOI22_X1 U15388 ( .A1(n15876), .A2(n13860), .B1(n13859), .B2(n15873), .ZN(
        n13861) );
  NAND2_X1 U15389 ( .A1(n13862), .A2(n13861), .ZN(n13947) );
  NAND2_X1 U15390 ( .A1(n13947), .A2(n15899), .ZN(n13867) );
  INV_X1 U15391 ( .A(n13943), .ZN(n13865) );
  OAI22_X1 U15392 ( .A1(n15899), .A2(n15767), .B1(n13863), .B2(n15892), .ZN(
        n13864) );
  AOI21_X1 U15393 ( .B1(n13865), .B2(n15399), .A(n13864), .ZN(n13866) );
  OAI211_X1 U15394 ( .C1(n13945), .C2(n13868), .A(n13867), .B(n13866), .ZN(
        P3_U3218) );
  OR2_X1 U15395 ( .A1(n15389), .A2(n13869), .ZN(n13871) );
  NAND2_X1 U15396 ( .A1(n13871), .A2(n13870), .ZN(n13873) );
  XNOR2_X1 U15397 ( .A(n13873), .B(n13872), .ZN(n13875) );
  OAI222_X1 U15398 ( .A1(n15390), .A2(n13877), .B1(n15392), .B2(n13876), .C1(
        n13875), .C2(n13874), .ZN(n13949) );
  INV_X1 U15399 ( .A(n13949), .ZN(n13889) );
  NAND2_X1 U15400 ( .A1(n13879), .A2(n13878), .ZN(n13881) );
  XNOR2_X1 U15401 ( .A(n13881), .B(n13880), .ZN(n13950) );
  NOR2_X1 U15402 ( .A1(n14014), .A2(n13882), .ZN(n13886) );
  OAI22_X1 U15403 ( .A1(n15899), .A2(n13884), .B1(n13883), .B2(n15892), .ZN(
        n13885) );
  AOI211_X1 U15404 ( .C1(n13950), .C2(n13887), .A(n13886), .B(n13885), .ZN(
        n13888) );
  OAI21_X1 U15405 ( .B1(n13889), .B2(n13853), .A(n13888), .ZN(P3_U3219) );
  NAND2_X1 U15406 ( .A1(n16155), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n13890) );
  NAND3_X1 U15407 ( .A1(n13960), .A2(n16101), .A3(n13959), .ZN(n16157) );
  OAI211_X1 U15408 ( .C1(n13962), .C2(n16154), .A(n13890), .B(n16157), .ZN(
        P3_U3490) );
  INV_X1 U15409 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13893) );
  AOI21_X1 U15410 ( .B1(n13892), .B2(n13955), .A(n13891), .ZN(n13963) );
  MUX2_X1 U15411 ( .A(n13893), .B(n13963), .S(n16101), .Z(n13894) );
  OAI21_X1 U15412 ( .B1(n13966), .B2(n16154), .A(n13894), .ZN(P3_U3487) );
  INV_X1 U15413 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13896) );
  MUX2_X1 U15414 ( .A(n13896), .B(n13895), .S(n16101), .Z(n13897) );
  OAI21_X1 U15415 ( .B1(n13898), .B2(n16154), .A(n13897), .ZN(P3_U3486) );
  AOI22_X1 U15416 ( .A1(n13900), .A2(n13955), .B1(n13954), .B2(n13899), .ZN(
        n13901) );
  NAND2_X1 U15417 ( .A1(n13902), .A2(n13901), .ZN(n13967) );
  MUX2_X1 U15418 ( .A(P3_REG1_REG_26__SCAN_IN), .B(n13967), .S(n16101), .Z(
        P3_U3485) );
  INV_X1 U15419 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13905) );
  AOI21_X1 U15420 ( .B1(n13904), .B2(n13955), .A(n13903), .ZN(n13968) );
  MUX2_X1 U15421 ( .A(n13905), .B(n13968), .S(n16101), .Z(n13906) );
  OAI21_X1 U15422 ( .B1(n13971), .B2(n16154), .A(n13906), .ZN(P3_U3484) );
  INV_X1 U15423 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13910) );
  AND2_X1 U15424 ( .A1(n13907), .A2(n13955), .ZN(n13908) );
  NOR2_X1 U15425 ( .A1(n13909), .A2(n13908), .ZN(n13972) );
  MUX2_X1 U15426 ( .A(n13910), .B(n13972), .S(n16101), .Z(n13911) );
  OAI21_X1 U15427 ( .B1(n13975), .B2(n16154), .A(n13911), .ZN(P3_U3483) );
  INV_X1 U15428 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13914) );
  AOI21_X1 U15429 ( .B1(n13913), .B2(n13955), .A(n13912), .ZN(n13976) );
  MUX2_X1 U15430 ( .A(n13914), .B(n13976), .S(n16101), .Z(n13915) );
  OAI21_X1 U15431 ( .B1(n13979), .B2(n16154), .A(n13915), .ZN(P3_U3482) );
  INV_X1 U15432 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13918) );
  AOI21_X1 U15433 ( .B1(n16082), .B2(n13917), .A(n13916), .ZN(n13980) );
  MUX2_X1 U15434 ( .A(n13918), .B(n13980), .S(n16101), .Z(n13919) );
  OAI21_X1 U15435 ( .B1(n13983), .B2(n16154), .A(n13919), .ZN(P3_U3481) );
  INV_X1 U15436 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13922) );
  AOI21_X1 U15437 ( .B1(n13955), .B2(n13921), .A(n13920), .ZN(n13984) );
  MUX2_X1 U15438 ( .A(n13922), .B(n13984), .S(n16101), .Z(n13923) );
  OAI21_X1 U15439 ( .B1(n13987), .B2(n16154), .A(n13923), .ZN(P3_U3480) );
  INV_X1 U15440 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13926) );
  AOI21_X1 U15441 ( .B1(n16082), .B2(n13925), .A(n13924), .ZN(n13988) );
  MUX2_X1 U15442 ( .A(n13926), .B(n13988), .S(n16101), .Z(n13927) );
  OAI21_X1 U15443 ( .B1(n13991), .B2(n16154), .A(n13927), .ZN(P3_U3479) );
  AOI21_X1 U15444 ( .B1(n13955), .B2(n13929), .A(n13928), .ZN(n13992) );
  MUX2_X1 U15445 ( .A(n13930), .B(n13992), .S(n16101), .Z(n13931) );
  OAI21_X1 U15446 ( .B1(n13995), .B2(n16154), .A(n13931), .ZN(P3_U3478) );
  AOI21_X1 U15447 ( .B1(n13933), .B2(n13955), .A(n13932), .ZN(n13996) );
  MUX2_X1 U15448 ( .A(n13934), .B(n13996), .S(n16101), .Z(n13935) );
  OAI21_X1 U15449 ( .B1(n13999), .B2(n16154), .A(n13935), .ZN(P3_U3477) );
  AOI21_X1 U15450 ( .B1(n13955), .B2(n13937), .A(n13936), .ZN(n14000) );
  MUX2_X1 U15451 ( .A(n15819), .B(n14000), .S(n16101), .Z(n13938) );
  OAI21_X1 U15452 ( .B1(n16154), .B2(n14003), .A(n13938), .ZN(P3_U3476) );
  AOI21_X1 U15453 ( .B1(n13955), .B2(n13940), .A(n13939), .ZN(n14004) );
  MUX2_X1 U15454 ( .A(n13941), .B(n14004), .S(n16101), .Z(n13942) );
  OAI21_X1 U15455 ( .B1(n14007), .B2(n16154), .A(n13942), .ZN(P3_U3475) );
  OAI22_X1 U15456 ( .A1(n13945), .A2(n13944), .B1(n16096), .B2(n13943), .ZN(
        n13946) );
  NOR2_X1 U15457 ( .A1(n13947), .A2(n13946), .ZN(n14008) );
  MUX2_X1 U15458 ( .A(n15778), .B(n14008), .S(n16101), .Z(n13948) );
  INV_X1 U15459 ( .A(n13948), .ZN(P3_U3474) );
  AOI21_X1 U15460 ( .B1(n13950), .B2(n13955), .A(n13949), .ZN(n14011) );
  MUX2_X1 U15461 ( .A(n13951), .B(n14011), .S(n16101), .Z(n13952) );
  OAI21_X1 U15462 ( .B1(n16154), .B2(n14014), .A(n13952), .ZN(P3_U3473) );
  AOI22_X1 U15463 ( .A1(n13956), .A2(n13955), .B1(n13954), .B2(n13953), .ZN(
        n13957) );
  NAND2_X1 U15464 ( .A1(n13958), .A2(n13957), .ZN(n14015) );
  MUX2_X1 U15465 ( .A(P3_REG1_REG_10__SCAN_IN), .B(n14015), .S(n16101), .Z(
        P3_U3469) );
  NAND2_X1 U15466 ( .A1(n16160), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n13961) );
  NAND3_X1 U15467 ( .A1(n13960), .A2(n16104), .A3(n13959), .ZN(n16163) );
  OAI211_X1 U15468 ( .C1(n13962), .C2(n16159), .A(n13961), .B(n16163), .ZN(
        P3_U3458) );
  INV_X1 U15469 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13964) );
  MUX2_X1 U15470 ( .A(n13964), .B(n13963), .S(n16104), .Z(n13965) );
  MUX2_X1 U15471 ( .A(P3_REG0_REG_26__SCAN_IN), .B(n13967), .S(n16104), .Z(
        P3_U3453) );
  INV_X1 U15472 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13969) );
  MUX2_X1 U15473 ( .A(n13969), .B(n13968), .S(n16104), .Z(n13970) );
  OAI21_X1 U15474 ( .B1(n13971), .B2(n16159), .A(n13970), .ZN(P3_U3452) );
  INV_X1 U15475 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13973) );
  MUX2_X1 U15476 ( .A(n13973), .B(n13972), .S(n16104), .Z(n13974) );
  OAI21_X1 U15477 ( .B1(n13975), .B2(n16159), .A(n13974), .ZN(P3_U3451) );
  INV_X1 U15478 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13977) );
  MUX2_X1 U15479 ( .A(n13977), .B(n13976), .S(n16104), .Z(n13978) );
  OAI21_X1 U15480 ( .B1(n13979), .B2(n16159), .A(n13978), .ZN(P3_U3450) );
  INV_X1 U15481 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13981) );
  MUX2_X1 U15482 ( .A(n13981), .B(n13980), .S(n16104), .Z(n13982) );
  OAI21_X1 U15483 ( .B1(n13983), .B2(n16159), .A(n13982), .ZN(P3_U3449) );
  INV_X1 U15484 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13985) );
  MUX2_X1 U15485 ( .A(n13985), .B(n13984), .S(n16104), .Z(n13986) );
  OAI21_X1 U15486 ( .B1(n13987), .B2(n16159), .A(n13986), .ZN(P3_U3448) );
  INV_X1 U15487 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13989) );
  MUX2_X1 U15488 ( .A(n13989), .B(n13988), .S(n16104), .Z(n13990) );
  OAI21_X1 U15489 ( .B1(n13991), .B2(n16159), .A(n13990), .ZN(P3_U3447) );
  MUX2_X1 U15490 ( .A(n13993), .B(n13992), .S(n16104), .Z(n13994) );
  OAI21_X1 U15491 ( .B1(n13995), .B2(n16159), .A(n13994), .ZN(P3_U3446) );
  MUX2_X1 U15492 ( .A(n13997), .B(n13996), .S(n16104), .Z(n13998) );
  OAI21_X1 U15493 ( .B1(n13999), .B2(n16159), .A(n13998), .ZN(P3_U3444) );
  INV_X1 U15494 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n14001) );
  MUX2_X1 U15495 ( .A(n14001), .B(n14000), .S(n16104), .Z(n14002) );
  OAI21_X1 U15496 ( .B1(n16159), .B2(n14003), .A(n14002), .ZN(P3_U3441) );
  INV_X1 U15497 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n14005) );
  MUX2_X1 U15498 ( .A(n14005), .B(n14004), .S(n16104), .Z(n14006) );
  OAI21_X1 U15499 ( .B1(n14007), .B2(n16159), .A(n14006), .ZN(P3_U3438) );
  INV_X1 U15500 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n14009) );
  MUX2_X1 U15501 ( .A(n14009), .B(n14008), .S(n16104), .Z(n14010) );
  INV_X1 U15502 ( .A(n14010), .ZN(P3_U3435) );
  INV_X1 U15503 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n14012) );
  MUX2_X1 U15504 ( .A(n14012), .B(n14011), .S(n16104), .Z(n14013) );
  OAI21_X1 U15505 ( .B1(n16159), .B2(n14014), .A(n14013), .ZN(P3_U3432) );
  MUX2_X1 U15506 ( .A(P3_REG0_REG_10__SCAN_IN), .B(n14015), .S(n16104), .Z(
        P3_U3420) );
  MUX2_X1 U15507 ( .A(n14017), .B(P3_D_REG_0__SCAN_IN), .S(n14016), .Z(
        P3_U3376) );
  NAND3_X1 U15508 ( .A1(n14018), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n14020) );
  OAI22_X1 U15509 ( .A1(n14021), .A2(n14020), .B1(n14019), .B2(n13083), .ZN(
        n14022) );
  AOI21_X1 U15510 ( .B1(n14023), .B2(n16149), .A(n14022), .ZN(n14024) );
  INV_X1 U15511 ( .A(n14024), .ZN(P3_U3264) );
  MUX2_X1 U15512 ( .A(n14025), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  NAND2_X1 U15513 ( .A1(n14174), .A2(n14416), .ZN(n14039) );
  INV_X1 U15514 ( .A(n14039), .ZN(n14042) );
  XNOR2_X1 U15515 ( .A(n14277), .B(n14043), .ZN(n14041) );
  AND2_X1 U15516 ( .A1(n14027), .A2(n14026), .ZN(n14028) );
  XNOR2_X1 U15517 ( .A(n14480), .B(n14043), .ZN(n14030) );
  XNOR2_X1 U15518 ( .A(n14475), .B(n14032), .ZN(n14105) );
  NAND2_X1 U15519 ( .A1(n14176), .A2(n14416), .ZN(n14033) );
  NOR2_X1 U15520 ( .A1(n14105), .A2(n14033), .ZN(n14038) );
  AOI21_X1 U15521 ( .B1(n14105), .B2(n14033), .A(n14038), .ZN(n14117) );
  XNOR2_X1 U15522 ( .A(n14470), .B(n14043), .ZN(n14034) );
  AND2_X1 U15523 ( .A1(n14175), .A2(n14416), .ZN(n14035) );
  NAND2_X1 U15524 ( .A1(n14034), .A2(n14035), .ZN(n14040) );
  INV_X1 U15525 ( .A(n14034), .ZN(n14153) );
  INV_X1 U15526 ( .A(n14035), .ZN(n14036) );
  NAND2_X1 U15527 ( .A1(n14153), .A2(n14036), .ZN(n14037) );
  AND2_X1 U15528 ( .A1(n14040), .A2(n14037), .ZN(n14102) );
  XNOR2_X1 U15529 ( .A(n14041), .B(n14039), .ZN(n14154) );
  XNOR2_X1 U15530 ( .A(n14463), .B(n14043), .ZN(n14072) );
  AND2_X1 U15531 ( .A1(n14173), .A2(n14416), .ZN(n14044) );
  NAND2_X1 U15532 ( .A1(n14072), .A2(n14044), .ZN(n14085) );
  OAI21_X1 U15533 ( .B1(n14072), .B2(n14044), .A(n14085), .ZN(n14045) );
  OR2_X1 U15534 ( .A1(n14047), .A2(n14356), .ZN(n14049) );
  NAND2_X1 U15535 ( .A1(n14174), .A2(n14137), .ZN(n14048) );
  NAND2_X1 U15536 ( .A1(n14049), .A2(n14048), .ZN(n14260) );
  OAI22_X1 U15537 ( .A1(n14267), .A2(n14161), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14050), .ZN(n14051) );
  AOI21_X1 U15538 ( .B1(n14260), .B2(n14165), .A(n14051), .ZN(n14052) );
  OAI211_X1 U15539 ( .C1(n7375), .C2(n14162), .A(n14053), .B(n14052), .ZN(
        P2_U3186) );
  INV_X1 U15540 ( .A(n14054), .ZN(n14061) );
  AOI22_X1 U15541 ( .A1(n14055), .A2(n14115), .B1(n14063), .B2(n14177), .ZN(
        n14060) );
  AOI22_X1 U15542 ( .A1(n14176), .A2(n14139), .B1(n14137), .B2(n14178), .ZN(
        n14320) );
  INV_X1 U15543 ( .A(n14056), .ZN(n14327) );
  AOI22_X1 U15544 ( .A1(n14327), .A2(n14141), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14057) );
  OAI21_X1 U15545 ( .B1(n14320), .B2(n14144), .A(n14057), .ZN(n14058) );
  AOI21_X1 U15546 ( .B1(n14480), .B2(n14150), .A(n14058), .ZN(n14059) );
  OAI21_X1 U15547 ( .B1(n14061), .B2(n14060), .A(n14059), .ZN(P2_U3188) );
  INV_X1 U15548 ( .A(n14570), .ZN(n14071) );
  OAI21_X1 U15549 ( .B1(n14145), .B2(n14062), .A(n14115), .ZN(n14066) );
  NAND3_X1 U15550 ( .A1(n14064), .A2(n14063), .A3(n14182), .ZN(n14065) );
  NAND2_X1 U15551 ( .A1(n14066), .A2(n14065), .ZN(n14067) );
  NAND2_X1 U15552 ( .A1(n14127), .A2(n14067), .ZN(n14070) );
  AND2_X1 U15553 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n14223) );
  AOI22_X1 U15554 ( .A1(n14180), .A2(n14139), .B1(n14137), .B2(n14182), .ZN(
        n14395) );
  NOR2_X1 U15555 ( .A1(n14395), .A2(n14144), .ZN(n14068) );
  AOI211_X1 U15556 ( .C1(n14141), .C2(n14386), .A(n14223), .B(n14068), .ZN(
        n14069) );
  OAI211_X1 U15557 ( .C1(n14071), .C2(n14162), .A(n14070), .B(n14069), .ZN(
        P2_U3191) );
  INV_X1 U15558 ( .A(n14072), .ZN(n14073) );
  NOR3_X1 U15559 ( .A1(n14073), .A2(n14159), .A3(n14152), .ZN(n14074) );
  AOI21_X1 U15560 ( .B1(n14075), .B2(n14115), .A(n14074), .ZN(n14090) );
  MUX2_X1 U15561 ( .A(n14076), .B(n14250), .S(n14416), .Z(n14077) );
  XNOR2_X1 U15562 ( .A(n14077), .B(n14043), .ZN(n14089) );
  OR2_X1 U15563 ( .A1(n14078), .A2(n14356), .ZN(n14080) );
  NAND2_X1 U15564 ( .A1(n14173), .A2(n14137), .ZN(n14079) );
  NAND2_X1 U15565 ( .A1(n14080), .A2(n14079), .ZN(n14247) );
  OAI22_X1 U15566 ( .A1(n14082), .A2(n14161), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14081), .ZN(n14084) );
  NOR2_X1 U15567 ( .A1(n14544), .A2(n14162), .ZN(n14083) );
  AOI211_X1 U15568 ( .C1(n14165), .C2(n14247), .A(n14084), .B(n14083), .ZN(
        n14088) );
  AOI21_X1 U15569 ( .B1(n7309), .B2(n7311), .A(n14168), .ZN(n14094) );
  NOR3_X1 U15570 ( .A1(n14091), .A2(n14353), .A3(n14152), .ZN(n14093) );
  OAI21_X1 U15571 ( .B1(n14094), .B2(n14093), .A(n14092), .ZN(n14101) );
  OAI22_X1 U15572 ( .A1(n14161), .A2(n14362), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14095), .ZN(n14098) );
  NOR2_X1 U15573 ( .A1(n14096), .A2(n14353), .ZN(n14097) );
  AOI211_X1 U15574 ( .C1(n14099), .C2(n14178), .A(n14098), .B(n14097), .ZN(
        n14100) );
  OAI211_X1 U15575 ( .C1(n14562), .C2(n14162), .A(n14101), .B(n14100), .ZN(
        P2_U3195) );
  INV_X1 U15576 ( .A(n14102), .ZN(n14103) );
  AOI21_X1 U15577 ( .B1(n7212), .B2(n14103), .A(n14168), .ZN(n14108) );
  NOR3_X1 U15578 ( .A1(n14105), .A2(n14104), .A3(n14152), .ZN(n14107) );
  OAI21_X1 U15579 ( .B1(n14108), .B2(n14107), .A(n14106), .ZN(n14114) );
  NAND2_X1 U15580 ( .A1(n14174), .A2(n14139), .ZN(n14110) );
  NAND2_X1 U15581 ( .A1(n14176), .A2(n14137), .ZN(n14109) );
  NAND2_X1 U15582 ( .A1(n14110), .A2(n14109), .ZN(n14291) );
  OAI22_X1 U15583 ( .A1(n14296), .A2(n14161), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14111), .ZN(n14112) );
  AOI21_X1 U15584 ( .B1(n14291), .B2(n14165), .A(n14112), .ZN(n14113) );
  OAI211_X1 U15585 ( .C1(n7693), .C2(n14162), .A(n14114), .B(n14113), .ZN(
        P2_U3197) );
  OAI211_X1 U15586 ( .C1(n14117), .C2(n14116), .A(n7212), .B(n14115), .ZN(
        n14123) );
  OAI22_X1 U15587 ( .A1(n14158), .A2(n14356), .B1(n14118), .B2(n14354), .ZN(
        n14307) );
  INV_X1 U15588 ( .A(n14313), .ZN(n14120) );
  OAI22_X1 U15589 ( .A1(n14120), .A2(n14161), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14119), .ZN(n14121) );
  AOI21_X1 U15590 ( .B1(n14307), .B2(n14165), .A(n14121), .ZN(n14122) );
  OAI211_X1 U15591 ( .C1(n7691), .C2(n14162), .A(n14123), .B(n14122), .ZN(
        P2_U3201) );
  NOR3_X1 U15592 ( .A1(n14125), .A2(n14124), .A3(n14152), .ZN(n14129) );
  AOI21_X1 U15593 ( .B1(n14127), .B2(n14126), .A(n14168), .ZN(n14128) );
  OAI21_X1 U15594 ( .B1(n14129), .B2(n14128), .A(n7309), .ZN(n14136) );
  NAND2_X1 U15595 ( .A1(n14179), .A2(n14139), .ZN(n14131) );
  NAND2_X1 U15596 ( .A1(n14181), .A2(n14137), .ZN(n14130) );
  NAND2_X1 U15597 ( .A1(n14131), .A2(n14130), .ZN(n14371) );
  INV_X1 U15598 ( .A(n14377), .ZN(n14133) );
  OAI22_X1 U15599 ( .A1(n14161), .A2(n14133), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14132), .ZN(n14134) );
  AOI21_X1 U15600 ( .B1(n14371), .B2(n14165), .A(n14134), .ZN(n14135) );
  OAI211_X1 U15601 ( .C1(n14567), .C2(n14162), .A(n14136), .B(n14135), .ZN(
        P2_U3205) );
  AND2_X1 U15602 ( .A1(n14183), .A2(n14137), .ZN(n14138) );
  AOI21_X1 U15603 ( .B1(n14181), .B2(n14139), .A(n14138), .ZN(n14410) );
  INV_X1 U15604 ( .A(n14414), .ZN(n14140) );
  NAND2_X1 U15605 ( .A1(n14141), .A2(n14140), .ZN(n14142) );
  OAI211_X1 U15606 ( .C1(n14144), .C2(n14410), .A(n14143), .B(n14142), .ZN(
        n14149) );
  AOI211_X1 U15607 ( .C1(n14147), .C2(n14146), .A(n14168), .B(n14145), .ZN(
        n14148) );
  AOI211_X1 U15608 ( .C1(n14511), .C2(n14150), .A(n14149), .B(n14148), .ZN(
        n14151) );
  INV_X1 U15609 ( .A(n14151), .ZN(P2_U3210) );
  NOR2_X1 U15610 ( .A1(n14106), .A2(n14168), .ZN(n14157) );
  NOR3_X1 U15611 ( .A1(n14153), .A2(n14158), .A3(n14152), .ZN(n14156) );
  INV_X1 U15612 ( .A(n14154), .ZN(n14155) );
  OAI21_X1 U15613 ( .B1(n14157), .B2(n14156), .A(n14155), .ZN(n14167) );
  OAI22_X1 U15614 ( .A1(n14159), .A2(n14356), .B1(n14158), .B2(n14354), .ZN(
        n14284) );
  OAI22_X1 U15615 ( .A1(n14278), .A2(n14161), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14160), .ZN(n14164) );
  NOR2_X1 U15616 ( .A1(n14551), .A2(n14162), .ZN(n14163) );
  AOI211_X1 U15617 ( .C1(n14165), .C2(n14284), .A(n14164), .B(n14163), .ZN(
        n14166) );
  OAI211_X1 U15618 ( .C1(n14169), .C2(n14168), .A(n14167), .B(n14166), .ZN(
        P2_U3212) );
  INV_X2 U15619 ( .A(P2_U3947), .ZN(n14192) );
  MUX2_X1 U15620 ( .A(n14236), .B(P2_DATAO_REG_31__SCAN_IN), .S(n14192), .Z(
        P2_U3562) );
  MUX2_X1 U15621 ( .A(n14170), .B(P2_DATAO_REG_30__SCAN_IN), .S(n14192), .Z(
        P2_U3561) );
  MUX2_X1 U15622 ( .A(n14171), .B(P2_DATAO_REG_29__SCAN_IN), .S(n14192), .Z(
        P2_U3560) );
  MUX2_X1 U15623 ( .A(n14172), .B(P2_DATAO_REG_28__SCAN_IN), .S(n14192), .Z(
        P2_U3559) );
  MUX2_X1 U15624 ( .A(n14173), .B(P2_DATAO_REG_27__SCAN_IN), .S(n14192), .Z(
        P2_U3558) );
  MUX2_X1 U15625 ( .A(n14174), .B(P2_DATAO_REG_26__SCAN_IN), .S(n14192), .Z(
        P2_U3557) );
  MUX2_X1 U15626 ( .A(n14175), .B(P2_DATAO_REG_25__SCAN_IN), .S(n14192), .Z(
        P2_U3556) );
  MUX2_X1 U15627 ( .A(n14176), .B(P2_DATAO_REG_24__SCAN_IN), .S(n14192), .Z(
        P2_U3555) );
  MUX2_X1 U15628 ( .A(n14177), .B(P2_DATAO_REG_23__SCAN_IN), .S(n14192), .Z(
        P2_U3554) );
  MUX2_X1 U15629 ( .A(n14178), .B(P2_DATAO_REG_22__SCAN_IN), .S(n14192), .Z(
        P2_U3553) );
  MUX2_X1 U15630 ( .A(n14179), .B(P2_DATAO_REG_21__SCAN_IN), .S(n14192), .Z(
        P2_U3552) );
  MUX2_X1 U15631 ( .A(n14180), .B(P2_DATAO_REG_20__SCAN_IN), .S(n14192), .Z(
        P2_U3551) );
  MUX2_X1 U15632 ( .A(n14181), .B(P2_DATAO_REG_19__SCAN_IN), .S(n14192), .Z(
        P2_U3550) );
  MUX2_X1 U15633 ( .A(n14182), .B(P2_DATAO_REG_18__SCAN_IN), .S(n14192), .Z(
        P2_U3549) );
  MUX2_X1 U15634 ( .A(n14183), .B(P2_DATAO_REG_17__SCAN_IN), .S(n14192), .Z(
        P2_U3548) );
  MUX2_X1 U15635 ( .A(n14184), .B(P2_DATAO_REG_16__SCAN_IN), .S(n14192), .Z(
        P2_U3547) );
  MUX2_X1 U15636 ( .A(n14185), .B(P2_DATAO_REG_15__SCAN_IN), .S(n14192), .Z(
        P2_U3546) );
  MUX2_X1 U15637 ( .A(n14186), .B(P2_DATAO_REG_14__SCAN_IN), .S(n14192), .Z(
        P2_U3545) );
  MUX2_X1 U15638 ( .A(n14187), .B(P2_DATAO_REG_13__SCAN_IN), .S(n14192), .Z(
        P2_U3544) );
  MUX2_X1 U15639 ( .A(n14188), .B(P2_DATAO_REG_12__SCAN_IN), .S(n14192), .Z(
        P2_U3543) );
  MUX2_X1 U15640 ( .A(n14189), .B(P2_DATAO_REG_11__SCAN_IN), .S(n14192), .Z(
        P2_U3542) );
  MUX2_X1 U15641 ( .A(n14190), .B(P2_DATAO_REG_10__SCAN_IN), .S(n14192), .Z(
        P2_U3541) );
  MUX2_X1 U15642 ( .A(n14191), .B(P2_DATAO_REG_9__SCAN_IN), .S(n14192), .Z(
        P2_U3540) );
  MUX2_X1 U15643 ( .A(n14193), .B(P2_DATAO_REG_8__SCAN_IN), .S(n14192), .Z(
        P2_U3539) );
  MUX2_X1 U15644 ( .A(n14194), .B(P2_DATAO_REG_7__SCAN_IN), .S(n14192), .Z(
        P2_U3538) );
  MUX2_X1 U15645 ( .A(n14195), .B(P2_DATAO_REG_6__SCAN_IN), .S(n14192), .Z(
        P2_U3537) );
  MUX2_X1 U15646 ( .A(n14196), .B(P2_DATAO_REG_5__SCAN_IN), .S(n14192), .Z(
        P2_U3536) );
  MUX2_X1 U15647 ( .A(n14197), .B(P2_DATAO_REG_4__SCAN_IN), .S(n14192), .Z(
        P2_U3535) );
  MUX2_X1 U15648 ( .A(n14198), .B(P2_DATAO_REG_3__SCAN_IN), .S(n14192), .Z(
        P2_U3534) );
  MUX2_X1 U15649 ( .A(n14199), .B(P2_DATAO_REG_2__SCAN_IN), .S(n14192), .Z(
        P2_U3533) );
  MUX2_X1 U15650 ( .A(n14200), .B(P2_DATAO_REG_1__SCAN_IN), .S(n14192), .Z(
        P2_U3532) );
  MUX2_X1 U15651 ( .A(n9773), .B(P2_DATAO_REG_0__SCAN_IN), .S(n14192), .Z(
        P2_U3531) );
  AOI22_X1 U15652 ( .A1(n15471), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n14212) );
  OAI211_X1 U15653 ( .C1(n14203), .C2(n14202), .A(n15473), .B(n14201), .ZN(
        n14211) );
  NAND2_X1 U15654 ( .A1(n14205), .A2(n14204), .ZN(n14210) );
  OAI211_X1 U15655 ( .C1(n14208), .C2(n14207), .A(n15477), .B(n14206), .ZN(
        n14209) );
  NAND4_X1 U15656 ( .A1(n14212), .A2(n14211), .A3(n14210), .A4(n14209), .ZN(
        P2_U3216) );
  AOI22_X1 U15657 ( .A1(n14215), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n14214), 
        .B2(n14213), .ZN(n14217) );
  XNOR2_X1 U15658 ( .A(n7183), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n14216) );
  XNOR2_X1 U15659 ( .A(n14217), .B(n14216), .ZN(n14231) );
  MUX2_X1 U15660 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n14388), .S(n7183), .Z(
        n14222) );
  NOR2_X1 U15661 ( .A1(n14220), .A2(n14219), .ZN(n14221) );
  XOR2_X1 U15662 ( .A(n14222), .B(n14221), .Z(n14228) );
  NAND2_X1 U15663 ( .A1(n15471), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n14225) );
  INV_X1 U15664 ( .A(n14223), .ZN(n14224) );
  OAI211_X1 U15665 ( .C1(n15466), .C2(n14226), .A(n14225), .B(n14224), .ZN(
        n14227) );
  AOI21_X1 U15666 ( .B1(n14228), .B2(n15477), .A(n14227), .ZN(n14229) );
  OAI21_X1 U15667 ( .B1(n14231), .B2(n14230), .A(n14229), .ZN(P2_U3233) );
  NAND2_X1 U15668 ( .A1(n14540), .A2(n14240), .ZN(n14239) );
  XNOR2_X1 U15669 ( .A(n14239), .B(n14233), .ZN(n14234) );
  NOR2_X2 U15670 ( .A1(n14234), .A2(n14416), .ZN(n14445) );
  NAND2_X1 U15671 ( .A1(n14445), .A2(n14438), .ZN(n14238) );
  AND2_X1 U15672 ( .A1(n14236), .A2(n14235), .ZN(n14444) );
  INV_X1 U15673 ( .A(n14444), .ZN(n14448) );
  NOR2_X1 U15674 ( .A1(n14378), .A2(n14448), .ZN(n14242) );
  AOI21_X1 U15675 ( .B1(n14378), .B2(P2_REG2_REG_31__SCAN_IN), .A(n14242), 
        .ZN(n14237) );
  OAI211_X1 U15676 ( .C1(n14536), .C2(n14366), .A(n14238), .B(n14237), .ZN(
        P2_U3234) );
  OAI211_X1 U15677 ( .C1(n14540), .C2(n14240), .A(n14397), .B(n14239), .ZN(
        n14449) );
  NOR2_X1 U15678 ( .A1(n14540), .A2(n14366), .ZN(n14241) );
  AOI211_X1 U15679 ( .C1(n14378), .C2(P2_REG2_REG_30__SCAN_IN), .A(n14242), 
        .B(n14241), .ZN(n14243) );
  OAI21_X1 U15680 ( .B1(n14420), .B2(n14449), .A(n14243), .ZN(P2_U3235) );
  NAND2_X1 U15681 ( .A1(n14244), .A2(n14250), .ZN(n14245) );
  NAND3_X1 U15682 ( .A1(n14246), .A2(n14393), .A3(n14245), .ZN(n14249) );
  INV_X1 U15683 ( .A(n14247), .ZN(n14248) );
  XNOR2_X1 U15684 ( .A(n14251), .B(n14250), .ZN(n14457) );
  NAND2_X1 U15685 ( .A1(n14457), .A2(n14436), .ZN(n14258) );
  NOR2_X1 U15686 ( .A1(n14544), .A2(n14264), .ZN(n14252) );
  AOI22_X1 U15687 ( .A1(n14254), .A2(n14376), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n14378), .ZN(n14255) );
  OAI21_X1 U15688 ( .B1(n14544), .B2(n14366), .A(n14255), .ZN(n14256) );
  AOI21_X1 U15689 ( .B1(n8180), .B2(n14438), .A(n14256), .ZN(n14257) );
  OAI211_X1 U15690 ( .C1(n7242), .C2(n14378), .A(n14258), .B(n14257), .ZN(
        P2_U3237) );
  XNOR2_X1 U15691 ( .A(n14259), .B(n14262), .ZN(n14261) );
  AOI21_X1 U15692 ( .B1(n14261), .B2(n14393), .A(n14260), .ZN(n14461) );
  XNOR2_X1 U15693 ( .A(n14263), .B(n14262), .ZN(n14459) );
  INV_X1 U15694 ( .A(n14264), .ZN(n14266) );
  NAND2_X1 U15695 ( .A1(n14274), .A2(n14463), .ZN(n14265) );
  NAND3_X1 U15696 ( .A1(n14266), .A2(n14397), .A3(n14265), .ZN(n14460) );
  NOR2_X1 U15697 ( .A1(n14460), .A2(n14420), .ZN(n14271) );
  INV_X1 U15698 ( .A(n14267), .ZN(n14268) );
  AOI22_X1 U15699 ( .A1(n14268), .A2(n14376), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n14378), .ZN(n14269) );
  OAI21_X1 U15700 ( .B1(n7375), .B2(n14366), .A(n14269), .ZN(n14270) );
  AOI211_X1 U15701 ( .C1(n14459), .C2(n14436), .A(n14271), .B(n14270), .ZN(
        n14272) );
  OAI21_X1 U15702 ( .B1(n14461), .B2(n14378), .A(n14272), .ZN(P2_U3238) );
  XNOR2_X1 U15703 ( .A(n14273), .B(n14282), .ZN(n14466) );
  INV_X1 U15704 ( .A(n14466), .ZN(n14289) );
  INV_X1 U15705 ( .A(n14300), .ZN(n14276) );
  INV_X1 U15706 ( .A(n14274), .ZN(n14275) );
  AOI211_X1 U15707 ( .C1(n14277), .C2(n14276), .A(n14416), .B(n14275), .ZN(
        n14464) );
  INV_X1 U15708 ( .A(n14278), .ZN(n14279) );
  AOI22_X1 U15709 ( .A1(n14279), .A2(n14376), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14378), .ZN(n14280) );
  OAI21_X1 U15710 ( .B1(n14551), .B2(n14366), .A(n14280), .ZN(n14281) );
  AOI21_X1 U15711 ( .B1(n14464), .B2(n14438), .A(n14281), .ZN(n14288) );
  XNOR2_X1 U15712 ( .A(n14283), .B(n14282), .ZN(n14286) );
  INV_X1 U15713 ( .A(n14284), .ZN(n14285) );
  OAI21_X1 U15714 ( .B1(n14286), .B2(n14413), .A(n14285), .ZN(n14465) );
  NAND2_X1 U15715 ( .A1(n14465), .A2(n14427), .ZN(n14287) );
  OAI211_X1 U15716 ( .C1(n14289), .C2(n14303), .A(n14288), .B(n14287), .ZN(
        P2_U3239) );
  XNOR2_X1 U15717 ( .A(n14290), .B(n14294), .ZN(n14292) );
  AOI21_X1 U15718 ( .B1(n14292), .B2(n14393), .A(n14291), .ZN(n14472) );
  AOI21_X1 U15719 ( .B1(n14294), .B2(n14293), .A(n7251), .ZN(n14473) );
  INV_X1 U15720 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n14295) );
  OAI22_X1 U15721 ( .A1(n14296), .A2(n14430), .B1(n14295), .B2(n14427), .ZN(
        n14297) );
  AOI21_X1 U15722 ( .B1(n14470), .B2(n14434), .A(n14297), .ZN(n14302) );
  NAND2_X1 U15723 ( .A1(n14470), .A2(n7220), .ZN(n14298) );
  NAND2_X1 U15724 ( .A1(n14298), .A2(n14397), .ZN(n14299) );
  NOR2_X1 U15725 ( .A1(n14300), .A2(n14299), .ZN(n14469) );
  NAND2_X1 U15726 ( .A1(n14469), .A2(n14438), .ZN(n14301) );
  OAI211_X1 U15727 ( .C1(n14473), .C2(n14303), .A(n14302), .B(n14301), .ZN(
        n14304) );
  INV_X1 U15728 ( .A(n14304), .ZN(n14305) );
  OAI21_X1 U15729 ( .B1(n14378), .B2(n14472), .A(n14305), .ZN(P2_U3240) );
  XNOR2_X1 U15730 ( .A(n14310), .B(n14306), .ZN(n14308) );
  AOI21_X1 U15731 ( .B1(n14308), .B2(n14393), .A(n14307), .ZN(n14477) );
  OAI21_X1 U15732 ( .B1(n14311), .B2(n14310), .A(n14309), .ZN(n14478) );
  INV_X1 U15733 ( .A(n14478), .ZN(n14317) );
  AOI21_X1 U15734 ( .B1(n14475), .B2(n14326), .A(n14416), .ZN(n14312) );
  AND2_X1 U15735 ( .A1(n14312), .A2(n7220), .ZN(n14474) );
  NAND2_X1 U15736 ( .A1(n14474), .A2(n14438), .ZN(n14315) );
  AOI22_X1 U15737 ( .A1(n14313), .A2(n14376), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n14378), .ZN(n14314) );
  OAI211_X1 U15738 ( .C1(n7691), .C2(n14366), .A(n14315), .B(n14314), .ZN(
        n14316) );
  AOI21_X1 U15739 ( .B1(n14317), .B2(n14436), .A(n14316), .ZN(n14318) );
  OAI21_X1 U15740 ( .B1(n14378), .B2(n14477), .A(n14318), .ZN(P2_U3241) );
  XNOR2_X1 U15741 ( .A(n14319), .B(n14324), .ZN(n14322) );
  INV_X1 U15742 ( .A(n14320), .ZN(n14321) );
  AOI21_X1 U15743 ( .B1(n14322), .B2(n14393), .A(n14321), .ZN(n14482) );
  AOI21_X1 U15744 ( .B1(n14324), .B2(n14323), .A(n7268), .ZN(n14484) );
  INV_X1 U15745 ( .A(n14484), .ZN(n14332) );
  INV_X1 U15746 ( .A(n14480), .ZN(n14330) );
  AOI21_X1 U15747 ( .B1(n14480), .B2(n14344), .A(n14416), .ZN(n14325) );
  AND2_X1 U15748 ( .A1(n14326), .A2(n14325), .ZN(n14479) );
  NAND2_X1 U15749 ( .A1(n14479), .A2(n14438), .ZN(n14329) );
  AOI22_X1 U15750 ( .A1(n14327), .A2(n14376), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n14378), .ZN(n14328) );
  OAI211_X1 U15751 ( .C1(n14330), .C2(n14366), .A(n14329), .B(n14328), .ZN(
        n14331) );
  AOI21_X1 U15752 ( .B1(n14332), .B2(n14436), .A(n14331), .ZN(n14333) );
  OAI21_X1 U15753 ( .B1(n14378), .B2(n14482), .A(n14333), .ZN(P2_U3242) );
  INV_X1 U15754 ( .A(n14334), .ZN(n14335) );
  AOI21_X1 U15755 ( .B1(n14340), .B2(n14336), .A(n14335), .ZN(n14488) );
  NAND2_X1 U15756 ( .A1(n14488), .A2(n14436), .ZN(n14349) );
  INV_X1 U15757 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n14338) );
  OAI22_X1 U15758 ( .A1(n14338), .A2(n14427), .B1(n14337), .B2(n14430), .ZN(
        n14339) );
  AOI21_X1 U15759 ( .B1(n14485), .B2(n14434), .A(n14339), .ZN(n14348) );
  XNOR2_X1 U15760 ( .A(n14341), .B(n14340), .ZN(n14343) );
  OAI21_X1 U15761 ( .B1(n14343), .B2(n14413), .A(n14342), .ZN(n14486) );
  NAND2_X1 U15762 ( .A1(n14486), .A2(n14427), .ZN(n14347) );
  AOI21_X1 U15763 ( .B1(n14485), .B2(n14359), .A(n14416), .ZN(n14345) );
  AND2_X1 U15764 ( .A1(n14345), .A2(n14344), .ZN(n14487) );
  NAND2_X1 U15765 ( .A1(n14487), .A2(n14438), .ZN(n14346) );
  NAND4_X1 U15766 ( .A1(n14349), .A2(n14348), .A3(n14347), .A4(n14346), .ZN(
        P2_U3243) );
  XNOR2_X1 U15767 ( .A(n14351), .B(n14350), .ZN(n14352) );
  OAI222_X1 U15768 ( .A1(n14356), .A2(n14355), .B1(n14354), .B2(n14353), .C1(
        n14352), .C2(n14413), .ZN(n14491) );
  INV_X1 U15769 ( .A(n14491), .ZN(n14369) );
  XNOR2_X1 U15770 ( .A(n14358), .B(n14357), .ZN(n14493) );
  INV_X1 U15771 ( .A(n14359), .ZN(n14360) );
  AOI211_X1 U15772 ( .C1(n14361), .C2(n14375), .A(n14416), .B(n14360), .ZN(
        n14492) );
  NAND2_X1 U15773 ( .A1(n14492), .A2(n14438), .ZN(n14365) );
  INV_X1 U15774 ( .A(n14362), .ZN(n14363) );
  AOI22_X1 U15775 ( .A1(n14378), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n14363), 
        .B2(n14376), .ZN(n14364) );
  OAI211_X1 U15776 ( .C1(n14562), .C2(n14366), .A(n14365), .B(n14364), .ZN(
        n14367) );
  AOI21_X1 U15777 ( .B1(n14436), .B2(n14493), .A(n14367), .ZN(n14368) );
  OAI21_X1 U15778 ( .B1(n14369), .B2(n14378), .A(n14368), .ZN(P2_U3244) );
  XNOR2_X1 U15779 ( .A(n14370), .B(n14373), .ZN(n14372) );
  AOI21_X1 U15780 ( .B1(n14372), .B2(n14393), .A(n14371), .ZN(n14499) );
  XNOR2_X1 U15781 ( .A(n14374), .B(n14373), .ZN(n14497) );
  OAI211_X1 U15782 ( .C1(n14400), .C2(n14567), .A(n14375), .B(n14397), .ZN(
        n14498) );
  AOI22_X1 U15783 ( .A1(n14378), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14377), 
        .B2(n14376), .ZN(n14380) );
  NAND2_X1 U15784 ( .A1(n14502), .A2(n14434), .ZN(n14379) );
  OAI211_X1 U15785 ( .C1(n14498), .C2(n14420), .A(n14380), .B(n14379), .ZN(
        n14381) );
  AOI21_X1 U15786 ( .B1(n14497), .B2(n14436), .A(n14381), .ZN(n14382) );
  OAI21_X1 U15787 ( .B1(n14378), .B2(n14499), .A(n14382), .ZN(P2_U3245) );
  OR2_X1 U15788 ( .A1(n14383), .A2(n14390), .ZN(n14384) );
  NAND2_X1 U15789 ( .A1(n14385), .A2(n14384), .ZN(n14506) );
  NAND2_X1 U15790 ( .A1(n14506), .A2(n14436), .ZN(n14404) );
  INV_X1 U15791 ( .A(n14386), .ZN(n14387) );
  OAI22_X1 U15792 ( .A1(n14427), .A2(n14388), .B1(n14387), .B2(n14430), .ZN(
        n14389) );
  AOI21_X1 U15793 ( .B1(n14570), .B2(n14434), .A(n14389), .ZN(n14403) );
  NAND2_X1 U15794 ( .A1(n14391), .A2(n14390), .ZN(n14392) );
  NAND3_X1 U15795 ( .A1(n14394), .A2(n14393), .A3(n14392), .ZN(n14396) );
  NAND2_X1 U15796 ( .A1(n14396), .A2(n14395), .ZN(n14505) );
  NAND2_X1 U15797 ( .A1(n14505), .A2(n14427), .ZN(n14402) );
  NAND2_X1 U15798 ( .A1(n14418), .A2(n14570), .ZN(n14398) );
  NAND2_X1 U15799 ( .A1(n14398), .A2(n14397), .ZN(n14399) );
  NOR2_X1 U15800 ( .A1(n14400), .A2(n14399), .ZN(n14504) );
  NAND2_X1 U15801 ( .A1(n14504), .A2(n14438), .ZN(n14401) );
  NAND4_X1 U15802 ( .A1(n14404), .A2(n14403), .A3(n14402), .A4(n14401), .ZN(
        P2_U3246) );
  OR2_X1 U15803 ( .A1(n14405), .A2(n14408), .ZN(n14407) );
  NAND2_X1 U15804 ( .A1(n14407), .A2(n14406), .ZN(n14512) );
  INV_X1 U15805 ( .A(n14512), .ZN(n14426) );
  XNOR2_X1 U15806 ( .A(n14409), .B(n7801), .ZN(n14412) );
  NAND2_X1 U15807 ( .A1(n14512), .A2(n15907), .ZN(n14411) );
  OAI211_X1 U15808 ( .C1(n14413), .C2(n14412), .A(n14411), .B(n14410), .ZN(
        n14516) );
  NAND2_X1 U15809 ( .A1(n14516), .A2(n14427), .ZN(n14424) );
  INV_X1 U15810 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n14415) );
  OAI22_X1 U15811 ( .A1(n14427), .A2(n14415), .B1(n14414), .B2(n14430), .ZN(
        n14422) );
  AOI21_X1 U15812 ( .B1(n14417), .B2(n14511), .A(n14416), .ZN(n14419) );
  NAND2_X1 U15813 ( .A1(n14419), .A2(n14418), .ZN(n14513) );
  NOR2_X1 U15814 ( .A1(n14513), .A2(n14420), .ZN(n14421) );
  AOI211_X1 U15815 ( .C1(n14434), .C2(n14511), .A(n14422), .B(n14421), .ZN(
        n14423) );
  OAI211_X1 U15816 ( .C1(n14426), .C2(n14425), .A(n14424), .B(n14423), .ZN(
        P2_U3247) );
  NAND2_X1 U15817 ( .A1(n14428), .A2(n14427), .ZN(n14443) );
  INV_X1 U15818 ( .A(n14429), .ZN(n14431) );
  OAI22_X1 U15819 ( .A1(n14427), .A2(n14432), .B1(n14431), .B2(n14430), .ZN(
        n14433) );
  AOI21_X1 U15820 ( .B1(n14435), .B2(n14434), .A(n14433), .ZN(n14442) );
  NAND2_X1 U15821 ( .A1(n14437), .A2(n14436), .ZN(n14441) );
  NAND2_X1 U15822 ( .A1(n14439), .A2(n14438), .ZN(n14440) );
  NAND4_X1 U15823 ( .A1(n14443), .A2(n14442), .A3(n14441), .A4(n14440), .ZN(
        P2_U3256) );
  INV_X1 U15824 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n14446) );
  NOR2_X1 U15825 ( .A1(n14445), .A2(n14444), .ZN(n14533) );
  MUX2_X1 U15826 ( .A(n14446), .B(n14533), .S(n16142), .Z(n14447) );
  INV_X1 U15827 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n14450) );
  AND2_X1 U15828 ( .A1(n14449), .A2(n14448), .ZN(n14537) );
  MUX2_X1 U15829 ( .A(n14450), .B(n14537), .S(n16142), .Z(n14451) );
  OAI21_X1 U15830 ( .B1(n14540), .B2(n14496), .A(n14451), .ZN(P2_U3529) );
  AOI21_X1 U15831 ( .B1(n15905), .B2(n14453), .A(n14452), .ZN(n14454) );
  OAI211_X1 U15832 ( .C1(n14483), .C2(n14456), .A(n14455), .B(n14454), .ZN(
        n14541) );
  MUX2_X1 U15833 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n14541), .S(n16142), .Z(
        P2_U3528) );
  OAI21_X1 U15834 ( .B1(n14544), .B2(n14496), .A(n14458), .ZN(P2_U3527) );
  NAND2_X1 U15835 ( .A1(n14459), .A2(n16140), .ZN(n14462) );
  INV_X1 U15836 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n14467) );
  AOI211_X1 U15837 ( .C1(n14466), .C2(n16140), .A(n14465), .B(n14464), .ZN(
        n14548) );
  MUX2_X1 U15838 ( .A(n14467), .B(n14548), .S(n16142), .Z(n14468) );
  OAI21_X1 U15839 ( .B1(n14551), .B2(n14496), .A(n14468), .ZN(P2_U3525) );
  AOI21_X1 U15840 ( .B1(n15905), .B2(n14470), .A(n14469), .ZN(n14471) );
  OAI211_X1 U15841 ( .C1(n14473), .C2(n14483), .A(n14472), .B(n14471), .ZN(
        n14552) );
  MUX2_X1 U15842 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14552), .S(n16142), .Z(
        P2_U3524) );
  AOI21_X1 U15843 ( .B1(n15905), .B2(n14475), .A(n14474), .ZN(n14476) );
  OAI211_X1 U15844 ( .C1(n14478), .C2(n14483), .A(n14477), .B(n14476), .ZN(
        n14553) );
  MUX2_X1 U15845 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14553), .S(n16142), .Z(
        P2_U3523) );
  AOI21_X1 U15846 ( .B1(n15905), .B2(n14480), .A(n14479), .ZN(n14481) );
  OAI211_X1 U15847 ( .C1(n14484), .C2(n14483), .A(n14482), .B(n14481), .ZN(
        n14554) );
  MUX2_X1 U15848 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14554), .S(n16142), .Z(
        P2_U3522) );
  INV_X1 U15849 ( .A(n14485), .ZN(n14558) );
  INV_X1 U15850 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n14489) );
  AOI211_X1 U15851 ( .C1(n14488), .C2(n16140), .A(n14487), .B(n14486), .ZN(
        n14555) );
  MUX2_X1 U15852 ( .A(n14489), .B(n14555), .S(n16142), .Z(n14490) );
  OAI21_X1 U15853 ( .B1(n14558), .B2(n14496), .A(n14490), .ZN(P2_U3521) );
  INV_X1 U15854 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n14494) );
  AOI211_X1 U15855 ( .C1(n14493), .C2(n16140), .A(n14492), .B(n14491), .ZN(
        n14559) );
  MUX2_X1 U15856 ( .A(n14494), .B(n14559), .S(n16142), .Z(n14495) );
  OAI21_X1 U15857 ( .B1(n14562), .B2(n14496), .A(n14495), .ZN(P2_U3520) );
  NAND2_X1 U15858 ( .A1(n14497), .A2(n16140), .ZN(n14500) );
  NAND3_X1 U15859 ( .A1(n14500), .A2(n14499), .A3(n14498), .ZN(n14563) );
  MUX2_X1 U15860 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14563), .S(n16142), .Z(
        n14501) );
  AOI21_X1 U15861 ( .B1(n14524), .B2(n14502), .A(n14501), .ZN(n14503) );
  INV_X1 U15862 ( .A(n14503), .ZN(P2_U3519) );
  NOR2_X1 U15863 ( .A1(n14505), .A2(n14504), .ZN(n14508) );
  NAND2_X1 U15864 ( .A1(n14506), .A2(n16140), .ZN(n14507) );
  NAND2_X1 U15865 ( .A1(n14508), .A2(n14507), .ZN(n14568) );
  MUX2_X1 U15866 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n14568), .S(n16142), .Z(
        n14509) );
  AOI21_X1 U15867 ( .B1(n14524), .B2(n14570), .A(n14509), .ZN(n14510) );
  INV_X1 U15868 ( .A(n14510), .ZN(P2_U3518) );
  NAND2_X1 U15869 ( .A1(n14512), .A2(n16092), .ZN(n14514) );
  OAI211_X1 U15870 ( .C1(n7683), .C2(n16136), .A(n14514), .B(n14513), .ZN(
        n14515) );
  NOR2_X1 U15871 ( .A1(n14516), .A2(n14515), .ZN(n14572) );
  INV_X1 U15872 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n14517) );
  MUX2_X1 U15873 ( .A(n14572), .B(n14517), .S(n16141), .Z(n14518) );
  INV_X1 U15874 ( .A(n14518), .ZN(P2_U3517) );
  NAND2_X1 U15875 ( .A1(n14519), .A2(n16140), .ZN(n14522) );
  NAND3_X1 U15876 ( .A1(n14522), .A2(n14521), .A3(n14520), .ZN(n14575) );
  MUX2_X1 U15877 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n14575), .S(n16142), .Z(
        n14523) );
  AOI21_X1 U15878 ( .B1(n14524), .B2(n14577), .A(n14523), .ZN(n14525) );
  INV_X1 U15879 ( .A(n14525), .ZN(P2_U3516) );
  NAND2_X1 U15880 ( .A1(n14526), .A2(n15905), .ZN(n14527) );
  NAND2_X1 U15881 ( .A1(n14528), .A2(n14527), .ZN(n14529) );
  AOI21_X1 U15882 ( .B1(n14530), .B2(n16092), .A(n14529), .ZN(n14531) );
  NAND2_X1 U15883 ( .A1(n14532), .A2(n14531), .ZN(n14580) );
  MUX2_X1 U15884 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14580), .S(n16142), .Z(
        P2_U3515) );
  MUX2_X1 U15885 ( .A(n14534), .B(n14533), .S(n16146), .Z(n14535) );
  MUX2_X1 U15886 ( .A(n14538), .B(n14537), .S(n16146), .Z(n14539) );
  OAI21_X1 U15887 ( .B1(n14540), .B2(n14566), .A(n14539), .ZN(P2_U3497) );
  MUX2_X1 U15888 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n14541), .S(n16146), .Z(
        P2_U3496) );
  MUX2_X1 U15889 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14545), .S(n16146), .Z(
        n14546) );
  INV_X1 U15890 ( .A(n14546), .ZN(n14547) );
  OAI21_X1 U15891 ( .B1(n7375), .B2(n14566), .A(n14547), .ZN(P2_U3494) );
  MUX2_X1 U15892 ( .A(n14549), .B(n14548), .S(n16146), .Z(n14550) );
  OAI21_X1 U15893 ( .B1(n14551), .B2(n14566), .A(n14550), .ZN(P2_U3493) );
  MUX2_X1 U15894 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14552), .S(n16146), .Z(
        P2_U3492) );
  MUX2_X1 U15895 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14553), .S(n16146), .Z(
        P2_U3491) );
  MUX2_X1 U15896 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14554), .S(n16146), .Z(
        P2_U3490) );
  MUX2_X1 U15897 ( .A(n14556), .B(n14555), .S(n16146), .Z(n14557) );
  OAI21_X1 U15898 ( .B1(n14558), .B2(n14566), .A(n14557), .ZN(P2_U3489) );
  MUX2_X1 U15899 ( .A(n14560), .B(n14559), .S(n16146), .Z(n14561) );
  OAI21_X1 U15900 ( .B1(n14562), .B2(n14566), .A(n14561), .ZN(P2_U3488) );
  MUX2_X1 U15901 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14563), .S(n16146), .Z(
        n14564) );
  INV_X1 U15902 ( .A(n14564), .ZN(n14565) );
  OAI21_X1 U15903 ( .B1(n14567), .B2(n14566), .A(n14565), .ZN(P2_U3487) );
  MUX2_X1 U15904 ( .A(n14568), .B(P2_REG0_REG_19__SCAN_IN), .S(n16143), .Z(
        n14569) );
  AOI21_X1 U15905 ( .B1(n14578), .B2(n14570), .A(n14569), .ZN(n14571) );
  INV_X1 U15906 ( .A(n14571), .ZN(P2_U3486) );
  MUX2_X1 U15907 ( .A(n14573), .B(n14572), .S(n16146), .Z(n14574) );
  INV_X1 U15908 ( .A(n14574), .ZN(P2_U3484) );
  MUX2_X1 U15909 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n14575), .S(n16146), .Z(
        n14576) );
  AOI21_X1 U15910 ( .B1(n14578), .B2(n14577), .A(n14576), .ZN(n14579) );
  INV_X1 U15911 ( .A(n14579), .ZN(P2_U3481) );
  MUX2_X1 U15912 ( .A(n14580), .B(P2_REG0_REG_16__SCAN_IN), .S(n16143), .Z(
        P2_U3478) );
  INV_X1 U15913 ( .A(n14581), .ZN(n15147) );
  NOR4_X1 U15914 ( .A1(n14583), .A2(P2_IR_REG_30__SCAN_IN), .A3(n14582), .A4(
        P2_U3088), .ZN(n14584) );
  AOI21_X1 U15915 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n14591), .A(n14584), 
        .ZN(n14585) );
  OAI21_X1 U15916 ( .B1(n15147), .B2(n14593), .A(n14585), .ZN(P2_U3296) );
  INV_X1 U15917 ( .A(n14586), .ZN(n15150) );
  OAI222_X1 U15918 ( .A1(n14588), .A2(n14587), .B1(n14593), .B2(n15150), .C1(
        n9578), .C2(P2_U3088), .ZN(P2_U3298) );
  INV_X1 U15919 ( .A(n14589), .ZN(n15152) );
  AOI21_X1 U15920 ( .B1(n14591), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n14590), 
        .ZN(n14592) );
  OAI21_X1 U15921 ( .B1(n15152), .B2(n14593), .A(n14592), .ZN(P2_U3299) );
  INV_X1 U15922 ( .A(n14594), .ZN(n15160) );
  OAI222_X1 U15923 ( .A1(P2_U3088), .A2(n14596), .B1(n14593), .B2(n15160), 
        .C1(n14595), .C2(n14588), .ZN(P2_U3301) );
  INV_X1 U15924 ( .A(n14598), .ZN(n15162) );
  OAI222_X1 U15925 ( .A1(n14588), .A2(n14600), .B1(n14593), .B2(n15162), .C1(
        n14599), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U15926 ( .A(n14601), .ZN(n15168) );
  OAI222_X1 U15927 ( .A1(n14588), .A2(n14603), .B1(n14593), .B2(n15168), .C1(
        P2_U3088), .C2(n14602), .ZN(P2_U3303) );
  INV_X1 U15928 ( .A(n14604), .ZN(n14605) );
  MUX2_X1 U15929 ( .A(n14605), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  AOI22_X1 U15930 ( .A1(n14870), .A2(n14728), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14608) );
  NAND2_X1 U15931 ( .A1(n14899), .A2(n14713), .ZN(n14607) );
  OAI211_X1 U15932 ( .C1(n14609), .C2(n16115), .A(n14608), .B(n14607), .ZN(
        n14610) );
  AOI21_X1 U15933 ( .B1(n14871), .B2(n16129), .A(n14610), .ZN(n14611) );
  OAI21_X1 U15934 ( .B1(n14612), .B2(n16123), .A(n14611), .ZN(P1_U3214) );
  XOR2_X1 U15935 ( .A(n14614), .B(n14613), .Z(n14620) );
  AND2_X1 U15936 ( .A1(n14961), .A2(n14978), .ZN(n14615) );
  AOI21_X1 U15937 ( .B1(n14900), .B2(n14980), .A(n14615), .ZN(n14931) );
  INV_X1 U15938 ( .A(n14616), .ZN(n14936) );
  AOI22_X1 U15939 ( .A1(n14936), .A2(n14728), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14617) );
  OAI21_X1 U15940 ( .B1(n14931), .B2(n14725), .A(n14617), .ZN(n14618) );
  AOI21_X1 U15941 ( .B1(n15069), .B2(n16129), .A(n14618), .ZN(n14619) );
  OAI21_X1 U15942 ( .B1(n14620), .B2(n16123), .A(n14619), .ZN(P1_U3216) );
  OAI21_X1 U15943 ( .B1(n14622), .B2(n14621), .A(n14680), .ZN(n14623) );
  NAND2_X1 U15944 ( .A1(n14623), .A2(n14719), .ZN(n14629) );
  OR2_X1 U15945 ( .A1(n14637), .A2(n15005), .ZN(n14625) );
  NAND2_X1 U15946 ( .A1(n14735), .A2(n14978), .ZN(n14624) );
  NAND2_X1 U15947 ( .A1(n14625), .A2(n14624), .ZN(n15094) );
  NOR2_X1 U15948 ( .A1(n14626), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14839) );
  NOR2_X1 U15949 ( .A1(n16133), .A2(n14993), .ZN(n14627) );
  AOI211_X1 U15950 ( .C1(n15094), .C2(n15927), .A(n14839), .B(n14627), .ZN(
        n14628) );
  OAI211_X1 U15951 ( .C1(n15097), .C2(n14731), .A(n14629), .B(n14628), .ZN(
        P1_U3219) );
  INV_X1 U15952 ( .A(n14630), .ZN(n14634) );
  AOI21_X1 U15953 ( .B1(n14681), .B2(n14632), .A(n14631), .ZN(n14633) );
  OAI21_X1 U15954 ( .B1(n14634), .B2(n14633), .A(n14719), .ZN(n14640) );
  INV_X1 U15955 ( .A(n14635), .ZN(n14963) );
  INV_X1 U15956 ( .A(n14713), .ZN(n16118) );
  INV_X1 U15957 ( .A(n16115), .ZN(n14684) );
  AOI22_X1 U15958 ( .A1(n14961), .A2(n14684), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14636) );
  OAI21_X1 U15959 ( .B1(n14637), .B2(n16118), .A(n14636), .ZN(n14638) );
  AOI21_X1 U15960 ( .B1(n14963), .B2(n14728), .A(n14638), .ZN(n14639) );
  OAI211_X1 U15961 ( .C1(n7609), .C2(n14731), .A(n14640), .B(n14639), .ZN(
        P1_U3223) );
  XOR2_X1 U15962 ( .A(n14642), .B(n14641), .Z(n14647) );
  AOI22_X1 U15963 ( .A1(n14903), .A2(n14728), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14644) );
  NAND2_X1 U15964 ( .A1(n14900), .A2(n14713), .ZN(n14643) );
  OAI211_X1 U15965 ( .C1(n14859), .C2(n16115), .A(n14644), .B(n14643), .ZN(
        n14645) );
  AOI21_X1 U15966 ( .B1(n15057), .B2(n16129), .A(n14645), .ZN(n14646) );
  OAI21_X1 U15967 ( .B1(n14647), .B2(n16123), .A(n14646), .ZN(P1_U3225) );
  INV_X1 U15968 ( .A(n14648), .ZN(n14649) );
  AOI21_X1 U15969 ( .B1(n14651), .B2(n14650), .A(n14649), .ZN(n14658) );
  NOR2_X1 U15970 ( .A1(n16133), .A2(n14652), .ZN(n14655) );
  OAI21_X1 U15971 ( .B1(n14725), .B2(n15114), .A(n14653), .ZN(n14654) );
  AOI211_X1 U15972 ( .C1(n14656), .C2(n16129), .A(n14655), .B(n14654), .ZN(
        n14657) );
  OAI21_X1 U15973 ( .B1(n14658), .B2(n16123), .A(n14657), .ZN(P1_U3226) );
  XNOR2_X1 U15974 ( .A(n14660), .B(n14659), .ZN(n14661) );
  XNOR2_X1 U15975 ( .A(n14662), .B(n14661), .ZN(n14671) );
  OAI21_X1 U15976 ( .B1(n16118), .B2(n14664), .A(n14663), .ZN(n14665) );
  AOI21_X1 U15977 ( .B1(n14684), .B2(n14735), .A(n14665), .ZN(n14666) );
  OAI21_X1 U15978 ( .B1(n14667), .B2(n16133), .A(n14666), .ZN(n14668) );
  AOI21_X1 U15979 ( .B1(n14669), .B2(n16129), .A(n14668), .ZN(n14670) );
  OAI21_X1 U15980 ( .B1(n14671), .B2(n16123), .A(n14670), .ZN(P1_U3228) );
  XOR2_X1 U15981 ( .A(n14673), .B(n14672), .Z(n14678) );
  AOI22_X1 U15982 ( .A1(n14951), .A2(n14713), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14675) );
  NAND2_X1 U15983 ( .A1(n14923), .A2(n14728), .ZN(n14674) );
  OAI211_X1 U15984 ( .C1(n14914), .C2(n16115), .A(n14675), .B(n14674), .ZN(
        n14676) );
  AOI21_X1 U15985 ( .B1(n15064), .B2(n16129), .A(n14676), .ZN(n14677) );
  OAI21_X1 U15986 ( .B1(n14678), .B2(n16123), .A(n14677), .ZN(P1_U3229) );
  AND2_X1 U15987 ( .A1(n14680), .A2(n14679), .ZN(n14683) );
  OAI211_X1 U15988 ( .C1(n14683), .C2(n14682), .A(n14719), .B(n14681), .ZN(
        n14688) );
  AOI22_X1 U15989 ( .A1(n14981), .A2(n14684), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14685) );
  OAI21_X1 U15990 ( .B1(n15006), .B2(n16118), .A(n14685), .ZN(n14686) );
  AOI21_X1 U15991 ( .B1(n14982), .B2(n14728), .A(n14686), .ZN(n14687) );
  OAI211_X1 U15992 ( .C1(n14976), .C2(n14731), .A(n14688), .B(n14687), .ZN(
        P1_U3233) );
  INV_X1 U15993 ( .A(n14692), .ZN(n14689) );
  NOR2_X1 U15994 ( .A1(n14690), .A2(n14689), .ZN(n14695) );
  AOI21_X1 U15995 ( .B1(n14693), .B2(n14692), .A(n14691), .ZN(n14694) );
  OAI21_X1 U15996 ( .B1(n14695), .B2(n14694), .A(n14719), .ZN(n14699) );
  AOI22_X1 U15997 ( .A1(n14981), .A2(n14713), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14696) );
  OAI21_X1 U15998 ( .B1(n14913), .B2(n16115), .A(n14696), .ZN(n14697) );
  AOI21_X1 U15999 ( .B1(n14954), .B2(n14728), .A(n14697), .ZN(n14698) );
  OAI211_X1 U16000 ( .C1(n14731), .C2(n15075), .A(n14699), .B(n14698), .ZN(
        P1_U3235) );
  INV_X1 U16001 ( .A(n14700), .ZN(n14701) );
  AOI21_X1 U16002 ( .B1(n14703), .B2(n14702), .A(n14701), .ZN(n14709) );
  OAI21_X1 U16003 ( .B1(n16115), .B2(n15006), .A(n14704), .ZN(n14705) );
  AOI21_X1 U16004 ( .B1(n14713), .B2(n14736), .A(n14705), .ZN(n14706) );
  OAI21_X1 U16005 ( .B1(n15017), .B2(n16133), .A(n14706), .ZN(n14707) );
  AOI21_X1 U16006 ( .B1(n15104), .B2(n16129), .A(n14707), .ZN(n14708) );
  OAI21_X1 U16007 ( .B1(n14709), .B2(n16123), .A(n14708), .ZN(P1_U3238) );
  XOR2_X1 U16008 ( .A(n14711), .B(n14710), .Z(n14718) );
  INV_X1 U16009 ( .A(n14712), .ZN(n14887) );
  AOI22_X1 U16010 ( .A1(n14887), .A2(n14728), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14715) );
  NAND2_X1 U16011 ( .A1(n14881), .A2(n14713), .ZN(n14714) );
  OAI211_X1 U16012 ( .C1(n7998), .C2(n16115), .A(n14715), .B(n14714), .ZN(
        n14716) );
  AOI21_X1 U16013 ( .B1(n15051), .B2(n16129), .A(n14716), .ZN(n14717) );
  OAI21_X1 U16014 ( .B1(n14718), .B2(n16123), .A(n14717), .ZN(P1_U3240) );
  OAI211_X1 U16015 ( .C1(n14722), .C2(n14721), .A(n14720), .B(n14719), .ZN(
        n14730) );
  OAI22_X1 U16016 ( .A1(n14725), .A2(n14724), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14723), .ZN(n14726) );
  AOI21_X1 U16017 ( .B1(n14728), .B2(n14727), .A(n14726), .ZN(n14729) );
  OAI211_X1 U16018 ( .C1(n14732), .C2(n14731), .A(n14730), .B(n14729), .ZN(
        P1_U3241) );
  MUX2_X1 U16019 ( .A(n14845), .B(P1_DATAO_REG_31__SCAN_IN), .S(n14752), .Z(
        P1_U3591) );
  MUX2_X1 U16020 ( .A(n14733), .B(P1_DATAO_REG_30__SCAN_IN), .S(n14752), .Z(
        P1_U3590) );
  MUX2_X1 U16021 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14734), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16022 ( .A(n14857), .B(P1_DATAO_REG_28__SCAN_IN), .S(n14752), .Z(
        P1_U3588) );
  MUX2_X1 U16023 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14882), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16024 ( .A(n14899), .B(P1_DATAO_REG_26__SCAN_IN), .S(n14752), .Z(
        P1_U3586) );
  MUX2_X1 U16025 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14881), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16026 ( .A(n14900), .B(P1_DATAO_REG_24__SCAN_IN), .S(n14752), .Z(
        P1_U3584) );
  MUX2_X1 U16027 ( .A(n14951), .B(P1_DATAO_REG_23__SCAN_IN), .S(n14752), .Z(
        P1_U3583) );
  MUX2_X1 U16028 ( .A(n14961), .B(P1_DATAO_REG_22__SCAN_IN), .S(n14752), .Z(
        P1_U3582) );
  MUX2_X1 U16029 ( .A(n14981), .B(P1_DATAO_REG_21__SCAN_IN), .S(n14752), .Z(
        P1_U3581) );
  MUX2_X1 U16030 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14962), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16031 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14979), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16032 ( .A(n14735), .B(P1_DATAO_REG_18__SCAN_IN), .S(n14752), .Z(
        P1_U3578) );
  MUX2_X1 U16033 ( .A(n14736), .B(P1_DATAO_REG_17__SCAN_IN), .S(n14752), .Z(
        P1_U3577) );
  MUX2_X1 U16034 ( .A(n14737), .B(P1_DATAO_REG_16__SCAN_IN), .S(n14752), .Z(
        P1_U3576) );
  MUX2_X1 U16035 ( .A(n14738), .B(P1_DATAO_REG_15__SCAN_IN), .S(n14752), .Z(
        P1_U3575) );
  MUX2_X1 U16036 ( .A(n14739), .B(P1_DATAO_REG_14__SCAN_IN), .S(n14752), .Z(
        P1_U3574) );
  MUX2_X1 U16037 ( .A(n14740), .B(P1_DATAO_REG_13__SCAN_IN), .S(n14752), .Z(
        P1_U3573) );
  MUX2_X1 U16038 ( .A(n14741), .B(P1_DATAO_REG_12__SCAN_IN), .S(n14752), .Z(
        P1_U3572) );
  MUX2_X1 U16039 ( .A(n14742), .B(P1_DATAO_REG_11__SCAN_IN), .S(n14752), .Z(
        P1_U3571) );
  MUX2_X1 U16040 ( .A(n14743), .B(P1_DATAO_REG_10__SCAN_IN), .S(n14752), .Z(
        P1_U3570) );
  MUX2_X1 U16041 ( .A(n14744), .B(P1_DATAO_REG_9__SCAN_IN), .S(n14752), .Z(
        P1_U3569) );
  MUX2_X1 U16042 ( .A(n14745), .B(P1_DATAO_REG_8__SCAN_IN), .S(n14752), .Z(
        P1_U3568) );
  MUX2_X1 U16043 ( .A(n14746), .B(P1_DATAO_REG_7__SCAN_IN), .S(n14752), .Z(
        P1_U3567) );
  MUX2_X1 U16044 ( .A(n14747), .B(P1_DATAO_REG_6__SCAN_IN), .S(n14752), .Z(
        P1_U3566) );
  MUX2_X1 U16045 ( .A(n14748), .B(P1_DATAO_REG_5__SCAN_IN), .S(n14752), .Z(
        P1_U3565) );
  MUX2_X1 U16046 ( .A(n14749), .B(P1_DATAO_REG_4__SCAN_IN), .S(n14752), .Z(
        P1_U3564) );
  MUX2_X1 U16047 ( .A(n14750), .B(P1_DATAO_REG_3__SCAN_IN), .S(n14752), .Z(
        P1_U3563) );
  MUX2_X1 U16048 ( .A(n14751), .B(P1_DATAO_REG_2__SCAN_IN), .S(n14752), .Z(
        P1_U3562) );
  MUX2_X1 U16049 ( .A(n14753), .B(P1_DATAO_REG_1__SCAN_IN), .S(n14752), .Z(
        P1_U3561) );
  MUX2_X1 U16050 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14754), .S(P1_U4016), .Z(
        P1_U3560) );
  AOI22_X1 U16051 ( .A1(n14797), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14766) );
  OAI211_X1 U16052 ( .C1(n14756), .C2(n14768), .A(n14833), .B(n14755), .ZN(
        n14765) );
  NAND2_X1 U16053 ( .A1(n14787), .A2(n14757), .ZN(n14764) );
  MUX2_X1 U16054 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n15859), .S(n14758), .Z(
        n14759) );
  OAI21_X1 U16055 ( .B1(n15836), .B2(n14760), .A(n14759), .ZN(n14761) );
  NAND3_X1 U16056 ( .A1(n14834), .A2(n14762), .A3(n14761), .ZN(n14763) );
  NAND4_X1 U16057 ( .A1(n14766), .A2(n14765), .A3(n14764), .A4(n14763), .ZN(
        P1_U3244) );
  MUX2_X1 U16058 ( .A(n14768), .B(n14767), .S(n15154), .Z(n14770) );
  NAND2_X1 U16059 ( .A1(n14770), .A2(n14769), .ZN(n14771) );
  OAI211_X1 U16060 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n14772), .A(n14771), .B(
        P1_U4016), .ZN(n14818) );
  AOI22_X1 U16061 ( .A1(n14797), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n14784) );
  OAI211_X1 U16062 ( .C1(n14774), .C2(n14773), .A(n14833), .B(n14790), .ZN(
        n14780) );
  INV_X1 U16063 ( .A(n14775), .ZN(n14777) );
  XNOR2_X1 U16064 ( .A(n14777), .B(n14776), .ZN(n14778) );
  NAND2_X1 U16065 ( .A1(n14834), .A2(n14778), .ZN(n14779) );
  AND2_X1 U16066 ( .A1(n14780), .A2(n14779), .ZN(n14783) );
  OR2_X1 U16067 ( .A1(n14828), .A2(n14781), .ZN(n14782) );
  NAND4_X1 U16068 ( .A1(n14818), .A2(n14784), .A3(n14783), .A4(n14782), .ZN(
        P1_U3245) );
  OAI211_X1 U16069 ( .C1(n14786), .C2(n14785), .A(n14834), .B(n14805), .ZN(
        n14796) );
  NAND2_X1 U16070 ( .A1(n14787), .A2(n14788), .ZN(n14795) );
  MUX2_X1 U16071 ( .A(n10627), .B(P1_REG2_REG_3__SCAN_IN), .S(n14788), .Z(
        n14791) );
  NAND3_X1 U16072 ( .A1(n14791), .A2(n14790), .A3(n14789), .ZN(n14792) );
  NAND3_X1 U16073 ( .A1(n14833), .A2(n14812), .A3(n14792), .ZN(n14794) );
  AND2_X1 U16074 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n15919) );
  AOI21_X1 U16075 ( .B1(n14797), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n15919), .ZN(
        n14793) );
  NAND4_X1 U16076 ( .A1(n14796), .A2(n14795), .A3(n14794), .A4(n14793), .ZN(
        P1_U3246) );
  NAND2_X1 U16077 ( .A1(n14797), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n14799) );
  OAI211_X1 U16078 ( .C1(n14828), .C2(n14800), .A(n14799), .B(n14798), .ZN(
        n14801) );
  INV_X1 U16079 ( .A(n14801), .ZN(n14817) );
  INV_X1 U16080 ( .A(n14802), .ZN(n14807) );
  NAND3_X1 U16081 ( .A1(n14805), .A2(n14804), .A3(n14803), .ZN(n14806) );
  NAND3_X1 U16082 ( .A1(n14834), .A2(n14807), .A3(n14806), .ZN(n14816) );
  MUX2_X1 U16083 ( .A(n14809), .B(P1_REG2_REG_4__SCAN_IN), .S(n14808), .Z(
        n14810) );
  NAND3_X1 U16084 ( .A1(n14812), .A2(n14811), .A3(n14810), .ZN(n14813) );
  NAND3_X1 U16085 ( .A1(n14833), .A2(n14814), .A3(n14813), .ZN(n14815) );
  NAND4_X1 U16086 ( .A1(n14818), .A2(n14817), .A3(n14816), .A4(n14815), .ZN(
        P1_U3247) );
  NAND2_X1 U16087 ( .A1(n14824), .A2(n14819), .ZN(n14820) );
  NAND2_X1 U16088 ( .A1(n14821), .A2(n14820), .ZN(n14822) );
  XOR2_X1 U16089 ( .A(n14822), .B(P1_REG1_REG_19__SCAN_IN), .Z(n14835) );
  INV_X1 U16090 ( .A(n14835), .ZN(n14831) );
  NAND2_X1 U16091 ( .A1(n14824), .A2(n14823), .ZN(n14825) );
  NAND2_X1 U16092 ( .A1(n14826), .A2(n14825), .ZN(n14827) );
  XOR2_X1 U16093 ( .A(n14827), .B(P1_REG2_REG_19__SCAN_IN), .Z(n14832) );
  OAI21_X1 U16094 ( .B1(n14832), .B2(n14829), .A(n14828), .ZN(n14830) );
  AOI21_X1 U16095 ( .B1(n14831), .B2(n14834), .A(n14830), .ZN(n14838) );
  AOI22_X1 U16096 ( .A1(n14835), .A2(n14834), .B1(n14833), .B2(n14832), .ZN(
        n14837) );
  MUX2_X1 U16097 ( .A(n14838), .B(n14837), .S(n14836), .Z(n14841) );
  INV_X1 U16098 ( .A(n14839), .ZN(n14840) );
  OAI211_X1 U16099 ( .C1(n14842), .C2(n7623), .A(n14841), .B(n14840), .ZN(
        P1_U3262) );
  INV_X1 U16100 ( .A(n14843), .ZN(n15840) );
  AND2_X1 U16101 ( .A1(n14845), .A2(n14844), .ZN(n15027) );
  INV_X1 U16102 ( .A(n15027), .ZN(n14846) );
  NOR2_X1 U16103 ( .A1(n16047), .A2(n14846), .ZN(n14853) );
  AOI21_X1 U16104 ( .B1(n16047), .B2(P1_REG2_REG_31__SCAN_IN), .A(n14853), 
        .ZN(n14848) );
  NAND2_X1 U16105 ( .A1(n15024), .A2(n15990), .ZN(n14847) );
  OAI211_X1 U16106 ( .C1(n15023), .C2(n15840), .A(n14848), .B(n14847), .ZN(
        P1_U3263) );
  OAI21_X1 U16107 ( .B1(n14850), .B2(n14851), .A(n14849), .ZN(n15030) );
  NOR2_X1 U16108 ( .A1(n14851), .A2(n16041), .ZN(n14852) );
  AOI211_X1 U16109 ( .C1(n16047), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14853), 
        .B(n14852), .ZN(n14854) );
  OAI21_X1 U16110 ( .B1(n15840), .B2(n15030), .A(n14854), .ZN(P1_U3264) );
  OAI21_X1 U16111 ( .B1(n14856), .B2(n14862), .A(n14855), .ZN(n14861) );
  NAND2_X1 U16112 ( .A1(n14857), .A2(n14980), .ZN(n14858) );
  OAI21_X1 U16113 ( .B1(n14859), .B2(n15003), .A(n14858), .ZN(n14860) );
  NAND2_X1 U16114 ( .A1(n14863), .A2(n14862), .ZN(n14864) );
  NAND2_X1 U16115 ( .A1(n14865), .A2(n14864), .ZN(n15046) );
  NAND2_X1 U16116 ( .A1(n15046), .A2(n16034), .ZN(n14866) );
  NAND2_X1 U16117 ( .A1(n14871), .A2(n14885), .ZN(n14867) );
  NAND2_X1 U16118 ( .A1(n14867), .A2(n15041), .ZN(n14868) );
  OR2_X1 U16119 ( .A1(n7185), .A2(n14868), .ZN(n15047) );
  AOI22_X1 U16120 ( .A1(n14870), .A2(n16037), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n15998), .ZN(n14873) );
  NAND2_X1 U16121 ( .A1(n14871), .A2(n15990), .ZN(n14872) );
  OAI211_X1 U16122 ( .C1(n15047), .C2(n14997), .A(n14873), .B(n14872), .ZN(
        n14874) );
  AOI21_X1 U16123 ( .B1(n15046), .B2(n16044), .A(n14874), .ZN(n14875) );
  OAI21_X1 U16124 ( .B1(n7293), .B2(n15998), .A(n14875), .ZN(P1_U3266) );
  XNOR2_X1 U16125 ( .A(n14876), .B(n14877), .ZN(n15054) );
  OAI21_X1 U16126 ( .B1(n14880), .B2(n14879), .A(n14878), .ZN(n14883) );
  AOI222_X1 U16127 ( .A1(n15955), .A2(n14883), .B1(n14882), .B2(n14980), .C1(
        n14881), .C2(n14978), .ZN(n15053) );
  INV_X1 U16128 ( .A(n15053), .ZN(n14891) );
  AOI21_X1 U16129 ( .B1(n15051), .B2(n14897), .A(n15952), .ZN(n14886) );
  AND2_X1 U16130 ( .A1(n14886), .A2(n14885), .ZN(n15050) );
  NAND2_X1 U16131 ( .A1(n15050), .A2(n16035), .ZN(n14889) );
  AOI22_X1 U16132 ( .A1(n14887), .A2(n16037), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n15998), .ZN(n14888) );
  OAI211_X1 U16133 ( .C1(n12164), .C2(n16041), .A(n14889), .B(n14888), .ZN(
        n14890) );
  AOI21_X1 U16134 ( .B1(n14891), .B2(n11899), .A(n14890), .ZN(n14892) );
  OAI21_X1 U16135 ( .B1(n14967), .B2(n15054), .A(n14892), .ZN(P1_U3267) );
  OAI21_X1 U16136 ( .B1(n7294), .B2(n14894), .A(n14893), .ZN(n15061) );
  OAI21_X1 U16137 ( .B1(n14896), .B2(n12103), .A(n14895), .ZN(n15058) );
  AOI21_X1 U16138 ( .B1(n15057), .B2(n14921), .A(n15952), .ZN(n14898) );
  AND2_X1 U16139 ( .A1(n14898), .A2(n14897), .ZN(n15055) );
  NAND2_X1 U16140 ( .A1(n15055), .A2(n16035), .ZN(n14908) );
  NAND2_X1 U16141 ( .A1(n15057), .A2(n15990), .ZN(n14907) );
  NAND2_X1 U16142 ( .A1(n14899), .A2(n14980), .ZN(n14902) );
  NAND2_X1 U16143 ( .A1(n14900), .A2(n14978), .ZN(n14901) );
  NAND2_X1 U16144 ( .A1(n14902), .A2(n14901), .ZN(n15056) );
  AND2_X1 U16145 ( .A1(n14903), .A2(n16037), .ZN(n14904) );
  OAI21_X1 U16146 ( .B1(n15056), .B2(n14904), .A(n11899), .ZN(n14906) );
  NAND2_X1 U16147 ( .A1(n15998), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n14905) );
  NAND4_X1 U16148 ( .A1(n14908), .A2(n14907), .A3(n14906), .A4(n14905), .ZN(
        n14909) );
  AOI21_X1 U16149 ( .B1(n15058), .B2(n14910), .A(n14909), .ZN(n14911) );
  OAI21_X1 U16150 ( .B1(n14967), .B2(n15061), .A(n14911), .ZN(P1_U3268) );
  OAI21_X1 U16151 ( .B1(n14918), .B2(n7272), .A(n14912), .ZN(n15062) );
  OAI22_X1 U16152 ( .A1(n14914), .A2(n15005), .B1(n14913), .B2(n15003), .ZN(
        n14920) );
  INV_X1 U16153 ( .A(n14915), .ZN(n14916) );
  AOI211_X1 U16154 ( .C1(n16034), .C2(n15062), .A(n14920), .B(n14919), .ZN(
        n15066) );
  INV_X1 U16155 ( .A(n15064), .ZN(n14926) );
  INV_X1 U16156 ( .A(n14921), .ZN(n14922) );
  AOI211_X1 U16157 ( .C1(n15064), .C2(n14934), .A(n15952), .B(n14922), .ZN(
        n15063) );
  NAND2_X1 U16158 ( .A1(n15063), .A2(n16035), .ZN(n14925) );
  AOI22_X1 U16159 ( .A1(n14923), .A2(n16037), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n15998), .ZN(n14924) );
  OAI211_X1 U16160 ( .C1(n14926), .C2(n16041), .A(n14925), .B(n14924), .ZN(
        n14927) );
  AOI21_X1 U16161 ( .B1(n16044), .B2(n15062), .A(n14927), .ZN(n14928) );
  OAI21_X1 U16162 ( .B1(n15066), .B2(n15998), .A(n14928), .ZN(P1_U3269) );
  OAI21_X1 U16163 ( .B1(n14930), .B2(n14939), .A(n14929), .ZN(n14933) );
  INV_X1 U16164 ( .A(n14931), .ZN(n14932) );
  AOI21_X1 U16165 ( .B1(n14933), .B2(n15955), .A(n14932), .ZN(n15071) );
  INV_X1 U16166 ( .A(n14934), .ZN(n14935) );
  AOI211_X1 U16167 ( .C1(n15069), .C2(n14949), .A(n15952), .B(n14935), .ZN(
        n15068) );
  INV_X1 U16168 ( .A(n15069), .ZN(n14938) );
  AOI22_X1 U16169 ( .A1(n14936), .A2(n16037), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n15998), .ZN(n14937) );
  OAI21_X1 U16170 ( .B1(n14938), .B2(n16041), .A(n14937), .ZN(n14943) );
  NAND2_X1 U16171 ( .A1(n14940), .A2(n14939), .ZN(n14941) );
  NAND2_X1 U16172 ( .A1(n7210), .A2(n14941), .ZN(n15072) );
  NOR2_X1 U16173 ( .A1(n15072), .A2(n14967), .ZN(n14942) );
  AOI211_X1 U16174 ( .C1(n15068), .C2(n16035), .A(n14943), .B(n14942), .ZN(
        n14944) );
  OAI21_X1 U16175 ( .B1(n16047), .B2(n15071), .A(n14944), .ZN(P1_U3270) );
  XNOR2_X1 U16176 ( .A(n14945), .B(n14947), .ZN(n15080) );
  OAI21_X1 U16177 ( .B1(n14948), .B2(n14947), .A(n14946), .ZN(n15078) );
  OAI21_X1 U16178 ( .B1(n15075), .B2(n7213), .A(n14949), .ZN(n15073) );
  AND2_X1 U16179 ( .A1(n14981), .A2(n14978), .ZN(n14950) );
  AOI21_X1 U16180 ( .B1(n14951), .B2(n14980), .A(n14950), .ZN(n15074) );
  OAI21_X1 U16181 ( .B1(n15073), .B2(n14952), .A(n15074), .ZN(n14953) );
  NAND2_X1 U16182 ( .A1(n14953), .A2(n11899), .ZN(n14956) );
  AOI22_X1 U16183 ( .A1(n14954), .A2(n16037), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n15998), .ZN(n14955) );
  OAI211_X1 U16184 ( .C1(n16041), .C2(n15075), .A(n14956), .B(n14955), .ZN(
        n14957) );
  AOI21_X1 U16185 ( .B1(n15078), .B2(n14999), .A(n14957), .ZN(n14958) );
  OAI21_X1 U16186 ( .B1(n15001), .B2(n15080), .A(n14958), .ZN(P1_U3271) );
  XOR2_X1 U16187 ( .A(n14966), .B(n14959), .Z(n14960) );
  AOI222_X1 U16188 ( .A1(n14962), .A2(n14978), .B1(n14961), .B2(n14980), .C1(
        n15955), .C2(n14960), .ZN(n15084) );
  AOI211_X1 U16189 ( .C1(n15082), .C2(n14975), .A(n15952), .B(n7213), .ZN(
        n15081) );
  AOI22_X1 U16190 ( .A1(n14963), .A2(n16037), .B1(n15998), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n14964) );
  OAI21_X1 U16191 ( .B1(n7609), .B2(n16041), .A(n14964), .ZN(n14969) );
  XOR2_X1 U16192 ( .A(n14966), .B(n14965), .Z(n15085) );
  NOR2_X1 U16193 ( .A1(n15085), .A2(n14967), .ZN(n14968) );
  AOI211_X1 U16194 ( .C1(n15081), .C2(n16035), .A(n14969), .B(n14968), .ZN(
        n14970) );
  OAI21_X1 U16195 ( .B1(n15084), .B2(n16047), .A(n14970), .ZN(P1_U3272) );
  OAI21_X1 U16196 ( .B1(n14972), .B2(n14974), .A(n14971), .ZN(n15093) );
  AOI21_X1 U16197 ( .B1(n14974), .B2(n14973), .A(n7249), .ZN(n15091) );
  INV_X1 U16198 ( .A(n14990), .ZN(n14977) );
  OAI21_X1 U16199 ( .B1(n14977), .B2(n14976), .A(n14975), .ZN(n15089) );
  AOI22_X1 U16200 ( .A1(n14981), .A2(n14980), .B1(n14979), .B2(n14978), .ZN(
        n15088) );
  AOI22_X1 U16201 ( .A1(n16047), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n14982), 
        .B2(n16037), .ZN(n14983) );
  OAI21_X1 U16202 ( .B1(n15088), .B2(n15998), .A(n14983), .ZN(n14984) );
  AOI21_X1 U16203 ( .B1(n15086), .B2(n15990), .A(n14984), .ZN(n14985) );
  OAI21_X1 U16204 ( .B1(n15089), .B2(n15840), .A(n14985), .ZN(n14986) );
  AOI21_X1 U16205 ( .B1(n15091), .B2(n14999), .A(n14986), .ZN(n14987) );
  OAI21_X1 U16206 ( .B1(n15001), .B2(n15093), .A(n14987), .ZN(P1_U3273) );
  XNOR2_X1 U16207 ( .A(n14988), .B(n12021), .ZN(n15101) );
  XNOR2_X1 U16208 ( .A(n14989), .B(n12021), .ZN(n15099) );
  OAI211_X1 U16209 ( .C1(n15013), .C2(n15097), .A(n15041), .B(n14990), .ZN(
        n15096) );
  NAND2_X1 U16210 ( .A1(n15094), .A2(n11899), .ZN(n14992) );
  NAND2_X1 U16211 ( .A1(n16047), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n14991) );
  OAI211_X1 U16212 ( .C1(n15016), .C2(n14993), .A(n14992), .B(n14991), .ZN(
        n14994) );
  AOI21_X1 U16213 ( .B1(n14995), .B2(n15990), .A(n14994), .ZN(n14996) );
  OAI21_X1 U16214 ( .B1(n15096), .B2(n14997), .A(n14996), .ZN(n14998) );
  AOI21_X1 U16215 ( .B1(n15099), .B2(n14999), .A(n14998), .ZN(n15000) );
  OAI21_X1 U16216 ( .B1(n15001), .B2(n15101), .A(n15000), .ZN(P1_U3274) );
  XNOR2_X1 U16217 ( .A(n15002), .B(n7955), .ZN(n15102) );
  OAI22_X1 U16218 ( .A1(n15006), .A2(n15005), .B1(n15004), .B2(n15003), .ZN(
        n15012) );
  INV_X1 U16219 ( .A(n15007), .ZN(n15008) );
  AOI211_X1 U16220 ( .C1(n15010), .C2(n15009), .A(n16060), .B(n15008), .ZN(
        n15011) );
  AOI211_X1 U16221 ( .C1(n16034), .C2(n15102), .A(n15012), .B(n15011), .ZN(
        n15106) );
  AOI211_X1 U16222 ( .C1(n15104), .C2(n15014), .A(n15952), .B(n15013), .ZN(
        n15103) );
  INV_X1 U16223 ( .A(n15104), .ZN(n15015) );
  NOR2_X1 U16224 ( .A1(n15015), .A2(n16041), .ZN(n15020) );
  OAI22_X1 U16225 ( .A1(n11899), .A2(n15018), .B1(n15017), .B2(n15016), .ZN(
        n15019) );
  AOI211_X1 U16226 ( .C1(n15103), .C2(n16035), .A(n15020), .B(n15019), .ZN(
        n15022) );
  NAND2_X1 U16227 ( .A1(n15102), .A2(n16044), .ZN(n15021) );
  OAI211_X1 U16228 ( .C1(n15106), .C2(n15998), .A(n15022), .B(n15021), .ZN(
        P1_U3275) );
  OR2_X1 U16229 ( .A1(n15023), .A2(n15952), .ZN(n15026) );
  AOI21_X1 U16230 ( .B1(n15024), .B2(n15948), .A(n15027), .ZN(n15025) );
  NAND2_X1 U16231 ( .A1(n15026), .A2(n15025), .ZN(n15126) );
  MUX2_X1 U16232 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15126), .S(n16067), .Z(
        P1_U3559) );
  AOI21_X1 U16233 ( .B1(n15028), .B2(n15948), .A(n15027), .ZN(n15029) );
  OAI21_X1 U16234 ( .B1(n15030), .B2(n15952), .A(n15029), .ZN(n15127) );
  MUX2_X1 U16235 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15127), .S(n16067), .Z(
        P1_U3558) );
  OAI211_X1 U16236 ( .C1(n7603), .C2(n16058), .A(n15033), .B(n15032), .ZN(
        n15034) );
  AOI21_X1 U16237 ( .B1(n15035), .B2(n15041), .A(n15034), .ZN(n15036) );
  INV_X1 U16238 ( .A(n15039), .ZN(n15045) );
  AOI22_X1 U16239 ( .A1(n15042), .A2(n15041), .B1(n15948), .B2(n15040), .ZN(
        n15043) );
  OAI211_X1 U16240 ( .C1(n15045), .C2(n15933), .A(n15044), .B(n15043), .ZN(
        n15129) );
  MUX2_X1 U16241 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15129), .S(n16067), .Z(
        P1_U3556) );
  NAND2_X1 U16242 ( .A1(n15046), .A2(n16017), .ZN(n15048) );
  OAI211_X1 U16243 ( .C1(n7999), .C2(n16058), .A(n15048), .B(n15047), .ZN(
        n15049) );
  AOI21_X1 U16244 ( .B1(n15948), .B2(n15051), .A(n15050), .ZN(n15052) );
  MUX2_X1 U16245 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15131), .S(n16067), .Z(
        P1_U3554) );
  AOI211_X1 U16246 ( .C1(n15948), .C2(n15057), .A(n15056), .B(n15055), .ZN(
        n15060) );
  NAND2_X1 U16247 ( .A1(n15058), .A2(n15955), .ZN(n15059) );
  OAI211_X1 U16248 ( .C1(n15061), .C2(n15933), .A(n15060), .B(n15059), .ZN(
        n15132) );
  MUX2_X1 U16249 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15132), .S(n16067), .Z(
        P1_U3553) );
  INV_X1 U16250 ( .A(n15062), .ZN(n15067) );
  AOI21_X1 U16251 ( .B1(n15948), .B2(n15064), .A(n15063), .ZN(n15065) );
  OAI211_X1 U16252 ( .C1(n15067), .C2(n15856), .A(n15066), .B(n15065), .ZN(
        n15133) );
  MUX2_X1 U16253 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15133), .S(n16067), .Z(
        P1_U3552) );
  AOI21_X1 U16254 ( .B1(n15948), .B2(n15069), .A(n15068), .ZN(n15070) );
  OAI211_X1 U16255 ( .C1(n15072), .C2(n15933), .A(n15071), .B(n15070), .ZN(
        n15134) );
  MUX2_X1 U16256 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15134), .S(n16067), .Z(
        P1_U3551) );
  NOR2_X1 U16257 ( .A1(n15073), .A2(n15952), .ZN(n15077) );
  OAI21_X1 U16258 ( .B1(n15075), .B2(n16058), .A(n15074), .ZN(n15076) );
  AOI211_X1 U16259 ( .C1(n15078), .C2(n16064), .A(n15077), .B(n15076), .ZN(
        n15079) );
  OAI21_X1 U16260 ( .B1(n16060), .B2(n15080), .A(n15079), .ZN(n15135) );
  MUX2_X1 U16261 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15135), .S(n16067), .Z(
        P1_U3550) );
  AOI21_X1 U16262 ( .B1(n15948), .B2(n15082), .A(n15081), .ZN(n15083) );
  OAI211_X1 U16263 ( .C1(n15933), .C2(n15085), .A(n15084), .B(n15083), .ZN(
        n15136) );
  MUX2_X1 U16264 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15136), .S(n16067), .Z(
        P1_U3549) );
  NAND2_X1 U16265 ( .A1(n15086), .A2(n15948), .ZN(n15087) );
  OAI211_X1 U16266 ( .C1(n15089), .C2(n15952), .A(n15088), .B(n15087), .ZN(
        n15090) );
  AOI21_X1 U16267 ( .B1(n15091), .B2(n16064), .A(n15090), .ZN(n15092) );
  OAI21_X1 U16268 ( .B1(n16060), .B2(n15093), .A(n15092), .ZN(n15137) );
  MUX2_X1 U16269 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15137), .S(n16067), .Z(
        P1_U3548) );
  INV_X1 U16270 ( .A(n15094), .ZN(n15095) );
  OAI211_X1 U16271 ( .C1(n15097), .C2(n16058), .A(n15096), .B(n15095), .ZN(
        n15098) );
  AOI21_X1 U16272 ( .B1(n15099), .B2(n16064), .A(n15098), .ZN(n15100) );
  OAI21_X1 U16273 ( .B1(n15101), .B2(n16060), .A(n15100), .ZN(n15138) );
  MUX2_X1 U16274 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15138), .S(n16067), .Z(
        P1_U3547) );
  INV_X1 U16275 ( .A(n15102), .ZN(n15107) );
  AOI21_X1 U16276 ( .B1(n15948), .B2(n15104), .A(n15103), .ZN(n15105) );
  OAI211_X1 U16277 ( .C1(n15107), .C2(n15856), .A(n15106), .B(n15105), .ZN(
        n15139) );
  MUX2_X1 U16278 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15139), .S(n16067), .Z(
        P1_U3546) );
  OAI21_X1 U16279 ( .B1(n7604), .B2(n16058), .A(n15108), .ZN(n15110) );
  AOI211_X1 U16280 ( .C1(n15955), .C2(n15111), .A(n15110), .B(n15109), .ZN(
        n15112) );
  OAI21_X1 U16281 ( .B1(n15933), .B2(n15113), .A(n15112), .ZN(n15140) );
  MUX2_X1 U16282 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15140), .S(n16067), .Z(
        P1_U3545) );
  OAI211_X1 U16283 ( .C1(n15116), .C2(n16058), .A(n15115), .B(n15114), .ZN(
        n15117) );
  AOI21_X1 U16284 ( .B1(n15118), .B2(n16064), .A(n15117), .ZN(n15119) );
  OAI21_X1 U16285 ( .B1(n15120), .B2(n16060), .A(n15119), .ZN(n15141) );
  MUX2_X1 U16286 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15141), .S(n16067), .Z(
        P1_U3544) );
  AOI21_X1 U16287 ( .B1(n15948), .B2(n15122), .A(n15121), .ZN(n15123) );
  OAI211_X1 U16288 ( .C1(n15933), .C2(n15125), .A(n15124), .B(n15123), .ZN(
        n15142) );
  MUX2_X1 U16289 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15142), .S(n16067), .Z(
        P1_U3543) );
  MUX2_X1 U16290 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15126), .S(n16071), .Z(
        P1_U3527) );
  MUX2_X1 U16291 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15127), .S(n16071), .Z(
        P1_U3526) );
  MUX2_X1 U16292 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n15129), .S(n16071), .Z(
        P1_U3524) );
  MUX2_X1 U16293 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15130), .S(n16071), .Z(
        P1_U3523) );
  MUX2_X1 U16294 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15131), .S(n16071), .Z(
        P1_U3522) );
  MUX2_X1 U16295 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15132), .S(n16071), .Z(
        P1_U3521) );
  MUX2_X1 U16296 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15133), .S(n16071), .Z(
        P1_U3520) );
  MUX2_X1 U16297 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15134), .S(n16071), .Z(
        P1_U3519) );
  MUX2_X1 U16298 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15135), .S(n16071), .Z(
        P1_U3518) );
  MUX2_X1 U16299 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15136), .S(n16071), .Z(
        P1_U3517) );
  MUX2_X1 U16300 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15137), .S(n16071), .Z(
        P1_U3516) );
  MUX2_X1 U16301 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15138), .S(n16071), .Z(
        P1_U3515) );
  MUX2_X1 U16302 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15139), .S(n16071), .Z(
        P1_U3513) );
  MUX2_X1 U16303 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15140), .S(n16071), .Z(
        P1_U3510) );
  MUX2_X1 U16304 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15141), .S(n16071), .Z(
        P1_U3507) );
  MUX2_X1 U16305 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15142), .S(n16071), .Z(
        P1_U3504) );
  MUX2_X1 U16306 ( .A(n15143), .B(P1_D_REG_1__SCAN_IN), .S(n15172), .Z(
        P1_U3446) );
  NOR4_X1 U16307 ( .A1(n15144), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n9069), .ZN(n15145) );
  AOI21_X1 U16308 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n15164), .A(n15145), 
        .ZN(n15146) );
  OAI21_X1 U16309 ( .B1(n15147), .B2(n15167), .A(n15146), .ZN(P1_U3324) );
  OAI222_X1 U16310 ( .A1(n15167), .A2(n15150), .B1(n15149), .B2(P1_U3086), 
        .C1(n15148), .C2(n15157), .ZN(P1_U3326) );
  OAI222_X1 U16311 ( .A1(n15157), .A2(n15153), .B1(n15167), .B2(n15152), .C1(
        P1_U3086), .C2(n15151), .ZN(P1_U3327) );
  OAI222_X1 U16312 ( .A1(n15157), .A2(n15156), .B1(n15167), .B2(n15155), .C1(
        P1_U3086), .C2(n15154), .ZN(P1_U3328) );
  OAI222_X1 U16313 ( .A1(n15167), .A2(n15160), .B1(P1_U3086), .B2(n15159), 
        .C1(n15158), .C2(n15157), .ZN(P1_U3329) );
  OAI222_X1 U16314 ( .A1(n15157), .A2(n15163), .B1(n15167), .B2(n15162), .C1(
        n15161), .C2(P1_U3086), .ZN(P1_U3330) );
  AOI22_X1 U16315 ( .A1(n15165), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n15164), .ZN(n15166) );
  OAI21_X1 U16316 ( .B1(n15168), .B2(n15167), .A(n15166), .ZN(P1_U3331) );
  MUX2_X1 U16317 ( .A(n15170), .B(n15169), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16318 ( .A(n15171), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AND2_X1 U16319 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15172), .ZN(P1_U3323) );
  AND2_X1 U16320 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15172), .ZN(P1_U3322) );
  AND2_X1 U16321 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15172), .ZN(P1_U3321) );
  AND2_X1 U16322 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15172), .ZN(P1_U3320) );
  AND2_X1 U16323 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15172), .ZN(P1_U3319) );
  AND2_X1 U16324 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15172), .ZN(P1_U3318) );
  AND2_X1 U16325 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15172), .ZN(P1_U3317) );
  AND2_X1 U16326 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15172), .ZN(P1_U3316) );
  AND2_X1 U16327 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15172), .ZN(P1_U3315) );
  AND2_X1 U16328 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15172), .ZN(P1_U3314) );
  AND2_X1 U16329 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15172), .ZN(P1_U3313) );
  AND2_X1 U16330 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15172), .ZN(P1_U3312) );
  AND2_X1 U16331 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15172), .ZN(P1_U3311) );
  AND2_X1 U16332 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15172), .ZN(P1_U3310) );
  AND2_X1 U16333 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15172), .ZN(P1_U3309) );
  AND2_X1 U16334 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15172), .ZN(P1_U3308) );
  AND2_X1 U16335 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15172), .ZN(P1_U3307) );
  AND2_X1 U16336 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15172), .ZN(P1_U3306) );
  AND2_X1 U16337 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15172), .ZN(P1_U3305) );
  AND2_X1 U16338 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15172), .ZN(P1_U3304) );
  AND2_X1 U16339 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15172), .ZN(P1_U3303) );
  AND2_X1 U16340 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15172), .ZN(P1_U3302) );
  AND2_X1 U16341 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15172), .ZN(P1_U3301) );
  AND2_X1 U16342 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15172), .ZN(P1_U3300) );
  AND2_X1 U16343 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15172), .ZN(P1_U3299) );
  AND2_X1 U16344 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15172), .ZN(P1_U3298) );
  AND2_X1 U16345 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15172), .ZN(P1_U3297) );
  AND2_X1 U16346 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15172), .ZN(P1_U3296) );
  AND2_X1 U16347 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15172), .ZN(P1_U3295) );
  AND2_X1 U16348 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15172), .ZN(P1_U3294) );
  INV_X1 U16349 ( .A(n15173), .ZN(n15174) );
  AOI21_X1 U16350 ( .B1(n15175), .B2(n15406), .A(n15174), .ZN(P2_U3417) );
  AND2_X1 U16351 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15177), .ZN(P2_U3295) );
  AND2_X1 U16352 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15177), .ZN(P2_U3294) );
  AND2_X1 U16353 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15177), .ZN(P2_U3293) );
  AND2_X1 U16354 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15177), .ZN(P2_U3292) );
  AND2_X1 U16355 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15177), .ZN(P2_U3291) );
  AND2_X1 U16356 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15177), .ZN(P2_U3290) );
  AND2_X1 U16357 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15177), .ZN(P2_U3289) );
  AND2_X1 U16358 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15177), .ZN(P2_U3288) );
  AND2_X1 U16359 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15177), .ZN(P2_U3287) );
  AND2_X1 U16360 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15177), .ZN(P2_U3286) );
  AND2_X1 U16361 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15177), .ZN(P2_U3285) );
  AND2_X1 U16362 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15177), .ZN(P2_U3284) );
  AND2_X1 U16363 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15177), .ZN(P2_U3283) );
  AND2_X1 U16364 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15177), .ZN(P2_U3282) );
  AND2_X1 U16365 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15177), .ZN(P2_U3281) );
  AND2_X1 U16366 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15177), .ZN(P2_U3280) );
  AND2_X1 U16367 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15177), .ZN(P2_U3279) );
  AND2_X1 U16368 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15177), .ZN(P2_U3278) );
  AND2_X1 U16369 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15177), .ZN(P2_U3277) );
  AND2_X1 U16370 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15177), .ZN(P2_U3276) );
  AND2_X1 U16371 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15177), .ZN(P2_U3275) );
  AND2_X1 U16372 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15177), .ZN(P2_U3274) );
  AND2_X1 U16373 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15177), .ZN(P2_U3273) );
  AND2_X1 U16374 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15177), .ZN(P2_U3272) );
  AND2_X1 U16375 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15177), .ZN(P2_U3271) );
  AND2_X1 U16376 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15177), .ZN(P2_U3270) );
  AND2_X1 U16377 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15177), .ZN(P2_U3269) );
  AND2_X1 U16378 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15177), .ZN(P2_U3268) );
  AND2_X1 U16379 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15177), .ZN(P2_U3267) );
  AND2_X1 U16380 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15177), .ZN(P2_U3266) );
  NOR2_X1 U16381 ( .A1(n15471), .A2(P2_U3947), .ZN(P2_U3087) );
  NOR2_X1 U16382 ( .A1(P3_U3897), .A2(n15771), .ZN(P3_U3150) );
  XOR2_X1 U16383 ( .A(keyinput_119), .B(P3_REG3_REG_20__SCAN_IN), .Z(n15270)
         );
  INV_X1 U16384 ( .A(keyinput_118), .ZN(n15266) );
  OAI22_X1 U16385 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(keyinput_105), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(keyinput_104), .ZN(n15178) );
  AOI221_X1 U16386 ( .B1(P3_REG3_REG_19__SCAN_IN), .B2(keyinput_105), .C1(
        keyinput_104), .C2(P3_REG3_REG_3__SCAN_IN), .A(n15178), .ZN(n15246) );
  INV_X1 U16387 ( .A(keyinput_103), .ZN(n15241) );
  INV_X1 U16388 ( .A(keyinput_102), .ZN(n15239) );
  INV_X1 U16389 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n15344) );
  INV_X1 U16390 ( .A(keyinput_98), .ZN(n15233) );
  AOI22_X1 U16391 ( .A1(n15181), .A2(keyinput_74), .B1(keyinput_77), .B2(
        n15180), .ZN(n15179) );
  OAI221_X1 U16392 ( .B1(n15181), .B2(keyinput_74), .C1(n15180), .C2(
        keyinput_77), .A(n15179), .ZN(n15186) );
  AOI22_X1 U16393 ( .A1(n15184), .A2(keyinput_78), .B1(n15183), .B2(
        keyinput_75), .ZN(n15182) );
  OAI221_X1 U16394 ( .B1(n15184), .B2(keyinput_78), .C1(n15183), .C2(
        keyinput_75), .A(n15182), .ZN(n15185) );
  AOI211_X1 U16395 ( .C1(keyinput_76), .C2(SI_20_), .A(n15186), .B(n15185), 
        .ZN(n15187) );
  OAI21_X1 U16396 ( .B1(keyinput_76), .B2(SI_20_), .A(n15187), .ZN(n15203) );
  OAI22_X1 U16397 ( .A1(n15287), .A2(keyinput_73), .B1(SI_25_), .B2(
        keyinput_71), .ZN(n15188) );
  AOI221_X1 U16398 ( .B1(n15287), .B2(keyinput_73), .C1(keyinput_71), .C2(
        SI_25_), .A(n15188), .ZN(n15199) );
  INV_X1 U16399 ( .A(keyinput_70), .ZN(n15197) );
  INV_X1 U16400 ( .A(keyinput_69), .ZN(n15195) );
  OAI22_X1 U16401 ( .A1(n15289), .A2(keyinput_67), .B1(keyinput_66), .B2(
        SI_30_), .ZN(n15189) );
  AOI221_X1 U16402 ( .B1(n15289), .B2(keyinput_67), .C1(SI_30_), .C2(
        keyinput_66), .A(n15189), .ZN(n15192) );
  AOI22_X1 U16403 ( .A1(P3_WR_REG_SCAN_IN), .A2(keyinput_64), .B1(SI_31_), 
        .B2(keyinput_65), .ZN(n15190) );
  OAI221_X1 U16404 ( .B1(P3_WR_REG_SCAN_IN), .B2(keyinput_64), .C1(SI_31_), 
        .C2(keyinput_65), .A(n15190), .ZN(n15191) );
  AOI22_X1 U16405 ( .A1(n15192), .A2(n15191), .B1(keyinput_68), .B2(SI_28_), 
        .ZN(n15193) );
  OAI21_X1 U16406 ( .B1(keyinput_68), .B2(SI_28_), .A(n15193), .ZN(n15194) );
  OAI221_X1 U16407 ( .B1(SI_27_), .B2(keyinput_69), .C1(n15297), .C2(n15195), 
        .A(n15194), .ZN(n15196) );
  OAI221_X1 U16408 ( .B1(SI_26_), .B2(n15197), .C1(n15301), .C2(keyinput_70), 
        .A(n15196), .ZN(n15198) );
  OAI211_X1 U16409 ( .C1(n15201), .C2(keyinput_72), .A(n15199), .B(n15198), 
        .ZN(n15200) );
  AOI21_X1 U16410 ( .B1(n15201), .B2(keyinput_72), .A(n15200), .ZN(n15202) );
  OAI22_X1 U16411 ( .A1(keyinput_79), .A2(n15205), .B1(n15203), .B2(n15202), 
        .ZN(n15204) );
  AOI21_X1 U16412 ( .B1(keyinput_79), .B2(n15205), .A(n15204), .ZN(n15223) );
  AOI22_X1 U16413 ( .A1(n15208), .A2(keyinput_85), .B1(n15207), .B2(
        keyinput_80), .ZN(n15206) );
  OAI221_X1 U16414 ( .B1(n15208), .B2(keyinput_85), .C1(n15207), .C2(
        keyinput_80), .A(n15206), .ZN(n15214) );
  XNOR2_X1 U16415 ( .A(SI_6_), .B(keyinput_90), .ZN(n15212) );
  XNOR2_X1 U16416 ( .A(SI_10_), .B(keyinput_86), .ZN(n15211) );
  XNOR2_X1 U16417 ( .A(SI_7_), .B(keyinput_89), .ZN(n15210) );
  XNOR2_X1 U16418 ( .A(SI_9_), .B(keyinput_87), .ZN(n15209) );
  NAND4_X1 U16419 ( .A1(n15212), .A2(n15211), .A3(n15210), .A4(n15209), .ZN(
        n15213) );
  NOR2_X1 U16420 ( .A1(n15214), .A2(n15213), .ZN(n15221) );
  OAI22_X1 U16421 ( .A1(SI_13_), .A2(keyinput_83), .B1(keyinput_88), .B2(SI_8_), .ZN(n15215) );
  AOI221_X1 U16422 ( .B1(SI_13_), .B2(keyinput_83), .C1(SI_8_), .C2(
        keyinput_88), .A(n15215), .ZN(n15220) );
  OAI22_X1 U16423 ( .A1(SI_14_), .A2(keyinput_82), .B1(SI_12_), .B2(
        keyinput_84), .ZN(n15216) );
  AOI221_X1 U16424 ( .B1(SI_14_), .B2(keyinput_82), .C1(keyinput_84), .C2(
        SI_12_), .A(n15216), .ZN(n15219) );
  OAI22_X1 U16425 ( .A1(SI_15_), .A2(keyinput_81), .B1(SI_5_), .B2(keyinput_91), .ZN(n15217) );
  AOI221_X1 U16426 ( .B1(SI_15_), .B2(keyinput_81), .C1(keyinput_91), .C2(
        SI_5_), .A(n15217), .ZN(n15218) );
  NAND4_X1 U16427 ( .A1(n15221), .A2(n15220), .A3(n15219), .A4(n15218), .ZN(
        n15222) );
  NOR2_X1 U16428 ( .A1(n15223), .A2(n15222), .ZN(n15231) );
  AOI22_X1 U16429 ( .A1(P3_RD_REG_SCAN_IN), .A2(keyinput_97), .B1(SI_1_), .B2(
        keyinput_95), .ZN(n15224) );
  OAI221_X1 U16430 ( .B1(P3_RD_REG_SCAN_IN), .B2(keyinput_97), .C1(SI_1_), 
        .C2(keyinput_95), .A(n15224), .ZN(n15230) );
  XOR2_X1 U16431 ( .A(SI_0_), .B(keyinput_96), .Z(n15228) );
  XNOR2_X1 U16432 ( .A(SI_3_), .B(keyinput_93), .ZN(n15227) );
  XNOR2_X1 U16433 ( .A(SI_4_), .B(keyinput_92), .ZN(n15226) );
  XNOR2_X1 U16434 ( .A(SI_2_), .B(keyinput_94), .ZN(n15225) );
  NAND4_X1 U16435 ( .A1(n15228), .A2(n15227), .A3(n15226), .A4(n15225), .ZN(
        n15229) );
  NOR3_X1 U16436 ( .A1(n15231), .A2(n15230), .A3(n15229), .ZN(n15232) );
  AOI221_X1 U16437 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n15233), .C1(P3_U3151), 
        .C2(keyinput_98), .A(n15232), .ZN(n15236) );
  AOI22_X1 U16438 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(keyinput_99), .B1(
        P3_REG3_REG_27__SCAN_IN), .B2(keyinput_100), .ZN(n15234) );
  OAI221_X1 U16439 ( .B1(P3_REG3_REG_7__SCAN_IN), .B2(keyinput_99), .C1(
        P3_REG3_REG_27__SCAN_IN), .C2(keyinput_100), .A(n15234), .ZN(n15235)
         );
  AOI211_X1 U16440 ( .C1(P3_REG3_REG_14__SCAN_IN), .C2(keyinput_101), .A(
        n15236), .B(n15235), .ZN(n15237) );
  OAI21_X1 U16441 ( .B1(P3_REG3_REG_14__SCAN_IN), .B2(keyinput_101), .A(n15237), .ZN(n15238) );
  OAI221_X1 U16442 ( .B1(P3_REG3_REG_23__SCAN_IN), .B2(n15239), .C1(n15344), 
        .C2(keyinput_102), .A(n15238), .ZN(n15240) );
  OAI221_X1 U16443 ( .B1(P3_REG3_REG_10__SCAN_IN), .B2(keyinput_103), .C1(
        n15347), .C2(n15241), .A(n15240), .ZN(n15245) );
  INV_X1 U16444 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n15243) );
  AOI22_X1 U16445 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(keyinput_107), .B1(n15243), .B2(keyinput_106), .ZN(n15242) );
  OAI221_X1 U16446 ( .B1(P3_REG3_REG_8__SCAN_IN), .B2(keyinput_107), .C1(
        n15243), .C2(keyinput_106), .A(n15242), .ZN(n15244) );
  AOI21_X1 U16447 ( .B1(n15246), .B2(n15245), .A(n15244), .ZN(n15259) );
  INV_X1 U16448 ( .A(keyinput_108), .ZN(n15247) );
  MUX2_X1 U16449 ( .A(n15247), .B(keyinput_108), .S(P3_REG3_REG_1__SCAN_IN), 
        .Z(n15258) );
  AOI22_X1 U16450 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(keyinput_110), .B1(
        P3_REG3_REG_17__SCAN_IN), .B2(keyinput_114), .ZN(n15248) );
  OAI221_X1 U16451 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_110), .C1(
        P3_REG3_REG_17__SCAN_IN), .C2(keyinput_114), .A(n15248), .ZN(n15256)
         );
  INV_X1 U16452 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n15251) );
  AOI22_X1 U16453 ( .A1(n15251), .A2(keyinput_112), .B1(n15250), .B2(
        keyinput_111), .ZN(n15249) );
  OAI221_X1 U16454 ( .B1(n15251), .B2(keyinput_112), .C1(n15250), .C2(
        keyinput_111), .A(n15249), .ZN(n15255) );
  AOI22_X1 U16455 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(keyinput_113), .B1(n15253), .B2(keyinput_109), .ZN(n15252) );
  OAI221_X1 U16456 ( .B1(P3_REG3_REG_5__SCAN_IN), .B2(keyinput_113), .C1(
        n15253), .C2(keyinput_109), .A(n15252), .ZN(n15254) );
  NOR3_X1 U16457 ( .A1(n15256), .A2(n15255), .A3(n15254), .ZN(n15257) );
  OAI21_X1 U16458 ( .B1(n15259), .B2(n15258), .A(n15257), .ZN(n15260) );
  INV_X1 U16459 ( .A(n15260), .ZN(n15263) );
  AOI22_X1 U16460 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(keyinput_115), .B1(
        n15365), .B2(keyinput_116), .ZN(n15261) );
  OAI221_X1 U16461 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput_115), .C1(
        n15365), .C2(keyinput_116), .A(n15261), .ZN(n15262) );
  AOI211_X1 U16462 ( .C1(P3_REG3_REG_9__SCAN_IN), .C2(keyinput_117), .A(n15263), .B(n15262), .ZN(n15264) );
  OAI21_X1 U16463 ( .B1(P3_REG3_REG_9__SCAN_IN), .B2(keyinput_117), .A(n15264), 
        .ZN(n15265) );
  OAI221_X1 U16464 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput_118), .C1(
        n15658), .C2(n15266), .A(n15265), .ZN(n15269) );
  INV_X1 U16465 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n15372) );
  AOI22_X1 U16466 ( .A1(n15891), .A2(keyinput_123), .B1(n15372), .B2(
        keyinput_121), .ZN(n15267) );
  OAI221_X1 U16467 ( .B1(n15891), .B2(keyinput_123), .C1(n15372), .C2(
        keyinput_121), .A(n15267), .ZN(n15268) );
  AOI21_X1 U16468 ( .B1(n15270), .B2(n15269), .A(n15268), .ZN(n15279) );
  OAI22_X1 U16469 ( .A1(n15272), .A2(keyinput_120), .B1(
        P3_REG3_REG_11__SCAN_IN), .B2(keyinput_122), .ZN(n15271) );
  AOI221_X1 U16470 ( .B1(n15272), .B2(keyinput_120), .C1(keyinput_122), .C2(
        P3_REG3_REG_11__SCAN_IN), .A(n15271), .ZN(n15278) );
  INV_X1 U16471 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n15381) );
  INV_X1 U16472 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n15382) );
  AOI22_X1 U16473 ( .A1(n15381), .A2(keyinput_126), .B1(keyinput_124), .B2(
        n15382), .ZN(n15273) );
  OAI221_X1 U16474 ( .B1(n15381), .B2(keyinput_126), .C1(n15382), .C2(
        keyinput_124), .A(n15273), .ZN(n15277) );
  AOI22_X1 U16475 ( .A1(P3_REG3_REG_15__SCAN_IN), .A2(keyinput_127), .B1(
        n15275), .B2(keyinput_125), .ZN(n15274) );
  OAI221_X1 U16476 ( .B1(P3_REG3_REG_15__SCAN_IN), .B2(keyinput_127), .C1(
        n15275), .C2(keyinput_125), .A(n15274), .ZN(n15276) );
  AOI211_X1 U16477 ( .C1(n15279), .C2(n15278), .A(n15277), .B(n15276), .ZN(
        n15386) );
  XNOR2_X1 U16478 ( .A(P3_REG3_REG_20__SCAN_IN), .B(keyinput_55), .ZN(n15378)
         );
  INV_X1 U16479 ( .A(keyinput_54), .ZN(n15370) );
  OAI22_X1 U16480 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(keyinput_41), .B1(
        keyinput_40), .B2(P3_REG3_REG_3__SCAN_IN), .ZN(n15280) );
  AOI221_X1 U16481 ( .B1(P3_REG3_REG_19__SCAN_IN), .B2(keyinput_41), .C1(
        P3_REG3_REG_3__SCAN_IN), .C2(keyinput_40), .A(n15280), .ZN(n15351) );
  INV_X1 U16482 ( .A(keyinput_39), .ZN(n15346) );
  INV_X1 U16483 ( .A(keyinput_38), .ZN(n15343) );
  INV_X1 U16484 ( .A(keyinput_34), .ZN(n15336) );
  AOI22_X1 U16485 ( .A1(SI_18_), .A2(keyinput_14), .B1(SI_19_), .B2(
        keyinput_13), .ZN(n15281) );
  OAI221_X1 U16486 ( .B1(SI_18_), .B2(keyinput_14), .C1(SI_19_), .C2(
        keyinput_13), .A(n15281), .ZN(n15284) );
  AOI22_X1 U16487 ( .A1(SI_20_), .A2(keyinput_12), .B1(SI_21_), .B2(
        keyinput_11), .ZN(n15282) );
  OAI221_X1 U16488 ( .B1(SI_20_), .B2(keyinput_12), .C1(SI_21_), .C2(
        keyinput_11), .A(n15282), .ZN(n15283) );
  AOI211_X1 U16489 ( .C1(keyinput_10), .C2(SI_22_), .A(n15284), .B(n15283), 
        .ZN(n15285) );
  OAI21_X1 U16490 ( .B1(keyinput_10), .B2(SI_22_), .A(n15285), .ZN(n15306) );
  OAI22_X1 U16491 ( .A1(n15287), .A2(keyinput_9), .B1(keyinput_7), .B2(SI_25_), 
        .ZN(n15286) );
  AOI221_X1 U16492 ( .B1(n15287), .B2(keyinput_9), .C1(SI_25_), .C2(keyinput_7), .A(n15286), .ZN(n15303) );
  INV_X1 U16493 ( .A(keyinput_6), .ZN(n15300) );
  INV_X1 U16494 ( .A(keyinput_5), .ZN(n15298) );
  AOI22_X1 U16495 ( .A1(n15290), .A2(keyinput_2), .B1(n15289), .B2(keyinput_3), 
        .ZN(n15288) );
  OAI221_X1 U16496 ( .B1(n15290), .B2(keyinput_2), .C1(n15289), .C2(keyinput_3), .A(n15288), .ZN(n15295) );
  OAI22_X1 U16497 ( .A1(SI_31_), .A2(keyinput_1), .B1(keyinput_0), .B2(
        P3_WR_REG_SCAN_IN), .ZN(n15291) );
  AOI221_X1 U16498 ( .B1(SI_31_), .B2(keyinput_1), .C1(P3_WR_REG_SCAN_IN), 
        .C2(keyinput_0), .A(n15291), .ZN(n15294) );
  NAND2_X1 U16499 ( .A1(n15293), .A2(keyinput_4), .ZN(n15292) );
  OAI221_X1 U16500 ( .B1(n15295), .B2(n15294), .C1(n15293), .C2(keyinput_4), 
        .A(n15292), .ZN(n15296) );
  OAI221_X1 U16501 ( .B1(SI_27_), .B2(n15298), .C1(n15297), .C2(keyinput_5), 
        .A(n15296), .ZN(n15299) );
  OAI221_X1 U16502 ( .B1(SI_26_), .B2(keyinput_6), .C1(n15301), .C2(n15300), 
        .A(n15299), .ZN(n15302) );
  OAI211_X1 U16503 ( .C1(SI_24_), .C2(keyinput_8), .A(n15303), .B(n15302), 
        .ZN(n15304) );
  AOI21_X1 U16504 ( .B1(SI_24_), .B2(keyinput_8), .A(n15304), .ZN(n15305) );
  OAI22_X1 U16505 ( .A1(n15306), .A2(n15305), .B1(keyinput_15), .B2(SI_17_), 
        .ZN(n15307) );
  AOI21_X1 U16506 ( .B1(keyinput_15), .B2(SI_17_), .A(n15307), .ZN(n15325) );
  OAI22_X1 U16507 ( .A1(SI_16_), .A2(keyinput_16), .B1(SI_15_), .B2(
        keyinput_17), .ZN(n15308) );
  AOI221_X1 U16508 ( .B1(SI_16_), .B2(keyinput_16), .C1(keyinput_17), .C2(
        SI_15_), .A(n15308), .ZN(n15316) );
  OAI22_X1 U16509 ( .A1(SI_11_), .A2(keyinput_21), .B1(keyinput_22), .B2(
        SI_10_), .ZN(n15309) );
  AOI221_X1 U16510 ( .B1(SI_11_), .B2(keyinput_21), .C1(SI_10_), .C2(
        keyinput_22), .A(n15309), .ZN(n15315) );
  OAI22_X1 U16511 ( .A1(n15311), .A2(keyinput_19), .B1(keyinput_23), .B2(SI_9_), .ZN(n15310) );
  AOI221_X1 U16512 ( .B1(n15311), .B2(keyinput_19), .C1(SI_9_), .C2(
        keyinput_23), .A(n15310), .ZN(n15314) );
  OAI22_X1 U16513 ( .A1(SI_8_), .A2(keyinput_24), .B1(keyinput_26), .B2(SI_6_), 
        .ZN(n15312) );
  AOI221_X1 U16514 ( .B1(SI_8_), .B2(keyinput_24), .C1(SI_6_), .C2(keyinput_26), .A(n15312), .ZN(n15313) );
  NAND4_X1 U16515 ( .A1(n15316), .A2(n15315), .A3(n15314), .A4(n15313), .ZN(
        n15324) );
  AOI22_X1 U16516 ( .A1(n15319), .A2(keyinput_20), .B1(n15318), .B2(
        keyinput_18), .ZN(n15317) );
  OAI221_X1 U16517 ( .B1(n15319), .B2(keyinput_20), .C1(n15318), .C2(
        keyinput_18), .A(n15317), .ZN(n15323) );
  XNOR2_X1 U16518 ( .A(SI_5_), .B(keyinput_27), .ZN(n15321) );
  XNOR2_X1 U16519 ( .A(SI_7_), .B(keyinput_25), .ZN(n15320) );
  NAND2_X1 U16520 ( .A1(n15321), .A2(n15320), .ZN(n15322) );
  NOR4_X1 U16521 ( .A1(n15325), .A2(n15324), .A3(n15323), .A4(n15322), .ZN(
        n15334) );
  INV_X1 U16522 ( .A(P3_RD_REG_SCAN_IN), .ZN(n15827) );
  AOI22_X1 U16523 ( .A1(n15827), .A2(keyinput_33), .B1(n9297), .B2(keyinput_32), .ZN(n15326) );
  OAI221_X1 U16524 ( .B1(n15827), .B2(keyinput_33), .C1(n9297), .C2(
        keyinput_32), .A(n15326), .ZN(n15333) );
  AOI22_X1 U16525 ( .A1(SI_3_), .A2(keyinput_29), .B1(n15328), .B2(keyinput_30), .ZN(n15327) );
  OAI221_X1 U16526 ( .B1(SI_3_), .B2(keyinput_29), .C1(n15328), .C2(
        keyinput_30), .A(n15327), .ZN(n15332) );
  XOR2_X1 U16527 ( .A(n8991), .B(keyinput_31), .Z(n15330) );
  XNOR2_X1 U16528 ( .A(SI_4_), .B(keyinput_28), .ZN(n15329) );
  NAND2_X1 U16529 ( .A1(n15330), .A2(n15329), .ZN(n15331) );
  NOR4_X1 U16530 ( .A1(n15334), .A2(n15333), .A3(n15332), .A4(n15331), .ZN(
        n15335) );
  AOI221_X1 U16531 ( .B1(P3_STATE_REG_SCAN_IN), .B2(keyinput_34), .C1(P3_U3151), .C2(n15336), .A(n15335), .ZN(n15340) );
  AOI22_X1 U16532 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(keyinput_37), .B1(n15338), .B2(keyinput_35), .ZN(n15337) );
  OAI221_X1 U16533 ( .B1(P3_REG3_REG_14__SCAN_IN), .B2(keyinput_37), .C1(
        n15338), .C2(keyinput_35), .A(n15337), .ZN(n15339) );
  AOI211_X1 U16534 ( .C1(P3_REG3_REG_27__SCAN_IN), .C2(keyinput_36), .A(n15340), .B(n15339), .ZN(n15341) );
  OAI21_X1 U16535 ( .B1(P3_REG3_REG_27__SCAN_IN), .B2(keyinput_36), .A(n15341), 
        .ZN(n15342) );
  OAI221_X1 U16536 ( .B1(P3_REG3_REG_23__SCAN_IN), .B2(keyinput_38), .C1(
        n15344), .C2(n15343), .A(n15342), .ZN(n15345) );
  OAI221_X1 U16537 ( .B1(P3_REG3_REG_10__SCAN_IN), .B2(keyinput_39), .C1(
        n15347), .C2(n15346), .A(n15345), .ZN(n15350) );
  AOI22_X1 U16538 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(keyinput_43), .B1(
        P3_REG3_REG_28__SCAN_IN), .B2(keyinput_42), .ZN(n15348) );
  OAI221_X1 U16539 ( .B1(P3_REG3_REG_8__SCAN_IN), .B2(keyinput_43), .C1(
        P3_REG3_REG_28__SCAN_IN), .C2(keyinput_42), .A(n15348), .ZN(n15349) );
  AOI21_X1 U16540 ( .B1(n15351), .B2(n15350), .A(n15349), .ZN(n15362) );
  INV_X1 U16541 ( .A(keyinput_44), .ZN(n15352) );
  MUX2_X1 U16542 ( .A(n15352), .B(keyinput_44), .S(P3_REG3_REG_1__SCAN_IN), 
        .Z(n15361) );
  AOI22_X1 U16543 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(keyinput_49), .B1(
        P3_REG3_REG_12__SCAN_IN), .B2(keyinput_46), .ZN(n15353) );
  OAI221_X1 U16544 ( .B1(P3_REG3_REG_5__SCAN_IN), .B2(keyinput_49), .C1(
        P3_REG3_REG_12__SCAN_IN), .C2(keyinput_46), .A(n15353), .ZN(n15359) );
  AOI22_X1 U16545 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(keyinput_48), .B1(
        P3_REG3_REG_25__SCAN_IN), .B2(keyinput_47), .ZN(n15354) );
  OAI221_X1 U16546 ( .B1(P3_REG3_REG_16__SCAN_IN), .B2(keyinput_48), .C1(
        P3_REG3_REG_25__SCAN_IN), .C2(keyinput_47), .A(n15354), .ZN(n15358) );
  AOI22_X1 U16547 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(keyinput_45), .B1(n15356), .B2(keyinput_50), .ZN(n15355) );
  OAI221_X1 U16548 ( .B1(P3_REG3_REG_21__SCAN_IN), .B2(keyinput_45), .C1(
        n15356), .C2(keyinput_50), .A(n15355), .ZN(n15357) );
  NOR3_X1 U16549 ( .A1(n15359), .A2(n15358), .A3(n15357), .ZN(n15360) );
  OAI21_X1 U16550 ( .B1(n15362), .B2(n15361), .A(n15360), .ZN(n15363) );
  INV_X1 U16551 ( .A(n15363), .ZN(n15367) );
  AOI22_X1 U16552 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(keyinput_53), .B1(n15365), 
        .B2(keyinput_52), .ZN(n15364) );
  OAI221_X1 U16553 ( .B1(P3_REG3_REG_9__SCAN_IN), .B2(keyinput_53), .C1(n15365), .C2(keyinput_52), .A(n15364), .ZN(n15366) );
  AOI211_X1 U16554 ( .C1(P3_REG3_REG_24__SCAN_IN), .C2(keyinput_51), .A(n15367), .B(n15366), .ZN(n15368) );
  OAI21_X1 U16555 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput_51), .A(n15368), 
        .ZN(n15369) );
  OAI221_X1 U16556 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput_54), .C1(n15658), .C2(n15370), .A(n15369), .ZN(n15377) );
  AOI22_X1 U16557 ( .A1(n15373), .A2(keyinput_58), .B1(n15372), .B2(
        keyinput_57), .ZN(n15371) );
  OAI221_X1 U16558 ( .B1(n15373), .B2(keyinput_58), .C1(n15372), .C2(
        keyinput_57), .A(n15371), .ZN(n15376) );
  AOI22_X1 U16559 ( .A1(P3_REG3_REG_13__SCAN_IN), .A2(keyinput_56), .B1(n15891), .B2(keyinput_59), .ZN(n15374) );
  OAI221_X1 U16560 ( .B1(P3_REG3_REG_13__SCAN_IN), .B2(keyinput_56), .C1(
        n15891), .C2(keyinput_59), .A(n15374), .ZN(n15375) );
  AOI211_X1 U16561 ( .C1(n15378), .C2(n15377), .A(n15376), .B(n15375), .ZN(
        n15385) );
  AOI22_X1 U16562 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(keyinput_61), .B1(n8195), 
        .B2(keyinput_63), .ZN(n15379) );
  OAI221_X1 U16563 ( .B1(P3_REG3_REG_6__SCAN_IN), .B2(keyinput_61), .C1(n8195), 
        .C2(keyinput_63), .A(n15379), .ZN(n15384) );
  AOI22_X1 U16564 ( .A1(n15382), .A2(keyinput_60), .B1(n15381), .B2(
        keyinput_62), .ZN(n15380) );
  OAI221_X1 U16565 ( .B1(n15382), .B2(keyinput_60), .C1(n15381), .C2(
        keyinput_62), .A(n15380), .ZN(n15383) );
  NOR4_X1 U16566 ( .A1(n15386), .A2(n15385), .A3(n15384), .A4(n15383), .ZN(
        n15405) );
  XNOR2_X1 U16567 ( .A(n7362), .B(n15388), .ZN(n16098) );
  XNOR2_X1 U16568 ( .A(n15389), .B(n15388), .ZN(n15395) );
  OAI22_X1 U16569 ( .A1(n15393), .A2(n15392), .B1(n15391), .B2(n15390), .ZN(
        n15394) );
  AOI21_X1 U16570 ( .B1(n15395), .B2(n15881), .A(n15394), .ZN(n15396) );
  OAI21_X1 U16571 ( .B1(n15886), .B2(n16098), .A(n15396), .ZN(n16100) );
  OAI22_X1 U16572 ( .A1(n15899), .A2(n8327), .B1(n15397), .B2(n15892), .ZN(
        n15398) );
  AOI21_X1 U16573 ( .B1(n15400), .B2(n15399), .A(n15398), .ZN(n15401) );
  OAI21_X1 U16574 ( .B1(n16098), .B2(n15402), .A(n15401), .ZN(n15403) );
  AOI21_X1 U16575 ( .B1(n16100), .B2(n15899), .A(n15403), .ZN(n15404) );
  XNOR2_X1 U16576 ( .A(n15405), .B(n15404), .ZN(P3_U3220) );
  INV_X1 U16577 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15407) );
  AOI22_X1 U16578 ( .A1(n15409), .A2(n15408), .B1(n15407), .B2(n15406), .ZN(
        P2_U3416) );
  OAI22_X1 U16579 ( .A1(n15466), .A2(n15410), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9585), .ZN(n15411) );
  AOI21_X1 U16580 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n15471), .A(n15411), .ZN(
        n15420) );
  OAI211_X1 U16581 ( .C1(n15414), .C2(n15413), .A(n15477), .B(n15412), .ZN(
        n15419) );
  OAI211_X1 U16582 ( .C1(n15417), .C2(n15416), .A(n15473), .B(n15415), .ZN(
        n15418) );
  NAND3_X1 U16583 ( .A1(n15420), .A2(n15419), .A3(n15418), .ZN(P2_U3217) );
  OAI21_X1 U16584 ( .B1(n15469), .B2(n15421), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15422) );
  OAI21_X1 U16585 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15422), .ZN(n15432) );
  OAI211_X1 U16586 ( .C1(n15425), .C2(n15424), .A(n15477), .B(n15423), .ZN(
        n15431) );
  OAI211_X1 U16587 ( .C1(n15428), .C2(n15427), .A(n15473), .B(n15426), .ZN(
        n15430) );
  NAND2_X1 U16588 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n15471), .ZN(n15429) );
  NAND4_X1 U16589 ( .A1(n15432), .A2(n15431), .A3(n15430), .A4(n15429), .ZN(
        P2_U3219) );
  OAI211_X1 U16590 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n15434), .A(n15477), 
        .B(n15433), .ZN(n15435) );
  NAND2_X1 U16591 ( .A1(n15436), .A2(n15435), .ZN(n15437) );
  AOI21_X1 U16592 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(n15471), .A(n15437), 
        .ZN(n15441) );
  OAI211_X1 U16593 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n15439), .A(n15473), 
        .B(n15438), .ZN(n15440) );
  OAI211_X1 U16594 ( .C1(n15466), .C2(n15442), .A(n15441), .B(n15440), .ZN(
        P2_U3229) );
  OAI211_X1 U16595 ( .C1(n15445), .C2(n15444), .A(n15477), .B(n15443), .ZN(
        n15446) );
  NAND2_X1 U16596 ( .A1(n15447), .A2(n15446), .ZN(n15448) );
  AOI21_X1 U16597 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(n15471), .A(n15448), 
        .ZN(n15453) );
  OAI211_X1 U16598 ( .C1(n15451), .C2(n15450), .A(n15473), .B(n15449), .ZN(
        n15452) );
  OAI211_X1 U16599 ( .C1(n15466), .C2(n15454), .A(n15453), .B(n15452), .ZN(
        P2_U3230) );
  OAI211_X1 U16600 ( .C1(n15457), .C2(n15456), .A(n15455), .B(n15477), .ZN(
        n15458) );
  NAND2_X1 U16601 ( .A1(n15459), .A2(n15458), .ZN(n15460) );
  AOI21_X1 U16602 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(n15471), .A(n15460), 
        .ZN(n15465) );
  OAI211_X1 U16603 ( .C1(n15463), .C2(n15462), .A(n15473), .B(n15461), .ZN(
        n15464) );
  OAI211_X1 U16604 ( .C1(n15467), .C2(n15466), .A(n15465), .B(n15464), .ZN(
        P2_U3231) );
  OAI21_X1 U16605 ( .B1(n15469), .B2(n15468), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15470) );
  OAI21_X1 U16606 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15470), .ZN(n15483) );
  NAND2_X1 U16607 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n15471), .ZN(n15482) );
  OAI211_X1 U16608 ( .C1(n15475), .C2(n15474), .A(n15473), .B(n15472), .ZN(
        n15481) );
  OAI211_X1 U16609 ( .C1(n15479), .C2(n15478), .A(n15477), .B(n15476), .ZN(
        n15480) );
  NAND4_X1 U16610 ( .A1(n15483), .A2(n15482), .A3(n15481), .A4(n15480), .ZN(
        P2_U3227) );
  INV_X1 U16611 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n15484) );
  NOR2_X1 U16612 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n15484), .ZN(n15490) );
  AOI21_X1 U16613 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n15484), .A(n15490), .ZN(
        n15486) );
  INV_X1 U16614 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15485) );
  NOR2_X1 U16615 ( .A1(n15486), .A2(n15485), .ZN(n15650) );
  AOI21_X1 U16616 ( .B1(n15486), .B2(n15485), .A(n15650), .ZN(SUB_1596_U53) );
  NAND2_X1 U16617 ( .A1(n15490), .A2(n15489), .ZN(n15487) );
  XNOR2_X1 U16618 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n15500), .ZN(n15495) );
  NAND2_X1 U16619 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n15491), .ZN(n15492) );
  XOR2_X1 U16620 ( .A(n15491), .B(P2_ADDR_REG_1__SCAN_IN), .Z(n15651) );
  NAND2_X1 U16621 ( .A1(n15495), .A2(n15494), .ZN(n15496) );
  OAI21_X1 U16622 ( .B1(n15495), .B2(n15494), .A(n15496), .ZN(n15493) );
  INV_X1 U16623 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n15497) );
  XOR2_X1 U16624 ( .A(n15493), .B(n15497), .Z(SUB_1596_U61) );
  NOR2_X1 U16625 ( .A1(n15495), .A2(n15494), .ZN(n15498) );
  NAND2_X1 U16626 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n15499), .ZN(n15501) );
  XNOR2_X1 U16627 ( .A(P3_ADDR_REG_3__SCAN_IN), .B(n15502), .ZN(n15503) );
  XNOR2_X1 U16628 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n15503), .ZN(n15506) );
  XNOR2_X1 U16629 ( .A(n15507), .B(n15506), .ZN(n15508) );
  XNOR2_X1 U16630 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15508), .ZN(SUB_1596_U60)
         );
  NAND2_X1 U16631 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n15502), .ZN(n15505) );
  NAND2_X1 U16632 ( .A1(n15505), .A2(n15504), .ZN(n15511) );
  XOR2_X1 U16633 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n15514), .Z(n15512) );
  XNOR2_X1 U16634 ( .A(n15511), .B(n15512), .ZN(n15516) );
  NOR2_X1 U16635 ( .A1(n15507), .A2(n15506), .ZN(n15510) );
  NOR2_X1 U16636 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(n15508), .ZN(n15509) );
  XOR2_X1 U16637 ( .A(n15518), .B(n15517), .Z(SUB_1596_U59) );
  XOR2_X1 U16638 ( .A(P3_ADDR_REG_5__SCAN_IN), .B(n15527), .Z(n15515) );
  NAND2_X1 U16639 ( .A1(n15512), .A2(n15511), .ZN(n15513) );
  XNOR2_X1 U16640 ( .A(n15515), .B(n15525), .ZN(n15521) );
  NAND2_X1 U16641 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n15516), .ZN(n15519) );
  XOR2_X1 U16642 ( .A(n15522), .B(P2_ADDR_REG_5__SCAN_IN), .Z(SUB_1596_U58) );
  NAND2_X1 U16643 ( .A1(n15521), .A2(n15520), .ZN(n15524) );
  NAND2_X1 U16644 ( .A1(n15522), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n15523) );
  NAND2_X1 U16645 ( .A1(n15524), .A2(n15523), .ZN(n15647) );
  XOR2_X1 U16646 ( .A(n15532), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n15528) );
  AND2_X1 U16647 ( .A1(n15527), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n15526) );
  XOR2_X1 U16648 ( .A(n15528), .B(n15530), .Z(n15646) );
  NOR2_X1 U16649 ( .A1(n15647), .A2(n15646), .ZN(n15529) );
  INV_X1 U16650 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n15648) );
  NAND2_X1 U16651 ( .A1(n15647), .A2(n15646), .ZN(n15645) );
  XNOR2_X1 U16652 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n15534), .ZN(n15535) );
  XNOR2_X1 U16653 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n15535), .ZN(n15539) );
  XNOR2_X1 U16654 ( .A(n15540), .B(n15539), .ZN(SUB_1596_U56) );
  XNOR2_X1 U16655 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(n15533), .ZN(n15548) );
  NAND2_X1 U16656 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n15534), .ZN(n15537) );
  XOR2_X1 U16657 ( .A(n15548), .B(n15547), .Z(n15542) );
  NOR2_X1 U16658 ( .A1(n15542), .A2(n15541), .ZN(n15546) );
  NOR2_X1 U16659 ( .A1(n15546), .A2(n15544), .ZN(n15543) );
  XOR2_X1 U16660 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n15543), .Z(SUB_1596_U55) );
  NOR2_X1 U16661 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n15544), .ZN(n15545) );
  INV_X1 U16662 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15550) );
  XNOR2_X1 U16663 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(n15551), .ZN(n15553) );
  XOR2_X1 U16664 ( .A(n15554), .B(n15553), .Z(n15556) );
  NAND2_X1 U16665 ( .A1(n15557), .A2(n15556), .ZN(n15558) );
  OAI21_X1 U16666 ( .B1(n15557), .B2(n15556), .A(n15558), .ZN(n15552) );
  XOR2_X1 U16667 ( .A(n15552), .B(n15559), .Z(SUB_1596_U54) );
  INV_X1 U16668 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n15692) );
  AOI21_X2 U16669 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n15692), .A(n15555), .ZN(
        n15562) );
  XOR2_X1 U16670 ( .A(n15564), .B(P1_ADDR_REG_10__SCAN_IN), .Z(n15561) );
  XNOR2_X1 U16671 ( .A(n15562), .B(n15561), .ZN(n15565) );
  AOI21_X1 U16672 ( .B1(n15565), .B2(n15566), .A(n15567), .ZN(n15560) );
  XOR2_X1 U16673 ( .A(n15560), .B(P2_ADDR_REG_10__SCAN_IN), .Z(SUB_1596_U70)
         );
  XOR2_X1 U16674 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n15575) );
  NAND2_X1 U16675 ( .A1(n15562), .A2(n15561), .ZN(n15563) );
  XOR2_X1 U16676 ( .A(n15575), .B(n15574), .Z(n15569) );
  NOR2_X1 U16677 ( .A1(n15573), .A2(n15571), .ZN(n15570) );
  XOR2_X1 U16678 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n15570), .Z(SUB_1596_U69)
         );
  NOR2_X1 U16679 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n15571), .ZN(n15572) );
  INV_X1 U16680 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n15700) );
  XOR2_X1 U16681 ( .A(n15585), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n15582) );
  XNOR2_X1 U16682 ( .A(n15583), .B(n15582), .ZN(n15577) );
  XNOR2_X1 U16683 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n15579), .ZN(SUB_1596_U68)
         );
  NOR2_X1 U16684 ( .A1(n15578), .A2(n15577), .ZN(n15581) );
  NOR2_X1 U16685 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n15579), .ZN(n15580) );
  INV_X1 U16686 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15730) );
  XOR2_X1 U16687 ( .A(n15730), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n15586) );
  NAND2_X1 U16688 ( .A1(n15583), .A2(n15582), .ZN(n15584) );
  XNOR2_X1 U16689 ( .A(n15586), .B(n15593), .ZN(n15588) );
  NAND2_X1 U16690 ( .A1(n15589), .A2(n15588), .ZN(n15590) );
  OAI21_X1 U16691 ( .B1(n15589), .B2(n15588), .A(n15590), .ZN(n15587) );
  INV_X1 U16692 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15591) );
  XOR2_X1 U16693 ( .A(n15587), .B(n15591), .Z(SUB_1596_U67) );
  NAND2_X1 U16694 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n15730), .ZN(n15592) );
  INV_X1 U16695 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15599) );
  XNOR2_X1 U16696 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(n15599), .ZN(n15596) );
  XNOR2_X1 U16697 ( .A(n15597), .B(n15596), .ZN(n15601) );
  NOR2_X1 U16698 ( .A1(n15601), .A2(n15600), .ZN(n15602) );
  AOI21_X1 U16699 ( .B1(n15600), .B2(n15601), .A(n15602), .ZN(n15595) );
  XOR2_X1 U16700 ( .A(n15595), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  NOR2_X1 U16701 ( .A1(n15597), .A2(n15596), .ZN(n15598) );
  AOI21_X1 U16702 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n15599), .A(n15598), 
        .ZN(n15607) );
  INV_X1 U16703 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15609) );
  XOR2_X1 U16704 ( .A(P3_ADDR_REG_15__SCAN_IN), .B(n15609), .Z(n15606) );
  XOR2_X1 U16705 ( .A(n15607), .B(n15606), .Z(n15610) );
  INV_X1 U16706 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15604) );
  NAND2_X1 U16707 ( .A1(n15601), .A2(n15600), .ZN(n15603) );
  NOR2_X1 U16708 ( .A1(n15611), .A2(n15610), .ZN(n15612) );
  AOI21_X1 U16709 ( .B1(n15610), .B2(n15611), .A(n15612), .ZN(n15605) );
  XOR2_X1 U16710 ( .A(n15605), .B(P2_ADDR_REG_15__SCAN_IN), .Z(SUB_1596_U65)
         );
  NAND2_X1 U16711 ( .A1(n15607), .A2(n15606), .ZN(n15608) );
  XOR2_X1 U16712 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n15616), .Z(n15617) );
  XNOR2_X1 U16713 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n15617), .ZN(n15620) );
  INV_X1 U16714 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15614) );
  NAND2_X1 U16715 ( .A1(n15611), .A2(n15610), .ZN(n15613) );
  NAND2_X1 U16716 ( .A1(n15621), .A2(n15620), .ZN(n15622) );
  OAI21_X1 U16717 ( .B1(n15620), .B2(n15621), .A(n15622), .ZN(n15615) );
  INV_X1 U16718 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15623) );
  XOR2_X1 U16719 ( .A(n15615), .B(n15623), .Z(SUB_1596_U64) );
  INV_X1 U16720 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n15807) );
  NOR2_X1 U16721 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n15616), .ZN(n15619) );
  XOR2_X1 U16722 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n15629), .Z(n15630) );
  XOR2_X1 U16723 ( .A(n15807), .B(n15630), .Z(n15625) );
  XOR2_X1 U16724 ( .A(n15625), .B(P2_ADDR_REG_17__SCAN_IN), .Z(n15627) );
  NOR2_X1 U16725 ( .A1(n15621), .A2(n15620), .ZN(n15624) );
  XOR2_X1 U16726 ( .A(n15627), .B(n15626), .Z(SUB_1596_U63) );
  NAND2_X1 U16727 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n15625), .ZN(n15628) );
  NOR2_X1 U16728 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n15629), .ZN(n15632) );
  AND2_X1 U16729 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n15630), .ZN(n15631) );
  NAND2_X1 U16730 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n15637), .ZN(n15633) );
  OAI21_X1 U16731 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n15637), .A(n15633), 
        .ZN(n15635) );
  XOR2_X1 U16732 ( .A(n15634), .B(n15635), .Z(n15639) );
  XOR2_X1 U16733 ( .A(n15640), .B(P2_ADDR_REG_18__SCAN_IN), .Z(SUB_1596_U62)
         );
  NOR2_X1 U16734 ( .A1(n15635), .A2(n15634), .ZN(n15636) );
  AOI21_X1 U16735 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n15637), .A(n15636), 
        .ZN(n15644) );
  NAND2_X1 U16736 ( .A1(n15639), .A2(n15638), .ZN(n15642) );
  NAND2_X1 U16737 ( .A1(n15640), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n15641) );
  XNOR2_X1 U16738 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n15643) );
  OAI21_X1 U16739 ( .B1(n15647), .B2(n15646), .A(n15645), .ZN(n15649) );
  XOR2_X1 U16740 ( .A(n15649), .B(n15648), .Z(SUB_1596_U57) );
  XOR2_X1 U16741 ( .A(n15651), .B(n15650), .Z(SUB_1596_U5) );
  NOR2_X1 U16742 ( .A1(n15652), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15654) );
  NAND3_X1 U16743 ( .A1(n15825), .A2(n15822), .A3(n15811), .ZN(n15653) );
  OAI21_X1 U16744 ( .B1(n15655), .B2(n15654), .A(n15653), .ZN(n15657) );
  AOI22_X1 U16745 ( .A1(n15817), .A2(P3_IR_REG_0__SCAN_IN), .B1(n15771), .B2(
        P3_ADDR_REG_0__SCAN_IN), .ZN(n15656) );
  OAI211_X1 U16746 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n15658), .A(n15657), .B(
        n15656), .ZN(P3_U3182) );
  AOI21_X1 U16747 ( .B1(n10760), .B2(n15660), .A(n15659), .ZN(n15664) );
  AOI21_X1 U16748 ( .B1(n10761), .B2(n15662), .A(n15661), .ZN(n15663) );
  OAI22_X1 U16749 ( .A1(n15664), .A2(n15822), .B1(n15663), .B2(n15825), .ZN(
        n15665) );
  AOI211_X1 U16750 ( .C1(P3_ADDR_REG_7__SCAN_IN), .C2(n15771), .A(n15666), .B(
        n15665), .ZN(n15674) );
  NAND2_X1 U16751 ( .A1(n15668), .A2(n15667), .ZN(n15669) );
  AOI21_X1 U16752 ( .B1(n15670), .B2(n15669), .A(n15811), .ZN(n15671) );
  AOI21_X1 U16753 ( .B1(n15817), .B2(n15672), .A(n15671), .ZN(n15673) );
  NAND2_X1 U16754 ( .A1(n15674), .A2(n15673), .ZN(P3_U3189) );
  AOI21_X1 U16755 ( .B1(n11319), .B2(n15676), .A(n15675), .ZN(n15677) );
  OR2_X1 U16756 ( .A1(n15677), .A2(n15822), .ZN(n15689) );
  AOI21_X1 U16757 ( .B1(n11320), .B2(n15679), .A(n15678), .ZN(n15680) );
  OR2_X1 U16758 ( .A1(n15680), .A2(n15825), .ZN(n15688) );
  NAND2_X1 U16759 ( .A1(n15682), .A2(n15681), .ZN(n15683) );
  NAND3_X1 U16760 ( .A1(n15684), .A2(n15775), .A3(n15683), .ZN(n15687) );
  NAND2_X1 U16761 ( .A1(n15817), .A2(n15685), .ZN(n15686) );
  OAI211_X1 U16762 ( .C1(n15692), .C2(n15808), .A(n15691), .B(n15690), .ZN(
        P3_U3191) );
  AOI21_X1 U16763 ( .B1(n11863), .B2(n15694), .A(n15693), .ZN(n15708) );
  XNOR2_X1 U16764 ( .A(n15696), .B(n15695), .ZN(n15702) );
  NAND2_X1 U16765 ( .A1(n15817), .A2(n15697), .ZN(n15699) );
  OAI211_X1 U16766 ( .C1(n15700), .C2(n15808), .A(n15699), .B(n15698), .ZN(
        n15701) );
  AOI21_X1 U16767 ( .B1(n15702), .B2(n15775), .A(n15701), .ZN(n15707) );
  AOI21_X1 U16768 ( .B1(n15704), .B2(n8487), .A(n15703), .ZN(n15705) );
  OR2_X1 U16769 ( .A1(n15822), .A2(n15705), .ZN(n15706) );
  OAI211_X1 U16770 ( .C1(n15708), .C2(n15825), .A(n15707), .B(n15706), .ZN(
        P3_U3193) );
  AOI21_X1 U16771 ( .B1(n15710), .B2(n15709), .A(n7223), .ZN(n15725) );
  INV_X1 U16772 ( .A(n15711), .ZN(n15718) );
  OAI21_X1 U16773 ( .B1(n15808), .B2(n15585), .A(n15712), .ZN(n15717) );
  INV_X1 U16774 ( .A(n15733), .ZN(n15713) );
  AOI211_X1 U16775 ( .C1(n15715), .C2(n15714), .A(n15811), .B(n15713), .ZN(
        n15716) );
  AOI211_X1 U16776 ( .C1(n15817), .C2(n15718), .A(n15717), .B(n15716), .ZN(
        n15724) );
  AOI21_X1 U16777 ( .B1(n15721), .B2(n15720), .A(n15719), .ZN(n15722) );
  OR2_X1 U16778 ( .A1(n15722), .A2(n15822), .ZN(n15723) );
  OAI211_X1 U16779 ( .C1(n15725), .C2(n15825), .A(n15724), .B(n15723), .ZN(
        P3_U3194) );
  AOI21_X1 U16780 ( .B1(n8327), .B2(n15727), .A(n15726), .ZN(n15745) );
  INV_X1 U16781 ( .A(n15728), .ZN(n15729) );
  OAI21_X1 U16782 ( .B1(n15808), .B2(n15730), .A(n15729), .ZN(n15738) );
  AOI21_X1 U16783 ( .B1(n15733), .B2(n15732), .A(n15731), .ZN(n15734) );
  INV_X1 U16784 ( .A(n15734), .ZN(n15736) );
  AOI21_X1 U16785 ( .B1(n15736), .B2(n15735), .A(n15811), .ZN(n15737) );
  AOI211_X1 U16786 ( .C1(n15817), .C2(n15739), .A(n15738), .B(n15737), .ZN(
        n15744) );
  AOI21_X1 U16787 ( .B1(n15741), .B2(n8325), .A(n15740), .ZN(n15742) );
  OR2_X1 U16788 ( .A1(n15822), .A2(n15742), .ZN(n15743) );
  OAI211_X1 U16789 ( .C1(n15745), .C2(n15825), .A(n15744), .B(n15743), .ZN(
        P3_U3195) );
  AOI21_X1 U16790 ( .B1(n15748), .B2(n15747), .A(n15746), .ZN(n15764) );
  INV_X1 U16791 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15750) );
  OAI21_X1 U16792 ( .B1(n15808), .B2(n15750), .A(n15749), .ZN(n15756) );
  OAI211_X1 U16793 ( .C1(n15753), .C2(n15752), .A(n15751), .B(n15775), .ZN(
        n15754) );
  INV_X1 U16794 ( .A(n15754), .ZN(n15755) );
  AOI211_X1 U16795 ( .C1(n15817), .C2(n15757), .A(n15756), .B(n15755), .ZN(
        n15763) );
  AOI21_X1 U16796 ( .B1(n15760), .B2(n15759), .A(n15758), .ZN(n15761) );
  OR2_X1 U16797 ( .A1(n15761), .A2(n15822), .ZN(n15762) );
  OAI211_X1 U16798 ( .C1(n15764), .C2(n15825), .A(n15763), .B(n15762), .ZN(
        P3_U3196) );
  AOI21_X1 U16799 ( .B1(n15767), .B2(n15766), .A(n15765), .ZN(n15783) );
  XOR2_X1 U16800 ( .A(n15769), .B(n15768), .Z(n15776) );
  AOI21_X1 U16801 ( .B1(n15771), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n15770), 
        .ZN(n15772) );
  OAI21_X1 U16802 ( .B1(n15773), .B2(n16152), .A(n15772), .ZN(n15774) );
  AOI21_X1 U16803 ( .B1(n15776), .B2(n15775), .A(n15774), .ZN(n15782) );
  AOI21_X1 U16804 ( .B1(n15779), .B2(n15778), .A(n15777), .ZN(n15780) );
  OR2_X1 U16805 ( .A1(n15822), .A2(n15780), .ZN(n15781) );
  OAI211_X1 U16806 ( .C1(n15783), .C2(n15825), .A(n15782), .B(n15781), .ZN(
        P3_U3197) );
  AOI21_X1 U16807 ( .B1(n15786), .B2(n15785), .A(n15784), .ZN(n15801) );
  INV_X1 U16808 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n15788) );
  OAI21_X1 U16809 ( .B1(n15808), .B2(n15788), .A(n15787), .ZN(n15794) );
  NAND2_X1 U16810 ( .A1(n15790), .A2(n15789), .ZN(n15791) );
  AOI21_X1 U16811 ( .B1(n15792), .B2(n15791), .A(n15811), .ZN(n15793) );
  AOI211_X1 U16812 ( .C1(n15817), .C2(n15795), .A(n15794), .B(n15793), .ZN(
        n15800) );
  AOI21_X1 U16813 ( .B1(n15797), .B2(n15796), .A(n7239), .ZN(n15798) );
  OR2_X1 U16814 ( .A1(n15798), .A2(n15822), .ZN(n15799) );
  OAI211_X1 U16815 ( .C1(n15801), .C2(n15825), .A(n15800), .B(n15799), .ZN(
        P3_U3198) );
  AOI21_X1 U16816 ( .B1(n15804), .B2(n15803), .A(n15802), .ZN(n15826) );
  INV_X1 U16817 ( .A(n15805), .ZN(n15806) );
  OAI21_X1 U16818 ( .B1(n15808), .B2(n15807), .A(n15806), .ZN(n15815) );
  INV_X1 U16819 ( .A(n15809), .ZN(n15810) );
  AOI211_X1 U16820 ( .C1(n15813), .C2(n15812), .A(n15811), .B(n15810), .ZN(
        n15814) );
  AOI211_X1 U16821 ( .C1(n15817), .C2(n15816), .A(n15815), .B(n15814), .ZN(
        n15824) );
  AOI21_X1 U16822 ( .B1(n15820), .B2(n15819), .A(n15818), .ZN(n15821) );
  OR2_X1 U16823 ( .A1(n15822), .A2(n15821), .ZN(n15823) );
  OAI211_X1 U16824 ( .C1(n15826), .C2(n15825), .A(n15824), .B(n15823), .ZN(
        P3_U3199) );
  INV_X1 U16825 ( .A(P1_RD_REG_SCAN_IN), .ZN(n15828) );
  OAI221_X1 U16826 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(
        n15829), .C2(n7622), .A(n15827), .ZN(U29) );
  INV_X1 U16827 ( .A(n15833), .ZN(n15842) );
  OAI21_X1 U16828 ( .B1(n16034), .B2(n15955), .A(n15842), .ZN(n15831) );
  AND2_X1 U16829 ( .A1(n15831), .A2(n15830), .ZN(n15845) );
  INV_X1 U16830 ( .A(n15845), .ZN(n15835) );
  OAI22_X1 U16831 ( .A1(n15833), .A2(n15856), .B1(n15839), .B2(n15832), .ZN(
        n15834) );
  NOR2_X1 U16832 ( .A1(n15835), .A2(n15834), .ZN(n15838) );
  AOI22_X1 U16833 ( .A1(n16067), .A2(n15838), .B1(n15836), .B2(n16066), .ZN(
        P1_U3528) );
  INV_X1 U16834 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15837) );
  AOI22_X1 U16835 ( .A1(n16071), .A2(n15838), .B1(n15837), .B2(n16068), .ZN(
        P1_U3459) );
  AOI22_X1 U16836 ( .A1(n16037), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n16047), 
        .B2(P1_REG2_REG_0__SCAN_IN), .ZN(n15844) );
  AOI21_X1 U16837 ( .B1(n16041), .B2(n15840), .A(n15839), .ZN(n15841) );
  AOI21_X1 U16838 ( .B1(n16044), .B2(n15842), .A(n15841), .ZN(n15843) );
  OAI211_X1 U16839 ( .C1(n16047), .C2(n15845), .A(n15844), .B(n15843), .ZN(
        P1_U3293) );
  OAI211_X1 U16840 ( .C1(n15848), .C2(n16106), .A(n15847), .B(n15846), .ZN(
        n15849) );
  INV_X1 U16841 ( .A(n15849), .ZN(n15851) );
  AOI22_X1 U16842 ( .A1(n16142), .A2(n15851), .B1(n15850), .B2(n16141), .ZN(
        P2_U3499) );
  AOI22_X1 U16843 ( .A1(n16146), .A2(n15851), .B1(n9621), .B2(n16143), .ZN(
        P2_U3430) );
  OAI211_X1 U16844 ( .C1(n15854), .C2(n16058), .A(n15853), .B(n15852), .ZN(
        n15858) );
  AOI21_X1 U16845 ( .B1(n15977), .B2(n15856), .A(n15855), .ZN(n15857) );
  NOR2_X1 U16846 ( .A1(n15858), .A2(n15857), .ZN(n15861) );
  AOI22_X1 U16847 ( .A1(n16067), .A2(n15861), .B1(n15859), .B2(n16066), .ZN(
        P1_U3529) );
  INV_X1 U16848 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15860) );
  AOI22_X1 U16849 ( .A1(n16071), .A2(n15861), .B1(n15860), .B2(n16068), .ZN(
        P1_U3462) );
  INV_X1 U16850 ( .A(n15862), .ZN(n15863) );
  AOI21_X1 U16851 ( .B1(n16107), .B2(n16106), .A(n15863), .ZN(n15868) );
  NOR2_X1 U16852 ( .A1(n15864), .A2(n16136), .ZN(n15866) );
  NOR4_X1 U16853 ( .A1(n15868), .A2(n15867), .A3(n15866), .A4(n15865), .ZN(
        n15869) );
  AOI22_X1 U16854 ( .A1(n16142), .A2(n15869), .B1(n9450), .B2(n16141), .ZN(
        P2_U3500) );
  AOI22_X1 U16855 ( .A1(n16146), .A2(n15869), .B1(n9579), .B2(n16143), .ZN(
        P2_U3433) );
  XNOR2_X1 U16856 ( .A(n15871), .B(n15870), .ZN(n15887) );
  INV_X1 U16857 ( .A(n15887), .ZN(n15897) );
  NOR2_X1 U16858 ( .A1(n15872), .A2(n16096), .ZN(n15890) );
  AOI22_X1 U16859 ( .A1(n15876), .A2(n15875), .B1(n15874), .B2(n15873), .ZN(
        n15885) );
  INV_X1 U16860 ( .A(n15877), .ZN(n15883) );
  AND3_X1 U16861 ( .A1(n15880), .A2(n15879), .A3(n15878), .ZN(n15882) );
  OAI21_X1 U16862 ( .B1(n15883), .B2(n15882), .A(n15881), .ZN(n15884) );
  OAI211_X1 U16863 ( .C1(n15887), .C2(n15886), .A(n15885), .B(n15884), .ZN(
        n15895) );
  AOI211_X1 U16864 ( .C1(n15897), .C2(n16082), .A(n15890), .B(n15895), .ZN(
        n15889) );
  AOI22_X1 U16865 ( .A1(n16101), .A2(n15889), .B1(n9825), .B2(n16155), .ZN(
        P3_U3461) );
  INV_X1 U16866 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15888) );
  AOI22_X1 U16867 ( .A1(n16104), .A2(n15889), .B1(n15888), .B2(n16160), .ZN(
        P3_U3396) );
  INV_X1 U16868 ( .A(n15890), .ZN(n15894) );
  OAI22_X1 U16869 ( .A1(n15894), .A2(n15893), .B1(n15892), .B2(n15891), .ZN(
        n15896) );
  AOI211_X1 U16870 ( .C1(n15898), .C2(n15897), .A(n15896), .B(n15895), .ZN(
        n15900) );
  AOI22_X1 U16871 ( .A1(n13853), .A2(n9826), .B1(n15900), .B2(n15899), .ZN(
        P3_U3231) );
  INV_X1 U16872 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n15901) );
  AOI22_X1 U16873 ( .A1(n16071), .A2(n15902), .B1(n15901), .B2(n16068), .ZN(
        P1_U3465) );
  AOI21_X1 U16874 ( .B1(n15905), .B2(n15904), .A(n15903), .ZN(n15910) );
  OAI21_X1 U16875 ( .B1(n15907), .B2(n16092), .A(n15906), .ZN(n15908) );
  AND3_X1 U16876 ( .A1(n15910), .A2(n15909), .A3(n15908), .ZN(n15911) );
  AOI22_X1 U16877 ( .A1(n16142), .A2(n15911), .B1(n9449), .B2(n16141), .ZN(
        P2_U3501) );
  AOI22_X1 U16878 ( .A1(n16146), .A2(n15911), .B1(n9601), .B2(n16143), .ZN(
        P2_U3436) );
  OAI22_X1 U16879 ( .A1(n15913), .A2(n16097), .B1(n16096), .B2(n15912), .ZN(
        n15914) );
  NOR2_X1 U16880 ( .A1(n15915), .A2(n15914), .ZN(n15917) );
  AOI22_X1 U16881 ( .A1(n16101), .A2(n15917), .B1(n9832), .B2(n16155), .ZN(
        P3_U3462) );
  INV_X1 U16882 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15916) );
  AOI22_X1 U16883 ( .A1(n16104), .A2(n15917), .B1(n15916), .B2(n16160), .ZN(
        P3_U3399) );
  NAND2_X1 U16884 ( .A1(n15918), .A2(n15948), .ZN(n15930) );
  INV_X1 U16885 ( .A(n15930), .ZN(n15920) );
  AOI21_X1 U16886 ( .B1(n15921), .B2(n15920), .A(n15919), .ZN(n15929) );
  AOI211_X1 U16887 ( .C1(n15924), .C2(n15923), .A(n16123), .B(n15922), .ZN(
        n15925) );
  AOI21_X1 U16888 ( .B1(n15927), .B2(n15926), .A(n15925), .ZN(n15928) );
  OAI211_X1 U16889 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n16133), .A(n15929), .B(
        n15928), .ZN(P1_U3218) );
  NAND3_X1 U16890 ( .A1(n15932), .A2(n15931), .A3(n15930), .ZN(n15936) );
  NOR2_X1 U16891 ( .A1(n15934), .A2(n15933), .ZN(n15935) );
  AOI211_X1 U16892 ( .C1(n15955), .C2(n15937), .A(n15936), .B(n15935), .ZN(
        n15939) );
  AOI22_X1 U16893 ( .A1(n16067), .A2(n15939), .B1(n9158), .B2(n16066), .ZN(
        P1_U3531) );
  INV_X1 U16894 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n15938) );
  AOI22_X1 U16895 ( .A1(n16071), .A2(n15939), .B1(n15938), .B2(n16068), .ZN(
        P1_U3468) );
  INV_X1 U16896 ( .A(n15940), .ZN(n15941) );
  AOI21_X1 U16897 ( .B1(n16107), .B2(n16106), .A(n15941), .ZN(n15946) );
  OAI211_X1 U16898 ( .C1(n15944), .C2(n16136), .A(n15943), .B(n15942), .ZN(
        n15945) );
  NOR2_X1 U16899 ( .A1(n15946), .A2(n15945), .ZN(n15947) );
  AOI22_X1 U16900 ( .A1(n16142), .A2(n15947), .B1(n9455), .B2(n16141), .ZN(
        P2_U3502) );
  AOI22_X1 U16901 ( .A1(n16146), .A2(n15947), .B1(n9586), .B2(n16143), .ZN(
        P2_U3439) );
  NAND2_X1 U16902 ( .A1(n15949), .A2(n15948), .ZN(n15950) );
  OAI211_X1 U16903 ( .C1(n15953), .C2(n15952), .A(n15951), .B(n15950), .ZN(
        n15958) );
  AND3_X1 U16904 ( .A1(n15956), .A2(n15955), .A3(n15954), .ZN(n15957) );
  AOI211_X1 U16905 ( .C1(n15959), .C2(n16064), .A(n15958), .B(n15957), .ZN(
        n15962) );
  AOI22_X1 U16906 ( .A1(n16067), .A2(n15962), .B1(n15960), .B2(n16066), .ZN(
        P1_U3532) );
  INV_X1 U16907 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n15961) );
  AOI22_X1 U16908 ( .A1(n16071), .A2(n15962), .B1(n15961), .B2(n16068), .ZN(
        P1_U3471) );
  INV_X1 U16909 ( .A(n15963), .ZN(n15965) );
  OAI211_X1 U16910 ( .C1(n15966), .C2(n16136), .A(n15965), .B(n15964), .ZN(
        n15969) );
  AOI21_X1 U16911 ( .B1(n16107), .B2(n16106), .A(n15967), .ZN(n15968) );
  NOR2_X1 U16912 ( .A1(n15969), .A2(n15968), .ZN(n15971) );
  AOI22_X1 U16913 ( .A1(n16142), .A2(n15971), .B1(n9456), .B2(n16141), .ZN(
        P2_U3503) );
  INV_X1 U16914 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15970) );
  AOI22_X1 U16915 ( .A1(n16146), .A2(n15971), .B1(n15970), .B2(n16143), .ZN(
        P2_U3442) );
  INV_X1 U16916 ( .A(n15976), .ZN(n15979) );
  NOR3_X1 U16917 ( .A1(n15974), .A2(n15973), .A3(n15972), .ZN(n15975) );
  OAI21_X1 U16918 ( .B1(n15977), .B2(n15976), .A(n15975), .ZN(n15978) );
  AOI21_X1 U16919 ( .B1(n16017), .B2(n15979), .A(n15978), .ZN(n15982) );
  AOI22_X1 U16920 ( .A1(n16067), .A2(n15982), .B1(n15980), .B2(n16066), .ZN(
        P1_U3533) );
  INV_X1 U16921 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15981) );
  AOI22_X1 U16922 ( .A1(n16071), .A2(n15982), .B1(n15981), .B2(n16068), .ZN(
        P1_U3474) );
  NOR2_X1 U16923 ( .A1(n15983), .A2(n16096), .ZN(n15985) );
  AOI211_X1 U16924 ( .C1(n15986), .C2(n16082), .A(n15985), .B(n15984), .ZN(
        n15988) );
  AOI22_X1 U16925 ( .A1(n16101), .A2(n15988), .B1(n10178), .B2(n16155), .ZN(
        P3_U3465) );
  INV_X1 U16926 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15987) );
  AOI22_X1 U16927 ( .A1(n16104), .A2(n15988), .B1(n15987), .B2(n16160), .ZN(
        P3_U3408) );
  AOI222_X1 U16928 ( .A1(n15991), .A2(n15990), .B1(P1_REG2_REG_6__SCAN_IN), 
        .B2(n15998), .C1(n16037), .C2(n15989), .ZN(n15996) );
  INV_X1 U16929 ( .A(n15992), .ZN(n15994) );
  AOI22_X1 U16930 ( .A1(n15994), .A2(n16044), .B1(n16035), .B2(n15993), .ZN(
        n15995) );
  OAI211_X1 U16931 ( .C1(n15998), .C2(n15997), .A(n15996), .B(n15995), .ZN(
        P1_U3287) );
  OAI22_X1 U16932 ( .A1(n16000), .A2(n16097), .B1(n16096), .B2(n15999), .ZN(
        n16001) );
  NOR2_X1 U16933 ( .A1(n16002), .A2(n16001), .ZN(n16004) );
  AOI22_X1 U16934 ( .A1(n16101), .A2(n16004), .B1(n10760), .B2(n16155), .ZN(
        P3_U3466) );
  INV_X1 U16935 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n16003) );
  AOI22_X1 U16936 ( .A1(n16104), .A2(n16004), .B1(n16003), .B2(n16160), .ZN(
        P3_U3411) );
  OAI22_X1 U16937 ( .A1(n16006), .A2(n16097), .B1(n16005), .B2(n16096), .ZN(
        n16007) );
  NOR2_X1 U16938 ( .A1(n16008), .A2(n16007), .ZN(n16010) );
  AOI22_X1 U16939 ( .A1(n16101), .A2(n16010), .B1(n8471), .B2(n16155), .ZN(
        P3_U3467) );
  INV_X1 U16940 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n16009) );
  AOI22_X1 U16941 ( .A1(n16104), .A2(n16010), .B1(n16009), .B2(n16160), .ZN(
        P3_U3414) );
  INV_X1 U16942 ( .A(n16011), .ZN(n16016) );
  INV_X1 U16943 ( .A(n16012), .ZN(n16013) );
  OAI21_X1 U16944 ( .B1(n7593), .B2(n16058), .A(n16013), .ZN(n16015) );
  AOI211_X1 U16945 ( .C1(n16017), .C2(n16016), .A(n16015), .B(n16014), .ZN(
        n16020) );
  AOI22_X1 U16946 ( .A1(n16067), .A2(n16020), .B1(n16018), .B2(n16066), .ZN(
        P1_U3536) );
  INV_X1 U16947 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n16019) );
  AOI22_X1 U16948 ( .A1(n16071), .A2(n16020), .B1(n16019), .B2(n16068), .ZN(
        P1_U3483) );
  OAI21_X1 U16949 ( .B1(n7681), .B2(n16136), .A(n16021), .ZN(n16022) );
  AOI211_X1 U16950 ( .C1(n16024), .C2(n16140), .A(n16023), .B(n16022), .ZN(
        n16025) );
  AOI22_X1 U16951 ( .A1(n16142), .A2(n16025), .B1(n9467), .B2(n16141), .ZN(
        P2_U3507) );
  AOI22_X1 U16952 ( .A1(n16146), .A2(n16025), .B1(n10348), .B2(n16143), .ZN(
        P2_U3454) );
  OAI22_X1 U16953 ( .A1(n16027), .A2(n16097), .B1(n16096), .B2(n16026), .ZN(
        n16028) );
  NOR2_X1 U16954 ( .A1(n16029), .A2(n16028), .ZN(n16031) );
  AOI22_X1 U16955 ( .A1(n16101), .A2(n16031), .B1(n11319), .B2(n16155), .ZN(
        P3_U3468) );
  INV_X1 U16956 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n16030) );
  AOI22_X1 U16957 ( .A1(n16104), .A2(n16031), .B1(n16030), .B2(n16160), .ZN(
        P3_U3417) );
  INV_X1 U16958 ( .A(n16032), .ZN(n16033) );
  AOI21_X1 U16959 ( .B1(n16034), .B2(n16043), .A(n16033), .ZN(n16046) );
  NAND2_X1 U16960 ( .A1(n16036), .A2(n16035), .ZN(n16040) );
  AOI22_X1 U16961 ( .A1(n16047), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n16038), 
        .B2(n16037), .ZN(n16039) );
  OAI211_X1 U16962 ( .C1(n7591), .C2(n16041), .A(n16040), .B(n16039), .ZN(
        n16042) );
  AOI21_X1 U16963 ( .B1(n16044), .B2(n16043), .A(n16042), .ZN(n16045) );
  OAI21_X1 U16964 ( .B1(n16047), .B2(n16046), .A(n16045), .ZN(P1_U3284) );
  INV_X1 U16965 ( .A(n16048), .ZN(n16053) );
  OAI21_X1 U16966 ( .B1(n16050), .B2(n16136), .A(n16049), .ZN(n16052) );
  AOI211_X1 U16967 ( .C1(n16092), .C2(n16053), .A(n16052), .B(n16051), .ZN(
        n16055) );
  AOI22_X1 U16968 ( .A1(n16142), .A2(n16055), .B1(n16054), .B2(n16141), .ZN(
        P2_U3509) );
  AOI22_X1 U16969 ( .A1(n16146), .A2(n16055), .B1(n10568), .B2(n16143), .ZN(
        P2_U3460) );
  OAI211_X1 U16970 ( .C1(n16059), .C2(n16058), .A(n16057), .B(n16056), .ZN(
        n16063) );
  NOR2_X1 U16971 ( .A1(n16061), .A2(n16060), .ZN(n16062) );
  AOI211_X1 U16972 ( .C1(n16065), .C2(n16064), .A(n16063), .B(n16062), .ZN(
        n16070) );
  AOI22_X1 U16973 ( .A1(n16067), .A2(n16070), .B1(n9400), .B2(n16066), .ZN(
        P1_U3539) );
  INV_X1 U16974 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n16069) );
  AOI22_X1 U16975 ( .A1(n16071), .A2(n16070), .B1(n16069), .B2(n16068), .ZN(
        P1_U3492) );
  OAI21_X1 U16976 ( .B1(n16073), .B2(n16136), .A(n16072), .ZN(n16075) );
  AOI211_X1 U16977 ( .C1(n16092), .C2(n16076), .A(n16075), .B(n16074), .ZN(
        n16077) );
  AOI22_X1 U16978 ( .A1(n16142), .A2(n16077), .B1(n9531), .B2(n16141), .ZN(
        P2_U3510) );
  AOI22_X1 U16979 ( .A1(n16146), .A2(n16077), .B1(n10699), .B2(n16143), .ZN(
        P2_U3463) );
  NOR2_X1 U16980 ( .A1(n16078), .A2(n16096), .ZN(n16080) );
  AOI211_X1 U16981 ( .C1(n16082), .C2(n16081), .A(n16080), .B(n16079), .ZN(
        n16085) );
  AOI22_X1 U16982 ( .A1(n16101), .A2(n16085), .B1(n16083), .B2(n16155), .ZN(
        P3_U3471) );
  INV_X1 U16983 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n16084) );
  AOI22_X1 U16984 ( .A1(n16104), .A2(n16085), .B1(n16084), .B2(n16160), .ZN(
        P3_U3426) );
  INV_X1 U16985 ( .A(n16086), .ZN(n16091) );
  OAI21_X1 U16986 ( .B1(n16088), .B2(n16136), .A(n16087), .ZN(n16090) );
  AOI211_X1 U16987 ( .C1(n16092), .C2(n16091), .A(n16090), .B(n16089), .ZN(
        n16094) );
  AOI22_X1 U16988 ( .A1(n16142), .A2(n16094), .B1(n16093), .B2(n16141), .ZN(
        P2_U3511) );
  AOI22_X1 U16989 ( .A1(n16146), .A2(n16094), .B1(n10709), .B2(n16143), .ZN(
        P2_U3466) );
  OAI22_X1 U16990 ( .A1(n16098), .A2(n16097), .B1(n16096), .B2(n16095), .ZN(
        n16099) );
  NOR2_X1 U16991 ( .A1(n16100), .A2(n16099), .ZN(n16103) );
  AOI22_X1 U16992 ( .A1(n16101), .A2(n16103), .B1(n8325), .B2(n16155), .ZN(
        P3_U3472) );
  INV_X1 U16993 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n16102) );
  AOI22_X1 U16994 ( .A1(n16104), .A2(n16103), .B1(n16102), .B2(n16160), .ZN(
        P3_U3429) );
  AOI21_X1 U16995 ( .B1(n16107), .B2(n16106), .A(n16105), .ZN(n16112) );
  NOR2_X1 U16996 ( .A1(n16108), .A2(n16136), .ZN(n16110) );
  NOR4_X1 U16997 ( .A1(n16112), .A2(n16111), .A3(n16110), .A4(n16109), .ZN(
        n16114) );
  AOI22_X1 U16998 ( .A1(n16142), .A2(n16114), .B1(n16113), .B2(n16141), .ZN(
        P2_U3512) );
  AOI22_X1 U16999 ( .A1(n16146), .A2(n16114), .B1(n11147), .B2(n16143), .ZN(
        P2_U3469) );
  OAI22_X1 U17000 ( .A1(n16118), .A2(n16117), .B1(n16116), .B2(n16115), .ZN(
        n16127) );
  AOI21_X1 U17001 ( .B1(n16121), .B2(n16120), .A(n16119), .ZN(n16122) );
  INV_X1 U17002 ( .A(n16122), .ZN(n16125) );
  AOI21_X1 U17003 ( .B1(n16125), .B2(n16124), .A(n16123), .ZN(n16126) );
  AOI211_X1 U17004 ( .C1(n16129), .C2(n16128), .A(n16127), .B(n16126), .ZN(
        n16131) );
  OAI211_X1 U17005 ( .C1(n16133), .C2(n16132), .A(n16131), .B(n16130), .ZN(
        P1_U3215) );
  OAI211_X1 U17006 ( .C1(n16137), .C2(n16136), .A(n16135), .B(n16134), .ZN(
        n16138) );
  AOI21_X1 U17007 ( .B1(n16140), .B2(n16139), .A(n16138), .ZN(n16145) );
  AOI22_X1 U17008 ( .A1(n16142), .A2(n16145), .B1(n10405), .B2(n16141), .ZN(
        P2_U3513) );
  INV_X1 U17009 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n16144) );
  AOI22_X1 U17010 ( .A1(n16146), .A2(n16145), .B1(n16144), .B2(n16143), .ZN(
        P2_U3472) );
  INV_X1 U17011 ( .A(n16147), .ZN(n16150) );
  AOI22_X1 U17012 ( .A1(n16150), .A2(n16149), .B1(SI_15_), .B2(n16148), .ZN(
        n16151) );
  OAI21_X1 U17013 ( .B1(P3_U3151), .B2(n16152), .A(n16151), .ZN(P3_U3280) );
  INV_X1 U17014 ( .A(n16154), .ZN(n16156) );
  AOI22_X1 U17015 ( .A1(n16162), .A2(n16156), .B1(P3_REG1_REG_30__SCAN_IN), 
        .B2(n16155), .ZN(n16158) );
  NAND2_X1 U17016 ( .A1(n16158), .A2(n16157), .ZN(P3_U3489) );
  INV_X1 U17017 ( .A(n16159), .ZN(n16161) );
  AOI22_X1 U17018 ( .A1(n16162), .A2(n16161), .B1(P3_REG0_REG_30__SCAN_IN), 
        .B2(n16160), .ZN(n16164) );
  NAND2_X1 U17019 ( .A1(n16164), .A2(n16163), .ZN(P3_U3457) );
  AOI21_X1 U17020 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n16165) );
  OAI21_X1 U17021 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n16165), 
        .ZN(U28) );
  NOR2_X1 U9484 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n7879) );
  AND3_X1 U11385 ( .A1(n9563), .A2(n9478), .A3(n9477), .ZN(n9482) );
  AND3_X1 U10853 ( .A1(n9085), .A2(n9084), .A3(n9083), .ZN(n15170) );
  INV_X2 U7396 ( .A(n12314), .ZN(n12342) );
  INV_X2 U7290 ( .A(n12884), .ZN(n12868) );
  NAND2_X1 U7350 ( .A1(n10387), .A2(n10386), .ZN(n10594) );
  NAND2_X1 U7349 ( .A1(n10600), .A2(n10599), .ZN(n10819) );
  INV_X1 U7397 ( .A(n8182), .ZN(n12314) );
  NAND2_X1 U9372 ( .A1(n7589), .A2(n9312), .ZN(n12802) );
  CLKBUF_X1 U7327 ( .A(n8298), .Z(n8754) );
  XNOR2_X1 U7361 ( .A(n9305), .B(n9304), .ZN(n9367) );
  NAND2_X2 U7480 ( .A1(n7181), .A2(n14952), .ZN(n12524) );
  CLKBUF_X2 U7481 ( .A(n14869), .Z(n7185) );
  CLKBUF_X1 U7568 ( .A(n11374), .Z(n14043) );
  CLKBUF_X1 U7569 ( .A(n8990), .Z(n9540) );
endmodule

