

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4367, n4368, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569;

  AOI211_X1 U4872 ( .C1(n10306), .C2(n10214), .A(n10213), .B(n10212), .ZN(
        n10215) );
  INV_X1 U4873 ( .A(n9521), .ZN(n9437) );
  AOI211_X1 U4874 ( .C1(n10294), .C2(n7504), .A(n10456), .B(n4494), .ZN(n10293) );
  INV_X2 U4875 ( .A(n9484), .ZN(n9538) );
  AND2_X1 U4876 ( .A1(n8171), .A2(n8170), .ZN(n8943) );
  OR2_X1 U4877 ( .A1(n10219), .A2(n9843), .ZN(n8506) );
  NAND2_X1 U4878 ( .A1(n6842), .A2(n6841), .ZN(n6813) );
  INV_X2 U4879 ( .A(n5828), .ZN(n5841) );
  INV_X1 U4880 ( .A(n5548), .ZN(n5672) );
  AND2_X1 U4881 ( .A1(n6718), .A2(n6717), .ZN(n7289) );
  NAND2_X1 U4882 ( .A1(n6051), .A2(n8825), .ZN(n5711) );
  OR2_X1 U4883 ( .A1(n6928), .A2(n7008), .ZN(n8210) );
  INV_X1 U4884 ( .A(n4606), .ZN(n10496) );
  NAND4_X1 U4885 ( .A1(n6413), .A2(n6414), .A3(n6415), .A4(n6416), .ZN(n9856)
         );
  NAND4_X1 U4886 ( .A1(n6370), .A2(n6368), .A3(n6369), .A4(n6367), .ZN(n9859)
         );
  NAND2_X2 U4887 ( .A1(n8283), .A2(n8438), .ZN(n7143) );
  NAND2_X1 U4888 ( .A1(n5192), .A2(n5209), .ZN(n5194) );
  NOR2_X1 U4889 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5992) );
  NOR2_X1 U4890 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n8773) );
  INV_X1 U4891 ( .A(n6402), .ZN(n4376) );
  NOR3_X1 U4892 ( .A1(n9341), .A2(n9326), .A3(n9548), .ZN(n7846) );
  NAND2_X1 U4893 ( .A1(n9792), .A2(n9793), .ZN(n8099) );
  NAND2_X1 U4894 ( .A1(n4584), .A2(n4515), .ZN(n9791) );
  INV_X1 U4895 ( .A(n8154), .ZN(n8935) );
  INV_X1 U4896 ( .A(n6516), .ZN(n7910) );
  AOI21_X1 U4897 ( .B1(n7254), .B2(n8228), .A(n8311), .ZN(n7460) );
  NAND2_X1 U4898 ( .A1(n10207), .A2(n8943), .ZN(n8498) );
  INV_X1 U4899 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8570) );
  INV_X1 U4901 ( .A(n6840), .ZN(n7415) );
  NAND2_X1 U4902 ( .A1(n7952), .A2(n7951), .ZN(n9823) );
  CLKBUF_X3 U4903 ( .A(n7872), .Z(n4368) );
  INV_X1 U4904 ( .A(n9857), .ZN(n6590) );
  CLKBUF_X3 U4905 ( .A(n8135), .Z(n8112) );
  NAND2_X1 U4906 ( .A1(n7704), .A2(n6023), .ZN(n6371) );
  NAND2_X1 U4907 ( .A1(n6017), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U4908 ( .A1(n5417), .A2(n5416), .ZN(n5401) );
  NOR2_X2 U4909 ( .A1(n5114), .A2(n5113), .ZN(n9179) );
  NAND2_X1 U4910 ( .A1(n7909), .A2(n7908), .ZN(n10207) );
  NAND2_X1 U4911 ( .A1(n6695), .A2(n6694), .ZN(n6883) );
  INV_X1 U4912 ( .A(n4379), .ZN(n4380) );
  XNOR2_X1 U4913 ( .A(n6188), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6296) );
  OAI21_X1 U4914 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10528), .ZN(n10557) );
  INV_X1 U4915 ( .A(n9529), .ZN(n6051) );
  INV_X1 U4916 ( .A(n5931), .ZN(n4822) );
  AND2_X1 U4917 ( .A1(n9816), .A2(n4392), .ZN(n8958) );
  NAND2_X1 U4918 ( .A1(n6363), .A2(n6358), .ZN(n10348) );
  BUF_X1 U4919 ( .A(n6293), .Z(n4373) );
  OR3_X2 U4921 ( .A1(n8436), .A2(n8435), .A3(n8434), .ZN(n4415) );
  XNOR2_X2 U4922 ( .A(n5191), .B(n5189), .ZN(n6624) );
  NAND4_X4 U4924 ( .A1(n5130), .A2(n5128), .A3(n5129), .A4(n5131), .ZN(n6045)
         );
  INV_X2 U4925 ( .A(n7322), .ZN(n8825) );
  OAI21_X2 U4926 ( .B1(n8524), .B2(n9196), .A(n6758), .ZN(n9202) );
  XNOR2_X2 U4927 ( .A(n5216), .B(n5233), .ZN(n6885) );
  BUF_X4 U4929 ( .A(n6700), .Z(n4367) );
  BUF_X4 U4930 ( .A(n6700), .Z(n8934) );
  NAND2_X4 U4931 ( .A1(n6402), .A2(n6352), .ZN(n8154) );
  AND2_X2 U4932 ( .A1(n8210), .A2(n8405), .ZN(n8294) );
  INV_X4 U4933 ( .A(n8882), .ZN(n8872) );
  INV_X1 U4934 ( .A(n6425), .ZN(n6572) );
  INV_X1 U4935 ( .A(n8190), .ZN(n4379) );
  NAND2_X2 U4936 ( .A1(n5065), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5063) );
  INV_X1 U4937 ( .A(n6622), .ZN(n7872) );
  NOR2_X2 U4938 ( .A1(n10554), .A2(n10367), .ZN(n10368) );
  INV_X1 U4939 ( .A(n6373), .ZN(n6444) );
  NAND2_X2 U4940 ( .A1(n6420), .A2(n6421), .ZN(n8217) );
  XNOR2_X2 U4941 ( .A(n5194), .B(n5212), .ZN(n6696) );
  NAND2_X1 U4942 ( .A1(n4882), .A2(n4880), .ZN(n7254) );
  BUF_X8 U4943 ( .A(n6398), .Z(n5627) );
  OAI21_X4 U4944 ( .B1(n7471), .B2(n7477), .A(n5890), .ZN(n7664) );
  NAND2_X2 U4945 ( .A1(n4969), .A2(n4967), .ZN(n7471) );
  XNOR2_X2 U4946 ( .A(n5401), .B(n5400), .ZN(n7864) );
  AOI211_X2 U4947 ( .C1(n5837), .C2(n5836), .A(n5835), .B(n5839), .ZN(n4589)
         );
  BUF_X2 U4951 ( .A(n8960), .Z(n4372) );
  NAND2_X1 U4952 ( .A1(n6365), .A2(n10348), .ZN(n6707) );
  XNOR2_X2 U4953 ( .A(n6357), .B(P1_IR_REG_30__SCAN_IN), .ZN(n6365) );
  AOI21_X2 U4954 ( .B1(n9059), .B2(n8864), .A(n8863), .ZN(n9028) );
  AOI21_X2 U4955 ( .B1(n8857), .B2(n4665), .A(n5035), .ZN(n9059) );
  OAI21_X2 U4956 ( .B1(n7664), .B2(n5898), .A(n5897), .ZN(n7683) );
  AOI22_X2 U4957 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .B1(n10359), .B2(n6661), .ZN(n10565) );
  INV_X2 U4958 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6661) );
  NAND2_X2 U4959 ( .A1(n7875), .A2(n7874), .ZN(n10253) );
  NOR2_X1 U4960 ( .A1(n9702), .A2(n9701), .ZN(n9768) );
  OR2_X1 U4961 ( .A1(n9341), .A2(n9326), .ZN(n9324) );
  INV_X2 U4962 ( .A(n8532), .ZN(n8535) );
  OR2_X1 U4963 ( .A1(n10207), .A2(n8943), .ZN(n8370) );
  NAND2_X1 U4964 ( .A1(n7901), .A2(n7900), .ZN(n10219) );
  NAND2_X1 U4965 ( .A1(n7897), .A2(n7896), .ZN(n10222) );
  NAND2_X1 U4966 ( .A1(n7892), .A2(n7891), .ZN(n10229) );
  NAND2_X1 U4967 ( .A1(n7884), .A2(n7883), .ZN(n10237) );
  AOI211_X1 U4968 ( .C1(n9629), .C2(n4959), .A(n9538), .B(n7723), .ZN(n9628)
         );
  NAND2_X1 U4969 ( .A1(n9623), .A2(n9014), .ZN(n7540) );
  INV_X2 U4970 ( .A(n9536), .ZN(n4374) );
  NAND2_X1 U4971 ( .A1(n9629), .A2(n7671), .ZN(n5743) );
  NAND2_X1 U4972 ( .A1(n6928), .A2(n7008), .ZN(n8405) );
  INV_X1 U4973 ( .A(n9855), .ZN(n6670) );
  NAND2_X1 U4974 ( .A1(n6934), .A2(n7174), .ZN(n8403) );
  INV_X2 U4975 ( .A(n6866), .ZN(n9176) );
  INV_X1 U4976 ( .A(n5104), .ZN(n8834) );
  INV_X1 U4977 ( .A(n8388), .ZN(n8381) );
  NAND4_X2 U4978 ( .A1(n6569), .A2(n6573), .A3(n6571), .A4(n6570), .ZN(n4505)
         );
  INV_X1 U4979 ( .A(n7399), .ZN(n10455) );
  CLKBUF_X2 U4980 ( .A(n5467), .Z(n5548) );
  INV_X1 U4981 ( .A(n5157), .ZN(n5615) );
  BUF_X2 U4982 ( .A(n6707), .Z(n8187) );
  NAND2_X1 U4983 ( .A1(n8933), .A2(n9683), .ZN(n5143) );
  INV_X1 U4984 ( .A(n8286), .ZN(n8438) );
  AND4_X1 U4985 ( .A1(n5153), .A2(n5311), .A3(n5310), .A4(n5059), .ZN(n4383)
         );
  INV_X1 U4986 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6002) );
  INV_X2 U4987 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X4 U4988 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9677) );
  OR2_X1 U4989 ( .A1(n9813), .A2(n8140), .ZN(n9816) );
  AND2_X1 U4990 ( .A1(n5882), .A2(n5881), .ZN(n4732) );
  OAI21_X1 U4991 ( .B1(n5861), .B2(n6037), .A(n4822), .ZN(n4588) );
  AND2_X1 U4992 ( .A1(n4857), .A2(n4414), .ZN(n8533) );
  OAI211_X1 U4993 ( .C1(n9560), .C2(n9627), .A(n9559), .B(n9558), .ZN(n9561)
         );
  AND2_X1 U4994 ( .A1(n8432), .A2(n4536), .ZN(n4535) );
  NOR2_X1 U4995 ( .A1(n9550), .A2(n4650), .ZN(n9552) );
  NOR2_X1 U4996 ( .A1(n4625), .A2(n4788), .ZN(n4624) );
  OR2_X1 U4997 ( .A1(n8536), .A2(n8535), .ZN(n5050) );
  NOR2_X1 U4998 ( .A1(n9126), .A2(n9127), .ZN(n9125) );
  AND2_X1 U4999 ( .A1(n4538), .A2(n4537), .ZN(n4536) );
  AND2_X1 U5000 ( .A1(n9299), .A2(n9544), .ZN(n5985) );
  XNOR2_X1 U5001 ( .A(n9300), .B(n5978), .ZN(n5979) );
  AOI21_X1 U5002 ( .B1(n4855), .B2(n4853), .A(n4433), .ZN(n4852) );
  NAND2_X1 U5003 ( .A1(n4686), .A2(n8371), .ZN(n8387) );
  NAND2_X1 U5004 ( .A1(n7937), .A2(n7936), .ZN(n9689) );
  CLKBUF_X1 U5005 ( .A(n10045), .Z(n4504) );
  OAI21_X1 U5006 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10531), .ZN(n10529) );
  NAND2_X1 U5007 ( .A1(n5578), .A2(n5577), .ZN(n9566) );
  OR2_X1 U5008 ( .A1(n10229), .A2(n10015), .ZN(n8487) );
  AND2_X1 U5009 ( .A1(n4783), .A2(n4473), .ZN(n9934) );
  INV_X1 U5010 ( .A(n8255), .ZN(n8360) );
  NOR2_X1 U5011 ( .A1(n8467), .A2(n8466), .ZN(n10125) );
  AND2_X1 U5012 ( .A1(n10232), .A2(n10004), .ZN(n8255) );
  OR2_X1 U5013 ( .A1(n10232), .A2(n10004), .ZN(n8486) );
  NAND2_X1 U5014 ( .A1(n7882), .A2(n7881), .ZN(n10243) );
  NAND2_X1 U5015 ( .A1(n5557), .A2(n5556), .ZN(n5573) );
  XNOR2_X1 U5016 ( .A(n5555), .B(n5554), .ZN(n7885) );
  NAND2_X1 U5017 ( .A1(n7879), .A2(n7878), .ZN(n10249) );
  NAND3_X1 U5018 ( .A1(n4571), .A2(n4569), .A3(n4573), .ZN(n6690) );
  NAND2_X1 U5019 ( .A1(n5462), .A2(n5461), .ZN(n9595) );
  XNOR2_X1 U5020 ( .A(n5492), .B(n5512), .ZN(n7880) );
  INV_X1 U5021 ( .A(n9969), .ZN(n9843) );
  INV_X1 U5022 ( .A(n7045), .ZN(n4848) );
  XNOR2_X1 U5023 ( .A(n5478), .B(n5477), .ZN(n7876) );
  NAND2_X1 U5024 ( .A1(n10112), .A2(n10131), .ZN(n4838) );
  AND2_X1 U5025 ( .A1(n8109), .A2(n8108), .ZN(n9993) );
  AND2_X2 U5026 ( .A1(n8131), .A2(n8130), .ZN(n9969) );
  NAND2_X1 U5027 ( .A1(n10273), .A2(n9760), .ZN(n8471) );
  AND2_X1 U5028 ( .A1(n8081), .A2(n8080), .ZN(n10015) );
  NAND2_X1 U5029 ( .A1(n10294), .A2(n7628), .ZN(n8318) );
  NAND2_X1 U5030 ( .A1(n5334), .A2(n5333), .ZN(n7805) );
  NAND2_X1 U5031 ( .A1(n7619), .A2(n7618), .ZN(n10288) );
  NAND2_X1 U5032 ( .A1(n7252), .A2(n7251), .ZN(n7507) );
  NAND3_X1 U5033 ( .A1(n5295), .A2(n4591), .A3(n4590), .ZN(n9623) );
  NAND2_X1 U5034 ( .A1(n7857), .A2(n7856), .ZN(n10283) );
  OAI21_X2 U5035 ( .B1(n6872), .B2(n6871), .A(n6062), .ZN(n6941) );
  NAND2_X1 U5036 ( .A1(n5316), .A2(n5315), .ZN(n7700) );
  NAND2_X1 U5037 ( .A1(n8022), .A2(n8021), .ZN(n10047) );
  OAI22_X1 U5038 ( .A1(n8294), .A2(n6996), .B1(n7368), .B2(n9853), .ZN(n7038)
         );
  AND2_X1 U5039 ( .A1(n5889), .A2(n4975), .ZN(n4974) );
  NAND2_X1 U5040 ( .A1(n7140), .A2(n7139), .ZN(n10305) );
  INV_X1 U5041 ( .A(n8294), .ZN(n4375) );
  NAND2_X1 U5042 ( .A1(n5357), .A2(n4394), .ZN(n4769) );
  INV_X1 U5043 ( .A(n6932), .ZN(n7368) );
  XNOR2_X1 U5044 ( .A(n5290), .B(n4666), .ZN(n7203) );
  INV_X1 U5045 ( .A(n7253), .ZN(n9850) );
  AND2_X1 U5046 ( .A1(n7525), .A2(n5848), .ZN(n5725) );
  AND2_X1 U5047 ( .A1(n7058), .A2(n7057), .ZN(n7253) );
  NAND2_X1 U5048 ( .A1(n6699), .A2(n6698), .ZN(n6928) );
  NAND2_X2 U5049 ( .A1(n6887), .A2(n6886), .ZN(n6999) );
  NAND2_X1 U5050 ( .A1(n5247), .A2(n5246), .ZN(n7449) );
  NAND2_X1 U5051 ( .A1(n6745), .A2(n4505), .ZN(n7004) );
  AND4_X1 U5052 ( .A1(n5265), .A2(n5264), .A3(n5263), .A4(n5262), .ZN(n7671)
         );
  NAND2_X1 U5053 ( .A1(n6442), .A2(n7143), .ZN(n8135) );
  OR2_X1 U5054 ( .A1(n6502), .A2(n4442), .ZN(n4798) );
  AND4_X1 U5055 ( .A1(n5188), .A2(n5187), .A3(n5186), .A4(n5185), .ZN(n7100)
         );
  INV_X1 U5056 ( .A(n6946), .ZN(n9177) );
  NAND2_X1 U5057 ( .A1(n10370), .A2(n10369), .ZN(n10371) );
  BUF_X1 U5058 ( .A(n6446), .Z(n9857) );
  AND4_X1 U5059 ( .A1(n5109), .A2(n5108), .A3(n5107), .A4(n5106), .ZN(n6946)
         );
  INV_X1 U5060 ( .A(n7131), .ZN(n6678) );
  AND3_X1 U5061 ( .A1(n6641), .A2(n6640), .A3(n6639), .ZN(n7008) );
  INV_X2 U5062 ( .A(n5636), .ZN(n5598) );
  OR2_X2 U5063 ( .A1(n5959), .A2(n9359), .ZN(n8835) );
  AND4_X1 U5064 ( .A1(n5147), .A2(n5146), .A3(n5145), .A4(n5144), .ZN(n9529)
         );
  XNOR2_X1 U5065 ( .A(n4919), .B(n6002), .ZN(n8960) );
  CLKBUF_X3 U5066 ( .A(n6714), .Z(n8186) );
  NOR2_X1 U5067 ( .A1(n10386), .A2(n10385), .ZN(n10388) );
  AND2_X1 U5068 ( .A1(n5396), .A2(n5379), .ZN(n4768) );
  CLKBUF_X1 U5069 ( .A(n7852), .Z(n7911) );
  AND2_X1 U5070 ( .A1(n6000), .A2(n5999), .ZN(n8283) );
  INV_X2 U5071 ( .A(n4370), .ZN(n4721) );
  INV_X2 U5072 ( .A(n6771), .ZN(n5460) );
  NAND2_X1 U5073 ( .A1(n6622), .A2(n6398), .ZN(n6516) );
  OAI21_X1 U5074 ( .B1(n5696), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5699) );
  NAND2_X1 U5075 ( .A1(n6358), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6357) );
  CLKBUF_X1 U5076 ( .A(n6248), .Z(n7916) );
  CLKBUF_X2 U5077 ( .A(n5065), .Z(n9678) );
  XNOR2_X1 U5078 ( .A(n6198), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6697) );
  NAND3_X1 U5079 ( .A1(n5077), .A2(n5076), .A3(n5075), .ZN(n6774) );
  OAI21_X1 U5080 ( .B1(n9183), .B2(n9182), .A(n9184), .ZN(n9186) );
  NAND2_X1 U5081 ( .A1(n5060), .A2(n4560), .ZN(n5873) );
  AND2_X1 U5082 ( .A1(n5402), .A2(n4807), .ZN(n5457) );
  NAND2_X1 U5083 ( .A1(n5060), .A2(n4561), .ZN(n5077) );
  AND2_X1 U5084 ( .A1(n4602), .A2(n4383), .ZN(n4560) );
  NOR2_X1 U5085 ( .A1(n6026), .A2(n6033), .ZN(n4823) );
  AND3_X1 U5086 ( .A1(n4602), .A2(n4383), .A3(n4398), .ZN(n4561) );
  AND2_X1 U5087 ( .A1(n4602), .A2(n4383), .ZN(n5402) );
  NAND3_X1 U5088 ( .A1(n4921), .A2(n5988), .A3(n6174), .ZN(n6026) );
  AND2_X1 U5089 ( .A1(n4417), .A2(n4601), .ZN(n4602) );
  OR2_X1 U5090 ( .A1(n6032), .A2(n6028), .ZN(n6010) );
  AND2_X1 U5091 ( .A1(n5154), .A2(n5080), .ZN(n5113) );
  AND2_X1 U5092 ( .A1(n5153), .A2(n5059), .ZN(n5154) );
  NAND2_X1 U5093 ( .A1(n5044), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n6361) );
  NAND2_X1 U5094 ( .A1(n6359), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6360) );
  NAND3_X1 U5095 ( .A1(n4664), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4662) );
  INV_X1 U5096 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5062) );
  INV_X1 U5097 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n8553) );
  INV_X1 U5098 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6030) );
  INV_X1 U5099 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5456) );
  INV_X1 U5100 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6177) );
  INV_X2 U5101 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8561) );
  NOR2_X1 U5102 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5056) );
  NOR3_X1 U5103 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .A3(
        P2_IR_REG_3__SCAN_IN), .ZN(n4601) );
  INV_X1 U5104 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5404) );
  NOR2_X2 U5105 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6174) );
  NOR2_X1 U5106 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5311) );
  NOR2_X1 U5107 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5310) );
  INV_X1 U5108 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8763) );
  NOR2_X1 U5109 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5989) );
  INV_X4 U5110 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U5111 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5055) );
  INV_X1 U5112 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6190) );
  NAND3_X1 U5113 ( .A1(n9954), .A2(n4661), .A3(n4660), .ZN(n4663) );
  NAND2_X1 U5114 ( .A1(n6622), .A2(n5133), .ZN(n7852) );
  NOR2_X2 U5115 ( .A1(n7504), .A2(n10294), .ZN(n4494) );
  INV_X1 U5116 ( .A(n6365), .ZN(n10343) );
  INV_X2 U5117 ( .A(n10348), .ZN(n6364) );
  XOR2_X2 U5118 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n10371), .Z(n10563) );
  AOI21_X2 U5119 ( .B1(n7683), .B2(n7686), .A(n5899), .ZN(n7545) );
  OAI22_X2 U5120 ( .A1(n10165), .A2(n10176), .B1(n10173), .B2(n9830), .ZN(
        n10121) );
  AND2_X2 U5121 ( .A1(n7051), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7149) );
  NOR2_X2 U5122 ( .A1(n7052), .A2(n8764), .ZN(n7051) );
  NAND2_X2 U5123 ( .A1(n6810), .A2(n6815), .ZN(n6809) );
  AND2_X1 U5124 ( .A1(n6771), .A2(n6398), .ZN(n4377) );
  OAI21_X2 U5125 ( .B1(n4848), .B2(n4846), .A(n4844), .ZN(n7459) );
  BUF_X4 U5126 ( .A(n5615), .Z(n4378) );
  NAND2_X1 U5127 ( .A1(n6835), .A2(n5886), .ZN(n6810) );
  XOR2_X2 U5128 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n10374), .Z(n10562) );
  NAND2_X2 U5129 ( .A1(n10373), .A2(n10372), .ZN(n10374) );
  NOR2_X2 U5130 ( .A1(n7472), .A2(n4956), .ZN(n7723) );
  NAND2_X2 U5131 ( .A1(n5845), .A2(n5846), .ZN(n5883) );
  NOR2_X2 U5132 ( .A1(n6637), .A2(n6636), .ZN(n6635) );
  AOI21_X2 U5133 ( .B1(n8446), .B2(n8445), .A(n4545), .ZN(n10165) );
  OAI22_X2 U5134 ( .A1(n7616), .A2(n7615), .B1(n7614), .B2(n7628), .ZN(n8446)
         );
  XNOR2_X2 U5135 ( .A(n8086), .B(P1_REG3_REG_23__SCAN_IN), .ZN(n10021) );
  XNOR2_X2 U5136 ( .A(n8183), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n8948) );
  NOR4_X2 U5137 ( .A1(n8386), .A2(n8385), .A3(n8425), .A4(n8384), .ZN(n8392)
         );
  AND2_X1 U5138 ( .A1(n9725), .A2(n8044), .ZN(n8047) );
  OR2_X1 U5139 ( .A1(n10201), .A2(n8947), .ZN(n8254) );
  INV_X1 U5140 ( .A(n4780), .ZN(n4779) );
  OAI21_X1 U5141 ( .B1(n5643), .B2(n4781), .A(n5659), .ZN(n4780) );
  NAND2_X1 U5142 ( .A1(n5450), .A2(n5449), .ZN(n4675) );
  INV_X1 U5143 ( .A(n5448), .ZN(n5449) );
  AND2_X1 U5144 ( .A1(n5584), .A2(n5806), .ZN(n5033) );
  NAND2_X1 U5145 ( .A1(n9388), .A2(n5553), .ZN(n5034) );
  AND2_X1 U5146 ( .A1(n9353), .A2(n4659), .ZN(n5584) );
  AND2_X1 U5147 ( .A1(n4418), .A2(n4835), .ZN(n4832) );
  NAND2_X1 U5148 ( .A1(n10243), .A2(n4836), .ZN(n4835) );
  NAND2_X1 U5149 ( .A1(n10046), .A2(n4720), .ZN(n10045) );
  XNOR2_X1 U5150 ( .A(n5431), .B(SI_17_), .ZN(n5429) );
  OR2_X1 U5151 ( .A1(n9570), .A2(n9160), .ZN(n5925) );
  XNOR2_X1 U5152 ( .A(n9901), .B(n9889), .ZN(n9878) );
  INV_X1 U5153 ( .A(n7630), .ZN(n8325) );
  INV_X1 U5154 ( .A(n8353), .ZN(n4718) );
  OR2_X1 U5155 ( .A1(n7717), .A2(n7449), .ZN(n5739) );
  OR2_X1 U5156 ( .A1(n8177), .A2(n9839), .ZN(n8380) );
  INV_X1 U5157 ( .A(n5817), .ZN(n4729) );
  NAND2_X1 U5158 ( .A1(n9353), .A2(n4731), .ZN(n4730) );
  AOI22_X1 U5159 ( .A1(n5809), .A2(n5808), .B1(n5841), .B2(n5807), .ZN(n4587)
         );
  AOI21_X1 U5160 ( .B1(n7840), .B2(n5820), .A(n5821), .ZN(n5008) );
  NAND2_X1 U5161 ( .A1(n5031), .A2(n7331), .ZN(n5029) );
  OR2_X1 U5162 ( .A1(n10253), .A2(n10063), .ZN(n8341) );
  NAND2_X1 U5163 ( .A1(n5647), .A2(n4471), .ZN(n4781) );
  NAND2_X1 U5164 ( .A1(n5328), .A2(n5327), .ZN(n5352) );
  INV_X1 U5165 ( .A(n5271), .ZN(n4492) );
  NAND2_X1 U5166 ( .A1(n5275), .A2(n5303), .ZN(n4667) );
  NAND2_X1 U5167 ( .A1(n4531), .A2(n4532), .ZN(n5254) );
  OR2_X1 U5168 ( .A1(n5627), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n4532) );
  NAND2_X1 U5169 ( .A1(n5627), .A2(n5252), .ZN(n4531) );
  NAND2_X1 U5170 ( .A1(n4534), .A2(n4533), .ZN(n5242) );
  OR2_X1 U5171 ( .A1(n5627), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n4534) );
  NAND2_X1 U5172 ( .A1(n5627), .A2(n6194), .ZN(n4533) );
  NAND2_X1 U5173 ( .A1(n5193), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n4508) );
  AND2_X1 U5174 ( .A1(n8986), .A2(n8851), .ZN(n8853) );
  AND2_X1 U5175 ( .A1(n8962), .A2(n5705), .ZN(n5828) );
  AND2_X1 U5176 ( .A1(n5838), .A2(n4463), .ZN(n5019) );
  INV_X1 U5177 ( .A(n9683), .ZN(n5070) );
  INV_X1 U5178 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5061) );
  OR2_X1 U5179 ( .A1(n9308), .A2(n7844), .ZN(n5832) );
  INV_X1 U5180 ( .A(n4995), .ZN(n4994) );
  OAI21_X1 U5181 ( .B1(n4554), .B2(n4553), .A(n5773), .ZN(n4552) );
  NAND2_X1 U5182 ( .A1(n4441), .A2(n5775), .ZN(n4553) );
  OR2_X1 U5183 ( .A1(n9623), .A2(n9014), .ZN(n5853) );
  NAND2_X1 U5184 ( .A1(n7088), .A2(n4606), .ZN(n5849) );
  NOR2_X1 U5185 ( .A1(n5870), .A2(n4437), .ZN(n4600) );
  NAND3_X1 U5186 ( .A1(n9828), .A2(n9823), .A3(n4462), .ZN(n4584) );
  INV_X1 U5187 ( .A(n4930), .ZN(n4924) );
  NOR2_X1 U5188 ( .A1(n6475), .A2(n4637), .ZN(n4636) );
  INV_X1 U5189 ( .A(n6472), .ZN(n4637) );
  NAND2_X1 U5190 ( .A1(n9917), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4787) );
  NAND2_X1 U5191 ( .A1(n4460), .A2(n4896), .ZN(n4895) );
  XNOR2_X1 U5192 ( .A(n6446), .B(n6445), .ZN(n6455) );
  NOR2_X1 U5193 ( .A1(n4767), .A2(n5472), .ZN(n4766) );
  INV_X1 U5194 ( .A(n5515), .ZN(n4767) );
  NAND2_X1 U5195 ( .A1(n4448), .A2(n4764), .ZN(n4763) );
  NAND2_X1 U5196 ( .A1(n4765), .A2(n5515), .ZN(n4764) );
  INV_X1 U5197 ( .A(n5490), .ZN(n4765) );
  INV_X1 U5198 ( .A(n5471), .ZN(n5474) );
  NAND2_X1 U5199 ( .A1(n4675), .A2(n5452), .ZN(n5471) );
  INV_X1 U5200 ( .A(n4672), .ZN(n4671) );
  OAI21_X1 U5201 ( .B1(n4768), .B2(n4407), .A(n5418), .ZN(n4672) );
  NAND2_X1 U5202 ( .A1(n5416), .A2(n5383), .ZN(n5395) );
  XNOR2_X1 U5203 ( .A(n4757), .B(n8578), .ZN(n5304) );
  AND2_X1 U5204 ( .A1(n8879), .A2(n8877), .ZN(n8898) );
  OR2_X1 U5205 ( .A1(n5579), .A2(n9029), .ZN(n5596) );
  NAND2_X1 U5206 ( .A1(n5560), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5579) );
  INV_X1 U5207 ( .A(n5561), .ZN(n5560) );
  INV_X1 U5208 ( .A(n5141), .ZN(n5636) );
  NAND2_X1 U5209 ( .A1(n4677), .A2(n4676), .ZN(n9126) );
  OR2_X1 U5210 ( .A1(n8866), .A2(n9026), .ZN(n4676) );
  NAND2_X1 U5211 ( .A1(n5863), .A2(n9359), .ZN(n6038) );
  NAND2_X1 U5212 ( .A1(n5832), .A2(n5833), .ZN(n5933) );
  OR2_X1 U5213 ( .A1(n5634), .A2(n5633), .ZN(n9307) );
  NAND2_X1 U5214 ( .A1(n4983), .A2(n4978), .ZN(n4977) );
  INV_X1 U5215 ( .A(n4412), .ZN(n4978) );
  AOI21_X2 U5216 ( .B1(n9460), .B2(n5507), .A(n5506), .ZN(n5508) );
  OR2_X1 U5217 ( .A1(n5036), .A2(n4419), .ZN(n5506) );
  NAND2_X1 U5218 ( .A1(n5423), .A2(n5422), .ZN(n9512) );
  CLKBUF_X1 U5219 ( .A(n9447), .Z(n9448) );
  NAND2_X2 U5220 ( .A1(n7757), .A2(n6774), .ZN(n6771) );
  AOI21_X1 U5221 ( .B1(n4943), .B2(n5047), .A(n4434), .ZN(n4942) );
  OR3_X2 U5222 ( .A1(n8532), .A2(n8280), .A3(n8507), .ZN(n8281) );
  NAND2_X1 U5223 ( .A1(n10343), .A2(n6364), .ZN(n6425) );
  NAND2_X1 U5224 ( .A1(n6296), .A2(n8682), .ZN(n4641) );
  OR2_X1 U5225 ( .A1(n6189), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n6192) );
  NAND2_X1 U5226 ( .A1(n4799), .A2(n10402), .ZN(n4797) );
  INV_X1 U5227 ( .A(n10409), .ZN(n4799) );
  NOR2_X1 U5228 ( .A1(n9866), .A2(n9865), .ZN(n9885) );
  NAND2_X1 U5229 ( .A1(n9877), .A2(n9876), .ZN(n9901) );
  NAND2_X1 U5230 ( .A1(n9899), .A2(n4787), .ZN(n4784) );
  OR2_X1 U5231 ( .A1(n9897), .A2(n4785), .ZN(n4783) );
  NAND2_X1 U5232 ( .A1(n4786), .A2(n4787), .ZN(n4785) );
  INV_X1 U5233 ( .A(n9896), .ZN(n4786) );
  INV_X1 U5234 ( .A(n10197), .ZN(n9956) );
  NAND2_X1 U5235 ( .A1(n9980), .A2(n4917), .ZN(n8540) );
  AND2_X1 U5236 ( .A1(n4393), .A2(n4918), .ZN(n4917) );
  NOR2_X2 U5237 ( .A1(n8540), .A2(n10201), .ZN(n9955) );
  NAND2_X1 U5238 ( .A1(n8100), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8124) );
  NAND2_X1 U5239 ( .A1(n8494), .A2(n8493), .ZN(n9989) );
  OR2_X1 U5240 ( .A1(n10229), .A2(n9844), .ZN(n8457) );
  AOI21_X1 U5241 ( .B1(n10045), .B2(n4408), .A(n4860), .ZN(n4859) );
  NAND2_X1 U5242 ( .A1(n4861), .A2(n8486), .ZN(n4860) );
  NAND2_X1 U5243 ( .A1(n4408), .A2(n4865), .ZN(n4861) );
  AOI21_X1 U5244 ( .B1(n4388), .B2(n4831), .A(n4443), .ZN(n4826) );
  AND2_X1 U5245 ( .A1(n10288), .A2(n9846), .ZN(n4545) );
  NAND2_X1 U5246 ( .A1(n9859), .A2(n6444), .ZN(n6448) );
  NOR2_X1 U5247 ( .A1(n6027), .A2(n6031), .ZN(n4824) );
  NOR2_X1 U5248 ( .A1(n6028), .A2(n6032), .ZN(n4825) );
  NAND2_X1 U5249 ( .A1(n5491), .A2(n5490), .ZN(n5516) );
  OR2_X1 U5250 ( .A1(n6192), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6202) );
  CLKBUF_X1 U5251 ( .A(n6027), .Z(n5990) );
  BUF_X4 U5252 ( .A(n5193), .Z(n6398) );
  INV_X1 U5253 ( .A(n4647), .ZN(n4646) );
  OAI21_X1 U5254 ( .B1(n10393), .B2(n4648), .A(n6273), .ZN(n4647) );
  AND2_X1 U5255 ( .A1(n4519), .A2(n9951), .ZN(n4625) );
  OAI21_X1 U5256 ( .B1(n9949), .B2(n9948), .A(n4391), .ZN(n4519) );
  NAND2_X1 U5257 ( .A1(n9950), .A2(n10427), .ZN(n4626) );
  OR2_X1 U5258 ( .A1(n4694), .A2(n4695), .ZN(n4692) );
  AND2_X1 U5259 ( .A1(n4698), .A2(n4696), .ZN(n4695) );
  NAND2_X1 U5260 ( .A1(n8292), .A2(n8388), .ZN(n4698) );
  NAND2_X1 U5261 ( .A1(n4697), .A2(n8381), .ZN(n4696) );
  NAND2_X1 U5262 ( .A1(n4381), .A2(n4432), .ZN(n4726) );
  INV_X1 U5263 ( .A(n5765), .ZN(n4723) );
  OAI21_X1 U5264 ( .B1(n8324), .B2(n8325), .A(n10177), .ZN(n4702) );
  NOR2_X1 U5265 ( .A1(n8325), .A2(n8321), .ZN(n4704) );
  INV_X1 U5266 ( .A(n8358), .ZN(n4719) );
  NOR2_X1 U5267 ( .A1(n4718), .A2(n4715), .ZN(n4714) );
  INV_X1 U5268 ( .A(n8349), .ZN(n4715) );
  OAI21_X1 U5269 ( .B1(n4716), .B2(n8358), .A(n8357), .ZN(n4713) );
  INV_X1 U5270 ( .A(n4717), .ZN(n4716) );
  OAI21_X1 U5271 ( .B1(n4718), .B2(n10060), .A(n4720), .ZN(n4717) );
  NAND2_X1 U5272 ( .A1(n4743), .A2(n4740), .ZN(n4739) );
  NOR2_X1 U5273 ( .A1(n4742), .A2(n4741), .ZN(n4740) );
  OAI21_X1 U5274 ( .B1(n5045), .B2(n5792), .A(n5791), .ZN(n4743) );
  NAND2_X1 U5275 ( .A1(n5796), .A2(n5841), .ZN(n4741) );
  INV_X1 U5276 ( .A(n5805), .ZN(n4738) );
  INV_X1 U5277 ( .A(n7536), .ZN(n4605) );
  NOR2_X1 U5278 ( .A1(n4609), .A2(n9496), .ZN(n4608) );
  NOR2_X1 U5279 ( .A1(n7796), .A2(n7742), .ZN(n4615) );
  NOR2_X1 U5280 ( .A1(n4611), .A2(n5854), .ZN(n4610) );
  INV_X1 U5281 ( .A(n4933), .ZN(n4929) );
  NAND2_X1 U5282 ( .A1(n8422), .A2(n4685), .ZN(n4684) );
  NOR2_X1 U5283 ( .A1(n8947), .A2(n8388), .ZN(n4685) );
  AND2_X1 U5284 ( .A1(n10193), .A2(n8381), .ZN(n8378) );
  INV_X1 U5285 ( .A(n5609), .ZN(n4772) );
  NAND2_X1 U5286 ( .A1(n5330), .A2(n5352), .ZN(n5346) );
  NAND2_X1 U5287 ( .A1(n4757), .A2(SI_11_), .ZN(n5343) );
  NAND2_X1 U5288 ( .A1(n4451), .A2(n4667), .ZN(n5347) );
  NAND2_X1 U5289 ( .A1(n4759), .A2(n4758), .ZN(n4757) );
  OR2_X1 U5290 ( .A1(n5627), .A2(n4760), .ZN(n4759) );
  NAND2_X1 U5291 ( .A1(n5627), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n4758) );
  INV_X1 U5292 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n4760) );
  AND2_X1 U5293 ( .A1(n5267), .A2(n4405), .ZN(n5268) );
  NAND2_X1 U5294 ( .A1(n5254), .A2(n5253), .ZN(n5271) );
  NAND2_X1 U5295 ( .A1(n4436), .A2(n8842), .ZN(n8854) );
  NAND2_X1 U5296 ( .A1(n4585), .A2(n4424), .ZN(n5827) );
  NAND2_X1 U5297 ( .A1(n4586), .A2(n4423), .ZN(n4585) );
  OR2_X1 U5298 ( .A1(n9548), .A2(n5828), .ZN(n4728) );
  NAND2_X1 U5299 ( .A1(n5007), .A2(n5833), .ZN(n5006) );
  AOI21_X1 U5300 ( .B1(n5019), .B2(n4395), .A(n5018), .ZN(n5017) );
  INV_X1 U5301 ( .A(n4444), .ZN(n5018) );
  OR2_X1 U5302 ( .A1(n5143), .A2(n5142), .ZN(n5144) );
  AND2_X1 U5303 ( .A1(n4999), .A2(n4996), .ZN(n4995) );
  NAND2_X1 U5304 ( .A1(n9642), .A2(n9129), .ZN(n5002) );
  OR2_X1 U5305 ( .A1(n9345), .A2(n8869), .ZN(n5815) );
  OR2_X1 U5306 ( .A1(n9566), .A2(n9128), .ZN(n5811) );
  NOR2_X1 U5307 ( .A1(n9570), .A2(n4961), .ZN(n4960) );
  INV_X1 U5308 ( .A(n4962), .ZN(n4961) );
  NOR2_X1 U5309 ( .A1(n9580), .A2(n9383), .ZN(n4962) );
  NAND2_X1 U5310 ( .A1(n5439), .A2(n4652), .ZN(n5481) );
  NOR2_X1 U5311 ( .A1(n9595), .A2(n9489), .ZN(n4952) );
  AND2_X1 U5312 ( .A1(n5022), .A2(n4456), .ZN(n4554) );
  AND2_X1 U5313 ( .A1(n5903), .A2(n7760), .ZN(n5904) );
  NAND2_X1 U5314 ( .A1(n5296), .A2(n4657), .ZN(n5368) );
  AND2_X1 U5315 ( .A1(n4658), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n4657) );
  NAND2_X1 U5316 ( .A1(n5296), .A2(n4658), .ZN(n5336) );
  NAND2_X1 U5317 ( .A1(n9177), .A2(n7415), .ZN(n5724) );
  AND2_X1 U5318 ( .A1(n5863), .A2(n5879), .ZN(n6096) );
  NAND2_X1 U5319 ( .A1(n9157), .A2(n9462), .ZN(n5938) );
  NOR2_X1 U5320 ( .A1(n7435), .A2(n4556), .ZN(n4555) );
  INV_X1 U5321 ( .A(n5736), .ZN(n4556) );
  AND2_X1 U5322 ( .A1(n5405), .A2(n5404), .ZN(n5406) );
  AND2_X1 U5323 ( .A1(n8160), .A2(n8159), .ZN(n8161) );
  AOI21_X1 U5324 ( .B1(n8047), .B2(n4923), .A(n5052), .ZN(n4922) );
  INV_X1 U5325 ( .A(n4926), .ZN(n4923) );
  NOR2_X1 U5326 ( .A1(n10193), .A2(n8374), .ZN(n8425) );
  AND2_X1 U5327 ( .A1(n8365), .A2(n9988), .ZN(n8496) );
  INV_X1 U5328 ( .A(n8366), .ZN(n8495) );
  OAI21_X1 U5329 ( .B1(n8451), .B2(n10074), .A(n8450), .ZN(n8452) );
  AND2_X1 U5330 ( .A1(n8341), .A2(n8344), .ZN(n8451) );
  OR2_X1 U5331 ( .A1(n10273), .A2(n9760), .ZN(n8332) );
  OR2_X1 U5332 ( .A1(n10277), .A2(n10185), .ZN(n8470) );
  OR2_X1 U5333 ( .A1(n10283), .A2(n9830), .ZN(n8465) );
  OR2_X1 U5334 ( .A1(n7260), .A2(n7259), .ZN(n7494) );
  OAI22_X1 U5335 ( .A1(n7246), .A2(n4843), .B1(n10305), .B2(n9850), .ZN(n4845)
         );
  NAND2_X1 U5336 ( .A1(n8305), .A2(n7141), .ZN(n4843) );
  NOR2_X1 U5337 ( .A1(n7060), .A2(n4886), .ZN(n4885) );
  INV_X1 U5338 ( .A(n7005), .ZN(n4886) );
  NAND2_X1 U5339 ( .A1(n7006), .A2(n4885), .ZN(n4884) );
  NAND2_X1 U5340 ( .A1(n4878), .A2(n8298), .ZN(n4881) );
  INV_X1 U5341 ( .A(n8258), .ZN(n4878) );
  NAND2_X1 U5342 ( .A1(n4848), .A2(n8258), .ZN(n7142) );
  INV_X1 U5343 ( .A(n6596), .ZN(n4908) );
  XNOR2_X1 U5344 ( .A(n9856), .B(n8217), .ZN(n8259) );
  NAND2_X1 U5345 ( .A1(n8442), .A2(n10053), .ZN(n6442) );
  AOI21_X1 U5346 ( .B1(n4779), .B2(n4781), .A(n5676), .ZN(n4776) );
  NAND2_X1 U5347 ( .A1(n6353), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U5348 ( .A1(n5626), .A2(n5625), .ZN(n5644) );
  AND2_X1 U5349 ( .A1(n5587), .A2(n5571), .ZN(n4773) );
  OR2_X1 U5350 ( .A1(n5573), .A2(n5572), .ZN(n4774) );
  XNOR2_X1 U5351 ( .A(n5451), .B(SI_18_), .ZN(n5448) );
  NAND2_X1 U5352 ( .A1(n5432), .A2(SI_17_), .ZN(n5433) );
  NAND2_X1 U5353 ( .A1(n5273), .A2(n5272), .ZN(n5303) );
  INV_X1 U5354 ( .A(n4667), .ZN(n4666) );
  NAND2_X1 U5355 ( .A1(n5242), .A2(n5241), .ZN(n5269) );
  INV_X1 U5356 ( .A(n5249), .ZN(n5267) );
  OR2_X1 U5357 ( .A1(n8843), .A2(n9095), .ZN(n8986) );
  NAND2_X1 U5358 ( .A1(n6089), .A2(n6088), .ZN(n4816) );
  AND2_X1 U5359 ( .A1(n8898), .A2(n4683), .ZN(n4682) );
  NAND2_X1 U5360 ( .A1(n8871), .A2(n9127), .ZN(n4683) );
  OR2_X1 U5361 ( .A1(n7098), .A2(n4810), .ZN(n4386) );
  INV_X1 U5362 ( .A(n6077), .ZN(n4810) );
  OR2_X1 U5363 ( .A1(n6771), .A2(n6170), .ZN(n5139) );
  AND2_X1 U5364 ( .A1(n9051), .A2(n4806), .ZN(n4805) );
  NAND2_X1 U5365 ( .A1(n6151), .A2(n6150), .ZN(n4806) );
  NAND2_X1 U5366 ( .A1(n8970), .A2(n6145), .ZN(n9037) );
  AND2_X1 U5367 ( .A1(n4815), .A2(n7514), .ZN(n4814) );
  INV_X1 U5368 ( .A(n6100), .ZN(n4815) );
  INV_X1 U5369 ( .A(n6122), .ZN(n4812) );
  AND2_X1 U5370 ( .A1(n6128), .A2(n6126), .ZN(n7779) );
  NAND2_X1 U5371 ( .A1(n4816), .A2(n4814), .ZN(n7781) );
  NAND2_X1 U5372 ( .A1(n6050), .A2(n7018), .ZN(n4802) );
  AND2_X1 U5373 ( .A1(n7087), .A2(n6862), .ZN(n4382) );
  OR2_X1 U5374 ( .A1(n6865), .A2(n6861), .ZN(n6071) );
  INV_X1 U5375 ( .A(n5858), .ZN(n4618) );
  NOR3_X1 U5376 ( .A1(n5857), .A2(n5933), .A3(n4620), .ZN(n4619) );
  AND2_X1 U5377 ( .A1(n5551), .A2(n5550), .ZN(n9108) );
  AOI21_X1 U5378 ( .B1(n9186), .B2(n8526), .A(n8525), .ZN(n8524) );
  AOI21_X1 U5379 ( .B1(n9202), .B2(n6921), .A(n6920), .ZN(n9214) );
  INV_X1 U5380 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5361) );
  NOR2_X1 U5381 ( .A1(n7178), .A2(n4469), .ZN(n7180) );
  NAND2_X1 U5382 ( .A1(n8909), .A2(n4479), .ZN(n9270) );
  NAND2_X1 U5383 ( .A1(n4953), .A2(n4954), .ZN(n9300) );
  NOR2_X1 U5384 ( .A1(n9548), .A2(n5693), .ZN(n4953) );
  NAND2_X1 U5385 ( .A1(n5595), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5634) );
  AOI22_X1 U5386 ( .A1(n4413), .A2(n5927), .B1(n9319), .B2(n5002), .ZN(n4999)
         );
  NAND2_X1 U5387 ( .A1(n9345), .A2(n8869), .ZN(n9320) );
  NAND2_X1 U5388 ( .A1(n8869), .A2(n9646), .ZN(n5003) );
  NAND2_X1 U5389 ( .A1(n5815), .A2(n9320), .ZN(n9336) );
  OR2_X1 U5390 ( .A1(n9570), .A2(n8983), .ZN(n9352) );
  AOI21_X1 U5391 ( .B1(n4986), .B2(n4396), .A(n4384), .ZN(n4985) );
  NOR2_X1 U5392 ( .A1(n5924), .A2(n4987), .ZN(n4986) );
  NOR2_X1 U5393 ( .A1(n4396), .A2(n5923), .ZN(n4987) );
  OR2_X1 U5394 ( .A1(n9580), .A2(n9005), .ZN(n9389) );
  OR2_X1 U5395 ( .A1(n5919), .A2(n5918), .ZN(n5920) );
  OR2_X1 U5396 ( .A1(n7833), .A2(n9047), .ZN(n9508) );
  NAND2_X1 U5397 ( .A1(n5021), .A2(n4554), .ZN(n4550) );
  NAND2_X1 U5398 ( .A1(n7769), .A2(n5943), .ZN(n7833) );
  AND2_X1 U5399 ( .A1(n9154), .A2(n8971), .ZN(n5943) );
  AOI21_X1 U5400 ( .B1(n7742), .B2(n5375), .A(n5023), .ZN(n5022) );
  NAND2_X1 U5401 ( .A1(n5296), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5318) );
  OR2_X1 U5402 ( .A1(n5284), .A2(n8720), .ZN(n5297) );
  NOR2_X1 U5403 ( .A1(n5027), .A2(n5026), .ZN(n5025) );
  AND4_X1 U5404 ( .A1(n5230), .A2(n5229), .A3(n5228), .A4(n5227), .ZN(n7717)
         );
  AND2_X1 U5405 ( .A1(n5727), .A2(n7475), .ZN(n7331) );
  NAND2_X1 U5406 ( .A1(n5848), .A2(n5849), .ZN(n7536) );
  INV_X1 U5407 ( .A(n9528), .ZN(n9464) );
  NAND2_X1 U5408 ( .A1(n4721), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5180) );
  INV_X1 U5409 ( .A(n9462), .ZN(n9531) );
  INV_X1 U5410 ( .A(n10507), .ZN(n9630) );
  INV_X1 U5411 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4744) );
  NAND2_X1 U5412 ( .A1(n5168), .A2(n5167), .ZN(n5196) );
  INV_X1 U5413 ( .A(n5166), .ZN(n5168) );
  INV_X1 U5414 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5080) );
  NAND2_X1 U5415 ( .A1(n5133), .A2(n5124), .ZN(n5132) );
  NAND2_X1 U5416 ( .A1(n10214), .A2(n4582), .ZN(n4581) );
  AND2_X1 U5417 ( .A1(n4946), .A2(n8099), .ZN(n9702) );
  NOR2_X1 U5418 ( .A1(n9697), .A2(n9699), .ZN(n4946) );
  OR2_X1 U5419 ( .A1(n9748), .A2(n9749), .ZN(n4933) );
  NAND2_X1 U5420 ( .A1(n9748), .A2(n9749), .ZN(n4932) );
  INV_X1 U5421 ( .A(n7645), .ZN(n4940) );
  INV_X1 U5422 ( .A(n4944), .ZN(n4943) );
  OAI21_X1 U5423 ( .B1(n5047), .B2(n7351), .A(n4945), .ZN(n4944) );
  NAND2_X1 U5424 ( .A1(n7149), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7260) );
  OR2_X1 U5425 ( .A1(n10389), .A2(n6309), .ZN(n6314) );
  AOI21_X1 U5426 ( .B1(n6481), .B2(n6480), .A(n6479), .ZN(n6502) );
  OR2_X1 U5427 ( .A1(n4636), .A2(n10405), .ZN(n4635) );
  NAND2_X1 U5428 ( .A1(n4410), .A2(n4797), .ZN(n4794) );
  INV_X1 U5429 ( .A(n4797), .ZN(n4795) );
  NAND2_X1 U5430 ( .A1(n6730), .A2(n4631), .ZN(n4630) );
  OR2_X1 U5431 ( .A1(n7138), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n4631) );
  NOR2_X1 U5432 ( .A1(n10419), .A2(n10418), .ZN(n10417) );
  NAND2_X1 U5433 ( .A1(n7110), .A2(n7111), .ZN(n7420) );
  NAND2_X1 U5434 ( .A1(n7489), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4790) );
  NOR2_X1 U5435 ( .A1(n9878), .A2(n9879), .ZN(n9902) );
  INV_X1 U5436 ( .A(n4784), .ZN(n4782) );
  OAI21_X1 U5437 ( .B1(n9675), .B2(n5133), .A(n4480), .ZN(n8177) );
  NAND2_X1 U5438 ( .A1(n5133), .A2(n5684), .ZN(n4770) );
  INV_X1 U5439 ( .A(n4874), .ZN(n4872) );
  OAI21_X1 U5440 ( .B1(n8499), .B2(n4876), .A(n4875), .ZN(n4874) );
  NOR2_X1 U5441 ( .A1(n8535), .A2(n4877), .ZN(n4876) );
  NAND2_X1 U5442 ( .A1(n8499), .A2(n8498), .ZN(n4875) );
  AND2_X1 U5443 ( .A1(n4452), .A2(n10117), .ZN(n4870) );
  OR2_X1 U5444 ( .A1(n9985), .A2(n7050), .ZN(n8131) );
  NAND2_X1 U5445 ( .A1(n10004), .A2(n10023), .ZN(n4544) );
  INV_X1 U5446 ( .A(n4866), .ZN(n4863) );
  NAND2_X1 U5447 ( .A1(n4866), .A2(n8484), .ZN(n4864) );
  INV_X1 U5448 ( .A(n8484), .ZN(n4865) );
  AOI21_X1 U5449 ( .B1(n4832), .B2(n4830), .A(n4445), .ZN(n4829) );
  INV_X1 U5450 ( .A(n8455), .ZN(n4830) );
  INV_X1 U5451 ( .A(n4832), .ZN(n4831) );
  NAND2_X1 U5452 ( .A1(n4887), .A2(n4889), .ZN(n10061) );
  NAND2_X1 U5453 ( .A1(n4888), .A2(n8344), .ZN(n4887) );
  NOR2_X1 U5455 ( .A1(n10077), .A2(n4891), .ZN(n4890) );
  INV_X1 U5456 ( .A(n8476), .ZN(n4891) );
  NAND2_X1 U5457 ( .A1(n8475), .A2(n4390), .ZN(n4892) );
  INV_X1 U5458 ( .A(n8451), .ZN(n10077) );
  OR2_X1 U5459 ( .A1(n7973), .A2(n7958), .ZN(n7974) );
  NOR2_X1 U5460 ( .A1(n7867), .A2(n4915), .ZN(n4493) );
  INV_X1 U5461 ( .A(n4841), .ZN(n4840) );
  OAI21_X1 U5462 ( .B1(n10137), .B2(n9760), .A(n8449), .ZN(n4841) );
  NAND2_X1 U5463 ( .A1(n7620), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7973) );
  AND2_X1 U5464 ( .A1(n7507), .A2(n9848), .ZN(n7508) );
  NAND2_X1 U5465 ( .A1(n4403), .A2(n6926), .ZN(n6930) );
  NAND2_X1 U5466 ( .A1(n4500), .A2(n6448), .ZN(n6587) );
  OR2_X1 U5467 ( .A1(n8434), .A2(n8929), .ZN(n10182) );
  OR2_X1 U5468 ( .A1(n8434), .A2(n6451), .ZN(n10184) );
  INV_X1 U5469 ( .A(n10117), .ZN(n10179) );
  INV_X1 U5470 ( .A(n10184), .ZN(n10148) );
  NAND2_X1 U5471 ( .A1(n7913), .A2(n7912), .ZN(n10201) );
  AND2_X1 U5472 ( .A1(n8540), .A2(n8539), .ZN(n10208) );
  NAND2_X1 U5473 ( .A1(n7898), .A2(n7910), .ZN(n7901) );
  INV_X1 U5474 ( .A(n10218), .ZN(n4503) );
  NAND2_X1 U5475 ( .A1(n7894), .A2(n7910), .ZN(n7897) );
  OR2_X1 U5476 ( .A1(n6610), .A2(n8286), .ZN(n10456) );
  CLKBUF_X1 U5477 ( .A(n6371), .Z(n6024) );
  XNOR2_X1 U5478 ( .A(n5644), .B(n5643), .ZN(n7907) );
  NAND2_X1 U5479 ( .A1(n4490), .A2(n4429), .ZN(n5555) );
  NAND2_X1 U5480 ( .A1(n4763), .A2(n4762), .ZN(n4761) );
  AND2_X1 U5481 ( .A1(n5556), .A2(n5540), .ZN(n5554) );
  XNOR2_X1 U5482 ( .A(n6346), .B(P1_IR_REG_20__SCAN_IN), .ZN(n8286) );
  INV_X1 U5483 ( .A(n5430), .ZN(n5419) );
  OAI21_X1 U5484 ( .B1(n4769), .B2(n4407), .A(n4671), .ZN(n5430) );
  NAND2_X1 U5485 ( .A1(n4769), .A2(n4768), .ZN(n5417) );
  NAND2_X1 U5486 ( .A1(n4769), .A2(n5379), .ZN(n5394) );
  AND2_X1 U5487 ( .A1(n6234), .A2(n6233), .ZN(n9864) );
  INV_X1 U5488 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4920) );
  INV_X1 U5489 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4664) );
  OR2_X1 U5490 ( .A1(n6174), .A2(n6218), .ZN(n6278) );
  INV_X1 U5491 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8548) );
  NAND2_X1 U5492 ( .A1(n10375), .A2(n10376), .ZN(n10377) );
  OAI21_X1 U5493 ( .B1(n9125), .B2(n8898), .A(n9105), .ZN(n4821) );
  NAND2_X1 U5494 ( .A1(n4678), .A2(n4682), .ZN(n8899) );
  NAND2_X1 U5495 ( .A1(n9126), .A2(n8871), .ZN(n4678) );
  AND2_X1 U5496 ( .A1(n9326), .A2(n9122), .ZN(n4818) );
  AND2_X1 U5497 ( .A1(n5487), .A2(n5486), .ZN(n9004) );
  AND2_X1 U5498 ( .A1(n5446), .A2(n5445), .ZN(n9500) );
  NAND2_X1 U5499 ( .A1(n5494), .A2(n5493), .ZN(n9414) );
  AND2_X1 U5500 ( .A1(n5596), .A2(n5580), .ZN(n9357) );
  NAND2_X1 U5501 ( .A1(n5170), .A2(n5171), .ZN(n4606) );
  AND3_X1 U5502 ( .A1(n5414), .A2(n5413), .A3(n5412), .ZN(n9499) );
  NAND2_X1 U5503 ( .A1(n5152), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n4590) );
  NAND2_X1 U5504 ( .A1(n9262), .A2(n5460), .ZN(n4591) );
  NAND2_X1 U5505 ( .A1(n6071), .A2(n4382), .ZN(n7085) );
  INV_X1 U5506 ( .A(n9143), .ZN(n9131) );
  OR2_X1 U5507 ( .A1(n9073), .A2(n9531), .ZN(n9145) );
  AND2_X1 U5508 ( .A1(n6103), .A2(n9485), .ZN(n9153) );
  NAND2_X1 U5509 ( .A1(n9252), .A2(n4750), .ZN(n7023) );
  OR2_X1 U5510 ( .A1(n9262), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4750) );
  NOR2_X1 U5511 ( .A1(n7182), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7604) );
  INV_X1 U5512 ( .A(n4991), .ZN(n4990) );
  AND2_X1 U5513 ( .A1(n5697), .A2(n5459), .ZN(n9359) );
  NAND2_X1 U5514 ( .A1(n4564), .A2(n9354), .ZN(n9564) );
  OAI21_X1 U5515 ( .B1(n4568), .B2(n4567), .A(n4565), .ZN(n4564) );
  NAND2_X1 U5516 ( .A1(n5926), .A2(n9352), .ZN(n4567) );
  INV_X1 U5517 ( .A(n9365), .ZN(n4568) );
  NAND2_X1 U5518 ( .A1(n7828), .A2(n5910), .ZN(n9505) );
  INV_X1 U5519 ( .A(n5982), .ZN(n5978) );
  NAND2_X1 U5520 ( .A1(n4497), .A2(n4496), .ZN(n4495) );
  INV_X1 U5521 ( .A(n9555), .ZN(n4496) );
  INV_X1 U5522 ( .A(n9554), .ZN(n4497) );
  OR2_X1 U5523 ( .A1(n9772), .A2(n7050), .ZN(n8081) );
  NAND2_X1 U5524 ( .A1(n9828), .A2(n9823), .ZN(n9751) );
  OR2_X1 U5525 ( .A1(n8459), .A2(n7050), .ZN(n8109) );
  INV_X1 U5526 ( .A(n8444), .ZN(n4512) );
  AND2_X1 U5527 ( .A1(n6193), .A2(n6202), .ZN(n7042) );
  NOR2_X1 U5528 ( .A1(n9891), .A2(n9890), .ZN(n9897) );
  XNOR2_X1 U5529 ( .A(n4638), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9947) );
  NAND2_X1 U5530 ( .A1(n9943), .A2(n4639), .ZN(n4638) );
  OR2_X1 U5531 ( .A1(n9944), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n4639) );
  INV_X1 U5532 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9954) );
  INV_X1 U5533 ( .A(n8177), .ZN(n10193) );
  NAND2_X1 U5534 ( .A1(n7854), .A2(n7853), .ZN(n10197) );
  NAND2_X1 U5535 ( .A1(n6012), .A2(n5996), .ZN(n4937) );
  NAND2_X1 U5536 ( .A1(n6000), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4919) );
  NAND2_X1 U5537 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6188) );
  XNOR2_X1 U5538 ( .A(n10377), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(n10561) );
  NOR2_X1 U5539 ( .A1(n10549), .A2(n4481), .ZN(n10548) );
  NOR2_X1 U5540 ( .A1(n10548), .A2(n10547), .ZN(n10546) );
  INV_X1 U5541 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4660) );
  NAND2_X1 U5542 ( .A1(n4746), .A2(n5828), .ZN(n4745) );
  NAND2_X1 U5543 ( .A1(n5849), .A2(n5716), .ZN(n4746) );
  INV_X1 U5544 ( .A(n8403), .ZN(n4697) );
  AND2_X1 U5545 ( .A1(n4692), .A2(n8305), .ZN(n4691) );
  INV_X1 U5546 ( .A(n8322), .ZN(n4705) );
  NAND2_X1 U5547 ( .A1(n4724), .A2(n4727), .ZN(n5772) );
  NAND2_X1 U5548 ( .A1(n8329), .A2(n4701), .ZN(n4700) );
  INV_X1 U5549 ( .A(n4702), .ZN(n4701) );
  INV_X1 U5550 ( .A(n5801), .ZN(n4742) );
  AOI21_X1 U5551 ( .B1(n4711), .B2(n4712), .A(n4539), .ZN(n8363) );
  INV_X1 U5552 ( .A(n4713), .ZN(n4712) );
  NAND2_X1 U5553 ( .A1(n4440), .A2(n5828), .ZN(n4736) );
  NAND2_X1 U5554 ( .A1(n5810), .A2(n5841), .ZN(n4731) );
  NAND2_X1 U5555 ( .A1(n4612), .A2(n4727), .ZN(n4611) );
  NOR2_X1 U5556 ( .A1(n4613), .A2(n7686), .ZN(n4612) );
  NAND2_X1 U5557 ( .A1(n4614), .A2(n5900), .ZN(n4613) );
  NOR2_X1 U5558 ( .A1(n4513), .A2(n7669), .ZN(n4614) );
  NOR2_X1 U5559 ( .A1(n5850), .A2(n4603), .ZN(n5852) );
  INV_X1 U5560 ( .A(n5849), .ZN(n5031) );
  NAND2_X1 U5561 ( .A1(n5008), .A2(n4996), .ZN(n5007) );
  NAND2_X1 U5562 ( .A1(n5694), .A2(n5879), .ZN(n5020) );
  OR2_X1 U5563 ( .A1(n5914), .A2(n5913), .ZN(n5916) );
  NOR2_X1 U5564 ( .A1(n8742), .A2(n9256), .ZN(n4658) );
  NOR2_X1 U5565 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5057) );
  AND2_X1 U5566 ( .A1(n5404), .A2(n5054), .ZN(n4807) );
  NAND2_X1 U5567 ( .A1(n4900), .A2(n4897), .ZN(n4896) );
  INV_X1 U5568 ( .A(n4903), .ZN(n4897) );
  OR2_X1 U5569 ( .A1(n8462), .A2(n8463), .ZN(n4905) );
  NAND2_X1 U5570 ( .A1(n7614), .A2(n9847), .ZN(n7630) );
  AND2_X1 U5571 ( .A1(n5511), .A2(n5514), .ZN(n5515) );
  AOI21_X1 U5572 ( .B1(n4671), .B2(n4407), .A(n4669), .ZN(n4668) );
  INV_X1 U5573 ( .A(n5429), .ZN(n4669) );
  OAI21_X1 U5574 ( .B1(n6398), .B2(n4517), .A(n4516), .ZN(n5238) );
  INV_X1 U5575 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n4517) );
  NAND2_X1 U5576 ( .A1(n6398), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n4516) );
  INV_X1 U5577 ( .A(n5440), .ZN(n5439) );
  NOR2_X1 U5578 ( .A1(n6163), .A2(n4653), .ZN(n4652) );
  INV_X1 U5579 ( .A(n5368), .ZN(n5366) );
  NOR2_X1 U5580 ( .A1(n9147), .A2(n5367), .ZN(n4655) );
  NOR2_X1 U5581 ( .A1(n5855), .A2(n4607), .ZN(n5856) );
  NAND2_X1 U5582 ( .A1(n4616), .A2(n4608), .ZN(n4607) );
  INV_X1 U5583 ( .A(n9439), .ZN(n4616) );
  NOR2_X1 U5584 ( .A1(n4622), .A2(n9336), .ZN(n4621) );
  NAND2_X1 U5585 ( .A1(n9319), .A2(n4659), .ZN(n4622) );
  NAND2_X1 U5586 ( .A1(n5366), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5388) );
  NOR2_X1 U5587 ( .A1(n9341), .A2(n4955), .ZN(n4954) );
  NAND2_X1 U5588 ( .A1(n5972), .A2(n9642), .ZN(n4955) );
  NOR2_X1 U5589 ( .A1(n4981), .A2(n4412), .ZN(n4980) );
  INV_X1 U5590 ( .A(n4986), .ZN(n4981) );
  AND2_X1 U5591 ( .A1(n9420), .A2(n9424), .ZN(n5503) );
  NOR2_X1 U5592 ( .A1(n5524), .A2(n5523), .ZN(n4649) );
  OR2_X1 U5593 ( .A1(n9433), .A2(n9004), .ZN(n9420) );
  NAND2_X1 U5594 ( .A1(n9497), .A2(n9504), .ZN(n9474) );
  NAND2_X1 U5595 ( .A1(n5439), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5463) );
  OR2_X1 U5596 ( .A1(n9512), .A2(n9479), .ZN(n9473) );
  AND2_X1 U5597 ( .A1(n5748), .A2(n5747), .ZN(n5900) );
  INV_X1 U5598 ( .A(n5297), .ZN(n5296) );
  NAND2_X1 U5599 ( .A1(n5892), .A2(n5891), .ZN(n5894) );
  AND2_X1 U5600 ( .A1(n4958), .A2(n10508), .ZN(n4957) );
  INV_X1 U5601 ( .A(n7449), .ZN(n4958) );
  INV_X1 U5602 ( .A(n5201), .ZN(n4651) );
  INV_X1 U5603 ( .A(n5887), .ZN(n4976) );
  NAND3_X1 U5604 ( .A1(n4822), .A2(n8962), .A3(n6878), .ZN(n5959) );
  OR2_X1 U5605 ( .A1(n5931), .A2(n6878), .ZN(n7318) );
  NAND2_X1 U5606 ( .A1(n5223), .A2(n5736), .ZN(n7436) );
  NAND2_X1 U5607 ( .A1(n5032), .A2(n5849), .ZN(n7330) );
  NAND2_X1 U5608 ( .A1(n7330), .A2(n7331), .ZN(n7476) );
  CLKBUF_X1 U5609 ( .A(n5402), .Z(n5405) );
  OR2_X1 U5610 ( .A1(n5313), .A2(n5312), .ZN(n5332) );
  NOR2_X1 U5611 ( .A1(n5196), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n4599) );
  NAND2_X1 U5612 ( .A1(n4931), .A2(n4932), .ZN(n4930) );
  INV_X1 U5613 ( .A(n8009), .ZN(n4931) );
  NOR2_X1 U5614 ( .A1(n4428), .A2(n4927), .ZN(n4926) );
  NOR2_X1 U5615 ( .A1(n8009), .A2(n4928), .ZN(n4927) );
  NAND2_X1 U5616 ( .A1(n4929), .A2(n4932), .ZN(n4928) );
  INV_X1 U5617 ( .A(n9964), .ZN(n8507) );
  AND2_X1 U5618 ( .A1(n8379), .A2(n8378), .ZN(n8386) );
  INV_X1 U5619 ( .A(n8498), .ZN(n4877) );
  AND2_X1 U5620 ( .A1(n8072), .A2(n8071), .ZN(n8100) );
  NAND2_X1 U5621 ( .A1(n10222), .A2(n9993), .ZN(n8493) );
  OR2_X1 U5622 ( .A1(n8485), .A2(n4867), .ZN(n4866) );
  INV_X1 U5623 ( .A(n8482), .ZN(n4867) );
  OR2_X1 U5624 ( .A1(n8030), .A2(n8029), .ZN(n8052) );
  AND2_X1 U5625 ( .A1(n7990), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8012) );
  NOR2_X1 U5626 ( .A1(n7974), .A2(n8634), .ZN(n7990) );
  NAND2_X1 U5627 ( .A1(n4916), .A2(n10161), .ZN(n4915) );
  NOR2_X2 U5628 ( .A1(n7622), .A2(n7621), .ZN(n7620) );
  NOR2_X1 U5629 ( .A1(n10283), .A2(n10288), .ZN(n4916) );
  NOR2_X1 U5630 ( .A1(n8232), .A2(n4901), .ZN(n4900) );
  NOR2_X1 U5631 ( .A1(n4910), .A2(n10301), .ZN(n4909) );
  INV_X1 U5632 ( .A(n4911), .ZN(n4910) );
  NOR2_X1 U5633 ( .A1(n7485), .A2(n8205), .ZN(n4901) );
  NAND2_X1 U5634 ( .A1(n7460), .A2(n4903), .ZN(n4902) );
  NOR2_X1 U5635 ( .A1(n10305), .A2(n7377), .ZN(n4911) );
  AND2_X1 U5636 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6565) );
  OR2_X1 U5637 ( .A1(n7852), .A2(n6397), .ZN(n6401) );
  OR2_X1 U5638 ( .A1(n6516), .A2(n6399), .ZN(n6400) );
  NAND2_X1 U5639 ( .A1(n8370), .A2(n8498), .ZN(n8532) );
  AND2_X1 U5640 ( .A1(n8507), .A2(n8505), .ZN(n4854) );
  AOI21_X1 U5641 ( .B1(n4775), .B2(n4402), .A(n4771), .ZN(n5624) );
  OAI21_X1 U5642 ( .B1(n4773), .B2(n4772), .A(n5608), .ZN(n4771) );
  INV_X1 U5643 ( .A(n5534), .ZN(n4762) );
  NAND2_X1 U5644 ( .A1(n4936), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6346) );
  AND2_X1 U5645 ( .A1(n5996), .A2(n4935), .ZN(n4934) );
  INV_X1 U5646 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4935) );
  NAND2_X1 U5647 ( .A1(n4675), .A2(n4674), .ZN(n5491) );
  AND2_X1 U5648 ( .A1(n5452), .A2(n5473), .ZN(n4674) );
  NAND2_X1 U5649 ( .A1(n5399), .A2(SI_16_), .ZN(n5418) );
  NAND2_X1 U5650 ( .A1(n5378), .A2(SI_14_), .ZN(n5379) );
  AND2_X1 U5651 ( .A1(n5992), .A2(n5991), .ZN(n6001) );
  AND2_X1 U5652 ( .A1(n5348), .A2(n5347), .ZN(n5349) );
  NOR2_X1 U5653 ( .A1(n5346), .A2(n5345), .ZN(n5348) );
  AOI21_X1 U5654 ( .B1(n5355), .B2(n5354), .A(n5353), .ZN(n5356) );
  INV_X1 U5655 ( .A(n5351), .ZN(n5354) );
  INV_X1 U5656 ( .A(n5346), .ZN(n5355) );
  NAND2_X1 U5657 ( .A1(n5255), .A2(SI_9_), .ZN(n4489) );
  NAND2_X1 U5658 ( .A1(n5269), .A2(n5244), .ZN(n5249) );
  INV_X1 U5659 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4661) );
  NAND2_X1 U5660 ( .A1(n8854), .A2(n4425), .ZN(n9000) );
  AND2_X1 U5661 ( .A1(n6134), .A2(n6132), .ZN(n9010) );
  NAND2_X1 U5662 ( .A1(n5366), .A2(n4655), .ZN(n5410) );
  OR2_X1 U5663 ( .A1(n5424), .A2(n9271), .ZN(n5440) );
  NAND2_X1 U5664 ( .A1(n4804), .A2(n4805), .ZN(n4665) );
  NAND2_X1 U5665 ( .A1(n4649), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U5666 ( .A1(n4673), .A2(n9002), .ZN(n9095) );
  INV_X1 U5667 ( .A(n9000), .ZN(n4673) );
  NAND2_X1 U5668 ( .A1(n5827), .A2(n4422), .ZN(n5829) );
  AND2_X1 U5669 ( .A1(n9638), .A2(n9155), .ZN(n5839) );
  NAND2_X1 U5670 ( .A1(n5017), .A2(n8923), .ZN(n5016) );
  AND2_X1 U5671 ( .A1(n5019), .A2(n9359), .ZN(n5015) );
  OAI21_X1 U5672 ( .B1(n5017), .B2(n9359), .A(n5012), .ZN(n5011) );
  NAND2_X1 U5673 ( .A1(n5017), .A2(n5013), .ZN(n5012) );
  NAND2_X1 U5674 ( .A1(n5014), .A2(n8923), .ZN(n5013) );
  INV_X1 U5675 ( .A(n5019), .ZN(n5014) );
  AOI21_X1 U5676 ( .B1(n9327), .B2(n5654), .A(n5620), .ZN(n9129) );
  AND2_X1 U5677 ( .A1(n5567), .A2(n5566), .ZN(n8983) );
  AND4_X1 U5678 ( .A1(n5207), .A2(n5206), .A3(n5205), .A4(n5204), .ZN(n7439)
         );
  NOR2_X2 U5679 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5153) );
  AND2_X1 U5680 ( .A1(n4748), .A2(n4747), .ZN(n9240) );
  INV_X1 U5681 ( .A(n9226), .ZN(n4747) );
  NOR2_X1 U5682 ( .A1(n7021), .A2(n4749), .ZN(n6764) );
  AND2_X1 U5683 ( .A1(n6800), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4749) );
  NAND2_X1 U5684 ( .A1(n9268), .A2(n4752), .ZN(n8914) );
  NAND2_X1 U5685 ( .A1(n8908), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4752) );
  NOR2_X1 U5686 ( .A1(n9677), .A2(n5061), .ZN(n4963) );
  AND2_X1 U5687 ( .A1(n4954), .A2(n5001), .ZN(n9301) );
  NOR2_X1 U5688 ( .A1(n4994), .A2(n9353), .ZN(n4992) );
  OAI21_X1 U5689 ( .B1(n4994), .B2(n5004), .A(n4993), .ZN(n4991) );
  AOI21_X1 U5690 ( .B1(n4995), .B2(n5000), .A(n4397), .ZN(n4993) );
  NAND2_X1 U5691 ( .A1(n7907), .A2(n4378), .ZN(n5630) );
  AND2_X1 U5692 ( .A1(n9334), .A2(n5604), .ZN(n5605) );
  NOR2_X1 U5693 ( .A1(n4566), .A2(n9442), .ZN(n4565) );
  AND2_X1 U5694 ( .A1(n9412), .A2(n4960), .ZN(n9367) );
  OAI21_X1 U5695 ( .B1(n5508), .B2(n4559), .A(n4557), .ZN(n9351) );
  INV_X1 U5696 ( .A(n4558), .ZN(n4557) );
  OAI21_X1 U5697 ( .B1(n4389), .B2(n4559), .A(n5806), .ZN(n4558) );
  INV_X1 U5698 ( .A(n5553), .ZN(n4559) );
  NAND2_X1 U5699 ( .A1(n9412), .A2(n4962), .ZN(n9381) );
  OR2_X1 U5700 ( .A1(n5496), .A2(n5495), .ZN(n5524) );
  INV_X1 U5701 ( .A(n4649), .ZN(n5544) );
  NAND2_X1 U5702 ( .A1(n9412), .A2(n4988), .ZN(n9400) );
  AND2_X1 U5703 ( .A1(n9507), .A2(n4399), .ZN(n9432) );
  NAND2_X1 U5704 ( .A1(n9507), .A2(n4952), .ZN(n9454) );
  AND2_X1 U5705 ( .A1(n5789), .A2(n9419), .ZN(n9461) );
  NAND2_X1 U5706 ( .A1(n9507), .A2(n9665), .ZN(n9483) );
  AND2_X1 U5707 ( .A1(n9473), .A2(n5779), .ZN(n9504) );
  NAND2_X1 U5708 ( .A1(n4488), .A2(n5907), .ZN(n7797) );
  NAND2_X1 U5709 ( .A1(n7765), .A2(n5375), .ZN(n7763) );
  NAND2_X1 U5710 ( .A1(n5024), .A2(n5342), .ZN(n7765) );
  INV_X1 U5711 ( .A(n7743), .ZN(n5024) );
  AND2_X1 U5712 ( .A1(n7750), .A2(n9092), .ZN(n7769) );
  INV_X1 U5713 ( .A(n5900), .ZN(n7546) );
  NAND2_X1 U5714 ( .A1(n4950), .A2(n4949), .ZN(n7690) );
  INV_X1 U5715 ( .A(n5894), .ZN(n7665) );
  NAND2_X1 U5716 ( .A1(n7714), .A2(n5743), .ZN(n7670) );
  OR2_X1 U5717 ( .A1(n5260), .A2(n5259), .ZN(n5284) );
  NAND2_X1 U5718 ( .A1(n7725), .A2(n4957), .ZN(n4956) );
  NAND2_X1 U5719 ( .A1(n7715), .A2(n7716), .ZN(n7714) );
  NAND2_X1 U5720 ( .A1(n7438), .A2(n5738), .ZN(n7715) );
  NAND2_X1 U5721 ( .A1(n4651), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5225) );
  INV_X1 U5722 ( .A(n7472), .ZN(n7474) );
  NAND2_X1 U5723 ( .A1(n7474), .A2(n10508), .ZN(n7473) );
  INV_X1 U5724 ( .A(n5851), .ZN(n7477) );
  NAND2_X1 U5725 ( .A1(n5181), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5201) );
  INV_X1 U5726 ( .A(n5182), .ZN(n5181) );
  NAND2_X1 U5727 ( .A1(n7531), .A2(n10501), .ZN(n7472) );
  AND2_X1 U5728 ( .A1(n7530), .A2(n10496), .ZN(n7531) );
  NAND3_X1 U5729 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5182) );
  NAND2_X1 U5730 ( .A1(n9176), .A2(n8834), .ZN(n7525) );
  NAND2_X1 U5731 ( .A1(n6824), .A2(n5713), .ZN(n6841) );
  OR2_X1 U5732 ( .A1(n9538), .A2(n8923), .ZN(n6104) );
  OR2_X1 U5733 ( .A1(n5548), .A2(n6756), .ZN(n5106) );
  NAND2_X1 U5734 ( .A1(n9519), .A2(n5884), .ZN(n6823) );
  INV_X1 U5735 ( .A(n8835), .ZN(n8880) );
  NAND2_X1 U5736 ( .A1(n5938), .A2(n5937), .ZN(n5939) );
  INV_X1 U5737 ( .A(n7337), .ZN(n10501) );
  NAND2_X1 U5738 ( .A1(n6768), .A2(n10480), .ZN(n10467) );
  AND2_X1 U5739 ( .A1(n5281), .A2(n5293), .ZN(n6796) );
  OAI21_X1 U5740 ( .B1(n5313), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5277) );
  NAND2_X1 U5741 ( .A1(n4599), .A2(n4598), .ZN(n5313) );
  INV_X1 U5742 ( .A(n4599), .ZN(n5218) );
  NAND2_X1 U5743 ( .A1(n5113), .A2(n5081), .ZN(n5166) );
  AND2_X1 U5744 ( .A1(n6896), .A2(n6895), .ZN(n7211) );
  AND2_X1 U5745 ( .A1(n8048), .A2(n8049), .ZN(n9728) );
  INV_X1 U5746 ( .A(n8117), .ZN(n9699) );
  OAI21_X1 U5747 ( .B1(n9751), .B2(n4930), .A(n4926), .ZN(n9782) );
  NAND2_X1 U5748 ( .A1(n4584), .A2(n4421), .ZN(n8063) );
  AND2_X1 U5749 ( .A1(n4922), .A2(n8069), .ZN(n4515) );
  AND2_X1 U5750 ( .A1(n6702), .A2(n6701), .ZN(n6882) );
  INV_X1 U5751 ( .A(n7951), .ZN(n4947) );
  NAND2_X1 U5752 ( .A1(n8437), .A2(n8438), .ZN(n4537) );
  OR2_X1 U5753 ( .A1(n8433), .A2(n8435), .ZN(n4538) );
  AND2_X1 U5754 ( .A1(n8193), .A2(n8192), .ZN(n8947) );
  AND3_X1 U5755 ( .A1(n7236), .A2(n7235), .A3(n7234), .ZN(n7506) );
  OR2_X1 U5756 ( .A1(n6707), .A2(n4642), .ZN(n6387) );
  NAND2_X1 U5757 ( .A1(n6572), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6369) );
  AND2_X1 U5758 ( .A1(n10422), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4520) );
  NAND2_X1 U5759 ( .A1(n4628), .A2(n4627), .ZN(n6733) );
  OR2_X1 U5760 ( .A1(n10422), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4627) );
  NAND2_X1 U5761 ( .A1(n4630), .A2(n4629), .ZN(n4628) );
  INV_X1 U5762 ( .A(n10425), .ZN(n4629) );
  NAND2_X1 U5763 ( .A1(n6733), .A2(n6732), .ZN(n7109) );
  NAND2_X1 U5764 ( .A1(n7420), .A2(n4468), .ZN(n7421) );
  NAND2_X1 U5765 ( .A1(n7421), .A2(n7422), .ZN(n9860) );
  OR2_X1 U5766 ( .A1(n7117), .A2(n7118), .ZN(n4791) );
  NAND2_X1 U5767 ( .A1(n9860), .A2(n4623), .ZN(n9874) );
  OR2_X1 U5768 ( .A1(n9864), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n4623) );
  NOR2_X1 U5769 ( .A1(n9925), .A2(n4640), .ZN(n9926) );
  AND2_X1 U5770 ( .A1(n9932), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n4640) );
  NAND2_X1 U5771 ( .A1(n9926), .A2(n9927), .ZN(n9943) );
  NOR2_X1 U5772 ( .A1(n4856), .A2(n4851), .ZN(n4850) );
  INV_X1 U5773 ( .A(n8506), .ZN(n4851) );
  INV_X1 U5774 ( .A(n4854), .ZN(n4853) );
  INV_X1 U5775 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5259) );
  OR2_X1 U5776 ( .A1(n10222), .A2(n9993), .ZN(n9988) );
  NOR2_X2 U5777 ( .A1(n10005), .A2(n10222), .ZN(n9980) );
  AND2_X1 U5778 ( .A1(n9988), .A2(n8493), .ZN(n8488) );
  AND2_X1 U5779 ( .A1(n8094), .A2(n8093), .ZN(n10004) );
  AND2_X1 U5780 ( .A1(n8487), .A2(n8359), .ZN(n9999) );
  NAND2_X1 U5781 ( .A1(n8456), .A2(n10013), .ZN(n10024) );
  NAND2_X1 U5782 ( .A1(n4912), .A2(n4834), .ZN(n10050) );
  NOR2_X1 U5783 ( .A1(n10050), .A2(n10237), .ZN(n10032) );
  OAI21_X1 U5784 ( .B1(n10061), .B2(n8481), .A(n8480), .ZN(n10046) );
  NAND2_X1 U5785 ( .A1(n8012), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n8030) );
  AND2_X1 U5786 ( .A1(n7999), .A2(n7998), .ZN(n10063) );
  NAND2_X1 U5787 ( .A1(n10097), .A2(n10087), .ZN(n10081) );
  AND2_X1 U5788 ( .A1(n10109), .A2(n10099), .ZN(n10097) );
  NAND2_X1 U5789 ( .A1(n8475), .A2(n8474), .ZN(n10114) );
  AND2_X1 U5790 ( .A1(n7983), .A2(n7982), .ZN(n10131) );
  AND2_X1 U5791 ( .A1(n8332), .A2(n8471), .ZN(n10128) );
  NOR2_X1 U5792 ( .A1(n7635), .A2(n4914), .ZN(n10167) );
  INV_X1 U5793 ( .A(n4916), .ZN(n4914) );
  NOR2_X1 U5794 ( .A1(n7635), .A2(n10288), .ZN(n10166) );
  AND2_X1 U5795 ( .A1(n8465), .A2(n8461), .ZN(n10176) );
  AND2_X1 U5796 ( .A1(n8468), .A2(n10177), .ZN(n8273) );
  INV_X1 U5797 ( .A(n8273), .ZN(n8445) );
  INV_X1 U5798 ( .A(n8270), .ZN(n7615) );
  NAND2_X1 U5799 ( .A1(n4902), .A2(n4899), .ZN(n7631) );
  INV_X1 U5800 ( .A(n4901), .ZN(n4899) );
  AND3_X1 U5801 ( .A1(n7264), .A2(n7263), .A3(n7262), .ZN(n7628) );
  OR2_X1 U5802 ( .A1(n7246), .A2(n4847), .ZN(n4846) );
  INV_X1 U5803 ( .A(n4845), .ZN(n4844) );
  INV_X1 U5804 ( .A(n7141), .ZN(n4847) );
  NAND2_X1 U5805 ( .A1(n4499), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7052) );
  INV_X1 U5806 ( .A(n6903), .ZN(n4499) );
  NAND2_X1 U5807 ( .A1(n7047), .A2(n4911), .ZN(n7464) );
  NAND2_X1 U5808 ( .A1(n4881), .A2(n8227), .ZN(n4880) );
  AND2_X1 U5809 ( .A1(n4885), .A2(n8227), .ZN(n4879) );
  NAND2_X1 U5810 ( .A1(n7142), .A2(n7141), .ZN(n7247) );
  NAND2_X1 U5811 ( .A1(n4884), .A2(n8298), .ZN(n7062) );
  AND2_X1 U5812 ( .A1(n4884), .A2(n4883), .ZN(n7144) );
  INV_X1 U5813 ( .A(n4881), .ZN(n4883) );
  NAND2_X1 U5814 ( .A1(n7047), .A2(n7290), .ZN(n7163) );
  NAND2_X1 U5815 ( .A1(n7003), .A2(n8225), .ZN(n7006) );
  NAND2_X1 U5816 ( .A1(n6748), .A2(n8401), .ZN(n7003) );
  NAND2_X1 U5817 ( .A1(n6933), .A2(n8403), .ZN(n8291) );
  OR2_X1 U5818 ( .A1(n6930), .A2(n7368), .ZN(n7001) );
  NAND2_X1 U5819 ( .A1(n4706), .A2(n4707), .ZN(n8296) );
  INV_X1 U5820 ( .A(n4708), .ZN(n4707) );
  OAI21_X1 U5821 ( .B1(n8399), .B2(n4709), .A(n8400), .ZN(n4708) );
  CLKBUF_X1 U5822 ( .A(n7036), .Z(n6998) );
  NAND2_X1 U5823 ( .A1(n6565), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6637) );
  NOR2_X1 U5824 ( .A1(n6678), .A2(n7399), .ZN(n4907) );
  NAND2_X1 U5825 ( .A1(n4710), .A2(n8399), .ZN(n6748) );
  NAND2_X1 U5826 ( .A1(n8408), .A2(n8261), .ZN(n4710) );
  NAND2_X1 U5827 ( .A1(n8262), .A2(n6672), .ZN(n6742) );
  INV_X1 U5828 ( .A(n6671), .ZN(n6672) );
  NAND2_X1 U5829 ( .A1(n6592), .A2(n6591), .ZN(n8220) );
  NAND2_X1 U5830 ( .A1(n7889), .A2(n7910), .ZN(n7892) );
  NAND2_X1 U5831 ( .A1(n7860), .A2(n7859), .ZN(n10277) );
  INV_X1 U5832 ( .A(n6928), .ZN(n6932) );
  OR2_X1 U5833 ( .A1(n8388), .A2(n8286), .ZN(n10311) );
  INV_X1 U5834 ( .A(n10456), .ZN(n10307) );
  INV_X1 U5835 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6355) );
  XNOR2_X1 U5836 ( .A(n5688), .B(n5687), .ZN(n9675) );
  XNOR2_X1 U5837 ( .A(n5678), .B(n5661), .ZN(n8931) );
  NAND2_X1 U5838 ( .A1(n6035), .A2(n6034), .ZN(n6362) );
  XNOR2_X1 U5839 ( .A(n5660), .B(n5648), .ZN(n9682) );
  NAND2_X1 U5840 ( .A1(n4778), .A2(n5647), .ZN(n5660) );
  NAND2_X1 U5841 ( .A1(n5644), .A2(n5643), .ZN(n4778) );
  XNOR2_X1 U5842 ( .A(n6362), .B(P1_IR_REG_28__SCAN_IN), .ZN(n6249) );
  XNOR2_X1 U5843 ( .A(n5624), .B(n5623), .ZN(n7903) );
  XNOR2_X1 U5844 ( .A(n5592), .B(n5591), .ZN(n7898) );
  NAND2_X1 U5845 ( .A1(n5610), .A2(n5607), .ZN(n5592) );
  NAND2_X1 U5846 ( .A1(n4774), .A2(n4773), .ZN(n5610) );
  NAND2_X1 U5847 ( .A1(n6021), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U5848 ( .A1(n4774), .A2(n5571), .ZN(n5585) );
  NAND2_X1 U5849 ( .A1(n6013), .A2(n6029), .ZN(n6021) );
  INV_X1 U5850 ( .A(n6019), .ZN(n6013) );
  AOI21_X1 U5851 ( .B1(n5474), .B2(n4766), .A(n4763), .ZN(n5535) );
  NAND2_X1 U5852 ( .A1(n5290), .A2(n4666), .ZN(n5291) );
  NAND2_X1 U5853 ( .A1(n5132), .A2(n4689), .ZN(n4688) );
  INV_X1 U5854 ( .A(n5134), .ZN(n4690) );
  INV_X1 U5855 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10358) );
  NOR2_X1 U5856 ( .A1(n10365), .A2(n10364), .ZN(n10366) );
  NOR2_X1 U5857 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10553), .ZN(n10367) );
  AND4_X1 U5858 ( .A1(n5341), .A2(n5340), .A3(n5339), .A4(n5338), .ZN(n8975)
         );
  NAND2_X1 U5859 ( .A1(n5542), .A2(n5541), .ZN(n9383) );
  INV_X1 U5860 ( .A(n6040), .ZN(n7730) );
  AND4_X1 U5861 ( .A1(n5302), .A2(n5301), .A3(n5300), .A4(n5299), .ZN(n9014)
         );
  NAND2_X1 U5862 ( .A1(n4816), .A2(n7514), .ZN(n6099) );
  INV_X1 U5863 ( .A(n4682), .ZN(n4681) );
  AOI21_X1 U5864 ( .B1(n4682), .B2(n8878), .A(n4680), .ZN(n4679) );
  INV_X1 U5865 ( .A(n8879), .ZN(n4680) );
  INV_X1 U5866 ( .A(n4809), .ZN(n4808) );
  OAI21_X1 U5867 ( .B1(n4382), .B2(n4386), .A(n4438), .ZN(n4809) );
  AND2_X1 U5868 ( .A1(n6048), .A2(n6049), .ZN(n6973) );
  NAND2_X1 U5869 ( .A1(n6973), .A2(n6972), .ZN(n6971) );
  NAND2_X1 U5870 ( .A1(n4803), .A2(n4802), .ZN(n6972) );
  INV_X1 U5871 ( .A(n9566), .ZN(n9030) );
  NAND2_X1 U5872 ( .A1(n5409), .A2(n5408), .ZN(n9047) );
  NAND2_X1 U5873 ( .A1(n4804), .A2(n4805), .ZN(n8858) );
  OAI21_X1 U5874 ( .B1(n9037), .B2(n6151), .A(n6150), .ZN(n9050) );
  NAND2_X1 U5875 ( .A1(n5559), .A2(n5558), .ZN(n9570) );
  AND4_X1 U5876 ( .A1(n5323), .A2(n5322), .A3(n5321), .A4(n5320), .ZN(n9086)
         );
  AND4_X1 U5877 ( .A1(n5289), .A2(n5288), .A3(n5287), .A4(n5286), .ZN(n7785)
         );
  AOI21_X1 U5878 ( .B1(n4814), .B2(n7515), .A(n4812), .ZN(n4811) );
  INV_X1 U5879 ( .A(n4814), .ZN(n4813) );
  NAND2_X1 U5880 ( .A1(n4800), .A2(n6049), .ZN(n8817) );
  AND2_X1 U5881 ( .A1(n5470), .A2(n5469), .ZN(n9480) );
  AND2_X1 U5882 ( .A1(n6071), .A2(n6862), .ZN(n7086) );
  NAND2_X1 U5883 ( .A1(n9126), .A2(n9127), .ZN(n4529) );
  OR2_X1 U5884 ( .A1(n5860), .A2(n5879), .ZN(n4735) );
  XNOR2_X1 U5885 ( .A(n4617), .B(n8923), .ZN(n5860) );
  AOI21_X1 U5886 ( .B1(n9357), .B2(n5654), .A(n5583), .ZN(n9128) );
  INV_X1 U5887 ( .A(n8983), .ZN(n9160) );
  INV_X1 U5888 ( .A(n9480), .ZN(n9164) );
  INV_X1 U5889 ( .A(n7100), .ZN(n9175) );
  XNOR2_X1 U5890 ( .A(n5138), .B(P2_IR_REG_1__SCAN_IN), .ZN(n6961) );
  NOR2_X1 U5891 ( .A1(n7079), .A2(n7080), .ZN(n9183) );
  INV_X1 U5892 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10359) );
  NOR2_X1 U5893 ( .A1(n5154), .A2(n4754), .ZN(n7083) );
  OAI21_X1 U5894 ( .B1(n5153), .B2(n4756), .A(n4755), .ZN(n4754) );
  NAND2_X1 U5895 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4756) );
  NAND2_X1 U5896 ( .A1(n9677), .A2(n5059), .ZN(n4755) );
  OAI21_X1 U5897 ( .B1(n9240), .B2(n9239), .A(n9238), .ZN(n9242) );
  AOI21_X1 U5898 ( .B1(n9242), .B2(n6849), .A(n6848), .ZN(n6860) );
  NOR2_X1 U5899 ( .A1(n7023), .A2(n7022), .ZN(n7021) );
  AND2_X1 U5900 ( .A1(n5384), .A2(n5363), .ZN(n6992) );
  NAND2_X1 U5901 ( .A1(n7181), .A2(n4753), .ZN(n7182) );
  NAND2_X1 U5902 ( .A1(n7180), .A2(n7597), .ZN(n4753) );
  INV_X1 U5903 ( .A(n9295), .ZN(n9258) );
  NAND3_X1 U5904 ( .A1(n7608), .A2(n7606), .A3(n4543), .ZN(n8909) );
  OR2_X1 U5905 ( .A1(n8902), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4543) );
  XNOR2_X1 U5906 ( .A(n8914), .B(n4751), .ZN(n9292) );
  AND2_X1 U5907 ( .A1(n5635), .A2(n9307), .ZN(n8892) );
  NAND2_X1 U5908 ( .A1(n7845), .A2(n8895), .ZN(n9550) );
  NAND2_X1 U5909 ( .A1(n7841), .A2(n4996), .ZN(n7842) );
  NAND2_X1 U5910 ( .A1(n7839), .A2(n7840), .ZN(n7843) );
  XNOR2_X1 U5911 ( .A(n4510), .B(n4996), .ZN(n9553) );
  NAND2_X1 U5912 ( .A1(n4997), .A2(n4999), .ZN(n4510) );
  NAND2_X1 U5913 ( .A1(n4984), .A2(n4985), .ZN(n9380) );
  AND2_X1 U5914 ( .A1(n4984), .A2(n4982), .ZN(n9379) );
  NAND2_X1 U5915 ( .A1(n9411), .A2(n4986), .ZN(n4984) );
  NAND2_X1 U5916 ( .A1(n5508), .A2(n5796), .ZN(n9405) );
  AOI21_X1 U5917 ( .B1(n9411), .B2(n5923), .A(n4396), .ZN(n9398) );
  NAND2_X1 U5918 ( .A1(n4550), .A2(n5775), .ZN(n7823) );
  AND2_X1 U5919 ( .A1(n5387), .A2(n5386), .ZN(n9154) );
  NAND2_X1 U5920 ( .A1(n5021), .A2(n5022), .ZN(n7793) );
  NAND2_X1 U5921 ( .A1(n4972), .A2(n4974), .ZN(n7326) );
  NAND2_X1 U5922 ( .A1(n4973), .A2(n5888), .ZN(n4972) );
  NAND2_X1 U5923 ( .A1(n6809), .A2(n5887), .ZN(n7537) );
  NAND2_X1 U5924 ( .A1(n9536), .A2(n7320), .ZN(n9495) );
  AND2_X1 U5925 ( .A1(n9536), .A2(n7321), .ZN(n9521) );
  NOR2_X1 U5926 ( .A1(n9564), .A2(n4562), .ZN(n9567) );
  OR2_X1 U5927 ( .A1(n9565), .A2(n4563), .ZN(n4562) );
  AND2_X1 U5928 ( .A1(n9566), .A2(n9630), .ZN(n4563) );
  INV_X1 U5929 ( .A(n9414), .ZN(n9657) );
  OR2_X1 U5930 ( .A1(n9609), .A2(n9608), .ZN(n9666) );
  AND2_X1 U5931 ( .A1(n6105), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10480) );
  NAND2_X1 U5932 ( .A1(n5077), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5064) );
  XNOR2_X1 U5933 ( .A(n5294), .B(P2_IR_REG_11__SCAN_IN), .ZN(n9262) );
  INV_X1 U5934 ( .A(n5113), .ZN(n5164) );
  AOI22_X1 U5935 ( .A1(n7873), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n4368), .B2(
        n10409), .ZN(n6886) );
  NAND2_X1 U5936 ( .A1(n6885), .A2(n7902), .ZN(n6887) );
  INV_X1 U5937 ( .A(n8140), .ZN(n4583) );
  OR2_X1 U5938 ( .A1(n9811), .A2(n9812), .ZN(n8140) );
  AND2_X1 U5939 ( .A1(n4392), .A2(n9815), .ZN(n4579) );
  OAI21_X1 U5940 ( .B1(n8163), .B2(n4387), .A(n4426), .ZN(n4577) );
  AND2_X1 U5941 ( .A1(n8946), .A2(n9815), .ZN(n4514) );
  NAND2_X1 U5942 ( .A1(n7907), .A2(n7910), .ZN(n7909) );
  NAND2_X1 U5943 ( .A1(n7880), .A2(n7910), .ZN(n7882) );
  AND3_X1 U5944 ( .A1(n7502), .A2(n7501), .A3(n7500), .ZN(n10183) );
  NAND2_X1 U5945 ( .A1(n4938), .A2(n4942), .ZN(n7646) );
  NAND2_X1 U5946 ( .A1(n7352), .A2(n4943), .ZN(n4938) );
  AND3_X1 U5947 ( .A1(n7945), .A2(n7944), .A3(n7943), .ZN(n10185) );
  CLKBUF_X1 U5948 ( .A(n6745), .Z(n6926) );
  NAND2_X1 U5949 ( .A1(n9751), .A2(n4933), .ZN(n4925) );
  NAND2_X1 U5950 ( .A1(n7863), .A2(n7862), .ZN(n10266) );
  AND2_X1 U5951 ( .A1(n4570), .A2(n6554), .ZN(n4569) );
  INV_X1 U5952 ( .A(n6561), .ZN(n4570) );
  NAND2_X1 U5953 ( .A1(n4571), .A2(n4478), .ZN(n6562) );
  OAI21_X1 U5954 ( .B1(n4942), .B2(n4940), .A(n4439), .ZN(n4939) );
  AND2_X1 U5955 ( .A1(n7156), .A2(n7155), .ZN(n7362) );
  NAND2_X1 U5956 ( .A1(n4941), .A2(n4943), .ZN(n7582) );
  OR2_X1 U5957 ( .A1(n7352), .A2(n5047), .ZN(n4941) );
  OR2_X1 U5958 ( .A1(n7852), .A2(n6417), .ZN(n6421) );
  OAI22_X1 U5959 ( .A1(n7851), .A2(n6649), .B1(n6418), .B2(n6516), .ZN(n6419)
         );
  INV_X1 U5960 ( .A(n9715), .ZN(n9804) );
  NAND2_X1 U5961 ( .A1(n7870), .A2(n7869), .ZN(n10258) );
  INV_X1 U5962 ( .A(n10219), .ZN(n9983) );
  AND3_X1 U5963 ( .A1(n7627), .A2(n7626), .A3(n7625), .ZN(n9830) );
  AND2_X1 U5964 ( .A1(n6385), .A2(n6384), .ZN(n9835) );
  INV_X1 U5965 ( .A(n10063), .ZN(n10094) );
  INV_X1 U5966 ( .A(n10079), .ZN(n10115) );
  AND2_X1 U5967 ( .A1(n6584), .A2(n6583), .ZN(n9760) );
  INV_X1 U5968 ( .A(n7628), .ZN(n9847) );
  INV_X1 U5969 ( .A(n7506), .ZN(n9848) );
  INV_X1 U5970 ( .A(n7362), .ZN(n9849) );
  BUF_X1 U5971 ( .A(P1_U4006), .Z(n9858) );
  NAND2_X1 U5972 ( .A1(n6321), .A2(n6320), .ZN(n10386) );
  NAND2_X1 U5973 ( .A1(n6473), .A2(n6472), .ZN(n6476) );
  NAND2_X1 U5974 ( .A1(n4633), .A2(n4385), .ZN(n10408) );
  OR2_X1 U5975 ( .A1(n6473), .A2(n10405), .ZN(n4633) );
  INV_X1 U5976 ( .A(n4798), .ZN(n10404) );
  NAND2_X1 U5977 ( .A1(n4796), .A2(n4797), .ZN(n6543) );
  AND2_X1 U5978 ( .A1(n4796), .A2(n4416), .ZN(n6542) );
  OR2_X1 U5979 ( .A1(n4798), .A2(n4410), .ZN(n4796) );
  NAND2_X1 U5980 ( .A1(n4632), .A2(n4634), .ZN(n6540) );
  NAND2_X1 U5981 ( .A1(n4385), .A2(n10405), .ZN(n4634) );
  NAND2_X1 U5982 ( .A1(n4793), .A2(n4435), .ZN(n4792) );
  OR2_X1 U5983 ( .A1(n6544), .A2(n4794), .ZN(n4793) );
  INV_X1 U5984 ( .A(n4630), .ZN(n10424) );
  OR2_X1 U5985 ( .A1(n7118), .A2(n7428), .ZN(n4789) );
  XNOR2_X1 U5986 ( .A(n9895), .B(n9889), .ZN(n9890) );
  NOR2_X1 U5987 ( .A1(n9897), .A2(n9896), .ZN(n9900) );
  NOR2_X1 U5988 ( .A1(n9902), .A2(n9903), .ZN(n9905) );
  NAND2_X1 U5989 ( .A1(n4783), .A2(n4784), .ZN(n9914) );
  XNOR2_X1 U5990 ( .A(n10193), .B(n7914), .ZN(n10195) );
  OAI211_X1 U5991 ( .C1(n8536), .C2(n4873), .A(n4871), .B(n4869), .ZN(n4868)
         );
  NAND2_X1 U5992 ( .A1(n4447), .A2(n10117), .ZN(n4873) );
  AOI21_X1 U5993 ( .B1(n4872), .B2(n10117), .A(n8502), .ZN(n4871) );
  AND2_X1 U5994 ( .A1(n8183), .A2(n8143), .ZN(n9973) );
  OR2_X1 U5995 ( .A1(n9969), .A2(n10182), .ZN(n4530) );
  XNOR2_X1 U5996 ( .A(n9962), .B(n9964), .ZN(n10216) );
  INV_X1 U5997 ( .A(n10229), .ZN(n10009) );
  OAI21_X1 U5998 ( .B1(n4504), .B2(n4865), .A(n4408), .ZN(n10017) );
  NAND2_X1 U5999 ( .A1(n4828), .A2(n4829), .ZN(n10031) );
  OR2_X1 U6000 ( .A1(n4518), .A2(n4831), .ZN(n4828) );
  AND2_X1 U6001 ( .A1(n4833), .A2(n4418), .ZN(n10044) );
  NAND2_X1 U6002 ( .A1(n4518), .A2(n8455), .ZN(n4833) );
  NAND2_X1 U6003 ( .A1(n4892), .A2(n8476), .ZN(n10076) );
  INV_X1 U6004 ( .A(n6448), .ZN(n6450) );
  OAI21_X1 U6006 ( .B1(n10199), .B2(n10456), .A(n10198), .ZN(n10315) );
  NOR2_X1 U6007 ( .A1(n10217), .A2(n4501), .ZN(n10220) );
  NAND2_X1 U6008 ( .A1(n4503), .A2(n4502), .ZN(n4501) );
  NAND2_X1 U6009 ( .A1(n10219), .A2(n10306), .ZN(n4502) );
  AND2_X1 U6010 ( .A1(n6024), .A2(n6344), .ZN(n10453) );
  CLKBUF_X1 U6011 ( .A(n6249), .Z(n8929) );
  INV_X1 U6012 ( .A(n9951), .ZN(n10053) );
  NOR2_X1 U6013 ( .A1(n6205), .A2(n6012), .ZN(n7138) );
  NAND2_X1 U6014 ( .A1(n6174), .A2(n4921), .ZN(n6171) );
  INV_X1 U6015 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n8176) );
  AOI22_X1 U6016 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .B1(n6305), .B2(n10358), .ZN(n10567) );
  AND2_X1 U6017 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10366), .ZN(n10553) );
  XOR2_X1 U6018 ( .A(n10368), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10552) );
  NOR2_X1 U6019 ( .A1(n10378), .A2(n10560), .ZN(n10551) );
  NOR2_X1 U6020 ( .A1(n10546), .A2(n4483), .ZN(n10545) );
  NAND2_X1 U6021 ( .A1(n10545), .A2(n10544), .ZN(n10543) );
  OAI21_X1 U6022 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10543), .ZN(n10541) );
  OAI21_X1 U6023 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10540), .ZN(n10538) );
  NAND2_X1 U6024 ( .A1(n10538), .A2(n10539), .ZN(n10537) );
  NAND2_X1 U6025 ( .A1(n10537), .A2(n4521), .ZN(n10535) );
  NAND2_X1 U6026 ( .A1(n4523), .A2(n4522), .ZN(n4521) );
  INV_X1 U6027 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n4522) );
  NAND2_X1 U6028 ( .A1(n7085), .A2(n6077), .ZN(n7099) );
  NOR2_X1 U6029 ( .A1(n8901), .A2(n4818), .ZN(n4817) );
  OR4_X1 U6030 ( .A1(n6168), .A2(n6167), .A3(n6166), .A4(n6165), .ZN(P2_U3221)
         );
  OAI21_X1 U6031 ( .B1(n4528), .B2(n9125), .A(n4526), .ZN(P2_U3242) );
  INV_X1 U6032 ( .A(n4527), .ZN(n4526) );
  NAND2_X1 U6033 ( .A1(n4529), .A2(n9105), .ZN(n4528) );
  OAI21_X1 U6034 ( .B1(n9646), .B2(n9153), .A(n9134), .ZN(n4527) );
  INV_X1 U6035 ( .A(n4548), .ZN(P2_U3557) );
  AOI21_X1 U6036 ( .B1(n9178), .B2(P2_DATAO_REG_5__SCAN_IN), .A(n4549), .ZN(
        n4548) );
  AOI21_X1 U6037 ( .B1(n8924), .B2(n8923), .A(n4541), .ZN(n4540) );
  NAND2_X1 U6038 ( .A1(n8925), .A2(n9359), .ZN(n4542) );
  OAI21_X1 U6039 ( .B1(n8927), .B2(n4660), .A(n8926), .ZN(n4541) );
  MUX2_X1 U6040 ( .A(n5985), .B(n5981), .S(n10519), .Z(n5983) );
  OAI21_X1 U6041 ( .B1(n9640), .B2(n10519), .A(n4486), .ZN(P2_U3547) );
  NOR2_X1 U6042 ( .A1(n4470), .A2(n4487), .ZN(n4486) );
  NOR2_X1 U6043 ( .A1(n10522), .A2(n9557), .ZN(n4487) );
  NAND2_X1 U6044 ( .A1(n9345), .A2(n7701), .ZN(n4485) );
  MUX2_X1 U6045 ( .A(n5985), .B(n5984), .S(n10512), .Z(n5986) );
  AOI21_X1 U6046 ( .B1(n9308), .B2(n5975), .A(n5974), .ZN(n5976) );
  NOR2_X1 U6047 ( .A1(n10513), .A2(n5973), .ZN(n5974) );
  INV_X1 U6048 ( .A(n4507), .ZN(n4506) );
  OAI22_X1 U6049 ( .A1(n9670), .A2(n9642), .B1(n10513), .B2(n9641), .ZN(n4507)
         );
  OAI211_X1 U6050 ( .C1(n9813), .C2(n4580), .A(n4578), .B(n4576), .ZN(P1_U3212) );
  AOI21_X1 U6051 ( .B1(n4579), .B2(n8140), .A(n4577), .ZN(n4576) );
  NAND2_X1 U6052 ( .A1(n4449), .A2(n9815), .ZN(n4580) );
  NAND2_X1 U6053 ( .A1(n9813), .A2(n4579), .ZN(n4578) );
  NAND2_X1 U6054 ( .A1(n4491), .A2(n4512), .ZN(n4511) );
  NAND2_X1 U6055 ( .A1(n6272), .A2(n4646), .ZN(n6274) );
  OAI21_X1 U6056 ( .B1(n9954), .B2(n10431), .A(n9953), .ZN(n4788) );
  AOI211_X1 U6057 ( .C1(n4484), .C2(n10460), .A(n7408), .B(n7407), .ZN(n7409)
         );
  OAI21_X1 U6058 ( .B1(n10350), .B2(n6397), .A(n4644), .ZN(P1_U3352) );
  OAI21_X1 U6059 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n10382), .A(n10556), .ZN(
        n10384) );
  NOR3_X1 U6060 ( .A1(n5746), .A2(n5745), .A3(n5751), .ZN(n4381) );
  AND2_X1 U6061 ( .A1(n4988), .A2(n9005), .ZN(n4384) );
  INV_X2 U6062 ( .A(n6516), .ZN(n7902) );
  INV_X2 U6063 ( .A(n5193), .ZN(n5133) );
  INV_X2 U6064 ( .A(n4376), .ZN(n8940) );
  INV_X1 U6065 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6218) );
  AND2_X1 U6066 ( .A1(n10406), .A2(n4635), .ZN(n4385) );
  OR2_X1 U6067 ( .A1(n8164), .A2(n9825), .ZN(n4387) );
  AND2_X1 U6068 ( .A1(n4829), .A2(n4427), .ZN(n4388) );
  AND2_X1 U6069 ( .A1(n5924), .A2(n5796), .ZN(n4389) );
  AND2_X1 U6070 ( .A1(n8474), .A2(n4893), .ZN(n4390) );
  AND2_X1 U6071 ( .A1(n4626), .A2(n10393), .ZN(n4391) );
  NOR2_X1 U6072 ( .A1(n8162), .A2(n8161), .ZN(n4392) );
  AND2_X1 U6073 ( .A1(n9976), .A2(n9983), .ZN(n4393) );
  OR2_X1 U6074 ( .A1(n9326), .A2(n9129), .ZN(n5819) );
  AND2_X1 U6075 ( .A1(n5356), .A2(n5376), .ZN(n4394) );
  AND2_X1 U6076 ( .A1(n5839), .A2(n5020), .ZN(n4395) );
  NOR2_X1 U6077 ( .A1(n9414), .A2(n9163), .ZN(n4396) );
  AND2_X1 U6078 ( .A1(n5001), .A2(n8881), .ZN(n4397) );
  NAND2_X1 U6079 ( .A1(n5819), .A2(n5822), .ZN(n9315) );
  INV_X1 U6080 ( .A(n10004), .ZN(n10039) );
  AND2_X1 U6081 ( .A1(n5061), .A2(n4966), .ZN(n4398) );
  AND2_X1 U6082 ( .A1(n4951), .A2(n4952), .ZN(n4399) );
  NAND2_X1 U6083 ( .A1(n5630), .A2(n5629), .ZN(n9548) );
  INV_X1 U6084 ( .A(n9548), .ZN(n5001) );
  AND2_X1 U6085 ( .A1(n5737), .A2(n5248), .ZN(n4400) );
  NAND2_X1 U6086 ( .A1(n9175), .A2(n7337), .ZN(n4401) );
  INV_X1 U6087 ( .A(n9580), .ZN(n4988) );
  INV_X1 U6088 ( .A(n10064), .ZN(n4836) );
  INV_X1 U6089 ( .A(n6038), .ZN(n6037) );
  AND2_X1 U6090 ( .A1(n5568), .A2(n5609), .ZN(n4402) );
  INV_X1 U6091 ( .A(n10243), .ZN(n4834) );
  NAND2_X1 U6092 ( .A1(n7906), .A2(n7905), .ZN(n10214) );
  INV_X1 U6093 ( .A(n6836), .ZN(n6842) );
  AND3_X1 U6094 ( .A1(n4908), .A2(n7563), .A3(n4907), .ZN(n4403) );
  AND2_X1 U6095 ( .A1(n4908), .A2(n7563), .ZN(n4404) );
  OAI211_X1 U6096 ( .C1(n6516), .C2(n8175), .A(n6518), .B(n6517), .ZN(n7399)
         );
  INV_X1 U6097 ( .A(n5143), .ZN(n5126) );
  AND2_X1 U6098 ( .A1(n4489), .A2(n5271), .ZN(n4405) );
  OR2_X1 U6099 ( .A1(n6745), .A2(n6934), .ZN(n4406) );
  NAND2_X1 U6100 ( .A1(n5416), .A2(n5415), .ZN(n4407) );
  AND2_X1 U6101 ( .A1(n10027), .A2(n4864), .ZN(n4408) );
  NOR2_X1 U6102 ( .A1(n8286), .A2(n9951), .ZN(n4409) );
  AND2_X1 U6103 ( .A1(n10409), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4410) );
  AND3_X1 U6104 ( .A1(n5178), .A2(n5177), .A3(n5179), .ZN(n4411) );
  AND2_X1 U6105 ( .A1(n9161), .A2(n9383), .ZN(n4412) );
  AND2_X1 U6106 ( .A1(n5002), .A2(n5003), .ZN(n4413) );
  OR2_X1 U6107 ( .A1(n10214), .A2(n9842), .ZN(n4414) );
  INV_X1 U6108 ( .A(n7377), .ZN(n7290) );
  NAND2_X1 U6109 ( .A1(n7044), .A2(n7043), .ZN(n7377) );
  NAND2_X1 U6110 ( .A1(n8458), .A2(n8457), .ZN(n8504) );
  INV_X1 U6111 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5695) );
  INV_X1 U6112 ( .A(n5743), .ZN(n5026) );
  NAND2_X1 U6113 ( .A1(n5617), .A2(n5616), .ZN(n9326) );
  INV_X1 U6114 ( .A(n9404), .ZN(n5924) );
  NAND2_X1 U6115 ( .A1(n6626), .A2(n6625), .ZN(n7174) );
  INV_X1 U6116 ( .A(n8477), .ZN(n4893) );
  NAND2_X1 U6117 ( .A1(n5438), .A2(n5437), .ZN(n9489) );
  INV_X1 U6118 ( .A(n5903), .ZN(n4727) );
  NOR2_X1 U6119 ( .A1(n6544), .A2(n4795), .ZN(n4416) );
  AND3_X1 U6120 ( .A1(n5058), .A2(n5057), .A3(n5056), .ZN(n4417) );
  NAND2_X1 U6121 ( .A1(n10249), .A2(n10047), .ZN(n4418) );
  NOR2_X1 U6122 ( .A1(n5505), .A2(n9421), .ZN(n4419) );
  AND2_X1 U6123 ( .A1(n8038), .A2(n8037), .ZN(n10064) );
  INV_X1 U6124 ( .A(n4868), .ZN(n10204) );
  NAND2_X1 U6125 ( .A1(n5522), .A2(n5521), .ZN(n9580) );
  AND2_X1 U6126 ( .A1(n4943), .A2(n7645), .ZN(n4420) );
  AND2_X1 U6127 ( .A1(n4922), .A2(n9727), .ZN(n4421) );
  AND2_X1 U6128 ( .A1(n5826), .A2(n4728), .ZN(n4422) );
  AND2_X1 U6129 ( .A1(n9319), .A2(n5816), .ZN(n4423) );
  NAND2_X1 U6130 ( .A1(n4925), .A2(n4932), .ZN(n9710) );
  INV_X1 U6131 ( .A(n5802), .ZN(n9390) );
  INV_X1 U6132 ( .A(n7435), .ZN(n5248) );
  AND2_X1 U6133 ( .A1(n5824), .A2(n5826), .ZN(n4424) );
  AOI21_X1 U6134 ( .B1(n4504), .B2(n4863), .A(n4865), .ZN(n4862) );
  AND2_X1 U6135 ( .A1(n5744), .A2(n5743), .ZN(n7716) );
  NAND2_X1 U6136 ( .A1(n9068), .A2(n8842), .ZN(n4425) );
  AND2_X1 U6137 ( .A1(n8174), .A2(n4581), .ZN(n4426) );
  OR2_X1 U6138 ( .A1(n10237), .A2(n10048), .ZN(n4427) );
  NAND2_X1 U6139 ( .A1(n8008), .A2(n8007), .ZN(n4428) );
  AND2_X1 U6140 ( .A1(n4761), .A2(n5533), .ZN(n4429) );
  NAND2_X1 U6141 ( .A1(n9335), .A2(n9334), .ZN(n4566) );
  INV_X1 U6142 ( .A(n4413), .ZN(n5000) );
  AND2_X1 U6143 ( .A1(n5663), .A2(n5662), .ZN(n9638) );
  INV_X1 U6144 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5059) );
  AND2_X1 U6145 ( .A1(n4892), .A2(n4890), .ZN(n4430) );
  AND3_X1 U6146 ( .A1(n5900), .A2(n5755), .A3(n5754), .ZN(n4431) );
  OR2_X1 U6147 ( .A1(n5026), .A2(n5742), .ZN(n4432) );
  NOR2_X1 U6148 ( .A1(n4918), .A2(n8943), .ZN(n4433) );
  NOR2_X1 U6149 ( .A1(n7581), .A2(n7580), .ZN(n4434) );
  OR2_X1 U6150 ( .A1(n9548), .A2(n8881), .ZN(n5818) );
  INV_X1 U6151 ( .A(n4856), .ZN(n4855) );
  NAND2_X1 U6152 ( .A1(n8532), .A2(n4414), .ZN(n4856) );
  INV_X1 U6153 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6902) );
  NAND2_X1 U6154 ( .A1(n7042), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4435) );
  OR2_X1 U6155 ( .A1(n8838), .A2(n9071), .ZN(n4436) );
  INV_X1 U6156 ( .A(n8205), .ZN(n8320) );
  OR2_X1 U6157 ( .A1(n10301), .A2(n7362), .ZN(n8205) );
  OR2_X1 U6158 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n4437) );
  OR2_X1 U6159 ( .A1(n6082), .A2(n6081), .ZN(n4438) );
  NAND2_X1 U6160 ( .A1(n7644), .A2(n7643), .ZN(n4439) );
  OR2_X1 U6161 ( .A1(n9373), .A2(n5804), .ZN(n4440) );
  INV_X1 U6162 ( .A(n5004), .ZN(n4998) );
  NAND2_X1 U6163 ( .A1(n9030), .A2(n9128), .ZN(n5004) );
  NAND2_X1 U6164 ( .A1(n9047), .A2(n9499), .ZN(n4441) );
  AND2_X1 U6165 ( .A1(n6697), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4442) );
  NOR2_X1 U6166 ( .A1(n10036), .A2(n10014), .ZN(n4443) );
  NAND2_X1 U6167 ( .A1(n5982), .A2(n5694), .ZN(n4444) );
  AND2_X1 U6168 ( .A1(n4834), .A2(n10064), .ZN(n4445) );
  AND2_X1 U6169 ( .A1(n5818), .A2(n5826), .ZN(n7840) );
  INV_X1 U6170 ( .A(n7840), .ZN(n4996) );
  OR2_X1 U6171 ( .A1(n4694), .A2(n8388), .ZN(n4446) );
  NAND2_X1 U6172 ( .A1(n5258), .A2(n5257), .ZN(n9629) );
  AND2_X1 U6173 ( .A1(n8508), .A2(n8498), .ZN(n4447) );
  AND2_X1 U6174 ( .A1(n8376), .A2(n8375), .ZN(n8422) );
  NAND2_X1 U6175 ( .A1(n5514), .A2(n5513), .ZN(n4448) );
  AND2_X1 U6176 ( .A1(n4583), .A2(n8162), .ZN(n4449) );
  NAND2_X1 U6177 ( .A1(n9352), .A2(n5808), .ZN(n9373) );
  INV_X1 U6178 ( .A(n9373), .ZN(n4659) );
  INV_X1 U6179 ( .A(n4983), .ZN(n4982) );
  NAND2_X1 U6180 ( .A1(n4985), .A2(n5802), .ZN(n4983) );
  OR2_X1 U6181 ( .A1(n5001), .A2(n10507), .ZN(n4450) );
  AND2_X1 U6182 ( .A1(n5304), .A2(n5303), .ZN(n4451) );
  AND2_X1 U6183 ( .A1(n8499), .A2(n8535), .ZN(n4452) );
  OR2_X1 U6184 ( .A1(n7772), .A2(n9146), .ZN(n5767) );
  INV_X1 U6185 ( .A(n5767), .ZN(n5023) );
  OR2_X1 U6186 ( .A1(n9175), .A2(n7337), .ZN(n4453) );
  INV_X1 U6187 ( .A(n8401), .ZN(n4709) );
  AND2_X1 U6188 ( .A1(n4766), .A2(n4762), .ZN(n4454) );
  INV_X1 U6189 ( .A(n10207), .ZN(n4918) );
  AND2_X1 U6190 ( .A1(n9496), .A2(n5910), .ZN(n4455) );
  NAND2_X1 U6191 ( .A1(n9154), .A2(n9166), .ZN(n4456) );
  NOR2_X1 U6192 ( .A1(n9900), .A2(n9899), .ZN(n4457) );
  INV_X1 U6193 ( .A(n9353), .ZN(n5926) );
  AND2_X1 U6194 ( .A1(n5811), .A2(n5812), .ZN(n9353) );
  AND2_X1 U6195 ( .A1(n8472), .A2(n10122), .ZN(n4458) );
  XNOR2_X1 U6196 ( .A(n5377), .B(SI_14_), .ZN(n5376) );
  AND2_X1 U6197 ( .A1(n9030), .A2(n4960), .ZN(n4459) );
  NOR2_X1 U6198 ( .A1(n10174), .A2(n4905), .ZN(n4460) );
  NOR2_X1 U6199 ( .A1(n10409), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n4461) );
  OR2_X1 U6200 ( .A1(n7377), .A2(n7305), .ZN(n8227) );
  AND2_X1 U6201 ( .A1(n8047), .A2(n4924), .ZN(n4462) );
  OR2_X1 U6202 ( .A1(n9638), .A2(n5020), .ZN(n4463) );
  AND2_X1 U6203 ( .A1(n4390), .A2(n8344), .ZN(n4464) );
  BUF_X1 U6204 ( .A(n6622), .Z(n7851) );
  AND2_X1 U6205 ( .A1(n4398), .A2(n4744), .ZN(n4465) );
  INV_X1 U6206 ( .A(n8869), .ZN(n9159) );
  AND2_X1 U6207 ( .A1(n5603), .A2(n5602), .ZN(n8869) );
  AND2_X1 U6208 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_8__SCAN_IN), 
        .ZN(n4466) );
  INV_X1 U6209 ( .A(n7507), .ZN(n7569) );
  AND2_X1 U6210 ( .A1(n5842), .A2(n5834), .ZN(n5838) );
  INV_X1 U6211 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4966) );
  INV_X1 U6212 ( .A(n10192), .ZN(n4524) );
  INV_X1 U6213 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n4642) );
  AND2_X1 U6214 ( .A1(n7047), .A2(n4909), .ZN(n4467) );
  AND2_X1 U6215 ( .A1(n5642), .A2(n5641), .ZN(n8881) );
  OR2_X1 U6216 ( .A1(n7489), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n4468) );
  NAND2_X1 U6217 ( .A1(n7006), .A2(n7005), .ZN(n7061) );
  INV_X1 U6218 ( .A(n4494), .ZN(n7635) );
  NAND2_X1 U6219 ( .A1(n7888), .A2(n7887), .ZN(n10232) );
  INV_X1 U6220 ( .A(n10232), .ZN(n10023) );
  AND2_X1 U6221 ( .A1(n5532), .A2(n5531), .ZN(n9005) );
  NAND2_X1 U6222 ( .A1(n7474), .A2(n4957), .ZN(n4959) );
  INV_X1 U6223 ( .A(n4912), .ZN(n10065) );
  NOR2_X1 U6224 ( .A1(n10081), .A2(n10249), .ZN(n4912) );
  AND2_X1 U6225 ( .A1(n7188), .A2(n7179), .ZN(n4469) );
  NOR2_X1 U6226 ( .A1(n9642), .A2(n9615), .ZN(n4470) );
  OR2_X1 U6227 ( .A1(n5658), .A2(SI_29_), .ZN(n4471) );
  INV_X1 U6228 ( .A(n4913), .ZN(n10154) );
  NOR2_X1 U6229 ( .A1(n7635), .A2(n4915), .ZN(n4913) );
  INV_X1 U6230 ( .A(n9345), .ZN(n9646) );
  NAND2_X1 U6231 ( .A1(n5594), .A2(n5593), .ZN(n9345) );
  INV_X1 U6232 ( .A(n9308), .ZN(n5972) );
  NAND2_X1 U6233 ( .A1(n5650), .A2(n5649), .ZN(n9308) );
  NAND2_X1 U6234 ( .A1(n4902), .A2(n4900), .ZN(n4906) );
  OR2_X1 U6235 ( .A1(n9670), .A2(n9646), .ZN(n4472) );
  AND2_X1 U6236 ( .A1(n5773), .A2(n4441), .ZN(n7831) );
  NOR2_X1 U6237 ( .A1(n9913), .A2(n4782), .ZN(n4473) );
  AND2_X1 U6238 ( .A1(n4652), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n4474) );
  AND2_X1 U6239 ( .A1(n4655), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n4475) );
  AND2_X1 U6240 ( .A1(n4791), .A2(n4790), .ZN(n4476) );
  AND2_X1 U6241 ( .A1(n6349), .A2(n10439), .ZN(n9838) );
  INV_X1 U6242 ( .A(n9838), .ZN(n4582) );
  NAND2_X1 U6243 ( .A1(n5480), .A2(n5479), .ZN(n9433) );
  INV_X1 U6244 ( .A(n9433), .ZN(n4951) );
  INV_X1 U6245 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n4653) );
  INV_X1 U6246 ( .A(n8259), .ZN(n6588) );
  XNOR2_X1 U6247 ( .A(n5671), .B(n5670), .ZN(n6878) );
  INV_X1 U6248 ( .A(n6878), .ZN(n5879) );
  INV_X1 U6249 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n4656) );
  INV_X1 U6250 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n4654) );
  AND2_X1 U6251 ( .A1(n8227), .A2(n8306), .ZN(n8305) );
  INV_X1 U6252 ( .A(n8305), .ZN(n8258) );
  AND2_X1 U6253 ( .A1(n6473), .A2(n4636), .ZN(n4477) );
  INV_X1 U6254 ( .A(n9623), .ZN(n4949) );
  NAND2_X1 U6255 ( .A1(n7525), .A2(n5716), .ZN(n6815) );
  INV_X1 U6256 ( .A(n6815), .ZN(n4604) );
  INV_X1 U6257 ( .A(n4547), .ZN(n7088) );
  AND2_X1 U6258 ( .A1(n4573), .A2(n6554), .ZN(n4478) );
  OR2_X1 U6259 ( .A1(n8911), .A2(n8910), .ZN(n4479) );
  AND2_X1 U6260 ( .A1(n7851), .A2(n4770), .ZN(n4480) );
  AND2_X1 U6261 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n4481) );
  NAND3_X1 U6262 ( .A1(n4908), .A2(n7563), .A3(n10455), .ZN(n4482) );
  AND2_X1 U6263 ( .A1(n6385), .A2(n6382), .ZN(n9815) );
  INV_X1 U6264 ( .A(n8913), .ZN(n4751) );
  INV_X1 U6265 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5867) );
  XNOR2_X1 U6266 ( .A(n5698), .B(P2_IR_REG_20__SCAN_IN), .ZN(n5931) );
  AND2_X1 U6267 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n4483) );
  INV_X1 U6268 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4598) );
  INV_X1 U6269 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10527) );
  INV_X1 U6270 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n4509) );
  INV_X1 U6271 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n4523) );
  AOI21_X1 U6272 ( .B1(n9340), .B2(n9524), .A(n9339), .ZN(n9559) );
  CLKBUF_X1 U6273 ( .A(n10163), .Z(n4484) );
  INV_X2 U6274 ( .A(n10340), .ZN(n10350) );
  NAND2_X1 U6275 ( .A1(n9563), .A2(n4485), .ZN(P2_U3546) );
  NAND2_X1 U6276 ( .A1(n9645), .A2(n4472), .ZN(P2_U3514) );
  NAND2_X2 U6277 ( .A1(n5909), .A2(n7822), .ZN(n7828) );
  AOI21_X2 U6278 ( .B1(n9431), .B2(n9439), .A(n5922), .ZN(n9411) );
  OR2_X1 U6279 ( .A1(n9530), .A2(n7018), .ZN(n9520) );
  NAND2_X1 U6280 ( .A1(n7795), .A2(n5908), .ZN(n7830) );
  OAI21_X1 U6281 ( .B1(n9333), .B2(n5927), .A(n5003), .ZN(n9316) );
  NAND2_X1 U6282 ( .A1(n7739), .A2(n5904), .ZN(n4488) );
  NAND2_X1 U6283 ( .A1(n5724), .A2(n6814), .ZN(n6836) );
  NAND2_X1 U6284 ( .A1(n5474), .A2(n4454), .ZN(n4490) );
  NAND3_X1 U6285 ( .A1(n4535), .A2(n8431), .A3(n4415), .ZN(n4491) );
  AOI21_X1 U6286 ( .B1(n4405), .B2(n5270), .A(n4492), .ZN(n5305) );
  NAND3_X1 U6287 ( .A1(n6005), .A2(n8773), .A3(n6004), .ZN(n6028) );
  NAND2_X1 U6288 ( .A1(n10032), .A2(n10023), .ZN(n10019) );
  AOI211_X1 U6289 ( .C1(n10214), .C2(n9972), .A(n10456), .B(n9971), .ZN(n10213) );
  NAND2_X2 U6290 ( .A1(n6249), .A2(n6248), .ZN(n6622) );
  NOR2_X4 U6291 ( .A1(n7001), .A2(n6999), .ZN(n7047) );
  AND2_X2 U6292 ( .A1(n4494), .A2(n4493), .ZN(n10109) );
  NAND2_X2 U6293 ( .A1(n7283), .A2(n7223), .ZN(n7352) );
  NAND2_X1 U6294 ( .A1(n8958), .A2(n4514), .ZN(n8956) );
  INV_X1 U6295 ( .A(n8099), .ZN(n9698) );
  NAND2_X1 U6296 ( .A1(n6823), .A2(n6827), .ZN(n6822) );
  NAND2_X1 U6297 ( .A1(n7797), .A2(n7796), .ZN(n7795) );
  NAND2_X2 U6298 ( .A1(n9372), .A2(n5925), .ZN(n9350) );
  INV_X2 U6299 ( .A(n5941), .ZN(n10488) );
  AOI21_X1 U6300 ( .B1(n9556), .B2(n10510), .A(n4495), .ZN(n9640) );
  INV_X1 U6301 ( .A(n5873), .ZN(n4965) );
  NAND2_X1 U6302 ( .A1(n6809), .A2(n4970), .ZN(n4969) );
  XNOR2_X1 U6303 ( .A(n4498), .B(n8815), .ZN(P1_U3263) );
  NAND3_X1 U6304 ( .A1(n5042), .A2(n8545), .A3(n8544), .ZN(n4498) );
  NAND2_X1 U6305 ( .A1(n9965), .A2(n9964), .ZN(n9963) );
  NAND2_X1 U6306 ( .A1(n10000), .A2(n9999), .ZN(n9998) );
  AOI21_X1 U6307 ( .B1(n8538), .B2(n10117), .A(n8537), .ZN(n10210) );
  INV_X1 U6308 ( .A(n6455), .ZN(n4500) );
  AOI21_X2 U6309 ( .B1(n7459), .B2(n8313), .A(n7248), .ZN(n7510) );
  NAND2_X2 U6310 ( .A1(n6434), .A2(n6433), .ZN(n9855) );
  AOI21_X2 U6311 ( .B1(n8504), .B2(n8503), .A(n5038), .ZN(n9979) );
  AND2_X4 U6312 ( .A1(n6364), .A2(n6365), .ZN(n8184) );
  OAI21_X2 U6313 ( .B1(n7050), .B2(P1_REG3_REG_3__SCAN_IN), .A(n6431), .ZN(
        n6432) );
  AOI21_X2 U6314 ( .B1(n7510), .B2(n7509), .A(n7508), .ZN(n7616) );
  NAND3_X1 U6315 ( .A1(n7397), .A2(n8262), .A3(n7401), .ZN(n6744) );
  NAND2_X1 U6316 ( .A1(n6669), .A2(n6668), .ZN(n7397) );
  NAND4_X1 U6317 ( .A1(n6389), .A2(n6390), .A3(n6387), .A4(n6388), .ZN(n6446)
         );
  NAND2_X1 U6318 ( .A1(n10024), .A2(n4544), .ZN(n9997) );
  OAI21_X1 U6319 ( .B1(n10108), .B2(n4839), .A(n4838), .ZN(n4837) );
  NAND2_X1 U6320 ( .A1(n4670), .A2(n4668), .ZN(n5434) );
  INV_X1 U6321 ( .A(n4890), .ZN(n4888) );
  INV_X1 U6322 ( .A(n4505), .ZN(n6934) );
  INV_X1 U6323 ( .A(n6419), .ZN(n6420) );
  NOR2_X1 U6324 ( .A1(n5212), .A2(n5211), .ZN(n5232) );
  OAI21_X2 U6325 ( .B1(n8533), .B2(n8532), .A(n8531), .ZN(n10211) );
  NAND2_X1 U6326 ( .A1(n5162), .A2(n5161), .ZN(n5231) );
  NAND2_X1 U6327 ( .A1(n4375), .A2(n4406), .ZN(n7034) );
  NAND2_X1 U6328 ( .A1(n4857), .A2(n4855), .ZN(n8531) );
  NAND2_X1 U6329 ( .A1(n9979), .A2(n8506), .ZN(n4858) );
  NAND2_X1 U6330 ( .A1(n8454), .A2(n8453), .ZN(n10059) );
  NAND2_X1 U6331 ( .A1(n5921), .A2(n5920), .ZN(n9431) );
  OAI21_X1 U6332 ( .B1(n9640), .B2(n10512), .A(n4506), .ZN(P2_U3515) );
  INV_X2 U6333 ( .A(n6045), .ZN(n6829) );
  INV_X1 U6334 ( .A(n7716), .ZN(n4513) );
  OAI21_X1 U6335 ( .B1(n5193), .B2(n4509), .A(n4508), .ZN(n5214) );
  INV_X1 U6336 ( .A(n7692), .ZN(n4950) );
  NAND2_X1 U6337 ( .A1(n9270), .A2(n9269), .ZN(n9268) );
  NAND2_X1 U6338 ( .A1(n4542), .A2(n4540), .ZN(P2_U3264) );
  NAND2_X1 U6339 ( .A1(n9551), .A2(n4450), .ZN(n4650) );
  NOR2_X2 U6340 ( .A1(n7604), .A2(n7605), .ZN(n7608) );
  NOR2_X4 U6341 ( .A1(n9508), .A2(n9512), .ZN(n9507) );
  NAND2_X1 U6342 ( .A1(n5888), .A2(n4976), .ZN(n4975) );
  INV_X1 U6343 ( .A(n4968), .ZN(n4967) );
  NAND2_X1 U6344 ( .A1(n4974), .A2(n4453), .ZN(n4971) );
  NAND2_X1 U6345 ( .A1(n4511), .A2(n8443), .ZN(P1_U3240) );
  NAND2_X1 U6346 ( .A1(n6635), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6903) );
  AND2_X2 U6347 ( .A1(n4600), .A2(n5053), .ZN(n5060) );
  NAND2_X2 U6348 ( .A1(n5079), .A2(n4964), .ZN(n7757) );
  NAND3_X1 U6349 ( .A1(n5248), .A2(n4513), .A3(n5893), .ZN(n5892) );
  NAND2_X1 U6350 ( .A1(n5998), .A2(n8570), .ZN(n6000) );
  NAND2_X1 U6351 ( .A1(n5357), .A2(n5356), .ZN(n5380) );
  INV_X1 U6352 ( .A(n4552), .ZN(n4551) );
  NAND3_X1 U6353 ( .A1(n5992), .A2(n5991), .A3(n6009), .ZN(n6033) );
  NAND2_X1 U6354 ( .A1(n6454), .A2(n6447), .ZN(n6592) );
  NAND2_X1 U6355 ( .A1(n4842), .A2(n4840), .ZN(n10108) );
  INV_X1 U6356 ( .A(n4837), .ZN(n10105) );
  NOR2_X2 U6357 ( .A1(n10417), .A2(n4520), .ZN(n6726) );
  NAND2_X1 U6358 ( .A1(n9887), .A2(n9886), .ZN(n9895) );
  OAI21_X1 U6359 ( .B1(n7250), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7116), .ZN(
        n7117) );
  NAND2_X1 U6360 ( .A1(n6324), .A2(n6323), .ZN(n6481) );
  NOR2_X1 U6361 ( .A1(n9934), .A2(n9933), .ZN(n9937) );
  OAI21_X1 U6362 ( .B1(n9952), .B2(n9951), .A(n4624), .ZN(P1_U3260) );
  NAND2_X1 U6363 ( .A1(n10121), .A2(n4458), .ZN(n4842) );
  NAND2_X1 U6364 ( .A1(n4525), .A2(n4524), .ZN(n8545) );
  INV_X1 U6365 ( .A(n10211), .ZN(n4525) );
  AOI21_X2 U6366 ( .B1(n9989), .B2(n8496), .A(n8495), .ZN(n9965) );
  NAND2_X1 U6367 ( .A1(n4979), .A2(n4977), .ZN(n9374) );
  NAND2_X1 U6368 ( .A1(n9333), .A2(n4413), .ZN(n4997) );
  INV_X1 U6369 ( .A(n4900), .ZN(n4898) );
  NAND3_X1 U6370 ( .A1(n9968), .A2(n9967), .A3(n4530), .ZN(n10212) );
  NAND2_X1 U6371 ( .A1(n5250), .A2(n5268), .ZN(n5306) );
  NAND2_X1 U6372 ( .A1(n4705), .A2(n4704), .ZN(n4703) );
  NOR2_X1 U6373 ( .A1(n8387), .A2(n4684), .ZN(n8384) );
  NAND2_X1 U6374 ( .A1(n4700), .A2(n8326), .ZN(n4699) );
  NAND2_X1 U6375 ( .A1(n4699), .A2(n8461), .ZN(n8327) );
  NAND3_X1 U6376 ( .A1(n8361), .A2(n8359), .A3(n8360), .ZN(n4539) );
  NAND2_X1 U6377 ( .A1(n9228), .A2(n9227), .ZN(n4748) );
  NAND2_X1 U6378 ( .A1(n9253), .A2(n9254), .ZN(n9252) );
  NAND3_X1 U6379 ( .A1(n5402), .A2(n5060), .A3(n4966), .ZN(n4964) );
  NAND2_X1 U6380 ( .A1(n4827), .A2(n4826), .ZN(n10026) );
  NAND2_X1 U6381 ( .A1(n4725), .A2(n4592), .ZN(n4724) );
  INV_X1 U6382 ( .A(n5726), .ZN(n5717) );
  NAND2_X1 U6383 ( .A1(n4745), .A2(n4546), .ZN(n5726) );
  OR2_X1 U6384 ( .A1(n5828), .A2(n5725), .ZN(n4546) );
  NAND2_X1 U6385 ( .A1(n4737), .A2(n4736), .ZN(n5809) );
  OAI21_X1 U6386 ( .B1(n4589), .B2(n5844), .A(n5843), .ZN(n5861) );
  OAI21_X1 U6387 ( .B1(n4587), .B2(n4730), .A(n4729), .ZN(n4586) );
  NAND2_X1 U6388 ( .A1(n4588), .A2(n4735), .ZN(n4734) );
  NAND2_X1 U6389 ( .A1(n4733), .A2(n4732), .ZN(P2_U3244) );
  NAND2_X1 U6390 ( .A1(n5730), .A2(n5729), .ZN(n4594) );
  NAND2_X1 U6391 ( .A1(n4594), .A2(n5734), .ZN(n4593) );
  NAND2_X1 U6392 ( .A1(n4547), .A2(n10496), .ZN(n5848) );
  NAND2_X2 U6393 ( .A1(n5180), .A2(n4411), .ZN(n4547) );
  NAND2_X1 U6394 ( .A1(n4547), .A2(n8835), .ZN(n6068) );
  NAND2_X1 U6395 ( .A1(n4606), .A2(n4547), .ZN(n5888) );
  AOI22_X1 U6396 ( .A1(n9464), .A2(n9174), .B1(n9462), .B2(n4547), .ZN(n7333)
         );
  AOI22_X1 U6397 ( .A1(n9464), .A2(n4547), .B1(n9177), .B2(n9462), .ZN(n6818)
         );
  NOR2_X1 U6398 ( .A1(n9178), .A2(n7088), .ZN(n4549) );
  OAI21_X2 U6399 ( .B1(n5021), .B2(n4553), .A(n4551), .ZN(n9497) );
  NAND2_X1 U6400 ( .A1(n5223), .A2(n4555), .ZN(n7438) );
  NAND2_X1 U6401 ( .A1(n5508), .A2(n4389), .ZN(n9388) );
  NAND2_X2 U6402 ( .A1(n5066), .A2(n9678), .ZN(n9683) );
  NOR2_X1 U6403 ( .A1(n9859), .A2(n6373), .ZN(n6454) );
  NAND2_X1 U6404 ( .A1(n6549), .A2(n4574), .ZN(n4573) );
  INV_X1 U6405 ( .A(n6515), .ZN(n4572) );
  NAND3_X1 U6406 ( .A1(n4572), .A2(n6549), .A3(n4575), .ZN(n4571) );
  OAI21_X1 U6407 ( .B1(n6515), .B2(n6514), .A(n6513), .ZN(n6550) );
  INV_X1 U6408 ( .A(n6513), .ZN(n4574) );
  INV_X1 U6409 ( .A(n6514), .ZN(n4575) );
  NAND4_X1 U6410 ( .A1(n4593), .A2(n5763), .A3(n4381), .A4(n4400), .ZN(n4592)
         );
  NAND3_X1 U6411 ( .A1(n4739), .A2(n4595), .A3(n4738), .ZN(n4737) );
  NAND2_X1 U6412 ( .A1(n4596), .A2(n5828), .ZN(n4595) );
  NAND2_X1 U6413 ( .A1(n4597), .A2(n5801), .ZN(n4596) );
  NAND3_X1 U6414 ( .A1(n5799), .A2(n5800), .A3(n9389), .ZN(n4597) );
  NAND3_X1 U6415 ( .A1(n4605), .A2(n6842), .A3(n4604), .ZN(n4603) );
  NAND4_X1 U6416 ( .A1(n7831), .A2(n4615), .A3(n4610), .A4(n9471), .ZN(n4609)
         );
  NAND3_X1 U6417 ( .A1(n5838), .A2(n4619), .A3(n4618), .ZN(n4617) );
  NAND3_X1 U6418 ( .A1(n7840), .A2(n4621), .A3(n9353), .ZN(n4620) );
  AOI21_X1 U6419 ( .B1(n4385), .B2(n6473), .A(n4461), .ZN(n4632) );
  OAI21_X1 U6420 ( .B1(n6296), .B2(n8682), .A(n4641), .ZN(n6267) );
  NAND2_X1 U6421 ( .A1(n6296), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6283) );
  XNOR2_X1 U6422 ( .A(n6296), .B(n4642), .ZN(n6295) );
  MUX2_X1 U6423 ( .A(n8682), .B(P1_REG1_REG_1__SCAN_IN), .S(n6296), .Z(n6270)
         );
  NAND3_X1 U6424 ( .A1(n6400), .A2(n6401), .A3(n4643), .ZN(n6445) );
  NAND2_X1 U6425 ( .A1(n7872), .A2(n6296), .ZN(n4643) );
  AOI21_X1 U6426 ( .B1(n6296), .B2(P1_STATE_REG_SCAN_IN), .A(n4645), .ZN(n4644) );
  NOR2_X1 U6427 ( .A1(n10347), .A2(n6399), .ZN(n4645) );
  INV_X1 U6428 ( .A(n6296), .ZN(n4648) );
  NAND2_X1 U6429 ( .A1(n4651), .A2(n4466), .ZN(n5260) );
  NAND2_X1 U6430 ( .A1(n5439), .A2(n4474), .ZN(n5496) );
  NAND2_X1 U6431 ( .A1(n5366), .A2(n4475), .ZN(n5424) );
  NAND2_X4 U6432 ( .A1(n4663), .A2(n4662), .ZN(n5193) );
  NAND2_X1 U6433 ( .A1(n4769), .A2(n4671), .ZN(n4670) );
  OR2_X1 U6434 ( .A1(n8867), .A2(n9025), .ZN(n4677) );
  OAI21_X2 U6435 ( .B1(n9126), .B2(n4681), .A(n4679), .ZN(n8891) );
  NAND3_X1 U6436 ( .A1(n4687), .A2(n8535), .A3(n8369), .ZN(n4686) );
  NAND3_X1 U6437 ( .A1(n8368), .A2(n9964), .A3(n8367), .ZN(n4687) );
  XNOR2_X1 U6438 ( .A(n4688), .B(n5135), .ZN(n5137) );
  NAND2_X1 U6439 ( .A1(n6398), .A2(n4690), .ZN(n4689) );
  INV_X1 U6440 ( .A(n8303), .ZN(n4694) );
  OAI211_X1 U6441 ( .C1(n6933), .C2(n4446), .A(n4693), .B(n4691), .ZN(n8316)
         );
  NAND2_X1 U6442 ( .A1(n8304), .A2(n8303), .ZN(n4693) );
  OR2_X1 U6443 ( .A1(n8323), .A2(n4703), .ZN(n8329) );
  NAND3_X1 U6444 ( .A1(n8408), .A2(n8261), .A3(n8401), .ZN(n4706) );
  NAND4_X1 U6445 ( .A1(n8350), .A2(n8351), .A3(n4719), .A4(n4714), .ZN(n4711)
         );
  INV_X1 U6446 ( .A(n8352), .ZN(n4720) );
  NAND2_X1 U6447 ( .A1(n4721), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5391) );
  NAND2_X1 U6448 ( .A1(n4721), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5265) );
  NAND2_X1 U6449 ( .A1(n4721), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U6450 ( .A1(n4721), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5302) );
  NAND2_X1 U6451 ( .A1(n4721), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U6452 ( .A1(n4721), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5372) );
  NAND2_X1 U6453 ( .A1(n4721), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5427) );
  NAND2_X1 U6454 ( .A1(n4721), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5341) );
  NAND2_X1 U6455 ( .A1(n4721), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5443) );
  NAND2_X1 U6456 ( .A1(n4721), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5466) );
  NAND2_X1 U6457 ( .A1(n4721), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U6458 ( .A1(n4721), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U6459 ( .A1(n4721), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5547) );
  NAND2_X1 U6460 ( .A1(n4721), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U6461 ( .A1(n4721), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U6462 ( .A1(n4721), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U6463 ( .A1(n4721), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U6464 ( .A1(n4721), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5639) );
  NAND2_X1 U6465 ( .A1(n4721), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5652) );
  NAND2_X1 U6466 ( .A1(n4721), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U6467 ( .A1(n4721), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5664) );
  AOI22_X1 U6468 ( .A1(n5672), .A2(P2_REG2_REG_16__SCAN_IN), .B1(
        P2_REG0_REG_16__SCAN_IN), .B2(n4721), .ZN(n5413) );
  OAI21_X1 U6469 ( .B1(n5763), .B2(n4723), .A(n4722), .ZN(n4725) );
  NAND3_X1 U6470 ( .A1(n4431), .A2(n4726), .A3(n5765), .ZN(n4722) );
  NAND3_X1 U6471 ( .A1(n4734), .A2(n5862), .A3(n7095), .ZN(n4733) );
  NAND2_X1 U6472 ( .A1(n4965), .A2(n4465), .ZN(n5065) );
  OAI21_X2 U6473 ( .B1(n9214), .B2(n9213), .A(n9212), .ZN(n9228) );
  INV_X1 U6474 ( .A(n5573), .ZN(n4775) );
  OAI21_X1 U6475 ( .B1(n5644), .B2(n4781), .A(n4779), .ZN(n5678) );
  NAND2_X1 U6476 ( .A1(n4777), .A2(n4776), .ZN(n5681) );
  NAND2_X1 U6477 ( .A1(n5644), .A2(n4779), .ZN(n4777) );
  OAI22_X1 U6478 ( .A1(n7117), .A2(n4789), .B1(n7428), .B2(n4790), .ZN(n9866)
         );
  INV_X1 U6479 ( .A(n4791), .ZN(n7426) );
  AOI21_X1 U6480 ( .B1(n4798), .B2(n4416), .A(n4792), .ZN(n6506) );
  OR4_X2 U6481 ( .A1(n8430), .A2(n9951), .A3(n8429), .A4(n8438), .ZN(n8431) );
  NAND2_X1 U6482 ( .A1(n5677), .A2(n5676), .ZN(n5683) );
  NAND2_X1 U6483 ( .A1(n5624), .A2(n5623), .ZN(n5626) );
  NAND2_X1 U6484 ( .A1(n5434), .A2(n5433), .ZN(n5450) );
  NOR2_X2 U6485 ( .A1(n7180), .A2(n7597), .ZN(n7605) );
  NOR2_X1 U6486 ( .A1(n10388), .A2(n6322), .ZN(n6324) );
  NOR2_X1 U6487 ( .A1(n6506), .A2(n6505), .ZN(n6725) );
  NAND2_X1 U6488 ( .A1(n6727), .A2(n6726), .ZN(n7116) );
  NAND2_X1 U6489 ( .A1(n6301), .A2(n6302), .ZN(n6321) );
  AOI21_X1 U6490 ( .B1(n7138), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6725), .ZN(
        n10419) );
  NOR4_X2 U6491 ( .A1(n8425), .A2(n8282), .A3(n8508), .A4(n8281), .ZN(n8285)
         );
  NAND2_X1 U6492 ( .A1(n4803), .A2(n4802), .ZN(n4801) );
  NAND2_X1 U6493 ( .A1(n7014), .A2(n10481), .ZN(n4803) );
  NAND2_X1 U6494 ( .A1(n6048), .A2(n4801), .ZN(n4800) );
  NAND2_X1 U6495 ( .A1(n8817), .A2(n8818), .ZN(n8816) );
  NAND2_X1 U6496 ( .A1(n9037), .A2(n6150), .ZN(n4804) );
  OR2_X1 U6497 ( .A1(n5406), .A2(n9677), .ZN(n5420) );
  OAI21_X2 U6498 ( .B1(n6071), .B2(n4386), .A(n4808), .ZN(n7276) );
  OAI21_X1 U6499 ( .B1(n6089), .B2(n4813), .A(n4811), .ZN(n6127) );
  NAND2_X1 U6500 ( .A1(n4819), .A2(n4817), .ZN(P2_U3216) );
  NAND2_X1 U6501 ( .A1(n8899), .A2(n4820), .ZN(n4819) );
  NAND2_X1 U6502 ( .A1(n4821), .A2(n8900), .ZN(n4820) );
  NAND2_X1 U6503 ( .A1(n6878), .A2(n8962), .ZN(n6101) );
  XNOR2_X2 U6504 ( .A(n5699), .B(n5695), .ZN(n8962) );
  NAND3_X1 U6505 ( .A1(n4823), .A2(n4825), .A3(n4824), .ZN(n6353) );
  NAND2_X1 U6506 ( .A1(n10059), .A2(n4388), .ZN(n4827) );
  AND2_X1 U6507 ( .A1(n10266), .A2(n10095), .ZN(n4839) );
  NAND2_X1 U6508 ( .A1(n4849), .A2(n4852), .ZN(n8509) );
  NAND2_X1 U6509 ( .A1(n9979), .A2(n4850), .ZN(n4849) );
  NAND2_X1 U6510 ( .A1(n4858), .A2(n4854), .ZN(n4857) );
  AND2_X1 U6511 ( .A1(n4858), .A2(n8505), .ZN(n9962) );
  INV_X1 U6512 ( .A(n4859), .ZN(n10000) );
  NAND2_X1 U6513 ( .A1(n4504), .A2(n8482), .ZN(n10037) );
  NAND2_X1 U6514 ( .A1(n8536), .A2(n4870), .ZN(n4869) );
  NAND2_X1 U6515 ( .A1(n8536), .A2(n8535), .ZN(n8534) );
  NAND2_X1 U6516 ( .A1(n7006), .A2(n4879), .ZN(n4882) );
  NAND2_X1 U6517 ( .A1(n8475), .A2(n4464), .ZN(n4889) );
  NOR2_X1 U6518 ( .A1(n7460), .A2(n4898), .ZN(n4894) );
  NOR2_X1 U6519 ( .A1(n4895), .A2(n4894), .ZN(n8467) );
  AOI21_X1 U6520 ( .B1(n7460), .B2(n8317), .A(n8320), .ZN(n7486) );
  NOR2_X1 U6521 ( .A1(n7485), .A2(n4904), .ZN(n4903) );
  INV_X1 U6522 ( .A(n8317), .ZN(n4904) );
  INV_X1 U6523 ( .A(n4906), .ZN(n8464) );
  NAND3_X1 U6524 ( .A1(n7569), .A2(n4909), .A3(n7047), .ZN(n7504) );
  NAND2_X1 U6525 ( .A1(n9980), .A2(n4393), .ZN(n9970) );
  AND2_X1 U6526 ( .A1(n9980), .A2(n9983), .ZN(n9981) );
  AND2_X2 U6527 ( .A1(n4920), .A2(n6280), .ZN(n4921) );
  NAND2_X1 U6528 ( .A1(n6012), .A2(n4934), .ZN(n4936) );
  NAND2_X1 U6529 ( .A1(n4937), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6347) );
  AOI21_X2 U6530 ( .B1(n7352), .B2(n4420), .A(n4939), .ZN(n7926) );
  AOI21_X1 U6531 ( .B1(n7352), .B2(n7351), .A(n5047), .ZN(n7358) );
  INV_X1 U6532 ( .A(n7357), .ZN(n4945) );
  NAND2_X1 U6533 ( .A1(n4948), .A2(n9689), .ZN(n7952) );
  NAND2_X1 U6534 ( .A1(n9688), .A2(n9691), .ZN(n4948) );
  NAND2_X1 U6535 ( .A1(n9824), .A2(n9822), .ZN(n9828) );
  NAND3_X1 U6536 ( .A1(n4948), .A2(n9689), .A3(n4947), .ZN(n9824) );
  NOR2_X2 U6537 ( .A1(n7690), .A2(n7700), .ZN(n7750) );
  INV_X1 U6538 ( .A(n4959), .ZN(n7722) );
  AND2_X2 U6539 ( .A1(n9412), .A2(n4459), .ZN(n9355) );
  NAND2_X1 U6540 ( .A1(n4964), .A2(n4963), .ZN(n5076) );
  NAND2_X1 U6541 ( .A1(n7828), .A2(n4455), .ZN(n9447) );
  INV_X1 U6542 ( .A(n4971), .ZN(n4970) );
  INV_X1 U6543 ( .A(n6809), .ZN(n4973) );
  OAI21_X1 U6544 ( .B1(n4971), .B2(n5888), .A(n4401), .ZN(n4968) );
  NAND2_X1 U6545 ( .A1(n9411), .A2(n4980), .ZN(n4979) );
  NAND2_X1 U6546 ( .A1(n4989), .A2(n4990), .ZN(n5928) );
  NAND2_X1 U6547 ( .A1(n9350), .A2(n4992), .ZN(n4989) );
  AOI21_X2 U6548 ( .B1(n9350), .B2(n5926), .A(n4998), .ZN(n9333) );
  NAND2_X1 U6549 ( .A1(n9317), .A2(n5819), .ZN(n7839) );
  OAI21_X1 U6550 ( .B1(n9317), .B2(n4996), .A(n5008), .ZN(n5934) );
  INV_X1 U6551 ( .A(n5005), .ZN(n5656) );
  AOI21_X1 U6552 ( .B1(n9317), .B2(n5008), .A(n5006), .ZN(n5005) );
  OR2_X1 U6553 ( .A1(n5675), .A2(n5016), .ZN(n5010) );
  NAND3_X1 U6554 ( .A1(n5010), .A2(n5009), .A3(n5011), .ZN(n5704) );
  NAND2_X1 U6555 ( .A1(n5675), .A2(n5015), .ZN(n5009) );
  NAND2_X1 U6556 ( .A1(n7743), .A2(n5375), .ZN(n5021) );
  NAND2_X1 U6557 ( .A1(n7714), .A2(n5025), .ZN(n7685) );
  INV_X1 U6558 ( .A(n5048), .ZN(n5027) );
  NAND2_X1 U6559 ( .A1(n7526), .A2(n5028), .ZN(n5030) );
  AND2_X1 U6560 ( .A1(n5725), .A2(n7331), .ZN(n5028) );
  NAND2_X1 U6561 ( .A1(n7526), .A2(n5725), .ZN(n5032) );
  NAND3_X1 U6562 ( .A1(n5030), .A2(n5222), .A3(n5029), .ZN(n5223) );
  NAND2_X1 U6563 ( .A1(n5034), .A2(n5033), .ZN(n9335) );
  XNOR2_X1 U6564 ( .A(n5585), .B(n5586), .ZN(n7894) );
  NAND2_X1 U6565 ( .A1(n7903), .A2(n7902), .ZN(n7906) );
  OR2_X1 U6566 ( .A1(n6047), .A2(n6046), .ZN(n6048) );
  NAND2_X1 U6567 ( .A1(n8259), .A2(n8220), .ZN(n6676) );
  NAND2_X1 U6568 ( .A1(n8534), .A2(n5050), .ZN(n8538) );
  NAND2_X1 U6569 ( .A1(n8184), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6389) );
  NAND2_X1 U6570 ( .A1(n5942), .A2(n7415), .ZN(n6811) );
  NOR2_X2 U6571 ( .A1(n6811), .A2(n5104), .ZN(n7530) );
  XNOR2_X1 U6572 ( .A(n5137), .B(n5136), .ZN(n6399) );
  MUX2_X2 U6573 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5078), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5079) );
  NAND2_X1 U6574 ( .A1(n4371), .A2(n4409), .ZN(n6352) );
  AND2_X1 U6575 ( .A1(n6377), .A2(n6376), .ZN(n6381) );
  AND2_X1 U6576 ( .A1(n10204), .A2(n10203), .ZN(n10205) );
  NAND2_X1 U6577 ( .A1(n7723), .A2(n7730), .ZN(n7692) );
  NAND2_X1 U6578 ( .A1(n9335), .A2(n5605), .ZN(n9318) );
  NAND2_X1 U6579 ( .A1(n5883), .A2(n9520), .ZN(n9519) );
  OR2_X1 U6580 ( .A1(n9368), .A2(n5598), .ZN(n5567) );
  INV_X1 U6581 ( .A(n4372), .ZN(n8442) );
  NAND2_X1 U6582 ( .A1(n9355), .A2(n9646), .ZN(n9341) );
  INV_X1 U6583 ( .A(n6445), .ZN(n6459) );
  INV_X1 U6584 ( .A(n6839), .ZN(n5942) );
  AOI211_X1 U6585 ( .C1(n6840), .C2(n6839), .A(n9538), .B(n6838), .ZN(n7413)
         );
  NOR2_X1 U6586 ( .A1(n9028), .A2(n8865), .ZN(n8867) );
  OAI222_X1 U6587 ( .A1(P2_U3152), .A2(n8933), .B1(n9684), .B2(n10344), .C1(
        n8932), .C2(n9686), .ZN(P2_U3328) );
  AND2_X2 U6588 ( .A1(n8933), .A2(n5070), .ZN(n5175) );
  INV_X1 U6589 ( .A(n8933), .ZN(n5069) );
  NAND2_X1 U6590 ( .A1(n8825), .A2(n9537), .ZN(n6839) );
  INV_X2 U6591 ( .A(n10512), .ZN(n10513) );
  NOR2_X1 U6592 ( .A1(n8856), .A2(n8985), .ZN(n5035) );
  NOR2_X1 U6593 ( .A1(n5504), .A2(n9419), .ZN(n5036) );
  NAND2_X1 U6594 ( .A1(n10513), .A2(n9630), .ZN(n9670) );
  OR2_X1 U6595 ( .A1(n5978), .A2(n9615), .ZN(n5037) );
  AND2_X1 U6596 ( .A1(n9747), .A2(n9993), .ZN(n5038) );
  OR2_X1 U6597 ( .A1(n10009), .A2(n10015), .ZN(n5039) );
  NOR2_X1 U6598 ( .A1(n5972), .A2(n9615), .ZN(n5040) );
  OR2_X1 U6599 ( .A1(n5978), .A2(n9670), .ZN(n5041) );
  OR2_X1 U6600 ( .A1(n10210), .A2(n10437), .ZN(n5042) );
  AND3_X1 U6601 ( .A1(n6355), .A2(n6354), .A3(n6359), .ZN(n5043) );
  NAND2_X1 U6602 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n5044) );
  AND2_X1 U6603 ( .A1(n5790), .A2(n5794), .ZN(n5045) );
  NAND2_X1 U6604 ( .A1(n5691), .A2(n5690), .ZN(n5982) );
  AND2_X1 U6605 ( .A1(n5209), .A2(n5208), .ZN(n5046) );
  NOR2_X1 U6606 ( .A1(n7350), .A2(n7349), .ZN(n5047) );
  NAND2_X1 U6607 ( .A1(n6040), .A2(n7785), .ZN(n5048) );
  OR2_X1 U6608 ( .A1(n6883), .A2(n6882), .ZN(n5049) );
  NAND2_X1 U6609 ( .A1(n8254), .A2(n8421), .ZN(n8508) );
  AND3_X1 U6610 ( .A1(n10128), .A2(n8470), .A3(n10124), .ZN(n5051) );
  NOR2_X1 U6611 ( .A1(n9728), .A2(n9779), .ZN(n5052) );
  AND2_X1 U6612 ( .A1(n5800), .A2(n9420), .ZN(n5791) );
  INV_X1 U6613 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6004) );
  INV_X1 U6614 ( .A(n6826), .ZN(n5158) );
  INV_X1 U6615 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6003) );
  OR2_X1 U6616 ( .A1(n5926), .A2(n9352), .ZN(n9334) );
  NAND2_X1 U6617 ( .A1(n5980), .A2(n9155), .ZN(n5937) );
  NAND2_X1 U6618 ( .A1(n6045), .A2(n10488), .ZN(n5846) );
  AND2_X1 U6619 ( .A1(n9727), .A2(n8068), .ZN(n8069) );
  INV_X1 U6620 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n8764) );
  INV_X1 U6621 ( .A(n8508), .ZN(n8499) );
  INV_X1 U6622 ( .A(n7034), .ZN(n6997) );
  INV_X1 U6623 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6359) );
  INV_X1 U6624 ( .A(n5586), .ZN(n5587) );
  AND2_X1 U6625 ( .A1(n5489), .A2(n5488), .ZN(n5490) );
  INV_X1 U6626 ( .A(n5472), .ZN(n5473) );
  INV_X1 U6627 ( .A(n5395), .ZN(n5396) );
  INV_X1 U6628 ( .A(n9301), .ZN(n5944) );
  AND2_X1 U6629 ( .A1(n9781), .A2(n9780), .ZN(n9725) );
  INV_X1 U6630 ( .A(n7174), .ZN(n6745) );
  INV_X1 U6631 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6636) );
  INV_X1 U6632 ( .A(n8184), .ZN(n7050) );
  INV_X1 U6633 ( .A(n9888), .ZN(n9889) );
  INV_X1 U6634 ( .A(n10128), .ZN(n8472) );
  XNOR2_X1 U6635 ( .A(n6035), .B(n6355), .ZN(n6248) );
  INV_X1 U6636 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6009) );
  INV_X1 U6637 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6491) );
  INV_X1 U6638 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U6639 ( .A1(n5193), .A2(n8176), .ZN(n5097) );
  OR2_X1 U6640 ( .A1(n9343), .A2(n5598), .ZN(n5603) );
  OR2_X1 U6641 ( .A1(n4370), .A2(n5067), .ZN(n5074) );
  NAND2_X1 U6642 ( .A1(n5061), .A2(n9677), .ZN(n5075) );
  OR2_X1 U6643 ( .A1(n7602), .A2(n7603), .ZN(n8904) );
  OR2_X1 U6644 ( .A1(n9278), .A2(n9279), .ZN(n9276) );
  INV_X1 U6645 ( .A(n5457), .ZN(n5435) );
  AND2_X1 U6646 ( .A1(n8116), .A2(n8115), .ZN(n9740) );
  OR2_X1 U6647 ( .A1(n9738), .A2(n9740), .ZN(n9766) );
  AND2_X1 U6648 ( .A1(n8139), .A2(n8138), .ZN(n9812) );
  OR2_X1 U6649 ( .A1(n6425), .A2(n8682), .ZN(n6390) );
  AND2_X1 U6650 ( .A1(n10392), .A2(n7128), .ZN(n6322) );
  INV_X1 U6651 ( .A(n8488), .ZN(n8503) );
  AND2_X1 U6652 ( .A1(n6522), .A2(n10453), .ZN(n7123) );
  OAI21_X1 U6653 ( .B1(n5193), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n5097), .ZN(
        n5098) );
  OR3_X1 U6654 ( .A1(n7343), .A2(n7708), .A3(n7577), .ZN(n6768) );
  INV_X1 U6655 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8720) );
  OR2_X1 U6656 ( .A1(n9073), .A2(n9528), .ZN(n9148) );
  AND2_X1 U6657 ( .A1(n6975), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9143) );
  INV_X1 U6658 ( .A(n9153), .ZN(n9122) );
  OR2_X1 U6659 ( .A1(n10467), .A2(n6104), .ZN(n9485) );
  AND2_X1 U6660 ( .A1(n5702), .A2(n7095), .ZN(n5703) );
  OR2_X1 U6661 ( .A1(n7025), .A2(n7024), .ZN(n7027) );
  INV_X1 U6662 ( .A(n9286), .ZN(n9263) );
  AND2_X1 U6663 ( .A1(n6775), .A2(n6773), .ZN(n9291) );
  AND2_X1 U6664 ( .A1(n6096), .A2(n6766), .ZN(n9462) );
  OR2_X1 U6665 ( .A1(n6037), .A2(n5935), .ZN(n9524) );
  INV_X1 U6666 ( .A(n9491), .ZN(n9540) );
  INV_X1 U6667 ( .A(n9495), .ZN(n9522) );
  INV_X1 U6668 ( .A(n9670), .ZN(n5975) );
  INV_X1 U6669 ( .A(n10510), .ZN(n9627) );
  OR2_X1 U6670 ( .A1(n5969), .A2(n5968), .ZN(n7314) );
  AND2_X1 U6671 ( .A1(n5948), .A2(n5947), .ZN(n10466) );
  AND2_X1 U6672 ( .A1(n8014), .A2(n7993), .ZN(n10084) );
  AND2_X1 U6673 ( .A1(n7965), .A2(n7964), .ZN(n10079) );
  OR2_X1 U6674 ( .A1(n6425), .A2(n6282), .ZN(n6415) );
  AND2_X1 U6675 ( .A1(n6266), .A2(n6257), .ZN(n10427) );
  INV_X1 U6676 ( .A(n10182), .ZN(n10147) );
  AND2_X1 U6677 ( .A1(n10071), .A2(n10307), .ZN(n10156) );
  INV_X1 U6678 ( .A(n6459), .ZN(n7195) );
  INV_X1 U6679 ( .A(n10260), .ZN(n10298) );
  AND2_X1 U6680 ( .A1(n7123), .A2(n6438), .ZN(n6605) );
  XNOR2_X1 U6681 ( .A(n5098), .B(SI_3_), .ZN(n5111) );
  INV_X1 U6682 ( .A(n8927), .ZN(n9289) );
  NAND2_X1 U6683 ( .A1(n6102), .A2(n6097), .ZN(n9138) );
  INV_X1 U6684 ( .A(n8881), .ZN(n9157) );
  INV_X1 U6685 ( .A(n9005), .ZN(n9162) );
  OR2_X1 U6686 ( .A1(n6805), .A2(n6804), .ZN(n9295) );
  NOR2_X1 U6687 ( .A1(n5040), .A2(n5964), .ZN(n5965) );
  INV_X1 U6688 ( .A(n10522), .ZN(n10519) );
  INV_X1 U6689 ( .A(n9326), .ZN(n9642) );
  INV_X1 U6690 ( .A(n9489), .ZN(n9665) );
  OR2_X1 U6691 ( .A1(n7314), .A2(n5971), .ZN(n10512) );
  INV_X1 U6692 ( .A(n10474), .ZN(n10477) );
  XNOR2_X1 U6693 ( .A(n5868), .B(n5867), .ZN(n7343) );
  INV_X1 U6694 ( .A(n9359), .ZN(n8923) );
  INV_X1 U6695 ( .A(n10214), .ZN(n9976) );
  INV_X1 U6696 ( .A(n10222), .ZN(n9747) );
  INV_X1 U6697 ( .A(n10237), .ZN(n10036) );
  INV_X1 U6698 ( .A(n9815), .ZN(n9825) );
  INV_X1 U6699 ( .A(n9994), .ZN(n9842) );
  INV_X1 U6700 ( .A(n10015), .ZN(n9844) );
  INV_X1 U6701 ( .A(n10183), .ZN(n9846) );
  OR2_X1 U6702 ( .A1(n9948), .A2(n8929), .ZN(n10416) );
  XNOR2_X1 U6703 ( .A(n9956), .B(n9955), .ZN(n10199) );
  OR2_X1 U6704 ( .A1(n10311), .A2(n6348), .ZN(n10439) );
  INV_X1 U6705 ( .A(n10448), .ZN(n10449) );
  INV_X1 U6706 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n8787) );
  NOR2_X1 U6707 ( .A1(n6501), .A2(n10561), .ZN(n10560) );
  NOR2_X1 U6708 ( .A1(n10551), .A2(n10550), .ZN(n10549) );
  AND2_X1 U6709 ( .A1(n5987), .A2(n10480), .ZN(P2_U3966) );
  NAND4_X1 U6710 ( .A1(n5867), .A2(n5668), .A3(n5456), .A4(n5695), .ZN(n5869)
         );
  INV_X1 U6711 ( .A(n5869), .ZN(n5053) );
  INV_X1 U6712 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5054) );
  NAND4_X1 U6713 ( .A1(n5055), .A2(n8561), .A3(n5054), .A4(n5404), .ZN(n5870)
         );
  NOR2_X1 U6714 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5058) );
  XNOR2_X2 U6715 ( .A(n5063), .B(n5062), .ZN(n8933) );
  MUX2_X1 U6716 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5064), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5066) );
  INV_X1 U6717 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5067) );
  NAND2_X2 U6718 ( .A1(n5069), .A2(n9683), .ZN(n5467) );
  INV_X1 U6719 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5068) );
  OR2_X1 U6720 ( .A1(n5548), .A2(n5068), .ZN(n5073) );
  NAND2_X2 U6721 ( .A1(n5069), .A2(n5070), .ZN(n5141) );
  XNOR2_X1 U6722 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8826) );
  OR2_X1 U6723 ( .A1(n5598), .A2(n8826), .ZN(n5072) );
  INV_X2 U6724 ( .A(n5175), .ZN(n5666) );
  INV_X1 U6725 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6787) );
  OR2_X1 U6726 ( .A1(n5666), .A2(n6787), .ZN(n5071) );
  AND4_X2 U6727 ( .A1(n5074), .A2(n5073), .A3(n5072), .A4(n5071), .ZN(n6866)
         );
  NAND2_X1 U6728 ( .A1(n5873), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5078) );
  NAND2_X1 U6729 ( .A1(n5164), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5082) );
  INV_X1 U6730 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5081) );
  XNOR2_X1 U6731 ( .A(n5082), .B(n5081), .ZN(n8530) );
  INV_X1 U6732 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U6733 ( .A1(n5193), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5083) );
  INV_X1 U6734 ( .A(SI_2_), .ZN(n5148) );
  OAI211_X1 U6735 ( .C1(n5193), .C2(n6183), .A(n5083), .B(n5148), .ZN(n5093)
         );
  NOR2_X1 U6736 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5086) );
  AND2_X1 U6737 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5124) );
  INV_X1 U6738 ( .A(n5124), .ZN(n5085) );
  NAND2_X1 U6739 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5084) );
  OAI21_X1 U6740 ( .B1(n5086), .B2(n5085), .A(n5084), .ZN(n5087) );
  NAND2_X1 U6741 ( .A1(n5133), .A2(n5087), .ZN(n5092) );
  NOR2_X1 U6742 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n5089) );
  NAND2_X1 U6743 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5134) );
  NAND2_X1 U6744 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n5088) );
  OAI21_X1 U6745 ( .B1(n5089), .B2(n5134), .A(n5088), .ZN(n5090) );
  NAND2_X1 U6746 ( .A1(n5193), .A2(n5090), .ZN(n5091) );
  NAND2_X1 U6747 ( .A1(n5092), .A2(n5091), .ZN(n5149) );
  NAND2_X1 U6748 ( .A1(n5093), .A2(n5149), .ZN(n5096) );
  INV_X1 U6749 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6417) );
  NAND2_X1 U6750 ( .A1(n5193), .A2(n6417), .ZN(n5094) );
  OAI211_X1 U6751 ( .C1(n6398), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n5094), .B(
        SI_2_), .ZN(n5095) );
  NAND2_X1 U6752 ( .A1(n5096), .A2(n5095), .ZN(n5110) );
  NAND2_X1 U6753 ( .A1(n5110), .A2(n5111), .ZN(n5101) );
  INV_X1 U6754 ( .A(n5098), .ZN(n5099) );
  NAND2_X1 U6755 ( .A1(n5099), .A2(SI_3_), .ZN(n5100) );
  NAND2_X1 U6756 ( .A1(n5101), .A2(n5100), .ZN(n5161) );
  MUX2_X1 U6757 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5193), .Z(n5163) );
  XNOR2_X1 U6758 ( .A(n5163), .B(SI_4_), .ZN(n5160) );
  XNOR2_X1 U6759 ( .A(n5161), .B(n5160), .ZN(n6555) );
  NAND2_X1 U6760 ( .A1(n6771), .A2(n5133), .ZN(n5157) );
  NAND2_X1 U6761 ( .A1(n6555), .A2(n5615), .ZN(n5103) );
  AND2_X2 U6762 ( .A1(n6771), .A2(n6398), .ZN(n5152) );
  NAND2_X1 U6763 ( .A1(n5152), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5102) );
  OAI211_X1 U6764 ( .C1(n6771), .C2(n8530), .A(n5103), .B(n5102), .ZN(n5104)
         );
  NAND2_X1 U6765 ( .A1(n6866), .A2(n5104), .ZN(n5716) );
  NAND2_X1 U6766 ( .A1(n5126), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5109) );
  OR2_X1 U6767 ( .A1(n5141), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5108) );
  INV_X1 U6768 ( .A(n5175), .ZN(n5105) );
  INV_X1 U6769 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6785) );
  OR2_X1 U6770 ( .A1(n5105), .A2(n6785), .ZN(n5107) );
  INV_X1 U6771 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6756) );
  XNOR2_X1 U6772 ( .A(n5111), .B(n5110), .ZN(n8175) );
  NAND2_X1 U6773 ( .A1(n5152), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5116) );
  NOR2_X1 U6774 ( .A1(n5154), .A2(n9677), .ZN(n5112) );
  MUX2_X1 U6775 ( .A(n9677), .B(n5112), .S(P2_IR_REG_3__SCAN_IN), .Z(n5114) );
  NAND2_X1 U6776 ( .A1(n5460), .A2(n9179), .ZN(n5115) );
  OAI211_X1 U6777 ( .C1(n5157), .C2(n8175), .A(n5116), .B(n5115), .ZN(n6840)
         );
  NAND2_X1 U6778 ( .A1(n6946), .A2(n6840), .ZN(n6814) );
  INV_X1 U6779 ( .A(n6814), .ZN(n5718) );
  NOR2_X1 U6780 ( .A1(n6815), .A2(n5718), .ZN(n5159) );
  NAND2_X1 U6781 ( .A1(n5175), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5121) );
  INV_X1 U6782 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n8758) );
  OR2_X1 U6783 ( .A1(n5467), .A2(n8758), .ZN(n5120) );
  INV_X1 U6784 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7555) );
  OR2_X1 U6785 ( .A1(n5141), .A2(n7555), .ZN(n5119) );
  INV_X1 U6786 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5117) );
  OR2_X1 U6787 ( .A1(n4370), .A2(n5117), .ZN(n5118) );
  AND4_X1 U6788 ( .A1(n5121), .A2(n5120), .A3(n5119), .A4(n5118), .ZN(n9530)
         );
  NAND2_X1 U6789 ( .A1(n5133), .A2(SI_0_), .ZN(n5123) );
  INV_X1 U6790 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5122) );
  NAND2_X1 U6791 ( .A1(n5123), .A2(n5122), .ZN(n5125) );
  AND2_X1 U6792 ( .A1(n5125), .A2(n5132), .ZN(n9687) );
  MUX2_X1 U6793 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9687), .S(n6771), .Z(n10481)
         );
  NAND2_X1 U6794 ( .A1(n9530), .A2(n10481), .ZN(n7554) );
  NAND2_X1 U6795 ( .A1(n5126), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5131) );
  INV_X1 U6796 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n5127) );
  OR2_X1 U6797 ( .A1(n5467), .A2(n5127), .ZN(n5130) );
  NAND2_X1 U6798 ( .A1(n5175), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5129) );
  INV_X1 U6799 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6953) );
  OR2_X1 U6800 ( .A1(n5141), .A2(n6953), .ZN(n5128) );
  INV_X1 U6801 ( .A(SI_1_), .ZN(n5135) );
  MUX2_X1 U6802 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n6398), .Z(n5136) );
  NAND2_X1 U6803 ( .A1(n4377), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5140) );
  NAND2_X1 U6804 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5138) );
  OAI211_X1 U6805 ( .C1(n5157), .C2(n6399), .A(n5140), .B(n5139), .ZN(n5941)
         );
  NAND2_X1 U6806 ( .A1(n6829), .A2(n5941), .ZN(n5845) );
  NAND2_X1 U6807 ( .A1(n7554), .A2(n5845), .ZN(n5707) );
  NAND2_X1 U6808 ( .A1(n5707), .A2(n5846), .ZN(n6826) );
  NAND2_X1 U6809 ( .A1(n5175), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5147) );
  INV_X1 U6810 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n8753) );
  OR2_X1 U6811 ( .A1(n5141), .A2(n8753), .ZN(n5146) );
  INV_X1 U6812 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6754) );
  OR2_X1 U6813 ( .A1(n5467), .A2(n6754), .ZN(n5145) );
  INV_X1 U6814 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5142) );
  XNOR2_X1 U6815 ( .A(n5149), .B(n5148), .ZN(n5151) );
  MUX2_X1 U6816 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5193), .Z(n5150) );
  XNOR2_X1 U6817 ( .A(n5151), .B(n5150), .ZN(n6418) );
  NAND2_X1 U6818 ( .A1(n5152), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5156) );
  NAND2_X1 U6819 ( .A1(n5460), .A2(n7083), .ZN(n5155) );
  OAI211_X1 U6820 ( .C1(n5157), .C2(n6418), .A(n5156), .B(n5155), .ZN(n7322)
         );
  NAND2_X1 U6821 ( .A1(n9529), .A2(n7322), .ZN(n5713) );
  NAND2_X1 U6822 ( .A1(n5713), .A2(n5711), .ZN(n6827) );
  INV_X1 U6823 ( .A(n6827), .ZN(n5847) );
  NAND2_X1 U6824 ( .A1(n5158), .A2(n5847), .ZN(n6824) );
  NAND2_X1 U6825 ( .A1(n5159), .A2(n6813), .ZN(n7526) );
  INV_X1 U6826 ( .A(n5160), .ZN(n5162) );
  NAND2_X1 U6827 ( .A1(n5163), .A2(SI_4_), .ZN(n5208) );
  MUX2_X1 U6828 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5193), .Z(n5210) );
  XNOR2_X1 U6829 ( .A(n5210), .B(SI_5_), .ZN(n5189) );
  NAND2_X1 U6830 ( .A1(n6624), .A2(n4378), .ZN(n5171) );
  NAND2_X1 U6831 ( .A1(n5166), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5165) );
  MUX2_X1 U6832 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5165), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5169) );
  INV_X1 U6833 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U6834 ( .A1(n5169), .A2(n5196), .ZN(n9197) );
  INV_X1 U6835 ( .A(n9197), .ZN(n9194) );
  AOI22_X1 U6836 ( .A1(n5152), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n5460), .B2(
        n9194), .ZN(n5170) );
  INV_X1 U6837 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6757) );
  OR2_X1 U6838 ( .A1(n5548), .A2(n6757), .ZN(n5179) );
  INV_X1 U6839 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5173) );
  NAND2_X1 U6840 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5172) );
  NAND2_X1 U6841 ( .A1(n5173), .A2(n5172), .ZN(n5174) );
  NAND2_X1 U6842 ( .A1(n5182), .A2(n5174), .ZN(n7533) );
  OR2_X1 U6843 ( .A1(n5598), .A2(n7533), .ZN(n5178) );
  INV_X1 U6844 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5176) );
  OR2_X1 U6845 ( .A1(n5105), .A2(n5176), .ZN(n5177) );
  NAND2_X1 U6846 ( .A1(n5175), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5188) );
  INV_X1 U6847 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6759) );
  OR2_X1 U6848 ( .A1(n5548), .A2(n6759), .ZN(n5187) );
  INV_X1 U6849 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8547) );
  NAND2_X1 U6850 ( .A1(n5182), .A2(n8547), .ZN(n5183) );
  NAND2_X1 U6851 ( .A1(n5201), .A2(n5183), .ZN(n7329) );
  OR2_X1 U6852 ( .A1(n5598), .A2(n7329), .ZN(n5186) );
  INV_X1 U6853 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5184) );
  OR2_X1 U6854 ( .A1(n4370), .A2(n5184), .ZN(n5185) );
  INV_X1 U6855 ( .A(n5189), .ZN(n5190) );
  NAND2_X1 U6856 ( .A1(n5191), .A2(n5190), .ZN(n5192) );
  NAND2_X1 U6857 ( .A1(n5210), .A2(SI_5_), .ZN(n5209) );
  XNOR2_X1 U6858 ( .A(n5214), .B(SI_6_), .ZN(n5212) );
  NAND2_X1 U6859 ( .A1(n6696), .A2(n4378), .ZN(n5199) );
  NAND2_X1 U6860 ( .A1(n5196), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5195) );
  MUX2_X1 U6861 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5195), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5197) );
  AND2_X1 U6862 ( .A1(n5197), .A2(n5218), .ZN(n6919) );
  AOI22_X1 U6863 ( .A1(n5152), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5460), .B2(
        n6919), .ZN(n5198) );
  NAND2_X1 U6864 ( .A1(n5199), .A2(n5198), .ZN(n7337) );
  OR2_X1 U6865 ( .A1(n7100), .A2(n7337), .ZN(n5727) );
  NAND2_X1 U6866 ( .A1(n7337), .A2(n7100), .ZN(n7475) );
  NAND2_X1 U6867 ( .A1(n5175), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5207) );
  INV_X1 U6868 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6761) );
  OR2_X1 U6869 ( .A1(n5548), .A2(n6761), .ZN(n5206) );
  INV_X1 U6870 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5200) );
  NAND2_X1 U6871 ( .A1(n5201), .A2(n5200), .ZN(n5202) );
  NAND2_X1 U6872 ( .A1(n5225), .A2(n5202), .ZN(n7480) );
  OR2_X1 U6873 ( .A1(n5598), .A2(n7480), .ZN(n5205) );
  INV_X1 U6874 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5203) );
  OR2_X1 U6875 ( .A1(n4370), .A2(n5203), .ZN(n5204) );
  NAND2_X1 U6876 ( .A1(n5231), .A2(n5046), .ZN(n5213) );
  NOR2_X1 U6877 ( .A1(n5210), .A2(SI_5_), .ZN(n5211) );
  NAND2_X1 U6878 ( .A1(n5213), .A2(n5232), .ZN(n5215) );
  NAND2_X1 U6879 ( .A1(n5214), .A2(SI_6_), .ZN(n5234) );
  XNOR2_X1 U6880 ( .A(n5238), .B(SI_7_), .ZN(n5233) );
  NAND2_X1 U6881 ( .A1(n6885), .A2(n4378), .ZN(n5221) );
  NAND2_X1 U6882 ( .A1(n5218), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5217) );
  MUX2_X1 U6883 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5217), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5219) );
  AND2_X1 U6884 ( .A1(n5219), .A2(n5313), .ZN(n9210) );
  AOI22_X1 U6885 ( .A1(n5152), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5460), .B2(
        n9210), .ZN(n5220) );
  NAND2_X1 U6886 ( .A1(n5221), .A2(n5220), .ZN(n6078) );
  OR2_X1 U6887 ( .A1(n7439), .A2(n6078), .ZN(n5736) );
  NAND2_X1 U6888 ( .A1(n7439), .A2(n6078), .ZN(n5735) );
  NAND2_X1 U6889 ( .A1(n5736), .A2(n5735), .ZN(n5851) );
  INV_X1 U6890 ( .A(n7475), .ZN(n5731) );
  NOR2_X1 U6891 ( .A1(n5851), .A2(n5731), .ZN(n5222) );
  NAND2_X1 U6892 ( .A1(n5672), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5230) );
  INV_X1 U6893 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n8597) );
  OR2_X1 U6894 ( .A1(n4370), .A2(n8597), .ZN(n5229) );
  INV_X1 U6895 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U6896 ( .A1(n5225), .A2(n5224), .ZN(n5226) );
  NAND2_X1 U6897 ( .A1(n5260), .A2(n5226), .ZN(n7453) );
  OR2_X1 U6898 ( .A1(n5598), .A2(n7453), .ZN(n5228) );
  INV_X1 U6899 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6792) );
  OR2_X1 U6900 ( .A1(n5666), .A2(n6792), .ZN(n5227) );
  NAND3_X1 U6901 ( .A1(n5231), .A2(n5046), .A3(n5234), .ZN(n5237) );
  INV_X1 U6902 ( .A(n5232), .ZN(n5235) );
  AOI21_X1 U6903 ( .B1(n5235), .B2(n5234), .A(n5233), .ZN(n5236) );
  NAND2_X1 U6904 ( .A1(n5237), .A2(n5236), .ZN(n5240) );
  NAND2_X1 U6905 ( .A1(n5238), .A2(SI_7_), .ZN(n5239) );
  NAND2_X1 U6906 ( .A1(n5240), .A2(n5239), .ZN(n5266) );
  INV_X1 U6907 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6196) );
  INV_X1 U6908 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6194) );
  INV_X1 U6909 ( .A(SI_8_), .ZN(n5241) );
  INV_X1 U6910 ( .A(n5242), .ZN(n5243) );
  NAND2_X1 U6911 ( .A1(n5243), .A2(SI_8_), .ZN(n5244) );
  XNOR2_X1 U6912 ( .A(n5266), .B(n5249), .ZN(n7041) );
  NAND2_X1 U6913 ( .A1(n7041), .A2(n4378), .ZN(n5247) );
  NAND2_X1 U6914 ( .A1(n5313), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5245) );
  XNOR2_X1 U6915 ( .A(n5245), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9223) );
  AOI22_X1 U6916 ( .A1(n5152), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5460), .B2(
        n9223), .ZN(n5246) );
  NAND2_X1 U6917 ( .A1(n7449), .A2(n7717), .ZN(n5738) );
  NAND2_X1 U6918 ( .A1(n5739), .A2(n5738), .ZN(n7435) );
  INV_X1 U6919 ( .A(n5266), .ZN(n5250) );
  NAND2_X1 U6920 ( .A1(n5250), .A2(n5267), .ZN(n5251) );
  NAND2_X1 U6921 ( .A1(n5251), .A2(n5269), .ZN(n5256) );
  INV_X1 U6922 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5252) );
  INV_X1 U6923 ( .A(SI_9_), .ZN(n5253) );
  INV_X1 U6924 ( .A(n5254), .ZN(n5255) );
  XNOR2_X1 U6925 ( .A(n5256), .B(n4405), .ZN(n7137) );
  NAND2_X1 U6926 ( .A1(n7137), .A2(n4378), .ZN(n5258) );
  XNOR2_X1 U6927 ( .A(n5277), .B(P2_IR_REG_9__SCAN_IN), .ZN(n9247) );
  AOI22_X1 U6928 ( .A1(n5460), .A2(n9247), .B1(n5152), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n5257) );
  INV_X1 U6929 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7721) );
  OR2_X1 U6930 ( .A1(n5467), .A2(n7721), .ZN(n5264) );
  NAND2_X1 U6931 ( .A1(n5260), .A2(n5259), .ZN(n5261) );
  NAND2_X1 U6932 ( .A1(n5284), .A2(n5261), .ZN(n7724) );
  OR2_X1 U6933 ( .A1(n5598), .A2(n7724), .ZN(n5263) );
  INV_X1 U6934 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8731) );
  OR2_X1 U6935 ( .A1(n5666), .A2(n8731), .ZN(n5262) );
  OR2_X1 U6936 ( .A1(n9629), .A2(n7671), .ZN(n5744) );
  INV_X1 U6937 ( .A(n5269), .ZN(n5270) );
  NAND2_X1 U6938 ( .A1(n5306), .A2(n5305), .ZN(n5290) );
  INV_X1 U6939 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6214) );
  INV_X1 U6940 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6212) );
  MUX2_X1 U6941 ( .A(n6214), .B(n6212), .S(n5627), .Z(n5273) );
  INV_X1 U6942 ( .A(SI_10_), .ZN(n5272) );
  INV_X1 U6943 ( .A(n5273), .ZN(n5274) );
  NAND2_X1 U6944 ( .A1(n5274), .A2(SI_10_), .ZN(n5275) );
  NAND2_X1 U6945 ( .A1(n7203), .A2(n4378), .ZN(n5283) );
  INV_X1 U6946 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5276) );
  AOI21_X1 U6947 ( .B1(n5277), .B2(n5276), .A(n9677), .ZN(n5278) );
  NAND2_X1 U6948 ( .A1(n5278), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5281) );
  INV_X1 U6949 ( .A(n5278), .ZN(n5280) );
  INV_X1 U6950 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5279) );
  NAND2_X1 U6951 ( .A1(n5280), .A2(n5279), .ZN(n5293) );
  AOI22_X1 U6952 ( .A1(n6796), .A2(n5460), .B1(n5152), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n5282) );
  NAND2_X1 U6953 ( .A1(n5283), .A2(n5282), .ZN(n6040) );
  INV_X1 U6954 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7676) );
  OR2_X1 U6955 ( .A1(n5548), .A2(n7676), .ZN(n5288) );
  NAND2_X1 U6956 ( .A1(n5284), .A2(n8720), .ZN(n5285) );
  NAND2_X1 U6957 ( .A1(n5297), .A2(n5285), .ZN(n7677) );
  OR2_X1 U6958 ( .A1(n5598), .A2(n7677), .ZN(n5287) );
  INV_X1 U6959 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6795) );
  OR2_X1 U6960 ( .A1(n5666), .A2(n6795), .ZN(n5286) );
  NAND2_X1 U6961 ( .A1(n5291), .A2(n5303), .ZN(n5292) );
  INV_X1 U6962 ( .A(SI_11_), .ZN(n8578) );
  XNOR2_X1 U6963 ( .A(n5292), .B(n5304), .ZN(n7249) );
  NAND2_X1 U6964 ( .A1(n7249), .A2(n4378), .ZN(n5295) );
  NAND2_X1 U6965 ( .A1(n5293), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5294) );
  INV_X1 U6966 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7689) );
  OR2_X1 U6967 ( .A1(n5548), .A2(n7689), .ZN(n5301) );
  INV_X1 U6968 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9256) );
  NAND2_X1 U6969 ( .A1(n5297), .A2(n9256), .ZN(n5298) );
  NAND2_X1 U6970 ( .A1(n5318), .A2(n5298), .ZN(n7786) );
  OR2_X1 U6971 ( .A1(n5598), .A2(n7786), .ZN(n5300) );
  INV_X1 U6972 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6798) );
  OR2_X1 U6973 ( .A1(n5666), .A2(n6798), .ZN(n5299) );
  OR2_X1 U6974 ( .A1(n6040), .A2(n7785), .ZN(n7684) );
  AND2_X1 U6975 ( .A1(n5853), .A2(n7684), .ZN(n5750) );
  NAND2_X1 U6976 ( .A1(n7685), .A2(n5750), .ZN(n7541) );
  NAND3_X1 U6977 ( .A1(n5306), .A2(n4451), .A3(n5305), .ZN(n5350) );
  AND2_X1 U6978 ( .A1(n5350), .A2(n5347), .ZN(n5307) );
  NAND2_X1 U6979 ( .A1(n5307), .A2(n5343), .ZN(n5326) );
  INV_X1 U6980 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6229) );
  INV_X1 U6981 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6227) );
  MUX2_X1 U6982 ( .A(n6229), .B(n6227), .S(n5627), .Z(n5308) );
  INV_X1 U6983 ( .A(SI_12_), .ZN(n8796) );
  NAND2_X1 U6984 ( .A1(n5308), .A2(n8796), .ZN(n5351) );
  INV_X1 U6985 ( .A(n5308), .ZN(n5309) );
  NAND2_X1 U6986 ( .A1(n5309), .A2(SI_12_), .ZN(n5344) );
  NAND2_X1 U6987 ( .A1(n5351), .A2(n5344), .ZN(n5325) );
  XNOR2_X1 U6988 ( .A(n5326), .B(n5325), .ZN(n7488) );
  NAND2_X1 U6989 ( .A1(n7488), .A2(n4378), .ZN(n5316) );
  NAND2_X1 U6990 ( .A1(n5311), .A2(n5310), .ZN(n5312) );
  NAND2_X1 U6991 ( .A1(n5332), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5314) );
  XNOR2_X1 U6992 ( .A(n5314), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6800) );
  AOI22_X1 U6993 ( .A1(n5460), .A2(n6800), .B1(n5152), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n5315) );
  INV_X1 U6994 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n5317) );
  OR2_X1 U6995 ( .A1(n5548), .A2(n5317), .ZN(n5322) );
  INV_X1 U6996 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8742) );
  NAND2_X1 U6997 ( .A1(n5318), .A2(n8742), .ZN(n5319) );
  NAND2_X1 U6998 ( .A1(n5336), .A2(n5319), .ZN(n7547) );
  OR2_X1 U6999 ( .A1(n5598), .A2(n7547), .ZN(n5321) );
  INV_X1 U7000 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8788) );
  OR2_X1 U7001 ( .A1(n5666), .A2(n8788), .ZN(n5320) );
  NAND2_X1 U7002 ( .A1(n7700), .A2(n9086), .ZN(n5747) );
  NAND3_X1 U7003 ( .A1(n7541), .A2(n5747), .A3(n7540), .ZN(n5324) );
  OR2_X1 U7004 ( .A1(n7700), .A2(n9086), .ZN(n5748) );
  NAND2_X1 U7005 ( .A1(n5324), .A2(n5748), .ZN(n7743) );
  OAI21_X1 U7006 ( .B1(n5326), .B2(n5325), .A(n5351), .ZN(n5331) );
  INV_X1 U7007 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6236) );
  INV_X1 U7008 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n8776) );
  MUX2_X1 U7009 ( .A(n6236), .B(n8776), .S(n5627), .Z(n5328) );
  INV_X1 U7010 ( .A(SI_13_), .ZN(n5327) );
  INV_X1 U7011 ( .A(n5328), .ZN(n5329) );
  NAND2_X1 U7012 ( .A1(n5329), .A2(SI_13_), .ZN(n5330) );
  XNOR2_X1 U7013 ( .A(n5331), .B(n5355), .ZN(n7617) );
  NAND2_X1 U7014 ( .A1(n7617), .A2(n4378), .ZN(n5334) );
  OAI21_X1 U7015 ( .B1(n5332), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5359) );
  XNOR2_X1 U7016 ( .A(n5359), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6983) );
  AOI22_X1 U7017 ( .A1(n6983), .A2(n5460), .B1(n5152), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n5333) );
  INV_X1 U7018 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7749) );
  OR2_X1 U7019 ( .A1(n5548), .A2(n7749), .ZN(n5340) );
  INV_X1 U7020 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5335) );
  NAND2_X1 U7021 ( .A1(n5336), .A2(n5335), .ZN(n5337) );
  NAND2_X1 U7022 ( .A1(n5368), .A2(n5337), .ZN(n9083) );
  OR2_X1 U7023 ( .A1(n5598), .A2(n9083), .ZN(n5339) );
  INV_X1 U7024 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8645) );
  OR2_X1 U7025 ( .A1(n5666), .A2(n8645), .ZN(n5338) );
  OR2_X1 U7026 ( .A1(n7805), .A2(n8975), .ZN(n5764) );
  NAND2_X1 U7027 ( .A1(n7805), .A2(n8975), .ZN(n7764) );
  NAND2_X1 U7028 ( .A1(n5764), .A2(n7764), .ZN(n7742) );
  INV_X1 U7029 ( .A(n7742), .ZN(n5342) );
  INV_X1 U7030 ( .A(n7764), .ZN(n5374) );
  NAND2_X1 U7031 ( .A1(n5344), .A2(n5343), .ZN(n5345) );
  NAND2_X1 U7032 ( .A1(n5350), .A2(n5349), .ZN(n5357) );
  INV_X1 U7033 ( .A(n5352), .ZN(n5353) );
  INV_X1 U7034 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6224) );
  MUX2_X1 U7035 ( .A(n6224), .B(n8787), .S(n5627), .Z(n5377) );
  XNOR2_X1 U7036 ( .A(n5380), .B(n5376), .ZN(n7855) );
  NAND2_X1 U7037 ( .A1(n7855), .A2(n4378), .ZN(n5365) );
  INV_X1 U7038 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5358) );
  NAND2_X1 U7039 ( .A1(n5359), .A2(n5358), .ZN(n5360) );
  NAND2_X1 U7040 ( .A1(n5360), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U7041 ( .A1(n5362), .A2(n5361), .ZN(n5384) );
  OR2_X1 U7042 ( .A1(n5362), .A2(n5361), .ZN(n5363) );
  AOI22_X1 U7043 ( .A1(n6992), .A2(n5460), .B1(n5152), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5364) );
  NAND2_X1 U7044 ( .A1(n5365), .A2(n5364), .ZN(n7772) );
  INV_X1 U7045 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5367) );
  NAND2_X1 U7046 ( .A1(n5368), .A2(n5367), .ZN(n5369) );
  NAND2_X1 U7047 ( .A1(n5388), .A2(n5369), .ZN(n7773) );
  OR2_X1 U7048 ( .A1(n7773), .A2(n5598), .ZN(n5373) );
  INV_X1 U7049 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7179) );
  OR2_X1 U7050 ( .A1(n5467), .A2(n7179), .ZN(n5371) );
  INV_X1 U7051 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8744) );
  OR2_X1 U7052 ( .A1(n5666), .A2(n8744), .ZN(n5370) );
  NAND4_X1 U7053 ( .A1(n5373), .A2(n5372), .A3(n5371), .A4(n5370), .ZN(n9167)
         );
  INV_X1 U7054 ( .A(n9167), .ZN(n9146) );
  NAND2_X1 U7055 ( .A1(n7772), .A2(n9146), .ZN(n5766) );
  NAND2_X1 U7056 ( .A1(n5767), .A2(n5766), .ZN(n5903) );
  NOR2_X1 U7057 ( .A1(n5374), .A2(n5903), .ZN(n5375) );
  INV_X1 U7058 ( .A(n5377), .ZN(n5378) );
  INV_X1 U7059 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n8635) );
  INV_X1 U7060 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6245) );
  MUX2_X1 U7061 ( .A(n8635), .B(n6245), .S(n5627), .Z(n5381) );
  INV_X1 U7062 ( .A(SI_15_), .ZN(n8598) );
  NAND2_X1 U7063 ( .A1(n5381), .A2(n8598), .ZN(n5416) );
  INV_X1 U7064 ( .A(n5381), .ZN(n5382) );
  NAND2_X1 U7065 ( .A1(n5382), .A2(SI_15_), .ZN(n5383) );
  XNOR2_X1 U7066 ( .A(n5394), .B(n5395), .ZN(n7858) );
  NAND2_X1 U7067 ( .A1(n7858), .A2(n4378), .ZN(n5387) );
  NAND2_X1 U7068 ( .A1(n5384), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5385) );
  XNOR2_X1 U7069 ( .A(n5385), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7597) );
  AOI22_X1 U7070 ( .A1(n7597), .A2(n5460), .B1(n5689), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5386) );
  INV_X1 U7071 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9147) );
  NAND2_X1 U7072 ( .A1(n5388), .A2(n9147), .ZN(n5389) );
  NAND2_X1 U7073 ( .A1(n5410), .A2(n5389), .ZN(n7800) );
  NAND2_X1 U7074 ( .A1(n5672), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5390) );
  AND2_X1 U7075 ( .A1(n5391), .A2(n5390), .ZN(n5393) );
  NAND2_X1 U7076 ( .A1(n5175), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5392) );
  OAI211_X1 U7077 ( .C1(n7800), .C2(n5598), .A(n5393), .B(n5392), .ZN(n9166)
         );
  INV_X1 U7078 ( .A(n9154), .ZN(n9618) );
  INV_X1 U7079 ( .A(n9166), .ZN(n9137) );
  NAND2_X1 U7080 ( .A1(n9618), .A2(n9137), .ZN(n5775) );
  INV_X1 U7081 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n8782) );
  INV_X1 U7082 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6265) );
  MUX2_X1 U7083 ( .A(n8782), .B(n6265), .S(n5627), .Z(n5398) );
  INV_X1 U7084 ( .A(SI_16_), .ZN(n5397) );
  NAND2_X1 U7085 ( .A1(n5398), .A2(n5397), .ZN(n5415) );
  INV_X1 U7086 ( .A(n5398), .ZN(n5399) );
  AND2_X1 U7087 ( .A1(n5415), .A2(n5418), .ZN(n5400) );
  NAND2_X1 U7088 ( .A1(n7864), .A2(n4378), .ZN(n5409) );
  NOR2_X1 U7089 ( .A1(n5405), .A2(n9677), .ZN(n5403) );
  MUX2_X1 U7090 ( .A(n9677), .B(n5403), .S(P2_IR_REG_16__SCAN_IN), .Z(n5407)
         );
  NOR2_X1 U7091 ( .A1(n5407), .A2(n5406), .ZN(n8902) );
  AOI22_X1 U7092 ( .A1(n5689), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5460), .B2(
        n8902), .ZN(n5408) );
  NAND2_X1 U7093 ( .A1(n5410), .A2(n4656), .ZN(n5411) );
  NAND2_X1 U7094 ( .A1(n5424), .A2(n5411), .ZN(n9045) );
  OR2_X1 U7095 ( .A1(n9045), .A2(n5598), .ZN(n5414) );
  NAND2_X1 U7096 ( .A1(n5175), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5412) );
  OR2_X1 U7097 ( .A1(n9047), .A2(n9499), .ZN(n5773) );
  INV_X1 U7098 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6487) );
  INV_X1 U7099 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6495) );
  MUX2_X1 U7100 ( .A(n6487), .B(n6495), .S(n5627), .Z(n5431) );
  XNOR2_X1 U7101 ( .A(n5419), .B(n5429), .ZN(n7861) );
  NAND2_X1 U7102 ( .A1(n7861), .A2(n4378), .ZN(n5423) );
  MUX2_X1 U7103 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5420), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5421) );
  AND2_X1 U7104 ( .A1(n5421), .A2(n5435), .ZN(n8908) );
  AOI22_X1 U7105 ( .A1(n5689), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5460), .B2(
        n8908), .ZN(n5422) );
  INV_X1 U7106 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9271) );
  NAND2_X1 U7107 ( .A1(n5424), .A2(n9271), .ZN(n5425) );
  AND2_X1 U7108 ( .A1(n5440), .A2(n5425), .ZN(n9511) );
  INV_X1 U7109 ( .A(n5598), .ZN(n5654) );
  INV_X1 U7110 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8912) );
  NAND2_X1 U7111 ( .A1(n5175), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5426) );
  OAI211_X1 U7112 ( .C1(n5548), .C2(n8912), .A(n5427), .B(n5426), .ZN(n5428)
         );
  AOI21_X1 U7113 ( .B1(n9511), .B2(n5654), .A(n5428), .ZN(n9479) );
  NAND2_X1 U7114 ( .A1(n9512), .A2(n9479), .ZN(n5779) );
  INV_X1 U7115 ( .A(n5431), .ZN(n5432) );
  MUX2_X1 U7116 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5627), .Z(n5451) );
  XNOR2_X1 U7117 ( .A(n5450), .B(n5448), .ZN(n7868) );
  NAND2_X1 U7118 ( .A1(n7868), .A2(n4378), .ZN(n5438) );
  NAND2_X1 U7119 ( .A1(n5435), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5436) );
  XNOR2_X1 U7120 ( .A(n5436), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8913) );
  AOI22_X1 U7121 ( .A1(n5689), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5460), .B2(
        n8913), .ZN(n5437) );
  NAND2_X1 U7122 ( .A1(n5440), .A2(n4653), .ZN(n5441) );
  NAND2_X1 U7123 ( .A1(n5463), .A2(n5441), .ZN(n9486) );
  OR2_X1 U7124 ( .A1(n9486), .A2(n5598), .ZN(n5446) );
  INV_X1 U7125 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9487) );
  NAND2_X1 U7126 ( .A1(n5175), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5442) );
  OAI211_X1 U7127 ( .C1(n5548), .C2(n9487), .A(n5443), .B(n5442), .ZN(n5444)
         );
  INV_X1 U7128 ( .A(n5444), .ZN(n5445) );
  OR2_X1 U7129 ( .A1(n9489), .A2(n9500), .ZN(n5788) );
  NAND2_X1 U7130 ( .A1(n9489), .A2(n9500), .ZN(n5787) );
  NAND2_X1 U7131 ( .A1(n5788), .A2(n5787), .ZN(n9475) );
  INV_X1 U7132 ( .A(n9475), .ZN(n9471) );
  AND2_X1 U7133 ( .A1(n9473), .A2(n9471), .ZN(n5447) );
  NAND2_X1 U7134 ( .A1(n9474), .A2(n5447), .ZN(n9478) );
  NAND2_X1 U7135 ( .A1(n9478), .A2(n5787), .ZN(n9460) );
  NAND2_X1 U7136 ( .A1(n5451), .A2(SI_18_), .ZN(n5452) );
  INV_X1 U7137 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6683) );
  INV_X1 U7138 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6685) );
  MUX2_X1 U7139 ( .A(n6683), .B(n6685), .S(n6398), .Z(n5453) );
  INV_X1 U7140 ( .A(SI_19_), .ZN(n8601) );
  NAND2_X1 U7141 ( .A1(n5453), .A2(n8601), .ZN(n5489) );
  INV_X1 U7142 ( .A(n5453), .ZN(n5454) );
  NAND2_X1 U7143 ( .A1(n5454), .A2(SI_19_), .ZN(n5455) );
  NAND2_X1 U7144 ( .A1(n5489), .A2(n5455), .ZN(n5472) );
  XNOR2_X1 U7145 ( .A(n5471), .B(n5472), .ZN(n7871) );
  NAND2_X1 U7146 ( .A1(n7871), .A2(n4378), .ZN(n5462) );
  NAND2_X1 U7147 ( .A1(n5457), .A2(n5456), .ZN(n5667) );
  NAND2_X1 U7148 ( .A1(n5667), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U7149 ( .A1(n5458), .A2(n8561), .ZN(n5697) );
  OR2_X1 U7150 ( .A1(n5458), .A2(n8561), .ZN(n5459) );
  AOI22_X1 U7151 ( .A1(n5689), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5460), .B2(
        n9359), .ZN(n5461) );
  INV_X1 U7152 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U7153 ( .A1(n5463), .A2(n6163), .ZN(n5464) );
  AND2_X1 U7154 ( .A1(n5481), .A2(n5464), .ZN(n6164) );
  NAND2_X1 U7155 ( .A1(n6164), .A2(n5636), .ZN(n5470) );
  INV_X1 U7156 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8916) );
  NAND2_X1 U7157 ( .A1(n5175), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5465) );
  OAI211_X1 U7158 ( .C1(n5467), .C2(n8916), .A(n5466), .B(n5465), .ZN(n5468)
         );
  INV_X1 U7159 ( .A(n5468), .ZN(n5469) );
  OR2_X1 U7160 ( .A1(n9595), .A2(n9480), .ZN(n5789) );
  NAND2_X1 U7161 ( .A1(n9595), .A2(n9480), .ZN(n9419) );
  NAND2_X1 U7162 ( .A1(n5491), .A2(n5489), .ZN(n5478) );
  INV_X1 U7163 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8730) );
  INV_X1 U7164 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7877) );
  MUX2_X1 U7165 ( .A(n8730), .B(n7877), .S(n5627), .Z(n5475) );
  INV_X1 U7166 ( .A(SI_20_), .ZN(n8607) );
  NAND2_X1 U7167 ( .A1(n5475), .A2(n8607), .ZN(n5488) );
  INV_X1 U7168 ( .A(n5475), .ZN(n5476) );
  NAND2_X1 U7169 ( .A1(n5476), .A2(SI_20_), .ZN(n5511) );
  AND2_X1 U7170 ( .A1(n5488), .A2(n5511), .ZN(n5477) );
  NAND2_X1 U7171 ( .A1(n7876), .A2(n4378), .ZN(n5480) );
  NAND2_X1 U7172 ( .A1(n5689), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U7173 ( .A1(n5481), .A2(n4654), .ZN(n5482) );
  NAND2_X1 U7174 ( .A1(n5496), .A2(n5482), .ZN(n9434) );
  OR2_X1 U7175 ( .A1(n9434), .A2(n5598), .ZN(n5487) );
  INV_X1 U7176 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9659) );
  NAND2_X1 U7177 ( .A1(n5175), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U7178 ( .A1(n5672), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5483) );
  OAI211_X1 U7179 ( .C1(n4370), .C2(n9659), .A(n5484), .B(n5483), .ZN(n5485)
         );
  INV_X1 U7180 ( .A(n5485), .ZN(n5486) );
  AND2_X1 U7181 ( .A1(n5516), .A2(n5511), .ZN(n5492) );
  INV_X1 U7182 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8795) );
  INV_X1 U7183 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8629) );
  MUX2_X1 U7184 ( .A(n8795), .B(n8629), .S(n5627), .Z(n5509) );
  XNOR2_X1 U7185 ( .A(n5509), .B(SI_21_), .ZN(n5512) );
  NAND2_X1 U7186 ( .A1(n7880), .A2(n4378), .ZN(n5494) );
  NAND2_X1 U7187 ( .A1(n5689), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5493) );
  INV_X1 U7188 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U7189 ( .A1(n5496), .A2(n5495), .ZN(n5497) );
  NAND2_X1 U7190 ( .A1(n5524), .A2(n5497), .ZN(n9415) );
  OR2_X1 U7191 ( .A1(n9415), .A2(n5598), .ZN(n5502) );
  INV_X1 U7192 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9587) );
  NAND2_X1 U7193 ( .A1(n5672), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5499) );
  OAI211_X1 U7194 ( .C1(n5666), .C2(n9587), .A(n5499), .B(n5498), .ZN(n5500)
         );
  INV_X1 U7195 ( .A(n5500), .ZN(n5501) );
  NAND2_X1 U7196 ( .A1(n5502), .A2(n5501), .ZN(n9163) );
  XNOR2_X1 U7197 ( .A(n9414), .B(n9163), .ZN(n9424) );
  AND2_X1 U7198 ( .A1(n9461), .A2(n5503), .ZN(n5507) );
  INV_X1 U7199 ( .A(n5503), .ZN(n5504) );
  INV_X1 U7200 ( .A(n9424), .ZN(n5505) );
  NAND2_X1 U7201 ( .A1(n9433), .A2(n9004), .ZN(n9421) );
  INV_X1 U7202 ( .A(n9163), .ZN(n9107) );
  NAND2_X1 U7203 ( .A1(n9414), .A2(n9107), .ZN(n5796) );
  INV_X1 U7204 ( .A(n5509), .ZN(n5510) );
  NAND2_X1 U7205 ( .A1(n5510), .A2(SI_21_), .ZN(n5514) );
  INV_X1 U7206 ( .A(n5512), .ZN(n5513) );
  INV_X1 U7207 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8965) );
  INV_X1 U7208 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8961) );
  MUX2_X1 U7209 ( .A(n8965), .B(n8961), .S(n5627), .Z(n5518) );
  INV_X1 U7210 ( .A(SI_22_), .ZN(n5517) );
  NAND2_X1 U7211 ( .A1(n5518), .A2(n5517), .ZN(n5533) );
  INV_X1 U7212 ( .A(n5518), .ZN(n5519) );
  NAND2_X1 U7213 ( .A1(n5519), .A2(SI_22_), .ZN(n5520) );
  NAND2_X1 U7214 ( .A1(n5533), .A2(n5520), .ZN(n5534) );
  XNOR2_X1 U7215 ( .A(n5535), .B(n5534), .ZN(n8959) );
  NAND2_X1 U7216 ( .A1(n8959), .A2(n4378), .ZN(n5522) );
  NAND2_X1 U7217 ( .A1(n5689), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5521) );
  INV_X1 U7218 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n5523) );
  NAND2_X1 U7219 ( .A1(n5524), .A2(n5523), .ZN(n5525) );
  NAND2_X1 U7220 ( .A1(n5544), .A2(n5525), .ZN(n9403) );
  INV_X1 U7221 ( .A(n9403), .ZN(n5526) );
  NAND2_X1 U7222 ( .A1(n5526), .A2(n5636), .ZN(n5532) );
  INV_X1 U7223 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U7224 ( .A1(n5672), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5528) );
  OAI211_X1 U7225 ( .C1(n5666), .C2(n5529), .A(n5528), .B(n5527), .ZN(n5530)
         );
  INV_X1 U7226 ( .A(n5530), .ZN(n5531) );
  NAND2_X1 U7227 ( .A1(n9580), .A2(n9005), .ZN(n5801) );
  NAND2_X1 U7228 ( .A1(n9389), .A2(n5801), .ZN(n9404) );
  INV_X1 U7229 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5536) );
  INV_X1 U7230 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7886) );
  MUX2_X1 U7231 ( .A(n5536), .B(n7886), .S(n5627), .Z(n5538) );
  INV_X1 U7232 ( .A(SI_23_), .ZN(n5537) );
  NAND2_X1 U7233 ( .A1(n5538), .A2(n5537), .ZN(n5556) );
  INV_X1 U7234 ( .A(n5538), .ZN(n5539) );
  NAND2_X1 U7235 ( .A1(n5539), .A2(SI_23_), .ZN(n5540) );
  NAND2_X1 U7236 ( .A1(n7885), .A2(n4378), .ZN(n5542) );
  NAND2_X1 U7237 ( .A1(n5689), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5541) );
  INV_X1 U7238 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5543) );
  NAND2_X1 U7239 ( .A1(n5544), .A2(n5543), .ZN(n5545) );
  NAND2_X1 U7240 ( .A1(n5561), .A2(n5545), .ZN(n9384) );
  OR2_X1 U7241 ( .A1(n9384), .A2(n5598), .ZN(n5551) );
  INV_X1 U7242 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8647) );
  NAND2_X1 U7243 ( .A1(n5175), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5546) );
  OAI211_X1 U7244 ( .C1(n5548), .C2(n8647), .A(n5547), .B(n5546), .ZN(n5549)
         );
  INV_X1 U7245 ( .A(n5549), .ZN(n5550) );
  OR2_X1 U7246 ( .A1(n9383), .A2(n9108), .ZN(n5803) );
  NAND2_X1 U7247 ( .A1(n9383), .A2(n9108), .ZN(n5806) );
  NAND2_X1 U7248 ( .A1(n5803), .A2(n5806), .ZN(n5802) );
  INV_X1 U7249 ( .A(n9389), .ZN(n5552) );
  NOR2_X1 U7250 ( .A1(n5802), .A2(n5552), .ZN(n5553) );
  NAND2_X1 U7251 ( .A1(n5555), .A2(n5554), .ZN(n5557) );
  INV_X1 U7252 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7341) );
  INV_X1 U7253 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7890) );
  MUX2_X1 U7254 ( .A(n7341), .B(n7890), .S(n5627), .Z(n5569) );
  XNOR2_X1 U7255 ( .A(n5569), .B(SI_24_), .ZN(n5568) );
  XNOR2_X1 U7256 ( .A(n5573), .B(n5568), .ZN(n7889) );
  NAND2_X1 U7257 ( .A1(n7889), .A2(n4378), .ZN(n5559) );
  NAND2_X1 U7258 ( .A1(n5689), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5558) );
  INV_X1 U7259 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8581) );
  NAND2_X1 U7260 ( .A1(n5561), .A2(n8581), .ZN(n5562) );
  NAND2_X1 U7261 ( .A1(n5579), .A2(n5562), .ZN(n9368) );
  INV_X1 U7262 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8560) );
  NAND2_X1 U7263 ( .A1(n5672), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5564) );
  OAI211_X1 U7264 ( .C1(n5105), .C2(n8560), .A(n5564), .B(n5563), .ZN(n5565)
         );
  INV_X1 U7265 ( .A(n5565), .ZN(n5566) );
  NAND2_X1 U7266 ( .A1(n9570), .A2(n8983), .ZN(n5808) );
  INV_X1 U7267 ( .A(n5568), .ZN(n5572) );
  INV_X1 U7268 ( .A(n5569), .ZN(n5570) );
  NAND2_X1 U7269 ( .A1(n5570), .A2(SI_24_), .ZN(n5571) );
  INV_X1 U7270 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7578) );
  INV_X1 U7271 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7895) );
  MUX2_X1 U7272 ( .A(n7578), .B(n7895), .S(n5627), .Z(n5574) );
  INV_X1 U7273 ( .A(SI_25_), .ZN(n8797) );
  NAND2_X1 U7274 ( .A1(n5574), .A2(n8797), .ZN(n5607) );
  INV_X1 U7275 ( .A(n5574), .ZN(n5575) );
  NAND2_X1 U7276 ( .A1(n5575), .A2(SI_25_), .ZN(n5576) );
  NAND2_X1 U7277 ( .A1(n5607), .A2(n5576), .ZN(n5586) );
  NAND2_X1 U7278 ( .A1(n7894), .A2(n4378), .ZN(n5578) );
  NAND2_X1 U7279 ( .A1(n5689), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5577) );
  INV_X1 U7280 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9029) );
  NAND2_X1 U7281 ( .A1(n5579), .A2(n9029), .ZN(n5580) );
  INV_X1 U7282 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8632) );
  NAND2_X1 U7283 ( .A1(n5672), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5581) );
  OAI211_X1 U7284 ( .C1(n8632), .C2(n5666), .A(n5582), .B(n5581), .ZN(n5583)
         );
  NAND2_X1 U7285 ( .A1(n9566), .A2(n9128), .ZN(n5812) );
  INV_X1 U7286 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7706) );
  INV_X1 U7287 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7899) );
  MUX2_X1 U7288 ( .A(n7706), .B(n7899), .S(n5627), .Z(n5589) );
  INV_X1 U7289 ( .A(SI_26_), .ZN(n5588) );
  NAND2_X1 U7290 ( .A1(n5589), .A2(n5588), .ZN(n5606) );
  INV_X1 U7291 ( .A(n5589), .ZN(n5590) );
  NAND2_X1 U7292 ( .A1(n5590), .A2(SI_26_), .ZN(n5608) );
  AND2_X1 U7293 ( .A1(n5606), .A2(n5608), .ZN(n5591) );
  NAND2_X1 U7294 ( .A1(n7898), .A2(n4378), .ZN(n5594) );
  NAND2_X1 U7295 ( .A1(n5689), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5593) );
  INV_X1 U7296 ( .A(n5596), .ZN(n5595) );
  INV_X1 U7297 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9130) );
  NAND2_X1 U7298 ( .A1(n5596), .A2(n9130), .ZN(n5597) );
  NAND2_X1 U7299 ( .A1(n5634), .A2(n5597), .ZN(n9343) );
  INV_X1 U7300 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9562) );
  NAND2_X1 U7301 ( .A1(n5672), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5599) );
  OAI211_X1 U7302 ( .C1(n9562), .C2(n5666), .A(n5600), .B(n5599), .ZN(n5601)
         );
  INV_X1 U7303 ( .A(n5601), .ZN(n5602) );
  INV_X1 U7304 ( .A(n5811), .ZN(n9337) );
  NOR2_X1 U7305 ( .A1(n9336), .A2(n9337), .ZN(n5604) );
  AND2_X1 U7306 ( .A1(n5607), .A2(n5606), .ZN(n5609) );
  INV_X1 U7307 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7759) );
  INV_X1 U7308 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7904) );
  MUX2_X1 U7309 ( .A(n7759), .B(n7904), .S(n5627), .Z(n5612) );
  INV_X1 U7310 ( .A(SI_27_), .ZN(n5611) );
  NAND2_X1 U7311 ( .A1(n5612), .A2(n5611), .ZN(n5625) );
  INV_X1 U7312 ( .A(n5612), .ZN(n5613) );
  NAND2_X1 U7313 ( .A1(n5613), .A2(SI_27_), .ZN(n5614) );
  AND2_X1 U7314 ( .A1(n5625), .A2(n5614), .ZN(n5623) );
  NAND2_X1 U7315 ( .A1(n7903), .A2(n4378), .ZN(n5617) );
  NAND2_X1 U7316 ( .A1(n5689), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5616) );
  XNOR2_X1 U7317 ( .A(n5634), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n9327) );
  INV_X1 U7318 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9557) );
  NAND2_X1 U7319 ( .A1(n5672), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5619) );
  OAI211_X1 U7320 ( .C1(n9557), .C2(n5666), .A(n5619), .B(n5618), .ZN(n5620)
         );
  NAND2_X1 U7321 ( .A1(n9326), .A2(n9129), .ZN(n5822) );
  INV_X1 U7322 ( .A(n9320), .ZN(n5621) );
  NOR2_X1 U7323 ( .A1(n9315), .A2(n5621), .ZN(n5622) );
  NAND2_X1 U7324 ( .A1(n9318), .A2(n5622), .ZN(n9317) );
  INV_X1 U7325 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5628) );
  INV_X1 U7326 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8930) );
  MUX2_X1 U7327 ( .A(n5628), .B(n8930), .S(n5627), .Z(n5646) );
  XNOR2_X1 U7328 ( .A(n5646), .B(SI_28_), .ZN(n5643) );
  NAND2_X1 U7329 ( .A1(n5689), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5629) );
  INV_X1 U7330 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5632) );
  INV_X1 U7331 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5631) );
  OAI21_X1 U7332 ( .B1(n5634), .B2(n5632), .A(n5631), .ZN(n5635) );
  NAND2_X1 U7333 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n5633) );
  NAND2_X1 U7334 ( .A1(n8892), .A2(n5636), .ZN(n5642) );
  INV_X1 U7335 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8789) );
  INV_X1 U7336 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n5637) );
  OR2_X1 U7337 ( .A1(n5548), .A2(n5637), .ZN(n5638) );
  OAI211_X1 U7338 ( .C1(n8789), .C2(n5105), .A(n5639), .B(n5638), .ZN(n5640)
         );
  INV_X1 U7339 ( .A(n5640), .ZN(n5641) );
  NAND2_X1 U7340 ( .A1(n9548), .A2(n8881), .ZN(n5826) );
  INV_X1 U7341 ( .A(SI_28_), .ZN(n5645) );
  NAND2_X1 U7342 ( .A1(n5646), .A2(n5645), .ZN(n5647) );
  INV_X1 U7343 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9685) );
  INV_X1 U7344 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10349) );
  MUX2_X1 U7345 ( .A(n9685), .B(n10349), .S(n6398), .Z(n5657) );
  XNOR2_X1 U7346 ( .A(n5657), .B(SI_29_), .ZN(n5648) );
  NAND2_X1 U7347 ( .A1(n9682), .A2(n4378), .ZN(n5650) );
  NAND2_X1 U7348 ( .A1(n5689), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5649) );
  INV_X1 U7349 ( .A(n9307), .ZN(n5655) );
  INV_X1 U7350 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8765) );
  NAND2_X1 U7351 ( .A1(n5672), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5651) );
  OAI211_X1 U7352 ( .C1(n8765), .C2(n5666), .A(n5652), .B(n5651), .ZN(n5653)
         );
  AOI21_X1 U7353 ( .B1(n5655), .B2(n5654), .A(n5653), .ZN(n7844) );
  NAND2_X1 U7354 ( .A1(n9308), .A2(n7844), .ZN(n5833) );
  NAND2_X1 U7355 ( .A1(n5656), .A2(n5832), .ZN(n5675) );
  INV_X1 U7356 ( .A(n5657), .ZN(n5658) );
  NAND2_X1 U7357 ( .A1(n5658), .A2(SI_29_), .ZN(n5659) );
  MUX2_X1 U7358 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n6398), .Z(n5679) );
  XNOR2_X1 U7359 ( .A(n5679), .B(SI_30_), .ZN(n5661) );
  NAND2_X1 U7360 ( .A1(n8931), .A2(n4378), .ZN(n5663) );
  NAND2_X1 U7361 ( .A1(n5689), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n5662) );
  INV_X1 U7362 ( .A(n9638), .ZN(n5693) );
  INV_X1 U7363 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9546) );
  NAND2_X1 U7364 ( .A1(n5672), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5665) );
  OAI211_X1 U7365 ( .C1(n5666), .C2(n9546), .A(n5665), .B(n5664), .ZN(n9155)
         );
  INV_X1 U7366 ( .A(n5667), .ZN(n5669) );
  INV_X1 U7367 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5668) );
  NAND3_X1 U7368 ( .A1(n5669), .A2(n5668), .A3(n8561), .ZN(n5696) );
  NAND2_X1 U7369 ( .A1(n5696), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5671) );
  INV_X1 U7370 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5670) );
  INV_X1 U7371 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7372 ( .A1(n5672), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5674) );
  OAI211_X1 U7373 ( .C1(n5105), .C2(n5981), .A(n5674), .B(n5673), .ZN(n6241)
         );
  INV_X1 U7374 ( .A(n5678), .ZN(n5677) );
  INV_X1 U7375 ( .A(SI_30_), .ZN(n5676) );
  INV_X1 U7376 ( .A(n5679), .ZN(n5680) );
  NAND2_X1 U7377 ( .A1(n5681), .A2(n5680), .ZN(n5682) );
  NAND2_X1 U7378 ( .A1(n5683), .A2(n5682), .ZN(n5688) );
  INV_X1 U7379 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5685) );
  INV_X1 U7380 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5684) );
  MUX2_X1 U7381 ( .A(n5685), .B(n5684), .S(n6398), .Z(n5686) );
  XNOR2_X1 U7382 ( .A(n5686), .B(SI_31_), .ZN(n5687) );
  NAND2_X1 U7383 ( .A1(n9675), .A2(n4378), .ZN(n5691) );
  NAND2_X1 U7384 ( .A1(n5689), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n5690) );
  INV_X1 U7385 ( .A(n6241), .ZN(n5694) );
  OR2_X1 U7386 ( .A1(n5982), .A2(n5694), .ZN(n5842) );
  INV_X1 U7387 ( .A(n9155), .ZN(n5692) );
  NAND2_X1 U7388 ( .A1(n5693), .A2(n5692), .ZN(n5834) );
  NAND2_X1 U7389 ( .A1(n5697), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5698) );
  AND2_X1 U7390 ( .A1(n5931), .A2(n5879), .ZN(n5935) );
  OR2_X1 U7391 ( .A1(n8880), .A2(n5935), .ZN(n5702) );
  NAND2_X1 U7392 ( .A1(n5699), .A2(n5695), .ZN(n5700) );
  NAND2_X1 U7393 ( .A1(n5700), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5865) );
  INV_X1 U7394 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5864) );
  XNOR2_X1 U7395 ( .A(n5865), .B(n5864), .ZN(n6105) );
  INV_X1 U7396 ( .A(n6105), .ZN(n5701) );
  AND2_X1 U7397 ( .A1(n5701), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7095) );
  NAND2_X1 U7398 ( .A1(n5704), .A2(n5703), .ZN(n5882) );
  INV_X1 U7399 ( .A(n9352), .ZN(n5810) );
  AND2_X1 U7400 ( .A1(n5879), .A2(n9359), .ZN(n5705) );
  INV_X1 U7401 ( .A(n9530), .ZN(n6976) );
  INV_X1 U7402 ( .A(n10481), .ZN(n7018) );
  NAND2_X1 U7403 ( .A1(n6976), .A2(n7018), .ZN(n7553) );
  AND2_X1 U7404 ( .A1(n7553), .A2(n5879), .ZN(n5706) );
  OAI211_X1 U7405 ( .C1(n5707), .C2(n5706), .A(n5711), .B(n5846), .ZN(n5708)
         );
  NAND3_X1 U7406 ( .A1(n5708), .A2(n5713), .A3(n5841), .ZN(n5709) );
  NAND3_X1 U7407 ( .A1(n5717), .A2(n6842), .A3(n5709), .ZN(n5721) );
  NAND2_X1 U7408 ( .A1(n5846), .A2(n7553), .ZN(n5710) );
  NAND2_X1 U7409 ( .A1(n5845), .A2(n5710), .ZN(n5712) );
  NAND2_X1 U7410 ( .A1(n5712), .A2(n5711), .ZN(n5714) );
  NAND2_X1 U7411 ( .A1(n5714), .A2(n5713), .ZN(n5715) );
  OAI21_X1 U7412 ( .B1(n5721), .B2(n5715), .A(n5828), .ZN(n5723) );
  INV_X1 U7413 ( .A(n5716), .ZN(n5719) );
  OAI21_X1 U7414 ( .B1(n5719), .B2(n5718), .A(n5717), .ZN(n5720) );
  NAND4_X1 U7415 ( .A1(n5721), .A2(n7475), .A3(n5849), .A4(n5720), .ZN(n5722)
         );
  NAND2_X1 U7416 ( .A1(n5723), .A2(n5722), .ZN(n5730) );
  AOI22_X1 U7417 ( .A1(n5726), .A2(n5848), .B1(n5725), .B2(n5724), .ZN(n5728)
         );
  INV_X1 U7418 ( .A(n5727), .ZN(n5732) );
  OAI21_X1 U7419 ( .B1(n5728), .B2(n5732), .A(n5828), .ZN(n5729) );
  MUX2_X1 U7420 ( .A(n5732), .B(n5731), .S(n5828), .Z(n5733) );
  NOR2_X1 U7421 ( .A1(n5733), .A2(n5851), .ZN(n5734) );
  MUX2_X1 U7422 ( .A(n5736), .B(n5735), .S(n5841), .Z(n5737) );
  INV_X1 U7423 ( .A(n5738), .ZN(n5741) );
  INV_X1 U7424 ( .A(n5739), .ZN(n5740) );
  MUX2_X1 U7425 ( .A(n5741), .B(n5740), .S(n5841), .Z(n5742) );
  AOI21_X1 U7426 ( .B1(n5048), .B2(n5743), .A(n5828), .ZN(n5746) );
  INV_X1 U7427 ( .A(n7684), .ZN(n5745) );
  INV_X1 U7428 ( .A(n5744), .ZN(n5751) );
  NAND2_X1 U7429 ( .A1(n7540), .A2(n5048), .ZN(n5749) );
  NAND2_X1 U7430 ( .A1(n5749), .A2(n5828), .ZN(n5755) );
  INV_X1 U7431 ( .A(n5750), .ZN(n5753) );
  AND2_X1 U7432 ( .A1(n5048), .A2(n5751), .ZN(n5752) );
  OAI21_X1 U7433 ( .B1(n5753), .B2(n5752), .A(n5841), .ZN(n5754) );
  AOI21_X1 U7434 ( .B1(n5853), .B2(n9086), .A(n5841), .ZN(n5756) );
  INV_X1 U7435 ( .A(n7700), .ZN(n9019) );
  NAND2_X1 U7436 ( .A1(n5756), .A2(n9019), .ZN(n5761) );
  INV_X1 U7437 ( .A(n9086), .ZN(n9169) );
  NAND2_X1 U7438 ( .A1(n7540), .A2(n9169), .ZN(n5757) );
  NAND3_X1 U7439 ( .A1(n7700), .A2(n5841), .A3(n5757), .ZN(n5760) );
  OR3_X1 U7440 ( .A1(n5853), .A2(n9086), .A3(n5841), .ZN(n5759) );
  OR3_X1 U7441 ( .A1(n7540), .A2(n5828), .A3(n9169), .ZN(n5758) );
  NAND4_X1 U7442 ( .A1(n5761), .A2(n5760), .A3(n5759), .A4(n5758), .ZN(n5762)
         );
  NOR2_X1 U7443 ( .A1(n7742), .A2(n5762), .ZN(n5763) );
  MUX2_X1 U7444 ( .A(n7764), .B(n5764), .S(n5841), .Z(n5765) );
  INV_X1 U7445 ( .A(n5766), .ZN(n5768) );
  MUX2_X1 U7446 ( .A(n5768), .B(n5023), .S(n5841), .Z(n5769) );
  INV_X1 U7447 ( .A(n5769), .ZN(n5771) );
  NAND2_X1 U7448 ( .A1(n4456), .A2(n5775), .ZN(n7796) );
  INV_X1 U7449 ( .A(n7796), .ZN(n5770) );
  NAND3_X1 U7450 ( .A1(n5772), .A2(n5771), .A3(n5770), .ZN(n5774) );
  NAND2_X1 U7451 ( .A1(n5774), .A2(n7831), .ZN(n5786) );
  NAND3_X1 U7452 ( .A1(n9473), .A2(n5828), .A3(n4456), .ZN(n5777) );
  NAND3_X1 U7453 ( .A1(n5779), .A2(n5775), .A3(n5841), .ZN(n5776) );
  AND2_X1 U7454 ( .A1(n5777), .A2(n5776), .ZN(n5785) );
  NAND2_X1 U7455 ( .A1(n5787), .A2(n5779), .ZN(n5778) );
  NAND2_X1 U7456 ( .A1(n5778), .A2(n5828), .ZN(n5784) );
  NAND4_X1 U7457 ( .A1(n9473), .A2(n9499), .A3(n5828), .A4(n9047), .ZN(n5781)
         );
  INV_X1 U7458 ( .A(n9047), .ZN(n9671) );
  INV_X1 U7459 ( .A(n9499), .ZN(n9165) );
  NAND4_X1 U7460 ( .A1(n5779), .A2(n9671), .A3(n9165), .A4(n5841), .ZN(n5780)
         );
  OAI211_X1 U7461 ( .C1(n5828), .C2(n9473), .A(n5781), .B(n5780), .ZN(n5782)
         );
  INV_X1 U7462 ( .A(n5782), .ZN(n5783) );
  OAI211_X1 U7463 ( .C1(n5786), .C2(n5785), .A(n5784), .B(n5783), .ZN(n5795)
         );
  NAND2_X1 U7464 ( .A1(n5795), .A2(n5787), .ZN(n5790) );
  AND2_X1 U7465 ( .A1(n5789), .A2(n5788), .ZN(n5794) );
  NAND2_X1 U7466 ( .A1(n9421), .A2(n9419), .ZN(n5792) );
  OR2_X1 U7467 ( .A1(n9414), .A2(n9107), .ZN(n5800) );
  INV_X1 U7468 ( .A(n9419), .ZN(n5793) );
  AOI21_X1 U7469 ( .B1(n5795), .B2(n5794), .A(n5793), .ZN(n5798) );
  INV_X1 U7470 ( .A(n9420), .ZN(n5797) );
  OAI211_X1 U7471 ( .C1(n5798), .C2(n5797), .A(n9421), .B(n5796), .ZN(n5799)
         );
  OAI21_X1 U7472 ( .B1(n5828), .B2(n9389), .A(n9390), .ZN(n5805) );
  INV_X1 U7473 ( .A(n5803), .ZN(n5804) );
  NAND2_X1 U7474 ( .A1(n5808), .A2(n5806), .ZN(n5807) );
  NAND2_X1 U7475 ( .A1(n5815), .A2(n5811), .ZN(n5814) );
  NAND2_X1 U7476 ( .A1(n9320), .A2(n5812), .ZN(n5813) );
  MUX2_X1 U7477 ( .A(n5814), .B(n5813), .S(n5841), .Z(n5817) );
  INV_X1 U7478 ( .A(n9315), .ZN(n9319) );
  MUX2_X1 U7479 ( .A(n9320), .B(n5815), .S(n5841), .Z(n5816) );
  INV_X1 U7480 ( .A(n5818), .ZN(n5821) );
  INV_X1 U7481 ( .A(n5819), .ZN(n5820) );
  NOR2_X1 U7482 ( .A1(n5821), .A2(n5820), .ZN(n5823) );
  MUX2_X1 U7483 ( .A(n5823), .B(n5822), .S(n5841), .Z(n5824) );
  AOI21_X1 U7484 ( .B1(n5827), .B2(n8881), .A(n5933), .ZN(n5831) );
  INV_X1 U7485 ( .A(n5832), .ZN(n5825) );
  NOR2_X1 U7486 ( .A1(n5825), .A2(n5841), .ZN(n5830) );
  OAI21_X1 U7487 ( .B1(n5831), .B2(n5830), .A(n5829), .ZN(n5837) );
  MUX2_X1 U7488 ( .A(n5833), .B(n5832), .S(n5841), .Z(n5836) );
  INV_X1 U7489 ( .A(n5834), .ZN(n5835) );
  INV_X1 U7490 ( .A(n5838), .ZN(n5859) );
  INV_X1 U7491 ( .A(n5839), .ZN(n5840) );
  NAND2_X1 U7492 ( .A1(n4444), .A2(n5840), .ZN(n5858) );
  MUX2_X1 U7493 ( .A(n5859), .B(n5858), .S(n5841), .Z(n5844) );
  MUX2_X1 U7494 ( .A(n4444), .B(n5842), .S(n5841), .Z(n5843) );
  INV_X1 U7495 ( .A(n8962), .ZN(n5863) );
  NAND2_X1 U7496 ( .A1(n9420), .A2(n9421), .ZN(n9439) );
  INV_X1 U7497 ( .A(n9461), .ZN(n5855) );
  INV_X1 U7498 ( .A(n9504), .ZN(n9496) );
  INV_X1 U7499 ( .A(n7831), .ZN(n7822) );
  INV_X1 U7500 ( .A(n7554), .ZN(n9523) );
  NOR2_X1 U7501 ( .A1(n5883), .A2(n9523), .ZN(n9527) );
  NAND4_X1 U7502 ( .A1(n9527), .A2(n5847), .A3(n5931), .A4(n7553), .ZN(n5850)
         );
  NAND4_X1 U7503 ( .A1(n5852), .A2(n7477), .A3(n5248), .A4(n7331), .ZN(n5854)
         );
  NAND2_X1 U7504 ( .A1(n5853), .A2(n7540), .ZN(n7686) );
  NAND2_X1 U7505 ( .A1(n7684), .A2(n5048), .ZN(n7669) );
  NAND4_X1 U7506 ( .A1(n9390), .A2(n5924), .A3(n5856), .A4(n9424), .ZN(n5857)
         );
  INV_X1 U7507 ( .A(n6101), .ZN(n10482) );
  OAI211_X1 U7508 ( .C1(n10482), .C2(n6037), .A(n5861), .B(n4822), .ZN(n5862)
         );
  INV_X1 U7509 ( .A(n7095), .ZN(n6767) );
  NAND2_X1 U7510 ( .A1(n5865), .A2(n5864), .ZN(n5866) );
  NAND2_X1 U7511 ( .A1(n5866), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5868) );
  NOR2_X1 U7512 ( .A1(n5870), .A2(n5869), .ZN(n5871) );
  NAND2_X1 U7513 ( .A1(n5405), .A2(n5871), .ZN(n5875) );
  OR2_X1 U7514 ( .A1(n5875), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U7515 ( .A1(n5877), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5872) );
  MUX2_X1 U7516 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5872), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5874) );
  NAND2_X1 U7517 ( .A1(n5874), .A2(n5873), .ZN(n7708) );
  NAND2_X1 U7518 ( .A1(n5875), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5876) );
  MUX2_X1 U7519 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5876), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5878) );
  NAND2_X1 U7520 ( .A1(n5878), .A2(n5877), .ZN(n7577) );
  NAND2_X1 U7521 ( .A1(n4822), .A2(n8923), .ZN(n5963) );
  NOR2_X1 U7522 ( .A1(n10467), .A2(n5963), .ZN(n6111) );
  INV_X1 U7523 ( .A(n7757), .ZN(n6804) );
  INV_X1 U7524 ( .A(n6774), .ZN(n6766) );
  NAND3_X1 U7525 ( .A1(n6111), .A2(n6804), .A3(n9462), .ZN(n5880) );
  OAI211_X1 U7526 ( .C1(n5863), .C2(n6767), .A(n5880), .B(P2_B_REG_SCAN_IN), 
        .ZN(n5881) );
  INV_X1 U7527 ( .A(n9108), .ZN(n9161) );
  NAND2_X1 U7528 ( .A1(n6829), .A2(n10488), .ZN(n5884) );
  NAND2_X1 U7529 ( .A1(n9529), .A2(n8825), .ZN(n5885) );
  NAND2_X1 U7530 ( .A1(n6822), .A2(n5885), .ZN(n6837) );
  NAND2_X1 U7531 ( .A1(n6837), .A2(n6836), .ZN(n6835) );
  NAND2_X1 U7532 ( .A1(n6946), .A2(n7415), .ZN(n5886) );
  NAND2_X1 U7533 ( .A1(n6866), .A2(n8834), .ZN(n5887) );
  NAND2_X1 U7534 ( .A1(n7088), .A2(n10496), .ZN(n5889) );
  INV_X1 U7535 ( .A(n6078), .ZN(n10508) );
  NAND2_X1 U7536 ( .A1(n10508), .A2(n7439), .ZN(n5890) );
  INV_X1 U7537 ( .A(n7717), .ZN(n9173) );
  NAND2_X1 U7538 ( .A1(n9173), .A2(n7449), .ZN(n5893) );
  INV_X1 U7539 ( .A(n7671), .ZN(n9172) );
  OR2_X1 U7540 ( .A1(n9629), .A2(n9172), .ZN(n5891) );
  NAND2_X1 U7541 ( .A1(n7665), .A2(n7669), .ZN(n5898) );
  INV_X1 U7542 ( .A(n5893), .ZN(n7711) );
  OR2_X1 U7543 ( .A1(n7716), .A2(n7711), .ZN(n7666) );
  NAND2_X1 U7544 ( .A1(n7669), .A2(n7666), .ZN(n5895) );
  OAI22_X1 U7545 ( .A1(n5895), .A2(n5894), .B1(n7730), .B2(n7785), .ZN(n5896)
         );
  INV_X1 U7546 ( .A(n5896), .ZN(n5897) );
  INV_X1 U7547 ( .A(n9014), .ZN(n9170) );
  AND2_X1 U7548 ( .A1(n9623), .A2(n9170), .ZN(n5899) );
  NAND2_X1 U7549 ( .A1(n7545), .A2(n7546), .ZN(n5902) );
  OR2_X1 U7550 ( .A1(n7700), .A2(n9169), .ZN(n5901) );
  NAND2_X1 U7551 ( .A1(n5902), .A2(n5901), .ZN(n7739) );
  INV_X1 U7552 ( .A(n8975), .ZN(n9168) );
  NAND2_X1 U7553 ( .A1(n7805), .A2(n9168), .ZN(n7760) );
  INV_X1 U7554 ( .A(n5904), .ZN(n5905) );
  OAI22_X1 U7555 ( .A1(n7742), .A2(n5905), .B1(n9167), .B2(n7772), .ZN(n5906)
         );
  INV_X1 U7556 ( .A(n5906), .ZN(n5907) );
  NAND2_X1 U7557 ( .A1(n9154), .A2(n9137), .ZN(n5908) );
  INV_X1 U7558 ( .A(n7830), .ZN(n5909) );
  NAND2_X1 U7559 ( .A1(n9047), .A2(n9165), .ZN(n5910) );
  INV_X1 U7560 ( .A(n9479), .ZN(n5911) );
  OR2_X1 U7561 ( .A1(n9512), .A2(n5911), .ZN(n9449) );
  NAND2_X1 U7562 ( .A1(n9595), .A2(n9164), .ZN(n5917) );
  INV_X1 U7563 ( .A(n5917), .ZN(n5914) );
  OR2_X1 U7564 ( .A1(n9595), .A2(n9164), .ZN(n5912) );
  INV_X1 U7565 ( .A(n9500), .ZN(n9463) );
  OR2_X1 U7566 ( .A1(n9489), .A2(n9463), .ZN(n9451) );
  AND2_X1 U7567 ( .A1(n5912), .A2(n9451), .ZN(n5913) );
  AND2_X1 U7568 ( .A1(n9449), .A2(n5916), .ZN(n5915) );
  NAND2_X1 U7569 ( .A1(n9447), .A2(n5915), .ZN(n5921) );
  INV_X1 U7570 ( .A(n5916), .ZN(n5919) );
  NAND2_X1 U7571 ( .A1(n9489), .A2(n9463), .ZN(n9450) );
  AND2_X1 U7572 ( .A1(n9450), .A2(n5917), .ZN(n5918) );
  INV_X1 U7573 ( .A(n9004), .ZN(n9465) );
  AND2_X1 U7574 ( .A1(n9433), .A2(n9465), .ZN(n5922) );
  NAND2_X1 U7575 ( .A1(n9414), .A2(n9163), .ZN(n5923) );
  NAND2_X1 U7576 ( .A1(n9374), .A2(n9373), .ZN(n9372) );
  INV_X1 U7577 ( .A(n9336), .ZN(n5927) );
  XNOR2_X1 U7578 ( .A(n5928), .B(n5933), .ZN(n9305) );
  NAND2_X1 U7579 ( .A1(n6096), .A2(n4822), .ZN(n5930) );
  AOI21_X1 U7580 ( .B1(n7318), .B2(n8962), .A(n9359), .ZN(n5929) );
  NAND2_X1 U7581 ( .A1(n5930), .A2(n5929), .ZN(n7741) );
  NOR2_X1 U7582 ( .A1(n5931), .A2(n8923), .ZN(n5932) );
  NAND2_X1 U7583 ( .A1(n5932), .A2(n8962), .ZN(n9634) );
  NAND2_X1 U7584 ( .A1(n7741), .A2(n9634), .ZN(n10510) );
  XNOR2_X1 U7585 ( .A(n5934), .B(n5933), .ZN(n5940) );
  NAND2_X1 U7586 ( .A1(n6096), .A2(n6774), .ZN(n9528) );
  INV_X1 U7587 ( .A(P2_B_REG_SCAN_IN), .ZN(n8781) );
  NOR2_X1 U7588 ( .A1(n7757), .A2(n8781), .ZN(n5936) );
  NOR2_X1 U7589 ( .A1(n9528), .A2(n5936), .ZN(n5980) );
  AOI21_X1 U7590 ( .B1(n5940), .B2(n9524), .A(n5939), .ZN(n9306) );
  NOR2_X2 U7591 ( .A1(n9539), .A2(n10481), .ZN(n9537) );
  INV_X1 U7592 ( .A(n9629), .ZN(n7725) );
  INV_X1 U7593 ( .A(n7805), .ZN(n9092) );
  INV_X1 U7594 ( .A(n7772), .ZN(n8971) );
  AND2_X2 U7595 ( .A1(n9432), .A2(n9657), .ZN(n9412) );
  INV_X1 U7596 ( .A(n5959), .ZN(n9484) );
  OAI211_X1 U7597 ( .C1(n7846), .C2(n5972), .A(n5944), .B(n9484), .ZN(n9310)
         );
  NAND2_X1 U7598 ( .A1(n9306), .A2(n9310), .ZN(n5945) );
  AOI21_X1 U7599 ( .B1(n9305), .B2(n10510), .A(n5945), .ZN(n5977) );
  INV_X1 U7600 ( .A(n7708), .ZN(n5948) );
  XOR2_X1 U7601 ( .A(n7343), .B(n8781), .Z(n5946) );
  NAND2_X1 U7602 ( .A1(n7577), .A2(n5946), .ZN(n5947) );
  INV_X1 U7603 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10475) );
  AND2_X1 U7604 ( .A1(n7343), .A2(n7708), .ZN(n10476) );
  AOI21_X1 U7605 ( .B1(n10466), .B2(n10475), .A(n10476), .ZN(n5969) );
  NOR4_X1 U7606 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n5952) );
  NOR4_X1 U7607 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5951) );
  NOR4_X1 U7608 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5950) );
  NOR4_X1 U7609 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5949) );
  NAND4_X1 U7610 ( .A1(n5952), .A2(n5951), .A3(n5950), .A4(n5949), .ZN(n5958)
         );
  NOR2_X1 U7611 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .ZN(
        n5956) );
  NOR4_X1 U7612 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5955) );
  NOR4_X1 U7613 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5954) );
  NOR4_X1 U7614 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n5953) );
  NAND4_X1 U7615 ( .A1(n5956), .A2(n5955), .A3(n5954), .A4(n5953), .ZN(n5957)
         );
  OAI21_X1 U7616 ( .B1(n5958), .B2(n5957), .A(n10466), .ZN(n5967) );
  AND2_X1 U7617 ( .A1(n5969), .A2(n5967), .ZN(n6095) );
  NOR2_X1 U7618 ( .A1(n10467), .A2(n6096), .ZN(n6770) );
  OR2_X1 U7619 ( .A1(n6111), .A2(n6770), .ZN(n5966) );
  INV_X1 U7620 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10478) );
  NAND2_X1 U7621 ( .A1(n10466), .A2(n10478), .ZN(n5961) );
  AND2_X1 U7622 ( .A1(n7708), .A2(n7577), .ZN(n10479) );
  INV_X1 U7623 ( .A(n10479), .ZN(n5960) );
  NAND2_X1 U7624 ( .A1(n5961), .A2(n5960), .ZN(n6094) );
  AND2_X1 U7625 ( .A1(n6104), .A2(n6094), .ZN(n5970) );
  AND2_X1 U7626 ( .A1(n5966), .A2(n5970), .ZN(n5962) );
  AND2_X2 U7627 ( .A1(n6095), .A2(n5962), .ZN(n10522) );
  INV_X1 U7628 ( .A(n5963), .ZN(n6106) );
  OR2_X1 U7629 ( .A1(n6106), .A2(n6101), .ZN(n10507) );
  NAND2_X1 U7630 ( .A1(n10522), .A2(n9630), .ZN(n9615) );
  NOR2_X1 U7631 ( .A1(n10522), .A2(n8765), .ZN(n5964) );
  OAI21_X1 U7632 ( .B1(n5977), .B2(n10519), .A(n5965), .ZN(P2_U3549) );
  NAND2_X1 U7633 ( .A1(n5967), .A2(n5966), .ZN(n5968) );
  INV_X1 U7634 ( .A(n5970), .ZN(n5971) );
  INV_X1 U7635 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5973) );
  OAI21_X1 U7636 ( .B1(n5977), .B2(n10512), .A(n5976), .ZN(P2_U3517) );
  NAND2_X1 U7637 ( .A1(n5979), .A2(n9484), .ZN(n9299) );
  NAND2_X1 U7638 ( .A1(n5980), .A2(n6241), .ZN(n9544) );
  NAND2_X1 U7639 ( .A1(n5983), .A2(n5037), .ZN(P2_U3551) );
  INV_X1 U7640 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U7641 ( .A1(n5986), .A2(n5041), .ZN(P2_U3519) );
  INV_X1 U7642 ( .A(n6768), .ZN(n5987) );
  BUF_X2 U7643 ( .A(n6026), .Z(n6181) );
  NAND4_X1 U7644 ( .A1(n5989), .A2(n6177), .A3(n6190), .A4(n8763), .ZN(n6027)
         );
  NOR2_X4 U7645 ( .A1(n6181), .A2(n5990), .ZN(n6012) );
  NOR2_X2 U7646 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5991) );
  NOR2_X1 U7647 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5994) );
  INV_X1 U7648 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6220) );
  INV_X1 U7649 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5993) );
  AND4_X1 U7650 ( .A1(n5994), .A2(n6220), .A3(n6004), .A4(n5993), .ZN(n5995)
         );
  AND2_X1 U7651 ( .A1(n6001), .A2(n5995), .ZN(n5996) );
  NAND2_X1 U7652 ( .A1(n6346), .A2(n6003), .ZN(n5997) );
  NAND2_X1 U7653 ( .A1(n5997), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5998) );
  OR2_X1 U7654 ( .A1(n5998), .A2(n8570), .ZN(n5999) );
  NAND2_X1 U7655 ( .A1(n8442), .A2(n8283), .ZN(n8434) );
  AND2_X1 U7656 ( .A1(n6001), .A2(n6012), .ZN(n6232) );
  NAND4_X1 U7657 ( .A1(n6491), .A2(n6003), .A3(n8570), .A4(n6002), .ZN(n6032)
         );
  NOR2_X1 U7658 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n6005) );
  INV_X1 U7659 ( .A(n6010), .ZN(n6006) );
  NAND2_X1 U7660 ( .A1(n6232), .A2(n6006), .ZN(n6007) );
  NAND2_X1 U7661 ( .A1(n6007), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6008) );
  XNOR2_X1 U7662 ( .A(n6008), .B(n6009), .ZN(n6521) );
  INV_X1 U7663 ( .A(n6521), .ZN(n7107) );
  OR2_X1 U7664 ( .A1(n8434), .A2(n7107), .ZN(n6025) );
  NOR2_X1 U7665 ( .A1(n6010), .A2(n6033), .ZN(n6011) );
  NAND2_X1 U7666 ( .A1(n6012), .A2(n6011), .ZN(n6019) );
  NAND2_X1 U7667 ( .A1(n6015), .A2(n6030), .ZN(n6017) );
  XNOR2_X2 U7668 ( .A(n6014), .B(P1_IR_REG_26__SCAN_IN), .ZN(n7704) );
  INV_X1 U7669 ( .A(n6015), .ZN(n6016) );
  NAND2_X1 U7670 ( .A1(n6016), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7671 ( .A1(n6018), .A2(n6017), .ZN(n6328) );
  NAND2_X1 U7672 ( .A1(n6019), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6020) );
  MUX2_X1 U7673 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6020), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n6022) );
  NAND2_X1 U7674 ( .A1(n6022), .A2(n6021), .ZN(n7340) );
  NOR2_X1 U7675 ( .A1(n6328), .A2(n7340), .ZN(n6023) );
  OR2_X1 U7676 ( .A1(n6024), .A2(n7107), .ZN(n6246) );
  AND2_X1 U7677 ( .A1(n6025), .A2(n6246), .ZN(n6266) );
  INV_X1 U7678 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6029) );
  NAND3_X1 U7679 ( .A1(n8553), .A2(n6030), .A3(n6029), .ZN(n6031) );
  NAND2_X1 U7680 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n6034) );
  NAND2_X1 U7681 ( .A1(n6266), .A2(n7851), .ZN(n6036) );
  NAND2_X1 U7682 ( .A1(n6036), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NOR2_X2 U7683 ( .A1(n6246), .A2(P1_U3084), .ZN(P1_U4006) );
  NAND3_X1 U7684 ( .A1(n6038), .A2(n6101), .A3(n6878), .ZN(n6039) );
  NAND2_X2 U7685 ( .A1(n6039), .A2(n7318), .ZN(n6050) );
  INV_X2 U7686 ( .A(n6050), .ZN(n8882) );
  INV_X2 U7687 ( .A(n8882), .ZN(n8868) );
  XNOR2_X1 U7688 ( .A(n6040), .B(n8868), .ZN(n6041) );
  INV_X1 U7689 ( .A(n7785), .ZN(n9171) );
  AND2_X1 U7690 ( .A1(n9171), .A2(n8835), .ZN(n6042) );
  NAND2_X1 U7691 ( .A1(n6041), .A2(n6042), .ZN(n6122) );
  INV_X1 U7692 ( .A(n6041), .ZN(n7782) );
  INV_X1 U7693 ( .A(n6042), .ZN(n6043) );
  NAND2_X1 U7694 ( .A1(n7782), .A2(n6043), .ZN(n6044) );
  NAND2_X1 U7695 ( .A1(n6122), .A2(n6044), .ZN(n6100) );
  XNOR2_X1 U7696 ( .A(n6050), .B(n10488), .ZN(n6047) );
  NAND2_X1 U7697 ( .A1(n6045), .A2(n8835), .ZN(n6046) );
  NAND2_X1 U7698 ( .A1(n6047), .A2(n6046), .ZN(n6049) );
  NAND2_X1 U7699 ( .A1(n6976), .A2(n8835), .ZN(n7014) );
  XNOR2_X1 U7700 ( .A(n6050), .B(n8825), .ZN(n6052) );
  NAND2_X1 U7701 ( .A1(n6051), .A2(n8835), .ZN(n6053) );
  NAND2_X1 U7702 ( .A1(n6052), .A2(n6053), .ZN(n6057) );
  INV_X1 U7703 ( .A(n6052), .ZN(n6055) );
  INV_X1 U7704 ( .A(n6053), .ZN(n6054) );
  NAND2_X1 U7705 ( .A1(n6055), .A2(n6054), .ZN(n6056) );
  AND2_X1 U7706 ( .A1(n6057), .A2(n6056), .ZN(n8818) );
  NAND2_X1 U7707 ( .A1(n8816), .A2(n6057), .ZN(n6872) );
  XNOR2_X1 U7708 ( .A(n6050), .B(n7415), .ZN(n6058) );
  NAND2_X1 U7709 ( .A1(n9177), .A2(n8835), .ZN(n6059) );
  XNOR2_X1 U7710 ( .A(n6058), .B(n6059), .ZN(n6871) );
  INV_X1 U7711 ( .A(n6058), .ZN(n6061) );
  INV_X1 U7712 ( .A(n6059), .ZN(n6060) );
  NAND2_X1 U7713 ( .A1(n6061), .A2(n6060), .ZN(n6062) );
  XNOR2_X1 U7714 ( .A(n8868), .B(n5104), .ZN(n6063) );
  AND2_X1 U7715 ( .A1(n9176), .A2(n8835), .ZN(n6064) );
  AND2_X1 U7716 ( .A1(n6063), .A2(n6064), .ZN(n6943) );
  INV_X1 U7717 ( .A(n6063), .ZN(n6066) );
  INV_X1 U7718 ( .A(n6064), .ZN(n6065) );
  NAND2_X1 U7719 ( .A1(n6066), .A2(n6065), .ZN(n6942) );
  OAI21_X1 U7720 ( .B1(n6941), .B2(n6943), .A(n6942), .ZN(n6865) );
  XNOR2_X1 U7721 ( .A(n8872), .B(n10496), .ZN(n6067) );
  AND2_X1 U7722 ( .A1(n6067), .A2(n6068), .ZN(n6861) );
  INV_X1 U7723 ( .A(n6067), .ZN(n6070) );
  INV_X1 U7724 ( .A(n6068), .ZN(n6069) );
  NAND2_X1 U7725 ( .A1(n6070), .A2(n6069), .ZN(n6862) );
  XNOR2_X1 U7726 ( .A(n10501), .B(n8868), .ZN(n6072) );
  NAND2_X1 U7727 ( .A1(n9175), .A2(n8835), .ZN(n6073) );
  NAND2_X1 U7728 ( .A1(n6072), .A2(n6073), .ZN(n6077) );
  INV_X1 U7729 ( .A(n6072), .ZN(n6075) );
  INV_X1 U7730 ( .A(n6073), .ZN(n6074) );
  NAND2_X1 U7731 ( .A1(n6075), .A2(n6074), .ZN(n6076) );
  AND2_X1 U7732 ( .A1(n6077), .A2(n6076), .ZN(n7087) );
  XNOR2_X1 U7733 ( .A(n8872), .B(n6078), .ZN(n6079) );
  INV_X1 U7734 ( .A(n7439), .ZN(n9174) );
  AND2_X1 U7735 ( .A1(n9174), .A2(n8835), .ZN(n6080) );
  XNOR2_X1 U7736 ( .A(n6079), .B(n6080), .ZN(n7098) );
  INV_X1 U7737 ( .A(n6079), .ZN(n6082) );
  INV_X1 U7738 ( .A(n6080), .ZN(n6081) );
  XNOR2_X1 U7739 ( .A(n8868), .B(n7449), .ZN(n6085) );
  NAND2_X1 U7740 ( .A1(n9173), .A2(n8835), .ZN(n6083) );
  XNOR2_X1 U7741 ( .A(n6085), .B(n6083), .ZN(n7275) );
  NAND2_X1 U7742 ( .A1(n7276), .A2(n7275), .ZN(n6087) );
  INV_X1 U7743 ( .A(n6083), .ZN(n6084) );
  NAND2_X1 U7744 ( .A1(n6085), .A2(n6084), .ZN(n6086) );
  NAND2_X1 U7745 ( .A1(n6087), .A2(n6086), .ZN(n7518) );
  INV_X1 U7746 ( .A(n7518), .ZN(n6089) );
  XNOR2_X1 U7747 ( .A(n9629), .B(n8872), .ZN(n6090) );
  AND2_X1 U7748 ( .A1(n9172), .A2(n8835), .ZN(n6091) );
  AND2_X1 U7749 ( .A1(n6090), .A2(n6091), .ZN(n7515) );
  INV_X1 U7750 ( .A(n7515), .ZN(n6088) );
  INV_X1 U7751 ( .A(n6090), .ZN(n6093) );
  INV_X1 U7752 ( .A(n6091), .ZN(n6092) );
  NAND2_X1 U7753 ( .A1(n6093), .A2(n6092), .ZN(n7514) );
  INV_X1 U7754 ( .A(n6094), .ZN(n7312) );
  NAND2_X1 U7755 ( .A1(n6095), .A2(n7312), .ZN(n6110) );
  NOR2_X1 U7756 ( .A1(n6110), .A2(n10467), .ZN(n6102) );
  INV_X1 U7757 ( .A(n6096), .ZN(n6237) );
  AND2_X1 U7758 ( .A1(n6237), .A2(n10507), .ZN(n6097) );
  INV_X1 U7759 ( .A(n7781), .ZN(n6098) );
  AOI211_X1 U7760 ( .C1(n6100), .C2(n6099), .A(n9138), .B(n6098), .ZN(n6116)
         );
  NOR2_X1 U7761 ( .A1(n6101), .A2(n4822), .ZN(n7321) );
  NAND2_X1 U7762 ( .A1(n6102), .A2(n7321), .ZN(n6103) );
  NOR2_X1 U7763 ( .A1(n9153), .A2(n7730), .ZN(n6115) );
  NAND2_X1 U7764 ( .A1(n6110), .A2(n6104), .ZN(n6109) );
  OAI211_X1 U7765 ( .C1(n6106), .C2(n6237), .A(n6768), .B(n6105), .ZN(n6107)
         );
  INV_X1 U7766 ( .A(n6107), .ZN(n6108) );
  NAND2_X1 U7767 ( .A1(n6109), .A2(n6108), .ZN(n6975) );
  INV_X1 U7768 ( .A(n6110), .ZN(n6112) );
  NAND2_X1 U7769 ( .A1(n6112), .A2(n6111), .ZN(n9073) );
  OAI22_X1 U7770 ( .A1(n9131), .A2(n7677), .B1(n7671), .B2(n9145), .ZN(n6114)
         );
  OAI22_X1 U7771 ( .A1(n9148), .A2(n9014), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8720), .ZN(n6113) );
  OR4_X1 U7772 ( .A1(n6116), .A2(n6115), .A3(n6114), .A4(n6113), .ZN(P2_U3219)
         );
  XNOR2_X1 U7773 ( .A(n9595), .B(n8872), .ZN(n6120) );
  INV_X1 U7774 ( .A(n6120), .ZN(n6118) );
  NOR2_X1 U7775 ( .A1(n9480), .A2(n8880), .ZN(n6119) );
  INV_X1 U7776 ( .A(n6119), .ZN(n6117) );
  NAND2_X1 U7777 ( .A1(n6118), .A2(n6117), .ZN(n9069) );
  INV_X1 U7778 ( .A(n9069), .ZN(n8838) );
  AND2_X1 U7779 ( .A1(n6120), .A2(n6119), .ZN(n8841) );
  NOR3_X1 U7780 ( .A1(n8838), .A2(n8841), .A3(n9138), .ZN(n6161) );
  OR2_X1 U7781 ( .A1(n9138), .A2(n8880), .ZN(n9136) );
  INV_X1 U7782 ( .A(n9136), .ZN(n9102) );
  NAND3_X1 U7783 ( .A1(n6120), .A2(n9102), .A3(n9164), .ZN(n6121) );
  OAI21_X1 U7784 ( .B1(n9069), .B2(n9138), .A(n6121), .ZN(n6160) );
  XNOR2_X1 U7785 ( .A(n9623), .B(n8872), .ZN(n6123) );
  AND2_X1 U7786 ( .A1(n9170), .A2(n8835), .ZN(n6124) );
  NAND2_X1 U7787 ( .A1(n6123), .A2(n6124), .ZN(n6128) );
  INV_X1 U7788 ( .A(n6123), .ZN(n9013) );
  INV_X1 U7789 ( .A(n6124), .ZN(n6125) );
  NAND2_X1 U7790 ( .A1(n9013), .A2(n6125), .ZN(n6126) );
  NAND2_X1 U7791 ( .A1(n6127), .A2(n7779), .ZN(n9012) );
  NAND2_X1 U7792 ( .A1(n9012), .A2(n6128), .ZN(n6133) );
  XNOR2_X1 U7793 ( .A(n7700), .B(n8868), .ZN(n6129) );
  AND2_X1 U7794 ( .A1(n9169), .A2(n8835), .ZN(n6130) );
  NAND2_X1 U7795 ( .A1(n6129), .A2(n6130), .ZN(n6134) );
  INV_X1 U7796 ( .A(n6129), .ZN(n9080) );
  INV_X1 U7797 ( .A(n6130), .ZN(n6131) );
  NAND2_X1 U7798 ( .A1(n9080), .A2(n6131), .ZN(n6132) );
  NAND2_X1 U7799 ( .A1(n6133), .A2(n9010), .ZN(n9015) );
  NAND2_X1 U7800 ( .A1(n9015), .A2(n6134), .ZN(n6139) );
  XNOR2_X1 U7801 ( .A(n7805), .B(n8868), .ZN(n6135) );
  AND2_X1 U7802 ( .A1(n9168), .A2(n8835), .ZN(n6136) );
  NAND2_X1 U7803 ( .A1(n6135), .A2(n6136), .ZN(n6140) );
  INV_X1 U7804 ( .A(n6135), .ZN(n8967) );
  INV_X1 U7805 ( .A(n6136), .ZN(n6137) );
  NAND2_X1 U7806 ( .A1(n8967), .A2(n6137), .ZN(n6138) );
  AND2_X1 U7807 ( .A1(n6140), .A2(n6138), .ZN(n9078) );
  NAND2_X1 U7808 ( .A1(n6139), .A2(n9078), .ZN(n8966) );
  XNOR2_X1 U7809 ( .A(n7772), .B(n8872), .ZN(n6142) );
  NAND2_X1 U7810 ( .A1(n8835), .A2(n9167), .ZN(n6143) );
  XNOR2_X1 U7811 ( .A(n6142), .B(n6143), .ZN(n8981) );
  AND2_X1 U7812 ( .A1(n8981), .A2(n6140), .ZN(n6141) );
  NAND2_X1 U7813 ( .A1(n8966), .A2(n6141), .ZN(n8970) );
  INV_X1 U7814 ( .A(n6142), .ZN(n6144) );
  NAND2_X1 U7815 ( .A1(n6144), .A2(n6143), .ZN(n6145) );
  XNOR2_X1 U7816 ( .A(n9047), .B(n8872), .ZN(n9040) );
  NOR2_X1 U7817 ( .A1(n9499), .A2(n8880), .ZN(n6146) );
  AND2_X1 U7818 ( .A1(n8835), .A2(n9166), .ZN(n9036) );
  XNOR2_X1 U7819 ( .A(n9154), .B(n8882), .ZN(n9035) );
  OAI22_X1 U7820 ( .A1(n9040), .A2(n6146), .B1(n9036), .B2(n9035), .ZN(n6151)
         );
  INV_X1 U7821 ( .A(n9035), .ZN(n9038) );
  INV_X1 U7822 ( .A(n9036), .ZN(n6147) );
  INV_X1 U7823 ( .A(n6146), .ZN(n9039) );
  OAI21_X1 U7824 ( .B1(n9038), .B2(n6147), .A(n9039), .ZN(n6149) );
  NOR2_X1 U7825 ( .A1(n9039), .A2(n6147), .ZN(n6148) );
  AOI22_X1 U7826 ( .A1(n6149), .A2(n9040), .B1(n6148), .B2(n9035), .ZN(n6150)
         );
  XNOR2_X1 U7827 ( .A(n9512), .B(n8872), .ZN(n6152) );
  NOR2_X1 U7828 ( .A1(n9479), .A2(n8880), .ZN(n6153) );
  NAND2_X1 U7829 ( .A1(n6152), .A2(n6153), .ZN(n8852) );
  INV_X1 U7830 ( .A(n6152), .ZN(n9116) );
  INV_X1 U7831 ( .A(n6153), .ZN(n6154) );
  NAND2_X1 U7832 ( .A1(n9116), .A2(n6154), .ZN(n6155) );
  AND2_X1 U7833 ( .A1(n8852), .A2(n6155), .ZN(n9051) );
  NAND2_X1 U7834 ( .A1(n8858), .A2(n8852), .ZN(n9094) );
  XNOR2_X1 U7835 ( .A(n9489), .B(n8872), .ZN(n6158) );
  NAND2_X1 U7836 ( .A1(n9463), .A2(n8835), .ZN(n6156) );
  XNOR2_X1 U7837 ( .A(n6158), .B(n6156), .ZN(n9114) );
  NAND2_X1 U7838 ( .A1(n9094), .A2(n9114), .ZN(n9117) );
  INV_X1 U7839 ( .A(n6156), .ZN(n6157) );
  NAND2_X1 U7840 ( .A1(n6158), .A2(n6157), .ZN(n8839) );
  NAND2_X1 U7841 ( .A1(n9117), .A2(n8839), .ZN(n6159) );
  MUX2_X1 U7842 ( .A(n6161), .B(n6160), .S(n6159), .Z(n6168) );
  INV_X1 U7843 ( .A(n9595), .ZN(n6162) );
  NOR2_X1 U7844 ( .A1(n6162), .A2(n9153), .ZN(n6167) );
  OAI22_X1 U7845 ( .A1(n9145), .A2(n9500), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6163), .ZN(n6166) );
  INV_X1 U7846 ( .A(n6164), .ZN(n9458) );
  OAI22_X1 U7847 ( .A1(n9131), .A2(n9458), .B1(n9004), .B2(n9148), .ZN(n6165)
         );
  INV_X1 U7848 ( .A(n6961), .ZN(n6170) );
  NAND2_X1 U7849 ( .A1(n5133), .A2(P2_U3152), .ZN(n8964) );
  INV_X1 U7850 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6169) );
  NOR2_X1 U7851 ( .A1(n5133), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9680) );
  INV_X1 U7852 ( .A(n9680), .ZN(n9686) );
  OAI222_X1 U7853 ( .A1(n6170), .A2(P2_U3152), .B1(n8964), .B2(n6399), .C1(
        n6169), .C2(n9686), .ZN(P2_U3357) );
  AND2_X1 U7854 ( .A1(n5133), .A2(P1_U3084), .ZN(n10340) );
  INV_X1 U7855 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6556) );
  AND2_X1 U7856 ( .A1(n6398), .A2(P1_U3084), .ZN(n7106) );
  INV_X2 U7857 ( .A(n7106), .ZN(n10347) );
  INV_X1 U7858 ( .A(n6555), .ZN(n6186) );
  NAND2_X1 U7859 ( .A1(n6171), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6172) );
  MUX2_X1 U7860 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6172), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n6173) );
  NAND2_X1 U7861 ( .A1(n6173), .A2(n6181), .ZN(n10392) );
  OAI222_X1 U7862 ( .A1(n10350), .A2(n6556), .B1(n10347), .B2(n6186), .C1(
        P1_U3084), .C2(n10392), .ZN(P1_U3349) );
  XNOR2_X1 U7863 ( .A(n6278), .B(n8548), .ZN(n6649) );
  OAI222_X1 U7864 ( .A1(n6649), .A2(P1_U3084), .B1(n10347), .B2(n6418), .C1(
        n6417), .C2(n10350), .ZN(P1_U3351) );
  CLKBUF_X1 U7865 ( .A(n8964), .Z(n9684) );
  AOI22_X1 U7866 ( .A1(n9179), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n9680), .ZN(n6175) );
  OAI21_X1 U7867 ( .B1(n8175), .B2(n9684), .A(n6175), .ZN(P2_U3355) );
  INV_X1 U7868 ( .A(n6885), .ZN(n6180) );
  AOI22_X1 U7869 ( .A1(n9210), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n9680), .ZN(n6176) );
  OAI21_X1 U7870 ( .B1(n6180), .B2(n9684), .A(n6176), .ZN(P2_U3351) );
  NOR2_X1 U7871 ( .A1(n6181), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n6197) );
  NAND2_X1 U7872 ( .A1(n6197), .A2(n6177), .ZN(n6189) );
  NAND2_X1 U7873 ( .A1(n6189), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6178) );
  XNOR2_X1 U7874 ( .A(n6178), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10409) );
  AOI22_X1 U7875 ( .A1(n10409), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10340), .ZN(n6179) );
  OAI21_X1 U7876 ( .B1(n6180), .B2(n10347), .A(n6179), .ZN(P1_U3346) );
  INV_X1 U7877 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n8576) );
  INV_X1 U7878 ( .A(n6624), .ZN(n6184) );
  NAND2_X1 U7879 ( .A1(n6181), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6182) );
  XNOR2_X1 U7880 ( .A(n6182), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6623) );
  INV_X1 U7881 ( .A(n6623), .ZN(n6317) );
  OAI222_X1 U7882 ( .A1(n10350), .A2(n8576), .B1(n10347), .B2(n6184), .C1(
        P1_U3084), .C2(n6317), .ZN(P1_U3348) );
  INV_X1 U7883 ( .A(n7083), .ZN(n6755) );
  OAI222_X1 U7884 ( .A1(n6755), .A2(P2_U3152), .B1(n9684), .B2(n6418), .C1(
        n6183), .C2(n9686), .ZN(P2_U3356) );
  INV_X1 U7885 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6185) );
  OAI222_X1 U7886 ( .A1(n9686), .A2(n6185), .B1(n9684), .B2(n6184), .C1(
        P2_U3152), .C2(n9197), .ZN(P2_U3353) );
  INV_X1 U7887 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6187) );
  OAI222_X1 U7888 ( .A1(n9686), .A2(n6187), .B1(n9684), .B2(n6186), .C1(
        P2_U3152), .C2(n8530), .ZN(P2_U3354) );
  INV_X1 U7889 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n8546) );
  INV_X1 U7890 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6397) );
  INV_X1 U7891 ( .A(n7041), .ZN(n6195) );
  NAND2_X1 U7892 ( .A1(n6192), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6191) );
  MUX2_X1 U7893 ( .A(n6191), .B(P1_IR_REG_31__SCAN_IN), .S(n6190), .Z(n6193)
         );
  INV_X1 U7894 ( .A(n7042), .ZN(n6541) );
  OAI222_X1 U7895 ( .A1(n10350), .A2(n6194), .B1(n10347), .B2(n6195), .C1(
        P1_U3084), .C2(n6541), .ZN(P1_U3345) );
  INV_X1 U7896 ( .A(n9223), .ZN(n6763) );
  OAI222_X1 U7897 ( .A1(n9686), .A2(n6196), .B1(n8964), .B2(n6195), .C1(
        P2_U3152), .C2(n6763), .ZN(P2_U3350) );
  INV_X1 U7898 ( .A(n6696), .ZN(n6200) );
  INV_X1 U7899 ( .A(n6919), .ZN(n6760) );
  OAI222_X1 U7900 ( .A1(n9686), .A2(n4509), .B1(n9684), .B2(n6200), .C1(
        P2_U3152), .C2(n6760), .ZN(P2_U3352) );
  INV_X1 U7901 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n8756) );
  OR2_X1 U7902 ( .A1(n6197), .A2(n6218), .ZN(n6198) );
  INV_X1 U7903 ( .A(n6697), .ZN(n6199) );
  OAI222_X1 U7904 ( .A1(n10350), .A2(n8756), .B1(n10347), .B2(n6200), .C1(
        P1_U3084), .C2(n6199), .ZN(P1_U3347) );
  INV_X1 U7905 ( .A(n7137), .ZN(n6207) );
  AOI22_X1 U7906 ( .A1(n9247), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n9680), .ZN(n6201) );
  OAI21_X1 U7907 ( .B1(n6207), .B2(n9684), .A(n6201), .ZN(P2_U3349) );
  NAND2_X1 U7908 ( .A1(n6202), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6203) );
  MUX2_X1 U7909 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6203), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n6204) );
  INV_X1 U7910 ( .A(n6204), .ZN(n6205) );
  AOI22_X1 U7911 ( .A1(n7138), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n10340), .ZN(n6206) );
  OAI21_X1 U7912 ( .B1(n6207), .B2(n10347), .A(n6206), .ZN(P1_U3344) );
  INV_X1 U7913 ( .A(n7249), .ZN(n6216) );
  AOI22_X1 U7914 ( .A1(n9262), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n9680), .ZN(n6208) );
  OAI21_X1 U7915 ( .B1(n6216), .B2(n9684), .A(n6208), .ZN(P2_U3347) );
  INV_X1 U7916 ( .A(n7203), .ZN(n6213) );
  NOR2_X1 U7917 ( .A1(n6012), .A2(n6218), .ZN(n6209) );
  MUX2_X1 U7918 ( .A(n6218), .B(n6209), .S(P1_IR_REG_10__SCAN_IN), .Z(n6211)
         );
  INV_X1 U7919 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n8554) );
  NAND2_X1 U7920 ( .A1(n6012), .A2(n8554), .ZN(n6225) );
  INV_X1 U7921 ( .A(n6225), .ZN(n6210) );
  OR2_X1 U7922 ( .A1(n6211), .A2(n6210), .ZN(n6729) );
  OAI222_X1 U7923 ( .A1(n10350), .A2(n6212), .B1(n10347), .B2(n6213), .C1(
        n6729), .C2(P1_U3084), .ZN(P1_U3343) );
  INV_X1 U7924 ( .A(n6796), .ZN(n6851) );
  OAI222_X1 U7925 ( .A1(n9686), .A2(n6214), .B1(n8964), .B2(n6213), .C1(n6851), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U7926 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7927 ( .A1(n6225), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6215) );
  XNOR2_X1 U7928 ( .A(n6215), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7250) );
  INV_X1 U7929 ( .A(n7250), .ZN(n6734) );
  OAI222_X1 U7930 ( .A1(n10350), .A2(n6217), .B1(n10347), .B2(n6216), .C1(
        n6734), .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U7931 ( .A(n7855), .ZN(n6223) );
  NOR2_X1 U7932 ( .A1(n6232), .A2(n6218), .ZN(n6219) );
  MUX2_X1 U7933 ( .A(n6218), .B(n6219), .S(P1_IR_REG_14__SCAN_IN), .Z(n6222)
         );
  NAND2_X1 U7934 ( .A1(n6232), .A2(n6220), .ZN(n6262) );
  INV_X1 U7935 ( .A(n6262), .ZN(n6221) );
  OR2_X1 U7936 ( .A1(n6222), .A2(n6221), .ZN(n9884) );
  OAI222_X1 U7937 ( .A1(n10350), .A2(n8787), .B1(n10347), .B2(n6223), .C1(
        n9884), .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U7938 ( .A(n6992), .ZN(n7188) );
  OAI222_X1 U7939 ( .A1(n9686), .A2(n6224), .B1(n8964), .B2(n6223), .C1(n7188), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U7940 ( .A(n7488), .ZN(n6228) );
  OR2_X1 U7941 ( .A1(n6225), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n6230) );
  NAND2_X1 U7942 ( .A1(n6230), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6226) );
  XNOR2_X1 U7943 ( .A(n6226), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7489) );
  INV_X1 U7944 ( .A(n7489), .ZN(n7114) );
  OAI222_X1 U7945 ( .A1(n10350), .A2(n6227), .B1(n10347), .B2(n6228), .C1(
        P1_U3084), .C2(n7114), .ZN(P1_U3341) );
  INV_X1 U7946 ( .A(n6800), .ZN(n7030) );
  OAI222_X1 U7947 ( .A1(n9686), .A2(n6229), .B1(n8964), .B2(n6228), .C1(
        P2_U3152), .C2(n7030), .ZN(P2_U3346) );
  INV_X1 U7948 ( .A(n7617), .ZN(n6235) );
  OAI21_X1 U7949 ( .B1(n6230), .B2(P1_IR_REG_12__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6231) );
  MUX2_X1 U7950 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6231), .S(
        P1_IR_REG_13__SCAN_IN), .Z(n6234) );
  INV_X1 U7951 ( .A(n6232), .ZN(n6233) );
  INV_X1 U7952 ( .A(n9864), .ZN(n7425) );
  OAI222_X1 U7953 ( .A1(n10350), .A2(n8776), .B1(n10347), .B2(n6235), .C1(
        n7425), .C2(P1_U3084), .ZN(P1_U3340) );
  INV_X1 U7954 ( .A(n6983), .ZN(n6777) );
  OAI222_X1 U7955 ( .A1(n9686), .A2(n6236), .B1(n8964), .B2(n6235), .C1(n6777), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  OAI21_X1 U7956 ( .B1(n10467), .B2(n6237), .A(n6771), .ZN(n6239) );
  NAND2_X1 U7957 ( .A1(n10467), .A2(n6767), .ZN(n6238) );
  NAND2_X1 U7958 ( .A1(n6239), .A2(n6238), .ZN(n8927) );
  NOR2_X1 U7959 ( .A1(n9289), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7960 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8705) );
  NAND2_X1 U7961 ( .A1(n6976), .A2(P2_U3966), .ZN(n6240) );
  OAI21_X1 U7962 ( .B1(n8705), .B2(P2_U3966), .A(n6240), .ZN(P2_U3552) );
  NAND2_X1 U7963 ( .A1(n6241), .A2(P2_U3966), .ZN(n6242) );
  OAI21_X1 U7964 ( .B1(n5684), .B2(P2_U3966), .A(n6242), .ZN(P2_U3583) );
  INV_X1 U7965 ( .A(n7858), .ZN(n6244) );
  INV_X1 U7966 ( .A(n7597), .ZN(n7183) );
  OAI222_X1 U7967 ( .A1(n9686), .A2(n8635), .B1(n8964), .B2(n6244), .C1(
        P2_U3152), .C2(n7183), .ZN(P2_U3343) );
  NAND2_X1 U7968 ( .A1(n6262), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6243) );
  XNOR2_X1 U7969 ( .A(n6243), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9888) );
  OAI222_X1 U7970 ( .A1(n10350), .A2(n6245), .B1(n10347), .B2(n6244), .C1(
        P1_U3084), .C2(n9889), .ZN(P1_U3338) );
  INV_X1 U7971 ( .A(n6246), .ZN(n6247) );
  OR2_X1 U7972 ( .A1(P1_U3083), .A2(n6247), .ZN(n10431) );
  INV_X1 U7973 ( .A(n10431), .ZN(n10410) );
  INV_X1 U7974 ( .A(n6266), .ZN(n6255) );
  NOR2_X1 U7975 ( .A1(n7916), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6250) );
  OR2_X1 U7976 ( .A1(n6250), .A2(n8929), .ZN(n6251) );
  INV_X1 U7977 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6374) );
  OR2_X1 U7978 ( .A1(n6251), .A2(n6374), .ZN(n6656) );
  NAND2_X1 U7979 ( .A1(n6251), .A2(n6374), .ZN(n6658) );
  INV_X1 U7980 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6380) );
  OAI21_X1 U7981 ( .B1(n8929), .B2(n6380), .A(n7916), .ZN(n6252) );
  NAND4_X1 U7982 ( .A1(n6656), .A2(P1_STATE_REG_SCAN_IN), .A3(n6658), .A4(
        n6252), .ZN(n6254) );
  INV_X1 U7983 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6253) );
  OAI22_X1 U7984 ( .A1(n6255), .A2(n6254), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6253), .ZN(n6259) );
  NAND2_X1 U7985 ( .A1(n7916), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6256) );
  NOR2_X1 U7986 ( .A1(n8929), .A2(n6256), .ZN(n6257) );
  INV_X1 U7987 ( .A(n10427), .ZN(n10394) );
  NOR3_X1 U7988 ( .A1(n10394), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n6374), .ZN(
        n6258) );
  AOI211_X1 U7989 ( .C1(P1_ADDR_REG_0__SCAN_IN), .C2(n10410), .A(n6259), .B(
        n6258), .ZN(n6260) );
  INV_X1 U7990 ( .A(n6260), .ZN(P1_U3241) );
  MUX2_X1 U7991 ( .A(n6495), .B(n9479), .S(P2_U3966), .Z(n6261) );
  INV_X1 U7992 ( .A(n6261), .ZN(P2_U3569) );
  INV_X1 U7993 ( .A(n7864), .ZN(n6264) );
  INV_X1 U7994 ( .A(n8902), .ZN(n8911) );
  OAI222_X1 U7995 ( .A1(n9686), .A2(n8782), .B1(n8964), .B2(n6264), .C1(n8911), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  OR2_X1 U7996 ( .A1(n6262), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n6488) );
  NAND2_X1 U7997 ( .A1(n6488), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6263) );
  XNOR2_X1 U7998 ( .A(n6263), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9917) );
  INV_X1 U7999 ( .A(n9917), .ZN(n9908) );
  OAI222_X1 U8000 ( .A1(n10350), .A2(n6265), .B1(n10347), .B2(n6264), .C1(
        n9908), .C2(P1_U3084), .ZN(P1_U3337) );
  INV_X1 U8001 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6277) );
  NOR2_X1 U8002 ( .A1(n7916), .A2(P1_U3084), .ZN(n7709) );
  NAND2_X1 U8003 ( .A1(n6266), .A2(n7709), .ZN(n9948) );
  INV_X1 U8004 ( .A(n10416), .ZN(n9946) );
  AND2_X1 U8005 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6294) );
  XOR2_X1 U8006 ( .A(n6295), .B(n6294), .Z(n6275) );
  INV_X1 U8007 ( .A(n8929), .ZN(n6451) );
  OR2_X1 U8008 ( .A1(n9948), .A2(n6451), .ZN(n10393) );
  NAND2_X1 U8009 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(P1_U3084), .ZN(n6273) );
  INV_X1 U8010 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n8682) );
  AND2_X1 U8011 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6268) );
  NAND2_X1 U8012 ( .A1(n6267), .A2(n6268), .ZN(n6284) );
  INV_X1 U8013 ( .A(n6268), .ZN(n6269) );
  NAND2_X1 U8014 ( .A1(n6270), .A2(n6269), .ZN(n6271) );
  NAND3_X1 U8015 ( .A1(n10427), .A2(n6284), .A3(n6271), .ZN(n6272) );
  AOI21_X1 U8016 ( .B1(n9946), .B2(n6275), .A(n6274), .ZN(n6276) );
  OAI21_X1 U8017 ( .B1(n10431), .B2(n6277), .A(n6276), .ZN(P1_U3242) );
  INV_X1 U8018 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6305) );
  NAND2_X1 U8019 ( .A1(n6278), .A2(n8548), .ZN(n6279) );
  NAND2_X1 U8020 ( .A1(n6279), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6281) );
  INV_X1 U8021 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n6280) );
  XNOR2_X1 U8022 ( .A(n6281), .B(n6280), .ZN(n6293) );
  NAND2_X1 U8023 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6526) );
  INV_X1 U8024 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6282) );
  MUX2_X1 U8025 ( .A(n6282), .B(P1_REG1_REG_2__SCAN_IN), .S(n6649), .Z(n6285)
         );
  NAND2_X1 U8026 ( .A1(n6284), .A2(n6283), .ZN(n6648) );
  NAND2_X1 U8027 ( .A1(n6285), .A2(n6648), .ZN(n6650) );
  INV_X1 U8028 ( .A(n6649), .ZN(n6655) );
  NAND2_X1 U8029 ( .A1(n6655), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U8030 ( .A1(n6650), .A2(n6288), .ZN(n6287) );
  INV_X1 U8031 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6428) );
  MUX2_X1 U8032 ( .A(n6428), .B(P1_REG1_REG_3__SCAN_IN), .S(n4373), .Z(n6286)
         );
  NAND2_X1 U8033 ( .A1(n6287), .A2(n6286), .ZN(n6307) );
  MUX2_X1 U8034 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6428), .S(n4373), .Z(n6289)
         );
  NAND3_X1 U8035 ( .A1(n6289), .A2(n6650), .A3(n6288), .ZN(n6290) );
  NAND3_X1 U8036 ( .A1(n10427), .A2(n6307), .A3(n6290), .ZN(n6291) );
  OAI211_X1 U8037 ( .C1(n10393), .C2(n4373), .A(n6526), .B(n6291), .ZN(n6292)
         );
  INV_X1 U8038 ( .A(n6292), .ZN(n6304) );
  INV_X1 U8039 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6430) );
  MUX2_X1 U8040 ( .A(n6430), .B(P1_REG2_REG_3__SCAN_IN), .S(n4373), .Z(n6302)
         );
  NAND2_X1 U8041 ( .A1(n6295), .A2(n6294), .ZN(n6298) );
  NAND2_X1 U8042 ( .A1(n6296), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6297) );
  NAND2_X1 U8043 ( .A1(n6298), .A2(n6297), .ZN(n6662) );
  XNOR2_X1 U8044 ( .A(n6649), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6663) );
  NAND2_X1 U8045 ( .A1(n6662), .A2(n6663), .ZN(n6300) );
  NAND2_X1 U8046 ( .A1(n6655), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6299) );
  NAND2_X1 U8047 ( .A1(n6300), .A2(n6299), .ZN(n6301) );
  OAI211_X1 U8048 ( .C1(n6302), .C2(n6301), .A(n9946), .B(n6321), .ZN(n6303)
         );
  OAI211_X1 U8049 ( .C1(n6305), .C2(n10431), .A(n6304), .B(n6303), .ZN(
        P1_U3244) );
  INV_X1 U8050 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6327) );
  NAND2_X1 U8051 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3084), .ZN(n6642) );
  INV_X1 U8052 ( .A(n4373), .ZN(n6319) );
  NAND2_X1 U8053 ( .A1(n6319), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U8054 ( .A1(n6307), .A2(n6306), .ZN(n10390) );
  INV_X1 U8055 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6308) );
  MUX2_X1 U8056 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6308), .S(n10392), .Z(n10391) );
  NOR2_X1 U8057 ( .A1(n10390), .A2(n10391), .ZN(n10389) );
  AND2_X1 U8058 ( .A1(n10392), .A2(n6308), .ZN(n6309) );
  INV_X1 U8059 ( .A(n6314), .ZN(n6312) );
  INV_X1 U8060 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6310) );
  MUX2_X1 U8061 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6310), .S(n6623), .Z(n6311)
         );
  NAND2_X1 U8062 ( .A1(n6312), .A2(n6311), .ZN(n6473) );
  MUX2_X1 U8063 ( .A(n6310), .B(P1_REG1_REG_5__SCAN_IN), .S(n6623), .Z(n6313)
         );
  NAND2_X1 U8064 ( .A1(n6314), .A2(n6313), .ZN(n6315) );
  NAND3_X1 U8065 ( .A1(n10427), .A2(n6473), .A3(n6315), .ZN(n6316) );
  OAI211_X1 U8066 ( .C1(n10393), .C2(n6317), .A(n6642), .B(n6316), .ZN(n6318)
         );
  INV_X1 U8067 ( .A(n6318), .ZN(n6326) );
  NAND2_X1 U8068 ( .A1(n6319), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6320) );
  INV_X1 U8069 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7128) );
  MUX2_X1 U8070 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7128), .S(n10392), .Z(n10385) );
  INV_X1 U8071 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7173) );
  MUX2_X1 U8072 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7173), .S(n6623), .Z(n6323)
         );
  OAI211_X1 U8073 ( .C1(n6324), .C2(n6323), .A(n9946), .B(n6481), .ZN(n6325)
         );
  OAI211_X1 U8074 ( .C1(n6327), .C2(n10431), .A(n6326), .B(n6325), .ZN(
        P1_U3246) );
  NAND2_X1 U8075 ( .A1(n6328), .A2(P1_B_REG_SCAN_IN), .ZN(n6329) );
  MUX2_X1 U8076 ( .A(P1_B_REG_SCAN_IN), .B(n6329), .S(n7340), .Z(n6330) );
  NAND2_X1 U8077 ( .A1(n6330), .A2(n7704), .ZN(n10337) );
  INV_X1 U8078 ( .A(n6328), .ZN(n6331) );
  OAI22_X1 U8079 ( .A1(n10337), .A2(P1_D_REG_1__SCAN_IN), .B1(n7704), .B2(
        n6331), .ZN(n7122) );
  NOR2_X1 U8080 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .ZN(
        n8740) );
  NOR4_X1 U8081 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6334) );
  NOR4_X1 U8082 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n6333) );
  NOR4_X1 U8083 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n6332) );
  AND4_X1 U8084 ( .A1(n8740), .A2(n6334), .A3(n6333), .A4(n6332), .ZN(n6340)
         );
  NOR4_X1 U8085 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6338) );
  NOR4_X1 U8086 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6337) );
  NOR4_X1 U8087 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n6336) );
  NOR4_X1 U8088 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n6335) );
  AND4_X1 U8089 ( .A1(n6338), .A2(n6337), .A3(n6336), .A4(n6335), .ZN(n6339)
         );
  NAND2_X1 U8090 ( .A1(n6340), .A2(n6339), .ZN(n6600) );
  INV_X1 U8091 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6341) );
  NOR2_X1 U8092 ( .A1(n6600), .A2(n6341), .ZN(n6343) );
  INV_X1 U8093 ( .A(n7340), .ZN(n6342) );
  OR2_X1 U8094 ( .A1(n7704), .A2(n6342), .ZN(n10338) );
  OAI21_X1 U8095 ( .B1(n10337), .B2(n6343), .A(n10338), .ZN(n6439) );
  OR2_X1 U8096 ( .A1(n7122), .A2(n6439), .ZN(n6520) );
  AND2_X1 U8097 ( .A1(n6521), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6344) );
  INV_X1 U8098 ( .A(n10453), .ZN(n6345) );
  NOR2_X1 U8099 ( .A1(n6520), .A2(n6345), .ZN(n6385) );
  INV_X1 U8100 ( .A(n8283), .ZN(n8426) );
  NAND2_X1 U8101 ( .A1(n4372), .A2(n8426), .ZN(n6610) );
  INV_X1 U8102 ( .A(n6610), .ZN(n6607) );
  AND2_X1 U8103 ( .A1(n6607), .A2(n8286), .ZN(n7129) );
  NAND2_X1 U8104 ( .A1(n6385), .A2(n7129), .ZN(n6349) );
  XNOR2_X2 U8105 ( .A(n6347), .B(P1_IR_REG_19__SCAN_IN), .ZN(n9951) );
  NAND2_X1 U8107 ( .A1(n10453), .A2(n8426), .ZN(n6348) );
  INV_X1 U8108 ( .A(SI_0_), .ZN(n6350) );
  NOR2_X1 U8109 ( .A1(n5133), .A2(n6350), .ZN(n6351) );
  XNOR2_X1 U8110 ( .A(n6351), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n10351) );
  MUX2_X1 U8111 ( .A(n6374), .B(n10351), .S(n7851), .Z(n6373) );
  AND2_X2 U8112 ( .A1(n7143), .A2(n6371), .ZN(n6402) );
  INV_X1 U8113 ( .A(n6353), .ZN(n6356) );
  INV_X1 U8114 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6354) );
  NAND2_X1 U8115 ( .A1(n6356), .A2(n5043), .ZN(n6358) );
  OAI21_X2 U8116 ( .B1(n6362), .B2(n6361), .A(n6360), .ZN(n6363) );
  NAND2_X1 U8117 ( .A1(n8184), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6370) );
  INV_X1 U8118 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n8757) );
  OR2_X1 U8119 ( .A1(n6707), .A2(n8757), .ZN(n6368) );
  NAND2_X2 U8120 ( .A1(n10348), .A2(n10343), .ZN(n6714) );
  INV_X1 U8121 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6366) );
  OR2_X1 U8122 ( .A1(n6714), .A2(n6366), .ZN(n6367) );
  INV_X1 U8123 ( .A(n9859), .ZN(n6458) );
  OR2_X1 U8124 ( .A1(n8154), .A2(n6458), .ZN(n6377) );
  INV_X1 U8125 ( .A(n6371), .ZN(n6372) );
  OR2_X4 U8126 ( .A1(n7143), .A2(n6372), .ZN(n8942) );
  OAI22_X1 U8127 ( .A1(n8942), .A2(n6373), .B1(n6374), .B2(n6024), .ZN(n6375)
         );
  INV_X1 U8128 ( .A(n6375), .ZN(n6376) );
  NAND2_X1 U8129 ( .A1(n6700), .A2(n9859), .ZN(n6379) );
  NAND2_X1 U8130 ( .A1(n6402), .A2(n6444), .ZN(n6378) );
  OAI211_X1 U8131 ( .C1(n6024), .C2(n6380), .A(n6379), .B(n6378), .ZN(n6393)
         );
  NAND2_X1 U8132 ( .A1(n6381), .A2(n6393), .ZN(n6396) );
  OAI21_X1 U8133 ( .B1(n6381), .B2(n6393), .A(n6396), .ZN(n6657) );
  OR2_X1 U8134 ( .A1(n6610), .A2(n4409), .ZN(n10454) );
  AND2_X1 U8135 ( .A1(n10454), .A2(n8434), .ZN(n6382) );
  AOI22_X1 U8136 ( .A1(n4582), .A2(n6444), .B1(n6657), .B2(n9815), .ZN(n6392)
         );
  OR2_X1 U8137 ( .A1(n10311), .A2(n8283), .ZN(n6438) );
  INV_X1 U8138 ( .A(n6438), .ZN(n6383) );
  INV_X1 U8139 ( .A(n6520), .ZN(n6424) );
  OR2_X1 U8140 ( .A1(n8434), .A2(n4409), .ZN(n6522) );
  OAI21_X1 U8141 ( .B1(n6383), .B2(n6424), .A(n7123), .ZN(n6468) );
  OR2_X1 U8142 ( .A1(n6442), .A2(n7143), .ZN(n7125) );
  NOR2_X1 U8143 ( .A1(n7125), .A2(n6451), .ZN(n6384) );
  INV_X1 U8144 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6386) );
  OR2_X1 U8145 ( .A1(n6714), .A2(n6386), .ZN(n6388) );
  AOI22_X1 U8146 ( .A1(n6468), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n9835), .B2(
        n9857), .ZN(n6391) );
  NAND2_X1 U8147 ( .A1(n6392), .A2(n6391), .ZN(P1_U3230) );
  INV_X1 U8148 ( .A(n6393), .ZN(n6394) );
  NAND2_X1 U8149 ( .A1(n6394), .A2(n8112), .ZN(n6395) );
  NAND2_X1 U8150 ( .A1(n6396), .A2(n6395), .ZN(n6406) );
  OAI22_X1 U8151 ( .A1(n6590), .A2(n8942), .B1(n6459), .B2(n4376), .ZN(n6403)
         );
  XNOR2_X1 U8153 ( .A(n6403), .B(n8938), .ZN(n6407) );
  NAND2_X1 U8154 ( .A1(n6406), .A2(n6407), .ZN(n6464) );
  OR2_X1 U8155 ( .A1(n8154), .A2(n6590), .ZN(n6405) );
  INV_X2 U8156 ( .A(n8942), .ZN(n6700) );
  NAND2_X1 U8157 ( .A1(n4367), .A2(n7195), .ZN(n6404) );
  NAND2_X1 U8158 ( .A1(n6405), .A2(n6404), .ZN(n6467) );
  NAND2_X1 U8159 ( .A1(n6464), .A2(n6467), .ZN(n6410) );
  INV_X1 U8160 ( .A(n6406), .ZN(n6409) );
  INV_X1 U8161 ( .A(n6407), .ZN(n6408) );
  NAND2_X1 U8162 ( .A1(n6409), .A2(n6408), .ZN(n6465) );
  NAND2_X1 U8163 ( .A1(n6410), .A2(n6465), .ZN(n6515) );
  INV_X1 U8164 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6411) );
  OR2_X1 U8165 ( .A1(n6714), .A2(n6411), .ZN(n6416) );
  NAND2_X1 U8166 ( .A1(n8184), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6414) );
  INV_X1 U8167 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6412) );
  OR2_X1 U8168 ( .A1(n6707), .A2(n6412), .ZN(n6413) );
  AOI22_X1 U8169 ( .A1(n8935), .A2(n9856), .B1(n8934), .B2(n8217), .ZN(n6511)
         );
  INV_X1 U8170 ( .A(n9856), .ZN(n8218) );
  INV_X1 U8171 ( .A(n8217), .ZN(n7563) );
  OAI22_X1 U8172 ( .A1(n8218), .A2(n8942), .B1(n7563), .B2(n4376), .ZN(n6422)
         );
  XNOR2_X1 U8173 ( .A(n6422), .B(n8938), .ZN(n6512) );
  XNOR2_X1 U8174 ( .A(n6511), .B(n6512), .ZN(n6514) );
  XOR2_X1 U8175 ( .A(n6515), .B(n6514), .Z(n6437) );
  NAND2_X1 U8176 ( .A1(n10453), .A2(n6451), .ZN(n6423) );
  NOR2_X1 U8177 ( .A1(n7125), .A2(n6423), .ZN(n8440) );
  NAND2_X1 U8178 ( .A1(n8440), .A2(n6424), .ZN(n9831) );
  INV_X1 U8179 ( .A(n9831), .ZN(n9785) );
  INV_X1 U8180 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6426) );
  OR2_X1 U8181 ( .A1(n6714), .A2(n6426), .ZN(n6427) );
  OAI21_X1 U8182 ( .B1(n8190), .B2(n6428), .A(n6427), .ZN(n6429) );
  INV_X1 U8183 ( .A(n6429), .ZN(n6434) );
  OR2_X1 U8184 ( .A1(n6707), .A2(n6430), .ZN(n6431) );
  INV_X1 U8185 ( .A(n6432), .ZN(n6433) );
  AOI22_X1 U8186 ( .A1(n9785), .A2(n9857), .B1(n9835), .B2(n9855), .ZN(n6436)
         );
  AOI22_X1 U8187 ( .A1(n4582), .A2(n8217), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n6468), .ZN(n6435) );
  OAI211_X1 U8188 ( .C1(n6437), .C2(n9825), .A(n6436), .B(n6435), .ZN(P1_U3235) );
  INV_X1 U8189 ( .A(n6439), .ZN(n6440) );
  AND2_X1 U8190 ( .A1(n6440), .A2(n7122), .ZN(n6441) );
  AND2_X2 U8191 ( .A1(n6605), .A2(n6441), .ZN(n10465) );
  NAND2_X1 U8192 ( .A1(n4372), .A2(n10053), .ZN(n6443) );
  MUX2_X1 U8193 ( .A(n6443), .B(n6442), .S(n7143), .Z(n7268) );
  NAND2_X1 U8194 ( .A1(n7268), .A2(n10311), .ZN(n10260) );
  CLKBUF_X1 U8195 ( .A(n6455), .Z(n6447) );
  INV_X1 U8196 ( .A(n6587), .ZN(n6449) );
  AOI21_X1 U8197 ( .B1(n6450), .B2(n6447), .A(n6449), .ZN(n7202) );
  NOR2_X1 U8198 ( .A1(n8426), .A2(n8438), .ZN(n8396) );
  INV_X1 U8199 ( .A(n8396), .ZN(n6453) );
  OR2_X1 U8200 ( .A1(n4372), .A2(n10053), .ZN(n6452) );
  NAND2_X1 U8201 ( .A1(n6453), .A2(n6452), .ZN(n10117) );
  INV_X1 U8202 ( .A(n6454), .ZN(n6606) );
  INV_X1 U8203 ( .A(n6592), .ZN(n6456) );
  AOI21_X1 U8204 ( .B1(n4500), .B2(n6606), .A(n6456), .ZN(n6457) );
  OAI222_X1 U8205 ( .A1(n10184), .A2(n8218), .B1(n10182), .B2(n6458), .C1(
        n10179), .C2(n6457), .ZN(n7199) );
  INV_X1 U8206 ( .A(n7199), .ZN(n6462) );
  INV_X2 U8207 ( .A(n10454), .ZN(n10306) );
  NAND2_X1 U8208 ( .A1(n6459), .A2(n6373), .ZN(n6596) );
  OAI211_X1 U8209 ( .C1(n6459), .C2(n6373), .A(n10307), .B(n6596), .ZN(n7197)
         );
  INV_X1 U8210 ( .A(n7197), .ZN(n6460) );
  AOI21_X1 U8211 ( .B1(n10306), .B2(n7195), .A(n6460), .ZN(n6461) );
  OAI211_X1 U8212 ( .C1(n10298), .C2(n7202), .A(n6462), .B(n6461), .ZN(n6612)
         );
  NAND2_X1 U8213 ( .A1(n6612), .A2(n10465), .ZN(n6463) );
  OAI21_X1 U8214 ( .B1(n10465), .B2(n8682), .A(n6463), .ZN(P1_U3524) );
  NAND2_X1 U8215 ( .A1(n6465), .A2(n6464), .ZN(n6466) );
  XOR2_X1 U8216 ( .A(n6467), .B(n6466), .Z(n6471) );
  AOI22_X1 U8217 ( .A1(n9785), .A2(n9859), .B1(n9835), .B2(n9856), .ZN(n6470)
         );
  AOI22_X1 U8218 ( .A1(n4582), .A2(n7195), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n6468), .ZN(n6469) );
  OAI211_X1 U8219 ( .C1(n6471), .C2(n9825), .A(n6470), .B(n6469), .ZN(P1_U3220) );
  INV_X1 U8220 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6486) );
  INV_X1 U8221 ( .A(n10393), .ZN(n10423) );
  NAND2_X1 U8222 ( .A1(n6623), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6472) );
  INV_X1 U8223 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6474) );
  MUX2_X1 U8224 ( .A(n6474), .B(P1_REG1_REG_6__SCAN_IN), .S(n6697), .Z(n6475)
         );
  AOI21_X1 U8225 ( .B1(n6476), .B2(n6475), .A(n4477), .ZN(n6477) );
  NAND2_X1 U8226 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3084), .ZN(n6719) );
  OAI21_X1 U8227 ( .B1(n10394), .B2(n6477), .A(n6719), .ZN(n6484) );
  NAND2_X1 U8228 ( .A1(n6623), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6480) );
  INV_X1 U8229 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6478) );
  MUX2_X1 U8230 ( .A(n6478), .B(P1_REG2_REG_6__SCAN_IN), .S(n6697), .Z(n6479)
         );
  AND3_X1 U8231 ( .A1(n6481), .A2(n6480), .A3(n6479), .ZN(n6482) );
  NOR3_X1 U8232 ( .A1(n10416), .A2(n6502), .A3(n6482), .ZN(n6483) );
  AOI211_X1 U8233 ( .C1(n10423), .C2(n6697), .A(n6484), .B(n6483), .ZN(n6485)
         );
  OAI21_X1 U8234 ( .B1(n10431), .B2(n6486), .A(n6485), .ZN(P1_U3247) );
  INV_X1 U8235 ( .A(n7861), .ZN(n6494) );
  INV_X1 U8236 ( .A(n8908), .ZN(n9275) );
  OAI222_X1 U8237 ( .A1(n9686), .A2(n6487), .B1(n8964), .B2(n6494), .C1(n9275), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  OR2_X1 U8238 ( .A1(n6488), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n6489) );
  NAND2_X1 U8239 ( .A1(n6489), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6492) );
  INV_X1 U8240 ( .A(n6492), .ZN(n6490) );
  NAND2_X1 U8241 ( .A1(n6490), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n6493) );
  NAND2_X1 U8242 ( .A1(n6492), .A2(n6491), .ZN(n6614) );
  AND2_X1 U8243 ( .A1(n6493), .A2(n6614), .ZN(n9932) );
  INV_X1 U8244 ( .A(n9932), .ZN(n9912) );
  OAI222_X1 U8245 ( .A1(n10350), .A2(n6495), .B1(n10347), .B2(n6494), .C1(
        n9912), .C2(P1_U3084), .ZN(P1_U3336) );
  XOR2_X1 U8246 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n7138), .Z(n6499) );
  INV_X1 U8247 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6496) );
  NOR2_X1 U8248 ( .A1(n6697), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10405) );
  INV_X1 U8249 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7011) );
  MUX2_X1 U8250 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n7011), .S(n10409), .Z(n10406) );
  OAI21_X1 U8251 ( .B1(n6496), .B2(n6541), .A(n6540), .ZN(n6497) );
  OAI21_X1 U8252 ( .B1(n7042), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6497), .ZN(
        n6498) );
  NAND2_X1 U8253 ( .A1(n6498), .A2(n6499), .ZN(n6730) );
  OAI21_X1 U8254 ( .B1(n6499), .B2(n6498), .A(n6730), .ZN(n6509) );
  INV_X1 U8255 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6501) );
  NAND2_X1 U8256 ( .A1(n10423), .A2(n7138), .ZN(n6500) );
  NAND2_X1 U8257 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7303) );
  OAI211_X1 U8258 ( .C1(n10431), .C2(n6501), .A(n6500), .B(n7303), .ZN(n6508)
         );
  INV_X1 U8259 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10402) );
  INV_X1 U8260 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6503) );
  MUX2_X1 U8261 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n6503), .S(n7042), .Z(n6504)
         );
  INV_X1 U8262 ( .A(n6504), .ZN(n6544) );
  INV_X1 U8263 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7161) );
  MUX2_X1 U8264 ( .A(n7161), .B(P1_REG2_REG_9__SCAN_IN), .S(n7138), .Z(n6505)
         );
  AOI211_X1 U8265 ( .C1(n6506), .C2(n6505), .A(n10416), .B(n6725), .ZN(n6507)
         );
  AOI211_X1 U8266 ( .C1(n10427), .C2(n6509), .A(n6508), .B(n6507), .ZN(n6510)
         );
  INV_X1 U8267 ( .A(n6510), .ZN(P1_U3250) );
  NAND2_X1 U8268 ( .A1(n6512), .A2(n6511), .ZN(n6513) );
  OR2_X1 U8269 ( .A1(n7851), .A2(n4373), .ZN(n6518) );
  OR2_X1 U8270 ( .A1(n7852), .A2(n8176), .ZN(n6517) );
  OAI22_X1 U8271 ( .A1(n6670), .A2(n8942), .B1(n4376), .B2(n10455), .ZN(n6519)
         );
  XNOR2_X1 U8272 ( .A(n6519), .B(n8135), .ZN(n6551) );
  AOI22_X1 U8273 ( .A1(n8935), .A2(n9855), .B1(n4367), .B2(n7399), .ZN(n6552)
         );
  XNOR2_X1 U8274 ( .A(n6551), .B(n6552), .ZN(n6549) );
  XOR2_X1 U8275 ( .A(n6550), .B(n6549), .Z(n6538) );
  INV_X1 U8276 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7398) );
  NAND2_X1 U8277 ( .A1(n6605), .A2(n6520), .ZN(n6525) );
  NAND3_X1 U8278 ( .A1(n6522), .A2(n6521), .A3(n6024), .ZN(n6523) );
  NAND2_X1 U8279 ( .A1(n6523), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6524) );
  NAND2_X1 U8280 ( .A1(n6525), .A2(n6524), .ZN(n9773) );
  INV_X1 U8281 ( .A(n6526), .ZN(n6527) );
  AOI21_X1 U8282 ( .B1(n9785), .B2(n9856), .A(n6527), .ZN(n6535) );
  NAND2_X1 U8283 ( .A1(n6572), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6533) );
  INV_X1 U8284 ( .A(n6565), .ZN(n6567) );
  OAI21_X1 U8285 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(P1_REG3_REG_4__SCAN_IN), 
        .A(n6567), .ZN(n7130) );
  INV_X1 U8286 ( .A(n7130), .ZN(n6528) );
  NAND2_X1 U8287 ( .A1(n8184), .A2(n6528), .ZN(n6532) );
  INV_X1 U8288 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6529) );
  OR2_X1 U8289 ( .A1(n6714), .A2(n6529), .ZN(n6531) );
  OR2_X1 U8290 ( .A1(n6707), .A2(n7128), .ZN(n6530) );
  NAND4_X1 U8291 ( .A1(n6533), .A2(n6532), .A3(n6531), .A4(n6530), .ZN(n9854)
         );
  NAND2_X1 U8292 ( .A1(n9835), .A2(n9854), .ZN(n6534) );
  OAI211_X1 U8293 ( .C1(n10455), .C2(n9838), .A(n6535), .B(n6534), .ZN(n6536)
         );
  AOI21_X1 U8294 ( .B1(n7398), .B2(n9773), .A(n6536), .ZN(n6537) );
  OAI21_X1 U8295 ( .B1(n6538), .B2(n9825), .A(n6537), .ZN(P1_U3216) );
  XNOR2_X1 U8296 ( .A(n7042), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n6539) );
  XNOR2_X1 U8297 ( .A(n6540), .B(n6539), .ZN(n6548) );
  NAND2_X1 U8298 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7287) );
  OAI21_X1 U8299 ( .B1(n10393), .B2(n6541), .A(n7287), .ZN(n6546) );
  AOI211_X1 U8300 ( .C1(n6544), .C2(n6543), .A(n10416), .B(n6542), .ZN(n6545)
         );
  AOI211_X1 U8301 ( .C1(n10410), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n6546), .B(
        n6545), .ZN(n6547) );
  OAI21_X1 U8302 ( .B1(n10394), .B2(n6548), .A(n6547), .ZN(P1_U3249) );
  INV_X1 U8303 ( .A(n9773), .ZN(n9832) );
  INV_X1 U8304 ( .A(n6551), .ZN(n6553) );
  NAND2_X1 U8305 ( .A1(n6553), .A2(n6552), .ZN(n6554) );
  INV_X1 U8306 ( .A(n9854), .ZN(n7402) );
  NAND2_X1 U8307 ( .A1(n6555), .A2(n7902), .ZN(n6559) );
  OR2_X1 U8308 ( .A1(n7851), .A2(n10392), .ZN(n6558) );
  OR2_X1 U8309 ( .A1(n7852), .A2(n6556), .ZN(n6557) );
  AND3_X2 U8310 ( .A1(n6559), .A2(n6558), .A3(n6557), .ZN(n7131) );
  OAI22_X1 U8311 ( .A1(n7402), .A2(n8942), .B1(n7131), .B2(n4376), .ZN(n6560)
         );
  XNOR2_X1 U8312 ( .A(n6560), .B(n8938), .ZN(n6621) );
  AOI22_X1 U8313 ( .A1(n8935), .A2(n9854), .B1(n8934), .B2(n6678), .ZN(n6620)
         );
  XNOR2_X1 U8314 ( .A(n6621), .B(n6620), .ZN(n6561) );
  AOI21_X1 U8315 ( .B1(n6562), .B2(n6561), .A(n9825), .ZN(n6563) );
  NAND2_X1 U8316 ( .A1(n6563), .A2(n6690), .ZN(n6577) );
  OR2_X1 U8317 ( .A1(n6707), .A2(n7173), .ZN(n6571) );
  INV_X1 U8318 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6564) );
  OR2_X1 U8319 ( .A1(n6714), .A2(n6564), .ZN(n6570) );
  INV_X1 U8320 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6566) );
  NAND2_X1 U8321 ( .A1(n6567), .A2(n6566), .ZN(n6568) );
  AND2_X1 U8322 ( .A1(n6637), .A2(n6568), .ZN(n7171) );
  NAND2_X1 U8323 ( .A1(n8184), .A2(n7171), .ZN(n6569) );
  NAND2_X1 U8324 ( .A1(n6572), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6573) );
  NAND2_X1 U8325 ( .A1(n9835), .A2(n4505), .ZN(n6574) );
  NAND2_X1 U8326 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3084), .ZN(n10399) );
  OAI211_X1 U8327 ( .C1(n6670), .C2(n9831), .A(n6574), .B(n10399), .ZN(n6575)
         );
  AOI21_X1 U8328 ( .B1(n6678), .B2(n4582), .A(n6575), .ZN(n6576) );
  OAI211_X1 U8329 ( .C1(n9832), .C2(n7130), .A(n6577), .B(n6576), .ZN(P1_U3228) );
  INV_X1 U8330 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7259) );
  INV_X1 U8331 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7493) );
  OR2_X2 U8332 ( .A1(n7494), .A2(n7493), .ZN(n7622) );
  INV_X1 U8333 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7621) );
  XNOR2_X1 U8334 ( .A(n7973), .B(P1_REG3_REG_16__SCAN_IN), .ZN(n10134) );
  NAND2_X1 U8335 ( .A1(n10134), .A2(n8184), .ZN(n6584) );
  INV_X1 U8336 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n6581) );
  INV_X1 U8337 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n8766) );
  OR2_X1 U8338 ( .A1(n8186), .A2(n8766), .ZN(n6580) );
  INV_X1 U8339 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n6578) );
  OR2_X1 U8340 ( .A1(n8187), .A2(n6578), .ZN(n6579) );
  OAI211_X1 U8341 ( .C1(n4380), .C2(n6581), .A(n6580), .B(n6579), .ZN(n6582)
         );
  INV_X1 U8342 ( .A(n6582), .ZN(n6583) );
  MUX2_X1 U8343 ( .A(n8782), .B(n9760), .S(n9858), .Z(n6585) );
  INV_X1 U8344 ( .A(n6585), .ZN(P1_U3571) );
  NAND2_X1 U8345 ( .A1(n6590), .A2(n6459), .ZN(n6586) );
  NAND2_X1 U8346 ( .A1(n6587), .A2(n6586), .ZN(n6589) );
  NAND2_X1 U8347 ( .A1(n6588), .A2(n6589), .ZN(n6669) );
  OAI21_X1 U8348 ( .B1(n6589), .B2(n6588), .A(n6669), .ZN(n7565) );
  INV_X1 U8349 ( .A(n7565), .ZN(n6598) );
  INV_X1 U8350 ( .A(n7268), .ZN(n10153) );
  OAI22_X1 U8351 ( .A1(n6590), .A2(n10182), .B1(n10184), .B2(n6670), .ZN(n6595) );
  NAND2_X1 U8352 ( .A1(n6590), .A2(n7195), .ZN(n6591) );
  XNOR2_X1 U8353 ( .A(n8220), .B(n6588), .ZN(n6593) );
  NOR2_X1 U8354 ( .A1(n6593), .A2(n10179), .ZN(n6594) );
  AOI211_X1 U8355 ( .C1(n10153), .C2(n7565), .A(n6595), .B(n6594), .ZN(n7567)
         );
  AOI21_X1 U8356 ( .B1(n8217), .B2(n6596), .A(n4404), .ZN(n7560) );
  AOI22_X1 U8357 ( .A1(n7560), .A2(n10307), .B1(n10306), .B2(n8217), .ZN(n6597) );
  OAI211_X1 U8358 ( .C1(n6598), .C2(n10311), .A(n7567), .B(n6597), .ZN(n6618)
         );
  NAND2_X1 U8359 ( .A1(n6618), .A2(n10465), .ZN(n6599) );
  OAI21_X1 U8360 ( .B1(n10465), .B2(n6282), .A(n6599), .ZN(P1_U3525) );
  INV_X1 U8361 ( .A(n10337), .ZN(n6601) );
  NAND2_X1 U8362 ( .A1(n6601), .A2(n6600), .ZN(n6603) );
  OAI21_X1 U8363 ( .B1(n10337), .B2(P1_D_REG_0__SCAN_IN), .A(n10338), .ZN(
        n6602) );
  AND2_X1 U8364 ( .A1(n6603), .A2(n6602), .ZN(n7387) );
  AND2_X1 U8365 ( .A1(n7387), .A2(n7122), .ZN(n6604) );
  NAND2_X1 U8366 ( .A1(n6605), .A2(n6604), .ZN(n10462) );
  INV_X2 U8367 ( .A(n10462), .ZN(n10335) );
  NAND2_X1 U8368 ( .A1(n9859), .A2(n6373), .ZN(n8215) );
  AND2_X1 U8369 ( .A1(n6606), .A2(n8215), .ZN(n8260) );
  INV_X1 U8370 ( .A(n7125), .ZN(n6608) );
  NOR3_X1 U8371 ( .A1(n8260), .A2(n6608), .A3(n6607), .ZN(n6609) );
  AOI21_X1 U8372 ( .B1(n10148), .B2(n9857), .A(n6609), .ZN(n10432) );
  OAI21_X1 U8373 ( .B1(n6373), .B2(n6610), .A(n10432), .ZN(n10313) );
  NAND2_X1 U8374 ( .A1(n10313), .A2(n10335), .ZN(n6611) );
  OAI21_X1 U8375 ( .B1(n10335), .B2(n6366), .A(n6611), .ZN(P1_U3454) );
  NAND2_X1 U8376 ( .A1(n6612), .A2(n10335), .ZN(n6613) );
  OAI21_X1 U8377 ( .B1(n10335), .B2(n6386), .A(n6613), .ZN(P1_U3457) );
  INV_X1 U8378 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n8786) );
  INV_X1 U8379 ( .A(n7868), .ZN(n6616) );
  OAI222_X1 U8380 ( .A1(n9686), .A2(n8786), .B1(n9684), .B2(n6616), .C1(
        P2_U3152), .C2(n4751), .ZN(P2_U3340) );
  INV_X1 U8381 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6617) );
  NAND2_X1 U8382 ( .A1(n6614), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6615) );
  XNOR2_X1 U8383 ( .A(n6615), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9944) );
  INV_X1 U8384 ( .A(n9944), .ZN(n9931) );
  OAI222_X1 U8385 ( .A1(n10350), .A2(n6617), .B1(n10347), .B2(n6616), .C1(
        P1_U3084), .C2(n9931), .ZN(P1_U3335) );
  NAND2_X1 U8386 ( .A1(n6618), .A2(n10335), .ZN(n6619) );
  OAI21_X1 U8387 ( .B1(n10335), .B2(n6411), .A(n6619), .ZN(P1_U3460) );
  OR2_X1 U8388 ( .A1(n6621), .A2(n6620), .ZN(n6688) );
  NAND2_X1 U8389 ( .A1(n6690), .A2(n6688), .ZN(n6631) );
  INV_X2 U8390 ( .A(n7852), .ZN(n7873) );
  AOI22_X1 U8391 ( .A1(n7873), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n4368), .B2(
        n6623), .ZN(n6626) );
  NAND2_X1 U8392 ( .A1(n6624), .A2(n7902), .ZN(n6625) );
  NAND2_X1 U8393 ( .A1(n8934), .A2(n4505), .ZN(n6627) );
  OAI21_X1 U8394 ( .B1(n6926), .B2(n4376), .A(n6627), .ZN(n6628) );
  XNOR2_X1 U8395 ( .A(n6628), .B(n8112), .ZN(n6691) );
  OR2_X1 U8396 ( .A1(n8154), .A2(n6934), .ZN(n6629) );
  OAI21_X1 U8397 ( .B1(n6926), .B2(n8942), .A(n6629), .ZN(n6686) );
  INV_X1 U8398 ( .A(n6686), .ZN(n6692) );
  XNOR2_X1 U8399 ( .A(n6691), .B(n6692), .ZN(n6630) );
  XNOR2_X1 U8400 ( .A(n6631), .B(n6630), .ZN(n6647) );
  OR2_X1 U8401 ( .A1(n6707), .A2(n6478), .ZN(n6634) );
  INV_X1 U8402 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6632) );
  OR2_X1 U8403 ( .A1(n6714), .A2(n6632), .ZN(n6633) );
  AND2_X1 U8404 ( .A1(n6634), .A2(n6633), .ZN(n6641) );
  INV_X1 U8405 ( .A(n6635), .ZN(n6711) );
  NAND2_X1 U8406 ( .A1(n6637), .A2(n6636), .ZN(n6638) );
  AND2_X1 U8407 ( .A1(n6711), .A2(n6638), .ZN(n7367) );
  NAND2_X1 U8408 ( .A1(n8184), .A2(n7367), .ZN(n6640) );
  NAND2_X1 U8409 ( .A1(n6572), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6639) );
  INV_X1 U8410 ( .A(n7008), .ZN(n9853) );
  NAND2_X1 U8411 ( .A1(n9835), .A2(n9853), .ZN(n6643) );
  OAI211_X1 U8412 ( .C1(n7402), .C2(n9831), .A(n6643), .B(n6642), .ZN(n6645)
         );
  NOR2_X1 U8413 ( .A1(n9838), .A2(n6926), .ZN(n6644) );
  AOI211_X1 U8414 ( .C1(n7171), .C2(n9773), .A(n6645), .B(n6644), .ZN(n6646)
         );
  OAI21_X1 U8415 ( .B1(n6647), .B2(n9825), .A(n6646), .ZN(P1_U3225) );
  INV_X1 U8416 ( .A(n6648), .ZN(n6653) );
  MUX2_X1 U8417 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6282), .S(n6649), .Z(n6652)
         );
  INV_X1 U8418 ( .A(n6650), .ZN(n6651) );
  AOI211_X1 U8419 ( .C1(n6653), .C2(n6652), .A(n6651), .B(n10394), .ZN(n6654)
         );
  AOI21_X1 U8420 ( .B1(n10423), .B2(n6655), .A(n6654), .ZN(n6660) );
  INV_X1 U8421 ( .A(n7916), .ZN(n8439) );
  MUX2_X1 U8422 ( .A(n6657), .B(n6656), .S(n8439), .Z(n6659) );
  OAI211_X1 U8423 ( .C1(n6659), .C2(n4368), .A(n9858), .B(n6658), .ZN(n10396)
         );
  OAI211_X1 U8424 ( .C1(n10431), .C2(n6661), .A(n6660), .B(n10396), .ZN(n6667)
         );
  INV_X1 U8425 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6665) );
  XNOR2_X1 U8426 ( .A(n6663), .B(n6662), .ZN(n6664) );
  OAI22_X1 U8427 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6665), .B1(n6664), .B2(
        n10416), .ZN(n6666) );
  OR2_X1 U8428 ( .A1(n6667), .A2(n6666), .ZN(P1_U3243) );
  NAND2_X1 U8429 ( .A1(n8218), .A2(n7563), .ZN(n6668) );
  NAND2_X2 U8430 ( .A1(n6670), .A2(n7399), .ZN(n8399) );
  NAND2_X1 U8431 ( .A1(n9855), .A2(n10455), .ZN(n8213) );
  NAND2_X2 U8432 ( .A1(n8399), .A2(n8213), .ZN(n7401) );
  NAND2_X1 U8433 ( .A1(n7397), .A2(n7401), .ZN(n7396) );
  NAND2_X1 U8434 ( .A1(n6670), .A2(n10455), .ZN(n6671) );
  NAND2_X1 U8435 ( .A1(n7396), .A2(n6671), .ZN(n6674) );
  NAND2_X1 U8436 ( .A1(n7402), .A2(n6678), .ZN(n8400) );
  NAND2_X1 U8437 ( .A1(n9854), .A2(n7131), .ZN(n8401) );
  NAND2_X2 U8438 ( .A1(n8400), .A2(n8401), .ZN(n8262) );
  AND2_X1 U8439 ( .A1(n6744), .A2(n6742), .ZN(n6673) );
  OAI21_X1 U8440 ( .B1(n6674), .B2(n8262), .A(n6673), .ZN(n6675) );
  INV_X1 U8441 ( .A(n6675), .ZN(n7136) );
  NAND2_X1 U8442 ( .A1(n8218), .A2(n8217), .ZN(n8221) );
  NAND2_X1 U8443 ( .A1(n6676), .A2(n8221), .ZN(n8408) );
  INV_X2 U8444 ( .A(n7401), .ZN(n8261) );
  XOR2_X1 U8445 ( .A(n6748), .B(n8262), .Z(n6677) );
  AOI222_X1 U8446 ( .A1(n10117), .A2(n6677), .B1(n4505), .B2(n10148), .C1(
        n9855), .C2(n10147), .ZN(n7127) );
  AOI21_X1 U8447 ( .B1(n6678), .B2(n4482), .A(n4403), .ZN(n7133) );
  AOI22_X1 U8448 ( .A1(n7133), .A2(n10307), .B1(n10306), .B2(n6678), .ZN(n6679) );
  OAI211_X1 U8449 ( .C1(n10298), .C2(n7136), .A(n7127), .B(n6679), .ZN(n6681)
         );
  NAND2_X1 U8450 ( .A1(n6681), .A2(n10465), .ZN(n6680) );
  OAI21_X1 U8451 ( .B1(n10465), .B2(n6308), .A(n6680), .ZN(P1_U3527) );
  NAND2_X1 U8452 ( .A1(n6681), .A2(n10335), .ZN(n6682) );
  OAI21_X1 U8453 ( .B1(n10335), .B2(n6529), .A(n6682), .ZN(P1_U3466) );
  INV_X1 U8454 ( .A(n7871), .ZN(n6684) );
  OAI222_X1 U8455 ( .A1(n9686), .A2(n6683), .B1(n9684), .B2(n6684), .C1(
        P2_U3152), .C2(n8923), .ZN(P2_U3339) );
  OAI222_X1 U8456 ( .A1(n10350), .A2(n6685), .B1(n10347), .B2(n6684), .C1(
        n10053), .C2(P1_U3084), .ZN(P1_U3334) );
  NAND2_X1 U8457 ( .A1(n6691), .A2(n6686), .ZN(n6687) );
  AND2_X1 U8458 ( .A1(n6688), .A2(n6687), .ZN(n6689) );
  NAND2_X1 U8459 ( .A1(n6690), .A2(n6689), .ZN(n6695) );
  INV_X1 U8460 ( .A(n6691), .ZN(n6693) );
  NAND2_X1 U8461 ( .A1(n6693), .A2(n6692), .ZN(n6694) );
  NAND2_X1 U8462 ( .A1(n6696), .A2(n7902), .ZN(n6699) );
  AOI22_X1 U8463 ( .A1(n7873), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n4368), .B2(
        n6697), .ZN(n6698) );
  NAND2_X1 U8464 ( .A1(n7368), .A2(n8934), .ZN(n6702) );
  NAND2_X1 U8465 ( .A1(n8935), .A2(n9853), .ZN(n6701) );
  NAND2_X1 U8466 ( .A1(n7368), .A2(n8940), .ZN(n6704) );
  NAND2_X1 U8467 ( .A1(n9853), .A2(n8934), .ZN(n6703) );
  NAND2_X1 U8468 ( .A1(n6704), .A2(n6703), .ZN(n6705) );
  XNOR2_X1 U8469 ( .A(n6705), .B(n8112), .ZN(n6880) );
  XOR2_X1 U8470 ( .A(n6882), .B(n6880), .Z(n6706) );
  XNOR2_X1 U8471 ( .A(n6883), .B(n6706), .ZN(n6724) );
  OR2_X1 U8472 ( .A1(n6707), .A2(n10402), .ZN(n6708) );
  OAI21_X1 U8473 ( .B1(n8190), .B2(n7011), .A(n6708), .ZN(n6709) );
  INV_X1 U8474 ( .A(n6709), .ZN(n6718) );
  INV_X1 U8475 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6710) );
  NAND2_X1 U8476 ( .A1(n6711), .A2(n6710), .ZN(n6712) );
  NAND2_X1 U8477 ( .A1(n6903), .A2(n6712), .ZN(n6899) );
  INV_X1 U8478 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6713) );
  OR2_X1 U8479 ( .A1(n6714), .A2(n6713), .ZN(n6715) );
  OAI21_X1 U8480 ( .B1(n7050), .B2(n6899), .A(n6715), .ZN(n6716) );
  INV_X1 U8481 ( .A(n6716), .ZN(n6717) );
  INV_X1 U8482 ( .A(n7289), .ZN(n9852) );
  NAND2_X1 U8483 ( .A1(n9835), .A2(n9852), .ZN(n6720) );
  OAI211_X1 U8484 ( .C1(n6934), .C2(n9831), .A(n6720), .B(n6719), .ZN(n6721)
         );
  AOI21_X1 U8485 ( .B1(n7367), .B2(n9773), .A(n6721), .ZN(n6723) );
  NAND2_X1 U8486 ( .A1(n4582), .A2(n7368), .ZN(n6722) );
  OAI211_X1 U8487 ( .C1(n6724), .C2(n9825), .A(n6723), .B(n6722), .ZN(P1_U3237) );
  INV_X1 U8488 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6740) );
  INV_X1 U8489 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n8579) );
  AOI22_X1 U8490 ( .A1(n7250), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8579), .B2(
        n6734), .ZN(n6727) );
  INV_X1 U8491 ( .A(n6729), .ZN(n10422) );
  INV_X1 U8492 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7145) );
  XNOR2_X1 U8493 ( .A(n6729), .B(n7145), .ZN(n10418) );
  OAI21_X1 U8494 ( .B1(n6727), .B2(n6726), .A(n7116), .ZN(n6728) );
  NAND2_X1 U8495 ( .A1(n6728), .A2(n9946), .ZN(n6739) );
  INV_X1 U8496 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7147) );
  XNOR2_X1 U8497 ( .A(n6729), .B(n7147), .ZN(n10425) );
  INV_X1 U8498 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6731) );
  AOI22_X1 U8499 ( .A1(n7250), .A2(P1_REG1_REG_11__SCAN_IN), .B1(n6731), .B2(
        n6734), .ZN(n6732) );
  OAI21_X1 U8500 ( .B1(n6733), .B2(n6732), .A(n7109), .ZN(n6737) );
  NAND2_X1 U8501 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7360) );
  INV_X1 U8502 ( .A(n7360), .ZN(n6736) );
  NOR2_X1 U8503 ( .A1(n10393), .A2(n6734), .ZN(n6735) );
  AOI211_X1 U8504 ( .C1(n10427), .C2(n6737), .A(n6736), .B(n6735), .ZN(n6738)
         );
  OAI211_X1 U8505 ( .C1(n10431), .C2(n6740), .A(n6739), .B(n6738), .ZN(
        P1_U3252) );
  NAND2_X1 U8506 ( .A1(n7402), .A2(n7131), .ZN(n6741) );
  AND2_X1 U8507 ( .A1(n6742), .A2(n6741), .ZN(n6743) );
  NAND2_X1 U8508 ( .A1(n6744), .A2(n6743), .ZN(n7036) );
  INV_X1 U8509 ( .A(n6998), .ZN(n6747) );
  AND2_X2 U8510 ( .A1(n7004), .A2(n8403), .ZN(n8265) );
  INV_X1 U8511 ( .A(n8265), .ZN(n6746) );
  OR2_X1 U8512 ( .A1(n6998), .A2(n8265), .ZN(n6927) );
  OAI21_X1 U8513 ( .B1(n6747), .B2(n6746), .A(n6927), .ZN(n7177) );
  XOR2_X1 U8514 ( .A(n8265), .B(n8296), .Z(n6749) );
  OAI222_X1 U8515 ( .A1(n10182), .A2(n7402), .B1(n10184), .B2(n7008), .C1(
        n6749), .C2(n10179), .ZN(n7169) );
  INV_X1 U8516 ( .A(n7169), .ZN(n6752) );
  OAI211_X1 U8517 ( .C1(n4403), .C2(n6926), .A(n10307), .B(n6930), .ZN(n7168)
         );
  INV_X1 U8518 ( .A(n7168), .ZN(n6750) );
  AOI21_X1 U8519 ( .B1(n10306), .B2(n7174), .A(n6750), .ZN(n6751) );
  OAI211_X1 U8520 ( .C1(n10298), .C2(n7177), .A(n6752), .B(n6751), .ZN(n6832)
         );
  NAND2_X1 U8521 ( .A1(n6832), .A2(n10465), .ZN(n6753) );
  OAI21_X1 U8522 ( .B1(n10465), .B2(n6310), .A(n6753), .ZN(P1_U3528) );
  NOR2_X1 U8523 ( .A1(n6983), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6986) );
  AOI21_X1 U8524 ( .B1(n6983), .B2(P2_REG2_REG_13__SCAN_IN), .A(n6986), .ZN(
        n6765) );
  MUX2_X1 U8525 ( .A(n6754), .B(P2_REG2_REG_2__SCAN_IN), .S(n7083), .Z(n7079)
         );
  XOR2_X1 U8526 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6961), .Z(n6952) );
  AND2_X1 U8527 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n6951) );
  AOI22_X1 U8528 ( .A1(n6952), .A2(n6951), .B1(P2_REG2_REG_1__SCAN_IN), .B2(
        n6961), .ZN(n7080) );
  NOR2_X1 U8529 ( .A1(n6755), .A2(n6754), .ZN(n9182) );
  MUX2_X1 U8530 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6756), .S(n9179), .Z(n9184)
         );
  NAND2_X1 U8531 ( .A1(n9179), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8526) );
  MUX2_X1 U8532 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n5068), .S(n8530), .Z(n8525)
         );
  NOR2_X1 U8533 ( .A1(n8530), .A2(n5068), .ZN(n9196) );
  MUX2_X1 U8534 ( .A(n6757), .B(P2_REG2_REG_5__SCAN_IN), .S(n9197), .Z(n6758)
         );
  NAND2_X1 U8535 ( .A1(n9194), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6921) );
  MUX2_X1 U8536 ( .A(n6759), .B(P2_REG2_REG_6__SCAN_IN), .S(n6919), .Z(n6920)
         );
  NOR2_X1 U8537 ( .A1(n6760), .A2(n6759), .ZN(n9213) );
  MUX2_X1 U8538 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6761), .S(n9210), .Z(n9212)
         );
  NAND2_X1 U8539 ( .A1(n9210), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9227) );
  INV_X1 U8540 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6762) );
  MUX2_X1 U8541 ( .A(n6762), .B(P2_REG2_REG_8__SCAN_IN), .S(n9223), .Z(n9226)
         );
  NOR2_X1 U8542 ( .A1(n6763), .A2(n6762), .ZN(n9239) );
  MUX2_X1 U8543 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7721), .S(n9247), .Z(n9238)
         );
  NAND2_X1 U8544 ( .A1(n9247), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6849) );
  MUX2_X1 U8545 ( .A(n7676), .B(P2_REG2_REG_10__SCAN_IN), .S(n6796), .Z(n6848)
         );
  AOI21_X1 U8546 ( .B1(n6796), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6860), .ZN(
        n9253) );
  MUX2_X1 U8547 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n7689), .S(n9262), .Z(n9254)
         );
  MUX2_X1 U8548 ( .A(n5317), .B(P2_REG2_REG_12__SCAN_IN), .S(n6800), .Z(n7022)
         );
  NAND2_X1 U8549 ( .A1(n6764), .A2(n6765), .ZN(n6989) );
  OAI21_X1 U8550 ( .B1(n6765), .B2(n6764), .A(n6989), .ZN(n6779) );
  NAND2_X1 U8551 ( .A1(n6766), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7792) );
  OAI21_X1 U8552 ( .B1(n6768), .B2(n7792), .A(n6767), .ZN(n6769) );
  OR2_X1 U8553 ( .A1(n6770), .A2(n6769), .ZN(n6772) );
  NAND2_X1 U8554 ( .A1(n6772), .A2(n6771), .ZN(n6805) );
  INV_X2 U8555 ( .A(P2_U3966), .ZN(n9178) );
  NAND2_X1 U8556 ( .A1(n6805), .A2(n9178), .ZN(n6775) );
  NOR2_X1 U8557 ( .A1(n6774), .A2(n7757), .ZN(n6773) );
  NAND2_X1 U8558 ( .A1(n6775), .A2(n6774), .ZN(n9286) );
  NAND2_X1 U8559 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9087) );
  NAND2_X1 U8560 ( .A1(n9289), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6776) );
  OAI211_X1 U8561 ( .C1(n9286), .C2(n6777), .A(n9087), .B(n6776), .ZN(n6778)
         );
  AOI21_X1 U8562 ( .B1(n6779), .B2(n9291), .A(n6778), .ZN(n6808) );
  XNOR2_X1 U8563 ( .A(n6983), .B(n8645), .ZN(n6803) );
  INV_X1 U8564 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6780) );
  XNOR2_X1 U8565 ( .A(n7083), .B(n6780), .ZN(n7076) );
  INV_X1 U8566 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6781) );
  XNOR2_X1 U8567 ( .A(n6961), .B(n6781), .ZN(n6954) );
  NAND2_X1 U8568 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n6958) );
  INV_X1 U8569 ( .A(n6958), .ZN(n6782) );
  NAND2_X1 U8570 ( .A1(n6954), .A2(n6782), .ZN(n6955) );
  NAND2_X1 U8571 ( .A1(n6961), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6783) );
  NAND2_X1 U8572 ( .A1(n6955), .A2(n6783), .ZN(n7075) );
  NAND2_X1 U8573 ( .A1(n7076), .A2(n7075), .ZN(n7074) );
  NAND2_X1 U8574 ( .A1(n7083), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6784) );
  NAND2_X1 U8575 ( .A1(n7074), .A2(n6784), .ZN(n9188) );
  XNOR2_X1 U8576 ( .A(n9179), .B(n6785), .ZN(n9189) );
  NAND2_X1 U8577 ( .A1(n9188), .A2(n9189), .ZN(n9187) );
  NAND2_X1 U8578 ( .A1(n9179), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6786) );
  NAND2_X1 U8579 ( .A1(n9187), .A2(n6786), .ZN(n8519) );
  MUX2_X1 U8580 ( .A(n6787), .B(P2_REG1_REG_4__SCAN_IN), .S(n8530), .Z(n8520)
         );
  NAND2_X1 U8581 ( .A1(n8519), .A2(n8520), .ZN(n8518) );
  OR2_X1 U8582 ( .A1(n8530), .A2(n6787), .ZN(n6788) );
  NAND2_X1 U8583 ( .A1(n8518), .A2(n6788), .ZN(n9204) );
  XNOR2_X1 U8584 ( .A(n9197), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n9205) );
  NAND2_X1 U8585 ( .A1(n9204), .A2(n9205), .ZN(n9203) );
  NAND2_X1 U8586 ( .A1(n9194), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6789) );
  NAND2_X1 U8587 ( .A1(n9203), .A2(n6789), .ZN(n6914) );
  INV_X1 U8588 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10517) );
  MUX2_X1 U8589 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10517), .S(n6919), .Z(n6915)
         );
  NAND2_X1 U8590 ( .A1(n6914), .A2(n6915), .ZN(n6913) );
  NAND2_X1 U8591 ( .A1(n6919), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6790) );
  NAND2_X1 U8592 ( .A1(n6913), .A2(n6790), .ZN(n9217) );
  INV_X1 U8593 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10520) );
  MUX2_X1 U8594 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10520), .S(n9210), .Z(n9218)
         );
  NAND2_X1 U8595 ( .A1(n9217), .A2(n9218), .ZN(n9216) );
  NAND2_X1 U8596 ( .A1(n9210), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6791) );
  NAND2_X1 U8597 ( .A1(n9216), .A2(n6791), .ZN(n9232) );
  XNOR2_X1 U8598 ( .A(n9223), .B(n6792), .ZN(n9233) );
  NAND2_X1 U8599 ( .A1(n9232), .A2(n9233), .ZN(n9231) );
  NAND2_X1 U8600 ( .A1(n9223), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6793) );
  NAND2_X1 U8601 ( .A1(n9231), .A2(n6793), .ZN(n9245) );
  XNOR2_X1 U8602 ( .A(n9247), .B(n8731), .ZN(n9246) );
  NAND2_X1 U8603 ( .A1(n9245), .A2(n9246), .ZN(n9244) );
  NAND2_X1 U8604 ( .A1(n9247), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6794) );
  NAND2_X1 U8605 ( .A1(n9244), .A2(n6794), .ZN(n6855) );
  XNOR2_X1 U8606 ( .A(n6796), .B(n6795), .ZN(n6856) );
  NAND2_X1 U8607 ( .A1(n6855), .A2(n6856), .ZN(n6854) );
  NAND2_X1 U8608 ( .A1(n6796), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6797) );
  NAND2_X1 U8609 ( .A1(n6854), .A2(n6797), .ZN(n9261) );
  XNOR2_X1 U8610 ( .A(n9262), .B(n6798), .ZN(n9260) );
  NAND2_X1 U8611 ( .A1(n9261), .A2(n9260), .ZN(n9259) );
  NAND2_X1 U8612 ( .A1(n9262), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6799) );
  NAND2_X1 U8613 ( .A1(n9259), .A2(n6799), .ZN(n7025) );
  XNOR2_X1 U8614 ( .A(n6800), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n7024) );
  NAND2_X1 U8615 ( .A1(n7030), .A2(n8788), .ZN(n6801) );
  NAND2_X1 U8616 ( .A1(n7027), .A2(n6801), .ZN(n6802) );
  NAND2_X1 U8617 ( .A1(n6802), .A2(n6803), .ZN(n6985) );
  OAI21_X1 U8618 ( .B1(n6803), .B2(n6802), .A(n6985), .ZN(n6806) );
  NAND2_X1 U8619 ( .A1(n6806), .A2(n9258), .ZN(n6807) );
  NAND2_X1 U8620 ( .A1(n6808), .A2(n6807), .ZN(P2_U3258) );
  OAI21_X1 U8621 ( .B1(n6810), .B2(n6815), .A(n6809), .ZN(n8831) );
  INV_X1 U8622 ( .A(n6811), .ZN(n6838) );
  INV_X1 U8623 ( .A(n7530), .ZN(n6812) );
  OAI21_X1 U8624 ( .B1(n8834), .B2(n6838), .A(n6812), .ZN(n8827) );
  OAI22_X1 U8625 ( .A1(n8827), .A2(n9538), .B1(n8834), .B2(n10507), .ZN(n6820)
         );
  NAND2_X1 U8626 ( .A1(n6813), .A2(n6814), .ZN(n6816) );
  XNOR2_X1 U8627 ( .A(n6816), .B(n4604), .ZN(n6817) );
  NAND2_X1 U8628 ( .A1(n6817), .A2(n9524), .ZN(n6819) );
  NAND2_X1 U8629 ( .A1(n6819), .A2(n6818), .ZN(n8830) );
  AOI211_X1 U8630 ( .C1(n10510), .C2(n8831), .A(n6820), .B(n8830), .ZN(n6981)
         );
  OR2_X1 U8631 ( .A1(n6981), .A2(n10519), .ZN(n6821) );
  OAI21_X1 U8632 ( .B1(n10522), .B2(n6787), .A(n6821), .ZN(P2_U3524) );
  OAI21_X1 U8633 ( .B1(n6823), .B2(n6827), .A(n6822), .ZN(n7323) );
  OAI21_X1 U8634 ( .B1(n9537), .B2(n8825), .A(n6839), .ZN(n7315) );
  OAI22_X1 U8635 ( .A1(n7315), .A2(n9538), .B1(n8825), .B2(n10507), .ZN(n6830)
         );
  INV_X1 U8636 ( .A(n9524), .ZN(n9442) );
  INV_X1 U8637 ( .A(n6824), .ZN(n6825) );
  AOI21_X1 U8638 ( .B1(n6827), .B2(n6826), .A(n6825), .ZN(n6828) );
  OAI222_X1 U8639 ( .A1(n9528), .A2(n6946), .B1(n9531), .B2(n6829), .C1(n9442), 
        .C2(n6828), .ZN(n7317) );
  AOI211_X1 U8640 ( .C1(n10510), .C2(n7323), .A(n6830), .B(n7317), .ZN(n6979)
         );
  OR2_X1 U8641 ( .A1(n6979), .A2(n10519), .ZN(n6831) );
  OAI21_X1 U8642 ( .B1(n10522), .B2(n6780), .A(n6831), .ZN(P2_U3522) );
  NAND2_X1 U8643 ( .A1(n6832), .A2(n10335), .ZN(n6833) );
  OAI21_X1 U8644 ( .B1(n10335), .B2(n6564), .A(n6833), .ZN(P1_U3469) );
  INV_X1 U8645 ( .A(n7876), .ZN(n6834) );
  OAI222_X1 U8646 ( .A1(n9686), .A2(n8730), .B1(n9684), .B2(n6834), .C1(n4822), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  OAI222_X1 U8647 ( .A1(P1_U3084), .A2(n8438), .B1(n10347), .B2(n6834), .C1(
        n7877), .C2(n10350), .ZN(P1_U3333) );
  INV_X1 U8648 ( .A(n9634), .ZN(n7735) );
  OAI21_X1 U8649 ( .B1(n6837), .B2(n6836), .A(n6835), .ZN(n7418) );
  INV_X1 U8650 ( .A(n7418), .ZN(n6845) );
  AOI22_X1 U8651 ( .A1(n9462), .A2(n6051), .B1(n9176), .B2(n9464), .ZN(n6873)
         );
  OAI21_X1 U8652 ( .B1(n6842), .B2(n6841), .A(n6813), .ZN(n6843) );
  NAND2_X1 U8653 ( .A1(n6843), .A2(n9524), .ZN(n6844) );
  OAI211_X1 U8654 ( .C1(n6845), .C2(n7741), .A(n6873), .B(n6844), .ZN(n7412)
         );
  AOI211_X1 U8655 ( .C1(n7735), .C2(n7418), .A(n7413), .B(n7412), .ZN(n7245)
         );
  OAI22_X1 U8656 ( .A1(n9615), .A2(n7415), .B1(n10522), .B2(n6785), .ZN(n6846)
         );
  INV_X1 U8657 ( .A(n6846), .ZN(n6847) );
  OAI21_X1 U8658 ( .B1(n7245), .B2(n10519), .A(n6847), .ZN(P2_U3523) );
  NAND3_X1 U8659 ( .A1(n9242), .A2(n6849), .A3(n6848), .ZN(n6850) );
  NAND2_X1 U8660 ( .A1(n6850), .A2(n9291), .ZN(n6859) );
  NOR2_X1 U8661 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8720), .ZN(n6853) );
  NOR2_X1 U8662 ( .A1(n9286), .A2(n6851), .ZN(n6852) );
  AOI211_X1 U8663 ( .C1(n9289), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n6853), .B(
        n6852), .ZN(n6858) );
  OAI211_X1 U8664 ( .C1(n6856), .C2(n6855), .A(n9258), .B(n6854), .ZN(n6857)
         );
  OAI211_X1 U8665 ( .C1(n6860), .C2(n6859), .A(n6858), .B(n6857), .ZN(P2_U3255) );
  INV_X1 U8666 ( .A(n6861), .ZN(n6863) );
  NAND2_X1 U8667 ( .A1(n6863), .A2(n6862), .ZN(n6864) );
  XNOR2_X1 U8668 ( .A(n6865), .B(n6864), .ZN(n6870) );
  INV_X1 U8669 ( .A(n9073), .ZN(n9133) );
  OAI22_X1 U8670 ( .A1(n9531), .A2(n6866), .B1(n7100), .B2(n9528), .ZN(n7528)
         );
  AOI22_X1 U8671 ( .A1(n9133), .A2(n7528), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n6867) );
  OAI21_X1 U8672 ( .B1(n9131), .B2(n7533), .A(n6867), .ZN(n6868) );
  AOI21_X1 U8673 ( .B1(n4606), .B2(n9122), .A(n6868), .ZN(n6869) );
  OAI21_X1 U8674 ( .B1(n9138), .B2(n6870), .A(n6869), .ZN(P2_U3229) );
  XNOR2_X1 U8675 ( .A(n6872), .B(n6871), .ZN(n6877) );
  INV_X1 U8676 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9180) );
  OAI22_X1 U8677 ( .A1(n9073), .A2(n6873), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9180), .ZN(n6875) );
  NOR2_X1 U8678 ( .A1(n9153), .A2(n7415), .ZN(n6874) );
  AOI211_X1 U8679 ( .C1(n9143), .C2(n9180), .A(n6875), .B(n6874), .ZN(n6876)
         );
  OAI21_X1 U8680 ( .B1(n6877), .B2(n9138), .A(n6876), .ZN(P2_U3220) );
  INV_X1 U8681 ( .A(n7880), .ZN(n6879) );
  OAI222_X1 U8682 ( .A1(n9686), .A2(n8795), .B1(n9684), .B2(n6879), .C1(n6878), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  OAI222_X1 U8683 ( .A1(P1_U3084), .A2(n8426), .B1(n10347), .B2(n6879), .C1(
        n8629), .C2(n10350), .ZN(P1_U3332) );
  NAND2_X1 U8684 ( .A1(n6883), .A2(n6882), .ZN(n6881) );
  NAND2_X1 U8685 ( .A1(n6881), .A2(n6880), .ZN(n6884) );
  NAND2_X1 U8686 ( .A1(n6884), .A2(n5049), .ZN(n7212) );
  NAND2_X1 U8687 ( .A1(n6999), .A2(n8940), .ZN(n6889) );
  NAND2_X1 U8688 ( .A1(n9852), .A2(n8934), .ZN(n6888) );
  NAND2_X1 U8689 ( .A1(n6889), .A2(n6888), .ZN(n6890) );
  XNOR2_X1 U8690 ( .A(n6890), .B(n8112), .ZN(n6896) );
  INV_X1 U8691 ( .A(n6896), .ZN(n6894) );
  NAND2_X1 U8692 ( .A1(n6999), .A2(n4367), .ZN(n6892) );
  OR2_X1 U8693 ( .A1(n8154), .A2(n7289), .ZN(n6891) );
  NAND2_X1 U8694 ( .A1(n6892), .A2(n6891), .ZN(n6895) );
  INV_X1 U8695 ( .A(n6895), .ZN(n6893) );
  NAND2_X1 U8696 ( .A1(n6894), .A2(n6893), .ZN(n7210) );
  INV_X1 U8697 ( .A(n7210), .ZN(n6897) );
  NOR2_X1 U8698 ( .A1(n6897), .A2(n7211), .ZN(n6898) );
  XNOR2_X1 U8699 ( .A(n7212), .B(n6898), .ZN(n6912) );
  INV_X1 U8700 ( .A(n6899), .ZN(n7386) );
  INV_X1 U8701 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n8694) );
  OR2_X1 U8702 ( .A1(n8186), .A2(n8694), .ZN(n6901) );
  OR2_X1 U8703 ( .A1(n8187), .A2(n6503), .ZN(n6900) );
  AND2_X1 U8704 ( .A1(n6901), .A2(n6900), .ZN(n6907) );
  NAND2_X1 U8705 ( .A1(n6903), .A2(n6902), .ZN(n6904) );
  AND2_X1 U8706 ( .A1(n7052), .A2(n6904), .ZN(n7376) );
  NAND2_X1 U8707 ( .A1(n8184), .A2(n7376), .ZN(n6906) );
  NAND2_X1 U8708 ( .A1(n4379), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6905) );
  AND3_X2 U8709 ( .A1(n6907), .A2(n6906), .A3(n6905), .ZN(n7305) );
  INV_X1 U8710 ( .A(n7305), .ZN(n9851) );
  NAND2_X1 U8711 ( .A1(n9835), .A2(n9851), .ZN(n6908) );
  NAND2_X1 U8712 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3084), .ZN(n10412) );
  OAI211_X1 U8713 ( .C1(n7008), .C2(n9831), .A(n6908), .B(n10412), .ZN(n6909)
         );
  AOI21_X1 U8714 ( .B1(n7386), .B2(n9773), .A(n6909), .ZN(n6911) );
  NAND2_X1 U8715 ( .A1(n4582), .A2(n6999), .ZN(n6910) );
  OAI211_X1 U8716 ( .C1(n6912), .C2(n9825), .A(n6911), .B(n6910), .ZN(P1_U3211) );
  INV_X1 U8717 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6917) );
  OAI211_X1 U8718 ( .C1(n6915), .C2(n6914), .A(n9258), .B(n6913), .ZN(n6916)
         );
  NAND2_X1 U8719 ( .A1(P2_U3152), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7090) );
  OAI211_X1 U8720 ( .C1(n8927), .C2(n6917), .A(n6916), .B(n7090), .ZN(n6918)
         );
  AOI21_X1 U8721 ( .B1(n6919), .B2(n9263), .A(n6918), .ZN(n6925) );
  INV_X1 U8722 ( .A(n9214), .ZN(n6923) );
  NAND3_X1 U8723 ( .A1(n9202), .A2(n6921), .A3(n6920), .ZN(n6922) );
  NAND3_X1 U8724 ( .A1(n9291), .A2(n6923), .A3(n6922), .ZN(n6924) );
  NAND2_X1 U8725 ( .A1(n6925), .A2(n6924), .ZN(P2_U3251) );
  INV_X1 U8726 ( .A(n10311), .ZN(n10461) );
  NAND2_X1 U8727 ( .A1(n6927), .A2(n4406), .ZN(n6929) );
  XNOR2_X1 U8728 ( .A(n6929), .B(n8294), .ZN(n7374) );
  NAND2_X1 U8729 ( .A1(n6930), .A2(n7368), .ZN(n6931) );
  NAND2_X1 U8730 ( .A1(n7001), .A2(n6931), .ZN(n7370) );
  OAI22_X1 U8731 ( .A1(n7370), .A2(n10456), .B1(n6932), .B2(n10454), .ZN(n6939) );
  NAND2_X1 U8732 ( .A1(n7374), .A2(n10153), .ZN(n6938) );
  NAND2_X1 U8733 ( .A1(n8296), .A2(n7004), .ZN(n6933) );
  XNOR2_X1 U8734 ( .A(n8291), .B(n8294), .ZN(n6936) );
  OAI22_X1 U8735 ( .A1(n7289), .A2(n10184), .B1(n10182), .B2(n6934), .ZN(n6935) );
  AOI21_X1 U8736 ( .B1(n6936), .B2(n10117), .A(n6935), .ZN(n6937) );
  NAND2_X1 U8737 ( .A1(n6938), .A2(n6937), .ZN(n7371) );
  AOI211_X1 U8738 ( .C1(n10461), .C2(n7374), .A(n6939), .B(n7371), .ZN(n7072)
         );
  INV_X1 U8739 ( .A(n10465), .ZN(n10463) );
  NAND2_X1 U8740 ( .A1(n10463), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6940) );
  OAI21_X1 U8741 ( .B1(n7072), .B2(n10463), .A(n6940), .ZN(P1_U3529) );
  INV_X1 U8742 ( .A(n6942), .ZN(n6944) );
  NOR2_X1 U8743 ( .A1(n6944), .A2(n6943), .ZN(n6945) );
  XNOR2_X1 U8744 ( .A(n6941), .B(n6945), .ZN(n6950) );
  NAND2_X1 U8745 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n8517) );
  OAI21_X1 U8746 ( .B1(n9148), .B2(n7088), .A(n8517), .ZN(n6948) );
  OAI22_X1 U8747 ( .A1(n9131), .A2(n8826), .B1(n6946), .B2(n9145), .ZN(n6947)
         );
  AOI211_X1 U8748 ( .C1(n5104), .C2(n9122), .A(n6948), .B(n6947), .ZN(n6949)
         );
  OAI21_X1 U8749 ( .B1(n6950), .B2(n9138), .A(n6949), .ZN(P2_U3232) );
  INV_X1 U8750 ( .A(n9291), .ZN(n8921) );
  XNOR2_X1 U8751 ( .A(n6952), .B(n6951), .ZN(n6963) );
  OAI22_X1 U8752 ( .A1(n8927), .A2(n10527), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6953), .ZN(n6960) );
  INV_X1 U8753 ( .A(n6954), .ZN(n6957) );
  INV_X1 U8754 ( .A(n6955), .ZN(n6956) );
  AOI211_X1 U8755 ( .C1(n6958), .C2(n6957), .A(n6956), .B(n9295), .ZN(n6959)
         );
  AOI211_X1 U8756 ( .C1(n9263), .C2(n6961), .A(n6960), .B(n6959), .ZN(n6962)
         );
  OAI21_X1 U8757 ( .B1(n8921), .B2(n6963), .A(n6962), .ZN(P2_U3246) );
  INV_X1 U8758 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6964) );
  OAI22_X1 U8759 ( .A1(n8921), .A2(n8758), .B1(n6964), .B2(n9295), .ZN(n6967)
         );
  NAND2_X1 U8760 ( .A1(n9291), .A2(n8758), .ZN(n6965) );
  OAI211_X1 U8761 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n9295), .A(n6965), .B(
        n9286), .ZN(n6966) );
  MUX2_X1 U8762 ( .A(n6967), .B(n6966), .S(P2_IR_REG_0__SCAN_IN), .Z(n6970) );
  INV_X1 U8763 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6968) );
  OAI22_X1 U8764 ( .A1(n8927), .A2(n6968), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7555), .ZN(n6969) );
  OR2_X1 U8765 ( .A1(n6970), .A2(n6969), .ZN(P2_U3245) );
  INV_X1 U8766 ( .A(n9138), .ZN(n9105) );
  OAI21_X1 U8767 ( .B1(n6973), .B2(n6972), .A(n6971), .ZN(n6974) );
  INV_X1 U8768 ( .A(n9148), .ZN(n8819) );
  AOI22_X1 U8769 ( .A1(n9105), .A2(n6974), .B1(n8819), .B2(n6051), .ZN(n6978)
         );
  INV_X1 U8770 ( .A(n9145), .ZN(n8822) );
  OR2_X1 U8771 ( .A1(n6975), .A2(P2_U3152), .ZN(n8821) );
  AOI22_X1 U8772 ( .A1(n8822), .A2(n6976), .B1(n8821), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n6977) );
  OAI211_X1 U8773 ( .C1(n10488), .C2(n9153), .A(n6978), .B(n6977), .ZN(
        P2_U3224) );
  OR2_X1 U8774 ( .A1(n6979), .A2(n10512), .ZN(n6980) );
  OAI21_X1 U8775 ( .B1(n10513), .B2(n5142), .A(n6980), .ZN(P2_U3457) );
  OR2_X1 U8776 ( .A1(n6981), .A2(n10512), .ZN(n6982) );
  OAI21_X1 U8777 ( .B1(n10513), .B2(n5067), .A(n6982), .ZN(P2_U3463) );
  XNOR2_X1 U8778 ( .A(n6992), .B(n8744), .ZN(n7186) );
  OR2_X1 U8779 ( .A1(n6983), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6984) );
  NAND2_X1 U8780 ( .A1(n6985), .A2(n6984), .ZN(n7187) );
  XOR2_X1 U8781 ( .A(n7186), .B(n7187), .Z(n6995) );
  INV_X1 U8782 ( .A(n6986), .ZN(n6987) );
  MUX2_X1 U8783 ( .A(n7179), .B(P2_REG2_REG_14__SCAN_IN), .S(n6992), .Z(n6988)
         );
  AOI21_X1 U8784 ( .B1(n6989), .B2(n6987), .A(n6988), .ZN(n7178) );
  AND3_X1 U8785 ( .A1(n6989), .A2(n6988), .A3(n6987), .ZN(n6990) );
  OAI21_X1 U8786 ( .B1(n7178), .B2(n6990), .A(n9291), .ZN(n6994) );
  NAND2_X1 U8787 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8972) );
  OAI21_X1 U8788 ( .B1(n8927), .B2(n4523), .A(n8972), .ZN(n6991) );
  AOI21_X1 U8789 ( .B1(n9263), .B2(n6992), .A(n6991), .ZN(n6993) );
  OAI211_X1 U8790 ( .C1(n6995), .C2(n9295), .A(n6994), .B(n6993), .ZN(P2_U3259) );
  NAND2_X1 U8791 ( .A1(n4406), .A2(n8265), .ZN(n6996) );
  AOI21_X1 U8792 ( .B1(n6998), .B2(n6997), .A(n7038), .ZN(n7000) );
  OR2_X2 U8793 ( .A1(n6999), .A2(n7289), .ZN(n8299) );
  NAND2_X2 U8794 ( .A1(n6999), .A2(n7289), .ZN(n8298) );
  AND2_X2 U8795 ( .A1(n8299), .A2(n8298), .ZN(n8293) );
  INV_X1 U8796 ( .A(n8293), .ZN(n7060) );
  XNOR2_X1 U8797 ( .A(n7000), .B(n7060), .ZN(n7390) );
  AOI211_X1 U8798 ( .C1(n6999), .C2(n7001), .A(n10456), .B(n7047), .ZN(n7393)
         );
  AND2_X1 U8799 ( .A1(n8400), .A2(n8403), .ZN(n7002) );
  AND2_X1 U8800 ( .A1(n8405), .A2(n7002), .ZN(n8225) );
  INV_X1 U8801 ( .A(n7004), .ZN(n8292) );
  NAND2_X1 U8802 ( .A1(n8405), .A2(n8292), .ZN(n8211) );
  AND2_X1 U8803 ( .A1(n8211), .A2(n8210), .ZN(n7005) );
  XNOR2_X1 U8804 ( .A(n7061), .B(n8293), .ZN(n7007) );
  OAI222_X1 U8805 ( .A1(n10184), .A2(n7305), .B1(n10182), .B2(n7008), .C1(
        n10179), .C2(n7007), .ZN(n7385) );
  AOI211_X1 U8806 ( .C1(n10306), .C2(n6999), .A(n7393), .B(n7385), .ZN(n7009)
         );
  OAI21_X1 U8807 ( .B1(n10298), .B2(n7390), .A(n7009), .ZN(n7012) );
  NAND2_X1 U8808 ( .A1(n7012), .A2(n10465), .ZN(n7010) );
  OAI21_X1 U8809 ( .B1(n10465), .B2(n7011), .A(n7010), .ZN(P1_U3530) );
  NAND2_X1 U8810 ( .A1(n7012), .A2(n10335), .ZN(n7013) );
  OAI21_X1 U8811 ( .B1(n10335), .B2(n6713), .A(n7013), .ZN(P1_U3475) );
  AOI21_X1 U8812 ( .B1(n9105), .B2(n7014), .A(n9122), .ZN(n7019) );
  AOI22_X1 U8813 ( .A1(n8819), .A2(n6045), .B1(n8821), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n7017) );
  INV_X1 U8814 ( .A(n7553), .ZN(n7015) );
  NAND2_X1 U8815 ( .A1(n9102), .A2(n7015), .ZN(n7016) );
  OAI211_X1 U8816 ( .C1(n7019), .C2(n7018), .A(n7017), .B(n7016), .ZN(P2_U3234) );
  NAND2_X1 U8817 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n9178), .ZN(n7020) );
  OAI21_X1 U8818 ( .B1(n9128), .B2(n9178), .A(n7020), .ZN(P2_U3577) );
  AOI211_X1 U8819 ( .C1(n7023), .C2(n7022), .A(n8921), .B(n7021), .ZN(n7033)
         );
  NAND2_X1 U8820 ( .A1(n7025), .A2(n7024), .ZN(n7026) );
  AOI21_X1 U8821 ( .B1(n7027), .B2(n7026), .A(n9295), .ZN(n7032) );
  NOR2_X1 U8822 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8742), .ZN(n7028) );
  AOI21_X1 U8823 ( .B1(n9289), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7028), .ZN(
        n7029) );
  OAI21_X1 U8824 ( .B1(n9286), .B2(n7030), .A(n7029), .ZN(n7031) );
  OR3_X1 U8825 ( .A1(n7033), .A2(n7032), .A3(n7031), .ZN(P2_U3257) );
  NOR2_X1 U8826 ( .A1(n7034), .A2(n8293), .ZN(n7035) );
  NAND2_X1 U8827 ( .A1(n7036), .A2(n7035), .ZN(n7040) );
  NOR2_X1 U8828 ( .A1(n6999), .A2(n9852), .ZN(n7037) );
  AOI21_X1 U8829 ( .B1(n7038), .B2(n7060), .A(n7037), .ZN(n7039) );
  NAND2_X1 U8830 ( .A1(n7040), .A2(n7039), .ZN(n7045) );
  NAND2_X1 U8831 ( .A1(n7041), .A2(n7910), .ZN(n7044) );
  AOI22_X1 U8832 ( .A1(n7873), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n4368), .B2(
        n7042), .ZN(n7043) );
  NAND2_X1 U8833 ( .A1(n7377), .A2(n7305), .ZN(n8306) );
  NAND2_X1 U8834 ( .A1(n7045), .A2(n8305), .ZN(n7046) );
  NAND2_X1 U8835 ( .A1(n7142), .A2(n7046), .ZN(n7067) );
  INV_X1 U8836 ( .A(n7067), .ZN(n7383) );
  OAI21_X1 U8837 ( .B1(n7047), .B2(n7290), .A(n7163), .ZN(n7379) );
  OAI22_X1 U8838 ( .A1(n7379), .A2(n10456), .B1(n7290), .B2(n10454), .ZN(n7068) );
  INV_X1 U8839 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n8684) );
  OR2_X1 U8840 ( .A1(n8187), .A2(n7161), .ZN(n7048) );
  OAI21_X1 U8841 ( .B1(n8190), .B2(n8684), .A(n7048), .ZN(n7049) );
  INV_X1 U8842 ( .A(n7049), .ZN(n7058) );
  INV_X1 U8843 ( .A(n7051), .ZN(n7151) );
  NAND2_X1 U8844 ( .A1(n7052), .A2(n8764), .ZN(n7053) );
  NAND2_X1 U8845 ( .A1(n7151), .A2(n7053), .ZN(n7302) );
  INV_X1 U8846 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7054) );
  OR2_X1 U8847 ( .A1(n8186), .A2(n7054), .ZN(n7055) );
  OAI21_X1 U8848 ( .B1(n7050), .B2(n7302), .A(n7055), .ZN(n7056) );
  INV_X1 U8849 ( .A(n7056), .ZN(n7057) );
  OAI22_X1 U8850 ( .A1(n7289), .A2(n10182), .B1(n10184), .B2(n7253), .ZN(n7059) );
  INV_X1 U8851 ( .A(n7059), .ZN(n7066) );
  NAND2_X1 U8852 ( .A1(n7062), .A2(n8258), .ZN(n7063) );
  NAND2_X1 U8853 ( .A1(n7063), .A2(n10117), .ZN(n7064) );
  OR2_X1 U8854 ( .A1(n7144), .A2(n7064), .ZN(n7065) );
  OAI211_X1 U8855 ( .C1(n7067), .C2(n7268), .A(n7066), .B(n7065), .ZN(n7380)
         );
  AOI211_X1 U8856 ( .C1(n10461), .C2(n7383), .A(n7068), .B(n7380), .ZN(n7071)
         );
  NAND2_X1 U8857 ( .A1(n10463), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7069) );
  OAI21_X1 U8858 ( .B1(n7071), .B2(n10463), .A(n7069), .ZN(P1_U3531) );
  NAND2_X1 U8859 ( .A1(n10462), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7070) );
  OAI21_X1 U8860 ( .B1(n7071), .B2(n10462), .A(n7070), .ZN(P1_U3478) );
  OR2_X1 U8861 ( .A1(n7072), .A2(n10462), .ZN(n7073) );
  OAI21_X1 U8862 ( .B1(n10335), .B2(n6632), .A(n7073), .ZN(P1_U3472) );
  OAI211_X1 U8863 ( .C1(n7076), .C2(n7075), .A(n9258), .B(n7074), .ZN(n7078)
         );
  NAND2_X1 U8864 ( .A1(P2_U3152), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7077) );
  OAI211_X1 U8865 ( .C1(n10359), .C2(n8927), .A(n7078), .B(n7077), .ZN(n7082)
         );
  AOI211_X1 U8866 ( .C1(n7080), .C2(n7079), .A(n9183), .B(n8921), .ZN(n7081)
         );
  AOI211_X1 U8867 ( .C1(n9263), .C2(n7083), .A(n7082), .B(n7081), .ZN(n7084)
         );
  INV_X1 U8868 ( .A(n7084), .ZN(P2_U3247) );
  OAI21_X1 U8869 ( .B1(n7087), .B2(n7086), .A(n7085), .ZN(n7093) );
  OAI22_X1 U8870 ( .A1(n9153), .A2(n10501), .B1(n7088), .B2(n9145), .ZN(n7092)
         );
  NAND2_X1 U8871 ( .A1(n8819), .A2(n9174), .ZN(n7089) );
  OAI211_X1 U8872 ( .C1(n9131), .C2(n7329), .A(n7090), .B(n7089), .ZN(n7091)
         );
  AOI211_X1 U8873 ( .C1(n7093), .C2(n9105), .A(n7092), .B(n7091), .ZN(n7094)
         );
  INV_X1 U8874 ( .A(n7094), .ZN(P2_U3241) );
  INV_X1 U8875 ( .A(n7885), .ZN(n7097) );
  AOI21_X1 U8876 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n9680), .A(n7095), .ZN(
        n7096) );
  OAI21_X1 U8877 ( .B1(n7097), .B2(n9684), .A(n7096), .ZN(P2_U3335) );
  XNOR2_X1 U8878 ( .A(n7099), .B(n7098), .ZN(n7105) );
  INV_X1 U8879 ( .A(n7480), .ZN(n7103) );
  OAI22_X1 U8880 ( .A1(n9148), .A2(n7717), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5200), .ZN(n7102) );
  OAI22_X1 U8881 ( .A1(n9153), .A2(n10508), .B1(n7100), .B2(n9145), .ZN(n7101)
         );
  AOI211_X1 U8882 ( .C1(n7103), .C2(n9143), .A(n7102), .B(n7101), .ZN(n7104)
         );
  OAI21_X1 U8883 ( .B1(n7105), .B2(n9138), .A(n7104), .ZN(P2_U3215) );
  NAND2_X1 U8884 ( .A1(n7885), .A2(n7106), .ZN(n7108) );
  NAND2_X1 U8885 ( .A1(n7107), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8444) );
  OAI211_X1 U8886 ( .C1(n7886), .C2(n10350), .A(n7108), .B(n8444), .ZN(
        P1_U3330) );
  XOR2_X1 U8887 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7489), .Z(n7111) );
  OAI21_X1 U8888 ( .B1(n7250), .B2(P1_REG1_REG_11__SCAN_IN), .A(n7109), .ZN(
        n7110) );
  OAI21_X1 U8889 ( .B1(n7111), .B2(n7110), .A(n7420), .ZN(n7112) );
  NOR2_X1 U8890 ( .A1(n7259), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7589) );
  AOI21_X1 U8891 ( .B1(n10427), .B2(n7112), .A(n7589), .ZN(n7113) );
  OAI21_X1 U8892 ( .B1(n7114), .B2(n10393), .A(n7113), .ZN(n7120) );
  NAND2_X1 U8893 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7489), .ZN(n7115) );
  OAI21_X1 U8894 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7489), .A(n7115), .ZN(
        n7118) );
  AOI211_X1 U8895 ( .C1(n7118), .C2(n7117), .A(n7426), .B(n10416), .ZN(n7119)
         );
  AOI211_X1 U8896 ( .C1(n10410), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n7120), .B(
        n7119), .ZN(n7121) );
  INV_X1 U8897 ( .A(n7121), .ZN(P1_U3253) );
  INV_X1 U8898 ( .A(n7122), .ZN(n10450) );
  AND2_X1 U8899 ( .A1(n7123), .A2(n10450), .ZN(n7388) );
  NAND2_X1 U8900 ( .A1(n7388), .A2(n7387), .ZN(n7124) );
  NAND2_X1 U8901 ( .A1(n7124), .A2(n10439), .ZN(n10011) );
  AND2_X1 U8902 ( .A1(n7125), .A2(n8112), .ZN(n7126) );
  NAND2_X1 U8903 ( .A1(n10139), .A2(n7126), .ZN(n10192) );
  MUX2_X1 U8904 ( .A(n7128), .B(n7127), .S(n10139), .Z(n7135) );
  AND2_X1 U8905 ( .A1(n10139), .A2(n10053), .ZN(n10071) );
  NAND2_X1 U8906 ( .A1(n10139), .A2(n7129), .ZN(n10433) );
  OAI22_X1 U8907 ( .A1(n10433), .A2(n7131), .B1(n10439), .B2(n7130), .ZN(n7132) );
  AOI21_X1 U8908 ( .B1(n10156), .B2(n7133), .A(n7132), .ZN(n7134) );
  OAI211_X1 U8909 ( .C1(n7136), .C2(n10192), .A(n7135), .B(n7134), .ZN(
        P1_U3287) );
  NAND2_X1 U8910 ( .A1(n7137), .A2(n7902), .ZN(n7140) );
  AOI22_X1 U8911 ( .A1(n7138), .A2(n4368), .B1(n7873), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n7139) );
  XNOR2_X1 U8912 ( .A(n10305), .B(n7253), .ZN(n8267) );
  NAND2_X1 U8913 ( .A1(n7377), .A2(n9851), .ZN(n7141) );
  XOR2_X1 U8914 ( .A(n8267), .B(n7247), .Z(n7160) );
  INV_X1 U8915 ( .A(n7160), .ZN(n10312) );
  INV_X2 U8916 ( .A(n10011), .ZN(n10437) );
  NOR3_X1 U8917 ( .A1(n10437), .A2(n7143), .A3(n10053), .ZN(n10163) );
  INV_X1 U8918 ( .A(n4484), .ZN(n7274) );
  XNOR2_X1 U8919 ( .A(n7254), .B(n8267), .ZN(n7158) );
  OR2_X1 U8920 ( .A1(n8187), .A2(n7145), .ZN(n7146) );
  OAI21_X1 U8921 ( .B1(n8190), .B2(n7147), .A(n7146), .ZN(n7148) );
  INV_X1 U8922 ( .A(n7148), .ZN(n7156) );
  INV_X1 U8923 ( .A(n7149), .ZN(n7232) );
  INV_X1 U8924 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7150) );
  NAND2_X1 U8925 ( .A1(n7151), .A2(n7150), .ZN(n7152) );
  NAND2_X1 U8926 ( .A1(n7232), .A2(n7152), .ZN(n7228) );
  INV_X1 U8927 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n8555) );
  OR2_X1 U8928 ( .A1(n8186), .A2(n8555), .ZN(n7153) );
  OAI21_X1 U8929 ( .B1(n7050), .B2(n7228), .A(n7153), .ZN(n7154) );
  INV_X1 U8930 ( .A(n7154), .ZN(n7155) );
  AOI22_X1 U8931 ( .A1(n10148), .A2(n9849), .B1(n10147), .B2(n9851), .ZN(n7157) );
  OAI21_X1 U8932 ( .B1(n7158), .B2(n10179), .A(n7157), .ZN(n7159) );
  AOI21_X1 U8933 ( .B1(n10153), .B2(n7160), .A(n7159), .ZN(n10310) );
  MUX2_X1 U8934 ( .A(n7161), .B(n10310), .S(n10139), .Z(n7167) );
  INV_X1 U8935 ( .A(n7464), .ZN(n7162) );
  AOI21_X1 U8936 ( .B1(n10305), .B2(n7163), .A(n7162), .ZN(n10308) );
  INV_X1 U8937 ( .A(n10305), .ZN(n7164) );
  OAI22_X1 U8938 ( .A1(n10433), .A2(n7164), .B1(n10439), .B2(n7302), .ZN(n7165) );
  AOI21_X1 U8939 ( .B1(n10308), .B2(n10156), .A(n7165), .ZN(n7166) );
  OAI211_X1 U8940 ( .C1(n10312), .C2(n7274), .A(n7167), .B(n7166), .ZN(
        P1_U3282) );
  INV_X1 U8941 ( .A(n10439), .ZN(n10170) );
  NOR2_X1 U8942 ( .A1(n7168), .A2(n9951), .ZN(n7170) );
  AOI211_X1 U8943 ( .C1(n10170), .C2(n7171), .A(n7170), .B(n7169), .ZN(n7172)
         );
  MUX2_X1 U8944 ( .A(n7173), .B(n7172), .S(n10139), .Z(n7176) );
  INV_X1 U8945 ( .A(n10433), .ZN(n9960) );
  NAND2_X1 U8946 ( .A1(n9960), .A2(n7174), .ZN(n7175) );
  OAI211_X1 U8947 ( .C1(n10192), .C2(n7177), .A(n7176), .B(n7175), .ZN(
        P1_U3286) );
  INV_X1 U8948 ( .A(n7605), .ZN(n7181) );
  AOI21_X1 U8949 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n7182), .A(n7604), .ZN(
        n7194) );
  NOR2_X1 U8950 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9147), .ZN(n7185) );
  NOR2_X1 U8951 ( .A1(n9286), .A2(n7183), .ZN(n7184) );
  AOI211_X1 U8952 ( .C1(n9289), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n7185), .B(
        n7184), .ZN(n7193) );
  NAND2_X1 U8953 ( .A1(n7187), .A2(n7186), .ZN(n7190) );
  NAND2_X1 U8954 ( .A1(n7188), .A2(n8744), .ZN(n7189) );
  NAND2_X1 U8955 ( .A1(n7190), .A2(n7189), .ZN(n7596) );
  XNOR2_X1 U8956 ( .A(n7596), .B(n7597), .ZN(n7191) );
  NAND2_X1 U8957 ( .A1(n7191), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n7600) );
  OAI211_X1 U8958 ( .C1(n7191), .C2(P2_REG1_REG_15__SCAN_IN), .A(n7600), .B(
        n9258), .ZN(n7192) );
  OAI211_X1 U8959 ( .C1(n7194), .C2(n8921), .A(n7193), .B(n7192), .ZN(P2_U3260) );
  AOI22_X1 U8960 ( .A1(n9960), .A2(n7195), .B1(n10437), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7201) );
  INV_X1 U8961 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7196) );
  OAI22_X1 U8962 ( .A1(n7197), .A2(n9951), .B1(n10439), .B2(n7196), .ZN(n7198)
         );
  OAI21_X1 U8963 ( .B1(n7199), .B2(n7198), .A(n10139), .ZN(n7200) );
  OAI211_X1 U8964 ( .C1(n10192), .C2(n7202), .A(n7201), .B(n7200), .ZN(
        P1_U3290) );
  NAND2_X1 U8965 ( .A1(n7203), .A2(n7902), .ZN(n7205) );
  AOI22_X1 U8966 ( .A1(n7873), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n4368), .B2(
        n10422), .ZN(n7204) );
  NAND2_X2 U8967 ( .A1(n7205), .A2(n7204), .ZN(n10301) );
  NAND2_X1 U8968 ( .A1(n10301), .A2(n8940), .ZN(n7207) );
  NAND2_X1 U8969 ( .A1(n9849), .A2(n4367), .ZN(n7206) );
  NAND2_X1 U8970 ( .A1(n7207), .A2(n7206), .ZN(n7208) );
  XNOR2_X1 U8971 ( .A(n7208), .B(n8112), .ZN(n7344) );
  NOR2_X1 U8972 ( .A1(n8154), .A2(n7362), .ZN(n7209) );
  AOI21_X1 U8973 ( .B1(n10301), .B2(n8934), .A(n7209), .ZN(n7345) );
  XNOR2_X1 U8974 ( .A(n7344), .B(n7345), .ZN(n7349) );
  OAI21_X2 U8975 ( .B1(n7212), .B2(n7211), .A(n7210), .ZN(n7283) );
  NAND2_X1 U8976 ( .A1(n10305), .A2(n8940), .ZN(n7214) );
  NAND2_X1 U8977 ( .A1(n9850), .A2(n8934), .ZN(n7213) );
  NAND2_X1 U8978 ( .A1(n7214), .A2(n7213), .ZN(n7215) );
  XNOR2_X1 U8979 ( .A(n7215), .B(n8112), .ZN(n7299) );
  NAND2_X1 U8980 ( .A1(n10305), .A2(n8934), .ZN(n7217) );
  NAND2_X1 U8981 ( .A1(n8935), .A2(n9850), .ZN(n7216) );
  NAND2_X1 U8982 ( .A1(n7217), .A2(n7216), .ZN(n7298) );
  NAND2_X1 U8983 ( .A1(n7377), .A2(n4367), .ZN(n7219) );
  NAND2_X1 U8984 ( .A1(n8935), .A2(n9851), .ZN(n7218) );
  NAND2_X1 U8985 ( .A1(n7219), .A2(n7218), .ZN(n7281) );
  NAND2_X1 U8986 ( .A1(n7377), .A2(n8940), .ZN(n7221) );
  NAND2_X1 U8987 ( .A1(n9851), .A2(n8934), .ZN(n7220) );
  NAND2_X1 U8988 ( .A1(n7221), .A2(n7220), .ZN(n7222) );
  XNOR2_X1 U8989 ( .A(n7222), .B(n8112), .ZN(n7297) );
  AOI22_X1 U8990 ( .A1(n7299), .A2(n7298), .B1(n7281), .B2(n7297), .ZN(n7223)
         );
  INV_X1 U8991 ( .A(n7299), .ZN(n7226) );
  OAI21_X1 U8992 ( .B1(n7297), .B2(n7281), .A(n7298), .ZN(n7225) );
  NOR2_X1 U8993 ( .A1(n7298), .A2(n7281), .ZN(n7224) );
  INV_X1 U8994 ( .A(n7297), .ZN(n7285) );
  AOI22_X1 U8995 ( .A1(n7226), .A2(n7225), .B1(n7224), .B2(n7285), .ZN(n7347)
         );
  NAND2_X1 U8996 ( .A1(n7352), .A2(n7347), .ZN(n7227) );
  XOR2_X1 U8997 ( .A(n7349), .B(n7227), .Z(n7241) );
  INV_X1 U8998 ( .A(n7228), .ZN(n7465) );
  INV_X1 U8999 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n8733) );
  OR2_X1 U9000 ( .A1(n8186), .A2(n8733), .ZN(n7230) );
  OR2_X1 U9001 ( .A1(n8187), .A2(n8579), .ZN(n7229) );
  AND2_X1 U9002 ( .A1(n7230), .A2(n7229), .ZN(n7236) );
  INV_X1 U9003 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7231) );
  NAND2_X1 U9004 ( .A1(n7232), .A2(n7231), .ZN(n7233) );
  AND2_X1 U9005 ( .A1(n7260), .A2(n7233), .ZN(n7364) );
  NAND2_X1 U9006 ( .A1(n8184), .A2(n7364), .ZN(n7235) );
  NAND2_X1 U9007 ( .A1(n4379), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7234) );
  NAND2_X1 U9008 ( .A1(n9835), .A2(n9848), .ZN(n7237) );
  NAND2_X1 U9009 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10415) );
  OAI211_X1 U9010 ( .C1(n7253), .C2(n9831), .A(n7237), .B(n10415), .ZN(n7238)
         );
  AOI21_X1 U9011 ( .B1(n7465), .B2(n9773), .A(n7238), .ZN(n7240) );
  NAND2_X1 U9012 ( .A1(n4582), .A2(n10301), .ZN(n7239) );
  OAI211_X1 U9013 ( .C1(n7241), .C2(n9825), .A(n7240), .B(n7239), .ZN(P1_U3215) );
  INV_X1 U9014 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7242) );
  OAI22_X1 U9015 ( .A1(n9670), .A2(n7415), .B1(n10513), .B2(n7242), .ZN(n7243)
         );
  INV_X1 U9016 ( .A(n7243), .ZN(n7244) );
  OAI21_X1 U9017 ( .B1(n7245), .B2(n10512), .A(n7244), .ZN(P2_U3460) );
  AND2_X1 U9018 ( .A1(n10305), .A2(n9850), .ZN(n7246) );
  NAND2_X1 U9019 ( .A1(n10301), .A2(n7362), .ZN(n8317) );
  NAND2_X1 U9020 ( .A1(n8205), .A2(n8317), .ZN(n8313) );
  NOR2_X1 U9021 ( .A1(n10301), .A2(n9849), .ZN(n7248) );
  NAND2_X1 U9022 ( .A1(n7249), .A2(n7902), .ZN(n7252) );
  AOI22_X1 U9023 ( .A1(n7873), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n4368), .B2(
        n7250), .ZN(n7251) );
  XNOR2_X1 U9024 ( .A(n7507), .B(n7506), .ZN(n8321) );
  XNOR2_X1 U9025 ( .A(n7510), .B(n8321), .ZN(n7568) );
  NOR2_X1 U9026 ( .A1(n10305), .A2(n7253), .ZN(n8310) );
  INV_X1 U9027 ( .A(n8310), .ZN(n8228) );
  AND2_X1 U9028 ( .A1(n10305), .A2(n7253), .ZN(n8311) );
  INV_X1 U9029 ( .A(n8321), .ZN(n8271) );
  XNOR2_X1 U9030 ( .A(n7486), .B(n8271), .ZN(n7266) );
  INV_X1 U9031 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7255) );
  OR2_X1 U9032 ( .A1(n8187), .A2(n7255), .ZN(n7258) );
  INV_X1 U9033 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7256) );
  OR2_X1 U9034 ( .A1(n8186), .A2(n7256), .ZN(n7257) );
  AND2_X1 U9035 ( .A1(n7258), .A2(n7257), .ZN(n7264) );
  NAND2_X1 U9036 ( .A1(n7260), .A2(n7259), .ZN(n7261) );
  AND2_X1 U9037 ( .A1(n7494), .A2(n7261), .ZN(n7590) );
  NAND2_X1 U9038 ( .A1(n8184), .A2(n7590), .ZN(n7263) );
  NAND2_X1 U9039 ( .A1(n4379), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7262) );
  OAI22_X1 U9040 ( .A1(n7628), .A2(n10184), .B1(n10182), .B2(n7362), .ZN(n7265) );
  AOI21_X1 U9041 ( .B1(n7266), .B2(n10117), .A(n7265), .ZN(n7267) );
  OAI21_X1 U9042 ( .B1(n7268), .B2(n7568), .A(n7267), .ZN(n7571) );
  NAND2_X1 U9043 ( .A1(n7571), .A2(n10011), .ZN(n7273) );
  INV_X1 U9044 ( .A(n7364), .ZN(n7269) );
  OAI22_X1 U9045 ( .A1(n10139), .A2(n8579), .B1(n7269), .B2(n10439), .ZN(n7271) );
  OAI21_X1 U9046 ( .B1(n4467), .B2(n7569), .A(n7504), .ZN(n7570) );
  INV_X1 U9047 ( .A(n10156), .ZN(n10434) );
  NOR2_X1 U9048 ( .A1(n7570), .A2(n10434), .ZN(n7270) );
  AOI211_X1 U9049 ( .C1(n9960), .C2(n7507), .A(n7271), .B(n7270), .ZN(n7272)
         );
  OAI211_X1 U9050 ( .C1(n7568), .C2(n7274), .A(n7273), .B(n7272), .ZN(P1_U3280) );
  XNOR2_X1 U9051 ( .A(n7276), .B(n7275), .ZN(n7280) );
  NAND2_X1 U9052 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n9224) );
  OAI21_X1 U9053 ( .B1(n9148), .B2(n7671), .A(n9224), .ZN(n7278) );
  OAI22_X1 U9054 ( .A1(n9131), .A2(n7453), .B1(n7439), .B2(n9145), .ZN(n7277)
         );
  AOI211_X1 U9055 ( .C1(n7449), .C2(n9122), .A(n7278), .B(n7277), .ZN(n7279)
         );
  OAI21_X1 U9056 ( .B1(n7280), .B2(n9138), .A(n7279), .ZN(P2_U3223) );
  INV_X1 U9057 ( .A(n7281), .ZN(n7282) );
  NOR2_X1 U9058 ( .A1(n7283), .A2(n7282), .ZN(n7295) );
  INV_X1 U9059 ( .A(n7295), .ZN(n7284) );
  NAND2_X1 U9060 ( .A1(n7283), .A2(n7282), .ZN(n7296) );
  NAND2_X1 U9061 ( .A1(n7284), .A2(n7296), .ZN(n7286) );
  XNOR2_X1 U9062 ( .A(n7286), .B(n7285), .ZN(n7294) );
  NAND2_X1 U9063 ( .A1(n9835), .A2(n9850), .ZN(n7288) );
  OAI211_X1 U9064 ( .C1(n7289), .C2(n9831), .A(n7288), .B(n7287), .ZN(n7292)
         );
  NOR2_X1 U9065 ( .A1(n9838), .A2(n7290), .ZN(n7291) );
  AOI211_X1 U9066 ( .C1(n7376), .C2(n9773), .A(n7292), .B(n7291), .ZN(n7293)
         );
  OAI21_X1 U9067 ( .B1(n7294), .B2(n9825), .A(n7293), .ZN(P1_U3219) );
  AOI21_X1 U9068 ( .B1(n7297), .B2(n7296), .A(n7295), .ZN(n7301) );
  XNOR2_X1 U9069 ( .A(n7299), .B(n7298), .ZN(n7300) );
  XNOR2_X1 U9070 ( .A(n7301), .B(n7300), .ZN(n7310) );
  INV_X1 U9071 ( .A(n7302), .ZN(n7307) );
  NAND2_X1 U9072 ( .A1(n9835), .A2(n9849), .ZN(n7304) );
  OAI211_X1 U9073 ( .C1(n7305), .C2(n9831), .A(n7304), .B(n7303), .ZN(n7306)
         );
  AOI21_X1 U9074 ( .B1(n7307), .B2(n9773), .A(n7306), .ZN(n7309) );
  NAND2_X1 U9075 ( .A1(n4582), .A2(n10305), .ZN(n7308) );
  OAI211_X1 U9076 ( .C1(n7310), .C2(n9825), .A(n7309), .B(n7308), .ZN(P1_U3229) );
  INV_X1 U9077 ( .A(n7314), .ZN(n7311) );
  NAND2_X1 U9078 ( .A1(n7311), .A2(n7312), .ZN(n7327) );
  NAND2_X2 U9079 ( .A1(n7327), .A2(n9485), .ZN(n9536) );
  NAND2_X1 U9080 ( .A1(n8880), .A2(n7312), .ZN(n7313) );
  NOR2_X1 U9081 ( .A1(n7314), .A2(n7313), .ZN(n7679) );
  INV_X1 U9082 ( .A(n7679), .ZN(n8828) );
  OAI22_X1 U9083 ( .A1(n8828), .A2(n7315), .B1(n8753), .B2(n9485), .ZN(n7316)
         );
  AOI21_X1 U9084 ( .B1(n9536), .B2(n7317), .A(n7316), .ZN(n7325) );
  INV_X1 U9085 ( .A(n7318), .ZN(n7319) );
  NAND2_X1 U9086 ( .A1(n7319), .A2(n9359), .ZN(n7410) );
  NAND2_X1 U9087 ( .A1(n7741), .A2(n7410), .ZN(n7320) );
  AOI22_X1 U9088 ( .A1(n9522), .A2(n7323), .B1(n9521), .B2(n7322), .ZN(n7324)
         );
  OAI211_X1 U9089 ( .C1(n6754), .C2(n9536), .A(n7325), .B(n7324), .ZN(P2_U3294) );
  XOR2_X1 U9090 ( .A(n7331), .B(n7326), .Z(n10504) );
  INV_X1 U9091 ( .A(n10504), .ZN(n7339) );
  INV_X1 U9092 ( .A(n7327), .ZN(n7328) );
  NAND2_X1 U9093 ( .A1(n7328), .A2(n8923), .ZN(n9491) );
  OAI211_X1 U9094 ( .C1(n7531), .C2(n10501), .A(n9484), .B(n7472), .ZN(n10500)
         );
  OAI22_X1 U9095 ( .A1(n9491), .A2(n10500), .B1(n7329), .B2(n9485), .ZN(n7336)
         );
  OAI21_X1 U9096 ( .B1(n7331), .B2(n7330), .A(n7476), .ZN(n7332) );
  NAND2_X1 U9097 ( .A1(n7332), .A2(n9524), .ZN(n7334) );
  NAND2_X1 U9098 ( .A1(n7334), .A2(n7333), .ZN(n10503) );
  MUX2_X1 U9099 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10503), .S(n9536), .Z(n7335)
         );
  AOI211_X1 U9100 ( .C1(n9521), .C2(n7337), .A(n7336), .B(n7335), .ZN(n7338)
         );
  OAI21_X1 U9101 ( .B1(n7339), .B2(n9495), .A(n7338), .ZN(P2_U3290) );
  INV_X1 U9102 ( .A(n7889), .ZN(n7342) );
  OAI222_X1 U9103 ( .A1(n7340), .A2(P1_U3084), .B1(n10347), .B2(n7342), .C1(
        n7890), .C2(n10350), .ZN(P1_U3329) );
  OAI222_X1 U9104 ( .A1(P2_U3152), .A2(n7343), .B1(n9684), .B2(n7342), .C1(
        n7341), .C2(n9686), .ZN(P2_U3334) );
  INV_X1 U9105 ( .A(n7344), .ZN(n7346) );
  NAND2_X1 U9106 ( .A1(n7346), .A2(n7345), .ZN(n7348) );
  AND2_X1 U9107 ( .A1(n7347), .A2(n7348), .ZN(n7351) );
  INV_X1 U9108 ( .A(n7348), .ZN(n7350) );
  NAND2_X1 U9109 ( .A1(n7507), .A2(n8940), .ZN(n7354) );
  NAND2_X1 U9110 ( .A1(n9848), .A2(n4367), .ZN(n7353) );
  NAND2_X1 U9111 ( .A1(n7354), .A2(n7353), .ZN(n7355) );
  XNOR2_X1 U9112 ( .A(n7355), .B(n8938), .ZN(n7581) );
  NOR2_X1 U9113 ( .A1(n8154), .A2(n7506), .ZN(n7356) );
  AOI21_X1 U9114 ( .B1(n7507), .B2(n4367), .A(n7356), .ZN(n7580) );
  XNOR2_X1 U9115 ( .A(n7581), .B(n7580), .ZN(n7357) );
  AOI21_X1 U9116 ( .B1(n7358), .B2(n7357), .A(n9825), .ZN(n7359) );
  NAND2_X1 U9117 ( .A1(n7359), .A2(n7582), .ZN(n7366) );
  NAND2_X1 U9118 ( .A1(n9835), .A2(n9847), .ZN(n7361) );
  OAI211_X1 U9119 ( .C1(n7362), .C2(n9831), .A(n7361), .B(n7360), .ZN(n7363)
         );
  AOI21_X1 U9120 ( .B1(n7364), .B2(n9773), .A(n7363), .ZN(n7365) );
  OAI211_X1 U9121 ( .C1(n7569), .C2(n9838), .A(n7366), .B(n7365), .ZN(P1_U3234) );
  AOI22_X1 U9122 ( .A1(n9960), .A2(n7368), .B1(n10170), .B2(n7367), .ZN(n7369)
         );
  OAI21_X1 U9123 ( .B1(n10434), .B2(n7370), .A(n7369), .ZN(n7373) );
  MUX2_X1 U9124 ( .A(n7371), .B(P1_REG2_REG_6__SCAN_IN), .S(n10437), .Z(n7372)
         );
  AOI211_X1 U9125 ( .C1(n7374), .C2(n4484), .A(n7373), .B(n7372), .ZN(n7375)
         );
  INV_X1 U9126 ( .A(n7375), .ZN(P1_U3285) );
  AOI22_X1 U9127 ( .A1(n9960), .A2(n7377), .B1(n10170), .B2(n7376), .ZN(n7378)
         );
  OAI21_X1 U9128 ( .B1(n7379), .B2(n10434), .A(n7378), .ZN(n7382) );
  MUX2_X1 U9129 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n7380), .S(n10139), .Z(n7381)
         );
  AOI211_X1 U9130 ( .C1(n7383), .C2(n4484), .A(n7382), .B(n7381), .ZN(n7384)
         );
  INV_X1 U9131 ( .A(n7384), .ZN(P1_U3283) );
  AOI21_X1 U9132 ( .B1(n7386), .B2(n10170), .A(n7385), .ZN(n7395) );
  AND3_X1 U9133 ( .A1(n7388), .A2(n7387), .A3(n10053), .ZN(n10190) );
  INV_X1 U9134 ( .A(n6999), .ZN(n7389) );
  OAI22_X1 U9135 ( .A1(n10433), .A2(n7389), .B1(n10402), .B2(n10139), .ZN(
        n7392) );
  NOR2_X1 U9136 ( .A1(n7390), .A2(n10192), .ZN(n7391) );
  AOI211_X1 U9137 ( .C1(n7393), .C2(n10190), .A(n7392), .B(n7391), .ZN(n7394)
         );
  OAI21_X1 U9138 ( .B1(n10437), .B2(n7395), .A(n7394), .ZN(P1_U3284) );
  OAI21_X1 U9139 ( .B1(n7397), .B2(n7401), .A(n7396), .ZN(n10460) );
  OAI21_X1 U9140 ( .B1(n10455), .B2(n4404), .A(n4482), .ZN(n10457) );
  AOI22_X1 U9141 ( .A1(n9960), .A2(n7399), .B1(n10170), .B2(n7398), .ZN(n7400)
         );
  OAI21_X1 U9142 ( .B1(n10434), .B2(n10457), .A(n7400), .ZN(n7408) );
  XNOR2_X1 U9143 ( .A(n7401), .B(n8408), .ZN(n7406) );
  NAND2_X1 U9144 ( .A1(n10460), .A2(n10153), .ZN(n7405) );
  OAI22_X1 U9145 ( .A1(n8218), .A2(n10182), .B1(n10184), .B2(n7402), .ZN(n7403) );
  INV_X1 U9146 ( .A(n7403), .ZN(n7404) );
  OAI211_X1 U9147 ( .C1(n10179), .C2(n7406), .A(n7405), .B(n7404), .ZN(n10458)
         );
  MUX2_X1 U9148 ( .A(n10458), .B(P1_REG2_REG_3__SCAN_IN), .S(n10437), .Z(n7407) );
  INV_X1 U9149 ( .A(n7409), .ZN(P1_U3288) );
  INV_X1 U9150 ( .A(n7410), .ZN(n7411) );
  NAND2_X1 U9151 ( .A1(n9536), .A2(n7411), .ZN(n7756) );
  INV_X1 U9152 ( .A(n7756), .ZN(n7455) );
  MUX2_X1 U9153 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7412), .S(n9536), .Z(n7417)
         );
  INV_X1 U9154 ( .A(n9485), .ZN(n9535) );
  AOI22_X1 U9155 ( .A1(n9540), .A2(n7413), .B1(n9535), .B2(n9180), .ZN(n7414)
         );
  OAI21_X1 U9156 ( .B1(n9437), .B2(n7415), .A(n7414), .ZN(n7416) );
  AOI211_X1 U9157 ( .C1(n7455), .C2(n7418), .A(n7417), .B(n7416), .ZN(n7419)
         );
  INV_X1 U9158 ( .A(n7419), .ZN(P2_U3293) );
  XOR2_X1 U9159 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9864), .Z(n7422) );
  OAI21_X1 U9160 ( .B1(n7422), .B2(n7421), .A(n9860), .ZN(n7423) );
  NOR2_X1 U9161 ( .A1(n7493), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7657) );
  AOI21_X1 U9162 ( .B1(n10427), .B2(n7423), .A(n7657), .ZN(n7424) );
  OAI21_X1 U9163 ( .B1(n7425), .B2(n10393), .A(n7424), .ZN(n7430) );
  NAND2_X1 U9164 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n9864), .ZN(n7427) );
  OAI21_X1 U9165 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9864), .A(n7427), .ZN(
        n7428) );
  AOI211_X1 U9166 ( .C1(n4476), .C2(n7428), .A(n9866), .B(n10416), .ZN(n7429)
         );
  AOI211_X1 U9167 ( .C1(n10410), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n7430), .B(
        n7429), .ZN(n7431) );
  INV_X1 U9168 ( .A(n7431), .ZN(P1_U3254) );
  NOR2_X1 U9169 ( .A1(n7664), .A2(n5248), .ZN(n7712) );
  AND2_X1 U9170 ( .A1(n7664), .A2(n5248), .ZN(n7432) );
  OR2_X1 U9171 ( .A1(n7712), .A2(n7432), .ZN(n7443) );
  INV_X1 U9172 ( .A(n7443), .ZN(n7456) );
  NAND2_X1 U9173 ( .A1(n7473), .A2(n7449), .ZN(n7433) );
  NAND2_X1 U9174 ( .A1(n7433), .A2(n9484), .ZN(n7434) );
  NOR2_X1 U9175 ( .A1(n7722), .A2(n7434), .ZN(n7450) );
  NAND2_X1 U9176 ( .A1(n7436), .A2(n7435), .ZN(n7437) );
  NAND2_X1 U9177 ( .A1(n7438), .A2(n7437), .ZN(n7441) );
  OAI22_X1 U9178 ( .A1(n9531), .A2(n7439), .B1(n7671), .B2(n9528), .ZN(n7440)
         );
  AOI21_X1 U9179 ( .B1(n7441), .B2(n9524), .A(n7440), .ZN(n7442) );
  OAI21_X1 U9180 ( .B1(n7443), .B2(n7741), .A(n7442), .ZN(n7447) );
  AOI211_X1 U9181 ( .C1(n7456), .C2(n7735), .A(n7450), .B(n7447), .ZN(n7446)
         );
  AOI22_X1 U9182 ( .A1(n5975), .A2(n7449), .B1(n10512), .B2(
        P2_REG0_REG_8__SCAN_IN), .ZN(n7444) );
  OAI21_X1 U9183 ( .B1(n7446), .B2(n10512), .A(n7444), .ZN(P2_U3475) );
  INV_X1 U9184 ( .A(n9615), .ZN(n7701) );
  AOI22_X1 U9185 ( .A1(n7701), .A2(n7449), .B1(P2_REG1_REG_8__SCAN_IN), .B2(
        n10519), .ZN(n7445) );
  OAI21_X1 U9186 ( .B1(n7446), .B2(n10519), .A(n7445), .ZN(P2_U3528) );
  MUX2_X1 U9187 ( .A(n7447), .B(P2_REG2_REG_8__SCAN_IN), .S(n4374), .Z(n7448)
         );
  INV_X1 U9188 ( .A(n7448), .ZN(n7458) );
  NAND2_X1 U9189 ( .A1(n9521), .A2(n7449), .ZN(n7452) );
  NAND2_X1 U9190 ( .A1(n9540), .A2(n7450), .ZN(n7451) );
  OAI211_X1 U9191 ( .C1(n9485), .C2(n7453), .A(n7452), .B(n7451), .ZN(n7454)
         );
  AOI21_X1 U9192 ( .B1(n7456), .B2(n7455), .A(n7454), .ZN(n7457) );
  NAND2_X1 U9193 ( .A1(n7458), .A2(n7457), .ZN(P2_U3288) );
  XNOR2_X1 U9194 ( .A(n7459), .B(n8313), .ZN(n10299) );
  XOR2_X1 U9195 ( .A(n7460), .B(n8313), .Z(n7462) );
  AOI22_X1 U9196 ( .A1(n10148), .A2(n9848), .B1(n10147), .B2(n9850), .ZN(n7461) );
  OAI21_X1 U9197 ( .B1(n7462), .B2(n10179), .A(n7461), .ZN(n7463) );
  AOI21_X1 U9198 ( .B1(n10153), .B2(n10299), .A(n7463), .ZN(n10303) );
  INV_X1 U9199 ( .A(n10301), .ZN(n7468) );
  AOI211_X1 U9200 ( .C1(n10301), .C2(n7464), .A(n10456), .B(n4467), .ZN(n10300) );
  NAND2_X1 U9201 ( .A1(n10300), .A2(n10190), .ZN(n7467) );
  AOI22_X1 U9202 ( .A1(n10437), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7465), .B2(
        n10170), .ZN(n7466) );
  OAI211_X1 U9203 ( .C1(n7468), .C2(n10433), .A(n7467), .B(n7466), .ZN(n7469)
         );
  AOI21_X1 U9204 ( .B1(n4484), .B2(n10299), .A(n7469), .ZN(n7470) );
  OAI21_X1 U9205 ( .B1(n10303), .B2(n10437), .A(n7470), .ZN(P1_U3281) );
  XNOR2_X1 U9206 ( .A(n7471), .B(n7477), .ZN(n10511) );
  OAI211_X1 U9207 ( .C1(n7474), .C2(n10508), .A(n9484), .B(n7473), .ZN(n10505)
         );
  OAI22_X1 U9208 ( .A1(n9437), .A2(n10508), .B1(n10505), .B2(n9491), .ZN(n7483) );
  NAND2_X1 U9209 ( .A1(n7476), .A2(n7475), .ZN(n7478) );
  XNOR2_X1 U9210 ( .A(n7478), .B(n7477), .ZN(n7479) );
  AOI222_X1 U9211 ( .A1(n9524), .A2(n7479), .B1(n9175), .B2(n9462), .C1(n9173), 
        .C2(n9464), .ZN(n10506) );
  OAI21_X1 U9212 ( .B1(n7480), .B2(n9485), .A(n10506), .ZN(n7481) );
  MUX2_X1 U9213 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7481), .S(n9536), .Z(n7482)
         );
  AOI211_X1 U9214 ( .C1(n9522), .C2(n10511), .A(n7483), .B(n7482), .ZN(n7484)
         );
  INV_X1 U9215 ( .A(n7484), .ZN(P2_U3289) );
  NAND2_X1 U9216 ( .A1(n7507), .A2(n7506), .ZN(n8204) );
  INV_X1 U9217 ( .A(n8204), .ZN(n7485) );
  OR2_X1 U9218 ( .A1(n7507), .A2(n7506), .ZN(n7629) );
  INV_X1 U9219 ( .A(n7629), .ZN(n7487) );
  NOR2_X1 U9220 ( .A1(n7631), .A2(n7487), .ZN(n7492) );
  NAND2_X1 U9221 ( .A1(n7488), .A2(n7910), .ZN(n7491) );
  AOI22_X1 U9222 ( .A1(n7873), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n4368), .B2(
        n7489), .ZN(n7490) );
  NAND2_X2 U9223 ( .A1(n7491), .A2(n7490), .ZN(n10294) );
  INV_X1 U9224 ( .A(n10294), .ZN(n7614) );
  NAND2_X1 U9225 ( .A1(n7630), .A2(n8318), .ZN(n8270) );
  XNOR2_X1 U9226 ( .A(n7492), .B(n7615), .ZN(n7503) );
  NAND2_X1 U9227 ( .A1(n7494), .A2(n7493), .ZN(n7495) );
  AND2_X1 U9228 ( .A1(n7622), .A2(n7495), .ZN(n7658) );
  NAND2_X1 U9229 ( .A1(n7658), .A2(n8184), .ZN(n7502) );
  INV_X1 U9230 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7496) );
  OR2_X1 U9231 ( .A1(n8186), .A2(n7496), .ZN(n7499) );
  INV_X1 U9232 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7497) );
  OR2_X1 U9233 ( .A1(n8187), .A2(n7497), .ZN(n7498) );
  AND2_X1 U9234 ( .A1(n7499), .A2(n7498), .ZN(n7501) );
  NAND2_X1 U9235 ( .A1(n4379), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7500) );
  AOI222_X1 U9236 ( .A1(n10117), .A2(n7503), .B1(n9846), .B2(n10148), .C1(
        n9848), .C2(n10147), .ZN(n10296) );
  AOI22_X1 U9237 ( .A1(n10437), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7590), .B2(
        n10170), .ZN(n7505) );
  OAI21_X1 U9238 ( .B1(n7614), .B2(n10433), .A(n7505), .ZN(n7512) );
  NAND2_X1 U9239 ( .A1(n7569), .A2(n7506), .ZN(n7509) );
  XNOR2_X1 U9240 ( .A(n7616), .B(n7615), .ZN(n10297) );
  NOR2_X1 U9241 ( .A1(n10297), .A2(n10192), .ZN(n7511) );
  AOI211_X1 U9242 ( .C1(n10293), .C2(n10190), .A(n7512), .B(n7511), .ZN(n7513)
         );
  OAI21_X1 U9243 ( .B1(n10296), .B2(n10437), .A(n7513), .ZN(P1_U3279) );
  INV_X1 U9244 ( .A(n7514), .ZN(n7516) );
  NOR2_X1 U9245 ( .A1(n7516), .A2(n7515), .ZN(n7517) );
  XNOR2_X1 U9246 ( .A(n7518), .B(n7517), .ZN(n7524) );
  INV_X1 U9247 ( .A(n7724), .ZN(n7522) );
  NOR2_X1 U9248 ( .A1(n5259), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9243) );
  INV_X1 U9249 ( .A(n9243), .ZN(n7519) );
  OAI21_X1 U9250 ( .B1(n9148), .B2(n7785), .A(n7519), .ZN(n7521) );
  OAI22_X1 U9251 ( .A1(n9153), .A2(n7725), .B1(n7717), .B2(n9145), .ZN(n7520)
         );
  AOI211_X1 U9252 ( .C1(n7522), .C2(n9143), .A(n7521), .B(n7520), .ZN(n7523)
         );
  OAI21_X1 U9253 ( .B1(n7524), .B2(n9138), .A(n7523), .ZN(P2_U3233) );
  NAND2_X1 U9254 ( .A1(n7526), .A2(n7525), .ZN(n7527) );
  XNOR2_X1 U9255 ( .A(n7527), .B(n7536), .ZN(n7529) );
  AOI21_X1 U9256 ( .B1(n7529), .B2(n9524), .A(n7528), .ZN(n10495) );
  OAI21_X1 U9257 ( .B1(n7530), .B2(n10496), .A(n9484), .ZN(n7532) );
  NOR2_X1 U9258 ( .A1(n7532), .A2(n7531), .ZN(n10493) );
  NAND2_X1 U9259 ( .A1(n9536), .A2(n8923), .ZN(n9515) );
  INV_X1 U9260 ( .A(n9515), .ZN(n9469) );
  OAI22_X1 U9261 ( .A1(n9536), .A2(n6757), .B1(n7533), .B2(n9485), .ZN(n7535)
         );
  NOR2_X1 U9262 ( .A1(n9437), .A2(n10496), .ZN(n7534) );
  AOI211_X1 U9263 ( .C1(n10493), .C2(n9469), .A(n7535), .B(n7534), .ZN(n7539)
         );
  XNOR2_X1 U9264 ( .A(n7537), .B(n7536), .ZN(n10498) );
  NAND2_X1 U9265 ( .A1(n9522), .A2(n10498), .ZN(n7538) );
  OAI211_X1 U9266 ( .C1(n4374), .C2(n10495), .A(n7539), .B(n7538), .ZN(
        P2_U3291) );
  NAND2_X1 U9267 ( .A1(n7541), .A2(n7540), .ZN(n7542) );
  XNOR2_X1 U9268 ( .A(n7542), .B(n7546), .ZN(n7544) );
  OAI22_X1 U9269 ( .A1(n9531), .A2(n9014), .B1(n8975), .B2(n9528), .ZN(n9018)
         );
  INV_X1 U9270 ( .A(n9018), .ZN(n7543) );
  OAI21_X1 U9271 ( .B1(n7544), .B2(n9442), .A(n7543), .ZN(n7696) );
  INV_X1 U9272 ( .A(n7696), .ZN(n7552) );
  XNOR2_X1 U9273 ( .A(n7545), .B(n7546), .ZN(n7698) );
  AOI211_X1 U9274 ( .C1(n7700), .C2(n7690), .A(n9538), .B(n7750), .ZN(n7697)
         );
  NAND2_X1 U9275 ( .A1(n7697), .A2(n9540), .ZN(n7549) );
  INV_X1 U9276 ( .A(n7547), .ZN(n9020) );
  AOI22_X1 U9277 ( .A1(n4374), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n9020), .B2(
        n9535), .ZN(n7548) );
  OAI211_X1 U9278 ( .C1(n9019), .C2(n9437), .A(n7549), .B(n7548), .ZN(n7550)
         );
  AOI21_X1 U9279 ( .B1(n9522), .B2(n7698), .A(n7550), .ZN(n7551) );
  OAI21_X1 U9280 ( .B1(n4374), .B2(n7552), .A(n7551), .ZN(P2_U3284) );
  NAND2_X1 U9281 ( .A1(n7554), .A2(n7553), .ZN(n10483) );
  INV_X1 U9282 ( .A(n10483), .ZN(n7559) );
  AOI22_X1 U9283 ( .A1(n10483), .A2(n9524), .B1(n9464), .B2(n6045), .ZN(n10485) );
  OAI22_X1 U9284 ( .A1(n4374), .A2(n10485), .B1(n7555), .B2(n9485), .ZN(n7556)
         );
  AOI21_X1 U9285 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n4374), .A(n7556), .ZN(
        n7558) );
  OAI21_X1 U9286 ( .B1(n9521), .B2(n7679), .A(n10481), .ZN(n7557) );
  OAI211_X1 U9287 ( .C1(n7559), .C2(n9495), .A(n7558), .B(n7557), .ZN(P2_U3296) );
  NAND2_X1 U9288 ( .A1(n10156), .A2(n7560), .ZN(n7562) );
  AOI22_X1 U9289 ( .A1(n10437), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10170), .ZN(n7561) );
  OAI211_X1 U9290 ( .C1(n7563), .C2(n10433), .A(n7562), .B(n7561), .ZN(n7564)
         );
  AOI21_X1 U9291 ( .B1(n4484), .B2(n7565), .A(n7564), .ZN(n7566) );
  OAI21_X1 U9292 ( .B1(n7567), .B2(n10437), .A(n7566), .ZN(P1_U3289) );
  INV_X1 U9293 ( .A(n7568), .ZN(n7573) );
  OAI22_X1 U9294 ( .A1(n7570), .A2(n10456), .B1(n7569), .B2(n10454), .ZN(n7572) );
  AOI211_X1 U9295 ( .C1(n10461), .C2(n7573), .A(n7572), .B(n7571), .ZN(n7576)
         );
  NAND2_X1 U9296 ( .A1(n10463), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7574) );
  OAI21_X1 U9297 ( .B1(n7576), .B2(n10463), .A(n7574), .ZN(P1_U3534) );
  NAND2_X1 U9298 ( .A1(n10462), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7575) );
  OAI21_X1 U9299 ( .B1(n7576), .B2(n10462), .A(n7575), .ZN(P1_U3487) );
  INV_X1 U9300 ( .A(n7894), .ZN(n7579) );
  OAI222_X1 U9301 ( .A1(n9686), .A2(n7578), .B1(n8964), .B2(n7579), .C1(
        P2_U3152), .C2(n7577), .ZN(P2_U3333) );
  OAI222_X1 U9302 ( .A1(n10350), .A2(n7895), .B1(n10347), .B2(n7579), .C1(
        n6328), .C2(P1_U3084), .ZN(P1_U3328) );
  NAND2_X1 U9303 ( .A1(n10294), .A2(n8940), .ZN(n7584) );
  NAND2_X1 U9304 ( .A1(n9847), .A2(n8934), .ZN(n7583) );
  NAND2_X1 U9305 ( .A1(n7584), .A2(n7583), .ZN(n7585) );
  XNOR2_X1 U9306 ( .A(n7585), .B(n8112), .ZN(n7644) );
  NAND2_X1 U9307 ( .A1(n10294), .A2(n4367), .ZN(n7587) );
  NAND2_X1 U9308 ( .A1(n8935), .A2(n9847), .ZN(n7586) );
  NAND2_X1 U9309 ( .A1(n7587), .A2(n7586), .ZN(n7643) );
  INV_X1 U9310 ( .A(n7643), .ZN(n7641) );
  XNOR2_X1 U9311 ( .A(n7644), .B(n7641), .ZN(n7588) );
  XNOR2_X1 U9312 ( .A(n7646), .B(n7588), .ZN(n7595) );
  INV_X1 U9313 ( .A(n9835), .ZN(n9775) );
  AOI21_X1 U9314 ( .B1(n9785), .B2(n9848), .A(n7589), .ZN(n7592) );
  NAND2_X1 U9315 ( .A1(n9773), .A2(n7590), .ZN(n7591) );
  OAI211_X1 U9316 ( .C1(n10183), .C2(n9775), .A(n7592), .B(n7591), .ZN(n7593)
         );
  AOI21_X1 U9317 ( .B1(n10294), .B2(n4582), .A(n7593), .ZN(n7594) );
  OAI21_X1 U9318 ( .B1(n7595), .B2(n9825), .A(n7594), .ZN(P1_U3222) );
  XNOR2_X1 U9319 ( .A(n8902), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n7603) );
  INV_X1 U9320 ( .A(n7596), .ZN(n7598) );
  NAND2_X1 U9321 ( .A1(n7598), .A2(n7597), .ZN(n7599) );
  NAND2_X1 U9322 ( .A1(n7600), .A2(n7599), .ZN(n7602) );
  INV_X1 U9323 ( .A(n8904), .ZN(n7601) );
  AOI21_X1 U9324 ( .B1(n7603), .B2(n7602), .A(n7601), .ZN(n7613) );
  INV_X1 U9325 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8910) );
  MUX2_X1 U9326 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n8910), .S(n8902), .Z(n7607)
         );
  NAND2_X1 U9327 ( .A1(n8902), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7606) );
  OAI211_X1 U9328 ( .C1(n7608), .C2(n7607), .A(n8909), .B(n9291), .ZN(n7612)
         );
  NOR2_X1 U9329 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4656), .ZN(n7610) );
  NOR2_X1 U9330 ( .A1(n9286), .A2(n8911), .ZN(n7609) );
  AOI211_X1 U9331 ( .C1(n9289), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n7610), .B(
        n7609), .ZN(n7611) );
  OAI211_X1 U9332 ( .C1(n7613), .C2(n9295), .A(n7612), .B(n7611), .ZN(P2_U3261) );
  NAND2_X1 U9333 ( .A1(n7617), .A2(n7910), .ZN(n7619) );
  AOI22_X1 U9334 ( .A1(n7873), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n9864), .B2(
        n4368), .ZN(n7618) );
  OR2_X1 U9335 ( .A1(n10288), .A2(n10183), .ZN(n8468) );
  NAND2_X1 U9336 ( .A1(n10288), .A2(n10183), .ZN(n10177) );
  XNOR2_X1 U9337 ( .A(n8446), .B(n8273), .ZN(n10287) );
  INV_X1 U9338 ( .A(n7620), .ZN(n7939) );
  NAND2_X1 U9339 ( .A1(n7622), .A2(n7621), .ZN(n7623) );
  NAND2_X1 U9340 ( .A1(n7939), .A2(n7623), .ZN(n10169) );
  OR2_X1 U9341 ( .A1(n10169), .A2(n7050), .ZN(n7627) );
  INV_X1 U9342 ( .A(n8187), .ZN(n7942) );
  AOI22_X1 U9343 ( .A1(n4379), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n7942), .B2(
        P1_REG2_REG_14__SCAN_IN), .ZN(n7626) );
  INV_X1 U9344 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n7624) );
  OR2_X1 U9345 ( .A1(n8186), .A2(n7624), .ZN(n7625) );
  OAI22_X1 U9346 ( .A1(n9830), .A2(n10184), .B1(n10182), .B2(n7628), .ZN(n7634) );
  NAND2_X1 U9347 ( .A1(n7630), .A2(n7629), .ZN(n8232) );
  INV_X1 U9348 ( .A(n8318), .ZN(n8462) );
  OAI21_X1 U9349 ( .B1(n8464), .B2(n8462), .A(n8273), .ZN(n10180) );
  NAND3_X1 U9350 ( .A1(n4906), .A2(n8318), .A3(n8445), .ZN(n7632) );
  AOI21_X1 U9351 ( .B1(n10180), .B2(n7632), .A(n10179), .ZN(n7633) );
  AOI211_X1 U9352 ( .C1(n10287), .C2(n10153), .A(n7634), .B(n7633), .ZN(n10291) );
  INV_X1 U9353 ( .A(n10288), .ZN(n7638) );
  AOI21_X1 U9354 ( .B1(n10288), .B2(n7635), .A(n10166), .ZN(n10289) );
  NAND2_X1 U9355 ( .A1(n10289), .A2(n10156), .ZN(n7637) );
  AOI22_X1 U9356 ( .A1(n10437), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7658), .B2(
        n10170), .ZN(n7636) );
  OAI211_X1 U9357 ( .C1(n7638), .C2(n10433), .A(n7637), .B(n7636), .ZN(n7639)
         );
  AOI21_X1 U9358 ( .B1(n10287), .B2(n4484), .A(n7639), .ZN(n7640) );
  OAI21_X1 U9359 ( .B1(n10291), .B2(n10437), .A(n7640), .ZN(P1_U3278) );
  INV_X1 U9360 ( .A(n7644), .ZN(n7642) );
  NAND2_X1 U9361 ( .A1(n7642), .A2(n7641), .ZN(n7645) );
  NAND2_X1 U9362 ( .A1(n10288), .A2(n8940), .ZN(n7648) );
  NAND2_X1 U9363 ( .A1(n9846), .A2(n4367), .ZN(n7647) );
  NAND2_X1 U9364 ( .A1(n7648), .A2(n7647), .ZN(n7649) );
  XNOR2_X1 U9365 ( .A(n7649), .B(n8112), .ZN(n7655) );
  INV_X1 U9366 ( .A(n7655), .ZN(n7653) );
  NAND2_X1 U9367 ( .A1(n10288), .A2(n8934), .ZN(n7651) );
  NAND2_X1 U9368 ( .A1(n8935), .A2(n9846), .ZN(n7650) );
  NAND2_X1 U9369 ( .A1(n7651), .A2(n7650), .ZN(n7654) );
  INV_X1 U9370 ( .A(n7654), .ZN(n7652) );
  NAND2_X1 U9371 ( .A1(n7653), .A2(n7652), .ZN(n7927) );
  NAND2_X1 U9372 ( .A1(n7655), .A2(n7654), .ZN(n7925) );
  NAND2_X1 U9373 ( .A1(n7927), .A2(n7925), .ZN(n7656) );
  XNOR2_X1 U9374 ( .A(n7926), .B(n7656), .ZN(n7663) );
  AOI21_X1 U9375 ( .B1(n9785), .B2(n9847), .A(n7657), .ZN(n7660) );
  NAND2_X1 U9376 ( .A1(n9773), .A2(n7658), .ZN(n7659) );
  OAI211_X1 U9377 ( .C1(n9830), .C2(n9775), .A(n7660), .B(n7659), .ZN(n7661)
         );
  AOI21_X1 U9378 ( .B1(n10288), .B2(n4582), .A(n7661), .ZN(n7662) );
  OAI21_X1 U9379 ( .B1(n7663), .B2(n9825), .A(n7662), .ZN(P1_U3232) );
  INV_X1 U9380 ( .A(n7664), .ZN(n7667) );
  OAI21_X1 U9381 ( .B1(n7667), .B2(n7666), .A(n7665), .ZN(n7668) );
  XOR2_X1 U9382 ( .A(n7669), .B(n7668), .Z(n7729) );
  XOR2_X1 U9383 ( .A(n7670), .B(n7669), .Z(n7673) );
  OAI22_X1 U9384 ( .A1(n9531), .A2(n7671), .B1(n9014), .B2(n9528), .ZN(n7672)
         );
  AOI21_X1 U9385 ( .B1(n7673), .B2(n9524), .A(n7672), .ZN(n7674) );
  OAI21_X1 U9386 ( .B1(n7729), .B2(n7741), .A(n7674), .ZN(n7732) );
  INV_X1 U9387 ( .A(n7732), .ZN(n7675) );
  MUX2_X1 U9388 ( .A(n7676), .B(n7675), .S(n9536), .Z(n7682) );
  OAI21_X1 U9389 ( .B1(n7723), .B2(n7730), .A(n7692), .ZN(n7731) );
  INV_X1 U9390 ( .A(n7731), .ZN(n7680) );
  OAI22_X1 U9391 ( .A1(n9437), .A2(n7730), .B1(n9485), .B2(n7677), .ZN(n7678)
         );
  AOI21_X1 U9392 ( .B1(n7680), .B2(n7679), .A(n7678), .ZN(n7681) );
  OAI211_X1 U9393 ( .C1(n7729), .C2(n7756), .A(n7682), .B(n7681), .ZN(P2_U3286) );
  XNOR2_X1 U9394 ( .A(n7683), .B(n7686), .ZN(n9626) );
  NAND2_X1 U9395 ( .A1(n7685), .A2(n7684), .ZN(n7687) );
  XNOR2_X1 U9396 ( .A(n7687), .B(n7686), .ZN(n7688) );
  AOI222_X1 U9397 ( .A1(n9524), .A2(n7688), .B1(n9169), .B2(n9464), .C1(n9171), 
        .C2(n9462), .ZN(n9625) );
  MUX2_X1 U9398 ( .A(n7689), .B(n9625), .S(n9536), .Z(n7695) );
  INV_X1 U9399 ( .A(n7690), .ZN(n7691) );
  AOI211_X1 U9400 ( .C1(n9623), .C2(n7692), .A(n9538), .B(n7691), .ZN(n9622)
         );
  OAI22_X1 U9401 ( .A1(n9437), .A2(n4949), .B1(n7786), .B2(n9485), .ZN(n7693)
         );
  AOI21_X1 U9402 ( .B1(n9622), .B2(n9540), .A(n7693), .ZN(n7694) );
  OAI211_X1 U9403 ( .C1(n9495), .C2(n9626), .A(n7695), .B(n7694), .ZN(P2_U3285) );
  AOI211_X1 U9404 ( .C1(n7698), .C2(n10510), .A(n7697), .B(n7696), .ZN(n7703)
         );
  AOI22_X1 U9405 ( .A1(n5975), .A2(n7700), .B1(n10512), .B2(
        P2_REG0_REG_12__SCAN_IN), .ZN(n7699) );
  OAI21_X1 U9406 ( .B1(n7703), .B2(n10512), .A(n7699), .ZN(P2_U3487) );
  AOI22_X1 U9407 ( .A1(n7701), .A2(n7700), .B1(P2_REG1_REG_12__SCAN_IN), .B2(
        n10519), .ZN(n7702) );
  OAI21_X1 U9408 ( .B1(n7703), .B2(n10519), .A(n7702), .ZN(P2_U3532) );
  INV_X1 U9409 ( .A(n7704), .ZN(n7705) );
  INV_X1 U9410 ( .A(n7898), .ZN(n7707) );
  OAI222_X1 U9411 ( .A1(n7705), .A2(P1_U3084), .B1(n10347), .B2(n7707), .C1(
        n7899), .C2(n10350), .ZN(P1_U3327) );
  OAI222_X1 U9412 ( .A1(P2_U3152), .A2(n7708), .B1(n9684), .B2(n7707), .C1(
        n7706), .C2(n9686), .ZN(P2_U3332) );
  INV_X1 U9413 ( .A(n7903), .ZN(n7758) );
  AOI21_X1 U9414 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(n10340), .A(n7709), .ZN(
        n7710) );
  OAI21_X1 U9415 ( .B1(n7758), .B2(n10347), .A(n7710), .ZN(P1_U3326) );
  NOR2_X1 U9416 ( .A1(n7712), .A2(n7711), .ZN(n7713) );
  XNOR2_X1 U9417 ( .A(n7713), .B(n7716), .ZN(n9633) );
  OAI21_X1 U9418 ( .B1(n7716), .B2(n7715), .A(n7714), .ZN(n7720) );
  OAI22_X1 U9419 ( .A1(n9531), .A2(n7717), .B1(n7785), .B2(n9528), .ZN(n7719)
         );
  NOR2_X1 U9420 ( .A1(n9633), .A2(n7741), .ZN(n7718) );
  AOI211_X1 U9421 ( .C1(n9524), .C2(n7720), .A(n7719), .B(n7718), .ZN(n9632)
         );
  MUX2_X1 U9422 ( .A(n7721), .B(n9632), .S(n9536), .Z(n7728) );
  OAI22_X1 U9423 ( .A1(n9437), .A2(n7725), .B1(n9485), .B2(n7724), .ZN(n7726)
         );
  AOI21_X1 U9424 ( .B1(n9628), .B2(n9540), .A(n7726), .ZN(n7727) );
  OAI211_X1 U9425 ( .C1(n9633), .C2(n7756), .A(n7728), .B(n7727), .ZN(P2_U3287) );
  INV_X1 U9426 ( .A(n7729), .ZN(n7734) );
  OAI22_X1 U9427 ( .A1(n7731), .A2(n9538), .B1(n7730), .B2(n10507), .ZN(n7733)
         );
  AOI211_X1 U9428 ( .C1(n7735), .C2(n7734), .A(n7733), .B(n7732), .ZN(n7738)
         );
  NAND2_X1 U9429 ( .A1(n10512), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7736) );
  OAI21_X1 U9430 ( .B1(n7738), .B2(n10512), .A(n7736), .ZN(P2_U3481) );
  NAND2_X1 U9431 ( .A1(n10519), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7737) );
  OAI21_X1 U9432 ( .B1(n7738), .B2(n10519), .A(n7737), .ZN(P2_U3530) );
  OR2_X1 U9433 ( .A1(n7739), .A2(n5342), .ZN(n7761) );
  NAND2_X1 U9434 ( .A1(n7739), .A2(n5342), .ZN(n7740) );
  NAND2_X1 U9435 ( .A1(n7761), .A2(n7740), .ZN(n7808) );
  OR2_X1 U9436 ( .A1(n7808), .A2(n7741), .ZN(n7748) );
  NAND2_X1 U9437 ( .A1(n7743), .A2(n7742), .ZN(n7744) );
  NAND2_X1 U9438 ( .A1(n7765), .A2(n7744), .ZN(n7746) );
  OAI22_X1 U9439 ( .A1(n9531), .A2(n9086), .B1(n9146), .B2(n9528), .ZN(n7745)
         );
  AOI21_X1 U9440 ( .B1(n7746), .B2(n9524), .A(n7745), .ZN(n7747) );
  NAND2_X1 U9441 ( .A1(n7748), .A2(n7747), .ZN(n7809) );
  NAND2_X1 U9442 ( .A1(n7809), .A2(n9536), .ZN(n7755) );
  OAI22_X1 U9443 ( .A1(n9536), .A2(n7749), .B1(n9083), .B2(n9485), .ZN(n7753)
         );
  OAI21_X1 U9444 ( .B1(n7750), .B2(n9092), .A(n9484), .ZN(n7751) );
  OR2_X1 U9445 ( .A1(n7751), .A2(n7769), .ZN(n7806) );
  NOR2_X1 U9446 ( .A1(n7806), .A2(n9491), .ZN(n7752) );
  AOI211_X1 U9447 ( .C1(n9521), .C2(n7805), .A(n7753), .B(n7752), .ZN(n7754)
         );
  OAI211_X1 U9448 ( .C1(n7808), .C2(n7756), .A(n7755), .B(n7754), .ZN(P2_U3283) );
  OAI222_X1 U9449 ( .A1(n9686), .A2(n7759), .B1(n9684), .B2(n7758), .C1(n7757), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  NAND2_X1 U9450 ( .A1(n7761), .A2(n7760), .ZN(n7762) );
  XNOR2_X1 U9451 ( .A(n7762), .B(n4727), .ZN(n7817) );
  INV_X1 U9452 ( .A(n7817), .ZN(n7778) );
  NAND2_X1 U9453 ( .A1(n7763), .A2(n9524), .ZN(n7768) );
  AOI21_X1 U9454 ( .B1(n7765), .B2(n7764), .A(n4727), .ZN(n7767) );
  AOI22_X1 U9455 ( .A1(n9168), .A2(n9462), .B1(n9166), .B2(n9464), .ZN(n7766)
         );
  OAI21_X1 U9456 ( .B1(n7768), .B2(n7767), .A(n7766), .ZN(n7815) );
  INV_X1 U9457 ( .A(n7769), .ZN(n7771) );
  NAND2_X1 U9458 ( .A1(n7769), .A2(n8971), .ZN(n7799) );
  INV_X1 U9459 ( .A(n7799), .ZN(n7770) );
  AOI211_X1 U9460 ( .C1(n7772), .C2(n7771), .A(n9538), .B(n7770), .ZN(n7816)
         );
  NAND2_X1 U9461 ( .A1(n7816), .A2(n9540), .ZN(n7775) );
  INV_X1 U9462 ( .A(n7773), .ZN(n8973) );
  AOI22_X1 U9463 ( .A1(n4374), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8973), .B2(
        n9535), .ZN(n7774) );
  OAI211_X1 U9464 ( .C1(n8971), .C2(n9437), .A(n7775), .B(n7774), .ZN(n7776)
         );
  AOI21_X1 U9465 ( .B1(n9536), .B2(n7815), .A(n7776), .ZN(n7777) );
  OAI21_X1 U9466 ( .B1(n9495), .B2(n7778), .A(n7777), .ZN(P2_U3282) );
  INV_X1 U9467 ( .A(n7779), .ZN(n7780) );
  AOI21_X1 U9468 ( .B1(n7781), .B2(n7780), .A(n9138), .ZN(n7784) );
  NOR3_X1 U9469 ( .A1(n9136), .A2(n7785), .A3(n7782), .ZN(n7783) );
  OAI21_X1 U9470 ( .B1(n7784), .B2(n7783), .A(n9012), .ZN(n7790) );
  OAI22_X1 U9471 ( .A1(n9148), .A2(n9086), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9256), .ZN(n7788) );
  OAI22_X1 U9472 ( .A1(n9131), .A2(n7786), .B1(n7785), .B2(n9145), .ZN(n7787)
         );
  AOI211_X1 U9473 ( .C1(n9623), .C2(n9122), .A(n7788), .B(n7787), .ZN(n7789)
         );
  NAND2_X1 U9474 ( .A1(n7790), .A2(n7789), .ZN(P2_U3238) );
  INV_X1 U9475 ( .A(n7907), .ZN(n8928) );
  NAND2_X1 U9476 ( .A1(n9680), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7791) );
  OAI211_X1 U9477 ( .C1(n8928), .C2(n9684), .A(n7792), .B(n7791), .ZN(P2_U3330) );
  XNOR2_X1 U9478 ( .A(n7793), .B(n7796), .ZN(n7794) );
  AOI222_X1 U9479 ( .A1(n9524), .A2(n7794), .B1(n9165), .B2(n9464), .C1(n9167), 
        .C2(n9462), .ZN(n9620) );
  OAI21_X1 U9480 ( .B1(n7797), .B2(n7796), .A(n7795), .ZN(n9616) );
  INV_X1 U9481 ( .A(n7833), .ZN(n7798) );
  AOI211_X1 U9482 ( .C1(n9618), .C2(n7799), .A(n9538), .B(n7798), .ZN(n9617)
         );
  NAND2_X1 U9483 ( .A1(n9617), .A2(n9540), .ZN(n7802) );
  INV_X1 U9484 ( .A(n7800), .ZN(n9142) );
  AOI22_X1 U9485 ( .A1(n4374), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n9142), .B2(
        n9535), .ZN(n7801) );
  OAI211_X1 U9486 ( .C1(n9154), .C2(n9437), .A(n7802), .B(n7801), .ZN(n7803)
         );
  AOI21_X1 U9487 ( .B1(n9522), .B2(n9616), .A(n7803), .ZN(n7804) );
  OAI21_X1 U9488 ( .B1(n9620), .B2(n4374), .A(n7804), .ZN(P2_U3281) );
  NAND2_X1 U9489 ( .A1(n7805), .A2(n9630), .ZN(n7807) );
  OAI211_X1 U9490 ( .C1(n7808), .C2(n9634), .A(n7807), .B(n7806), .ZN(n7810)
         );
  NOR2_X1 U9491 ( .A1(n7810), .A2(n7809), .ZN(n7813) );
  INV_X1 U9492 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7811) );
  MUX2_X1 U9493 ( .A(n7813), .B(n7811), .S(n10512), .Z(n7812) );
  INV_X1 U9494 ( .A(n7812), .ZN(P2_U3490) );
  MUX2_X1 U9495 ( .A(n7813), .B(n8645), .S(n10519), .Z(n7814) );
  INV_X1 U9496 ( .A(n7814), .ZN(P2_U3533) );
  INV_X1 U9497 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7818) );
  AOI211_X1 U9498 ( .C1(n7817), .C2(n10510), .A(n7816), .B(n7815), .ZN(n7820)
         );
  MUX2_X1 U9499 ( .A(n7818), .B(n7820), .S(n10513), .Z(n7819) );
  OAI21_X1 U9500 ( .B1(n8971), .B2(n9670), .A(n7819), .ZN(P2_U3493) );
  MUX2_X1 U9501 ( .A(n8744), .B(n7820), .S(n10522), .Z(n7821) );
  OAI21_X1 U9502 ( .B1(n8971), .B2(n9615), .A(n7821), .ZN(P2_U3534) );
  XNOR2_X1 U9503 ( .A(n7823), .B(n7822), .ZN(n7827) );
  OR2_X1 U9504 ( .A1(n9479), .A2(n9528), .ZN(n7825) );
  NAND2_X1 U9505 ( .A1(n9166), .A2(n9462), .ZN(n7824) );
  NAND2_X1 U9506 ( .A1(n7825), .A2(n7824), .ZN(n9043) );
  INV_X1 U9507 ( .A(n9043), .ZN(n7826) );
  OAI21_X1 U9508 ( .B1(n7827), .B2(n9442), .A(n7826), .ZN(n9610) );
  INV_X1 U9509 ( .A(n9610), .ZN(n7838) );
  INV_X1 U9510 ( .A(n7828), .ZN(n7829) );
  AOI21_X1 U9511 ( .B1(n7831), .B2(n7830), .A(n7829), .ZN(n9612) );
  NAND2_X1 U9512 ( .A1(n9612), .A2(n9522), .ZN(n7837) );
  INV_X1 U9513 ( .A(n9508), .ZN(n7832) );
  AOI211_X1 U9514 ( .C1(n9047), .C2(n7833), .A(n9538), .B(n7832), .ZN(n9611)
         );
  NOR2_X1 U9515 ( .A1(n9437), .A2(n9671), .ZN(n7835) );
  OAI22_X1 U9516 ( .A1(n9536), .A2(n8910), .B1(n9045), .B2(n9485), .ZN(n7834)
         );
  AOI211_X1 U9517 ( .C1(n9611), .C2(n9540), .A(n7835), .B(n7834), .ZN(n7836)
         );
  OAI211_X1 U9518 ( .C1(n7838), .C2(n4374), .A(n7837), .B(n7836), .ZN(P2_U3280) );
  INV_X1 U9519 ( .A(n7839), .ZN(n7841) );
  NAND3_X1 U9520 ( .A1(n7843), .A2(n7842), .A3(n9524), .ZN(n7845) );
  INV_X1 U9521 ( .A(n9129), .ZN(n9158) );
  INV_X1 U9522 ( .A(n7844), .ZN(n9156) );
  AOI22_X1 U9523 ( .A1(n9158), .A2(n9462), .B1(n9156), .B2(n9464), .ZN(n8895)
         );
  AOI211_X1 U9524 ( .C1(n9548), .C2(n9324), .A(n9538), .B(n7846), .ZN(n9549)
         );
  NAND2_X1 U9525 ( .A1(n9549), .A2(n9540), .ZN(n7848) );
  AOI22_X1 U9526 ( .A1(n8892), .A2(n9535), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n4374), .ZN(n7847) );
  OAI211_X1 U9527 ( .C1(n5001), .C2(n9437), .A(n7848), .B(n7847), .ZN(n7849)
         );
  AOI21_X1 U9528 ( .B1(n9550), .B2(n9536), .A(n7849), .ZN(n7850) );
  OAI21_X1 U9529 ( .B1(n9553), .B2(n9495), .A(n7850), .ZN(P2_U3268) );
  NAND2_X1 U9530 ( .A1(n8931), .A2(n7902), .ZN(n7854) );
  INV_X1 U9531 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10345) );
  OR2_X1 U9532 ( .A1(n7911), .A2(n10345), .ZN(n7853) );
  NAND2_X1 U9533 ( .A1(n7855), .A2(n7910), .ZN(n7857) );
  INV_X1 U9534 ( .A(n9884), .ZN(n9867) );
  AOI22_X1 U9535 ( .A1(n7873), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n9867), .B2(
        n4368), .ZN(n7856) );
  INV_X1 U9536 ( .A(n10283), .ZN(n10173) );
  NAND2_X1 U9537 ( .A1(n7858), .A2(n7902), .ZN(n7860) );
  AOI22_X1 U9538 ( .A1(n7873), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n4368), .B2(
        n9888), .ZN(n7859) );
  INV_X1 U9539 ( .A(n10277), .ZN(n10161) );
  NAND2_X1 U9540 ( .A1(n7861), .A2(n7902), .ZN(n7863) );
  AOI22_X1 U9541 ( .A1(n9932), .A2(n4368), .B1(n7873), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n7862) );
  NAND2_X1 U9542 ( .A1(n7864), .A2(n7910), .ZN(n7866) );
  AOI22_X1 U9543 ( .A1(n7873), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9917), .B2(
        n4368), .ZN(n7865) );
  NAND2_X2 U9544 ( .A1(n7866), .A2(n7865), .ZN(n10273) );
  OR2_X1 U9545 ( .A1(n10266), .A2(n10273), .ZN(n7867) );
  NAND2_X1 U9546 ( .A1(n7868), .A2(n7902), .ZN(n7870) );
  AOI22_X1 U9547 ( .A1(n9944), .A2(n4368), .B1(n7873), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n7869) );
  INV_X1 U9548 ( .A(n10258), .ZN(n10099) );
  NAND2_X1 U9549 ( .A1(n7871), .A2(n7910), .ZN(n7875) );
  AOI22_X1 U9550 ( .A1(n7873), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n4368), .B2(
        n9951), .ZN(n7874) );
  INV_X1 U9551 ( .A(n10253), .ZN(n10087) );
  NAND2_X1 U9552 ( .A1(n7876), .A2(n7902), .ZN(n7879) );
  OR2_X1 U9553 ( .A1(n7911), .A2(n7877), .ZN(n7878) );
  OR2_X1 U9554 ( .A1(n7911), .A2(n8629), .ZN(n7881) );
  NAND2_X1 U9555 ( .A1(n8959), .A2(n7910), .ZN(n7884) );
  OR2_X1 U9556 ( .A1(n7911), .A2(n8961), .ZN(n7883) );
  NAND2_X1 U9557 ( .A1(n7885), .A2(n7910), .ZN(n7888) );
  OR2_X1 U9558 ( .A1(n7911), .A2(n7886), .ZN(n7887) );
  OR2_X1 U9559 ( .A1(n7911), .A2(n7890), .ZN(n7891) );
  NOR2_X2 U9560 ( .A1(n10019), .A2(n10229), .ZN(n7893) );
  INV_X1 U9561 ( .A(n7893), .ZN(n10005) );
  OR2_X1 U9562 ( .A1(n7911), .A2(n7895), .ZN(n7896) );
  OR2_X1 U9563 ( .A1(n7911), .A2(n7899), .ZN(n7900) );
  OR2_X1 U9564 ( .A1(n7911), .A2(n7904), .ZN(n7905) );
  OR2_X1 U9565 ( .A1(n7911), .A2(n8930), .ZN(n7908) );
  NAND2_X1 U9566 ( .A1(n9682), .A2(n7910), .ZN(n7913) );
  OR2_X1 U9567 ( .A1(n7911), .A2(n10349), .ZN(n7912) );
  NAND2_X1 U9568 ( .A1(n9956), .A2(n9955), .ZN(n7914) );
  INV_X1 U9569 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n7922) );
  INV_X1 U9570 ( .A(P1_B_REG_SCAN_IN), .ZN(n7915) );
  NOR2_X1 U9571 ( .A1(n7916), .A2(n7915), .ZN(n7917) );
  OR2_X1 U9572 ( .A1(n10184), .A2(n7917), .ZN(n8500) );
  INV_X1 U9573 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n7921) );
  OR2_X1 U9574 ( .A1(n8187), .A2(n7922), .ZN(n7920) );
  INV_X1 U9575 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n7918) );
  OR2_X1 U9576 ( .A1(n8186), .A2(n7918), .ZN(n7919) );
  OAI211_X1 U9577 ( .C1(n4380), .C2(n7921), .A(n7920), .B(n7919), .ZN(n9839)
         );
  INV_X1 U9578 ( .A(n9839), .ZN(n8374) );
  NOR2_X1 U9579 ( .A1(n8500), .A2(n8374), .ZN(n10196) );
  NAND2_X1 U9580 ( .A1(n10139), .A2(n10196), .ZN(n9957) );
  OAI21_X1 U9581 ( .B1(n10139), .B2(n7922), .A(n9957), .ZN(n7923) );
  AOI21_X1 U9582 ( .B1(n10193), .B2(n9960), .A(n7923), .ZN(n7924) );
  OAI21_X1 U9583 ( .B1(n10195), .B2(n10434), .A(n7924), .ZN(P1_U3261) );
  NAND2_X1 U9584 ( .A1(n7926), .A2(n7925), .ZN(n7928) );
  NAND2_X1 U9585 ( .A1(n7928), .A2(n7927), .ZN(n7934) );
  NAND2_X1 U9586 ( .A1(n10283), .A2(n8940), .ZN(n7930) );
  INV_X1 U9587 ( .A(n9830), .ZN(n10146) );
  NAND2_X1 U9588 ( .A1(n10146), .A2(n8934), .ZN(n7929) );
  NAND2_X1 U9589 ( .A1(n7930), .A2(n7929), .ZN(n7931) );
  XNOR2_X1 U9590 ( .A(n7931), .B(n8938), .ZN(n7935) );
  NAND2_X1 U9591 ( .A1(n7934), .A2(n7935), .ZN(n9688) );
  NAND2_X1 U9592 ( .A1(n10283), .A2(n8934), .ZN(n7933) );
  NAND2_X1 U9593 ( .A1(n10146), .A2(n8935), .ZN(n7932) );
  NAND2_X1 U9594 ( .A1(n7933), .A2(n7932), .ZN(n9691) );
  INV_X1 U9595 ( .A(n7934), .ZN(n7937) );
  INV_X1 U9596 ( .A(n7935), .ZN(n7936) );
  NAND2_X1 U9597 ( .A1(n10277), .A2(n8940), .ZN(n7947) );
  INV_X1 U9598 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7938) );
  NAND2_X1 U9599 ( .A1(n7939), .A2(n7938), .ZN(n7940) );
  NAND2_X1 U9600 ( .A1(n7973), .A2(n7940), .ZN(n10157) );
  OR2_X1 U9601 ( .A1(n10157), .A2(n7050), .ZN(n7945) );
  INV_X1 U9602 ( .A(n8186), .ZN(n7941) );
  AOI22_X1 U9603 ( .A1(n7942), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n7941), .B2(
        P1_REG0_REG_15__SCAN_IN), .ZN(n7944) );
  NAND2_X1 U9604 ( .A1(n4379), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n7943) );
  OR2_X1 U9605 ( .A1(n10185), .A2(n8942), .ZN(n7946) );
  NAND2_X1 U9606 ( .A1(n7947), .A2(n7946), .ZN(n7948) );
  XNOR2_X1 U9607 ( .A(n7948), .B(n8112), .ZN(n7951) );
  NAND2_X1 U9608 ( .A1(n10277), .A2(n4367), .ZN(n7950) );
  OR2_X1 U9609 ( .A1(n10185), .A2(n8154), .ZN(n7949) );
  NAND2_X1 U9610 ( .A1(n7950), .A2(n7949), .ZN(n9822) );
  NAND2_X1 U9611 ( .A1(n10273), .A2(n8940), .ZN(n7954) );
  OR2_X1 U9612 ( .A1(n9760), .A2(n8942), .ZN(n7953) );
  NAND2_X1 U9613 ( .A1(n7954), .A2(n7953), .ZN(n7955) );
  XNOR2_X1 U9614 ( .A(n7955), .B(n8112), .ZN(n9748) );
  NAND2_X1 U9615 ( .A1(n10273), .A2(n4367), .ZN(n7957) );
  OR2_X1 U9616 ( .A1(n9760), .A2(n8154), .ZN(n7956) );
  NAND2_X1 U9617 ( .A1(n7957), .A2(n7956), .ZN(n9749) );
  NAND2_X1 U9618 ( .A1(n10258), .A2(n8940), .ZN(n7967) );
  NAND2_X1 U9619 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_REG3_REG_16__SCAN_IN), 
        .ZN(n7958) );
  INV_X1 U9620 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8634) );
  INV_X1 U9621 ( .A(n7990), .ZN(n7992) );
  NAND2_X1 U9622 ( .A1(n7974), .A2(n8634), .ZN(n7959) );
  NAND2_X1 U9623 ( .A1(n7992), .A2(n7959), .ZN(n10100) );
  OR2_X1 U9624 ( .A1(n10100), .A2(n7050), .ZN(n7965) );
  INV_X1 U9625 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9924) );
  INV_X1 U9626 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10101) );
  OR2_X1 U9627 ( .A1(n8187), .A2(n10101), .ZN(n7962) );
  INV_X1 U9628 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n7960) );
  OR2_X1 U9629 ( .A1(n8186), .A2(n7960), .ZN(n7961) );
  OAI211_X1 U9630 ( .C1(n4380), .C2(n9924), .A(n7962), .B(n7961), .ZN(n7963)
         );
  INV_X1 U9631 ( .A(n7963), .ZN(n7964) );
  NAND2_X1 U9632 ( .A1(n10115), .A2(n8934), .ZN(n7966) );
  NAND2_X1 U9633 ( .A1(n7967), .A2(n7966), .ZN(n7968) );
  XNOR2_X1 U9634 ( .A(n7968), .B(n8938), .ZN(n9713) );
  NAND2_X1 U9635 ( .A1(n10258), .A2(n4367), .ZN(n7970) );
  NAND2_X1 U9636 ( .A1(n10115), .A2(n8935), .ZN(n7969) );
  NAND2_X1 U9637 ( .A1(n7970), .A2(n7969), .ZN(n9715) );
  NAND2_X1 U9638 ( .A1(n10266), .A2(n8940), .ZN(n7985) );
  INV_X1 U9639 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7972) );
  INV_X1 U9640 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n7971) );
  OAI21_X1 U9641 ( .B1(n7973), .B2(n7972), .A(n7971), .ZN(n7975) );
  AND2_X1 U9642 ( .A1(n7975), .A2(n7974), .ZN(n10110) );
  NAND2_X1 U9643 ( .A1(n10110), .A2(n8184), .ZN(n7983) );
  INV_X1 U9644 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n7980) );
  INV_X1 U9645 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n7976) );
  OR2_X1 U9646 ( .A1(n8187), .A2(n7976), .ZN(n7979) );
  INV_X1 U9647 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n7977) );
  OR2_X1 U9648 ( .A1(n8186), .A2(n7977), .ZN(n7978) );
  OAI211_X1 U9649 ( .C1(n4380), .C2(n7980), .A(n7979), .B(n7978), .ZN(n7981)
         );
  INV_X1 U9650 ( .A(n7981), .ZN(n7982) );
  INV_X1 U9651 ( .A(n10131), .ZN(n10095) );
  NAND2_X1 U9652 ( .A1(n10095), .A2(n8934), .ZN(n7984) );
  NAND2_X1 U9653 ( .A1(n7985), .A2(n7984), .ZN(n7986) );
  XNOR2_X1 U9654 ( .A(n7986), .B(n8938), .ZN(n8005) );
  INV_X1 U9655 ( .A(n8005), .ZN(n7989) );
  NOR2_X1 U9656 ( .A1(n10131), .A2(n8154), .ZN(n7987) );
  AOI21_X1 U9657 ( .B1(n10266), .B2(n4367), .A(n7987), .ZN(n8004) );
  INV_X1 U9658 ( .A(n8004), .ZN(n7988) );
  NAND2_X1 U9659 ( .A1(n7989), .A2(n7988), .ZN(n9711) );
  OAI21_X1 U9660 ( .B1(n9713), .B2(n9804), .A(n9711), .ZN(n8009) );
  NAND2_X1 U9661 ( .A1(n10253), .A2(n8940), .ZN(n8001) );
  INV_X1 U9662 ( .A(n8012), .ZN(n8014) );
  INV_X1 U9663 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7991) );
  NAND2_X1 U9664 ( .A1(n7992), .A2(n7991), .ZN(n7993) );
  NAND2_X1 U9665 ( .A1(n10084), .A2(n8184), .ZN(n7999) );
  INV_X1 U9666 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9945) );
  INV_X1 U9667 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n7994) );
  OR2_X1 U9668 ( .A1(n8187), .A2(n7994), .ZN(n7996) );
  INV_X1 U9669 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n8631) );
  OR2_X1 U9670 ( .A1(n8186), .A2(n8631), .ZN(n7995) );
  OAI211_X1 U9671 ( .C1(n4380), .C2(n9945), .A(n7996), .B(n7995), .ZN(n7997)
         );
  INV_X1 U9672 ( .A(n7997), .ZN(n7998) );
  NAND2_X1 U9673 ( .A1(n10094), .A2(n8934), .ZN(n8000) );
  NAND2_X1 U9674 ( .A1(n8001), .A2(n8000), .ZN(n8002) );
  XNOR2_X1 U9675 ( .A(n8002), .B(n8938), .ZN(n9717) );
  NOR2_X1 U9676 ( .A1(n10063), .A2(n8154), .ZN(n8003) );
  AOI21_X1 U9677 ( .B1(n10253), .B2(n8934), .A(n8003), .ZN(n9716) );
  NAND2_X1 U9678 ( .A1(n9717), .A2(n9716), .ZN(n8008) );
  NAND2_X1 U9679 ( .A1(n8005), .A2(n8004), .ZN(n9712) );
  NAND2_X1 U9680 ( .A1(n9712), .A2(n9715), .ZN(n8006) );
  INV_X1 U9681 ( .A(n9712), .ZN(n9758) );
  AOI22_X1 U9682 ( .A1(n9713), .A2(n8006), .B1(n9758), .B2(n9804), .ZN(n8007)
         );
  INV_X1 U9683 ( .A(n9717), .ZN(n8011) );
  INV_X1 U9684 ( .A(n9716), .ZN(n8010) );
  NAND2_X1 U9685 ( .A1(n8011), .A2(n8010), .ZN(n9781) );
  NAND2_X1 U9686 ( .A1(n10249), .A2(n8940), .ZN(n8024) );
  INV_X1 U9687 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8013) );
  NAND2_X1 U9688 ( .A1(n8014), .A2(n8013), .ZN(n8015) );
  NAND2_X1 U9689 ( .A1(n8030), .A2(n8015), .ZN(n10067) );
  OR2_X1 U9690 ( .A1(n10067), .A2(n7050), .ZN(n8022) );
  INV_X1 U9691 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n8019) );
  INV_X1 U9692 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n10068) );
  OR2_X1 U9693 ( .A1(n8187), .A2(n10068), .ZN(n8018) );
  INV_X1 U9694 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n8016) );
  OR2_X1 U9695 ( .A1(n8186), .A2(n8016), .ZN(n8017) );
  OAI211_X1 U9696 ( .C1(n4380), .C2(n8019), .A(n8018), .B(n8017), .ZN(n8020)
         );
  INV_X1 U9697 ( .A(n8020), .ZN(n8021) );
  NAND2_X1 U9698 ( .A1(n10047), .A2(n4367), .ZN(n8023) );
  NAND2_X1 U9699 ( .A1(n8024), .A2(n8023), .ZN(n8025) );
  XNOR2_X1 U9700 ( .A(n8025), .B(n8938), .ZN(n8046) );
  INV_X1 U9701 ( .A(n8046), .ZN(n8028) );
  AND2_X1 U9702 ( .A1(n10047), .A2(n8935), .ZN(n8026) );
  AOI21_X1 U9703 ( .B1(n10249), .B2(n4367), .A(n8026), .ZN(n8045) );
  INV_X1 U9704 ( .A(n8045), .ZN(n8027) );
  NAND2_X1 U9705 ( .A1(n8028), .A2(n8027), .ZN(n9780) );
  NAND2_X1 U9706 ( .A1(n10243), .A2(n8940), .ZN(n8040) );
  INV_X1 U9707 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8029) );
  NAND2_X1 U9708 ( .A1(n8030), .A2(n8029), .ZN(n8031) );
  AND2_X1 U9709 ( .A1(n8052), .A2(n8031), .ZN(n10052) );
  NAND2_X1 U9710 ( .A1(n10052), .A2(n8184), .ZN(n8038) );
  INV_X1 U9711 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n8035) );
  INV_X1 U9712 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n10055) );
  OR2_X1 U9713 ( .A1(n8187), .A2(n10055), .ZN(n8034) );
  INV_X1 U9714 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n8032) );
  OR2_X1 U9715 ( .A1(n8186), .A2(n8032), .ZN(n8033) );
  OAI211_X1 U9716 ( .C1(n4380), .C2(n8035), .A(n8034), .B(n8033), .ZN(n8036)
         );
  INV_X1 U9717 ( .A(n8036), .ZN(n8037) );
  OR2_X1 U9718 ( .A1(n10064), .A2(n8942), .ZN(n8039) );
  NAND2_X1 U9719 ( .A1(n8040), .A2(n8039), .ZN(n8041) );
  XNOR2_X1 U9720 ( .A(n8041), .B(n8112), .ZN(n8048) );
  NAND2_X1 U9721 ( .A1(n10243), .A2(n4367), .ZN(n8043) );
  OR2_X1 U9722 ( .A1(n10064), .A2(n8154), .ZN(n8042) );
  NAND2_X1 U9723 ( .A1(n8043), .A2(n8042), .ZN(n8049) );
  INV_X1 U9724 ( .A(n9728), .ZN(n8044) );
  NAND2_X1 U9725 ( .A1(n8046), .A2(n8045), .ZN(n9779) );
  INV_X1 U9726 ( .A(n8048), .ZN(n8051) );
  INV_X1 U9727 ( .A(n8049), .ZN(n8050) );
  NAND2_X1 U9728 ( .A1(n8051), .A2(n8050), .ZN(n9727) );
  INV_X1 U9729 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9796) );
  NOR2_X2 U9730 ( .A1(n8052), .A2(n9796), .ZN(n8072) );
  INV_X1 U9731 ( .A(n8072), .ZN(n8086) );
  NAND2_X1 U9732 ( .A1(n8052), .A2(n9796), .ZN(n8053) );
  NAND2_X1 U9733 ( .A1(n8086), .A2(n8053), .ZN(n10033) );
  OR2_X1 U9734 ( .A1(n10033), .A2(n7050), .ZN(n8061) );
  INV_X1 U9735 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n8058) );
  INV_X1 U9736 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n8054) );
  OR2_X1 U9737 ( .A1(n8186), .A2(n8054), .ZN(n8057) );
  INV_X1 U9738 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n8055) );
  OR2_X1 U9739 ( .A1(n8187), .A2(n8055), .ZN(n8056) );
  OAI211_X1 U9740 ( .C1(n4380), .C2(n8058), .A(n8057), .B(n8056), .ZN(n8059)
         );
  INV_X1 U9741 ( .A(n8059), .ZN(n8060) );
  AND2_X2 U9742 ( .A1(n8061), .A2(n8060), .ZN(n10014) );
  NOR2_X1 U9743 ( .A1(n10014), .A2(n8154), .ZN(n8062) );
  AOI21_X1 U9744 ( .B1(n10237), .B2(n4367), .A(n8062), .ZN(n8067) );
  NAND2_X1 U9745 ( .A1(n8063), .A2(n8067), .ZN(n9792) );
  NAND2_X1 U9746 ( .A1(n10237), .A2(n8940), .ZN(n8065) );
  OR2_X1 U9747 ( .A1(n10014), .A2(n8942), .ZN(n8064) );
  NAND2_X1 U9748 ( .A1(n8065), .A2(n8064), .ZN(n8066) );
  XNOR2_X1 U9749 ( .A(n8066), .B(n8112), .ZN(n9793) );
  INV_X1 U9750 ( .A(n8067), .ZN(n8068) );
  NAND2_X1 U9751 ( .A1(n8099), .A2(n9791), .ZN(n9700) );
  NAND2_X1 U9752 ( .A1(n10229), .A2(n8940), .ZN(n8083) );
  INV_X1 U9753 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9705) );
  INV_X1 U9754 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8070) );
  OAI21_X1 U9755 ( .B1(n8086), .B2(n9705), .A(n8070), .ZN(n8073) );
  AND2_X1 U9756 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .ZN(n8071) );
  INV_X1 U9757 ( .A(n8100), .ZN(n8102) );
  NAND2_X1 U9758 ( .A1(n8073), .A2(n8102), .ZN(n9772) );
  INV_X1 U9759 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n8078) );
  INV_X1 U9760 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n8074) );
  OR2_X1 U9761 ( .A1(n8186), .A2(n8074), .ZN(n8077) );
  INV_X1 U9762 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n8075) );
  OR2_X1 U9763 ( .A1(n8187), .A2(n8075), .ZN(n8076) );
  OAI211_X1 U9764 ( .C1(n4380), .C2(n8078), .A(n8077), .B(n8076), .ZN(n8079)
         );
  INV_X1 U9765 ( .A(n8079), .ZN(n8080) );
  NAND2_X1 U9766 ( .A1(n9844), .A2(n8934), .ZN(n8082) );
  NAND2_X1 U9767 ( .A1(n8083), .A2(n8082), .ZN(n8084) );
  XNOR2_X1 U9768 ( .A(n8084), .B(n8938), .ZN(n8116) );
  NOR2_X1 U9769 ( .A1(n10015), .A2(n8154), .ZN(n8085) );
  AOI21_X1 U9770 ( .B1(n10229), .B2(n4367), .A(n8085), .ZN(n8115) );
  INV_X1 U9771 ( .A(n9740), .ZN(n8098) );
  NAND2_X1 U9772 ( .A1(n10232), .A2(n8940), .ZN(n8096) );
  NAND2_X1 U9773 ( .A1(n10021), .A2(n8184), .ZN(n8094) );
  INV_X1 U9774 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n8091) );
  INV_X1 U9775 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n8087) );
  OR2_X1 U9776 ( .A1(n8187), .A2(n8087), .ZN(n8090) );
  INV_X1 U9777 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n8088) );
  OR2_X1 U9778 ( .A1(n8186), .A2(n8088), .ZN(n8089) );
  OAI211_X1 U9779 ( .C1(n4380), .C2(n8091), .A(n8090), .B(n8089), .ZN(n8092)
         );
  INV_X1 U9780 ( .A(n8092), .ZN(n8093) );
  OR2_X1 U9781 ( .A1(n10004), .A2(n8942), .ZN(n8095) );
  NAND2_X1 U9782 ( .A1(n8096), .A2(n8095), .ZN(n8097) );
  XNOR2_X1 U9783 ( .A(n8097), .B(n8938), .ZN(n8117) );
  NAND3_X1 U9784 ( .A1(n9700), .A2(n8098), .A3(n9699), .ZN(n8123) );
  NAND2_X1 U9785 ( .A1(n10222), .A2(n8940), .ZN(n8111) );
  INV_X1 U9786 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8101) );
  NAND2_X1 U9787 ( .A1(n8102), .A2(n8101), .ZN(n8103) );
  NAND2_X1 U9788 ( .A1(n8124), .A2(n8103), .ZN(n8459) );
  INV_X1 U9789 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n8728) );
  INV_X1 U9790 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n8600) );
  OR2_X1 U9791 ( .A1(n8186), .A2(n8600), .ZN(n8106) );
  INV_X1 U9792 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n8104) );
  OR2_X1 U9793 ( .A1(n8187), .A2(n8104), .ZN(n8105) );
  OAI211_X1 U9794 ( .C1(n4380), .C2(n8728), .A(n8106), .B(n8105), .ZN(n8107)
         );
  INV_X1 U9795 ( .A(n8107), .ZN(n8108) );
  INV_X1 U9796 ( .A(n9993), .ZN(n10001) );
  NAND2_X1 U9797 ( .A1(n10001), .A2(n8934), .ZN(n8110) );
  NAND2_X1 U9798 ( .A1(n8111), .A2(n8110), .ZN(n8113) );
  XNOR2_X1 U9799 ( .A(n8113), .B(n8112), .ZN(n8137) );
  NOR2_X1 U9800 ( .A1(n9993), .A2(n8154), .ZN(n8114) );
  AOI21_X1 U9801 ( .B1(n10222), .B2(n4367), .A(n8114), .ZN(n8138) );
  XNOR2_X1 U9802 ( .A(n8137), .B(n8138), .ZN(n9739) );
  OR2_X1 U9803 ( .A1(n8116), .A2(n8115), .ZN(n9737) );
  NAND4_X1 U9804 ( .A1(n9791), .A2(n9739), .A3(n8117), .A4(n9737), .ZN(n8121)
         );
  NOR2_X1 U9805 ( .A1(n10004), .A2(n8154), .ZN(n8118) );
  AOI21_X1 U9806 ( .B1(n10232), .B2(n8934), .A(n8118), .ZN(n9701) );
  AOI21_X1 U9807 ( .B1(n9701), .B2(n9737), .A(n9740), .ZN(n8120) );
  INV_X1 U9808 ( .A(n9739), .ZN(n8119) );
  OAI22_X1 U9809 ( .A1(n9698), .A2(n8121), .B1(n8120), .B2(n8119), .ZN(n8122)
         );
  AND2_X2 U9810 ( .A1(n8123), .A2(n8122), .ZN(n9813) );
  INV_X1 U9811 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9817) );
  OR2_X2 U9812 ( .A1(n8124), .A2(n9817), .ZN(n8142) );
  NAND2_X1 U9813 ( .A1(n8124), .A2(n9817), .ZN(n8125) );
  NAND2_X1 U9814 ( .A1(n8142), .A2(n8125), .ZN(n9985) );
  INV_X1 U9815 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n8128) );
  INV_X1 U9816 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n8696) );
  OR2_X1 U9817 ( .A1(n8186), .A2(n8696), .ZN(n8127) );
  INV_X1 U9818 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9984) );
  OR2_X1 U9819 ( .A1(n8187), .A2(n9984), .ZN(n8126) );
  OAI211_X1 U9820 ( .C1(n4380), .C2(n8128), .A(n8127), .B(n8126), .ZN(n8129)
         );
  INV_X1 U9821 ( .A(n8129), .ZN(n8130) );
  NOR2_X1 U9822 ( .A1(n9969), .A2(n8154), .ZN(n8132) );
  AOI21_X1 U9823 ( .B1(n10219), .B2(n4367), .A(n8132), .ZN(n8158) );
  NAND2_X1 U9824 ( .A1(n10219), .A2(n8940), .ZN(n8134) );
  NAND2_X1 U9825 ( .A1(n9843), .A2(n8934), .ZN(n8133) );
  NAND2_X1 U9826 ( .A1(n8134), .A2(n8133), .ZN(n8136) );
  XNOR2_X1 U9827 ( .A(n8136), .B(n8112), .ZN(n8160) );
  XOR2_X1 U9828 ( .A(n8158), .B(n8160), .Z(n9811) );
  INV_X1 U9829 ( .A(n8137), .ZN(n8139) );
  NAND2_X1 U9830 ( .A1(n10214), .A2(n8940), .ZN(n8152) );
  INV_X1 U9831 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8141) );
  OR2_X2 U9832 ( .A1(n8142), .A2(n8141), .ZN(n8183) );
  NAND2_X1 U9833 ( .A1(n8142), .A2(n8141), .ZN(n8143) );
  NAND2_X1 U9834 ( .A1(n9973), .A2(n8184), .ZN(n8150) );
  INV_X1 U9835 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8147) );
  INV_X1 U9836 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n8699) );
  OR2_X1 U9837 ( .A1(n8186), .A2(n8699), .ZN(n8146) );
  INV_X1 U9838 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n8144) );
  OR2_X1 U9839 ( .A1(n8187), .A2(n8144), .ZN(n8145) );
  OAI211_X1 U9840 ( .C1(n4380), .C2(n8147), .A(n8146), .B(n8145), .ZN(n8148)
         );
  INV_X1 U9841 ( .A(n8148), .ZN(n8149) );
  AND2_X2 U9842 ( .A1(n8150), .A2(n8149), .ZN(n9994) );
  NAND2_X1 U9843 ( .A1(n9842), .A2(n4367), .ZN(n8151) );
  NAND2_X1 U9844 ( .A1(n8152), .A2(n8151), .ZN(n8153) );
  XNOR2_X1 U9845 ( .A(n8153), .B(n8938), .ZN(n8157) );
  NOR2_X1 U9846 ( .A1(n9994), .A2(n8154), .ZN(n8155) );
  AOI21_X1 U9847 ( .B1(n10214), .B2(n8934), .A(n8155), .ZN(n8156) );
  NAND2_X1 U9848 ( .A1(n8157), .A2(n8156), .ZN(n8951) );
  OAI21_X1 U9849 ( .B1(n8157), .B2(n8156), .A(n8951), .ZN(n8162) );
  INV_X1 U9850 ( .A(n8158), .ZN(n8159) );
  INV_X1 U9851 ( .A(n8161), .ZN(n8164) );
  INV_X1 U9852 ( .A(n8162), .ZN(n8163) );
  NAND2_X1 U9853 ( .A1(n8948), .A2(n8184), .ZN(n8171) );
  INV_X1 U9854 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n8168) );
  INV_X1 U9855 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n8755) );
  OR2_X1 U9856 ( .A1(n8187), .A2(n8755), .ZN(n8167) );
  INV_X1 U9857 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n8165) );
  OR2_X1 U9858 ( .A1(n8186), .A2(n8165), .ZN(n8166) );
  OAI211_X1 U9859 ( .C1(n4380), .C2(n8168), .A(n8167), .B(n8166), .ZN(n8169)
         );
  INV_X1 U9860 ( .A(n8169), .ZN(n8170) );
  INV_X1 U9861 ( .A(n8943), .ZN(n9966) );
  AOI22_X1 U9862 ( .A1(n9973), .A2(n9773), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8172) );
  OAI21_X1 U9863 ( .B1(n9969), .B2(n9831), .A(n8172), .ZN(n8173) );
  AOI21_X1 U9864 ( .B1(n9966), .B2(n9835), .A(n8173), .ZN(n8174) );
  OAI222_X1 U9865 ( .A1(n10350), .A2(n8176), .B1(n10347), .B2(n8175), .C1(
        P1_U3084), .C2(n4373), .ZN(P1_U3350) );
  INV_X1 U9866 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8643) );
  INV_X1 U9867 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9958) );
  OR2_X1 U9868 ( .A1(n8187), .A2(n9958), .ZN(n8180) );
  INV_X1 U9869 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n8178) );
  OR2_X1 U9870 ( .A1(n8186), .A2(n8178), .ZN(n8179) );
  OAI211_X1 U9871 ( .C1(n4380), .C2(n8643), .A(n8180), .B(n8179), .ZN(n9840)
         );
  INV_X1 U9872 ( .A(n9840), .ZN(n8501) );
  OR2_X1 U9873 ( .A1(n10197), .A2(n8501), .ZN(n8181) );
  NAND2_X1 U9874 ( .A1(n8380), .A2(n8181), .ZN(n8379) );
  INV_X1 U9875 ( .A(n8379), .ZN(n8284) );
  NAND2_X1 U9876 ( .A1(n10214), .A2(n9994), .ZN(n8287) );
  OR2_X2 U9877 ( .A1(n10214), .A2(n9994), .ZN(n8497) );
  NAND2_X1 U9878 ( .A1(n10219), .A2(n9969), .ZN(n8366) );
  NAND2_X1 U9879 ( .A1(n8497), .A2(n8495), .ZN(n8182) );
  NAND3_X1 U9880 ( .A1(n8498), .A2(n8287), .A3(n8182), .ZN(n8419) );
  OR2_X1 U9881 ( .A1(n10219), .A2(n9969), .ZN(n8365) );
  OR2_X1 U9882 ( .A1(n8419), .A2(n8496), .ZN(n8194) );
  INV_X1 U9883 ( .A(n8183), .ZN(n8510) );
  NAND3_X1 U9884 ( .A1(n8510), .A2(n8184), .A3(P1_REG3_REG_28__SCAN_IN), .ZN(
        n8193) );
  INV_X1 U9885 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n8614) );
  INV_X1 U9886 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8185) );
  OR2_X1 U9887 ( .A1(n8186), .A2(n8185), .ZN(n8189) );
  INV_X1 U9888 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8513) );
  OR2_X1 U9889 ( .A1(n8187), .A2(n8513), .ZN(n8188) );
  OAI211_X1 U9890 ( .C1(n4380), .C2(n8614), .A(n8189), .B(n8188), .ZN(n8191)
         );
  INV_X1 U9891 ( .A(n8191), .ZN(n8192) );
  NAND3_X1 U9892 ( .A1(n8194), .A2(n8370), .A3(n8254), .ZN(n8423) );
  AND2_X2 U9893 ( .A1(n8497), .A2(n8287), .ZN(n9964) );
  NAND2_X1 U9894 ( .A1(n8487), .A2(n8486), .ZN(n8288) );
  INV_X1 U9895 ( .A(n8288), .ZN(n8361) );
  OR2_X1 U9896 ( .A1(n10243), .A2(n10064), .ZN(n8354) );
  INV_X1 U9897 ( .A(n8354), .ZN(n8199) );
  NAND2_X1 U9898 ( .A1(n10253), .A2(n10063), .ZN(n8344) );
  INV_X1 U9899 ( .A(n8344), .ZN(n8478) );
  NOR2_X1 U9900 ( .A1(n10258), .A2(n10079), .ZN(n8345) );
  INV_X1 U9901 ( .A(n8345), .ZN(n8257) );
  OR2_X1 U9902 ( .A1(n10266), .A2(n10131), .ZN(n10091) );
  NAND2_X1 U9903 ( .A1(n8257), .A2(n10091), .ZN(n8195) );
  NAND2_X1 U9904 ( .A1(n10258), .A2(n10079), .ZN(n8256) );
  NAND2_X1 U9905 ( .A1(n8195), .A2(n8256), .ZN(n8476) );
  INV_X1 U9906 ( .A(n10047), .ZN(n10080) );
  OR2_X1 U9907 ( .A1(n10249), .A2(n10080), .ZN(n8479) );
  OAI211_X1 U9908 ( .C1(n8478), .C2(n8476), .A(n8479), .B(n8341), .ZN(n8198)
         );
  NAND2_X1 U9909 ( .A1(n10237), .A2(n10014), .ZN(n8483) );
  NAND2_X1 U9910 ( .A1(n10243), .A2(n10064), .ZN(n8482) );
  NAND2_X1 U9911 ( .A1(n8483), .A2(n8482), .ZN(n8355) );
  INV_X1 U9912 ( .A(n8355), .ZN(n8197) );
  NAND2_X1 U9913 ( .A1(n10249), .A2(n10080), .ZN(n8480) );
  INV_X1 U9914 ( .A(n8480), .ZN(n8196) );
  NAND2_X1 U9915 ( .A1(n8354), .A2(n8196), .ZN(n8202) );
  OAI211_X1 U9916 ( .C1(n8199), .C2(n8198), .A(n8197), .B(n8202), .ZN(n8200)
         );
  OR2_X2 U9917 ( .A1(n10237), .A2(n10014), .ZN(n8484) );
  AND2_X1 U9918 ( .A1(n8200), .A2(n8484), .ZN(n8201) );
  NAND2_X1 U9919 ( .A1(n8361), .A2(n8201), .ZN(n8417) );
  INV_X1 U9920 ( .A(n8417), .ZN(n8248) );
  INV_X1 U9921 ( .A(n8202), .ZN(n8203) );
  OR3_X1 U9922 ( .A1(n8355), .A2(n8203), .A3(n8478), .ZN(n8412) );
  INV_X1 U9923 ( .A(n8412), .ZN(n8244) );
  NAND2_X1 U9924 ( .A1(n10266), .A2(n10131), .ZN(n10090) );
  NAND2_X1 U9925 ( .A1(n8256), .A2(n10090), .ZN(n8477) );
  NAND2_X1 U9926 ( .A1(n10277), .A2(n10185), .ZN(n10126) );
  AND2_X1 U9927 ( .A1(n8318), .A2(n8204), .ZN(n8324) );
  NAND2_X1 U9928 ( .A1(n10126), .A2(n8324), .ZN(n8229) );
  NAND2_X1 U9929 ( .A1(n8306), .A2(n8298), .ZN(n8209) );
  NAND2_X1 U9930 ( .A1(n10283), .A2(n9830), .ZN(n8461) );
  NAND2_X1 U9931 ( .A1(n10177), .A2(n8461), .ZN(n8469) );
  INV_X1 U9932 ( .A(n8311), .ZN(n8307) );
  NAND2_X1 U9933 ( .A1(n8317), .A2(n8307), .ZN(n8206) );
  AND2_X1 U9934 ( .A1(n8206), .A2(n8205), .ZN(n8207) );
  NOR2_X1 U9935 ( .A1(n8469), .A2(n8207), .ZN(n8226) );
  NAND2_X1 U9936 ( .A1(n8226), .A2(n8471), .ZN(n8208) );
  OR4_X1 U9937 ( .A1(n8477), .A2(n8229), .A3(n8209), .A4(n8208), .ZN(n8397) );
  NAND2_X1 U9938 ( .A1(n8210), .A2(n8299), .ZN(n8297) );
  INV_X1 U9939 ( .A(n8297), .ZN(n8212) );
  NAND2_X1 U9940 ( .A1(n8212), .A2(n8211), .ZN(n8398) );
  NAND2_X1 U9941 ( .A1(n8401), .A2(n8213), .ZN(n8214) );
  NOR2_X1 U9942 ( .A1(n8398), .A2(n8214), .ZN(n8409) );
  AOI21_X1 U9943 ( .B1(n9857), .B2(n6459), .A(n8426), .ZN(n8216) );
  AND2_X1 U9944 ( .A1(n8216), .A2(n8215), .ZN(n8219) );
  OAI22_X1 U9945 ( .A1(n8220), .A2(n8219), .B1(n8218), .B2(n8217), .ZN(n8222)
         );
  NAND3_X1 U9946 ( .A1(n8222), .A2(n8399), .A3(n8221), .ZN(n8223) );
  NAND2_X1 U9947 ( .A1(n8409), .A2(n8223), .ZN(n8224) );
  OAI21_X1 U9948 ( .B1(n8225), .B2(n8398), .A(n8224), .ZN(n8242) );
  INV_X1 U9949 ( .A(n8226), .ZN(n8239) );
  AND2_X1 U9950 ( .A1(n8228), .A2(n8227), .ZN(n8308) );
  INV_X1 U9951 ( .A(n8308), .ZN(n8231) );
  INV_X1 U9952 ( .A(n8229), .ZN(n8230) );
  OAI21_X1 U9953 ( .B1(n8320), .B2(n8231), .A(n8230), .ZN(n8238) );
  NAND2_X1 U9954 ( .A1(n8332), .A2(n8470), .ZN(n8331) );
  INV_X1 U9955 ( .A(n8331), .ZN(n8237) );
  AND2_X1 U9956 ( .A1(n8468), .A2(n8465), .ZN(n8326) );
  INV_X1 U9957 ( .A(n8326), .ZN(n8234) );
  AND2_X1 U9958 ( .A1(n8232), .A2(n8318), .ZN(n8233) );
  NOR2_X1 U9959 ( .A1(n8234), .A2(n8233), .ZN(n8328) );
  INV_X1 U9960 ( .A(n8328), .ZN(n8235) );
  NAND2_X1 U9961 ( .A1(n8469), .A2(n8465), .ZN(n8330) );
  NAND3_X1 U9962 ( .A1(n8235), .A2(n8330), .A3(n10126), .ZN(n8236) );
  OAI211_X1 U9963 ( .C1(n8239), .C2(n8238), .A(n8237), .B(n8236), .ZN(n8240)
         );
  NAND2_X1 U9964 ( .A1(n8240), .A2(n8471), .ZN(n8241) );
  OR2_X1 U9965 ( .A1(n8477), .A2(n8241), .ZN(n8414) );
  OAI21_X1 U9966 ( .B1(n8397), .B2(n8242), .A(n8414), .ZN(n8243) );
  NAND2_X1 U9967 ( .A1(n8244), .A2(n8243), .ZN(n8247) );
  NAND2_X1 U9968 ( .A1(n8487), .A2(n8255), .ZN(n8245) );
  NAND2_X1 U9969 ( .A1(n10229), .A2(n10015), .ZN(n8359) );
  AND2_X1 U9970 ( .A1(n8245), .A2(n8359), .ZN(n8246) );
  NAND2_X1 U9971 ( .A1(n8493), .A2(n8246), .ZN(n8415) );
  AOI21_X1 U9972 ( .B1(n8248), .B2(n8247), .A(n8415), .ZN(n8249) );
  NOR2_X1 U9973 ( .A1(n8507), .A2(n8249), .ZN(n8250) );
  NOR2_X1 U9974 ( .A1(n8419), .A2(n8250), .ZN(n8251) );
  NAND2_X1 U9975 ( .A1(n10197), .A2(n8501), .ZN(n8376) );
  NAND2_X1 U9976 ( .A1(n10201), .A2(n8947), .ZN(n8421) );
  OAI211_X1 U9977 ( .C1(n8423), .C2(n8251), .A(n8376), .B(n8421), .ZN(n8252)
         );
  AOI21_X1 U9978 ( .B1(n8284), .B2(n8252), .A(n8425), .ZN(n8253) );
  XNOR2_X1 U9979 ( .A(n8253), .B(n9951), .ZN(n8437) );
  INV_X1 U9980 ( .A(n8376), .ZN(n8282) );
  NAND2_X1 U9981 ( .A1(n10219), .A2(n9843), .ZN(n8505) );
  NAND2_X1 U9982 ( .A1(n8506), .A2(n8505), .ZN(n9990) );
  NAND2_X2 U9983 ( .A1(n8360), .A2(n8486), .ZN(n10013) );
  XNOR2_X1 U9984 ( .A(n10237), .B(n10014), .ZN(n10038) );
  XNOR2_X1 U9985 ( .A(n10243), .B(n10064), .ZN(n8352) );
  NAND2_X1 U9986 ( .A1(n8257), .A2(n8256), .ZN(n10104) );
  AND2_X1 U9987 ( .A1(n10091), .A2(n10090), .ZN(n10113) );
  NOR2_X1 U9988 ( .A1(n8258), .A2(n4375), .ZN(n8266) );
  NAND4_X1 U9989 ( .A1(n8259), .A2(n8260), .A3(n8261), .A4(n6447), .ZN(n8263)
         );
  NOR2_X1 U9990 ( .A1(n8263), .A2(n8262), .ZN(n8264) );
  NAND4_X1 U9991 ( .A1(n8266), .A2(n8293), .A3(n8265), .A4(n8264), .ZN(n8268)
         );
  OR3_X1 U9992 ( .A1(n8268), .A2(n8313), .A3(n8267), .ZN(n8269) );
  NOR2_X1 U9993 ( .A1(n8270), .A2(n8269), .ZN(n8272) );
  NAND4_X1 U9994 ( .A1(n8273), .A2(n10176), .A3(n8272), .A4(n8271), .ZN(n8274)
         );
  NAND2_X1 U9995 ( .A1(n8470), .A2(n10126), .ZN(n10145) );
  NOR2_X1 U9996 ( .A1(n8274), .A2(n10145), .ZN(n8275) );
  NAND3_X1 U9997 ( .A1(n10113), .A2(n10128), .A3(n8275), .ZN(n8276) );
  NOR2_X1 U9998 ( .A1(n10104), .A2(n8276), .ZN(n8277) );
  XNOR2_X1 U9999 ( .A(n10249), .B(n10047), .ZN(n10060) );
  NAND4_X1 U10000 ( .A1(n4720), .A2(n8451), .A3(n8277), .A4(n10060), .ZN(n8278) );
  NOR3_X1 U10001 ( .A1(n10013), .A2(n10038), .A3(n8278), .ZN(n8279) );
  NAND4_X1 U10002 ( .A1(n9990), .A2(n8488), .A3(n9999), .A4(n8279), .ZN(n8280)
         );
  AOI21_X1 U10003 ( .B1(n8285), .B2(n8284), .A(n8283), .ZN(n8430) );
  INV_X1 U10004 ( .A(n8430), .ZN(n8433) );
  NAND2_X1 U10005 ( .A1(n8286), .A2(n9951), .ZN(n8435) );
  MUX2_X1 U10006 ( .A(n8497), .B(n8287), .S(n8388), .Z(n8369) );
  NAND2_X1 U10007 ( .A1(n8288), .A2(n8359), .ZN(n8289) );
  NAND2_X1 U10008 ( .A1(n9988), .A2(n8289), .ZN(n8290) );
  MUX2_X1 U10009 ( .A(n8415), .B(n8290), .S(n8388), .Z(n8364) );
  NAND2_X1 U10010 ( .A1(n8403), .A2(n8388), .ZN(n8295) );
  OAI211_X1 U10011 ( .C1(n8296), .C2(n8295), .A(n8294), .B(n8293), .ZN(n8304)
         );
  NAND2_X1 U10012 ( .A1(n8297), .A2(n8298), .ZN(n8302) );
  NAND2_X1 U10013 ( .A1(n8405), .A2(n8298), .ZN(n8300) );
  NAND2_X1 U10014 ( .A1(n8300), .A2(n8299), .ZN(n8301) );
  MUX2_X1 U10015 ( .A(n8302), .B(n8301), .S(n8388), .Z(n8303) );
  AND2_X1 U10016 ( .A1(n8307), .A2(n8306), .ZN(n8309) );
  MUX2_X1 U10017 ( .A(n8309), .B(n8308), .S(n8381), .Z(n8315) );
  MUX2_X1 U10018 ( .A(n8311), .B(n8310), .S(n8388), .Z(n8312) );
  OR2_X1 U10019 ( .A1(n8313), .A2(n8312), .ZN(n8314) );
  AOI21_X1 U10020 ( .B1(n8316), .B2(n8315), .A(n8314), .ZN(n8323) );
  NAND2_X1 U10021 ( .A1(n8318), .A2(n8317), .ZN(n8319) );
  MUX2_X1 U10022 ( .A(n8320), .B(n8319), .S(n8388), .Z(n8322) );
  NAND4_X1 U10023 ( .A1(n8327), .A2(n8381), .A3(n8332), .A4(n8470), .ZN(n8340)
         );
  NAND2_X1 U10024 ( .A1(n8329), .A2(n8328), .ZN(n8338) );
  AND4_X1 U10025 ( .A1(n8471), .A2(n8388), .A3(n8330), .A4(n10126), .ZN(n8337)
         );
  NAND3_X1 U10026 ( .A1(n8331), .A2(n8388), .A3(n8471), .ZN(n8335) );
  NAND2_X1 U10027 ( .A1(n8471), .A2(n10126), .ZN(n8333) );
  NAND3_X1 U10028 ( .A1(n8333), .A2(n8381), .A3(n8332), .ZN(n8334) );
  NAND2_X1 U10029 ( .A1(n8335), .A2(n8334), .ZN(n8336) );
  AOI21_X1 U10030 ( .B1(n8338), .B2(n8337), .A(n8336), .ZN(n8339) );
  NAND2_X1 U10031 ( .A1(n8340), .A2(n8339), .ZN(n8343) );
  NAND2_X1 U10032 ( .A1(n8343), .A2(n4893), .ZN(n8342) );
  NAND4_X1 U10033 ( .A1(n8342), .A2(n8388), .A3(n8476), .A4(n8341), .ZN(n8351)
         );
  AOI21_X1 U10034 ( .B1(n8343), .B2(n10091), .A(n8477), .ZN(n8346) );
  OAI211_X1 U10035 ( .C1(n8346), .C2(n8345), .A(n8381), .B(n8344), .ZN(n8350)
         );
  AND2_X1 U10036 ( .A1(n10094), .A2(n8381), .ZN(n8348) );
  OAI21_X1 U10037 ( .B1(n8381), .B2(n10094), .A(n10253), .ZN(n8347) );
  OAI21_X1 U10038 ( .B1(n8348), .B2(n10253), .A(n8347), .ZN(n8349) );
  MUX2_X1 U10039 ( .A(n8479), .B(n8480), .S(n8388), .Z(n8353) );
  NAND2_X1 U10040 ( .A1(n8484), .A2(n8354), .ZN(n8356) );
  MUX2_X1 U10041 ( .A(n8356), .B(n8355), .S(n8388), .Z(n8358) );
  MUX2_X1 U10042 ( .A(n8483), .B(n8484), .S(n8388), .Z(n8357) );
  MUX2_X1 U10043 ( .A(n9988), .B(n8493), .S(n8388), .Z(n8362) );
  OAI211_X1 U10044 ( .C1(n8364), .C2(n8363), .A(n8362), .B(n9990), .ZN(n8368)
         );
  MUX2_X1 U10045 ( .A(n8366), .B(n8365), .S(n8388), .Z(n8367) );
  MUX2_X1 U10046 ( .A(n8370), .B(n8498), .S(n8381), .Z(n8371) );
  NAND2_X1 U10047 ( .A1(n8387), .A2(n8947), .ZN(n8372) );
  MUX2_X1 U10048 ( .A(n8372), .B(n8388), .S(n10201), .Z(n8373) );
  OAI21_X1 U10049 ( .B1(n8381), .B2(n8947), .A(n8373), .ZN(n8394) );
  NAND2_X1 U10050 ( .A1(n8379), .A2(n10193), .ZN(n8428) );
  INV_X1 U10051 ( .A(n8428), .ZN(n8377) );
  NAND2_X1 U10052 ( .A1(n10197), .A2(n8374), .ZN(n8375) );
  INV_X1 U10053 ( .A(n8422), .ZN(n8383) );
  NOR2_X1 U10054 ( .A1(n8377), .A2(n8383), .ZN(n8390) );
  INV_X1 U10055 ( .A(n8390), .ZN(n8393) );
  INV_X1 U10056 ( .A(n8380), .ZN(n8382) );
  NOR3_X1 U10057 ( .A1(n8382), .A2(n8422), .A3(n8381), .ZN(n8385) );
  INV_X1 U10058 ( .A(n8387), .ZN(n8389) );
  NAND4_X1 U10059 ( .A1(n8390), .A2(n8389), .A3(n8388), .A4(n10201), .ZN(n8391) );
  OAI211_X1 U10060 ( .C1(n8394), .C2(n8393), .A(n8392), .B(n8391), .ZN(n8436)
         );
  INV_X1 U10061 ( .A(n8425), .ZN(n8395) );
  NAND4_X1 U10062 ( .A1(n8436), .A2(n8396), .A3(n4372), .A4(n8395), .ZN(n8432)
         );
  INV_X1 U10063 ( .A(n8397), .ZN(n8411) );
  INV_X1 U10064 ( .A(n8398), .ZN(n8407) );
  NAND2_X1 U10065 ( .A1(n8400), .A2(n8399), .ZN(n8402) );
  NAND2_X1 U10066 ( .A1(n8402), .A2(n8401), .ZN(n8404) );
  NAND3_X1 U10067 ( .A1(n8405), .A2(n8404), .A3(n8403), .ZN(n8406) );
  AOI22_X1 U10068 ( .A1(n8409), .A2(n8408), .B1(n8407), .B2(n8406), .ZN(n8410)
         );
  NAND2_X1 U10069 ( .A1(n8411), .A2(n8410), .ZN(n8413) );
  AOI21_X1 U10070 ( .B1(n8414), .B2(n8413), .A(n8412), .ZN(n8418) );
  INV_X1 U10071 ( .A(n8415), .ZN(n8416) );
  OAI21_X1 U10072 ( .B1(n8418), .B2(n8417), .A(n8416), .ZN(n8420) );
  AOI21_X1 U10073 ( .B1(n8497), .B2(n8420), .A(n8419), .ZN(n8424) );
  OAI211_X1 U10074 ( .C1(n8424), .C2(n8423), .A(n8422), .B(n8421), .ZN(n8427)
         );
  AOI211_X1 U10075 ( .C1(n8428), .C2(n8427), .A(n8426), .B(n8425), .ZN(n8429)
         );
  NAND2_X1 U10076 ( .A1(n8440), .A2(n8439), .ZN(n8441) );
  OAI211_X1 U10077 ( .C1(n8442), .C2(n8444), .A(n8441), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8443) );
  INV_X1 U10078 ( .A(n10266), .ZN(n10112) );
  INV_X1 U10079 ( .A(n10273), .ZN(n10137) );
  INV_X1 U10080 ( .A(n10185), .ZN(n9845) );
  OR2_X1 U10081 ( .A1(n10277), .A2(n9845), .ZN(n10122) );
  INV_X1 U10082 ( .A(n10122), .ZN(n8447) );
  NOR2_X1 U10083 ( .A1(n10145), .A2(n8447), .ZN(n8448) );
  NAND2_X1 U10084 ( .A1(n8472), .A2(n8448), .ZN(n8449) );
  NAND3_X1 U10085 ( .A1(n10105), .A2(n10077), .A3(n10104), .ZN(n8454) );
  NAND2_X1 U10086 ( .A1(n10258), .A2(n10115), .ZN(n10074) );
  NAND2_X1 U10087 ( .A1(n10253), .A2(n10094), .ZN(n8450) );
  INV_X1 U10088 ( .A(n8452), .ZN(n8453) );
  INV_X1 U10089 ( .A(n10249), .ZN(n10066) );
  NAND2_X1 U10090 ( .A1(n10066), .A2(n10080), .ZN(n8455) );
  INV_X1 U10091 ( .A(n10014), .ZN(n10048) );
  INV_X1 U10092 ( .A(n10026), .ZN(n8456) );
  NAND2_X1 U10093 ( .A1(n9997), .A2(n5039), .ZN(n8458) );
  XNOR2_X1 U10094 ( .A(n8504), .B(n8488), .ZN(n10226) );
  AOI21_X1 U10095 ( .B1(n10222), .B2(n10005), .A(n9980), .ZN(n10223) );
  INV_X1 U10096 ( .A(n8459), .ZN(n9742) );
  AOI22_X1 U10097 ( .A1(n9742), .A2(n10170), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10437), .ZN(n8460) );
  OAI21_X1 U10098 ( .B1(n9747), .B2(n10433), .A(n8460), .ZN(n8491) );
  INV_X1 U10099 ( .A(n8461), .ZN(n8463) );
  INV_X1 U10100 ( .A(n10177), .ZN(n10174) );
  INV_X1 U10101 ( .A(n8465), .ZN(n8466) );
  OR2_X1 U10102 ( .A1(n8469), .A2(n8468), .ZN(n10124) );
  NAND2_X1 U10103 ( .A1(n10125), .A2(n5051), .ZN(n8475) );
  OAI21_X1 U10104 ( .B1(n8472), .B2(n10126), .A(n8471), .ZN(n8473) );
  INV_X1 U10105 ( .A(n8473), .ZN(n8474) );
  INV_X1 U10106 ( .A(n8479), .ZN(n8481) );
  INV_X1 U10107 ( .A(n8483), .ZN(n8485) );
  INV_X1 U10108 ( .A(n10013), .ZN(n10027) );
  NAND2_X1 U10109 ( .A1(n9998), .A2(n8487), .ZN(n8494) );
  XNOR2_X1 U10110 ( .A(n8494), .B(n8503), .ZN(n8489) );
  AOI222_X1 U10111 ( .A1(n10117), .A2(n8489), .B1(n9844), .B2(n10147), .C1(
        n9843), .C2(n10148), .ZN(n10225) );
  NOR2_X1 U10112 ( .A1(n10225), .A2(n10437), .ZN(n8490) );
  AOI211_X1 U10113 ( .C1(n10223), .C2(n10156), .A(n8491), .B(n8490), .ZN(n8492) );
  OAI21_X1 U10114 ( .B1(n10226), .B2(n10192), .A(n8492), .ZN(P1_U3266) );
  AND2_X2 U10115 ( .A1(n9963), .A2(n8497), .ZN(n8536) );
  OAI22_X1 U10116 ( .A1(n8943), .A2(n10182), .B1(n8501), .B2(n8500), .ZN(n8502) );
  XNOR2_X1 U10117 ( .A(n8509), .B(n8499), .ZN(n10200) );
  NAND2_X1 U10118 ( .A1(n10200), .A2(n4524), .ZN(n8516) );
  AOI21_X1 U10119 ( .B1(n10201), .B2(n8540), .A(n9955), .ZN(n10202) );
  NAND2_X1 U10120 ( .A1(n10201), .A2(n9960), .ZN(n8512) );
  NAND3_X1 U10121 ( .A1(n8510), .A2(P1_REG3_REG_28__SCAN_IN), .A3(n10170), 
        .ZN(n8511) );
  OAI211_X1 U10122 ( .C1(n10139), .C2(n8513), .A(n8512), .B(n8511), .ZN(n8514)
         );
  AOI21_X1 U10123 ( .B1(n10202), .B2(n10156), .A(n8514), .ZN(n8515) );
  OAI211_X1 U10124 ( .C1(n10204), .C2(n10437), .A(n8516), .B(n8515), .ZN(
        P1_U3355) );
  INV_X1 U10125 ( .A(n8517), .ZN(n8523) );
  OAI211_X1 U10126 ( .C1(n8520), .C2(n8519), .A(n9258), .B(n8518), .ZN(n8521)
         );
  INV_X1 U10127 ( .A(n8521), .ZN(n8522) );
  AOI211_X1 U10128 ( .C1(n9289), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n8523), .B(
        n8522), .ZN(n8529) );
  INV_X1 U10129 ( .A(n8524), .ZN(n9200) );
  NAND3_X1 U10130 ( .A1(n9186), .A2(n8526), .A3(n8525), .ZN(n8527) );
  NAND3_X1 U10131 ( .A1(n9291), .A2(n9200), .A3(n8527), .ZN(n8528) );
  OAI211_X1 U10132 ( .C1(n9286), .C2(n8530), .A(n8529), .B(n8528), .ZN(
        P2_U3249) );
  OAI22_X1 U10133 ( .A1(n9994), .A2(n10182), .B1(n8947), .B2(n10184), .ZN(
        n8537) );
  NAND2_X1 U10134 ( .A1(n9970), .A2(n10207), .ZN(n8539) );
  NAND2_X1 U10135 ( .A1(n10208), .A2(n10156), .ZN(n8542) );
  AOI22_X1 U10136 ( .A1(n8948), .A2(n10170), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n10437), .ZN(n8541) );
  OAI211_X1 U10137 ( .C1(n4918), .C2(n10433), .A(n8542), .B(n8541), .ZN(n8543)
         );
  INV_X1 U10138 ( .A(n8543), .ZN(n8544) );
  XNOR2_X1 U10139 ( .A(n8546), .B(keyinput17), .ZN(n8552) );
  XOR2_X1 U10140 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput85), .Z(n8551) );
  XNOR2_X1 U10141 ( .A(n8547), .B(keyinput15), .ZN(n8550) );
  XNOR2_X1 U10142 ( .A(n8548), .B(keyinput44), .ZN(n8549) );
  NOR4_X1 U10143 ( .A1(n8552), .A2(n8551), .A3(n8550), .A4(n8549), .ZN(n8574)
         );
  XNOR2_X1 U10144 ( .A(n8553), .B(keyinput36), .ZN(n8559) );
  XNOR2_X1 U10145 ( .A(n8554), .B(keyinput121), .ZN(n8558) );
  XNOR2_X1 U10146 ( .A(n4598), .B(keyinput101), .ZN(n8557) );
  XNOR2_X1 U10147 ( .A(n8555), .B(keyinput18), .ZN(n8556) );
  NOR4_X1 U10148 ( .A1(n8559), .A2(n8558), .A3(n8557), .A4(n8556), .ZN(n8573)
         );
  XOR2_X1 U10149 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput70), .Z(n8565) );
  XOR2_X1 U10150 ( .A(P2_REG0_REG_24__SCAN_IN), .B(keyinput59), .Z(n8564) );
  XNOR2_X1 U10151 ( .A(n8560), .B(keyinput94), .ZN(n8563) );
  XNOR2_X1 U10152 ( .A(n8561), .B(keyinput106), .ZN(n8562) );
  NOR4_X1 U10153 ( .A1(n8565), .A2(n8564), .A3(n8563), .A4(n8562), .ZN(n8572)
         );
  XNOR2_X1 U10154 ( .A(SI_25_), .B(keyinput41), .ZN(n8567) );
  XNOR2_X1 U10155 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput21), .ZN(n8566) );
  NAND2_X1 U10156 ( .A1(n8567), .A2(n8566), .ZN(n8569) );
  XOR2_X1 U10157 ( .A(SI_5_), .B(keyinput60), .Z(n8568) );
  AOI211_X1 U10158 ( .C1(keyinput12), .C2(n8570), .A(n8569), .B(n8568), .ZN(
        n8571) );
  NAND4_X1 U10159 ( .A1(n8574), .A2(n8573), .A3(n8572), .A4(n8571), .ZN(n8585)
         );
  AOI22_X1 U10160 ( .A1(n8576), .A2(keyinput77), .B1(keyinput43), .B2(n6474), 
        .ZN(n8575) );
  OAI221_X1 U10161 ( .B1(n8576), .B2(keyinput77), .C1(n6474), .C2(keyinput43), 
        .A(n8575), .ZN(n8584) );
  AOI22_X1 U10162 ( .A1(n8579), .A2(keyinput71), .B1(n8578), .B2(keyinput45), 
        .ZN(n8577) );
  OAI221_X1 U10163 ( .B1(n8579), .B2(keyinput71), .C1(n8578), .C2(keyinput45), 
        .A(n8577), .ZN(n8583) );
  INV_X1 U10164 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10446) );
  AOI22_X1 U10165 ( .A1(n10446), .A2(keyinput14), .B1(keyinput119), .B2(n8581), 
        .ZN(n8580) );
  OAI221_X1 U10166 ( .B1(n10446), .B2(keyinput14), .C1(n8581), .C2(keyinput119), .A(n8580), .ZN(n8582) );
  NOR4_X1 U10167 ( .A1(n8585), .A2(n8584), .A3(n8583), .A4(n8582), .ZN(n8627)
         );
  AOI22_X1 U10168 ( .A1(n6917), .A2(keyinput20), .B1(n6661), .B2(keyinput103), 
        .ZN(n8586) );
  OAI221_X1 U10169 ( .B1(n6917), .B2(keyinput20), .C1(n6661), .C2(keyinput103), 
        .A(n8586), .ZN(n8594) );
  INV_X1 U10170 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n8588) );
  AOI22_X1 U10171 ( .A1(n8588), .A2(keyinput90), .B1(keyinput73), .B2(n9029), 
        .ZN(n8587) );
  OAI221_X1 U10172 ( .B1(n8588), .B2(keyinput90), .C1(n9029), .C2(keyinput73), 
        .A(n8587), .ZN(n8593) );
  INV_X1 U10173 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10444) );
  AOI22_X1 U10174 ( .A1(n8776), .A2(keyinput98), .B1(keyinput95), .B2(n10444), 
        .ZN(n8589) );
  OAI221_X1 U10175 ( .B1(n8776), .B2(keyinput98), .C1(n10444), .C2(keyinput95), 
        .A(n8589), .ZN(n8592) );
  INV_X1 U10176 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n10473) );
  AOI22_X1 U10177 ( .A1(n8742), .A2(keyinput57), .B1(n10473), .B2(keyinput91), 
        .ZN(n8590) );
  OAI221_X1 U10178 ( .B1(n8742), .B2(keyinput57), .C1(n10473), .C2(keyinput91), 
        .A(n8590), .ZN(n8591) );
  NOR4_X1 U10179 ( .A1(n8594), .A2(n8593), .A3(n8592), .A4(n8591), .ZN(n8626)
         );
  AOI22_X1 U10180 ( .A1(n8787), .A2(keyinput96), .B1(keyinput31), .B2(n9487), 
        .ZN(n8595) );
  OAI221_X1 U10181 ( .B1(n8787), .B2(keyinput96), .C1(n9487), .C2(keyinput31), 
        .A(n8595), .ZN(n8604) );
  AOI22_X1 U10182 ( .A1(n8598), .A2(keyinput99), .B1(keyinput56), .B2(n8597), 
        .ZN(n8596) );
  OAI221_X1 U10183 ( .B1(n8598), .B2(keyinput99), .C1(n8597), .C2(keyinput56), 
        .A(n8596), .ZN(n8603) );
  AOI22_X1 U10184 ( .A1(n8601), .A2(keyinput83), .B1(keyinput13), .B2(n8600), 
        .ZN(n8599) );
  OAI221_X1 U10185 ( .B1(n8601), .B2(keyinput83), .C1(n8600), .C2(keyinput13), 
        .A(n8599), .ZN(n8602) );
  OR3_X1 U10186 ( .A1(n8604), .A2(n8603), .A3(n8602), .ZN(n8610) );
  INV_X1 U10187 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n10468) );
  AOI22_X1 U10188 ( .A1(n10468), .A2(keyinput0), .B1(keyinput9), .B2(n10517), 
        .ZN(n8605) );
  OAI221_X1 U10189 ( .B1(n10468), .B2(keyinput0), .C1(n10517), .C2(keyinput9), 
        .A(n8605), .ZN(n8609) );
  AOI22_X1 U10190 ( .A1(n8607), .A2(keyinput89), .B1(keyinput127), .B2(n5173), 
        .ZN(n8606) );
  OAI221_X1 U10191 ( .B1(n8607), .B2(keyinput89), .C1(n5173), .C2(keyinput127), 
        .A(n8606), .ZN(n8608) );
  NOR3_X1 U10192 ( .A1(n8610), .A2(n8609), .A3(n8608), .ZN(n8625) );
  INV_X1 U10193 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n8612) );
  AOI22_X1 U10194 ( .A1(n8612), .A2(keyinput26), .B1(n7676), .B2(keyinput74), 
        .ZN(n8611) );
  OAI221_X1 U10195 ( .B1(n8612), .B2(keyinput26), .C1(n7676), .C2(keyinput74), 
        .A(n8611), .ZN(n8618) );
  AOI22_X1 U10196 ( .A1(n5637), .A2(keyinput32), .B1(n8614), .B2(keyinput7), 
        .ZN(n8613) );
  OAI221_X1 U10197 ( .B1(n5637), .B2(keyinput32), .C1(n8614), .C2(keyinput7), 
        .A(n8613), .ZN(n8617) );
  INV_X1 U10198 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8932) );
  AOI22_X1 U10199 ( .A1(n8795), .A2(keyinput63), .B1(keyinput8), .B2(n8932), 
        .ZN(n8615) );
  OAI221_X1 U10200 ( .B1(n8795), .B2(keyinput63), .C1(n8932), .C2(keyinput8), 
        .A(n8615), .ZN(n8616) );
  OR3_X1 U10201 ( .A1(n8618), .A2(n8617), .A3(n8616), .ZN(n8623) );
  AOI22_X1 U10202 ( .A1(n9180), .A2(keyinput69), .B1(keyinput104), .B2(n6756), 
        .ZN(n8619) );
  OAI221_X1 U10203 ( .B1(n9180), .B2(keyinput69), .C1(n6756), .C2(keyinput104), 
        .A(n8619), .ZN(n8622) );
  INV_X1 U10204 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10558) );
  AOI22_X1 U10205 ( .A1(n6277), .A2(keyinput109), .B1(keyinput80), .B2(n10558), 
        .ZN(n8620) );
  OAI221_X1 U10206 ( .B1(n6277), .B2(keyinput109), .C1(n10558), .C2(keyinput80), .A(n8620), .ZN(n8621) );
  NOR3_X1 U10207 ( .A1(n8623), .A2(n8622), .A3(n8621), .ZN(n8624) );
  AND4_X1 U10208 ( .A1(n8627), .A2(n8626), .A3(n8625), .A4(n8624), .ZN(n8717)
         );
  AOI22_X1 U10209 ( .A1(P2_U3152), .A2(keyinput11), .B1(n8629), .B2(
        keyinput118), .ZN(n8628) );
  OAI221_X1 U10210 ( .B1(P2_U3152), .B2(keyinput11), .C1(n8629), .C2(
        keyinput118), .A(n8628), .ZN(n8640) );
  AOI22_X1 U10211 ( .A1(n8632), .A2(keyinput52), .B1(n8631), .B2(keyinput66), 
        .ZN(n8630) );
  OAI221_X1 U10212 ( .B1(n8632), .B2(keyinput52), .C1(n8631), .C2(keyinput66), 
        .A(n8630), .ZN(n8639) );
  AOI22_X1 U10213 ( .A1(n8635), .A2(keyinput75), .B1(keyinput22), .B2(n8634), 
        .ZN(n8633) );
  OAI221_X1 U10214 ( .B1(n8635), .B2(keyinput75), .C1(n8634), .C2(keyinput22), 
        .A(n8633), .ZN(n8638) );
  AOI22_X1 U10215 ( .A1(n9659), .A2(keyinput5), .B1(keyinput65), .B2(n10520), 
        .ZN(n8636) );
  OAI221_X1 U10216 ( .B1(n9659), .B2(keyinput5), .C1(n10520), .C2(keyinput65), 
        .A(n8636), .ZN(n8637) );
  NOR4_X1 U10217 ( .A1(n8640), .A2(n8639), .A3(n8638), .A4(n8637), .ZN(n8716)
         );
  INV_X1 U10218 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U10219 ( .A1(n10472), .A2(keyinput53), .B1(n8786), .B2(keyinput125), 
        .ZN(n8641) );
  OAI221_X1 U10220 ( .B1(n10472), .B2(keyinput53), .C1(n8786), .C2(keyinput125), .A(n8641), .ZN(n8651) );
  AOI22_X1 U10221 ( .A1(n8643), .A2(keyinput120), .B1(n5203), .B2(keyinput79), 
        .ZN(n8642) );
  OAI221_X1 U10222 ( .B1(n8643), .B2(keyinput120), .C1(n5203), .C2(keyinput79), 
        .A(n8642), .ZN(n8650) );
  INV_X1 U10223 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10443) );
  AOI22_X1 U10224 ( .A1(n10443), .A2(keyinput58), .B1(keyinput27), .B2(n8645), 
        .ZN(n8644) );
  OAI221_X1 U10225 ( .B1(n10443), .B2(keyinput58), .C1(n8645), .C2(keyinput27), 
        .A(n8644), .ZN(n8649) );
  AOI22_X1 U10226 ( .A1(n8647), .A2(keyinput92), .B1(keyinput39), .B2(n9958), 
        .ZN(n8646) );
  OAI221_X1 U10227 ( .B1(n8647), .B2(keyinput92), .C1(n9958), .C2(keyinput39), 
        .A(n8646), .ZN(n8648) );
  NOR4_X1 U10228 ( .A1(n8651), .A2(n8650), .A3(n8649), .A4(n8648), .ZN(n8715)
         );
  INV_X1 U10229 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10445) );
  AOI22_X1 U10230 ( .A1(n8781), .A2(keyinput62), .B1(n10445), .B2(keyinput117), 
        .ZN(n8652) );
  OAI221_X1 U10231 ( .B1(n8781), .B2(keyinput62), .C1(n10445), .C2(keyinput117), .A(n8652), .ZN(n8659) );
  INV_X1 U10232 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10471) );
  INV_X1 U10233 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10442) );
  AOI22_X1 U10234 ( .A1(n10471), .A2(keyinput3), .B1(n10442), .B2(keyinput40), 
        .ZN(n8653) );
  OAI221_X1 U10235 ( .B1(n10471), .B2(keyinput3), .C1(n10442), .C2(keyinput40), 
        .A(n8653), .ZN(n8658) );
  AOI22_X1 U10236 ( .A1(n10358), .A2(keyinput34), .B1(n6253), .B2(keyinput33), 
        .ZN(n8654) );
  OAI221_X1 U10237 ( .B1(n10358), .B2(keyinput34), .C1(n6253), .C2(keyinput33), 
        .A(n8654), .ZN(n8657) );
  INV_X1 U10238 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10447) );
  AOI22_X1 U10239 ( .A1(n9817), .A2(keyinput116), .B1(n10447), .B2(keyinput35), 
        .ZN(n8655) );
  OAI221_X1 U10240 ( .B1(n9817), .B2(keyinput116), .C1(n10447), .C2(keyinput35), .A(n8655), .ZN(n8656) );
  NOR4_X1 U10241 ( .A1(n8659), .A2(n8658), .A3(n8657), .A4(n8656), .ZN(n8713)
         );
  XNOR2_X1 U10242 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput126), .ZN(n8663)
         );
  XNOR2_X1 U10243 ( .A(P2_REG1_REG_29__SCAN_IN), .B(keyinput37), .ZN(n8662) );
  XNOR2_X1 U10244 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput122), .ZN(n8661) );
  XNOR2_X1 U10245 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput64), .ZN(n8660) );
  NAND4_X1 U10246 ( .A1(n8663), .A2(n8662), .A3(n8661), .A4(n8660), .ZN(n8679)
         );
  XNOR2_X1 U10247 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput105), .ZN(n8667) );
  XNOR2_X1 U10248 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput87), .ZN(n8666) );
  XNOR2_X1 U10249 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput97), .ZN(n8665) );
  XNOR2_X1 U10250 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput76), .ZN(n8664) );
  NAND4_X1 U10251 ( .A1(n8667), .A2(n8666), .A3(n8665), .A4(n8664), .ZN(n8678)
         );
  XNOR2_X1 U10252 ( .A(P2_REG2_REG_0__SCAN_IN), .B(keyinput84), .ZN(n8671) );
  XNOR2_X1 U10253 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput48), .ZN(n8670) );
  XNOR2_X1 U10254 ( .A(P1_REG2_REG_1__SCAN_IN), .B(keyinput68), .ZN(n8669) );
  XNOR2_X1 U10255 ( .A(P2_REG0_REG_25__SCAN_IN), .B(keyinput30), .ZN(n8668) );
  NAND4_X1 U10256 ( .A1(n8671), .A2(n8670), .A3(n8669), .A4(n8668), .ZN(n8677)
         );
  XNOR2_X1 U10257 ( .A(SI_30_), .B(keyinput42), .ZN(n8675) );
  XNOR2_X1 U10258 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput25), .ZN(n8674) );
  XNOR2_X1 U10259 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput4), .ZN(n8673) );
  XNOR2_X1 U10260 ( .A(P1_REG2_REG_0__SCAN_IN), .B(keyinput19), .ZN(n8672) );
  NAND4_X1 U10261 ( .A1(n8675), .A2(n8674), .A3(n8673), .A4(n8672), .ZN(n8676)
         );
  NOR4_X1 U10262 ( .A1(n8679), .A2(n8678), .A3(n8677), .A4(n8676), .ZN(n8712)
         );
  AOI22_X1 U10263 ( .A1(n7161), .A2(keyinput72), .B1(n10068), .B2(keyinput100), 
        .ZN(n8680) );
  OAI221_X1 U10264 ( .B1(n7161), .B2(keyinput72), .C1(n10068), .C2(keyinput100), .A(n8680), .ZN(n8692) );
  AOI22_X1 U10265 ( .A1(n8682), .A2(keyinput50), .B1(n8796), .B2(keyinput78), 
        .ZN(n8681) );
  OAI221_X1 U10266 ( .B1(n8682), .B2(keyinput50), .C1(n8796), .C2(keyinput78), 
        .A(n8681), .ZN(n8691) );
  AOI22_X1 U10267 ( .A1(n7976), .A2(keyinput2), .B1(keyinput93), .B2(n8684), 
        .ZN(n8683) );
  OAI221_X1 U10268 ( .B1(n7976), .B2(keyinput2), .C1(n8684), .C2(keyinput93), 
        .A(n8683), .ZN(n8690) );
  XOR2_X1 U10269 ( .A(n8755), .B(keyinput86), .Z(n8688) );
  INV_X1 U10270 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8743) );
  XOR2_X1 U10271 ( .A(n8743), .B(keyinput107), .Z(n8687) );
  XOR2_X1 U10272 ( .A(n8055), .B(keyinput16), .Z(n8686) );
  XNOR2_X1 U10273 ( .A(SI_0_), .B(keyinput1), .ZN(n8685) );
  NAND4_X1 U10274 ( .A1(n8688), .A2(n8687), .A3(n8686), .A4(n8685), .ZN(n8689)
         );
  NOR4_X1 U10275 ( .A1(n8692), .A2(n8691), .A3(n8690), .A4(n8689), .ZN(n8711)
         );
  AOI22_X1 U10276 ( .A1(n8744), .A2(keyinput113), .B1(n8694), .B2(keyinput54), 
        .ZN(n8693) );
  OAI221_X1 U10277 ( .B1(n8744), .B2(keyinput113), .C1(n8694), .C2(keyinput54), 
        .A(n8693), .ZN(n8703) );
  AOI22_X1 U10278 ( .A1(n9256), .A2(keyinput102), .B1(n8696), .B2(keyinput114), 
        .ZN(n8695) );
  OAI221_X1 U10279 ( .B1(n9256), .B2(keyinput102), .C1(n8696), .C2(keyinput114), .A(n8695), .ZN(n8702) );
  AOI22_X1 U10280 ( .A1(n8764), .A2(keyinput123), .B1(n9796), .B2(keyinput108), 
        .ZN(n8697) );
  OAI221_X1 U10281 ( .B1(n8764), .B2(keyinput123), .C1(n9796), .C2(keyinput108), .A(n8697), .ZN(n8701) );
  AOI22_X1 U10282 ( .A1(n8699), .A2(keyinput49), .B1(n8782), .B2(keyinput112), 
        .ZN(n8698) );
  OAI221_X1 U10283 ( .B1(n8699), .B2(keyinput49), .C1(n8782), .C2(keyinput112), 
        .A(n8698), .ZN(n8700) );
  OR4_X1 U10284 ( .A1(n8703), .A2(n8702), .A3(n8701), .A4(n8700), .ZN(n8709)
         );
  AOI22_X1 U10285 ( .A1(n8766), .A2(keyinput61), .B1(n8705), .B2(keyinput55), 
        .ZN(n8704) );
  OAI221_X1 U10286 ( .B1(n8766), .B2(keyinput61), .C1(n8705), .C2(keyinput55), 
        .A(n8704), .ZN(n8708) );
  INV_X1 U10287 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10440) );
  AOI22_X1 U10288 ( .A1(n10440), .A2(keyinput88), .B1(keyinput111), .B2(n5867), 
        .ZN(n8706) );
  OAI221_X1 U10289 ( .B1(n10440), .B2(keyinput88), .C1(n5867), .C2(keyinput111), .A(n8706), .ZN(n8707) );
  NOR3_X1 U10290 ( .A1(n8709), .A2(n8708), .A3(n8707), .ZN(n8710) );
  AND4_X1 U10291 ( .A1(n8713), .A2(n8712), .A3(n8711), .A4(n8710), .ZN(n8714)
         );
  AND4_X1 U10292 ( .A1(n8717), .A2(n8716), .A3(n8715), .A4(n8714), .ZN(n8814)
         );
  INV_X1 U10293 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10469) );
  AOI22_X1 U10294 ( .A1(n10527), .A2(keyinput23), .B1(n10469), .B2(keyinput115), .ZN(n8718) );
  OAI221_X1 U10295 ( .B1(n10527), .B2(keyinput23), .C1(n10469), .C2(
        keyinput115), .A(n8718), .ZN(n8726) );
  INV_X1 U10296 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10430) );
  AOI22_X1 U10297 ( .A1(n8720), .A2(keyinput28), .B1(keyinput124), .B2(n10430), 
        .ZN(n8719) );
  OAI221_X1 U10298 ( .B1(n8720), .B2(keyinput28), .C1(n10430), .C2(keyinput124), .A(n8719), .ZN(n8725) );
  INV_X1 U10299 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10441) );
  INV_X1 U10300 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8741) );
  AOI22_X1 U10301 ( .A1(n10441), .A2(keyinput82), .B1(keyinput6), .B2(n8741), 
        .ZN(n8721) );
  OAI221_X1 U10302 ( .B1(n10441), .B2(keyinput82), .C1(n8741), .C2(keyinput6), 
        .A(n8721), .ZN(n8724) );
  INV_X1 U10303 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n10470) );
  AOI22_X1 U10304 ( .A1(n10470), .A2(keyinput110), .B1(keyinput51), .B2(n5259), 
        .ZN(n8722) );
  OAI221_X1 U10305 ( .B1(n10470), .B2(keyinput110), .C1(n5259), .C2(keyinput51), .A(n8722), .ZN(n8723) );
  NOR4_X1 U10306 ( .A1(n8726), .A2(n8725), .A3(n8724), .A4(n8723), .ZN(n8813)
         );
  AOI22_X1 U10307 ( .A1(n8728), .A2(keyinput67), .B1(keyinput46), .B2(n8789), 
        .ZN(n8727) );
  OAI221_X1 U10308 ( .B1(n8728), .B2(keyinput67), .C1(n8789), .C2(keyinput46), 
        .A(n8727), .ZN(n8738) );
  AOI22_X1 U10309 ( .A1(n8731), .A2(keyinput24), .B1(n8730), .B2(keyinput38), 
        .ZN(n8729) );
  OAI221_X1 U10310 ( .B1(n8731), .B2(keyinput24), .C1(n8730), .C2(keyinput38), 
        .A(n8729), .ZN(n8737) );
  AOI22_X1 U10311 ( .A1(n8733), .A2(keyinput10), .B1(keyinput47), .B2(n8912), 
        .ZN(n8732) );
  OAI221_X1 U10312 ( .B1(n8733), .B2(keyinput10), .C1(n8912), .C2(keyinput47), 
        .A(n8732), .ZN(n8736) );
  AOI22_X1 U10313 ( .A1(n8788), .A2(keyinput29), .B1(keyinput81), .B2(n10345), 
        .ZN(n8734) );
  OAI221_X1 U10314 ( .B1(n8788), .B2(keyinput29), .C1(n10345), .C2(keyinput81), 
        .A(n8734), .ZN(n8735) );
  NOR4_X1 U10315 ( .A1(n8738), .A2(n8737), .A3(n8736), .A4(n8735), .ZN(n8812)
         );
  NAND4_X1 U10316 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_REG3_REG_0__SCAN_IN), 
        .A3(P2_REG3_REG_24__SCAN_IN), .A4(P2_REG3_REG_17__SCAN_IN), .ZN(n8739)
         );
  NOR3_X1 U10317 ( .A1(P2_REG2_REG_28__SCAN_IN), .A2(n7676), .A3(n8739), .ZN(
        n8752) );
  NAND4_X1 U10318 ( .A1(n8740), .A2(P1_IR_REG_10__SCAN_IN), .A3(
        P2_ADDR_REG_3__SCAN_IN), .A4(n6661), .ZN(n8750) );
  NOR4_X1 U10319 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .A3(P1_ADDR_REG_10__SCAN_IN), .A4(n8741), .ZN(n8748) );
  NOR4_X1 U10320 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_1__SCAN_IN), 
        .A3(P1_ADDR_REG_18__SCAN_IN), .A4(n6277), .ZN(n8747) );
  NOR4_X1 U10321 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(n10473), .A3(n9029), .A4(
        n8742), .ZN(n8746) );
  NOR4_X1 U10322 ( .A1(P1_REG0_REG_8__SCAN_IN), .A2(P2_REG0_REG_24__SCAN_IN), 
        .A3(n8744), .A4(n8743), .ZN(n8745) );
  NAND4_X1 U10323 ( .A1(n8748), .A2(n8747), .A3(n8746), .A4(n8745), .ZN(n8749)
         );
  NOR4_X1 U10324 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        n8750), .A4(n8749), .ZN(n8751) );
  NAND4_X1 U10325 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .A3(n8752), .A4(n8751), .ZN(n8808) );
  INV_X1 U10326 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n8754) );
  NOR4_X1 U10327 ( .A1(n8754), .A2(P2_U3152), .A3(n8753), .A4(
        P2_IR_REG_24__SCAN_IN), .ZN(n8762) );
  NOR4_X1 U10328 ( .A1(n8757), .A2(n8756), .A3(n8755), .A4(
        P1_REG1_REG_29__SCAN_IN), .ZN(n8761) );
  NOR4_X1 U10329 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG0_REG_25__SCAN_IN), 
        .A3(P2_REG0_REG_8__SCAN_IN), .A4(P2_REG1_REG_13__SCAN_IN), .ZN(n8760)
         );
  NOR4_X1 U10330 ( .A1(n8758), .A2(n5676), .A3(P1_D_REG_27__SCAN_IN), .A4(
        P2_D_REG_15__SCAN_IN), .ZN(n8759) );
  NAND4_X1 U10331 ( .A1(n8762), .A2(n8761), .A3(n8760), .A4(n8759), .ZN(n8780)
         );
  NOR4_X1 U10332 ( .A1(n8763), .A2(P1_IR_REG_8__SCAN_IN), .A3(SI_11_), .A4(
        SI_0_), .ZN(n8775) );
  NOR4_X1 U10333 ( .A1(n4642), .A2(P1_IR_REG_23__SCAN_IN), .A3(
        P1_REG2_REG_11__SCAN_IN), .A4(P1_REG0_REG_26__SCAN_IN), .ZN(n8774) );
  NOR4_X1 U10334 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(n8764), .A3(n9796), .A4(
        n8055), .ZN(n8770) );
  NOR4_X1 U10335 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(P2_DATAO_REG_0__SCAN_IN), 
        .A3(n8766), .A4(n8765), .ZN(n8769) );
  NOR4_X1 U10336 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(P1_DATAO_REG_15__SCAN_IN), .A3(P1_REG0_REG_19__SCAN_IN), .A4(P2_REG1_REG_25__SCAN_IN), .ZN(n8768) );
  NOR4_X1 U10337 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG1_REG_25__SCAN_IN), 
        .A3(P2_REG1_REG_7__SCAN_IN), .A4(n9659), .ZN(n8767) );
  NAND4_X1 U10338 ( .A1(n8770), .A2(n8769), .A3(n8768), .A4(n8767), .ZN(n8771)
         );
  NOR3_X1 U10339 ( .A1(n10442), .A2(SI_19_), .A3(n8771), .ZN(n8772) );
  NAND4_X1 U10340 ( .A1(n8775), .A2(n8774), .A3(n8773), .A4(n8772), .ZN(n8779)
         );
  NOR4_X1 U10341 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P1_REG0_REG_25__SCAN_IN), 
        .A3(P2_REG2_REG_3__SCAN_IN), .A4(n8776), .ZN(n8777) );
  NAND3_X1 U10342 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(SI_15_), .A3(n8777), .ZN(
        n8778) );
  NOR3_X1 U10343 ( .A1(n8780), .A2(n8779), .A3(n8778), .ZN(n8785) );
  NAND4_X1 U10344 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_REG0_REG_27__SCAN_IN), 
        .A3(n8782), .A4(n8781), .ZN(n8783) );
  NOR3_X1 U10345 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .A3(
        n8783), .ZN(n8784) );
  NAND2_X1 U10346 ( .A1(n8785), .A2(n8784), .ZN(n8807) );
  NAND4_X1 U10347 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_REG2_REG_23__SCAN_IN), 
        .A3(n8786), .A4(n9958), .ZN(n8793) );
  NAND4_X1 U10348 ( .A1(P1_REG1_REG_30__SCAN_IN), .A2(n8787), .A3(n9487), .A4(
        n5203), .ZN(n8792) );
  NAND4_X1 U10349 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(SI_5_), .A3(
        P2_DATAO_REG_30__SCAN_IN), .A4(n8788), .ZN(n8791) );
  NAND4_X1 U10350 ( .A1(P1_REG0_REG_11__SCAN_IN), .A2(P1_DATAO_REG_20__SCAN_IN), .A3(P2_REG1_REG_9__SCAN_IN), .A4(n8789), .ZN(n8790) );
  OR4_X1 U10351 ( .A1(n8793), .A2(n8792), .A3(n8791), .A4(n8790), .ZN(n8806)
         );
  NAND4_X1 U10352 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(P1_REG1_REG_6__SCAN_IN), 
        .A3(P1_REG1_REG_1__SCAN_IN), .A4(P2_REG3_REG_5__SCAN_IN), .ZN(n8794)
         );
  NOR3_X1 U10353 ( .A1(P2_REG1_REG_24__SCAN_IN), .A2(n8795), .A3(n8794), .ZN(
        n8804) );
  NAND4_X1 U10354 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), 
        .A3(P2_REG3_REG_9__SCAN_IN), .A4(n7976), .ZN(n8802) );
  NAND4_X1 U10355 ( .A1(P1_REG2_REG_20__SCAN_IN), .A2(P1_REG2_REG_9__SCAN_IN), 
        .A3(n8797), .A4(n8796), .ZN(n8798) );
  NOR2_X1 U10356 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(n8798), .ZN(n8799) );
  NAND4_X1 U10357 ( .A1(n8799), .A2(P2_REG3_REG_10__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n8801) );
  NAND4_X1 U10358 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_REG3_REG_26__SCAN_IN), 
        .A3(P1_REG0_REG_10__SCAN_IN), .A4(P2_REG1_REG_6__SCAN_IN), .ZN(n8800)
         );
  NOR3_X1 U10359 ( .A1(n8802), .A2(n8801), .A3(n8800), .ZN(n8803) );
  NAND4_X1 U10360 ( .A1(SI_20_), .A2(P1_DATAO_REG_30__SCAN_IN), .A3(n8804), 
        .A4(n8803), .ZN(n8805) );
  NOR4_X1 U10361 ( .A1(n8808), .A2(n8807), .A3(n8806), .A4(n8805), .ZN(n8810)
         );
  INV_X1 U10362 ( .A(keyinput12), .ZN(n8809) );
  OAI21_X1 U10363 ( .B1(n8810), .B2(P1_IR_REG_21__SCAN_IN), .A(n8809), .ZN(
        n8811) );
  NAND4_X1 U10364 ( .A1(n8814), .A2(n8813), .A3(n8812), .A4(n8811), .ZN(n8815)
         );
  OAI21_X1 U10365 ( .B1(n8818), .B2(n8817), .A(n8816), .ZN(n8820) );
  AOI22_X1 U10366 ( .A1(n9105), .A2(n8820), .B1(n8819), .B2(n9177), .ZN(n8824)
         );
  AOI22_X1 U10367 ( .A1(n8822), .A2(n6045), .B1(n8821), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n8823) );
  OAI211_X1 U10368 ( .C1(n8825), .C2(n9153), .A(n8824), .B(n8823), .ZN(
        P2_U3239) );
  OAI22_X1 U10369 ( .A1(n8828), .A2(n8827), .B1(n8826), .B2(n9485), .ZN(n8829)
         );
  AOI21_X1 U10370 ( .B1(n4374), .B2(P2_REG2_REG_4__SCAN_IN), .A(n8829), .ZN(
        n8833) );
  AOI22_X1 U10371 ( .A1(n9522), .A2(n8831), .B1(n9536), .B2(n8830), .ZN(n8832)
         );
  OAI211_X1 U10372 ( .C1(n8834), .C2(n9437), .A(n8833), .B(n8832), .ZN(
        P2_U3292) );
  XNOR2_X1 U10373 ( .A(n9580), .B(n8882), .ZN(n9100) );
  NAND2_X1 U10374 ( .A1(n9162), .A2(n8835), .ZN(n9104) );
  NAND2_X1 U10375 ( .A1(n9100), .A2(n9104), .ZN(n8855) );
  INV_X1 U10376 ( .A(n8855), .ZN(n8843) );
  XNOR2_X1 U10377 ( .A(n9414), .B(n8872), .ZN(n8848) );
  NAND2_X1 U10378 ( .A1(n9163), .A2(n8835), .ZN(n8844) );
  XNOR2_X1 U10379 ( .A(n8848), .B(n8844), .ZN(n9002) );
  XNOR2_X1 U10380 ( .A(n9433), .B(n8868), .ZN(n8837) );
  NOR2_X1 U10381 ( .A1(n9004), .A2(n8880), .ZN(n8836) );
  NAND2_X1 U10382 ( .A1(n8837), .A2(n8836), .ZN(n8842) );
  XNOR2_X1 U10383 ( .A(n8837), .B(n8836), .ZN(n9071) );
  INV_X1 U10384 ( .A(n8839), .ZN(n8840) );
  NOR2_X1 U10385 ( .A1(n8841), .A2(n8840), .ZN(n9068) );
  NOR2_X1 U10386 ( .A1(n9108), .A2(n8880), .ZN(n8860) );
  XNOR2_X1 U10387 ( .A(n9383), .B(n8872), .ZN(n8859) );
  INV_X1 U10388 ( .A(n9100), .ZN(n8846) );
  INV_X1 U10389 ( .A(n8844), .ZN(n8847) );
  NAND2_X1 U10390 ( .A1(n8848), .A2(n8847), .ZN(n9097) );
  NAND2_X1 U10391 ( .A1(n9097), .A2(n9104), .ZN(n8845) );
  NAND2_X1 U10392 ( .A1(n8846), .A2(n8845), .ZN(n8850) );
  NAND3_X1 U10393 ( .A1(n8848), .A2(n8847), .A3(n9162), .ZN(n8849) );
  NAND2_X1 U10394 ( .A1(n8850), .A2(n8849), .ZN(n8988) );
  AOI21_X1 U10395 ( .B1(n8860), .B2(n8859), .A(n8988), .ZN(n8851) );
  AND2_X1 U10396 ( .A1(n8852), .A2(n8853), .ZN(n8857) );
  INV_X1 U10397 ( .A(n8853), .ZN(n8856) );
  AND2_X1 U10398 ( .A1(n9114), .A2(n8854), .ZN(n8999) );
  AND2_X1 U10399 ( .A1(n8999), .A2(n9002), .ZN(n9093) );
  AND2_X1 U10400 ( .A1(n9093), .A2(n8855), .ZN(n8985) );
  XNOR2_X1 U10401 ( .A(n9570), .B(n8882), .ZN(n9060) );
  NAND2_X1 U10402 ( .A1(n9160), .A2(n8835), .ZN(n8861) );
  INV_X1 U10403 ( .A(n8859), .ZN(n8991) );
  INV_X1 U10404 ( .A(n8860), .ZN(n8995) );
  AND2_X1 U10405 ( .A1(n8991), .A2(n8995), .ZN(n9057) );
  AOI21_X1 U10406 ( .B1(n9060), .B2(n8861), .A(n9057), .ZN(n8864) );
  INV_X1 U10407 ( .A(n9060), .ZN(n8862) );
  INV_X1 U10408 ( .A(n8861), .ZN(n9062) );
  AND2_X1 U10409 ( .A1(n8862), .A2(n9062), .ZN(n8863) );
  XNOR2_X1 U10410 ( .A(n9566), .B(n8882), .ZN(n8865) );
  NOR2_X1 U10411 ( .A1(n9128), .A2(n8880), .ZN(n9025) );
  INV_X1 U10412 ( .A(n8865), .ZN(n9026) );
  INV_X1 U10413 ( .A(n9028), .ZN(n8866) );
  XNOR2_X1 U10414 ( .A(n9345), .B(n8868), .ZN(n8897) );
  NOR2_X1 U10415 ( .A1(n8869), .A2(n8880), .ZN(n8870) );
  NAND2_X1 U10416 ( .A1(n8897), .A2(n8870), .ZN(n8871) );
  OAI21_X1 U10417 ( .B1(n8897), .B2(n8870), .A(n8871), .ZN(n9127) );
  INV_X1 U10418 ( .A(n8871), .ZN(n8878) );
  XNOR2_X1 U10419 ( .A(n9326), .B(n8872), .ZN(n8873) );
  NOR2_X1 U10420 ( .A1(n9129), .A2(n8880), .ZN(n8874) );
  NAND2_X1 U10421 ( .A1(n8873), .A2(n8874), .ZN(n8879) );
  INV_X1 U10422 ( .A(n8873), .ZN(n8876) );
  INV_X1 U10423 ( .A(n8874), .ZN(n8875) );
  NAND2_X1 U10424 ( .A1(n8876), .A2(n8875), .ZN(n8877) );
  NOR2_X1 U10425 ( .A1(n8881), .A2(n8880), .ZN(n8883) );
  XNOR2_X1 U10426 ( .A(n8883), .B(n8882), .ZN(n8886) );
  NOR3_X1 U10427 ( .A1(n5001), .A2(n8886), .A3(n9122), .ZN(n8884) );
  AOI21_X1 U10428 ( .B1(n5001), .B2(n8886), .A(n8884), .ZN(n8890) );
  NAND3_X1 U10429 ( .A1(n9548), .A2(n9153), .A3(n8886), .ZN(n8885) );
  OAI21_X1 U10430 ( .B1(n9548), .B2(n8886), .A(n8885), .ZN(n8887) );
  NAND2_X1 U10431 ( .A1(n8891), .A2(n8887), .ZN(n8889) );
  OAI21_X1 U10432 ( .B1(n5001), .B2(n9153), .A(n9138), .ZN(n8888) );
  OAI211_X1 U10433 ( .C1(n8891), .C2(n8890), .A(n8889), .B(n8888), .ZN(n8894)
         );
  AOI22_X1 U10434 ( .A1(n8892), .A2(n9143), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8893) );
  OAI211_X1 U10435 ( .C1(n8895), .C2(n9073), .A(n8894), .B(n8893), .ZN(
        P2_U3222) );
  AOI22_X1 U10436 ( .A1(n9157), .A2(n9464), .B1(n9462), .B2(n9159), .ZN(n9321)
         );
  AOI22_X1 U10437 ( .A1(n9327), .A2(n9143), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8896) );
  OAI21_X1 U10438 ( .B1(n9321), .B2(n9073), .A(n8896), .ZN(n8901) );
  NAND3_X1 U10439 ( .A1(n8897), .A2(n9102), .A3(n9159), .ZN(n8900) );
  OR2_X1 U10440 ( .A1(n8902), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8903) );
  NAND2_X1 U10441 ( .A1(n8904), .A2(n8903), .ZN(n9278) );
  XNOR2_X1 U10442 ( .A(n8908), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n9279) );
  NAND2_X1 U10443 ( .A1(n8908), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8905) );
  NAND2_X1 U10444 ( .A1(n9276), .A2(n8905), .ZN(n9284) );
  XNOR2_X1 U10445 ( .A(n8913), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n9285) );
  OR2_X1 U10446 ( .A1(n9284), .A2(n9285), .ZN(n9282) );
  OR2_X1 U10447 ( .A1(n8913), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8906) );
  NAND2_X1 U10448 ( .A1(n9282), .A2(n8906), .ZN(n8907) );
  XNOR2_X1 U10449 ( .A(n8907), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8919) );
  AOI22_X1 U10450 ( .A1(n8908), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8912), .B2(
        n9275), .ZN(n9269) );
  NAND2_X1 U10451 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n9292), .ZN(n9290) );
  NAND2_X1 U10452 ( .A1(n8914), .A2(n8913), .ZN(n8915) );
  NAND2_X1 U10453 ( .A1(n9290), .A2(n8915), .ZN(n8917) );
  XOR2_X1 U10454 ( .A(n8917), .B(n8916), .Z(n8922) );
  NAND2_X1 U10455 ( .A1(n8922), .A2(n9291), .ZN(n8918) );
  OAI211_X1 U10456 ( .C1(n8919), .C2(n9295), .A(n8918), .B(n9286), .ZN(n8925)
         );
  INV_X1 U10457 ( .A(n8919), .ZN(n8920) );
  OAI22_X1 U10458 ( .A1(n8922), .A2(n8921), .B1(n8920), .B2(n9295), .ZN(n8924)
         );
  NAND2_X1 U10459 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8926) );
  OAI222_X1 U10460 ( .A1(n10350), .A2(n8930), .B1(P1_U3084), .B2(n8929), .C1(
        n10347), .C2(n8928), .ZN(P1_U3325) );
  INV_X1 U10461 ( .A(n8931), .ZN(n10344) );
  NAND2_X1 U10462 ( .A1(n10207), .A2(n8934), .ZN(n8937) );
  NAND2_X1 U10463 ( .A1(n9966), .A2(n8935), .ZN(n8936) );
  NAND2_X1 U10464 ( .A1(n8937), .A2(n8936), .ZN(n8939) );
  XNOR2_X1 U10465 ( .A(n8939), .B(n8938), .ZN(n8945) );
  NAND2_X1 U10466 ( .A1(n10207), .A2(n8940), .ZN(n8941) );
  OAI21_X1 U10467 ( .B1(n8943), .B2(n8942), .A(n8941), .ZN(n8944) );
  XNOR2_X1 U10468 ( .A(n8945), .B(n8944), .ZN(n8946) );
  INV_X1 U10469 ( .A(n8946), .ZN(n8952) );
  NAND3_X1 U10470 ( .A1(n8952), .A2(n9815), .A3(n8951), .ZN(n8957) );
  INV_X1 U10471 ( .A(n8947), .ZN(n9841) );
  AOI22_X1 U10472 ( .A1(n9841), .A2(n9835), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8950) );
  NAND2_X1 U10473 ( .A1(n8948), .A2(n9773), .ZN(n8949) );
  OAI211_X1 U10474 ( .C1(n9994), .C2(n9831), .A(n8950), .B(n8949), .ZN(n8954)
         );
  NOR3_X1 U10475 ( .A1(n8952), .A2(n8951), .A3(n9825), .ZN(n8953) );
  AOI211_X1 U10476 ( .C1(n10207), .C2(n4582), .A(n8954), .B(n8953), .ZN(n8955)
         );
  OAI211_X1 U10477 ( .C1(n8958), .C2(n8957), .A(n8956), .B(n8955), .ZN(
        P1_U3218) );
  INV_X1 U10478 ( .A(n8959), .ZN(n8963) );
  OAI222_X1 U10479 ( .A1(n10350), .A2(n8961), .B1(n10347), .B2(n8963), .C1(
        n4372), .C2(P1_U3084), .ZN(P1_U3331) );
  OAI222_X1 U10480 ( .A1(n9686), .A2(n8965), .B1(n8964), .B2(n8963), .C1(
        P2_U3152), .C2(n8962), .ZN(P2_U3336) );
  INV_X1 U10481 ( .A(n8966), .ZN(n8969) );
  NOR3_X1 U10482 ( .A1(n9136), .A2(n8967), .A3(n8975), .ZN(n8968) );
  AOI21_X1 U10483 ( .B1(n8969), .B2(n9105), .A(n8968), .ZN(n8982) );
  NOR2_X1 U10484 ( .A1(n8970), .A2(n9138), .ZN(n8979) );
  NOR2_X1 U10485 ( .A1(n9153), .A2(n8971), .ZN(n8978) );
  OAI21_X1 U10486 ( .B1(n9148), .B2(n9137), .A(n8972), .ZN(n8977) );
  NAND2_X1 U10487 ( .A1(n9143), .A2(n8973), .ZN(n8974) );
  OAI21_X1 U10488 ( .B1(n8975), .B2(n9145), .A(n8974), .ZN(n8976) );
  NOR4_X1 U10489 ( .A1(n8979), .A2(n8978), .A3(n8977), .A4(n8976), .ZN(n8980)
         );
  OAI21_X1 U10490 ( .B1(n8982), .B2(n8981), .A(n8980), .ZN(P2_U3217) );
  OAI22_X1 U10491 ( .A1(n8983), .A2(n9528), .B1(n9005), .B2(n9531), .ZN(n9392)
         );
  AOI22_X1 U10492 ( .A1(n9392), .A2(n9133), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8984) );
  OAI21_X1 U10493 ( .B1(n9384), .B2(n9131), .A(n8984), .ZN(n8994) );
  NAND2_X1 U10494 ( .A1(n9094), .A2(n8985), .ZN(n8987) );
  AND2_X1 U10495 ( .A1(n8987), .A2(n8986), .ZN(n8990) );
  INV_X1 U10496 ( .A(n8988), .ZN(n8989) );
  NAND2_X1 U10497 ( .A1(n8990), .A2(n8989), .ZN(n8992) );
  XNOR2_X1 U10498 ( .A(n8992), .B(n8991), .ZN(n8996) );
  NOR3_X1 U10499 ( .A1(n8996), .A2(n9108), .A3(n9136), .ZN(n8993) );
  AOI211_X1 U10500 ( .C1(n9383), .C2(n9122), .A(n8994), .B(n8993), .ZN(n8998)
         );
  NAND3_X1 U10501 ( .A1(n8996), .A2(n9105), .A3(n8995), .ZN(n8997) );
  NAND2_X1 U10502 ( .A1(n8998), .A2(n8997), .ZN(P2_U3218) );
  NAND2_X1 U10503 ( .A1(n9094), .A2(n8999), .ZN(n9001) );
  NAND2_X1 U10504 ( .A1(n9001), .A2(n9000), .ZN(n9003) );
  XNOR2_X1 U10505 ( .A(n9003), .B(n9002), .ZN(n9009) );
  OAI22_X1 U10506 ( .A1(n9005), .A2(n9528), .B1(n9004), .B2(n9531), .ZN(n9425)
         );
  AOI22_X1 U10507 ( .A1(n9425), .A2(n9133), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n9006) );
  OAI21_X1 U10508 ( .B1(n9415), .B2(n9131), .A(n9006), .ZN(n9007) );
  AOI21_X1 U10509 ( .B1(n9414), .B2(n9122), .A(n9007), .ZN(n9008) );
  OAI21_X1 U10510 ( .B1(n9009), .B2(n9138), .A(n9008), .ZN(P2_U3225) );
  INV_X1 U10511 ( .A(n9010), .ZN(n9011) );
  AOI21_X1 U10512 ( .B1(n9012), .B2(n9011), .A(n9138), .ZN(n9017) );
  NOR3_X1 U10513 ( .A1(n9136), .A2(n9014), .A3(n9013), .ZN(n9016) );
  OAI21_X1 U10514 ( .B1(n9017), .B2(n9016), .A(n9015), .ZN(n9024) );
  AOI22_X1 U10515 ( .A1(n9133), .A2(n9018), .B1(P2_REG3_REG_12__SCAN_IN), .B2(
        P2_U3152), .ZN(n9023) );
  OR2_X1 U10516 ( .A1(n9153), .A2(n9019), .ZN(n9022) );
  NAND2_X1 U10517 ( .A1(n9143), .A2(n9020), .ZN(n9021) );
  NAND4_X1 U10518 ( .A1(n9024), .A2(n9023), .A3(n9022), .A4(n9021), .ZN(
        P2_U3226) );
  XNOR2_X1 U10519 ( .A(n9026), .B(n9025), .ZN(n9027) );
  XNOR2_X1 U10520 ( .A(n9028), .B(n9027), .ZN(n9034) );
  AOI22_X1 U10521 ( .A1(n9159), .A2(n9464), .B1(n9462), .B2(n9160), .ZN(n9354)
         );
  OAI22_X1 U10522 ( .A1(n9354), .A2(n9073), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9029), .ZN(n9032) );
  NOR2_X1 U10523 ( .A1(n9030), .A2(n9153), .ZN(n9031) );
  AOI211_X1 U10524 ( .C1(n9143), .C2(n9357), .A(n9032), .B(n9031), .ZN(n9033)
         );
  OAI21_X1 U10525 ( .B1(n9034), .B2(n9138), .A(n9033), .ZN(P2_U3227) );
  XNOR2_X1 U10526 ( .A(n9037), .B(n9035), .ZN(n9135) );
  NAND2_X1 U10527 ( .A1(n9135), .A2(n9036), .ZN(n9140) );
  OAI21_X1 U10528 ( .B1(n9038), .B2(n9037), .A(n9140), .ZN(n9042) );
  XNOR2_X1 U10529 ( .A(n9040), .B(n9039), .ZN(n9041) );
  XNOR2_X1 U10530 ( .A(n9042), .B(n9041), .ZN(n9049) );
  AOI22_X1 U10531 ( .A1(n9133), .A2(n9043), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3152), .ZN(n9044) );
  OAI21_X1 U10532 ( .B1(n9131), .B2(n9045), .A(n9044), .ZN(n9046) );
  AOI21_X1 U10533 ( .B1(n9047), .B2(n9122), .A(n9046), .ZN(n9048) );
  OAI21_X1 U10534 ( .B1(n9049), .B2(n9138), .A(n9048), .ZN(P2_U3228) );
  INV_X1 U10535 ( .A(n9512), .ZN(n9607) );
  OAI211_X1 U10536 ( .C1(n9051), .C2(n9050), .A(n8858), .B(n9105), .ZN(n9055)
         );
  NOR2_X1 U10537 ( .A1(n9145), .A2(n9499), .ZN(n9053) );
  OAI22_X1 U10538 ( .A1(n9148), .A2(n9500), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9271), .ZN(n9052) );
  AOI211_X1 U10539 ( .C1(n9143), .C2(n9511), .A(n9053), .B(n9052), .ZN(n9054)
         );
  OAI211_X1 U10540 ( .C1(n9607), .C2(n9153), .A(n9055), .B(n9054), .ZN(
        P2_U3230) );
  OAI22_X1 U10541 ( .A1(n9128), .A2(n9528), .B1(n9108), .B2(n9531), .ZN(n9364)
         );
  AOI22_X1 U10542 ( .A1(n9364), .A2(n9133), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n9056) );
  OAI21_X1 U10543 ( .B1(n9368), .B2(n9131), .A(n9056), .ZN(n9064) );
  INV_X1 U10544 ( .A(n9057), .ZN(n9058) );
  NAND2_X1 U10545 ( .A1(n9059), .A2(n9058), .ZN(n9061) );
  XNOR2_X1 U10546 ( .A(n9061), .B(n9060), .ZN(n9065) );
  NOR3_X1 U10547 ( .A1(n9065), .A2(n9062), .A3(n9138), .ZN(n9063) );
  AOI211_X1 U10548 ( .C1(n9570), .C2(n9122), .A(n9064), .B(n9063), .ZN(n9067)
         );
  NAND3_X1 U10549 ( .A1(n9065), .A2(n9102), .A3(n9160), .ZN(n9066) );
  NAND2_X1 U10550 ( .A1(n9067), .A2(n9066), .ZN(P2_U3231) );
  NAND2_X1 U10551 ( .A1(n9068), .A2(n9117), .ZN(n9070) );
  NAND2_X1 U10552 ( .A1(n9070), .A2(n9069), .ZN(n9072) );
  XNOR2_X1 U10553 ( .A(n9072), .B(n9071), .ZN(n9077) );
  NOR2_X1 U10554 ( .A1(n9131), .A2(n9434), .ZN(n9075) );
  AOI22_X1 U10555 ( .A1(n9163), .A2(n9464), .B1(n9164), .B2(n9462), .ZN(n9441)
         );
  OAI22_X1 U10556 ( .A1(n9073), .A2(n9441), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n4654), .ZN(n9074) );
  AOI211_X1 U10557 ( .C1(n9433), .C2(n9122), .A(n9075), .B(n9074), .ZN(n9076)
         );
  OAI21_X1 U10558 ( .B1(n9077), .B2(n9138), .A(n9076), .ZN(P2_U3235) );
  INV_X1 U10559 ( .A(n9078), .ZN(n9079) );
  AOI21_X1 U10560 ( .B1(n9015), .B2(n9079), .A(n9138), .ZN(n9082) );
  NOR3_X1 U10561 ( .A1(n9136), .A2(n9086), .A3(n9080), .ZN(n9081) );
  OAI21_X1 U10562 ( .B1(n9082), .B2(n9081), .A(n8966), .ZN(n9091) );
  INV_X1 U10563 ( .A(n9083), .ZN(n9084) );
  NAND2_X1 U10564 ( .A1(n9143), .A2(n9084), .ZN(n9085) );
  OAI21_X1 U10565 ( .B1(n9086), .B2(n9145), .A(n9085), .ZN(n9089) );
  OAI21_X1 U10566 ( .B1(n9148), .B2(n9146), .A(n9087), .ZN(n9088) );
  NOR2_X1 U10567 ( .A1(n9089), .A2(n9088), .ZN(n9090) );
  OAI211_X1 U10568 ( .C1(n9092), .C2(n9153), .A(n9091), .B(n9090), .ZN(
        P2_U3236) );
  NAND2_X1 U10569 ( .A1(n9094), .A2(n9093), .ZN(n9096) );
  NAND2_X1 U10570 ( .A1(n9096), .A2(n9095), .ZN(n9099) );
  INV_X1 U10571 ( .A(n9097), .ZN(n9098) );
  NOR2_X1 U10572 ( .A1(n9099), .A2(n9098), .ZN(n9101) );
  XNOR2_X1 U10573 ( .A(n9101), .B(n9100), .ZN(n9103) );
  NAND3_X1 U10574 ( .A1(n9103), .A2(n9102), .A3(n9162), .ZN(n9113) );
  INV_X1 U10575 ( .A(n9103), .ZN(n9106) );
  NAND3_X1 U10576 ( .A1(n9106), .A2(n9105), .A3(n9104), .ZN(n9112) );
  OAI22_X1 U10577 ( .A1(n9108), .A2(n9528), .B1(n9107), .B2(n9531), .ZN(n9406)
         );
  AOI22_X1 U10578 ( .A1(n9406), .A2(n9133), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n9109) );
  OAI21_X1 U10579 ( .B1(n9403), .B2(n9131), .A(n9109), .ZN(n9110) );
  AOI21_X1 U10580 ( .B1(n9580), .B2(n9122), .A(n9110), .ZN(n9111) );
  NAND3_X1 U10581 ( .A1(n9113), .A2(n9112), .A3(n9111), .ZN(P2_U3237) );
  INV_X1 U10582 ( .A(n9114), .ZN(n9115) );
  AOI21_X1 U10583 ( .B1(n8858), .B2(n9115), .A(n9138), .ZN(n9119) );
  NOR3_X1 U10584 ( .A1(n9116), .A2(n9479), .A3(n9136), .ZN(n9118) );
  OAI21_X1 U10585 ( .B1(n9119), .B2(n9118), .A(n9117), .ZN(n9124) );
  OAI22_X1 U10586 ( .A1(n9148), .A2(n9480), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n4653), .ZN(n9121) );
  OAI22_X1 U10587 ( .A1(n9131), .A2(n9486), .B1(n9479), .B2(n9145), .ZN(n9120)
         );
  AOI211_X1 U10588 ( .C1(n9489), .C2(n9122), .A(n9121), .B(n9120), .ZN(n9123)
         );
  NAND2_X1 U10589 ( .A1(n9124), .A2(n9123), .ZN(P2_U3240) );
  OAI22_X1 U10590 ( .A1(n9129), .A2(n9528), .B1(n9128), .B2(n9531), .ZN(n9339)
         );
  OAI22_X1 U10591 ( .A1(n9131), .A2(n9343), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9130), .ZN(n9132) );
  AOI21_X1 U10592 ( .B1(n9339), .B2(n9133), .A(n9132), .ZN(n9134) );
  INV_X1 U10593 ( .A(n9135), .ZN(n9139) );
  OAI22_X1 U10594 ( .A1(n9139), .A2(n9138), .B1(n9137), .B2(n9136), .ZN(n9141)
         );
  NAND2_X1 U10595 ( .A1(n9141), .A2(n9140), .ZN(n9152) );
  NAND2_X1 U10596 ( .A1(n9143), .A2(n9142), .ZN(n9144) );
  OAI21_X1 U10597 ( .B1(n9146), .B2(n9145), .A(n9144), .ZN(n9150) );
  OAI22_X1 U10598 ( .A1(n9148), .A2(n9499), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9147), .ZN(n9149) );
  NOR2_X1 U10599 ( .A1(n9150), .A2(n9149), .ZN(n9151) );
  OAI211_X1 U10600 ( .C1(n9154), .C2(n9153), .A(n9152), .B(n9151), .ZN(
        P2_U3243) );
  MUX2_X1 U10601 ( .A(n9155), .B(P2_DATAO_REG_30__SCAN_IN), .S(n9178), .Z(
        P2_U3582) );
  MUX2_X1 U10602 ( .A(n9156), .B(P2_DATAO_REG_29__SCAN_IN), .S(n9178), .Z(
        P2_U3581) );
  MUX2_X1 U10603 ( .A(n9157), .B(P2_DATAO_REG_28__SCAN_IN), .S(n9178), .Z(
        P2_U3580) );
  MUX2_X1 U10604 ( .A(n9158), .B(P2_DATAO_REG_27__SCAN_IN), .S(n9178), .Z(
        P2_U3579) );
  MUX2_X1 U10605 ( .A(n9159), .B(P2_DATAO_REG_26__SCAN_IN), .S(n9178), .Z(
        P2_U3578) );
  MUX2_X1 U10606 ( .A(n9160), .B(P2_DATAO_REG_24__SCAN_IN), .S(n9178), .Z(
        P2_U3576) );
  MUX2_X1 U10607 ( .A(n9161), .B(P2_DATAO_REG_23__SCAN_IN), .S(n9178), .Z(
        P2_U3575) );
  MUX2_X1 U10608 ( .A(n9162), .B(P2_DATAO_REG_22__SCAN_IN), .S(n9178), .Z(
        P2_U3574) );
  MUX2_X1 U10609 ( .A(n9163), .B(P2_DATAO_REG_21__SCAN_IN), .S(n9178), .Z(
        P2_U3573) );
  MUX2_X1 U10610 ( .A(n9465), .B(P2_DATAO_REG_20__SCAN_IN), .S(n9178), .Z(
        P2_U3572) );
  MUX2_X1 U10611 ( .A(n9164), .B(P2_DATAO_REG_19__SCAN_IN), .S(n9178), .Z(
        P2_U3571) );
  MUX2_X1 U10612 ( .A(n9463), .B(P2_DATAO_REG_18__SCAN_IN), .S(n9178), .Z(
        P2_U3570) );
  MUX2_X1 U10613 ( .A(n9165), .B(P2_DATAO_REG_16__SCAN_IN), .S(n9178), .Z(
        P2_U3568) );
  MUX2_X1 U10614 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9166), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10615 ( .A(n9167), .B(P2_DATAO_REG_14__SCAN_IN), .S(n9178), .Z(
        P2_U3566) );
  MUX2_X1 U10616 ( .A(n9168), .B(P2_DATAO_REG_13__SCAN_IN), .S(n9178), .Z(
        P2_U3565) );
  MUX2_X1 U10617 ( .A(n9169), .B(P2_DATAO_REG_12__SCAN_IN), .S(n9178), .Z(
        P2_U3564) );
  MUX2_X1 U10618 ( .A(n9170), .B(P2_DATAO_REG_11__SCAN_IN), .S(n9178), .Z(
        P2_U3563) );
  MUX2_X1 U10619 ( .A(n9171), .B(P2_DATAO_REG_10__SCAN_IN), .S(n9178), .Z(
        P2_U3562) );
  MUX2_X1 U10620 ( .A(n9172), .B(P2_DATAO_REG_9__SCAN_IN), .S(n9178), .Z(
        P2_U3561) );
  MUX2_X1 U10621 ( .A(n9173), .B(P2_DATAO_REG_8__SCAN_IN), .S(n9178), .Z(
        P2_U3560) );
  MUX2_X1 U10622 ( .A(n9174), .B(P2_DATAO_REG_7__SCAN_IN), .S(n9178), .Z(
        P2_U3559) );
  MUX2_X1 U10623 ( .A(n9175), .B(P2_DATAO_REG_6__SCAN_IN), .S(n9178), .Z(
        P2_U3558) );
  MUX2_X1 U10624 ( .A(n9176), .B(P2_DATAO_REG_4__SCAN_IN), .S(n9178), .Z(
        P2_U3556) );
  MUX2_X1 U10625 ( .A(n9177), .B(P2_DATAO_REG_3__SCAN_IN), .S(n9178), .Z(
        P2_U3555) );
  MUX2_X1 U10626 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n6051), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U10627 ( .A(n6045), .B(P2_DATAO_REG_1__SCAN_IN), .S(n9178), .Z(
        P2_U3553) );
  NAND2_X1 U10628 ( .A1(n9263), .A2(n9179), .ZN(n9193) );
  NOR2_X1 U10629 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9180), .ZN(n9181) );
  AOI21_X1 U10630 ( .B1(n9289), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n9181), .ZN(
        n9192) );
  OR3_X1 U10631 ( .A1(n9184), .A2(n9183), .A3(n9182), .ZN(n9185) );
  NAND3_X1 U10632 ( .A1(n9291), .A2(n9186), .A3(n9185), .ZN(n9191) );
  OAI211_X1 U10633 ( .C1(n9189), .C2(n9188), .A(n9258), .B(n9187), .ZN(n9190)
         );
  NAND4_X1 U10634 ( .A1(n9193), .A2(n9192), .A3(n9191), .A4(n9190), .ZN(
        P2_U3248) );
  NAND2_X1 U10635 ( .A1(n9263), .A2(n9194), .ZN(n9209) );
  NOR2_X1 U10636 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5173), .ZN(n9195) );
  AOI21_X1 U10637 ( .B1(n9289), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n9195), .ZN(
        n9208) );
  INV_X1 U10638 ( .A(n9196), .ZN(n9199) );
  MUX2_X1 U10639 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n6757), .S(n9197), .Z(n9198)
         );
  NAND3_X1 U10640 ( .A1(n9200), .A2(n9199), .A3(n9198), .ZN(n9201) );
  NAND3_X1 U10641 ( .A1(n9291), .A2(n9202), .A3(n9201), .ZN(n9207) );
  OAI211_X1 U10642 ( .C1(n9205), .C2(n9204), .A(n9258), .B(n9203), .ZN(n9206)
         );
  NAND4_X1 U10643 ( .A1(n9209), .A2(n9208), .A3(n9207), .A4(n9206), .ZN(
        P2_U3250) );
  NAND2_X1 U10644 ( .A1(n9263), .A2(n9210), .ZN(n9222) );
  NOR2_X1 U10645 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5200), .ZN(n9211) );
  AOI21_X1 U10646 ( .B1(n9289), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n9211), .ZN(
        n9221) );
  OR3_X1 U10647 ( .A1(n9214), .A2(n9213), .A3(n9212), .ZN(n9215) );
  NAND3_X1 U10648 ( .A1(n9291), .A2(n9228), .A3(n9215), .ZN(n9220) );
  OAI211_X1 U10649 ( .C1(n9218), .C2(n9217), .A(n9258), .B(n9216), .ZN(n9219)
         );
  NAND4_X1 U10650 ( .A1(n9222), .A2(n9221), .A3(n9220), .A4(n9219), .ZN(
        P2_U3252) );
  NAND2_X1 U10651 ( .A1(n9263), .A2(n9223), .ZN(n9237) );
  INV_X1 U10652 ( .A(n9224), .ZN(n9225) );
  AOI21_X1 U10653 ( .B1(n9289), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n9225), .ZN(
        n9236) );
  INV_X1 U10654 ( .A(n9240), .ZN(n9230) );
  NAND3_X1 U10655 ( .A1(n9228), .A2(n9227), .A3(n9226), .ZN(n9229) );
  NAND3_X1 U10656 ( .A1(n9291), .A2(n9230), .A3(n9229), .ZN(n9235) );
  OAI211_X1 U10657 ( .C1(n9233), .C2(n9232), .A(n9258), .B(n9231), .ZN(n9234)
         );
  NAND4_X1 U10658 ( .A1(n9237), .A2(n9236), .A3(n9235), .A4(n9234), .ZN(
        P2_U3253) );
  OR3_X1 U10659 ( .A1(n9240), .A2(n9239), .A3(n9238), .ZN(n9241) );
  NAND3_X1 U10660 ( .A1(n9242), .A2(n9291), .A3(n9241), .ZN(n9251) );
  AOI21_X1 U10661 ( .B1(n9289), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n9243), .ZN(
        n9250) );
  OAI211_X1 U10662 ( .C1(n9246), .C2(n9245), .A(n9258), .B(n9244), .ZN(n9249)
         );
  NAND2_X1 U10663 ( .A1(n9263), .A2(n9247), .ZN(n9248) );
  NAND4_X1 U10664 ( .A1(n9251), .A2(n9250), .A3(n9249), .A4(n9248), .ZN(
        P2_U3254) );
  OAI21_X1 U10665 ( .B1(n9254), .B2(n9253), .A(n9252), .ZN(n9255) );
  NAND2_X1 U10666 ( .A1(n9255), .A2(n9291), .ZN(n9267) );
  NOR2_X1 U10667 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9256), .ZN(n9257) );
  AOI21_X1 U10668 ( .B1(n9289), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n9257), .ZN(
        n9266) );
  OAI211_X1 U10669 ( .C1(n9261), .C2(n9260), .A(n9259), .B(n9258), .ZN(n9265)
         );
  NAND2_X1 U10670 ( .A1(n9263), .A2(n9262), .ZN(n9264) );
  NAND4_X1 U10671 ( .A1(n9267), .A2(n9266), .A3(n9265), .A4(n9264), .ZN(
        P2_U3256) );
  OAI211_X1 U10672 ( .C1(n9270), .C2(n9269), .A(n9268), .B(n9291), .ZN(n9274)
         );
  NOR2_X1 U10673 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9271), .ZN(n9272) );
  AOI21_X1 U10674 ( .B1(n9289), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n9272), .ZN(
        n9273) );
  OAI211_X1 U10675 ( .C1(n9286), .C2(n9275), .A(n9274), .B(n9273), .ZN(n9281)
         );
  INV_X1 U10676 ( .A(n9276), .ZN(n9277) );
  AOI211_X1 U10677 ( .C1(n9279), .C2(n9278), .A(n9295), .B(n9277), .ZN(n9280)
         );
  OR2_X1 U10678 ( .A1(n9281), .A2(n9280), .ZN(P2_U3262) );
  INV_X1 U10679 ( .A(n9282), .ZN(n9283) );
  AOI21_X1 U10680 ( .B1(n9285), .B2(n9284), .A(n9283), .ZN(n9296) );
  NOR2_X1 U10681 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4653), .ZN(n9288) );
  NOR2_X1 U10682 ( .A1(n9286), .A2(n4751), .ZN(n9287) );
  AOI211_X1 U10683 ( .C1(n9289), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n9288), .B(
        n9287), .ZN(n9294) );
  OAI211_X1 U10684 ( .C1(P2_REG2_REG_18__SCAN_IN), .C2(n9292), .A(n9291), .B(
        n9290), .ZN(n9293) );
  OAI211_X1 U10685 ( .C1(n9296), .C2(n9295), .A(n9294), .B(n9293), .ZN(
        P2_U3263) );
  NOR2_X1 U10686 ( .A1(n4374), .A2(n9544), .ZN(n9303) );
  NOR2_X1 U10687 ( .A1(n5978), .A2(n9437), .ZN(n9297) );
  AOI211_X1 U10688 ( .C1(n4374), .C2(P2_REG2_REG_31__SCAN_IN), .A(n9303), .B(
        n9297), .ZN(n9298) );
  OAI21_X1 U10689 ( .B1(n9299), .B2(n9491), .A(n9298), .ZN(P2_U3265) );
  OAI211_X1 U10690 ( .C1(n9301), .C2(n9638), .A(n9484), .B(n9300), .ZN(n9545)
         );
  NOR2_X1 U10691 ( .A1(n9638), .A2(n9437), .ZN(n9302) );
  AOI211_X1 U10692 ( .C1(n4374), .C2(P2_REG2_REG_30__SCAN_IN), .A(n9303), .B(
        n9302), .ZN(n9304) );
  OAI21_X1 U10693 ( .B1(n9491), .B2(n9545), .A(n9304), .ZN(P2_U3266) );
  INV_X1 U10694 ( .A(n9305), .ZN(n9314) );
  OAI21_X1 U10695 ( .B1(n9307), .B2(n9485), .A(n9306), .ZN(n9312) );
  AOI22_X1 U10696 ( .A1(n9308), .A2(n9521), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n4374), .ZN(n9309) );
  OAI21_X1 U10697 ( .B1(n9310), .B2(n9491), .A(n9309), .ZN(n9311) );
  AOI21_X1 U10698 ( .B1(n9312), .B2(n9536), .A(n9311), .ZN(n9313) );
  OAI21_X1 U10699 ( .B1(n9314), .B2(n9495), .A(n9313), .ZN(P2_U3267) );
  XNOR2_X1 U10700 ( .A(n9316), .B(n9315), .ZN(n9556) );
  INV_X1 U10701 ( .A(n9556), .ZN(n9332) );
  NAND2_X1 U10702 ( .A1(n9317), .A2(n9524), .ZN(n9323) );
  AOI21_X1 U10703 ( .B1(n9318), .B2(n9320), .A(n9319), .ZN(n9322) );
  OAI21_X1 U10704 ( .B1(n9323), .B2(n9322), .A(n9321), .ZN(n9554) );
  INV_X1 U10705 ( .A(n9324), .ZN(n9325) );
  AOI211_X1 U10706 ( .C1(n9326), .C2(n9341), .A(n9538), .B(n9325), .ZN(n9555)
         );
  NAND2_X1 U10707 ( .A1(n9555), .A2(n9540), .ZN(n9329) );
  AOI22_X1 U10708 ( .A1(n9327), .A2(n9535), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n4374), .ZN(n9328) );
  OAI211_X1 U10709 ( .C1(n9642), .C2(n9437), .A(n9329), .B(n9328), .ZN(n9330)
         );
  AOI21_X1 U10710 ( .B1(n9554), .B2(n9536), .A(n9330), .ZN(n9331) );
  OAI21_X1 U10711 ( .B1(n9332), .B2(n9495), .A(n9331), .ZN(P2_U3269) );
  XNOR2_X1 U10712 ( .A(n9333), .B(n9336), .ZN(n9560) );
  OAI21_X1 U10713 ( .B1(n4566), .B2(n9337), .A(n9336), .ZN(n9338) );
  NAND2_X1 U10714 ( .A1(n9338), .A2(n9318), .ZN(n9340) );
  INV_X1 U10715 ( .A(n9559), .ZN(n9348) );
  OAI211_X1 U10716 ( .C1(n9355), .C2(n9646), .A(n9484), .B(n9341), .ZN(n9558)
         );
  INV_X1 U10717 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9342) );
  OAI22_X1 U10718 ( .A1(n9343), .A2(n9485), .B1(n9342), .B2(n9536), .ZN(n9344)
         );
  AOI21_X1 U10719 ( .B1(n9345), .B2(n9521), .A(n9344), .ZN(n9346) );
  OAI21_X1 U10720 ( .B1(n9558), .B2(n9515), .A(n9346), .ZN(n9347) );
  AOI21_X1 U10721 ( .B1(n9348), .B2(n9536), .A(n9347), .ZN(n9349) );
  OAI21_X1 U10722 ( .B1(n9560), .B2(n9495), .A(n9349), .ZN(P2_U3270) );
  XNOR2_X1 U10723 ( .A(n9350), .B(n9353), .ZN(n9568) );
  AOI22_X1 U10724 ( .A1(n9566), .A2(n9521), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n4374), .ZN(n9363) );
  OR2_X1 U10725 ( .A1(n9351), .A2(n9373), .ZN(n9365) );
  INV_X1 U10726 ( .A(n9367), .ZN(n9356) );
  AOI211_X1 U10727 ( .C1(n9566), .C2(n9356), .A(n9538), .B(n9355), .ZN(n9565)
         );
  INV_X1 U10728 ( .A(n9565), .ZN(n9360) );
  INV_X1 U10729 ( .A(n9357), .ZN(n9358) );
  OAI22_X1 U10730 ( .A1(n9360), .A2(n9359), .B1(n9485), .B2(n9358), .ZN(n9361)
         );
  OAI21_X1 U10731 ( .B1(n9564), .B2(n9361), .A(n9536), .ZN(n9362) );
  OAI211_X1 U10732 ( .C1(n9568), .C2(n9495), .A(n9363), .B(n9362), .ZN(
        P2_U3271) );
  AOI21_X1 U10733 ( .B1(n9351), .B2(n9373), .A(n9442), .ZN(n9366) );
  AOI21_X1 U10734 ( .B1(n9366), .B2(n9365), .A(n9364), .ZN(n9572) );
  AOI211_X1 U10735 ( .C1(n9570), .C2(n9381), .A(n9538), .B(n9367), .ZN(n9569)
         );
  INV_X1 U10736 ( .A(n9570), .ZN(n9371) );
  INV_X1 U10737 ( .A(n9368), .ZN(n9369) );
  AOI22_X1 U10738 ( .A1(n4374), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n9369), .B2(
        n9535), .ZN(n9370) );
  OAI21_X1 U10739 ( .B1(n9371), .B2(n9437), .A(n9370), .ZN(n9377) );
  OAI21_X1 U10740 ( .B1(n9374), .B2(n9373), .A(n9372), .ZN(n9375) );
  INV_X1 U10741 ( .A(n9375), .ZN(n9573) );
  NOR2_X1 U10742 ( .A1(n9573), .A2(n9495), .ZN(n9376) );
  AOI211_X1 U10743 ( .C1(n9569), .C2(n9540), .A(n9377), .B(n9376), .ZN(n9378)
         );
  OAI21_X1 U10744 ( .B1(n4374), .B2(n9572), .A(n9378), .ZN(P2_U3272) );
  AOI21_X1 U10745 ( .B1(n9390), .B2(n9380), .A(n9379), .ZN(n9576) );
  INV_X1 U10746 ( .A(n9576), .ZN(n9397) );
  INV_X1 U10747 ( .A(n9381), .ZN(n9382) );
  AOI211_X1 U10748 ( .C1(n9383), .C2(n9400), .A(n9538), .B(n9382), .ZN(n9575)
         );
  INV_X1 U10749 ( .A(n9383), .ZN(n9652) );
  INV_X1 U10750 ( .A(n9384), .ZN(n9385) );
  AOI22_X1 U10751 ( .A1(n4374), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n9385), .B2(
        n9535), .ZN(n9386) );
  OAI21_X1 U10752 ( .B1(n9652), .B2(n9437), .A(n9386), .ZN(n9387) );
  AOI21_X1 U10753 ( .B1(n9575), .B2(n9540), .A(n9387), .ZN(n9396) );
  NAND2_X1 U10754 ( .A1(n9388), .A2(n9389), .ZN(n9391) );
  XNOR2_X1 U10755 ( .A(n9391), .B(n9390), .ZN(n9394) );
  INV_X1 U10756 ( .A(n9392), .ZN(n9393) );
  OAI21_X1 U10757 ( .B1(n9394), .B2(n9442), .A(n9393), .ZN(n9574) );
  NAND2_X1 U10758 ( .A1(n9574), .A2(n9536), .ZN(n9395) );
  OAI211_X1 U10759 ( .C1(n9397), .C2(n9495), .A(n9396), .B(n9395), .ZN(
        P2_U3273) );
  XNOR2_X1 U10760 ( .A(n9398), .B(n9404), .ZN(n9583) );
  OR2_X1 U10761 ( .A1(n9412), .A2(n4988), .ZN(n9399) );
  AND3_X1 U10762 ( .A1(n9400), .A2(n9399), .A3(n9484), .ZN(n9579) );
  NAND2_X1 U10763 ( .A1(n9580), .A2(n9521), .ZN(n9402) );
  NAND2_X1 U10764 ( .A1(n4374), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n9401) );
  OAI211_X1 U10765 ( .C1(n9485), .C2(n9403), .A(n9402), .B(n9401), .ZN(n9409)
         );
  AOI21_X1 U10766 ( .B1(n9405), .B2(n9404), .A(n9442), .ZN(n9407) );
  AOI21_X1 U10767 ( .B1(n9407), .B2(n9388), .A(n9406), .ZN(n9582) );
  NOR2_X1 U10768 ( .A1(n9582), .A2(n4374), .ZN(n9408) );
  AOI211_X1 U10769 ( .C1(n9579), .C2(n9540), .A(n9409), .B(n9408), .ZN(n9410)
         );
  OAI21_X1 U10770 ( .B1(n9583), .B2(n9495), .A(n9410), .ZN(P2_U3274) );
  XOR2_X1 U10771 ( .A(n9411), .B(n9424), .Z(n9586) );
  INV_X1 U10772 ( .A(n9586), .ZN(n9430) );
  INV_X1 U10773 ( .A(n9432), .ZN(n9413) );
  AOI211_X1 U10774 ( .C1(n9414), .C2(n9413), .A(n9538), .B(n9412), .ZN(n9585)
         );
  INV_X1 U10775 ( .A(n9415), .ZN(n9416) );
  AOI22_X1 U10776 ( .A1(n4374), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9416), .B2(
        n9535), .ZN(n9417) );
  OAI21_X1 U10777 ( .B1(n9657), .B2(n9437), .A(n9417), .ZN(n9418) );
  AOI21_X1 U10778 ( .B1(n9585), .B2(n9540), .A(n9418), .ZN(n9429) );
  NAND2_X1 U10779 ( .A1(n9460), .A2(n9461), .ZN(n9459) );
  NAND2_X1 U10780 ( .A1(n9459), .A2(n9419), .ZN(n9440) );
  NAND2_X1 U10781 ( .A1(n9440), .A2(n9420), .ZN(n9422) );
  NAND2_X1 U10782 ( .A1(n9422), .A2(n9421), .ZN(n9423) );
  XOR2_X1 U10783 ( .A(n9424), .B(n9423), .Z(n9427) );
  INV_X1 U10784 ( .A(n9425), .ZN(n9426) );
  OAI21_X1 U10785 ( .B1(n9427), .B2(n9442), .A(n9426), .ZN(n9584) );
  NAND2_X1 U10786 ( .A1(n9584), .A2(n9536), .ZN(n9428) );
  OAI211_X1 U10787 ( .C1(n9430), .C2(n9495), .A(n9429), .B(n9428), .ZN(
        P2_U3275) );
  XOR2_X1 U10788 ( .A(n9439), .B(n9431), .Z(n9591) );
  INV_X1 U10789 ( .A(n9591), .ZN(n9446) );
  AOI211_X1 U10790 ( .C1(n9433), .C2(n9454), .A(n9538), .B(n9432), .ZN(n9590)
         );
  INV_X1 U10791 ( .A(n9434), .ZN(n9435) );
  AOI22_X1 U10792 ( .A1(n4374), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9435), .B2(
        n9535), .ZN(n9436) );
  OAI21_X1 U10793 ( .B1(n4951), .B2(n9437), .A(n9436), .ZN(n9438) );
  AOI21_X1 U10794 ( .B1(n9590), .B2(n9540), .A(n9438), .ZN(n9445) );
  XNOR2_X1 U10795 ( .A(n9440), .B(n9439), .ZN(n9443) );
  OAI21_X1 U10796 ( .B1(n9443), .B2(n9442), .A(n9441), .ZN(n9589) );
  NAND2_X1 U10797 ( .A1(n9589), .A2(n9536), .ZN(n9444) );
  OAI211_X1 U10798 ( .C1(n9446), .C2(n9495), .A(n9445), .B(n9444), .ZN(
        P2_U3276) );
  NAND2_X1 U10799 ( .A1(n9448), .A2(n9449), .ZN(n9472) );
  NAND2_X1 U10800 ( .A1(n9472), .A2(n9450), .ZN(n9452) );
  NAND2_X1 U10801 ( .A1(n9452), .A2(n9451), .ZN(n9453) );
  XNOR2_X1 U10802 ( .A(n9453), .B(n9461), .ZN(n9598) );
  AOI21_X1 U10803 ( .B1(n9483), .B2(n9595), .A(n9538), .ZN(n9455) );
  AND2_X1 U10804 ( .A1(n9455), .A2(n9454), .ZN(n9594) );
  NAND2_X1 U10805 ( .A1(n9595), .A2(n9521), .ZN(n9457) );
  NAND2_X1 U10806 ( .A1(n4374), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n9456) );
  OAI211_X1 U10807 ( .C1(n9485), .C2(n9458), .A(n9457), .B(n9456), .ZN(n9468)
         );
  OAI21_X1 U10808 ( .B1(n9461), .B2(n9460), .A(n9459), .ZN(n9466) );
  AOI222_X1 U10809 ( .A1(n9524), .A2(n9466), .B1(n9465), .B2(n9464), .C1(n9463), .C2(n9462), .ZN(n9597) );
  NOR2_X1 U10810 ( .A1(n9597), .A2(n4374), .ZN(n9467) );
  AOI211_X1 U10811 ( .C1(n9594), .C2(n9469), .A(n9468), .B(n9467), .ZN(n9470)
         );
  OAI21_X1 U10812 ( .B1(n9598), .B2(n9495), .A(n9470), .ZN(P2_U3277) );
  XNOR2_X1 U10813 ( .A(n9472), .B(n9471), .ZN(n9601) );
  NAND2_X1 U10814 ( .A1(n9474), .A2(n9473), .ZN(n9476) );
  NAND2_X1 U10815 ( .A1(n9476), .A2(n9475), .ZN(n9477) );
  NAND2_X1 U10816 ( .A1(n9478), .A2(n9477), .ZN(n9482) );
  OAI22_X1 U10817 ( .A1(n9480), .A2(n9528), .B1(n9479), .B2(n9531), .ZN(n9481)
         );
  AOI21_X1 U10818 ( .B1(n9482), .B2(n9524), .A(n9481), .ZN(n9600) );
  INV_X1 U10819 ( .A(n9600), .ZN(n9493) );
  OAI211_X1 U10820 ( .C1(n9507), .C2(n9665), .A(n9484), .B(n9483), .ZN(n9599)
         );
  OAI22_X1 U10821 ( .A1(n9536), .A2(n9487), .B1(n9486), .B2(n9485), .ZN(n9488)
         );
  AOI21_X1 U10822 ( .B1(n9489), .B2(n9521), .A(n9488), .ZN(n9490) );
  OAI21_X1 U10823 ( .B1(n9599), .B2(n9491), .A(n9490), .ZN(n9492) );
  AOI21_X1 U10824 ( .B1(n9493), .B2(n9536), .A(n9492), .ZN(n9494) );
  OAI21_X1 U10825 ( .B1(n9601), .B2(n9495), .A(n9494), .ZN(P2_U3278) );
  XNOR2_X1 U10826 ( .A(n9497), .B(n9496), .ZN(n9498) );
  NAND2_X1 U10827 ( .A1(n9498), .A2(n9524), .ZN(n9503) );
  OAI22_X1 U10828 ( .A1(n9500), .A2(n9528), .B1(n9499), .B2(n9531), .ZN(n9501)
         );
  INV_X1 U10829 ( .A(n9501), .ZN(n9502) );
  NAND2_X1 U10830 ( .A1(n9503), .A2(n9502), .ZN(n9608) );
  INV_X1 U10831 ( .A(n9608), .ZN(n9518) );
  NAND2_X1 U10832 ( .A1(n9505), .A2(n9504), .ZN(n9506) );
  NAND2_X1 U10833 ( .A1(n9448), .A2(n9506), .ZN(n9604) );
  INV_X1 U10834 ( .A(n9507), .ZN(n9510) );
  AOI21_X1 U10835 ( .B1(n9508), .B2(n9512), .A(n9538), .ZN(n9509) );
  NAND2_X1 U10836 ( .A1(n9510), .A2(n9509), .ZN(n9605) );
  AOI22_X1 U10837 ( .A1(n4374), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n9511), .B2(
        n9535), .ZN(n9514) );
  NAND2_X1 U10838 ( .A1(n9512), .A2(n9521), .ZN(n9513) );
  OAI211_X1 U10839 ( .C1(n9605), .C2(n9515), .A(n9514), .B(n9513), .ZN(n9516)
         );
  AOI21_X1 U10840 ( .B1(n9604), .B2(n9522), .A(n9516), .ZN(n9517) );
  OAI21_X1 U10841 ( .B1(n9518), .B2(n4374), .A(n9517), .ZN(P2_U3279) );
  OAI21_X1 U10842 ( .B1(n5883), .B2(n9520), .A(n9519), .ZN(n10491) );
  INV_X1 U10843 ( .A(n10488), .ZN(n9539) );
  AOI22_X1 U10844 ( .A1(n9522), .A2(n10491), .B1(n9521), .B2(n9539), .ZN(n9543) );
  NAND2_X1 U10845 ( .A1(n5883), .A2(n9523), .ZN(n9525) );
  NAND2_X1 U10846 ( .A1(n9525), .A2(n9524), .ZN(n9526) );
  OR2_X1 U10847 ( .A1(n9527), .A2(n9526), .ZN(n9534) );
  OAI22_X1 U10848 ( .A1(n9531), .A2(n9530), .B1(n9529), .B2(n9528), .ZN(n9532)
         );
  INV_X1 U10849 ( .A(n9532), .ZN(n9533) );
  NAND2_X1 U10850 ( .A1(n9534), .A2(n9533), .ZN(n10490) );
  AOI22_X1 U10851 ( .A1(n9536), .A2(n10490), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9535), .ZN(n9542) );
  AOI211_X1 U10852 ( .C1(n10481), .C2(n9539), .A(n9538), .B(n9537), .ZN(n10486) );
  AOI22_X1 U10853 ( .A1(n9540), .A2(n10486), .B1(n4374), .B2(
        P2_REG2_REG_1__SCAN_IN), .ZN(n9541) );
  NAND3_X1 U10854 ( .A1(n9543), .A2(n9542), .A3(n9541), .ZN(P2_U3295) );
  AND2_X1 U10855 ( .A1(n9545), .A2(n9544), .ZN(n9635) );
  MUX2_X1 U10856 ( .A(n9546), .B(n9635), .S(n10522), .Z(n9547) );
  OAI21_X1 U10857 ( .B1(n9638), .B2(n9615), .A(n9547), .ZN(P2_U3550) );
  INV_X1 U10858 ( .A(n9549), .ZN(n9551) );
  OAI21_X1 U10859 ( .B1(n9553), .B2(n9627), .A(n9552), .ZN(n9639) );
  MUX2_X1 U10860 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9639), .S(n10522), .Z(
        P2_U3548) );
  INV_X1 U10861 ( .A(n9561), .ZN(n9643) );
  MUX2_X1 U10862 ( .A(n9562), .B(n9643), .S(n10522), .Z(n9563) );
  OAI21_X1 U10863 ( .B1(n9568), .B2(n9627), .A(n9567), .ZN(n9647) );
  MUX2_X1 U10864 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9647), .S(n10522), .Z(
        P2_U3545) );
  AOI21_X1 U10865 ( .B1(n9630), .B2(n9570), .A(n9569), .ZN(n9571) );
  OAI211_X1 U10866 ( .C1(n9573), .C2(n9627), .A(n9572), .B(n9571), .ZN(n9648)
         );
  MUX2_X1 U10867 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9648), .S(n10522), .Z(
        P2_U3544) );
  INV_X1 U10868 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9577) );
  AOI211_X1 U10869 ( .C1(n9576), .C2(n10510), .A(n9575), .B(n9574), .ZN(n9649)
         );
  MUX2_X1 U10870 ( .A(n9577), .B(n9649), .S(n10522), .Z(n9578) );
  OAI21_X1 U10871 ( .B1(n9652), .B2(n9615), .A(n9578), .ZN(P2_U3543) );
  AOI21_X1 U10872 ( .B1(n9630), .B2(n9580), .A(n9579), .ZN(n9581) );
  OAI211_X1 U10873 ( .C1(n9583), .C2(n9627), .A(n9582), .B(n9581), .ZN(n9653)
         );
  MUX2_X1 U10874 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9653), .S(n10522), .Z(
        P2_U3542) );
  AOI211_X1 U10875 ( .C1(n10510), .C2(n9586), .A(n9585), .B(n9584), .ZN(n9654)
         );
  MUX2_X1 U10876 ( .A(n9587), .B(n9654), .S(n10522), .Z(n9588) );
  OAI21_X1 U10877 ( .B1(n9657), .B2(n9615), .A(n9588), .ZN(P2_U3541) );
  INV_X1 U10878 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9592) );
  AOI211_X1 U10879 ( .C1(n9591), .C2(n10510), .A(n9590), .B(n9589), .ZN(n9658)
         );
  MUX2_X1 U10880 ( .A(n9592), .B(n9658), .S(n10522), .Z(n9593) );
  OAI21_X1 U10881 ( .B1(n4951), .B2(n9615), .A(n9593), .ZN(P2_U3540) );
  AOI21_X1 U10882 ( .B1(n9630), .B2(n9595), .A(n9594), .ZN(n9596) );
  OAI211_X1 U10883 ( .C1(n9627), .C2(n9598), .A(n9597), .B(n9596), .ZN(n9661)
         );
  MUX2_X1 U10884 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9661), .S(n10522), .Z(
        P2_U3539) );
  OAI211_X1 U10885 ( .C1(n9627), .C2(n9601), .A(n9600), .B(n9599), .ZN(n9662)
         );
  MUX2_X1 U10886 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9662), .S(n10522), .Z(
        n9602) );
  INV_X1 U10887 ( .A(n9602), .ZN(n9603) );
  OAI21_X1 U10888 ( .B1(n9665), .B2(n9615), .A(n9603), .ZN(P2_U3538) );
  NAND2_X1 U10889 ( .A1(n9604), .A2(n10510), .ZN(n9606) );
  OAI211_X1 U10890 ( .C1(n9607), .C2(n10507), .A(n9606), .B(n9605), .ZN(n9609)
         );
  MUX2_X1 U10891 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9666), .S(n10522), .Z(
        P2_U3537) );
  INV_X1 U10892 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9613) );
  AOI211_X1 U10893 ( .C1(n9612), .C2(n10510), .A(n9611), .B(n9610), .ZN(n9667)
         );
  MUX2_X1 U10894 ( .A(n9613), .B(n9667), .S(n10522), .Z(n9614) );
  OAI21_X1 U10895 ( .B1(n9671), .B2(n9615), .A(n9614), .ZN(P2_U3536) );
  INV_X1 U10896 ( .A(n9616), .ZN(n9621) );
  AOI21_X1 U10897 ( .B1(n9630), .B2(n9618), .A(n9617), .ZN(n9619) );
  OAI211_X1 U10898 ( .C1(n9627), .C2(n9621), .A(n9620), .B(n9619), .ZN(n9672)
         );
  MUX2_X1 U10899 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9672), .S(n10522), .Z(
        P2_U3535) );
  AOI21_X1 U10900 ( .B1(n9630), .B2(n9623), .A(n9622), .ZN(n9624) );
  OAI211_X1 U10901 ( .C1(n9627), .C2(n9626), .A(n9625), .B(n9624), .ZN(n9673)
         );
  MUX2_X1 U10902 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9673), .S(n10522), .Z(
        P2_U3531) );
  AOI21_X1 U10903 ( .B1(n9630), .B2(n9629), .A(n9628), .ZN(n9631) );
  OAI211_X1 U10904 ( .C1(n9634), .C2(n9633), .A(n9632), .B(n9631), .ZN(n9674)
         );
  MUX2_X1 U10905 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n9674), .S(n10522), .Z(
        P2_U3529) );
  INV_X1 U10906 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9636) );
  MUX2_X1 U10907 ( .A(n9636), .B(n9635), .S(n10513), .Z(n9637) );
  OAI21_X1 U10908 ( .B1(n9638), .B2(n9670), .A(n9637), .ZN(P2_U3518) );
  MUX2_X1 U10909 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9639), .S(n10513), .Z(
        P2_U3516) );
  INV_X1 U10910 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9641) );
  INV_X1 U10911 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9644) );
  MUX2_X1 U10912 ( .A(n9644), .B(n9643), .S(n10513), .Z(n9645) );
  MUX2_X1 U10913 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9647), .S(n10513), .Z(
        P2_U3513) );
  MUX2_X1 U10914 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9648), .S(n10513), .Z(
        P2_U3512) );
  INV_X1 U10915 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9650) );
  MUX2_X1 U10916 ( .A(n9650), .B(n9649), .S(n10513), .Z(n9651) );
  OAI21_X1 U10917 ( .B1(n9652), .B2(n9670), .A(n9651), .ZN(P2_U3511) );
  MUX2_X1 U10918 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9653), .S(n10513), .Z(
        P2_U3510) );
  INV_X1 U10919 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9655) );
  MUX2_X1 U10920 ( .A(n9655), .B(n9654), .S(n10513), .Z(n9656) );
  OAI21_X1 U10921 ( .B1(n9657), .B2(n9670), .A(n9656), .ZN(P2_U3509) );
  MUX2_X1 U10922 ( .A(n9659), .B(n9658), .S(n10513), .Z(n9660) );
  OAI21_X1 U10923 ( .B1(n4951), .B2(n9670), .A(n9660), .ZN(P2_U3508) );
  MUX2_X1 U10924 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9661), .S(n10513), .Z(
        P2_U3507) );
  MUX2_X1 U10925 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9662), .S(n10513), .Z(
        n9663) );
  INV_X1 U10926 ( .A(n9663), .ZN(n9664) );
  OAI21_X1 U10927 ( .B1(n9665), .B2(n9670), .A(n9664), .ZN(P2_U3505) );
  MUX2_X1 U10928 ( .A(n9666), .B(P2_REG0_REG_17__SCAN_IN), .S(n10512), .Z(
        P2_U3502) );
  INV_X1 U10929 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9668) );
  MUX2_X1 U10930 ( .A(n9668), .B(n9667), .S(n10513), .Z(n9669) );
  OAI21_X1 U10931 ( .B1(n9671), .B2(n9670), .A(n9669), .ZN(P2_U3499) );
  MUX2_X1 U10932 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9672), .S(n10513), .Z(
        P2_U3496) );
  MUX2_X1 U10933 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n9673), .S(n10513), .Z(
        P2_U3484) );
  MUX2_X1 U10934 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n9674), .S(n10513), .Z(
        P2_U3478) );
  INV_X1 U10935 ( .A(n9675), .ZN(n10342) );
  NOR4_X1 U10936 ( .A1(n9678), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9677), .A4(
        P2_U3152), .ZN(n9679) );
  AOI21_X1 U10937 ( .B1(n9680), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9679), .ZN(
        n9681) );
  OAI21_X1 U10938 ( .B1(n10342), .B2(n9684), .A(n9681), .ZN(P2_U3327) );
  INV_X1 U10939 ( .A(n9682), .ZN(n10346) );
  OAI222_X1 U10940 ( .A1(n9686), .A2(n9685), .B1(n9684), .B2(n10346), .C1(
        n9683), .C2(P2_U3152), .ZN(P2_U3329) );
  MUX2_X1 U10941 ( .A(n9687), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U10942 ( .A1(n9689), .A2(n9688), .ZN(n9690) );
  XOR2_X1 U10943 ( .A(n9691), .B(n9690), .Z(n9696) );
  NAND2_X1 U10944 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9863) );
  OAI21_X1 U10945 ( .B1(n9831), .B2(n10183), .A(n9863), .ZN(n9692) );
  AOI21_X1 U10946 ( .B1(n9835), .B2(n9845), .A(n9692), .ZN(n9693) );
  OAI21_X1 U10947 ( .B1(n9832), .B2(n10169), .A(n9693), .ZN(n9694) );
  AOI21_X1 U10948 ( .B1(n10283), .B2(n4582), .A(n9694), .ZN(n9695) );
  OAI21_X1 U10949 ( .B1(n9696), .B2(n9825), .A(n9695), .ZN(P1_U3213) );
  INV_X1 U10950 ( .A(n9791), .ZN(n9697) );
  INV_X1 U10951 ( .A(n9768), .ZN(n9704) );
  AND2_X2 U10952 ( .A1(n9700), .A2(n9699), .ZN(n9767) );
  OAI21_X1 U10953 ( .B1(n9702), .B2(n9767), .A(n9701), .ZN(n9703) );
  OAI211_X1 U10954 ( .C1(n9704), .C2(n9767), .A(n9815), .B(n9703), .ZN(n9709)
         );
  OAI22_X1 U10955 ( .A1(n10014), .A2(n9831), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9705), .ZN(n9707) );
  NOR2_X1 U10956 ( .A1(n10015), .A2(n9775), .ZN(n9706) );
  AOI211_X1 U10957 ( .C1(n10021), .C2(n9773), .A(n9707), .B(n9706), .ZN(n9708)
         );
  OAI211_X1 U10958 ( .C1(n10023), .C2(n9838), .A(n9709), .B(n9708), .ZN(
        P1_U3214) );
  INV_X1 U10959 ( .A(n9711), .ZN(n9757) );
  OAI21_X1 U10960 ( .B1(n9710), .B2(n9757), .A(n9712), .ZN(n9714) );
  NOR2_X1 U10961 ( .A1(n9714), .A2(n9713), .ZN(n9801) );
  NAND2_X1 U10962 ( .A1(n9714), .A2(n9713), .ZN(n9802) );
  OAI21_X1 U10963 ( .B1(n9801), .B2(n9715), .A(n9802), .ZN(n9719) );
  XNOR2_X1 U10964 ( .A(n9717), .B(n9716), .ZN(n9718) );
  XNOR2_X1 U10965 ( .A(n9719), .B(n9718), .ZN(n9724) );
  NAND2_X1 U10966 ( .A1(n10047), .A2(n9835), .ZN(n9720) );
  NAND2_X1 U10967 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9953) );
  OAI211_X1 U10968 ( .C1(n10079), .C2(n9831), .A(n9720), .B(n9953), .ZN(n9722)
         );
  NOR2_X1 U10969 ( .A1(n10087), .A2(n9838), .ZN(n9721) );
  AOI211_X1 U10970 ( .C1(n10084), .C2(n9773), .A(n9722), .B(n9721), .ZN(n9723)
         );
  OAI21_X1 U10971 ( .B1(n9724), .B2(n9825), .A(n9723), .ZN(P1_U3217) );
  NAND2_X1 U10972 ( .A1(n9782), .A2(n9725), .ZN(n9726) );
  AND2_X1 U10973 ( .A1(n9726), .A2(n9779), .ZN(n9731) );
  INV_X1 U10974 ( .A(n9727), .ZN(n9729) );
  NOR2_X1 U10975 ( .A1(n9729), .A2(n9728), .ZN(n9730) );
  XNOR2_X1 U10976 ( .A(n9731), .B(n9730), .ZN(n9736) );
  AOI22_X1 U10977 ( .A1(n10047), .A2(n9785), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9733) );
  NAND2_X1 U10978 ( .A1(n10052), .A2(n9773), .ZN(n9732) );
  OAI211_X1 U10979 ( .C1(n10014), .C2(n9775), .A(n9733), .B(n9732), .ZN(n9734)
         );
  AOI21_X1 U10980 ( .B1(n10243), .B2(n4582), .A(n9734), .ZN(n9735) );
  OAI21_X1 U10981 ( .B1(n9736), .B2(n9825), .A(n9735), .ZN(P1_U3221) );
  INV_X1 U10982 ( .A(n9737), .ZN(n9738) );
  NOR3_X2 U10983 ( .A1(n9768), .A2(n9767), .A3(n9766), .ZN(n9771) );
  NOR3_X1 U10984 ( .A1(n9771), .A2(n9740), .A3(n9739), .ZN(n9741) );
  OAI21_X1 U10985 ( .B1(n9741), .B2(n9813), .A(n9815), .ZN(n9746) );
  AOI22_X1 U10986 ( .A1(n9742), .A2(n9773), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9743) );
  OAI21_X1 U10987 ( .B1(n10015), .B2(n9831), .A(n9743), .ZN(n9744) );
  AOI21_X1 U10988 ( .B1(n9843), .B2(n9835), .A(n9744), .ZN(n9745) );
  OAI211_X1 U10989 ( .C1(n9747), .C2(n9838), .A(n9746), .B(n9745), .ZN(
        P1_U3223) );
  XOR2_X1 U10990 ( .A(n9749), .B(n9748), .Z(n9750) );
  XNOR2_X1 U10991 ( .A(n9751), .B(n9750), .ZN(n9756) );
  NAND2_X1 U10992 ( .A1(n10095), .A2(n9835), .ZN(n9752) );
  NAND2_X1 U10993 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9906) );
  OAI211_X1 U10994 ( .C1(n10185), .C2(n9831), .A(n9752), .B(n9906), .ZN(n9754)
         );
  NOR2_X1 U10995 ( .A1(n10137), .A2(n9838), .ZN(n9753) );
  AOI211_X1 U10996 ( .C1(n10134), .C2(n9773), .A(n9754), .B(n9753), .ZN(n9755)
         );
  OAI21_X1 U10997 ( .B1(n9756), .B2(n9825), .A(n9755), .ZN(P1_U3224) );
  NOR2_X1 U10998 ( .A1(n9758), .A2(n9757), .ZN(n9759) );
  XNOR2_X1 U10999 ( .A(n9710), .B(n9759), .ZN(n9765) );
  INV_X1 U11000 ( .A(n9760), .ZN(n10149) );
  AND2_X1 U11001 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9921) );
  AOI21_X1 U11002 ( .B1(n9785), .B2(n10149), .A(n9921), .ZN(n9762) );
  NAND2_X1 U11003 ( .A1(n9773), .A2(n10110), .ZN(n9761) );
  OAI211_X1 U11004 ( .C1(n10079), .C2(n9775), .A(n9762), .B(n9761), .ZN(n9763)
         );
  AOI21_X1 U11005 ( .B1(n10266), .B2(n4582), .A(n9763), .ZN(n9764) );
  OAI21_X1 U11006 ( .B1(n9765), .B2(n9825), .A(n9764), .ZN(P1_U3226) );
  OAI21_X1 U11007 ( .B1(n9768), .B2(n9767), .A(n9766), .ZN(n9769) );
  INV_X1 U11008 ( .A(n9769), .ZN(n9770) );
  OAI21_X1 U11009 ( .B1(n9771), .B2(n9770), .A(n9815), .ZN(n9778) );
  INV_X1 U11010 ( .A(n9772), .ZN(n10006) );
  AOI22_X1 U11011 ( .A1(n10006), .A2(n9773), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9774) );
  OAI21_X1 U11012 ( .B1(n9993), .B2(n9775), .A(n9774), .ZN(n9776) );
  AOI21_X1 U11013 ( .B1(n9785), .B2(n10039), .A(n9776), .ZN(n9777) );
  OAI211_X1 U11014 ( .C1(n10009), .C2(n9838), .A(n9778), .B(n9777), .ZN(
        P1_U3227) );
  NAND2_X1 U11015 ( .A1(n9780), .A2(n9779), .ZN(n9784) );
  NAND2_X1 U11016 ( .A1(n9782), .A2(n9781), .ZN(n9783) );
  XOR2_X1 U11017 ( .A(n9784), .B(n9783), .Z(n9790) );
  NAND2_X1 U11018 ( .A1(n4836), .A2(n9835), .ZN(n9787) );
  AOI22_X1 U11019 ( .A1(n10094), .A2(n9785), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9786) );
  OAI211_X1 U11020 ( .C1(n9832), .C2(n10067), .A(n9787), .B(n9786), .ZN(n9788)
         );
  AOI21_X1 U11021 ( .B1(n10249), .B2(n4582), .A(n9788), .ZN(n9789) );
  OAI21_X1 U11022 ( .B1(n9790), .B2(n9825), .A(n9789), .ZN(P1_U3231) );
  NAND2_X1 U11023 ( .A1(n9792), .A2(n9791), .ZN(n9794) );
  XNOR2_X1 U11024 ( .A(n9794), .B(n9793), .ZN(n9795) );
  NAND2_X1 U11025 ( .A1(n9795), .A2(n9815), .ZN(n9800) );
  NOR2_X1 U11026 ( .A1(n10033), .A2(n9832), .ZN(n9798) );
  OAI22_X1 U11027 ( .A1(n10064), .A2(n9831), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9796), .ZN(n9797) );
  AOI211_X1 U11028 ( .C1(n10039), .C2(n9835), .A(n9798), .B(n9797), .ZN(n9799)
         );
  OAI211_X1 U11029 ( .C1(n10036), .C2(n9838), .A(n9800), .B(n9799), .ZN(
        P1_U3233) );
  INV_X1 U11030 ( .A(n9801), .ZN(n9803) );
  NAND2_X1 U11031 ( .A1(n9803), .A2(n9802), .ZN(n9805) );
  XNOR2_X1 U11032 ( .A(n9805), .B(n9804), .ZN(n9810) );
  NAND2_X1 U11033 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9930) );
  OAI21_X1 U11034 ( .B1(n10131), .B2(n9831), .A(n9930), .ZN(n9806) );
  AOI21_X1 U11035 ( .B1(n10094), .B2(n9835), .A(n9806), .ZN(n9807) );
  OAI21_X1 U11036 ( .B1(n9832), .B2(n10100), .A(n9807), .ZN(n9808) );
  AOI21_X1 U11037 ( .B1(n10258), .B2(n4582), .A(n9808), .ZN(n9809) );
  OAI21_X1 U11038 ( .B1(n9810), .B2(n9825), .A(n9809), .ZN(P1_U3236) );
  OAI21_X1 U11039 ( .B1(n9813), .B2(n9812), .A(n9811), .ZN(n9814) );
  NAND3_X1 U11040 ( .A1(n9816), .A2(n9815), .A3(n9814), .ZN(n9821) );
  NOR2_X1 U11041 ( .A1(n9993), .A2(n9831), .ZN(n9819) );
  OAI22_X1 U11042 ( .A1(n9985), .A2(n9832), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9817), .ZN(n9818) );
  AOI211_X1 U11043 ( .C1(n9842), .C2(n9835), .A(n9819), .B(n9818), .ZN(n9820)
         );
  OAI211_X1 U11044 ( .C1(n9983), .C2(n9838), .A(n9821), .B(n9820), .ZN(
        P1_U3238) );
  INV_X1 U11045 ( .A(n9823), .ZN(n9829) );
  AOI21_X1 U11046 ( .B1(n9824), .B2(n9823), .A(n9822), .ZN(n9826) );
  NOR2_X1 U11047 ( .A1(n9826), .A2(n9825), .ZN(n9827) );
  OAI21_X1 U11048 ( .B1(n9829), .B2(n9828), .A(n9827), .ZN(n9837) );
  NAND2_X1 U11049 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9883) );
  OAI21_X1 U11050 ( .B1(n9831), .B2(n9830), .A(n9883), .ZN(n9834) );
  NOR2_X1 U11051 ( .A1(n9832), .A2(n10157), .ZN(n9833) );
  AOI211_X1 U11052 ( .C1(n9835), .C2(n10149), .A(n9834), .B(n9833), .ZN(n9836)
         );
  OAI211_X1 U11053 ( .C1(n10161), .C2(n9838), .A(n9837), .B(n9836), .ZN(
        P1_U3239) );
  MUX2_X1 U11054 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9839), .S(n9858), .Z(
        P1_U3586) );
  MUX2_X1 U11055 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9840), .S(n9858), .Z(
        P1_U3585) );
  MUX2_X1 U11056 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9841), .S(n9858), .Z(
        P1_U3584) );
  MUX2_X1 U11057 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9966), .S(n9858), .Z(
        P1_U3583) );
  MUX2_X1 U11058 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9842), .S(n9858), .Z(
        P1_U3582) );
  MUX2_X1 U11059 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9843), .S(n9858), .Z(
        P1_U3581) );
  MUX2_X1 U11060 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n10001), .S(n9858), .Z(
        P1_U3580) );
  MUX2_X1 U11061 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9844), .S(n9858), .Z(
        P1_U3579) );
  MUX2_X1 U11062 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n10039), .S(n9858), .Z(
        P1_U3578) );
  MUX2_X1 U11063 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n10048), .S(n9858), .Z(
        P1_U3577) );
  MUX2_X1 U11064 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n4836), .S(n9858), .Z(
        P1_U3576) );
  MUX2_X1 U11065 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n10047), .S(n9858), .Z(
        P1_U3575) );
  MUX2_X1 U11066 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n10094), .S(n9858), .Z(
        P1_U3574) );
  MUX2_X1 U11067 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n10115), .S(n9858), .Z(
        P1_U3573) );
  MUX2_X1 U11068 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n10095), .S(n9858), .Z(
        P1_U3572) );
  MUX2_X1 U11069 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9845), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U11070 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n10146), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U11071 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9846), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U11072 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9847), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U11073 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9848), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U11074 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9849), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U11075 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9850), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U11076 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9851), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U11077 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9852), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U11078 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9853), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U11079 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n4505), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U11080 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9854), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U11081 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9855), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U11082 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9856), .S(n9858), .Z(
        P1_U3557) );
  MUX2_X1 U11083 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9857), .S(n9858), .Z(
        P1_U3556) );
  MUX2_X1 U11084 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9859), .S(n9858), .Z(
        P1_U3555) );
  XNOR2_X1 U11085 ( .A(n9884), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9873) );
  XNOR2_X1 U11086 ( .A(n9874), .B(n9873), .ZN(n9861) );
  NAND2_X1 U11087 ( .A1(n10427), .A2(n9861), .ZN(n9862) );
  OAI211_X1 U11088 ( .C1(n10393), .C2(n9884), .A(n9863), .B(n9862), .ZN(n9871)
         );
  AND2_X1 U11089 ( .A1(n9864), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9865) );
  XNOR2_X1 U11090 ( .A(n9885), .B(n9867), .ZN(n9869) );
  INV_X1 U11091 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9868) );
  NAND2_X1 U11092 ( .A1(n9869), .A2(n9868), .ZN(n9887) );
  AOI221_X1 U11093 ( .B1(n9869), .B2(n9887), .C1(n9868), .C2(n9887), .A(n10416), .ZN(n9870) );
  AOI211_X1 U11094 ( .C1(n10410), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n9871), .B(
        n9870), .ZN(n9872) );
  INV_X1 U11095 ( .A(n9872), .ZN(P1_U3255) );
  NAND2_X1 U11096 ( .A1(n9874), .A2(n9873), .ZN(n9877) );
  INV_X1 U11097 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9875) );
  NAND2_X1 U11098 ( .A1(n9884), .A2(n9875), .ZN(n9876) );
  INV_X1 U11099 ( .A(n9878), .ZN(n9881) );
  INV_X1 U11100 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9879) );
  INV_X1 U11101 ( .A(n9902), .ZN(n9880) );
  OAI211_X1 U11102 ( .C1(n9881), .C2(P1_REG1_REG_15__SCAN_IN), .A(n10427), .B(
        n9880), .ZN(n9882) );
  OAI211_X1 U11103 ( .C1(n10393), .C2(n9889), .A(n9883), .B(n9882), .ZN(n9893)
         );
  INV_X1 U11104 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9891) );
  NAND2_X1 U11105 ( .A1(n9885), .A2(n9884), .ZN(n9886) );
  AOI211_X1 U11106 ( .C1(n9891), .C2(n9890), .A(n9897), .B(n10416), .ZN(n9892)
         );
  AOI211_X1 U11107 ( .C1(n10410), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n9893), .B(
        n9892), .ZN(n9894) );
  INV_X1 U11108 ( .A(n9894), .ZN(P1_U3256) );
  NOR2_X1 U11109 ( .A1(n9889), .A2(n9895), .ZN(n9896) );
  NAND2_X1 U11110 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9917), .ZN(n9898) );
  OAI21_X1 U11111 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9917), .A(n9898), .ZN(
        n9899) );
  AOI211_X1 U11112 ( .C1(n9900), .C2(n9899), .A(n4457), .B(n10416), .ZN(n9911)
         );
  NOR2_X1 U11113 ( .A1(n9889), .A2(n9901), .ZN(n9903) );
  XNOR2_X1 U11114 ( .A(n9917), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9904) );
  NOR2_X1 U11115 ( .A1(n9905), .A2(n9904), .ZN(n9916) );
  AOI211_X1 U11116 ( .C1(n9905), .C2(n9904), .A(n9916), .B(n10394), .ZN(n9910)
         );
  NAND2_X1 U11117 ( .A1(n10410), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9907) );
  OAI211_X1 U11118 ( .C1(n10393), .C2(n9908), .A(n9907), .B(n9906), .ZN(n9909)
         );
  OR3_X1 U11119 ( .A1(n9911), .A2(n9910), .A3(n9909), .ZN(P1_U3257) );
  AOI22_X1 U11120 ( .A1(n9932), .A2(n7976), .B1(P1_REG2_REG_17__SCAN_IN), .B2(
        n9912), .ZN(n9913) );
  AOI211_X1 U11121 ( .C1(n9914), .C2(n9913), .A(n9934), .B(n10416), .ZN(n9915)
         );
  INV_X1 U11122 ( .A(n9915), .ZN(n9923) );
  AOI21_X1 U11123 ( .B1(n9917), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9916), .ZN(
        n9919) );
  XNOR2_X1 U11124 ( .A(n9932), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9918) );
  NOR2_X1 U11125 ( .A1(n9919), .A2(n9918), .ZN(n9925) );
  AOI211_X1 U11126 ( .C1(n9919), .C2(n9918), .A(n9925), .B(n10394), .ZN(n9920)
         );
  AOI211_X1 U11127 ( .C1(n10423), .C2(n9932), .A(n9921), .B(n9920), .ZN(n9922)
         );
  OAI211_X1 U11128 ( .C1(n10431), .C2(n8612), .A(n9923), .B(n9922), .ZN(
        P1_U3258) );
  XNOR2_X1 U11129 ( .A(n9944), .B(n9924), .ZN(n9927) );
  OAI21_X1 U11130 ( .B1(n9927), .B2(n9926), .A(n9943), .ZN(n9928) );
  NAND2_X1 U11131 ( .A1(n10427), .A2(n9928), .ZN(n9929) );
  OAI211_X1 U11132 ( .C1(n10393), .C2(n9931), .A(n9930), .B(n9929), .ZN(n9939)
         );
  AND2_X1 U11133 ( .A1(n9932), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9933) );
  NAND2_X1 U11134 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n9944), .ZN(n9935) );
  OAI21_X1 U11135 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9944), .A(n9935), .ZN(
        n9936) );
  NOR2_X1 U11136 ( .A1(n9937), .A2(n9936), .ZN(n9941) );
  AOI211_X1 U11137 ( .C1(n9937), .C2(n9936), .A(n9941), .B(n10416), .ZN(n9938)
         );
  AOI211_X1 U11138 ( .C1(n10410), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9939), .B(
        n9938), .ZN(n9940) );
  INV_X1 U11139 ( .A(n9940), .ZN(P1_U3259) );
  AOI21_X1 U11140 ( .B1(n9944), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9941), .ZN(
        n9942) );
  XNOR2_X1 U11141 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9942), .ZN(n9949) );
  AOI22_X1 U11142 ( .A1(n9949), .A2(n9946), .B1(n10427), .B2(n9947), .ZN(n9952) );
  INV_X1 U11143 ( .A(n9947), .ZN(n9950) );
  OAI21_X1 U11144 ( .B1(n10139), .B2(n9958), .A(n9957), .ZN(n9959) );
  AOI21_X1 U11145 ( .B1(n10197), .B2(n9960), .A(n9959), .ZN(n9961) );
  OAI21_X1 U11146 ( .B1(n10199), .B2(n10434), .A(n9961), .ZN(P1_U3262) );
  OAI211_X1 U11147 ( .C1(n9965), .C2(n9964), .A(n9963), .B(n10117), .ZN(n9968)
         );
  NAND2_X1 U11148 ( .A1(n9966), .A2(n10148), .ZN(n9967) );
  INV_X1 U11149 ( .A(n9981), .ZN(n9972) );
  INV_X1 U11150 ( .A(n9970), .ZN(n9971) );
  NAND2_X1 U11151 ( .A1(n10213), .A2(n10071), .ZN(n9975) );
  AOI22_X1 U11152 ( .A1(n9973), .A2(n10170), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10437), .ZN(n9974) );
  OAI211_X1 U11153 ( .C1(n9976), .C2(n10433), .A(n9975), .B(n9974), .ZN(n9977)
         );
  AOI21_X1 U11154 ( .B1(n10212), .B2(n10139), .A(n9977), .ZN(n9978) );
  OAI21_X1 U11155 ( .B1(n10216), .B2(n10192), .A(n9978), .ZN(P1_U3264) );
  XOR2_X1 U11156 ( .A(n9979), .B(n9990), .Z(n10221) );
  INV_X1 U11157 ( .A(n9980), .ZN(n9982) );
  AOI211_X1 U11158 ( .C1(n10219), .C2(n9982), .A(n10456), .B(n9981), .ZN(
        n10218) );
  NOR2_X1 U11159 ( .A1(n9983), .A2(n10433), .ZN(n9987) );
  OAI22_X1 U11160 ( .A1(n9985), .A2(n10439), .B1(n9984), .B2(n10139), .ZN(
        n9986) );
  AOI211_X1 U11161 ( .C1(n10218), .C2(n10071), .A(n9987), .B(n9986), .ZN(n9996) );
  NAND2_X1 U11162 ( .A1(n9989), .A2(n9988), .ZN(n9991) );
  XNOR2_X1 U11163 ( .A(n9991), .B(n9990), .ZN(n9992) );
  OAI222_X1 U11164 ( .A1(n10184), .A2(n9994), .B1(n10182), .B2(n9993), .C1(
        n9992), .C2(n10179), .ZN(n10217) );
  NAND2_X1 U11165 ( .A1(n10217), .A2(n10011), .ZN(n9995) );
  OAI211_X1 U11166 ( .C1(n10221), .C2(n10192), .A(n9996), .B(n9995), .ZN(
        P1_U3265) );
  XNOR2_X1 U11167 ( .A(n9997), .B(n9999), .ZN(n10231) );
  OAI211_X1 U11168 ( .C1(n10000), .C2(n9999), .A(n9998), .B(n10117), .ZN(
        n10003) );
  NAND2_X1 U11169 ( .A1(n10001), .A2(n10148), .ZN(n10002) );
  OAI211_X1 U11170 ( .C1(n10004), .C2(n10182), .A(n10003), .B(n10002), .ZN(
        n10227) );
  AOI211_X1 U11171 ( .C1(n10229), .C2(n10019), .A(n10456), .B(n7893), .ZN(
        n10228) );
  NAND2_X1 U11172 ( .A1(n10228), .A2(n10071), .ZN(n10008) );
  AOI22_X1 U11173 ( .A1(n10006), .A2(n10170), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10437), .ZN(n10007) );
  OAI211_X1 U11174 ( .C1(n10009), .C2(n10433), .A(n10008), .B(n10007), .ZN(
        n10010) );
  AOI21_X1 U11175 ( .B1(n10227), .B2(n10011), .A(n10010), .ZN(n10012) );
  OAI21_X1 U11176 ( .B1(n10231), .B2(n10192), .A(n10012), .ZN(P1_U3267) );
  AOI21_X1 U11177 ( .B1(n4862), .B2(n10013), .A(n10179), .ZN(n10018) );
  OAI22_X1 U11178 ( .A1(n10015), .A2(n10184), .B1(n10014), .B2(n10182), .ZN(
        n10016) );
  AOI21_X1 U11179 ( .B1(n10018), .B2(n10017), .A(n10016), .ZN(n10235) );
  OR2_X1 U11180 ( .A1(n10032), .A2(n10023), .ZN(n10020) );
  AND2_X1 U11181 ( .A1(n10020), .A2(n10019), .ZN(n10233) );
  AOI22_X1 U11182 ( .A1(n10021), .A2(n10170), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10437), .ZN(n10022) );
  OAI21_X1 U11183 ( .B1(n10023), .B2(n10433), .A(n10022), .ZN(n10029) );
  INV_X1 U11184 ( .A(n10024), .ZN(n10025) );
  AOI21_X1 U11185 ( .B1(n10027), .B2(n10026), .A(n10025), .ZN(n10236) );
  NOR2_X1 U11186 ( .A1(n10236), .A2(n10192), .ZN(n10028) );
  AOI211_X1 U11187 ( .C1(n10233), .C2(n10156), .A(n10029), .B(n10028), .ZN(
        n10030) );
  OAI21_X1 U11188 ( .B1(n10437), .B2(n10235), .A(n10030), .ZN(P1_U3268) );
  XOR2_X1 U11189 ( .A(n10031), .B(n10038), .Z(n10241) );
  AOI21_X1 U11190 ( .B1(n10237), .B2(n10050), .A(n10032), .ZN(n10238) );
  INV_X1 U11191 ( .A(n10033), .ZN(n10034) );
  AOI22_X1 U11192 ( .A1(n10034), .A2(n10170), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10437), .ZN(n10035) );
  OAI21_X1 U11193 ( .B1(n10036), .B2(n10433), .A(n10035), .ZN(n10042) );
  XOR2_X1 U11194 ( .A(n10038), .B(n10037), .Z(n10040) );
  AOI222_X1 U11195 ( .A1(n10117), .A2(n10040), .B1(n10039), .B2(n10148), .C1(
        n4836), .C2(n10147), .ZN(n10240) );
  NOR2_X1 U11196 ( .A1(n10240), .A2(n10437), .ZN(n10041) );
  AOI211_X1 U11197 ( .C1(n10238), .C2(n10156), .A(n10042), .B(n10041), .ZN(
        n10043) );
  OAI21_X1 U11198 ( .B1(n10192), .B2(n10241), .A(n10043), .ZN(P1_U3269) );
  XNOR2_X1 U11199 ( .A(n10044), .B(n4720), .ZN(n10246) );
  OAI21_X1 U11200 ( .B1(n10046), .B2(n4720), .A(n4504), .ZN(n10049) );
  AOI222_X1 U11201 ( .A1(n10117), .A2(n10049), .B1(n10048), .B2(n10148), .C1(
        n10047), .C2(n10147), .ZN(n10245) );
  AOI21_X1 U11202 ( .B1(n10065), .B2(n10243), .A(n10456), .ZN(n10051) );
  AND2_X1 U11203 ( .A1(n10051), .A2(n10050), .ZN(n10242) );
  AOI22_X1 U11204 ( .A1(n10242), .A2(n10053), .B1(n10170), .B2(n10052), .ZN(
        n10054) );
  AOI21_X1 U11205 ( .B1(n10245), .B2(n10054), .A(n10437), .ZN(n10057) );
  OAI22_X1 U11206 ( .A1(n4834), .A2(n10433), .B1(n10139), .B2(n10055), .ZN(
        n10056) );
  NOR2_X1 U11207 ( .A1(n10057), .A2(n10056), .ZN(n10058) );
  OAI21_X1 U11208 ( .B1(n10246), .B2(n10192), .A(n10058), .ZN(P1_U3270) );
  XOR2_X1 U11209 ( .A(n4518), .B(n10060), .Z(n10251) );
  XNOR2_X1 U11210 ( .A(n10061), .B(n10060), .ZN(n10062) );
  OAI222_X1 U11211 ( .A1(n10184), .A2(n10064), .B1(n10182), .B2(n10063), .C1(
        n10179), .C2(n10062), .ZN(n10247) );
  NAND2_X1 U11212 ( .A1(n10247), .A2(n10139), .ZN(n10073) );
  AOI211_X1 U11213 ( .C1(n10249), .C2(n10081), .A(n10456), .B(n4912), .ZN(
        n10248) );
  NOR2_X1 U11214 ( .A1(n10066), .A2(n10433), .ZN(n10070) );
  OAI22_X1 U11215 ( .A1(n10068), .A2(n10139), .B1(n10067), .B2(n10439), .ZN(
        n10069) );
  AOI211_X1 U11216 ( .C1(n10248), .C2(n10071), .A(n10070), .B(n10069), .ZN(
        n10072) );
  OAI211_X1 U11217 ( .C1(n10251), .C2(n10192), .A(n10073), .B(n10072), .ZN(
        P1_U3271) );
  NAND2_X1 U11218 ( .A1(n10105), .A2(n10104), .ZN(n10261) );
  NAND2_X1 U11219 ( .A1(n10261), .A2(n10074), .ZN(n10075) );
  XNOR2_X1 U11220 ( .A(n10075), .B(n10077), .ZN(n10257) );
  AOI21_X1 U11221 ( .B1(n10077), .B2(n10076), .A(n4430), .ZN(n10078) );
  OAI222_X1 U11222 ( .A1(n10184), .A2(n10080), .B1(n10182), .B2(n10079), .C1(
        n10179), .C2(n10078), .ZN(n10252) );
  INV_X1 U11223 ( .A(n10097), .ZN(n10083) );
  INV_X1 U11224 ( .A(n10081), .ZN(n10082) );
  AOI21_X1 U11225 ( .B1(n10253), .B2(n10083), .A(n10082), .ZN(n10254) );
  NAND2_X1 U11226 ( .A1(n10254), .A2(n10156), .ZN(n10086) );
  AOI22_X1 U11227 ( .A1(n10437), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n10084), 
        .B2(n10170), .ZN(n10085) );
  OAI211_X1 U11228 ( .C1(n10087), .C2(n10433), .A(n10086), .B(n10085), .ZN(
        n10088) );
  AOI21_X1 U11229 ( .B1(n10252), .B2(n10139), .A(n10088), .ZN(n10089) );
  OAI21_X1 U11230 ( .B1(n10192), .B2(n10257), .A(n10089), .ZN(P1_U3272) );
  INV_X1 U11231 ( .A(n10090), .ZN(n10092) );
  OAI21_X1 U11232 ( .B1(n10114), .B2(n10092), .A(n10091), .ZN(n10093) );
  XNOR2_X1 U11233 ( .A(n10093), .B(n10104), .ZN(n10096) );
  AOI222_X1 U11234 ( .A1(n10117), .A2(n10096), .B1(n10095), .B2(n10147), .C1(
        n10094), .C2(n10148), .ZN(n10265) );
  INV_X1 U11235 ( .A(n10109), .ZN(n10098) );
  AOI21_X1 U11236 ( .B1(n10258), .B2(n10098), .A(n10097), .ZN(n10259) );
  NOR2_X1 U11237 ( .A1(n10099), .A2(n10433), .ZN(n10103) );
  OAI22_X1 U11238 ( .A1(n10139), .A2(n10101), .B1(n10100), .B2(n10439), .ZN(
        n10102) );
  AOI211_X1 U11239 ( .C1(n10259), .C2(n10156), .A(n10103), .B(n10102), .ZN(
        n10107) );
  OR2_X1 U11240 ( .A1(n10105), .A2(n10104), .ZN(n10262) );
  NAND3_X1 U11241 ( .A1(n10262), .A2(n10261), .A3(n4524), .ZN(n10106) );
  OAI211_X1 U11242 ( .C1(n10265), .C2(n10437), .A(n10107), .B(n10106), .ZN(
        P1_U3273) );
  XOR2_X1 U11243 ( .A(n10108), .B(n10113), .Z(n10270) );
  OR2_X1 U11244 ( .A1(n10154), .A2(n10273), .ZN(n10132) );
  AOI21_X1 U11245 ( .B1(n10266), .B2(n10132), .A(n10109), .ZN(n10267) );
  AOI22_X1 U11246 ( .A1(n10437), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n10110), 
        .B2(n10170), .ZN(n10111) );
  OAI21_X1 U11247 ( .B1(n10112), .B2(n10433), .A(n10111), .ZN(n10119) );
  XNOR2_X1 U11248 ( .A(n10114), .B(n10113), .ZN(n10116) );
  AOI222_X1 U11249 ( .A1(n10117), .A2(n10116), .B1(n10115), .B2(n10148), .C1(
        n10149), .C2(n10147), .ZN(n10269) );
  NOR2_X1 U11250 ( .A1(n10269), .A2(n10437), .ZN(n10118) );
  AOI211_X1 U11251 ( .C1(n10267), .C2(n10156), .A(n10119), .B(n10118), .ZN(
        n10120) );
  OAI21_X1 U11252 ( .B1(n10192), .B2(n10270), .A(n10120), .ZN(P1_U3274) );
  INV_X1 U11253 ( .A(n10121), .ZN(n10142) );
  NAND2_X1 U11254 ( .A1(n10142), .A2(n10145), .ZN(n10141) );
  NAND2_X1 U11255 ( .A1(n10141), .A2(n10122), .ZN(n10123) );
  XNOR2_X1 U11256 ( .A(n10123), .B(n10128), .ZN(n10275) );
  NAND2_X1 U11257 ( .A1(n10125), .A2(n10124), .ZN(n10144) );
  NOR2_X1 U11258 ( .A1(n10144), .A2(n10145), .ZN(n10143) );
  INV_X1 U11259 ( .A(n10126), .ZN(n10127) );
  NOR2_X1 U11260 ( .A1(n10143), .A2(n10127), .ZN(n10129) );
  XNOR2_X1 U11261 ( .A(n10129), .B(n10128), .ZN(n10130) );
  OAI222_X1 U11262 ( .A1(n10184), .A2(n10131), .B1(n10182), .B2(n10185), .C1(
        n10130), .C2(n10179), .ZN(n10271) );
  INV_X1 U11263 ( .A(n10132), .ZN(n10133) );
  AOI211_X1 U11264 ( .C1(n10273), .C2(n10154), .A(n10456), .B(n10133), .ZN(
        n10272) );
  NAND2_X1 U11265 ( .A1(n10272), .A2(n10190), .ZN(n10136) );
  AOI22_X1 U11266 ( .A1(n10437), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n10134), 
        .B2(n10170), .ZN(n10135) );
  OAI211_X1 U11267 ( .C1(n10137), .C2(n10433), .A(n10136), .B(n10135), .ZN(
        n10138) );
  AOI21_X1 U11268 ( .B1(n10271), .B2(n10139), .A(n10138), .ZN(n10140) );
  OAI21_X1 U11269 ( .B1(n10275), .B2(n10192), .A(n10140), .ZN(P1_U3275) );
  OAI21_X1 U11270 ( .B1(n10142), .B2(n10145), .A(n10141), .ZN(n10276) );
  AOI21_X1 U11271 ( .B1(n10145), .B2(n10144), .A(n10143), .ZN(n10151) );
  AOI22_X1 U11272 ( .A1(n10149), .A2(n10148), .B1(n10147), .B2(n10146), .ZN(
        n10150) );
  OAI21_X1 U11273 ( .B1(n10151), .B2(n10179), .A(n10150), .ZN(n10152) );
  AOI21_X1 U11274 ( .B1(n10153), .B2(n10276), .A(n10152), .ZN(n10280) );
  INV_X1 U11275 ( .A(n10167), .ZN(n10155) );
  AOI21_X1 U11276 ( .B1(n10277), .B2(n10155), .A(n4913), .ZN(n10278) );
  NAND2_X1 U11277 ( .A1(n10278), .A2(n10156), .ZN(n10160) );
  INV_X1 U11278 ( .A(n10157), .ZN(n10158) );
  AOI22_X1 U11279 ( .A1(n10437), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n10158), 
        .B2(n10170), .ZN(n10159) );
  OAI211_X1 U11280 ( .C1(n10161), .C2(n10433), .A(n10160), .B(n10159), .ZN(
        n10162) );
  AOI21_X1 U11281 ( .B1(n10276), .B2(n4484), .A(n10162), .ZN(n10164) );
  OAI21_X1 U11282 ( .B1(n10280), .B2(n10437), .A(n10164), .ZN(P1_U3276) );
  XNOR2_X1 U11283 ( .A(n10165), .B(n10176), .ZN(n10286) );
  INV_X1 U11284 ( .A(n10166), .ZN(n10168) );
  AOI211_X1 U11285 ( .C1(n10283), .C2(n10168), .A(n10456), .B(n10167), .ZN(
        n10282) );
  INV_X1 U11286 ( .A(n10169), .ZN(n10171) );
  AOI22_X1 U11287 ( .A1(n10437), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n10171), 
        .B2(n10170), .ZN(n10172) );
  OAI21_X1 U11288 ( .B1(n10173), .B2(n10433), .A(n10172), .ZN(n10189) );
  INV_X1 U11289 ( .A(n10176), .ZN(n10175) );
  NOR2_X1 U11290 ( .A1(n10175), .A2(n10174), .ZN(n10181) );
  AOI21_X1 U11291 ( .B1(n10180), .B2(n10177), .A(n10176), .ZN(n10178) );
  AOI211_X1 U11292 ( .C1(n10181), .C2(n10180), .A(n10179), .B(n10178), .ZN(
        n10187) );
  OAI22_X1 U11293 ( .A1(n10185), .A2(n10184), .B1(n10183), .B2(n10182), .ZN(
        n10186) );
  NOR2_X1 U11294 ( .A1(n10187), .A2(n10186), .ZN(n10285) );
  NOR2_X1 U11295 ( .A1(n10285), .A2(n10437), .ZN(n10188) );
  AOI211_X1 U11296 ( .C1(n10190), .C2(n10282), .A(n10189), .B(n10188), .ZN(
        n10191) );
  OAI21_X1 U11297 ( .B1(n10192), .B2(n10286), .A(n10191), .ZN(P1_U3277) );
  AOI21_X1 U11298 ( .B1(n10193), .B2(n10306), .A(n10196), .ZN(n10194) );
  OAI21_X1 U11299 ( .B1(n10195), .B2(n10456), .A(n10194), .ZN(n10314) );
  MUX2_X1 U11300 ( .A(n10314), .B(P1_REG1_REG_31__SCAN_IN), .S(n10463), .Z(
        P1_U3554) );
  AOI21_X1 U11301 ( .B1(n10197), .B2(n10306), .A(n10196), .ZN(n10198) );
  MUX2_X1 U11302 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10315), .S(n10465), .Z(
        P1_U3553) );
  NAND2_X1 U11303 ( .A1(n10200), .A2(n10260), .ZN(n10206) );
  AOI22_X1 U11304 ( .A1(n10202), .A2(n10307), .B1(n10306), .B2(n10201), .ZN(
        n10203) );
  NAND2_X1 U11305 ( .A1(n10206), .A2(n10205), .ZN(n10316) );
  MUX2_X1 U11306 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10316), .S(n10465), .Z(
        P1_U3552) );
  AOI22_X1 U11307 ( .A1(n10208), .A2(n10307), .B1(n10306), .B2(n10207), .ZN(
        n10209) );
  OAI211_X1 U11308 ( .C1(n10211), .C2(n10298), .A(n10210), .B(n10209), .ZN(
        n10317) );
  MUX2_X1 U11309 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10317), .S(n10465), .Z(
        P1_U3551) );
  OAI21_X1 U11310 ( .B1(n10298), .B2(n10216), .A(n10215), .ZN(n10318) );
  MUX2_X1 U11311 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10318), .S(n10465), .Z(
        P1_U3550) );
  OAI21_X1 U11312 ( .B1(n10298), .B2(n10221), .A(n10220), .ZN(n10319) );
  MUX2_X1 U11313 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10319), .S(n10465), .Z(
        P1_U3549) );
  AOI22_X1 U11314 ( .A1(n10223), .A2(n10307), .B1(n10306), .B2(n10222), .ZN(
        n10224) );
  OAI211_X1 U11315 ( .C1(n10298), .C2(n10226), .A(n10225), .B(n10224), .ZN(
        n10320) );
  MUX2_X1 U11316 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10320), .S(n10465), .Z(
        P1_U3548) );
  AOI211_X1 U11317 ( .C1(n10306), .C2(n10229), .A(n10228), .B(n10227), .ZN(
        n10230) );
  OAI21_X1 U11318 ( .B1(n10298), .B2(n10231), .A(n10230), .ZN(n10321) );
  MUX2_X1 U11319 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10321), .S(n10465), .Z(
        P1_U3547) );
  AOI22_X1 U11320 ( .A1(n10233), .A2(n10307), .B1(n10306), .B2(n10232), .ZN(
        n10234) );
  OAI211_X1 U11321 ( .C1(n10236), .C2(n10298), .A(n10235), .B(n10234), .ZN(
        n10322) );
  MUX2_X1 U11322 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10322), .S(n10465), .Z(
        P1_U3546) );
  AOI22_X1 U11323 ( .A1(n10238), .A2(n10307), .B1(n10306), .B2(n10237), .ZN(
        n10239) );
  OAI211_X1 U11324 ( .C1(n10298), .C2(n10241), .A(n10240), .B(n10239), .ZN(
        n10323) );
  MUX2_X1 U11325 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10323), .S(n10465), .Z(
        P1_U3545) );
  AOI21_X1 U11326 ( .B1(n10306), .B2(n10243), .A(n10242), .ZN(n10244) );
  OAI211_X1 U11327 ( .C1(n10298), .C2(n10246), .A(n10245), .B(n10244), .ZN(
        n10324) );
  MUX2_X1 U11328 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10324), .S(n10465), .Z(
        P1_U3544) );
  AOI211_X1 U11329 ( .C1(n10306), .C2(n10249), .A(n10248), .B(n10247), .ZN(
        n10250) );
  OAI21_X1 U11330 ( .B1(n10298), .B2(n10251), .A(n10250), .ZN(n10325) );
  MUX2_X1 U11331 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10325), .S(n10465), .Z(
        P1_U3543) );
  INV_X1 U11332 ( .A(n10252), .ZN(n10256) );
  AOI22_X1 U11333 ( .A1(n10254), .A2(n10307), .B1(n10306), .B2(n10253), .ZN(
        n10255) );
  OAI211_X1 U11334 ( .C1(n10298), .C2(n10257), .A(n10256), .B(n10255), .ZN(
        n10326) );
  MUX2_X1 U11335 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10326), .S(n10465), .Z(
        P1_U3542) );
  AOI22_X1 U11336 ( .A1(n10259), .A2(n10307), .B1(n10306), .B2(n10258), .ZN(
        n10264) );
  NAND3_X1 U11337 ( .A1(n10262), .A2(n10261), .A3(n10260), .ZN(n10263) );
  NAND3_X1 U11338 ( .A1(n10265), .A2(n10264), .A3(n10263), .ZN(n10327) );
  MUX2_X1 U11339 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10327), .S(n10465), .Z(
        P1_U3541) );
  AOI22_X1 U11340 ( .A1(n10267), .A2(n10307), .B1(n10306), .B2(n10266), .ZN(
        n10268) );
  OAI211_X1 U11341 ( .C1(n10298), .C2(n10270), .A(n10269), .B(n10268), .ZN(
        n10328) );
  MUX2_X1 U11342 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10328), .S(n10465), .Z(
        P1_U3540) );
  AOI211_X1 U11343 ( .C1(n10306), .C2(n10273), .A(n10272), .B(n10271), .ZN(
        n10274) );
  OAI21_X1 U11344 ( .B1(n10298), .B2(n10275), .A(n10274), .ZN(n10329) );
  MUX2_X1 U11345 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10329), .S(n10465), .Z(
        P1_U3539) );
  INV_X1 U11346 ( .A(n10276), .ZN(n10281) );
  AOI22_X1 U11347 ( .A1(n10278), .A2(n10307), .B1(n10306), .B2(n10277), .ZN(
        n10279) );
  OAI211_X1 U11348 ( .C1(n10281), .C2(n10311), .A(n10280), .B(n10279), .ZN(
        n10330) );
  MUX2_X1 U11349 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10330), .S(n10465), .Z(
        P1_U3538) );
  AOI21_X1 U11350 ( .B1(n10306), .B2(n10283), .A(n10282), .ZN(n10284) );
  OAI211_X1 U11351 ( .C1(n10298), .C2(n10286), .A(n10285), .B(n10284), .ZN(
        n10331) );
  MUX2_X1 U11352 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10331), .S(n10465), .Z(
        P1_U3537) );
  INV_X1 U11353 ( .A(n10287), .ZN(n10292) );
  AOI22_X1 U11354 ( .A1(n10289), .A2(n10307), .B1(n10306), .B2(n10288), .ZN(
        n10290) );
  OAI211_X1 U11355 ( .C1(n10311), .C2(n10292), .A(n10291), .B(n10290), .ZN(
        n10332) );
  MUX2_X1 U11356 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10332), .S(n10465), .Z(
        P1_U3536) );
  AOI21_X1 U11357 ( .B1(n10306), .B2(n10294), .A(n10293), .ZN(n10295) );
  OAI211_X1 U11358 ( .C1(n10298), .C2(n10297), .A(n10296), .B(n10295), .ZN(
        n10333) );
  MUX2_X1 U11359 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10333), .S(n10465), .Z(
        P1_U3535) );
  INV_X1 U11360 ( .A(n10299), .ZN(n10304) );
  AOI21_X1 U11361 ( .B1(n10306), .B2(n10301), .A(n10300), .ZN(n10302) );
  OAI211_X1 U11362 ( .C1(n10304), .C2(n10311), .A(n10303), .B(n10302), .ZN(
        n10334) );
  MUX2_X1 U11363 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n10334), .S(n10465), .Z(
        P1_U3533) );
  AOI22_X1 U11364 ( .A1(n10308), .A2(n10307), .B1(n10306), .B2(n10305), .ZN(
        n10309) );
  OAI211_X1 U11365 ( .C1(n10312), .C2(n10311), .A(n10310), .B(n10309), .ZN(
        n10336) );
  MUX2_X1 U11366 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10336), .S(n10465), .Z(
        P1_U3532) );
  MUX2_X1 U11367 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n10313), .S(n10465), .Z(
        P1_U3523) );
  MUX2_X1 U11368 ( .A(n10314), .B(P1_REG0_REG_31__SCAN_IN), .S(n10462), .Z(
        P1_U3522) );
  MUX2_X1 U11369 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10315), .S(n10335), .Z(
        P1_U3521) );
  MUX2_X1 U11370 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10316), .S(n10335), .Z(
        P1_U3520) );
  MUX2_X1 U11371 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10317), .S(n10335), .Z(
        P1_U3519) );
  MUX2_X1 U11372 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10318), .S(n10335), .Z(
        P1_U3518) );
  MUX2_X1 U11373 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10319), .S(n10335), .Z(
        P1_U3517) );
  MUX2_X1 U11374 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10320), .S(n10335), .Z(
        P1_U3516) );
  MUX2_X1 U11375 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10321), .S(n10335), .Z(
        P1_U3515) );
  MUX2_X1 U11376 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10322), .S(n10335), .Z(
        P1_U3514) );
  MUX2_X1 U11377 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10323), .S(n10335), .Z(
        P1_U3513) );
  MUX2_X1 U11378 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10324), .S(n10335), .Z(
        P1_U3512) );
  MUX2_X1 U11379 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10325), .S(n10335), .Z(
        P1_U3511) );
  MUX2_X1 U11380 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10326), .S(n10335), .Z(
        P1_U3510) );
  MUX2_X1 U11381 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10327), .S(n10335), .Z(
        P1_U3508) );
  MUX2_X1 U11382 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10328), .S(n10335), .Z(
        P1_U3505) );
  MUX2_X1 U11383 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10329), .S(n10335), .Z(
        P1_U3502) );
  MUX2_X1 U11384 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10330), .S(n10335), .Z(
        P1_U3499) );
  MUX2_X1 U11385 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10331), .S(n10335), .Z(
        P1_U3496) );
  MUX2_X1 U11386 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n10332), .S(n10335), .Z(
        P1_U3493) );
  MUX2_X1 U11387 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n10333), .S(n10335), .Z(
        P1_U3490) );
  MUX2_X1 U11388 ( .A(P1_REG0_REG_10__SCAN_IN), .B(n10334), .S(n10335), .Z(
        P1_U3484) );
  MUX2_X1 U11389 ( .A(P1_REG0_REG_9__SCAN_IN), .B(n10336), .S(n10335), .Z(
        P1_U3481) );
  AND2_X1 U11390 ( .A1(n10453), .A2(n10337), .ZN(n10448) );
  MUX2_X1 U11391 ( .A(P1_D_REG_0__SCAN_IN), .B(n10338), .S(n10448), .Z(
        P1_U3440) );
  NOR4_X1 U11392 ( .A1(n6358), .A2(P1_IR_REG_30__SCAN_IN), .A3(n6218), .A4(
        P1_U3084), .ZN(n10339) );
  AOI21_X1 U11393 ( .B1(n10340), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10339), 
        .ZN(n10341) );
  OAI21_X1 U11394 ( .B1(n10342), .B2(n10347), .A(n10341), .ZN(P1_U3322) );
  OAI222_X1 U11395 ( .A1(n10350), .A2(n10345), .B1(n10347), .B2(n10344), .C1(
        n10343), .C2(P1_U3084), .ZN(P1_U3323) );
  OAI222_X1 U11396 ( .A1(n10350), .A2(n10349), .B1(P1_U3084), .B2(n10348), 
        .C1(n10347), .C2(n10346), .ZN(P1_U3324) );
  INV_X1 U11397 ( .A(n10351), .ZN(n10352) );
  MUX2_X1 U11398 ( .A(n10352), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NOR2_X1 U11399 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(P2_ADDR_REG_17__SCAN_IN), 
        .ZN(n10353) );
  AOI21_X1 U11400 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10353), .ZN(n10530) );
  NOR2_X1 U11401 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10354) );
  AOI21_X1 U11402 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10354), .ZN(n10533) );
  NOR2_X1 U11403 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10355) );
  AOI21_X1 U11404 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10355), .ZN(n10536) );
  NOR2_X1 U11405 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10356) );
  AOI21_X1 U11406 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10356), .ZN(n10539) );
  NOR2_X1 U11407 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10357) );
  AOI21_X1 U11408 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10357), .ZN(n10542) );
  NOR2_X1 U11409 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10365) );
  XNOR2_X1 U11410 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10569) );
  NAND2_X1 U11411 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n10363) );
  NAND2_X1 U11412 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10361) );
  AOI21_X1 U11413 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10523) );
  NAND3_X1 U11414 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10525) );
  OAI21_X1 U11415 ( .B1(n10523), .B2(n10527), .A(n10525), .ZN(n10564) );
  NAND2_X1 U11416 ( .A1(n10565), .A2(n10564), .ZN(n10360) );
  NAND2_X1 U11417 ( .A1(n10361), .A2(n10360), .ZN(n10566) );
  NAND2_X1 U11418 ( .A1(n10567), .A2(n10566), .ZN(n10362) );
  NAND2_X1 U11419 ( .A1(n10363), .A2(n10362), .ZN(n10568) );
  NOR2_X1 U11420 ( .A1(n10569), .A2(n10568), .ZN(n10364) );
  NOR2_X1 U11421 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10366), .ZN(n10554) );
  NAND2_X1 U11422 ( .A1(n10368), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n10370) );
  NAND2_X1 U11423 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10552), .ZN(n10369) );
  NAND2_X1 U11424 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n10371), .ZN(n10373) );
  NAND2_X1 U11425 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10563), .ZN(n10372) );
  NAND2_X1 U11426 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n10374), .ZN(n10376) );
  NAND2_X1 U11427 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10562), .ZN(n10375) );
  AND2_X1 U11428 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10377), .ZN(n10378) );
  NAND2_X1 U11429 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n10379) );
  OAI21_X1 U11430 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10379), .ZN(n10550) );
  NAND2_X1 U11431 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n10380) );
  OAI21_X1 U11432 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10380), .ZN(n10547) );
  NOR2_X1 U11433 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10381) );
  AOI21_X1 U11434 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10381), .ZN(n10544) );
  NAND2_X1 U11435 ( .A1(n10542), .A2(n10541), .ZN(n10540) );
  NAND2_X1 U11436 ( .A1(n10536), .A2(n10535), .ZN(n10534) );
  OAI21_X1 U11437 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10534), .ZN(n10532) );
  NAND2_X1 U11438 ( .A1(n10533), .A2(n10532), .ZN(n10531) );
  NAND2_X1 U11439 ( .A1(n10530), .A2(n10529), .ZN(n10528) );
  NOR2_X1 U11440 ( .A1(n10558), .A2(n10557), .ZN(n10382) );
  NAND2_X1 U11441 ( .A1(n10558), .A2(n10557), .ZN(n10556) );
  XNOR2_X1 U11442 ( .A(n4660), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n10383) );
  XNOR2_X1 U11443 ( .A(n10384), .B(n10383), .ZN(ADD_1071_U4) );
  XNOR2_X1 U11444 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11445 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  AND2_X1 U11446 ( .A1(n10386), .A2(n10385), .ZN(n10387) );
  NOR2_X1 U11447 ( .A1(n10388), .A2(n10387), .ZN(n10401) );
  AOI21_X1 U11448 ( .B1(n10391), .B2(n10390), .A(n10389), .ZN(n10395) );
  OAI22_X1 U11449 ( .A1(n10395), .A2(n10394), .B1(n10393), .B2(n10392), .ZN(
        n10398) );
  INV_X1 U11450 ( .A(n10396), .ZN(n10397) );
  AOI211_X1 U11451 ( .C1(n10410), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n10398), .B(
        n10397), .ZN(n10400) );
  OAI211_X1 U11452 ( .C1(n10401), .C2(n10416), .A(n10400), .B(n10399), .ZN(
        P1_U3245) );
  XOR2_X1 U11453 ( .A(n10402), .B(n10409), .Z(n10403) );
  XNOR2_X1 U11454 ( .A(n10404), .B(n10403), .ZN(n10414) );
  OR3_X1 U11455 ( .A1(n4477), .A2(n10406), .A3(n10405), .ZN(n10407) );
  NAND2_X1 U11456 ( .A1(n10408), .A2(n10407), .ZN(n10411) );
  AOI222_X1 U11457 ( .A1(n10411), .A2(n10427), .B1(n10410), .B2(
        P1_ADDR_REG_7__SCAN_IN), .C1(n10409), .C2(n10423), .ZN(n10413) );
  OAI211_X1 U11458 ( .C1(n10416), .C2(n10414), .A(n10413), .B(n10412), .ZN(
        P1_U3248) );
  INV_X1 U11459 ( .A(n10415), .ZN(n10421) );
  AOI211_X1 U11460 ( .C1(n10419), .C2(n10418), .A(n10417), .B(n10416), .ZN(
        n10420) );
  AOI211_X1 U11461 ( .C1(n10423), .C2(n10422), .A(n10421), .B(n10420), .ZN(
        n10429) );
  XNOR2_X1 U11462 ( .A(n10425), .B(n10424), .ZN(n10426) );
  NAND2_X1 U11463 ( .A1(n10427), .A2(n10426), .ZN(n10428) );
  OAI211_X1 U11464 ( .C1(n10431), .C2(n10430), .A(n10429), .B(n10428), .ZN(
        P1_U3251) );
  NOR2_X1 U11465 ( .A1(n10432), .A2(n10437), .ZN(n10436) );
  AOI21_X1 U11466 ( .B1(n10434), .B2(n10433), .A(n6373), .ZN(n10435) );
  AOI211_X1 U11467 ( .C1(n10437), .C2(P1_REG2_REG_0__SCAN_IN), .A(n10436), .B(
        n10435), .ZN(n10438) );
  OAI21_X1 U11468 ( .B1(n10439), .B2(n6253), .A(n10438), .ZN(P1_U3291) );
  AND2_X1 U11469 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10449), .ZN(P1_U3292) );
  AND2_X1 U11470 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10449), .ZN(P1_U3293) );
  AND2_X1 U11471 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10449), .ZN(P1_U3294) );
  AND2_X1 U11472 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10449), .ZN(P1_U3295) );
  NOR2_X1 U11473 ( .A1(n10448), .A2(n10440), .ZN(P1_U3296) );
  AND2_X1 U11474 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10449), .ZN(P1_U3297) );
  AND2_X1 U11475 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10449), .ZN(P1_U3298) );
  AND2_X1 U11476 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10449), .ZN(P1_U3299) );
  AND2_X1 U11477 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10449), .ZN(P1_U3300) );
  AND2_X1 U11478 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10449), .ZN(P1_U3301) );
  AND2_X1 U11479 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10449), .ZN(P1_U3302) );
  AND2_X1 U11480 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10449), .ZN(P1_U3303) );
  NOR2_X1 U11481 ( .A1(n10448), .A2(n10441), .ZN(P1_U3304) );
  AND2_X1 U11482 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10449), .ZN(P1_U3305) );
  AND2_X1 U11483 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10449), .ZN(P1_U3306) );
  AND2_X1 U11484 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10449), .ZN(P1_U3307) );
  NOR2_X1 U11485 ( .A1(n10448), .A2(n10442), .ZN(P1_U3308) );
  AND2_X1 U11486 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10449), .ZN(P1_U3309) );
  AND2_X1 U11487 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10449), .ZN(P1_U3310) );
  NOR2_X1 U11488 ( .A1(n10448), .A2(n10443), .ZN(P1_U3311) );
  AND2_X1 U11489 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10449), .ZN(P1_U3312) );
  NOR2_X1 U11490 ( .A1(n10448), .A2(n10444), .ZN(P1_U3313) );
  AND2_X1 U11491 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10449), .ZN(P1_U3314) );
  NOR2_X1 U11492 ( .A1(n10448), .A2(n10445), .ZN(P1_U3315) );
  AND2_X1 U11493 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10449), .ZN(P1_U3316) );
  AND2_X1 U11494 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10449), .ZN(P1_U3317) );
  NOR2_X1 U11495 ( .A1(n10448), .A2(n10446), .ZN(P1_U3318) );
  NOR2_X1 U11496 ( .A1(n10448), .A2(n10447), .ZN(P1_U3319) );
  AND2_X1 U11497 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10449), .ZN(P1_U3320) );
  AND2_X1 U11498 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10449), .ZN(P1_U3321) );
  INV_X1 U11499 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10452) );
  NAND2_X1 U11500 ( .A1(n10450), .A2(n10453), .ZN(n10451) );
  OAI21_X1 U11501 ( .B1(n10453), .B2(n10452), .A(n10451), .ZN(P1_U3441) );
  OAI22_X1 U11502 ( .A1(n10457), .A2(n10456), .B1(n10455), .B2(n10454), .ZN(
        n10459) );
  AOI211_X1 U11503 ( .C1(n10461), .C2(n10460), .A(n10459), .B(n10458), .ZN(
        n10464) );
  AOI22_X1 U11504 ( .A1(n10335), .A2(n10464), .B1(n6426), .B2(n10462), .ZN(
        P1_U3463) );
  AOI22_X1 U11505 ( .A1(n10465), .A2(n10464), .B1(n6428), .B2(n10463), .ZN(
        P1_U3526) );
  NOR2_X1 U11506 ( .A1(n10467), .A2(n10466), .ZN(n10474) );
  AND2_X1 U11507 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10477), .ZN(P2_U3297) );
  AND2_X1 U11508 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10477), .ZN(P2_U3298) );
  AND2_X1 U11509 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10477), .ZN(P2_U3299) );
  AND2_X1 U11510 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10477), .ZN(P2_U3300) );
  AND2_X1 U11511 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10477), .ZN(P2_U3301) );
  AND2_X1 U11512 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10477), .ZN(P2_U3302) );
  AND2_X1 U11513 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10477), .ZN(P2_U3303) );
  NOR2_X1 U11514 ( .A1(n10474), .A2(n10468), .ZN(P2_U3304) );
  NOR2_X1 U11515 ( .A1(n10474), .A2(n10469), .ZN(P2_U3305) );
  AND2_X1 U11516 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10477), .ZN(P2_U3306) );
  AND2_X1 U11517 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10477), .ZN(P2_U3307) );
  AND2_X1 U11518 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10477), .ZN(P2_U3308) );
  NOR2_X1 U11519 ( .A1(n10474), .A2(n10470), .ZN(P2_U3309) );
  AND2_X1 U11520 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10477), .ZN(P2_U3310) );
  AND2_X1 U11521 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10477), .ZN(P2_U3311) );
  AND2_X1 U11522 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10477), .ZN(P2_U3312) );
  NOR2_X1 U11523 ( .A1(n10474), .A2(n10471), .ZN(P2_U3313) );
  AND2_X1 U11524 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10477), .ZN(P2_U3314) );
  AND2_X1 U11525 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10477), .ZN(P2_U3315) );
  AND2_X1 U11526 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10477), .ZN(P2_U3316) );
  AND2_X1 U11527 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10477), .ZN(P2_U3317) );
  AND2_X1 U11528 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10477), .ZN(P2_U3318) );
  AND2_X1 U11529 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10477), .ZN(P2_U3319) );
  NOR2_X1 U11530 ( .A1(n10474), .A2(n10472), .ZN(P2_U3320) );
  AND2_X1 U11531 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10477), .ZN(P2_U3321) );
  AND2_X1 U11532 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10477), .ZN(P2_U3322) );
  AND2_X1 U11533 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10477), .ZN(P2_U3323) );
  AND2_X1 U11534 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10477), .ZN(P2_U3324) );
  AND2_X1 U11535 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10477), .ZN(P2_U3325) );
  NOR2_X1 U11536 ( .A1(n10474), .A2(n10473), .ZN(P2_U3326) );
  AOI22_X1 U11537 ( .A1(n10480), .A2(n10476), .B1(n10475), .B2(n10477), .ZN(
        P2_U3437) );
  AOI22_X1 U11538 ( .A1(n10480), .A2(n10479), .B1(n10478), .B2(n10477), .ZN(
        P2_U3438) );
  AOI22_X1 U11539 ( .A1(n10483), .A2(n10510), .B1(n10482), .B2(n10481), .ZN(
        n10484) );
  AND2_X1 U11540 ( .A1(n10485), .A2(n10484), .ZN(n10514) );
  AOI22_X1 U11541 ( .A1(n10513), .A2(n10514), .B1(n5117), .B2(n10512), .ZN(
        P2_U3451) );
  INV_X1 U11542 ( .A(n10486), .ZN(n10487) );
  OAI21_X1 U11543 ( .B1(n10488), .B2(n10507), .A(n10487), .ZN(n10489) );
  AOI211_X1 U11544 ( .C1(n10510), .C2(n10491), .A(n10490), .B(n10489), .ZN(
        n10515) );
  INV_X1 U11545 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10492) );
  AOI22_X1 U11546 ( .A1(n10513), .A2(n10515), .B1(n10492), .B2(n10512), .ZN(
        P2_U3454) );
  INV_X1 U11547 ( .A(n10493), .ZN(n10494) );
  OAI211_X1 U11548 ( .C1(n10496), .C2(n10507), .A(n10495), .B(n10494), .ZN(
        n10497) );
  AOI21_X1 U11549 ( .B1(n10510), .B2(n10498), .A(n10497), .ZN(n10516) );
  INV_X1 U11550 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U11551 ( .A1(n10513), .A2(n10516), .B1(n10499), .B2(n10512), .ZN(
        P2_U3466) );
  OAI21_X1 U11552 ( .B1(n10501), .B2(n10507), .A(n10500), .ZN(n10502) );
  AOI211_X1 U11553 ( .C1(n10504), .C2(n10510), .A(n10503), .B(n10502), .ZN(
        n10518) );
  AOI22_X1 U11554 ( .A1(n10513), .A2(n10518), .B1(n5184), .B2(n10512), .ZN(
        P2_U3469) );
  OAI211_X1 U11555 ( .C1(n10508), .C2(n10507), .A(n10506), .B(n10505), .ZN(
        n10509) );
  AOI21_X1 U11556 ( .B1(n10511), .B2(n10510), .A(n10509), .ZN(n10521) );
  AOI22_X1 U11557 ( .A1(n10513), .A2(n10521), .B1(n5203), .B2(n10512), .ZN(
        P2_U3472) );
  AOI22_X1 U11558 ( .A1(n10522), .A2(n10514), .B1(n6964), .B2(n10519), .ZN(
        P2_U3520) );
  AOI22_X1 U11559 ( .A1(n10522), .A2(n10515), .B1(n6781), .B2(n10519), .ZN(
        P2_U3521) );
  AOI22_X1 U11560 ( .A1(n10522), .A2(n10516), .B1(n5176), .B2(n10519), .ZN(
        P2_U3525) );
  AOI22_X1 U11561 ( .A1(n10522), .A2(n10518), .B1(n10517), .B2(n10519), .ZN(
        P2_U3526) );
  AOI22_X1 U11562 ( .A1(n10522), .A2(n10521), .B1(n10520), .B2(n10519), .ZN(
        P2_U3527) );
  INV_X1 U11563 ( .A(n10523), .ZN(n10524) );
  NAND2_X1 U11564 ( .A1(n10525), .A2(n10524), .ZN(n10526) );
  XOR2_X1 U11565 ( .A(n10527), .B(n10526), .Z(ADD_1071_U5) );
  XOR2_X1 U11566 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11567 ( .B1(n10530), .B2(n10529), .A(n10528), .ZN(ADD_1071_U56) );
  OAI21_X1 U11568 ( .B1(n10533), .B2(n10532), .A(n10531), .ZN(ADD_1071_U57) );
  OAI21_X1 U11569 ( .B1(n10536), .B2(n10535), .A(n10534), .ZN(ADD_1071_U58) );
  OAI21_X1 U11570 ( .B1(n10539), .B2(n10538), .A(n10537), .ZN(ADD_1071_U59) );
  OAI21_X1 U11571 ( .B1(n10542), .B2(n10541), .A(n10540), .ZN(ADD_1071_U60) );
  OAI21_X1 U11572 ( .B1(n10545), .B2(n10544), .A(n10543), .ZN(ADD_1071_U61) );
  AOI21_X1 U11573 ( .B1(n10548), .B2(n10547), .A(n10546), .ZN(ADD_1071_U62) );
  AOI21_X1 U11574 ( .B1(n10551), .B2(n10550), .A(n10549), .ZN(ADD_1071_U63) );
  XOR2_X1 U11575 ( .A(n10552), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11576 ( .A1(n10554), .A2(n10553), .ZN(n10555) );
  XOR2_X1 U11577 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10555), .Z(ADD_1071_U51) );
  OAI21_X1 U11578 ( .B1(n10558), .B2(n10557), .A(n10556), .ZN(n10559) );
  XNOR2_X1 U11579 ( .A(n10559), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11580 ( .B1(n6501), .B2(n10561), .A(n10560), .ZN(ADD_1071_U47) );
  XOR2_X1 U11581 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10562), .Z(ADD_1071_U48) );
  XOR2_X1 U11582 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10563), .Z(ADD_1071_U49) );
  XOR2_X1 U11583 ( .A(n10565), .B(n10564), .Z(ADD_1071_U54) );
  XOR2_X1 U11584 ( .A(n10567), .B(n10566), .Z(ADD_1071_U53) );
  XNOR2_X1 U11585 ( .A(n10569), .B(n10568), .ZN(ADD_1071_U52) );
  NAND2_X1 U4923 ( .A1(n5231), .A2(n5208), .ZN(n5191) );
  NAND2_X1 U8106 ( .A1(n4372), .A2(n9951), .ZN(n8388) );
  INV_X2 U8152 ( .A(n8135), .ZN(n8938) );
  CLKBUF_X1 U4900 ( .A(n8960), .Z(n4371) );
  CLKBUF_X1 U4920 ( .A(n5143), .Z(n4370) );
  CLKBUF_X1 U4928 ( .A(n6425), .Z(n8190) );
  CLKBUF_X1 U4948 ( .A(n5152), .Z(n5689) );
  NAND2_X1 U4949 ( .A1(n5215), .A2(n5234), .ZN(n5216) );
  CLKBUF_X1 U4950 ( .A(n10059), .Z(n4518) );
  CLKBUF_X1 U5454 ( .A(n10011), .Z(n10139) );
endmodule

