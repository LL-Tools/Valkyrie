

module b21_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006;

  INV_X4 U5102 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X4 U5103 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  XNOR2_X1 U5104 ( .A(n6651), .B(P1_IR_REG_26__SCAN_IN), .ZN(n10574) );
  AND2_X4 U5105 ( .A1(n6817), .A2(n6814), .ZN(n7099) );
  INV_X1 U5106 ( .A(n6542), .ZN(n6531) );
  INV_X1 U5107 ( .A(n6310), .ZN(n6214) );
  BUF_X1 U5108 ( .A(n5727), .Z(n6414) );
  INV_X2 U5109 ( .A(n7250), .ZN(n8793) );
  INV_X1 U5110 ( .A(n6948), .ZN(n5052) );
  INV_X1 U5111 ( .A(n8582), .ZN(n7269) );
  INV_X1 U5112 ( .A(n6436), .ZN(n6434) );
  NAND2_X1 U5113 ( .A1(n5662), .A2(n5661), .ZN(n9546) );
  NAND2_X1 U5114 ( .A1(n9063), .A2(n10568), .ZN(n5037) );
  MUX2_X2 U5115 ( .A(n9039), .B(n9038), .S(n9037), .Z(n9046) );
  NAND2_X1 U5116 ( .A1(n8857), .A2(n8859), .ZN(n8992) );
  AND2_X2 U5117 ( .A1(n7169), .A2(n7415), .ZN(n7250) );
  OAI222_X1 U5118 ( .A1(n10575), .A2(n9145), .B1(P1_U3084), .B2(n6753), .C1(
        n9147), .C2(n5044), .ZN(P1_U3325) );
  NAND2_X2 U5119 ( .A1(n6753), .A2(n6751), .ZN(n7113) );
  INV_X1 U5120 ( .A(n6433), .ZN(n7674) );
  NAND3_X2 U5121 ( .A1(n5683), .A2(n5639), .A3(n5682), .ZN(n6433) );
  OR2_X2 U5122 ( .A1(n6434), .A2(n5045), .ZN(n5712) );
  NAND2_X2 U5123 ( .A1(n5731), .A2(n5065), .ZN(n9281) );
  OR2_X2 U5124 ( .A1(n7509), .A2(n7184), .ZN(n7188) );
  INV_X2 U5125 ( .A(n6947), .ZN(n5038) );
  INV_X2 U5126 ( .A(n6947), .ZN(n5039) );
  NAND4_X1 U5127 ( .A1(n7159), .A2(n7160), .A3(n7158), .A4(n7161), .ZN(n9829)
         );
  OAI22_X2 U5128 ( .A1(n6234), .A2(n6233), .B1(n6232), .B2(n6231), .ZN(n6240)
         );
  XNOR2_X2 U5129 ( .A(n6210), .B(n6209), .ZN(n8599) );
  OAI21_X2 U5130 ( .B1(n8499), .B2(n5526), .A(n5524), .ZN(n8530) );
  NAND2_X2 U5131 ( .A1(n8275), .A2(n8274), .ZN(n8499) );
  AOI21_X2 U5132 ( .B1(n9484), .B2(n6609), .A(n6608), .ZN(n9467) );
  AOI21_X2 U5133 ( .B1(n9490), .B2(n6606), .A(n6605), .ZN(n9484) );
  OR2_X1 U5134 ( .A1(n9370), .A2(n5444), .ZN(n5443) );
  NOR2_X1 U5135 ( .A1(n9083), .A2(n9376), .ZN(n9364) );
  NAND2_X2 U5136 ( .A1(n8530), .A2(n8529), .ZN(n8533) );
  OR2_X1 U5137 ( .A1(n8302), .A2(n8511), .ZN(n8391) );
  OAI21_X1 U5138 ( .B1(n7713), .B2(n7714), .A(n6574), .ZN(n7670) );
  NAND2_X1 U5139 ( .A1(n6441), .A2(n6440), .ZN(n7713) );
  INV_X2 U5140 ( .A(n6628), .ZN(n9101) );
  NAND2_X1 U5141 ( .A1(n5666), .A2(n7147), .ZN(n5047) );
  CLKBUF_X2 U5142 ( .A(n7250), .Z(n8724) );
  INV_X4 U5144 ( .A(n7961), .ZN(n5040) );
  AND2_X1 U5145 ( .A1(n6957), .A2(n8061), .ZN(n7111) );
  INV_X2 U5146 ( .A(n7012), .ZN(n5041) );
  OR2_X2 U5147 ( .A1(n5657), .A2(n5651), .ZN(n6076) );
  NAND2_X1 U5148 ( .A1(n5479), .A2(n5478), .ZN(n9163) );
  OR3_X1 U5149 ( .A1(n10098), .A2(n10097), .A3(n10096), .ZN(n10552) );
  AOI21_X1 U5150 ( .B1(n5342), .B2(n10980), .A(n5339), .ZN(n10091) );
  NAND2_X1 U5151 ( .A1(n5185), .A2(n6616), .ZN(n9371) );
  OAI22_X1 U5152 ( .A1(n9898), .A2(n9904), .B1(n9915), .B2(n10088), .ZN(n9118)
         );
  NAND2_X1 U5153 ( .A1(n9190), .A2(n9189), .ZN(n5477) );
  NAND2_X1 U5154 ( .A1(n5229), .A2(n8534), .ZN(n5512) );
  AND2_X1 U5155 ( .A1(n8544), .A2(n5071), .ZN(n5229) );
  INV_X1 U5156 ( .A(n9447), .ZN(n9443) );
  OAI21_X1 U5157 ( .B1(n8499), .B2(n5533), .A(n5531), .ZN(n8529) );
  AND2_X1 U5158 ( .A1(n5183), .A2(n5182), .ZN(n9508) );
  INV_X1 U5159 ( .A(n9983), .ZN(n10114) );
  NAND2_X1 U5160 ( .A1(n5396), .A2(n9121), .ZN(n10038) );
  AND2_X1 U5161 ( .A1(n8681), .A2(n8680), .ZN(n9983) );
  NAND2_X1 U5162 ( .A1(n5280), .A2(n5278), .ZN(n8460) );
  AOI21_X1 U5163 ( .B1(n5464), .B2(n5463), .A(n5462), .ZN(n6602) );
  NAND2_X1 U5164 ( .A1(n10973), .A2(n10974), .ZN(n10972) );
  NAND2_X1 U5165 ( .A1(n8665), .A2(n8664), .ZN(n10120) );
  AND2_X1 U5166 ( .A1(n7966), .A2(n7967), .ZN(n5208) );
  NAND2_X1 U5167 ( .A1(n5994), .A2(n5993), .ZN(n9664) );
  NAND2_X1 U5168 ( .A1(n7515), .A2(n8999), .ZN(n7856) );
  NAND2_X1 U5169 ( .A1(n5985), .A2(n5984), .ZN(n6009) );
  INV_X2 U5170 ( .A(n10803), .ZN(n7664) );
  INV_X2 U5171 ( .A(n9220), .ZN(n5042) );
  NAND2_X2 U5172 ( .A1(n10808), .A2(n9279), .ZN(n6578) );
  NOR2_X1 U5173 ( .A1(n7326), .A2(n7199), .ZN(n7497) );
  AND2_X1 U5174 ( .A1(n5766), .A2(n5765), .ZN(n10775) );
  OAI211_X2 U5175 ( .C1(n7510), .C2(n9850), .A(n7188), .B(n7187), .ZN(n7199)
         );
  INV_X4 U5176 ( .A(n7104), .ZN(n7961) );
  AND2_X2 U5177 ( .A1(n8795), .A2(n5508), .ZN(n8790) );
  NAND4_X1 U5178 ( .A1(n7134), .A2(n7133), .A3(n7132), .A4(n7131), .ZN(n9827)
         );
  OAI211_X1 U5179 ( .C1(n7012), .C2(n7056), .A(n5749), .B(n5748), .ZN(n7681)
         );
  INV_X1 U5180 ( .A(n7111), .ZN(n7415) );
  NAND2_X1 U5181 ( .A1(n6652), .A2(n10574), .ZN(n7208) );
  INV_X2 U5182 ( .A(n6948), .ZN(n7351) );
  INV_X4 U5183 ( .A(n5037), .ZN(n5051) );
  CLKBUF_X3 U5184 ( .A(n5767), .Z(n6403) );
  CLKBUF_X1 U5185 ( .A(n6355), .Z(n6635) );
  NAND2_X1 U5186 ( .A1(n5703), .A2(n5680), .ZN(n5762) );
  AND2_X1 U5187 ( .A1(n9694), .A2(n9062), .ZN(n5768) );
  NAND2_X1 U5188 ( .A1(n6650), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6651) );
  INV_X1 U5189 ( .A(n9063), .ZN(n6817) );
  NAND2_X1 U5191 ( .A1(n6365), .A2(n6634), .ZN(n5703) );
  NAND2_X1 U5192 ( .A1(n5688), .A2(n5691), .ZN(n9062) );
  NAND2_X1 U5193 ( .A1(n6813), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6808) );
  NAND2_X1 U5194 ( .A1(n5688), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5687) );
  XNOR2_X1 U5195 ( .A(n6931), .B(n6653), .ZN(n9958) );
  INV_X2 U5196 ( .A(n8353), .ZN(n5043) );
  INV_X2 U5197 ( .A(n8350), .ZN(n5044) );
  AND2_X1 U5198 ( .A1(n5053), .A2(n5282), .ZN(n5281) );
  CLKBUF_X3 U5199 ( .A(n5720), .Z(n6789) );
  NAND2_X1 U5200 ( .A1(n6654), .A2(n5285), .ZN(n6646) );
  NOR2_X1 U5201 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(n5490), .ZN(n5440) );
  AND3_X1 U5202 ( .A1(n6928), .A2(n6672), .A3(n6645), .ZN(n6654) );
  AND2_X1 U5203 ( .A1(n6656), .A2(n6653), .ZN(n5285) );
  AND4_X1 U5204 ( .A1(n6686), .A2(n10318), .A3(n10319), .A4(n10325), .ZN(n5053) );
  NAND3_X1 U5205 ( .A1(n5337), .A2(n5338), .A3(n5336), .ZN(n5249) );
  NAND3_X1 U5206 ( .A1(n5407), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5248) );
  AND4_X1 U5207 ( .A1(n6642), .A2(n6718), .A3(n6691), .A4(n10301), .ZN(n6644)
         );
  AND3_X1 U5208 ( .A1(n6641), .A2(n6640), .A3(n6639), .ZN(n6693) );
  INV_X1 U5209 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6327) );
  NOR2_X1 U5210 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n6640) );
  INV_X1 U5211 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5337) );
  INV_X1 U5212 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n10325) );
  INV_X1 U5213 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n10318) );
  INV_X1 U5214 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n10319) );
  INV_X1 U5215 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6686) );
  NOR2_X1 U5216 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n6642) );
  INV_X1 U5217 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n10301) );
  NOR2_X1 U5218 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n6641) );
  NOR2_X1 U5219 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n6639) );
  INV_X1 U5220 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6718) );
  NOR2_X1 U5221 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6724) );
  INV_X1 U5222 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n6807) );
  INV_X1 U5223 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6691) );
  INV_X1 U5224 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5407) );
  INV_X1 U5225 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5336) );
  INV_X1 U5226 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5338) );
  INV_X1 U5227 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5948) );
  NOR2_X1 U5228 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5643) );
  INV_X1 U5229 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5990) );
  NOR2_X1 U5230 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5647) );
  NOR2_X1 U5231 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5648) );
  AND2_X1 U5232 ( .A1(n5699), .A2(n5698), .ZN(n5045) );
  OAI21_X2 U5233 ( .B1(n9508), .B2(n9507), .A(n5181), .ZN(n9490) );
  OAI21_X2 U5234 ( .B1(n9735), .B2(n5253), .A(n5252), .ZN(n5545) );
  NAND2_X1 U5235 ( .A1(n5666), .A2(n7147), .ZN(n5046) );
  NAND4_X2 U5236 ( .A1(n7103), .A2(n7102), .A3(n7101), .A4(n7100), .ZN(n9828)
         );
  XNOR2_X1 U5237 ( .A(n5713), .B(n5712), .ZN(n9179) );
  INV_X1 U5238 ( .A(n6751), .ZN(n5049) );
  INV_X1 U5239 ( .A(n5049), .ZN(n5050) );
  XNOR2_X2 U5240 ( .A(n6812), .B(P1_IR_REG_28__SCAN_IN), .ZN(n6753) );
  INV_X1 U5241 ( .A(n7199), .ZN(n7441) );
  NAND2_X1 U5242 ( .A1(n7493), .A2(n7199), .ZN(n8857) );
  INV_X1 U5243 ( .A(n7272), .ZN(n7274) );
  OR2_X1 U5244 ( .A1(n7275), .A2(n7272), .ZN(n7326) );
  OAI211_X2 U5245 ( .C1(n7510), .C2(n7109), .A(n7108), .B(n7107), .ZN(n7272)
         );
  AND2_X1 U5246 ( .A1(n6418), .A2(n6539), .ZN(n6626) );
  AND2_X1 U5247 ( .A1(n5109), .A2(n5192), .ZN(n5191) );
  NAND2_X1 U5248 ( .A1(n9443), .A2(n6611), .ZN(n5192) );
  OR2_X1 U5249 ( .A1(n9612), .A2(n9197), .ZN(n6612) );
  AOI21_X1 U5250 ( .B1(n5567), .B2(n5565), .A(n5094), .ZN(n5564) );
  INV_X1 U5251 ( .A(n5067), .ZN(n5565) );
  NOR2_X1 U5252 ( .A1(n9002), .A2(n5577), .ZN(n5576) );
  INV_X1 U5253 ( .A(n7855), .ZN(n5577) );
  NOR2_X1 U5254 ( .A1(n5938), .A2(n5412), .ZN(n5411) );
  INV_X1 U5255 ( .A(n5935), .ZN(n5938) );
  INV_X1 U5256 ( .A(n5916), .ZN(n5412) );
  CLKBUF_X1 U5257 ( .A(n5737), .Z(n6217) );
  INV_X1 U5258 ( .A(n5605), .ZN(n5604) );
  OAI21_X1 U5259 ( .B1(n9082), .B2(n5609), .A(n9081), .ZN(n5605) );
  OR2_X1 U5260 ( .A1(n9592), .A2(n9393), .ZN(n9081) );
  OR2_X1 U5261 ( .A1(n9482), .A2(n9266), .ZN(n5640) );
  OR2_X1 U5262 ( .A1(n8511), .A2(n8390), .ZN(n8922) );
  XNOR2_X1 U5263 ( .A(n6400), .B(n6399), .ZN(n9687) );
  INV_X1 U5264 ( .A(n9076), .ZN(n5616) );
  OR2_X1 U5265 ( .A1(n9629), .A2(n9266), .ZN(n6609) );
  OR2_X1 U5266 ( .A1(n9651), .A2(n9066), .ZN(n6603) );
  INV_X1 U5267 ( .A(n8424), .ZN(n5626) );
  OR2_X1 U5268 ( .A1(n9655), .A2(n9540), .ZN(n6600) );
  OR2_X1 U5269 ( .A1(n5955), .A2(n7790), .ZN(n5975) );
  NAND2_X1 U5270 ( .A1(n6445), .A2(n7681), .ZN(n6575) );
  XNOR2_X1 U5271 ( .A(n10790), .B(n10775), .ZN(n7750) );
  INV_X1 U5272 ( .A(n5491), .ZN(n5439) );
  NOR2_X1 U5273 ( .A1(n9809), .A2(n5242), .ZN(n5241) );
  INV_X1 U5274 ( .A(n8721), .ZN(n5242) );
  OR2_X1 U5275 ( .A1(n8231), .A2(n8295), .ZN(n8820) );
  NAND2_X1 U5276 ( .A1(n5267), .A2(n5265), .ZN(n8133) );
  NAND2_X1 U5277 ( .A1(n5433), .A2(n5432), .ZN(n6420) );
  AOI21_X1 U5278 ( .B1(n5434), .B2(n5436), .A(n5123), .ZN(n5432) );
  INV_X1 U5279 ( .A(n6646), .ZN(n5283) );
  NAND2_X1 U5280 ( .A1(n5415), .A2(n5413), .ZN(n6234) );
  AOI21_X1 U5281 ( .B1(n5416), .B2(n5418), .A(n5414), .ZN(n5413) );
  NAND2_X1 U5282 ( .A1(n5231), .A2(n5230), .ZN(n5415) );
  INV_X1 U5283 ( .A(n6211), .ZN(n5414) );
  OAI21_X1 U5284 ( .B1(n6094), .B2(n5428), .A(n5425), .ZN(n6126) );
  AOI21_X1 U5285 ( .B1(n6092), .B2(n5427), .A(n5426), .ZN(n5425) );
  INV_X1 U5286 ( .A(n6119), .ZN(n5426) );
  AND2_X1 U5287 ( .A1(n5409), .A2(n5937), .ZN(n5408) );
  INV_X1 U5288 ( .A(n5944), .ZN(n5409) );
  OAI21_X1 U5289 ( .B1(n5335), .B2(n5778), .A(n5801), .ZN(n5332) );
  INV_X1 U5290 ( .A(n5781), .ZN(n5335) );
  INV_X1 U5291 ( .A(n5883), .ZN(n5882) );
  NAND2_X1 U5292 ( .A1(n9241), .A2(n5962), .ZN(n8561) );
  INV_X1 U5293 ( .A(n5424), .ZN(n5423) );
  OAI21_X1 U5294 ( .B1(n6572), .B2(n5697), .A(n8174), .ZN(n5424) );
  AND2_X1 U5295 ( .A1(n6223), .A2(n6222), .ZN(n9197) );
  INV_X1 U5296 ( .A(n6414), .ZN(n6360) );
  AND2_X1 U5297 ( .A1(n6635), .A2(n6435), .ZN(n6855) );
  AND2_X1 U5298 ( .A1(n5187), .A2(n5143), .ZN(n5184) );
  OAI21_X1 U5299 ( .B1(n9398), .B2(n9401), .A(n5162), .ZN(n9384) );
  INV_X1 U5300 ( .A(n5164), .ZN(n5162) );
  AOI21_X1 U5301 ( .B1(n9412), .B2(n9420), .A(n9079), .ZN(n9398) );
  NOR2_X1 U5302 ( .A1(n9608), .A2(n9078), .ZN(n9079) );
  AND2_X1 U5303 ( .A1(n9618), .A2(n9468), .ZN(n9076) );
  NAND2_X1 U5304 ( .A1(n6612), .A2(n6550), .ZN(n9435) );
  NAND2_X1 U5305 ( .A1(n5171), .A2(n5059), .ZN(n9458) );
  NAND2_X1 U5306 ( .A1(n9496), .A2(n5172), .ZN(n5171) );
  NAND2_X1 U5307 ( .A1(n5172), .A2(n5174), .ZN(n5170) );
  OAI21_X1 U5308 ( .B1(n9496), .B2(n5174), .A(n5172), .ZN(n9474) );
  NOR2_X1 U5309 ( .A1(n9664), .A2(n10938), .ZN(n5305) );
  NAND2_X1 U5310 ( .A1(n6317), .A2(n6316), .ZN(n9592) );
  INV_X1 U5311 ( .A(n6055), .ZN(n5197) );
  INV_X1 U5312 ( .A(n5527), .ZN(n5526) );
  AOI21_X1 U5313 ( .B1(n5527), .B2(n5076), .A(n5525), .ZN(n5524) );
  NOR2_X1 U5314 ( .A1(n8516), .A2(n5528), .ZN(n5527) );
  NOR2_X1 U5315 ( .A1(n9933), .A2(n5319), .ZN(n9892) );
  NAND2_X1 U5316 ( .A1(n5321), .A2(n5320), .ZN(n5319) );
  NOR2_X1 U5317 ( .A1(n10078), .A2(n9922), .ZN(n5320) );
  NOR2_X1 U5318 ( .A1(n9118), .A2(n9130), .ZN(n9149) );
  NOR2_X1 U5319 ( .A1(n9933), .A2(n9922), .ZN(n9924) );
  NAND2_X1 U5320 ( .A1(n5260), .A2(n5562), .ZN(n9898) );
  AOI21_X1 U5321 ( .B1(n5564), .B2(n5566), .A(n5095), .ZN(n5562) );
  NAND2_X1 U5322 ( .A1(n9947), .A2(n5564), .ZN(n5260) );
  OR2_X1 U5323 ( .A1(n10105), .A2(n9971), .ZN(n9116) );
  OAI21_X1 U5324 ( .B1(n9110), .B2(n5276), .A(n5274), .ZN(n9976) );
  INV_X1 U5325 ( .A(n5275), .ZN(n5274) );
  OAI21_X1 U5326 ( .B1(n5068), .B2(n5276), .A(n9977), .ZN(n5275) );
  INV_X1 U5327 ( .A(n9111), .ZN(n5276) );
  OAI21_X1 U5328 ( .B1(n8254), .B2(n5324), .A(n5322), .ZN(n10973) );
  AOI21_X1 U5329 ( .B1(n9007), .B2(n5325), .A(n5323), .ZN(n5322) );
  INV_X1 U5330 ( .A(n5325), .ZN(n5324) );
  INV_X1 U5331 ( .A(n8925), .ZN(n5323) );
  AOI21_X1 U5332 ( .B1(n9007), .B2(n5571), .A(n5090), .ZN(n5570) );
  INV_X1 U5333 ( .A(n8241), .ZN(n5571) );
  INV_X1 U5334 ( .A(n7510), .ZN(n8637) );
  NAND2_X1 U5336 ( .A1(n9118), .A2(n9130), .ZN(n5590) );
  NAND2_X1 U5337 ( .A1(n6402), .A2(n6401), .ZN(n9580) );
  XNOR2_X1 U5338 ( .A(n10073), .B(n10072), .ZN(n10071) );
  INV_X1 U5339 ( .A(n9149), .ZN(n5591) );
  INV_X1 U5340 ( .A(n10733), .ZN(n10068) );
  OAI21_X1 U5341 ( .B1(n10159), .B2(n5381), .A(n10160), .ZN(n5380) );
  XNOR2_X1 U5342 ( .A(keyinput_134), .B(SI_26_), .ZN(n5381) );
  XNOR2_X1 U5343 ( .A(n10161), .B(n5379), .ZN(n5378) );
  INV_X1 U5344 ( .A(keyinput_137), .ZN(n5379) );
  AOI21_X1 U5345 ( .B1(n10190), .B2(n10191), .A(n5386), .ZN(n5385) );
  XNOR2_X1 U5346 ( .A(SI_5_), .B(keyinput_155), .ZN(n5386) );
  NAND2_X1 U5347 ( .A1(n10200), .A2(n10201), .ZN(n5383) );
  OR2_X1 U5348 ( .A1(n10208), .A2(n5353), .ZN(n5352) );
  NAND2_X1 U5349 ( .A1(n10209), .A2(n5354), .ZN(n5353) );
  NAND2_X1 U5350 ( .A1(keyinput_170), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5354)
         );
  NOR2_X1 U5351 ( .A1(n10217), .A2(n5351), .ZN(n5350) );
  XNOR2_X1 U5352 ( .A(n10210), .B(keyinput_172), .ZN(n5351) );
  AOI21_X1 U5353 ( .B1(n10224), .B2(n10223), .A(n5347), .ZN(n5346) );
  OAI22_X1 U5354 ( .A1(n10225), .A2(keyinput_182), .B1(n10226), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n5347) );
  INV_X1 U5355 ( .A(n5345), .ZN(n5344) );
  OAI22_X1 U5356 ( .A1(n10231), .A2(n10230), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(keyinput_184), .ZN(n5345) );
  NOR2_X1 U5357 ( .A1(n5975), .A2(n10231), .ZN(n5137) );
  NAND2_X1 U5358 ( .A1(n6438), .A2(n5597), .ZN(n6441) );
  NAND2_X1 U5359 ( .A1(n7313), .A2(n7272), .ZN(n8852) );
  AND2_X1 U5360 ( .A1(n6159), .A2(n6142), .ZN(n5232) );
  INV_X1 U5361 ( .A(n6117), .ZN(n5429) );
  NAND2_X1 U5362 ( .A1(n5872), .A2(n10186), .ZN(n5895) );
  AOI21_X1 U5363 ( .B1(n8557), .B2(n5474), .A(n5074), .ZN(n5473) );
  INV_X1 U5364 ( .A(n5965), .ZN(n5474) );
  INV_X1 U5365 ( .A(n6617), .ZN(n5442) );
  AOI21_X1 U5366 ( .B1(n6547), .B2(n6546), .A(n6545), .ZN(n6572) );
  OR2_X1 U5367 ( .A1(n9083), .A2(n9374), .ZN(n6618) );
  OR2_X1 U5368 ( .A1(n9597), .A2(n9375), .ZN(n6616) );
  NOR2_X1 U5369 ( .A1(n6244), .A2(n10213), .ZN(n5142) );
  OR2_X1 U5370 ( .A1(n9612), .A2(n9445), .ZN(n9077) );
  OR2_X1 U5371 ( .A1(n9618), .A2(n9436), .ZN(n6551) );
  INV_X1 U5372 ( .A(n9071), .ZN(n5174) );
  AND2_X1 U5373 ( .A1(n9475), .A2(n5173), .ZN(n5172) );
  NAND2_X1 U5374 ( .A1(n6606), .A2(n9071), .ZN(n5173) );
  INV_X1 U5375 ( .A(n5628), .ZN(n5625) );
  AND2_X1 U5376 ( .A1(n5305), .A2(n5304), .ZN(n5303) );
  INV_X1 U5377 ( .A(n5137), .ZN(n5996) );
  NOR2_X1 U5378 ( .A1(n7943), .A2(n7813), .ZN(n5302) );
  INV_X1 U5379 ( .A(n6579), .ZN(n5454) );
  NOR2_X1 U5380 ( .A1(n6580), .A2(n5452), .ZN(n5455) );
  INV_X1 U5381 ( .A(n6577), .ZN(n5452) );
  NOR2_X1 U5382 ( .A1(n9641), .A2(n9519), .ZN(n9511) );
  NOR2_X1 U5383 ( .A1(n6055), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n5657) );
  OR2_X1 U5384 ( .A1(n10083), .A2(n8841), .ZN(n9155) );
  OR2_X1 U5385 ( .A1(n9922), .A2(n9738), .ZN(n8879) );
  NAND2_X1 U5386 ( .A1(n9913), .A2(n9914), .ZN(n9912) );
  NOR2_X1 U5387 ( .A1(n10114), .A2(n5315), .ZN(n5314) );
  INV_X1 U5388 ( .A(n5316), .ZN(n5315) );
  OR2_X1 U5389 ( .A1(n8554), .A2(n8496), .ZN(n8926) );
  NAND2_X1 U5390 ( .A1(n8233), .A2(n8232), .ZN(n8292) );
  AND2_X1 U5391 ( .A1(n10891), .A2(n5062), .ZN(n5309) );
  INV_X1 U5392 ( .A(n7938), .ZN(n5311) );
  AND2_X1 U5393 ( .A1(n8013), .A2(n5272), .ZN(n5271) );
  NAND2_X1 U5394 ( .A1(n5070), .A2(n5273), .ZN(n5272) );
  AND2_X1 U5395 ( .A1(n5102), .A2(n8882), .ZN(n8862) );
  NAND2_X1 U5396 ( .A1(n7489), .A2(n8860), .ZN(n7527) );
  NAND2_X1 U5397 ( .A1(n5100), .A2(n5256), .ZN(n9158) );
  NAND2_X1 U5398 ( .A1(n5393), .A2(n5392), .ZN(n5391) );
  AOI21_X1 U5399 ( .B1(n5357), .B2(n5359), .A(n5132), .ZN(n5356) );
  AOI21_X1 U5400 ( .B1(n5237), .B2(n5235), .A(n5234), .ZN(n5233) );
  INV_X1 U5401 ( .A(n5237), .ZN(n5236) );
  INV_X1 U5402 ( .A(n6278), .ZN(n5234) );
  NAND2_X1 U5403 ( .A1(n5240), .A2(n5239), .ZN(n6257) );
  INV_X1 U5404 ( .A(n6239), .ZN(n5239) );
  INV_X1 U5405 ( .A(n6240), .ZN(n5240) );
  OAI21_X1 U5406 ( .B1(n6075), .B2(n6074), .A(n6073), .ZN(n6094) );
  NAND2_X1 U5407 ( .A1(n5211), .A2(n5209), .ZN(n6075) );
  AOI21_X1 U5408 ( .B1(n5213), .B2(n5216), .A(n5210), .ZN(n5209) );
  NAND2_X1 U5409 ( .A1(n6009), .A2(n5213), .ZN(n5211) );
  INV_X1 U5410 ( .A(n6053), .ZN(n5210) );
  OR2_X1 U5411 ( .A1(n6708), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6710) );
  NAND2_X1 U5412 ( .A1(n5848), .A2(n5847), .ZN(n5870) );
  NAND2_X1 U5413 ( .A1(n5868), .A2(n5852), .ZN(n5869) );
  AND2_X1 U5414 ( .A1(n5758), .A2(n5781), .ZN(n5333) );
  OAI21_X1 U5415 ( .B1(n6789), .B2(n5761), .A(n5760), .ZN(n5780) );
  NAND2_X1 U5416 ( .A1(n6789), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5760) );
  AND2_X1 U5417 ( .A1(n9254), .A2(n5482), .ZN(n5481) );
  OR2_X1 U5418 ( .A1(n9195), .A2(n5483), .ZN(n5482) );
  INV_X1 U5419 ( .A(n6255), .ZN(n5483) );
  INV_X1 U5420 ( .A(n9098), .ZN(n7148) );
  INV_X1 U5421 ( .A(n5768), .ZN(n6109) );
  INV_X1 U5422 ( .A(n5925), .ZN(n5924) );
  OR2_X1 U5423 ( .A1(n5904), .A2(n10140), .ZN(n5925) );
  NAND2_X1 U5424 ( .A1(n5489), .A2(n5487), .ZN(n9241) );
  AND2_X1 U5425 ( .A1(n9235), .A2(n5488), .ZN(n5487) );
  NAND2_X1 U5426 ( .A1(n7845), .A2(n5914), .ZN(n5488) );
  AND2_X1 U5427 ( .A1(n6068), .A2(n6049), .ZN(n5485) );
  NAND2_X1 U5428 ( .A1(n8371), .A2(n8174), .ZN(n6573) );
  XNOR2_X1 U5429 ( .A(n6572), .B(n5421), .ZN(n5420) );
  INV_X1 U5430 ( .A(n7146), .ZN(n5421) );
  NOR4_X1 U5431 ( .A1(n6569), .A2(n6568), .A3(n9372), .A4(n6567), .ZN(n6570)
         );
  AND4_X1 U5432 ( .A1(n5862), .A2(n5861), .A3(n5860), .A4(n5859), .ZN(n7603)
         );
  NAND2_X1 U5433 ( .A1(n5768), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5730) );
  NAND2_X1 U5434 ( .A1(n8052), .A2(n8053), .ZN(n8198) );
  NAND2_X1 U5435 ( .A1(n8201), .A2(n8200), .ZN(n9296) );
  OR2_X1 U5436 ( .A1(n9300), .A2(n9299), .ZN(n5157) );
  AOI21_X1 U5437 ( .B1(n5191), .B2(n5188), .A(n5099), .ZN(n5187) );
  INV_X1 U5438 ( .A(n6611), .ZN(n5188) );
  OR2_X1 U5439 ( .A1(n5458), .A2(n6615), .ZN(n5457) );
  INV_X1 U5440 ( .A(n5191), .ZN(n5189) );
  OR2_X1 U5441 ( .A1(n9608), .A2(n9437), .ZN(n9399) );
  INV_X1 U5442 ( .A(n5142), .ZN(n6265) );
  NAND2_X1 U5443 ( .A1(n9399), .A2(n6521), .ZN(n9420) );
  NAND2_X1 U5444 ( .A1(n5190), .A2(n6611), .ZN(n9434) );
  OR2_X1 U5445 ( .A1(n9444), .A2(n9443), .ZN(n5190) );
  NOR2_X1 U5446 ( .A1(n9434), .A2(n9435), .ZN(n9433) );
  XNOR2_X1 U5447 ( .A(n9624), .B(n9485), .ZN(n9466) );
  OR2_X1 U5448 ( .A1(n9629), .A2(n9498), .ZN(n9477) );
  OR2_X1 U5449 ( .A1(n9069), .A2(n9068), .ZN(n5634) );
  NAND2_X1 U5450 ( .A1(n9496), .A2(n9495), .ZN(n9494) );
  OR2_X1 U5451 ( .A1(n9641), .A2(n9068), .ZN(n5181) );
  NAND2_X1 U5452 ( .A1(n6102), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6131) );
  INV_X1 U5453 ( .A(n6104), .ZN(n6102) );
  OR2_X1 U5454 ( .A1(n6040), .A2(n6039), .ZN(n6059) );
  INV_X1 U5455 ( .A(n5136), .ZN(n6079) );
  NOR2_X1 U5456 ( .A1(n5468), .A2(n6595), .ZN(n5463) );
  NAND2_X1 U5457 ( .A1(n5627), .A2(n5626), .ZN(n5623) );
  INV_X1 U5458 ( .A(n5623), .ZN(n9065) );
  OR2_X1 U5459 ( .A1(n9659), .A2(n8422), .ZN(n8416) );
  AOI21_X1 U5460 ( .B1(n8421), .B2(n9052), .A(n8420), .ZN(n8441) );
  NAND2_X1 U5461 ( .A1(n8357), .A2(n5081), .ZN(n8359) );
  AOI21_X1 U5462 ( .B1(n8073), .B2(n8081), .A(n6593), .ZN(n8092) );
  AND2_X1 U5463 ( .A1(n8039), .A2(n8038), .ZN(n8083) );
  AND2_X1 U5464 ( .A1(n8083), .A2(n10920), .ZN(n8101) );
  AND2_X1 U5465 ( .A1(n5302), .A2(n5301), .ZN(n5300) );
  AND3_X1 U5466 ( .A1(n5300), .A2(n5299), .A3(n9565), .ZN(n8039) );
  NOR2_X1 U5467 ( .A1(n7948), .A2(n5619), .ZN(n5618) );
  INV_X1 U5468 ( .A(n7944), .ZN(n5619) );
  NAND2_X1 U5469 ( .A1(n9569), .A2(n5629), .ZN(n7808) );
  AND2_X1 U5470 ( .A1(n7809), .A2(n7777), .ZN(n5629) );
  AND2_X1 U5471 ( .A1(n6467), .A2(n6583), .ZN(n7807) );
  AND4_X1 U5472 ( .A1(n5836), .A2(n5835), .A3(n5834), .A4(n5833), .ZN(n9560)
         );
  NAND2_X1 U5473 ( .A1(n5455), .A2(n7742), .ZN(n5453) );
  NOR2_X1 U5474 ( .A1(n10783), .A2(n10795), .ZN(n10786) );
  NAND2_X1 U5475 ( .A1(n6578), .A2(n6579), .ZN(n10787) );
  NAND2_X1 U5476 ( .A1(n7669), .A2(n7748), .ZN(n5178) );
  AND4_X1 U5477 ( .A1(n5796), .A2(n5795), .A3(n5794), .A4(n5793), .ZN(n9562)
         );
  OR2_X1 U5478 ( .A1(n7141), .A2(n6367), .ZN(n9559) );
  OR2_X1 U5479 ( .A1(n7141), .A2(n6366), .ZN(n9561) );
  AOI21_X1 U5480 ( .B1(n7670), .B2(n7669), .A(n6576), .ZN(n7744) );
  INV_X1 U5481 ( .A(n9561), .ZN(n10789) );
  NAND2_X1 U5482 ( .A1(n7680), .A2(n7679), .ZN(n7749) );
  XNOR2_X1 U5483 ( .A(n10752), .B(n9281), .ZN(n7714) );
  INV_X1 U5484 ( .A(n5292), .ZN(n5289) );
  AND2_X1 U5485 ( .A1(n6354), .A2(n5698), .ZN(n10939) );
  NOR2_X1 U5486 ( .A1(n5673), .A2(n5054), .ZN(n5196) );
  NAND2_X1 U5487 ( .A1(n5661), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U5488 ( .A1(n7692), .A2(n7693), .ZN(n7834) );
  NAND2_X1 U5489 ( .A1(n5530), .A2(n5529), .ZN(n8517) );
  XNOR2_X1 U5490 ( .A(n7191), .B(n8793), .ZN(n7238) );
  INV_X1 U5491 ( .A(n5519), .ZN(n5518) );
  OAI21_X1 U5492 ( .B1(n5522), .B2(n7693), .A(n7830), .ZN(n5519) );
  NOR2_X1 U5493 ( .A1(n9763), .A2(n5560), .ZN(n5559) );
  INV_X1 U5494 ( .A(n5561), .ZN(n5560) );
  NOR2_X1 U5495 ( .A1(n8687), .A2(n8686), .ZN(n9702) );
  NAND2_X1 U5496 ( .A1(n9831), .A2(n8790), .ZN(n6960) );
  NAND2_X1 U5497 ( .A1(n5556), .A2(n9764), .ZN(n5555) );
  INV_X1 U5498 ( .A(n5559), .ZN(n5556) );
  NOR2_X1 U5499 ( .A1(n5557), .A2(n5551), .ZN(n5550) );
  INV_X1 U5500 ( .A(n9714), .ZN(n5551) );
  NAND2_X1 U5501 ( .A1(n5558), .A2(n9764), .ZN(n5557) );
  INV_X1 U5502 ( .A(n9723), .ZN(n5558) );
  XNOR2_X1 U5503 ( .A(n8793), .B(n5250), .ZN(n7194) );
  OAI21_X1 U5504 ( .B1(n7961), .B2(n7313), .A(n7110), .ZN(n5250) );
  NAND2_X1 U5505 ( .A1(n5228), .A2(n5226), .ZN(n5225) );
  NAND2_X1 U5506 ( .A1(n5228), .A2(n8546), .ZN(n5227) );
  NOR2_X1 U5507 ( .A1(n5504), .A2(n5503), .ZN(n5502) );
  NAND2_X1 U5508 ( .A1(n5504), .A2(n5503), .ZN(n5222) );
  NAND2_X1 U5509 ( .A1(n7207), .A2(n5509), .ZN(n5508) );
  NAND2_X1 U5510 ( .A1(n7351), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6949) );
  NAND2_X1 U5511 ( .A1(n8746), .A2(n8745), .ZN(n9893) );
  INV_X1 U5512 ( .A(n5321), .ZN(n5318) );
  NAND2_X1 U5513 ( .A1(n9912), .A2(n9903), .ZN(n5343) );
  NAND2_X1 U5514 ( .A1(n9905), .A2(n10977), .ZN(n5341) );
  AND2_X1 U5515 ( .A1(n8963), .A2(n9129), .ZN(n9904) );
  NAND2_X1 U5516 ( .A1(n5101), .A2(n5055), .ZN(n5567) );
  NAND2_X1 U5517 ( .A1(n5069), .A2(n9116), .ZN(n5568) );
  AND2_X1 U5518 ( .A1(n8879), .A2(n9903), .ZN(n9914) );
  INV_X1 U5519 ( .A(n9117), .ZN(n9941) );
  NAND2_X1 U5520 ( .A1(n9115), .A2(n9114), .ZN(n9947) );
  INV_X1 U5521 ( .A(n10003), .ZN(n5277) );
  AND2_X1 U5522 ( .A1(n8940), .A2(n9124), .ZN(n10003) );
  NOR2_X1 U5523 ( .A1(n5092), .A2(n5574), .ZN(n5573) );
  INV_X1 U5524 ( .A(n9108), .ZN(n5574) );
  NOR2_X1 U5525 ( .A1(n10031), .A2(n5397), .ZN(n5396) );
  OR2_X1 U5526 ( .A1(n10541), .A2(n9793), .ZN(n10059) );
  OR2_X1 U5527 ( .A1(n10982), .A2(n10541), .ZN(n10048) );
  NOR2_X2 U5528 ( .A1(n10048), .A2(n10534), .ZN(n10047) );
  OAI21_X1 U5529 ( .B1(n10970), .B2(n5596), .A(n5592), .ZN(n10046) );
  AOI21_X1 U5530 ( .B1(n5595), .B2(n10974), .A(n5088), .ZN(n5592) );
  INV_X1 U5531 ( .A(n10968), .ZN(n5594) );
  AND2_X1 U5532 ( .A1(n10059), .A2(n10057), .ZN(n10054) );
  NAND2_X1 U5533 ( .A1(n10970), .A2(n10969), .ZN(n10968) );
  NOR2_X2 U5534 ( .A1(n8391), .A2(n8554), .ZN(n10983) );
  NAND2_X1 U5535 ( .A1(n8240), .A2(n5569), .ZN(n5280) );
  NOR2_X1 U5536 ( .A1(n5572), .A2(n8991), .ZN(n5569) );
  NAND2_X1 U5537 ( .A1(n5399), .A2(n8917), .ZN(n5398) );
  NAND2_X1 U5538 ( .A1(n9004), .A2(n8917), .ZN(n5401) );
  NAND2_X1 U5539 ( .A1(n8254), .A2(n5572), .ZN(n8388) );
  OR2_X1 U5540 ( .A1(n7974), .A2(n8120), .ZN(n5273) );
  NAND2_X1 U5541 ( .A1(n7884), .A2(n7858), .ZN(n7918) );
  NAND2_X1 U5542 ( .A1(n7527), .A2(n8862), .ZN(n5394) );
  NAND2_X1 U5543 ( .A1(n5395), .A2(n8882), .ZN(n8865) );
  NAND2_X1 U5544 ( .A1(n7508), .A2(n7507), .ZN(n7515) );
  AND2_X1 U5545 ( .A1(n7135), .A2(n7506), .ZN(n10975) );
  NAND2_X1 U5546 ( .A1(n7163), .A2(n7164), .ZN(n7271) );
  NAND2_X1 U5547 ( .A1(n8748), .A2(n8747), .ZN(n10078) );
  OR2_X1 U5548 ( .A1(n9924), .A2(n9923), .ZN(n10095) );
  NAND2_X1 U5549 ( .A1(n8612), .A2(n8611), .ZN(n10130) );
  NAND3_X1 U5550 ( .A1(n5284), .A2(n5283), .A3(n5281), .ZN(n6802) );
  NOR2_X1 U5551 ( .A1(n5093), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5282) );
  NOR2_X1 U5552 ( .A1(n5264), .A2(n6811), .ZN(n5263) );
  NAND2_X1 U5553 ( .A1(n5637), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n6811) );
  INV_X1 U5554 ( .A(n6680), .ZN(n5264) );
  NAND2_X1 U5555 ( .A1(n6315), .A2(n6284), .ZN(n8789) );
  OR2_X1 U5556 ( .A1(n6283), .A2(n6282), .ZN(n6284) );
  XNOR2_X1 U5557 ( .A(n6277), .B(n6276), .ZN(n9697) );
  NAND2_X1 U5558 ( .A1(n6257), .A2(n6256), .ZN(n6277) );
  NAND2_X1 U5559 ( .A1(n6143), .A2(n6142), .ZN(n6161) );
  NAND2_X1 U5560 ( .A1(n5431), .A2(n6030), .ZN(n6050) );
  NAND2_X1 U5561 ( .A1(n5212), .A2(n5215), .ZN(n5431) );
  OAI21_X1 U5562 ( .B1(n6009), .B2(n5218), .A(n6008), .ZN(n6028) );
  NAND2_X1 U5563 ( .A1(n5410), .A2(n5937), .ZN(n5945) );
  XNOR2_X1 U5564 ( .A(n5803), .B(n5782), .ZN(n5801) );
  XNOR2_X1 U5565 ( .A(n5780), .B(n10193), .ZN(n5778) );
  XNOR2_X1 U5566 ( .A(n5757), .B(n5747), .ZN(n5755) );
  NAND2_X1 U5567 ( .A1(n5204), .A2(n5746), .ZN(n5756) );
  AND2_X1 U5568 ( .A1(n6272), .A2(n6271), .ZN(n9198) );
  OR2_X1 U5569 ( .A1(n9408), .A2(n6357), .ZN(n6272) );
  OAI21_X1 U5570 ( .B1(n5633), .B2(n6312), .A(n5495), .ZN(n5494) );
  NAND2_X1 U5571 ( .A1(n5499), .A2(n6312), .ZN(n5495) );
  OAI21_X1 U5572 ( .B1(n5633), .B2(n6311), .A(n5498), .ZN(n5497) );
  NAND2_X1 U5573 ( .A1(n5499), .A2(n6311), .ZN(n5498) );
  AND2_X1 U5574 ( .A1(n9592), .A2(n5500), .ZN(n5499) );
  NAND2_X1 U5575 ( .A1(n9099), .A2(n5042), .ZN(n5500) );
  NAND2_X1 U5576 ( .A1(n6298), .A2(n6297), .ZN(n6313) );
  NAND2_X1 U5577 ( .A1(n6228), .A2(n6227), .ZN(n9196) );
  NAND2_X1 U5578 ( .A1(n5974), .A2(n5973), .ZN(n10938) );
  AND2_X1 U5579 ( .A1(n6154), .A2(n6153), .ZN(n9266) );
  NAND2_X1 U5580 ( .A1(n6308), .A2(n6307), .ZN(n9393) );
  OR2_X1 U5581 ( .A1(n6368), .A2(n6357), .ZN(n6308) );
  INV_X1 U5582 ( .A(n9198), .ZN(n9392) );
  NAND2_X1 U5583 ( .A1(n5768), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5695) );
  AND2_X1 U5584 ( .A1(n6010), .A2(n5992), .ZN(n8199) );
  NOR2_X1 U5585 ( .A1(n9365), .A2(n9580), .ZN(n5294) );
  OR2_X1 U5586 ( .A1(n9364), .A2(n5293), .ZN(n5290) );
  INV_X1 U5587 ( .A(n9580), .ZN(n5293) );
  NAND2_X1 U5588 ( .A1(n9365), .A2(n9580), .ZN(n5292) );
  NAND2_X1 U5589 ( .A1(n5601), .A2(n5083), .ZN(n5600) );
  INV_X1 U5590 ( .A(n9384), .ZN(n5601) );
  OAI21_X1 U5591 ( .B1(n9088), .B2(n5604), .A(n5603), .ZN(n5602) );
  OAI21_X1 U5592 ( .B1(n5606), .B2(n9088), .A(n5604), .ZN(n5603) );
  XNOR2_X1 U5593 ( .A(n9090), .B(n9089), .ZN(n5202) );
  NAND2_X1 U5594 ( .A1(n5203), .A2(n5199), .ZN(n5198) );
  NAND2_X1 U5595 ( .A1(n9095), .A2(n5200), .ZN(n5199) );
  AOI21_X1 U5596 ( .B1(n9587), .B2(n9568), .A(n9096), .ZN(n5203) );
  XNOR2_X1 U5597 ( .A(n5169), .B(n9082), .ZN(n9596) );
  OAI21_X1 U5598 ( .B1(n9398), .B2(n5165), .A(n5163), .ZN(n5169) );
  AOI21_X1 U5599 ( .B1(n9080), .B2(n5164), .A(n5607), .ZN(n5163) );
  NAND2_X1 U5600 ( .A1(n9080), .A2(n5166), .ZN(n5165) );
  NAND2_X1 U5601 ( .A1(n5614), .A2(n5611), .ZN(n9428) );
  OR2_X1 U5602 ( .A1(n5762), .A2(n7114), .ZN(n5682) );
  NOR3_X1 U5603 ( .A1(n5673), .A2(n5054), .A3(P2_IR_REG_29__SCAN_IN), .ZN(
        n5195) );
  AND2_X1 U5604 ( .A1(n8729), .A2(n5548), .ZN(n5541) );
  NAND2_X1 U5605 ( .A1(n5542), .A2(n5535), .ZN(n5534) );
  NOR2_X1 U5606 ( .A1(n5548), .A2(n5540), .ZN(n5535) );
  AOI21_X1 U5607 ( .B1(n5056), .B2(n9744), .A(n5539), .ZN(n5538) );
  NAND2_X1 U5608 ( .A1(n8741), .A2(n8742), .ZN(n5539) );
  AND2_X1 U5609 ( .A1(n9733), .A2(n9732), .ZN(n5253) );
  NAND2_X1 U5610 ( .A1(n8706), .A2(n8705), .ZN(n5252) );
  NAND2_X1 U5611 ( .A1(n8245), .A2(n8244), .ZN(n8511) );
  XNOR2_X1 U5612 ( .A(n7238), .B(n7239), .ZN(n7236) );
  NAND2_X1 U5613 ( .A1(n5251), .A2(n5506), .ZN(n8273) );
  OR2_X1 U5614 ( .A1(n8221), .A2(n8220), .ZN(n5506) );
  OAI21_X1 U5615 ( .B1(n9755), .B2(n9756), .A(n5254), .ZN(n9735) );
  NAND2_X1 U5616 ( .A1(n8703), .A2(n5255), .ZN(n5254) );
  INV_X1 U5617 ( .A(n8704), .ZN(n5255) );
  NAND2_X1 U5618 ( .A1(n8690), .A2(n8689), .ZN(n10105) );
  INV_X1 U5619 ( .A(n5545), .ZN(n9803) );
  AOI21_X1 U5620 ( .B1(n5406), .B2(n10980), .A(n5259), .ZN(n10081) );
  INV_X1 U5621 ( .A(n5404), .ZN(n5259) );
  XNOR2_X1 U5622 ( .A(n9159), .B(n5073), .ZN(n5406) );
  AOI21_X1 U5623 ( .B1(n9905), .B2(n10975), .A(n5405), .ZN(n5404) );
  XNOR2_X1 U5624 ( .A(n9150), .B(n5073), .ZN(n10082) );
  NOR2_X1 U5625 ( .A1(n9149), .A2(n9148), .ZN(n9150) );
  AND2_X1 U5626 ( .A1(n10083), .A2(n9905), .ZN(n9148) );
  OR2_X1 U5627 ( .A1(n9149), .A2(n5583), .ZN(n10087) );
  INV_X1 U5628 ( .A(n5590), .ZN(n5583) );
  OR2_X1 U5629 ( .A1(n7185), .A2(n7114), .ZN(n7115) );
  INV_X1 U5630 ( .A(n7207), .ZN(n7418) );
  AOI21_X1 U5631 ( .B1(n10071), .B2(n10981), .A(n5308), .ZN(n5307) );
  NAND2_X1 U5632 ( .A1(n10990), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U5633 ( .A1(n5591), .A2(n5082), .ZN(n5586) );
  AOI22_X1 U5634 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_128), .B1(SI_31_), 
        .B2(keyinput_129), .ZN(n10148) );
  NAND2_X1 U5635 ( .A1(n5380), .A2(n5378), .ZN(n10164) );
  NAND2_X1 U5636 ( .A1(n5368), .A2(n10183), .ZN(n5367) );
  NAND2_X1 U5637 ( .A1(n10175), .A2(n10174), .ZN(n5368) );
  NOR2_X1 U5638 ( .A1(n10182), .A2(n10181), .ZN(n5366) );
  AOI21_X1 U5639 ( .B1(n5365), .B2(n5364), .A(n5363), .ZN(n10188) );
  XNOR2_X1 U5640 ( .A(SI_11_), .B(keyinput_149), .ZN(n5363) );
  INV_X1 U5641 ( .A(n10184), .ZN(n5364) );
  NAND2_X1 U5642 ( .A1(n5367), .A2(n5366), .ZN(n5365) );
  NAND2_X1 U5643 ( .A1(n5384), .A2(n5382), .ZN(n10206) );
  NOR2_X1 U5644 ( .A1(n5383), .A2(n10205), .ZN(n5382) );
  OAI21_X1 U5645 ( .B1(n5385), .B2(n10194), .A(n5121), .ZN(n5384) );
  NAND2_X1 U5646 ( .A1(n5349), .A2(n5348), .ZN(n10221) );
  AND2_X1 U5647 ( .A1(n10216), .A2(n10215), .ZN(n5348) );
  NAND2_X1 U5648 ( .A1(n5352), .A2(n5350), .ZN(n5349) );
  OAI21_X1 U5649 ( .B1(n5346), .B2(n10229), .A(n5344), .ZN(n10236) );
  NAND2_X1 U5650 ( .A1(keyinput_217), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n5376)
         );
  INV_X1 U5651 ( .A(n5372), .ZN(n5371) );
  OAI21_X1 U5652 ( .B1(n5373), .B2(n10291), .A(n5374), .ZN(n5372) );
  INV_X1 U5653 ( .A(n10298), .ZN(n5374) );
  AOI21_X1 U5654 ( .B1(n5128), .B2(n10288), .A(n5375), .ZN(n5373) );
  AOI221_X1 U5655 ( .B1(n10276), .B2(n10275), .C1(keyinput_206), .C2(n10274), 
        .A(n10273), .ZN(n10285) );
  AOI21_X1 U5656 ( .B1(n5371), .B2(n5064), .A(n5129), .ZN(n5370) );
  AND2_X1 U5657 ( .A1(n5130), .A2(n5362), .ZN(n5361) );
  OR2_X1 U5658 ( .A1(n10322), .A2(n5063), .ZN(n5362) );
  AOI21_X1 U5659 ( .B1(n5361), .B2(n5063), .A(n5131), .ZN(n5360) );
  OAI21_X1 U5660 ( .B1(n9580), .B2(n6531), .A(n5437), .ZN(n6544) );
  NAND2_X1 U5661 ( .A1(n6543), .A2(n6531), .ZN(n5437) );
  INV_X1 U5662 ( .A(n9914), .ZN(n5392) );
  AND2_X1 U5663 ( .A1(n9904), .A2(n9903), .ZN(n5393) );
  OAI211_X1 U5664 ( .C1(n10314), .C2(n10313), .A(n10312), .B(n10311), .ZN(
        n10323) );
  AOI21_X1 U5665 ( .B1(n5360), .B2(n5358), .A(n5133), .ZN(n5357) );
  INV_X1 U5666 ( .A(n5361), .ZN(n5358) );
  INV_X1 U5667 ( .A(n5360), .ZN(n5359) );
  INV_X1 U5668 ( .A(n5435), .ZN(n5434) );
  OAI21_X1 U5669 ( .B1(n6282), .B2(n5436), .A(n6380), .ZN(n5435) );
  INV_X1 U5670 ( .A(n6314), .ZN(n5436) );
  INV_X1 U5671 ( .A(SI_28_), .ZN(n10153) );
  AND2_X1 U5672 ( .A1(n5238), .A2(n6276), .ZN(n5237) );
  NAND2_X1 U5673 ( .A1(n6239), .A2(n6256), .ZN(n5238) );
  INV_X1 U5674 ( .A(n6256), .ZN(n5235) );
  AND2_X1 U5675 ( .A1(n5416), .A2(n5115), .ZN(n5230) );
  INV_X1 U5676 ( .A(n5417), .ZN(n5416) );
  OAI21_X1 U5677 ( .B1(n6167), .B2(n5418), .A(n6209), .ZN(n5417) );
  INV_X1 U5678 ( .A(n6189), .ZN(n5418) );
  AOI21_X1 U5679 ( .B1(n5215), .B2(n5214), .A(n5119), .ZN(n5213) );
  INV_X1 U5680 ( .A(n6008), .ZN(n5214) );
  NAND2_X1 U5681 ( .A1(n5218), .A2(n6008), .ZN(n5217) );
  INV_X1 U5682 ( .A(n6026), .ZN(n6027) );
  NAND2_X1 U5683 ( .A1(n5941), .A2(n10146), .ZN(n5966) );
  NOR2_X1 U5684 ( .A1(n6147), .A2(n5141), .ZN(n5140) );
  NAND2_X1 U5685 ( .A1(n9580), .A2(n6543), .ZN(n6624) );
  OR2_X1 U5686 ( .A1(n9603), .A2(n9198), .ZN(n6549) );
  NOR2_X1 U5687 ( .A1(n5085), .A2(n9420), .ZN(n5458) );
  NAND2_X1 U5688 ( .A1(n5096), .A2(n5297), .ZN(n5296) );
  INV_X1 U5689 ( .A(n5298), .ZN(n5297) );
  NAND2_X1 U5690 ( .A1(n9454), .A2(n9074), .ZN(n5298) );
  OR2_X1 U5691 ( .A1(n9634), .A2(n9510), .ZN(n6604) );
  INV_X1 U5692 ( .A(n6016), .ZN(n6014) );
  NOR2_X1 U5693 ( .A1(n6059), .A2(n9319), .ZN(n5136) );
  INV_X1 U5694 ( .A(n8416), .ZN(n5468) );
  OR2_X1 U5695 ( .A1(n6599), .A2(n6598), .ZN(n5462) );
  NOR2_X1 U5696 ( .A1(n8364), .A2(n5466), .ZN(n5465) );
  NAND2_X1 U5697 ( .A1(n5137), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6016) );
  AND2_X1 U5698 ( .A1(n6481), .A2(n6592), .ZN(n8081) );
  NAND2_X1 U5699 ( .A1(n9280), .A2(n10759), .ZN(n6449) );
  NAND2_X1 U5700 ( .A1(n6434), .A2(n6433), .ZN(n5597) );
  OR2_X1 U5701 ( .A1(n9592), .A2(n9385), .ZN(n9376) );
  NAND2_X1 U5702 ( .A1(n6319), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6323) );
  NOR2_X1 U5703 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5644) );
  INV_X1 U5704 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5949) );
  OR2_X1 U5705 ( .A1(n5827), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5853) );
  AND2_X1 U5706 ( .A1(n8498), .A2(n8497), .ZN(n5528) );
  INV_X1 U5707 ( .A(n8506), .ZN(n5525) );
  INV_X1 U5708 ( .A(n7832), .ZN(n5522) );
  NOR2_X1 U5709 ( .A1(n5522), .A2(n5523), .ZN(n5521) );
  INV_X1 U5710 ( .A(n7690), .ZN(n5523) );
  NAND2_X1 U5711 ( .A1(n5511), .A2(n8647), .ZN(n5228) );
  NAND2_X1 U5712 ( .A1(n5071), .A2(n8647), .ZN(n5226) );
  AND2_X1 U5713 ( .A1(n7255), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7352) );
  AND3_X1 U5714 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n7255) );
  OR2_X1 U5715 ( .A1(n10078), .A2(n9133), .ZN(n9014) );
  NOR2_X1 U5716 ( .A1(n10088), .A2(n10083), .ZN(n5321) );
  INV_X1 U5717 ( .A(n5567), .ZN(n5566) );
  INV_X1 U5718 ( .A(n8603), .ZN(n7367) );
  NOR2_X1 U5719 ( .A1(n10120), .A2(n10126), .ZN(n5316) );
  NOR2_X1 U5720 ( .A1(n8470), .A2(n5326), .ZN(n5325) );
  INV_X1 U5721 ( .A(n8922), .ZN(n5326) );
  AND2_X1 U5722 ( .A1(n8255), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6847) );
  OR2_X1 U5723 ( .A1(n8247), .A2(n8246), .ZN(n8257) );
  NAND2_X1 U5724 ( .A1(n8991), .A2(n8820), .ZN(n5399) );
  NOR2_X1 U5725 ( .A1(n7518), .A2(n7517), .ZN(n6823) );
  AND2_X1 U5726 ( .A1(n9155), .A2(n9157), .ZN(n9130) );
  NAND2_X1 U5727 ( .A1(n8789), .A2(n8749), .ZN(n5243) );
  OAI21_X1 U5728 ( .B1(n10038), .B2(n5330), .A(n5327), .ZN(n9996) );
  AOI21_X1 U5729 ( .B1(n10012), .B2(n5329), .A(n5328), .ZN(n5327) );
  INV_X1 U5730 ( .A(n9122), .ZN(n5329) );
  NAND2_X1 U5731 ( .A1(n10011), .A2(n10012), .ZN(n10010) );
  NAND2_X1 U5732 ( .A1(n5509), .A2(n10021), .ZN(n8972) );
  INV_X1 U5733 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6656) );
  NAND2_X1 U5734 ( .A1(n5284), .A2(n5517), .ZN(n6669) );
  AND2_X1 U5735 ( .A1(n5053), .A2(n6653), .ZN(n5517) );
  INV_X1 U5736 ( .A(n6005), .ZN(n5218) );
  XNOR2_X1 U5737 ( .A(n5936), .B(n5918), .ZN(n5935) );
  AND2_X1 U5738 ( .A1(n5895), .A2(n5874), .ZN(n5875) );
  XNOR2_X1 U5739 ( .A(n5846), .B(SI_7_), .ZN(n5843) );
  NAND2_X1 U5740 ( .A1(n5139), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5857) );
  INV_X1 U5741 ( .A(n5831), .ZN(n5139) );
  OR2_X1 U5742 ( .A1(n6131), .A2(n10228), .ZN(n6147) );
  NAND2_X1 U5743 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5791) );
  AND2_X1 U5744 ( .A1(n5754), .A2(n5736), .ZN(n5484) );
  INV_X1 U5745 ( .A(n7733), .ZN(n5754) );
  OR2_X1 U5746 ( .A1(n5857), .A2(n7650), .ZN(n5883) );
  NAND2_X1 U5747 ( .A1(n5140), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6196) );
  INV_X1 U5748 ( .A(n5140), .ZN(n6174) );
  NAND2_X1 U5749 ( .A1(n5477), .A2(n5476), .ZN(n9226) );
  AND2_X1 U5750 ( .A1(n6187), .A2(n6158), .ZN(n5476) );
  OR2_X1 U5751 ( .A1(n7844), .A2(n7845), .ZN(n9237) );
  CLKBUF_X1 U5752 ( .A(n7566), .Z(n9182) );
  AND2_X1 U5753 ( .A1(n5471), .A2(n8766), .ZN(n5470) );
  NAND2_X1 U5754 ( .A1(n5473), .A2(n5475), .ZN(n5471) );
  OR2_X1 U5755 ( .A1(n6995), .A2(n6994), .ZN(n5145) );
  AND2_X1 U5756 ( .A1(n7794), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5147) );
  NAND2_X1 U5757 ( .A1(n5072), .A2(n9283), .ZN(n9282) );
  NOR2_X1 U5758 ( .A1(n7906), .A2(n5155), .ZN(n7910) );
  AND2_X1 U5759 ( .A1(n7907), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5155) );
  NAND2_X1 U5760 ( .A1(n7910), .A2(n7909), .ZN(n8050) );
  NAND2_X1 U5761 ( .A1(n8050), .A2(n5154), .ZN(n8052) );
  OR2_X1 U5762 ( .A1(n8051), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5154) );
  NOR2_X1 U5763 ( .A1(n9082), .A2(n5143), .ZN(n5606) );
  AND2_X1 U5764 ( .A1(n9592), .A2(n9166), .ZN(n5444) );
  INV_X1 U5765 ( .A(n9401), .ZN(n5166) );
  NOR2_X1 U5766 ( .A1(n9392), .A2(n9603), .ZN(n5164) );
  AND2_X1 U5767 ( .A1(n6301), .A2(n6289), .ZN(n9388) );
  NOR3_X1 U5768 ( .A1(n9603), .A2(n9477), .A3(n5296), .ZN(n9405) );
  AND2_X1 U5769 ( .A1(n6549), .A2(n6614), .ZN(n9401) );
  NOR2_X1 U5770 ( .A1(n9477), .A2(n5296), .ZN(n9413) );
  NAND2_X1 U5771 ( .A1(n5610), .A2(n5612), .ZN(n9412) );
  INV_X1 U5772 ( .A(n5613), .ZN(n5612) );
  OAI21_X1 U5773 ( .B1(n5615), .B2(n9443), .A(n9077), .ZN(n5613) );
  OR2_X1 U5774 ( .A1(n9415), .A2(n6357), .ZN(n6251) );
  AND2_X1 U5775 ( .A1(n6203), .A2(n6202), .ZN(n9436) );
  NOR2_X1 U5776 ( .A1(n9477), .A2(n5298), .ZN(n9449) );
  NOR2_X1 U5777 ( .A1(n9477), .A2(n9624), .ZN(n9461) );
  NAND2_X1 U5778 ( .A1(n5136), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U5779 ( .A1(n9524), .A2(n9268), .ZN(n5182) );
  NAND2_X1 U5780 ( .A1(n9526), .A2(n9517), .ZN(n5183) );
  AOI21_X1 U5781 ( .B1(n9518), .B2(n9525), .A(n5175), .ZN(n9506) );
  NOR2_X1 U5782 ( .A1(n9644), .A2(n9268), .ZN(n5175) );
  OR2_X1 U5783 ( .A1(n9644), .A2(n9521), .ZN(n9519) );
  NAND2_X1 U5784 ( .A1(n5176), .A2(n5621), .ZN(n9518) );
  INV_X1 U5785 ( .A(n5622), .ZN(n5621) );
  NAND2_X1 U5786 ( .A1(n8423), .A2(n5620), .ZN(n5176) );
  OAI21_X1 U5787 ( .B1(n5624), .B2(n5626), .A(n9067), .ZN(n5622) );
  AND3_X1 U5788 ( .A1(n8430), .A2(n5303), .A3(n8101), .ZN(n9534) );
  OAI22_X1 U5789 ( .A1(n8441), .A2(n8445), .B1(n9270), .B2(n9659), .ZN(n8423)
         );
  AND2_X1 U5790 ( .A1(n6600), .A2(n6596), .ZN(n8424) );
  AND4_X1 U5791 ( .A1(n6021), .A2(n6020), .A3(n6019), .A4(n6018), .ZN(n8422)
         );
  AND2_X1 U5792 ( .A1(n6594), .A2(n6491), .ZN(n8360) );
  NOR2_X1 U5793 ( .A1(n8359), .A2(n8360), .ZN(n8420) );
  NAND2_X1 U5794 ( .A1(n8101), .A2(n8358), .ZN(n8429) );
  AND4_X1 U5795 ( .A1(n5980), .A2(n5979), .A3(n5978), .A4(n5977), .ZN(n8767)
         );
  NAND2_X1 U5796 ( .A1(n8033), .A2(n8032), .ZN(n8080) );
  AND4_X1 U5797 ( .A1(n5909), .A2(n5908), .A3(n5907), .A4(n5906), .ZN(n9239)
         );
  AND4_X1 U5798 ( .A1(n5960), .A2(n5959), .A3(n5958), .A4(n5957), .ZN(n8559)
         );
  NAND2_X1 U5799 ( .A1(n7985), .A2(n6589), .ZN(n8035) );
  AND4_X1 U5800 ( .A1(n5888), .A2(n5887), .A3(n5886), .A4(n5885), .ZN(n7986)
         );
  NAND2_X1 U5801 ( .A1(n9565), .A2(n5302), .ZN(n7992) );
  AOI21_X1 U5802 ( .B1(n7763), .B2(n7779), .A(n6586), .ZN(n7949) );
  NAND2_X1 U5803 ( .A1(n9565), .A2(n10830), .ZN(n7811) );
  NAND2_X1 U5804 ( .A1(n6581), .A2(n5454), .ZN(n5450) );
  AND3_X1 U5805 ( .A1(n6578), .A2(n7774), .A3(n6579), .ZN(n5177) );
  NAND2_X1 U5806 ( .A1(n5809), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5831) );
  INV_X1 U5807 ( .A(n5811), .ZN(n5809) );
  NAND2_X1 U5808 ( .A1(n5138), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5811) );
  INV_X1 U5809 ( .A(n5791), .ZN(n5138) );
  OR2_X1 U5810 ( .A1(n7752), .A2(n9214), .ZN(n10783) );
  NAND2_X1 U5811 ( .A1(n7710), .A2(n10759), .ZN(n7752) );
  NAND2_X1 U5812 ( .A1(n7717), .A2(n7678), .ZN(n7680) );
  AND2_X1 U5813 ( .A1(n10752), .A2(n5287), .ZN(n7710) );
  INV_X1 U5814 ( .A(n7711), .ZN(n5287) );
  NAND2_X1 U5815 ( .A1(n7674), .A2(n9102), .ZN(n7711) );
  NAND2_X1 U5816 ( .A1(n7144), .A2(n9180), .ZN(n7676) );
  AND2_X1 U5817 ( .A1(n6349), .A2(n6348), .ZN(n7288) );
  NAND2_X1 U5818 ( .A1(n6423), .A2(n6422), .ZN(n9083) );
  NAND2_X1 U5819 ( .A1(n6058), .A2(n6057), .ZN(n9651) );
  NAND2_X1 U5820 ( .A1(n7749), .A2(n7748), .ZN(n7751) );
  AND2_X1 U5821 ( .A1(n6660), .A2(n10694), .ZN(n10614) );
  XNOR2_X1 U5822 ( .A(n5675), .B(n5685), .ZN(n6365) );
  NAND2_X1 U5823 ( .A1(n5674), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5675) );
  XNOR2_X1 U5824 ( .A(n5677), .B(n5684), .ZN(n6634) );
  NAND2_X1 U5825 ( .A1(n5676), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5677) );
  XNOR2_X1 U5826 ( .A(n6323), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6355) );
  XNOR2_X1 U5827 ( .A(n5664), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6435) );
  NOR2_X1 U5828 ( .A1(n8114), .A2(n5516), .ZN(n5515) );
  INV_X1 U5829 ( .A(n8109), .ZN(n5516) );
  INV_X1 U5830 ( .A(n9802), .ZN(n5548) );
  XNOR2_X1 U5831 ( .A(n7119), .B(n8793), .ZN(n7126) );
  NAND2_X1 U5832 ( .A1(n7118), .A2(n7117), .ZN(n7119) );
  NAND2_X1 U5833 ( .A1(n9743), .A2(n5514), .ZN(n5513) );
  OR2_X1 U5834 ( .A1(n8650), .A2(n8649), .ZN(n5561) );
  NAND2_X1 U5835 ( .A1(n5502), .A2(n5222), .ZN(n5220) );
  NAND2_X1 U5836 ( .A1(n8985), .A2(n6957), .ZN(n7205) );
  NAND2_X1 U5837 ( .A1(n10078), .A2(n9133), .ZN(n9024) );
  OR2_X1 U5838 ( .A1(n6916), .A2(n6915), .ZN(n6913) );
  AND2_X1 U5839 ( .A1(n9160), .A2(n9816), .ZN(n5405) );
  AOI21_X1 U5840 ( .B1(n9158), .B2(n9157), .A(n9156), .ZN(n9159) );
  AND2_X1 U5841 ( .A1(n8734), .A2(n8733), .ZN(n9138) );
  AND2_X1 U5842 ( .A1(n9924), .A2(n9902), .ZN(n9899) );
  NAND2_X1 U5843 ( .A1(n9938), .A2(n9955), .ZN(n9933) );
  AND2_X1 U5844 ( .A1(n8956), .A2(n9127), .ZN(n9952) );
  AND2_X1 U5845 ( .A1(n8953), .A2(n9126), .ZN(n9970) );
  AND2_X1 U5846 ( .A1(n10032), .A2(n5061), .ZN(n9965) );
  NAND2_X1 U5847 ( .A1(n10032), .A2(n5316), .ZN(n9993) );
  NAND2_X1 U5848 ( .A1(n10032), .A2(n5314), .ZN(n9979) );
  NOR2_X1 U5849 ( .A1(n8615), .A2(n8614), .ZN(n8613) );
  AND2_X1 U5850 ( .A1(n10047), .A2(n10037), .ZN(n10032) );
  AND2_X1 U5851 ( .A1(n8813), .A2(n8936), .ZN(n9120) );
  NAND2_X1 U5852 ( .A1(n8942), .A2(n9122), .ZN(n10031) );
  AND2_X1 U5853 ( .A1(n8936), .A2(n8935), .ZN(n10060) );
  NOR2_X1 U5854 ( .A1(n9009), .A2(n5279), .ZN(n5278) );
  INV_X1 U5855 ( .A(n5570), .ZN(n5279) );
  NAND2_X1 U5856 ( .A1(n8240), .A2(n8239), .ZN(n8290) );
  NAND2_X1 U5857 ( .A1(n5311), .A2(n5058), .ZN(n8302) );
  NAND2_X1 U5858 ( .A1(n8253), .A2(n5402), .ZN(n8293) );
  INV_X1 U5859 ( .A(n5399), .ZN(n5402) );
  AND2_X1 U5860 ( .A1(n8253), .A2(n8820), .ZN(n8294) );
  INV_X1 U5861 ( .A(n5387), .ZN(n8138) );
  AOI21_X1 U5862 ( .B1(n7935), .B2(n8902), .A(n5388), .ZN(n5387) );
  NAND2_X1 U5863 ( .A1(n5389), .A2(n8905), .ZN(n5388) );
  OR2_X1 U5864 ( .A1(n8139), .A2(n8135), .ZN(n8253) );
  NAND2_X1 U5865 ( .A1(n5311), .A2(n5309), .ZN(n8300) );
  OR2_X1 U5866 ( .A1(n7923), .A2(n7922), .ZN(n7925) );
  NOR2_X1 U5867 ( .A1(n7938), .A2(n10872), .ZN(n8023) );
  NOR3_X1 U5868 ( .A1(n7938), .A2(n8170), .A3(n10872), .ZN(n8150) );
  AOI21_X1 U5869 ( .B1(n5271), .B2(n5269), .A(n5089), .ZN(n5268) );
  INV_X1 U5870 ( .A(n5273), .ZN(n5269) );
  INV_X1 U5871 ( .A(n5271), .ZN(n5270) );
  NAND2_X1 U5872 ( .A1(n8019), .A2(n8902), .ZN(n8137) );
  OR2_X1 U5873 ( .A1(n7867), .A2(n7866), .ZN(n7923) );
  NAND2_X1 U5874 ( .A1(n5390), .A2(n9003), .ZN(n8019) );
  INV_X1 U5875 ( .A(n7935), .ZN(n5390) );
  NAND2_X1 U5876 ( .A1(n7862), .A2(n7861), .ZN(n7974) );
  OR2_X1 U5877 ( .A1(n7894), .A2(n7974), .ZN(n7938) );
  NAND2_X1 U5878 ( .A1(n7856), .A2(n7855), .ZN(n7886) );
  AND2_X1 U5879 ( .A1(n7531), .A2(n7854), .ZN(n7893) );
  AND2_X1 U5880 ( .A1(n7552), .A2(n7447), .ZN(n7449) );
  NAND2_X1 U5881 ( .A1(n7449), .A2(n7448), .ZN(n7508) );
  NOR2_X1 U5882 ( .A1(n7543), .A2(n7472), .ZN(n7531) );
  OR2_X1 U5883 ( .A1(n7545), .A2(n7558), .ZN(n7543) );
  NAND2_X1 U5884 ( .A1(n7491), .A2(n8993), .ZN(n7490) );
  NAND2_X1 U5885 ( .A1(n7279), .A2(n7278), .ZN(n8856) );
  OAI221_X1 U5886 ( .B1(n10347), .B2(n10346), .C1(n10583), .C2(keyinput_254), 
        .A(n10345), .ZN(n10349) );
  NAND2_X1 U5887 ( .A1(n8640), .A2(n8639), .ZN(n10534) );
  NAND2_X1 U5888 ( .A1(n8468), .A2(n8467), .ZN(n10541) );
  XNOR2_X1 U5889 ( .A(n6410), .B(n6409), .ZN(n9693) );
  XNOR2_X1 U5890 ( .A(n6420), .B(n6419), .ZN(n9060) );
  XNOR2_X1 U5891 ( .A(n6381), .B(n6380), .ZN(n9144) );
  NAND2_X1 U5892 ( .A1(n6315), .A2(n6314), .ZN(n6381) );
  INV_X1 U5893 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6678) );
  INV_X1 U5894 ( .A(n6930), .ZN(n5578) );
  INV_X1 U5895 ( .A(n6162), .ZN(n6168) );
  INV_X1 U5896 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6672) );
  INV_X1 U5897 ( .A(n6126), .ZN(n6123) );
  OR2_X1 U5898 ( .A1(n6710), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n6706) );
  OR2_X1 U5899 ( .A1(n6706), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6742) );
  NAND2_X1 U5900 ( .A1(n5206), .A2(n5804), .ZN(n5823) );
  INV_X1 U5901 ( .A(n5332), .ZN(n5331) );
  NOR2_X1 U5902 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n6643) );
  NAND2_X1 U5903 ( .A1(n5205), .A2(n5719), .ZN(n5743) );
  NAND2_X1 U5904 ( .A1(n7588), .A2(n5821), .ZN(n7593) );
  AND2_X1 U5905 ( .A1(n5841), .A2(n5821), .ZN(n5486) );
  AOI21_X1 U5906 ( .B1(n5481), .B2(n5483), .A(n5117), .ZN(n5478) );
  NAND2_X1 U5907 ( .A1(n6287), .A2(n6286), .ZN(n9597) );
  NAND2_X1 U5908 ( .A1(n8789), .A2(n6421), .ZN(n6287) );
  NAND2_X1 U5909 ( .A1(n6195), .A2(n6194), .ZN(n9618) );
  NAND2_X1 U5910 ( .A1(n7570), .A2(n5736), .ZN(n7732) );
  NAND2_X1 U5911 ( .A1(n6146), .A2(n6145), .ZN(n9629) );
  AND4_X1 U5912 ( .A1(n5930), .A2(n5929), .A3(n5928), .A4(n5927), .ZN(n8075)
         );
  NAND2_X1 U5913 ( .A1(n6243), .A2(n6242), .ZN(n9608) );
  AND3_X1 U5914 ( .A1(n6044), .A2(n6043), .A3(n6042), .ZN(n9540) );
  NAND2_X1 U5915 ( .A1(n8197), .A2(n6049), .ZN(n6663) );
  NAND2_X1 U5916 ( .A1(n6213), .A2(n6212), .ZN(n9612) );
  AND2_X1 U5917 ( .A1(n6112), .A2(n6111), .ZN(n9068) );
  NAND2_X1 U5918 ( .A1(n5472), .A2(n8557), .ZN(n8771) );
  NAND2_X1 U5919 ( .A1(n8561), .A2(n5965), .ZN(n5472) );
  AND2_X1 U5920 ( .A1(n9257), .A2(n10789), .ZN(n9247) );
  AND4_X1 U5921 ( .A1(n5741), .A2(n5740), .A3(n5739), .A4(n5738), .ZN(n6445)
         );
  AND3_X1 U5922 ( .A1(n6063), .A2(n6062), .A3(n6061), .ZN(n9066) );
  AND2_X1 U5923 ( .A1(n6375), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9246) );
  NAND2_X1 U5924 ( .A1(n5480), .A2(n6255), .ZN(n9253) );
  NAND2_X1 U5925 ( .A1(n9196), .A2(n9195), .ZN(n5480) );
  AND4_X1 U5926 ( .A1(n6001), .A2(n6000), .A3(n5999), .A4(n5998), .ZN(n9052)
         );
  CLKBUF_X1 U5927 ( .A(n8190), .Z(n9059) );
  INV_X1 U5928 ( .A(n9247), .ZN(n9230) );
  NAND2_X1 U5929 ( .A1(n6571), .A2(n5423), .ZN(n5422) );
  INV_X1 U5930 ( .A(n9436), .ZN(n9468) );
  OR2_X1 U5931 ( .A1(n6989), .A2(n6661), .ZN(n9267) );
  NAND4_X2 U5932 ( .A1(n5772), .A2(n5771), .A3(n5770), .A4(n5769), .ZN(n10790)
         );
  NAND3_X1 U5933 ( .A1(n5702), .A2(n5193), .A3(n5701), .ZN(n9098) );
  AND2_X1 U5934 ( .A1(n5700), .A2(n5194), .ZN(n5193) );
  NOR2_X1 U5935 ( .A1(n10719), .A2(n5158), .ZN(n10722) );
  INV_X1 U5936 ( .A(n5159), .ZN(n5158) );
  AOI21_X1 U5937 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n10723), .A(n5160), .ZN(
        n7048) );
  NOR2_X1 U5938 ( .A1(n7061), .A2(n7060), .ZN(n7059) );
  NOR2_X1 U5939 ( .A1(n7059), .A2(n5146), .ZN(n6995) );
  AND2_X1 U5940 ( .A1(n6998), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5146) );
  INV_X1 U5941 ( .A(n5145), .ZN(n7084) );
  AND2_X1 U5942 ( .A1(n5145), .A2(n5144), .ZN(n7088) );
  NAND2_X1 U5943 ( .A1(n7085), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5144) );
  NOR2_X1 U5944 ( .A1(n7376), .A2(n5148), .ZN(n7381) );
  AND2_X1 U5945 ( .A1(n7377), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5148) );
  NOR2_X1 U5946 ( .A1(n7381), .A2(n7380), .ZN(n7793) );
  NAND2_X1 U5947 ( .A1(n9296), .A2(n9297), .ZN(n9300) );
  INV_X1 U5948 ( .A(n5157), .ZN(n9315) );
  AND2_X1 U5949 ( .A1(n5157), .A2(n5156), .ZN(n9317) );
  NAND2_X1 U5950 ( .A1(n9316), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5156) );
  NAND2_X1 U5951 ( .A1(n9345), .A2(n5152), .ZN(n5151) );
  NAND2_X1 U5952 ( .A1(n5153), .A2(n6083), .ZN(n5152) );
  NAND2_X1 U5953 ( .A1(n5186), .A2(n5187), .ZN(n9391) );
  NOR2_X1 U5954 ( .A1(n9433), .A2(n6613), .ZN(n9421) );
  INV_X1 U5955 ( .A(n9448), .ZN(n5617) );
  NAND2_X1 U5956 ( .A1(n9474), .A2(n5640), .ZN(n9460) );
  NAND2_X1 U5957 ( .A1(n9494), .A2(n9071), .ZN(n9476) );
  NAND2_X1 U5958 ( .A1(n6101), .A2(n6100), .ZN(n9641) );
  NAND2_X1 U5959 ( .A1(n5623), .A2(n5620), .ZN(n9541) );
  NOR2_X1 U5960 ( .A1(n9065), .A2(n5628), .ZN(n9543) );
  NAND2_X1 U5961 ( .A1(n8101), .A2(n5305), .ZN(n8442) );
  NAND2_X1 U5962 ( .A1(n5300), .A2(n9565), .ZN(n7993) );
  NAND2_X1 U5963 ( .A1(n10846), .A2(n7944), .ZN(n7946) );
  NAND2_X1 U5964 ( .A1(n7808), .A2(n5179), .ZN(n10846) );
  NOR2_X1 U5965 ( .A1(n7779), .A2(n5180), .ZN(n5179) );
  INV_X1 U5966 ( .A(n7778), .ZN(n5180) );
  NAND2_X1 U5967 ( .A1(n7808), .A2(n7778), .ZN(n7780) );
  AND2_X1 U5968 ( .A1(n9569), .A2(n7777), .ZN(n5630) );
  NAND2_X1 U5969 ( .A1(n5453), .A2(n6579), .ZN(n9558) );
  NAND2_X1 U5970 ( .A1(n7773), .A2(n7772), .ZN(n10782) );
  OR2_X1 U5971 ( .A1(n5722), .A2(n6790), .ZN(n5748) );
  INV_X1 U5972 ( .A(n10752), .ZN(n7728) );
  NAND2_X1 U5973 ( .A1(n7012), .A2(n9701), .ZN(n5708) );
  INV_X1 U5974 ( .A(n9363), .ZN(n9568) );
  NOR2_X1 U5975 ( .A1(n5289), .A2(n10921), .ZN(n5288) );
  AND2_X1 U5976 ( .A1(n9595), .A2(n9594), .ZN(n5167) );
  OR2_X1 U5977 ( .A1(n9596), .A2(n10904), .ZN(n5168) );
  MUX2_X1 U5978 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5690), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5691) );
  NAND2_X1 U5979 ( .A1(n5197), .A2(n5196), .ZN(n5689) );
  CLKBUF_X1 U5980 ( .A(n6365), .Z(n6366) );
  CLKBUF_X1 U5981 ( .A(n6634), .Z(n9091) );
  INV_X1 U5982 ( .A(n6435), .ZN(n8174) );
  INV_X1 U5983 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6831) );
  XNOR2_X1 U5984 ( .A(n5678), .B(n5161), .ZN(n10709) );
  NAND2_X1 U5985 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5161) );
  INV_X1 U5986 ( .A(n7126), .ZN(n8573) );
  NAND2_X1 U5987 ( .A1(n5552), .A2(n9764), .ZN(n9725) );
  NAND2_X1 U5988 ( .A1(n9713), .A2(n5559), .ZN(n5552) );
  NAND2_X1 U5989 ( .A1(n8130), .A2(n8129), .ZN(n8231) );
  NAND2_X1 U5990 ( .A1(n8588), .A2(n8587), .ZN(n10099) );
  NAND2_X1 U5991 ( .A1(n7965), .A2(n7966), .ZN(n7969) );
  NAND2_X1 U5992 ( .A1(n9713), .A2(n5561), .ZN(n9767) );
  NAND2_X1 U5993 ( .A1(n8273), .A2(n8272), .ZN(n8275) );
  INV_X1 U5994 ( .A(n5554), .ZN(n5553) );
  OAI21_X1 U5995 ( .B1(n9723), .B2(n5555), .A(n9721), .ZN(n5554) );
  CLKBUF_X1 U5996 ( .A(n7193), .Z(n7130) );
  OAI21_X1 U5997 ( .B1(n5502), .B2(n7468), .A(n5222), .ZN(n5221) );
  NAND2_X1 U5998 ( .A1(n8708), .A2(n8707), .ZN(n9922) );
  NAND2_X1 U5999 ( .A1(n9697), .A2(n8749), .ZN(n8708) );
  OR2_X1 U6000 ( .A1(n7080), .A2(n7076), .ZN(n9808) );
  NAND2_X1 U6001 ( .A1(n8376), .A2(n8375), .ZN(n8554) );
  OR2_X1 U6002 ( .A1(n6947), .A2(n7417), .ZN(n7131) );
  NAND2_X1 U6003 ( .A1(n5051), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n7101) );
  NAND2_X1 U6004 ( .A1(n5051), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6950) );
  AND2_X1 U6005 ( .A1(n6716), .A2(n6715), .ZN(n6842) );
  OR2_X1 U6006 ( .A1(n6879), .A2(n6878), .ZN(n6876) );
  INV_X1 U6007 ( .A(n6906), .ZN(n10679) );
  AOI21_X1 U6008 ( .B1(n9687), .B2(n8749), .A(n8744), .ZN(n10072) );
  INV_X1 U6009 ( .A(n9893), .ZN(n10077) );
  NAND2_X1 U6010 ( .A1(n5341), .A2(n5340), .ZN(n5339) );
  XNOR2_X1 U6011 ( .A(n5343), .B(n9904), .ZN(n5342) );
  NAND2_X1 U6012 ( .A1(n9942), .A2(n10975), .ZN(n5340) );
  NAND2_X1 U6013 ( .A1(n5563), .A2(n5567), .ZN(n9911) );
  NAND2_X1 U6014 ( .A1(n9947), .A2(n5067), .ZN(n5563) );
  OAI21_X1 U6015 ( .B1(n9947), .B2(n5069), .A(n9116), .ZN(n9932) );
  NAND2_X1 U6016 ( .A1(n10002), .A2(n9111), .ZN(n9978) );
  NAND2_X1 U6017 ( .A1(n9110), .A2(n9109), .ZN(n10004) );
  NAND2_X1 U6018 ( .A1(n5575), .A2(n9108), .ZN(n10008) );
  NAND2_X1 U6019 ( .A1(n10968), .A2(n5595), .ZN(n9106) );
  NOR2_X1 U6020 ( .A1(n5594), .A2(n5593), .ZN(n8469) );
  INV_X1 U6021 ( .A(n8465), .ZN(n5593) );
  NAND2_X1 U6022 ( .A1(n8464), .A2(n8463), .ZN(n10997) );
  NAND2_X1 U6023 ( .A1(n8388), .A2(n8922), .ZN(n8471) );
  AND2_X1 U6024 ( .A1(n7822), .A2(n7821), .ZN(n7898) );
  NAND2_X1 U6025 ( .A1(n5394), .A2(n8865), .ZN(n7863) );
  INV_X1 U6026 ( .A(n10734), .ZN(n10996) );
  OR2_X1 U6027 ( .A1(n7074), .A2(n10580), .ZN(n10741) );
  NAND2_X1 U6029 ( .A1(n6813), .A2(n5261), .ZN(n9063) );
  NAND2_X1 U6030 ( .A1(n5262), .A2(n6810), .ZN(n5261) );
  NAND2_X1 U6031 ( .A1(n6681), .A2(n5263), .ZN(n5262) );
  NAND2_X1 U6032 ( .A1(n6681), .A2(n6680), .ZN(n6812) );
  XNOR2_X1 U6033 ( .A(n6649), .B(n10330), .ZN(n8400) );
  OAI21_X1 U6034 ( .B1(n6930), .B2(n6646), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6649) );
  NAND2_X1 U6035 ( .A1(n6190), .A2(n6189), .ZN(n6210) );
  NAND2_X1 U6036 ( .A1(n6930), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6931) );
  INV_X1 U6037 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6908) );
  INV_X1 U6038 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6872) );
  NAND2_X1 U6039 ( .A1(n5334), .A2(n5781), .ZN(n5802) );
  NAND2_X1 U6040 ( .A1(n5779), .A2(n5778), .ZN(n5334) );
  AOI21_X1 U6041 ( .B1(n5499), .B2(n9248), .A(n5118), .ZN(n5493) );
  INV_X1 U6042 ( .A(n5497), .ZN(n5496) );
  AND2_X1 U6043 ( .A1(n9580), .A2(n9573), .ZN(n9361) );
  AOI21_X1 U6044 ( .B1(n5202), .B2(n5201), .A(n5198), .ZN(n9097) );
  OAI211_X1 U6045 ( .C1(n5545), .C2(n5537), .A(n5536), .B(n5091), .ZN(P1_U3212) );
  NAND2_X1 U6046 ( .A1(n5542), .A2(n9744), .ZN(n5537) );
  INV_X1 U6047 ( .A(n5257), .ZN(n9162) );
  OAI21_X1 U6048 ( .B1(n10081), .B2(n10738), .A(n5258), .ZN(n5257) );
  AOI21_X1 U6049 ( .B1(n10079), .B2(n10068), .A(n9161), .ZN(n5258) );
  AND2_X1 U6050 ( .A1(n5588), .A2(n5581), .ZN(n10086) );
  AOI211_X1 U6051 ( .C1(n10068), .C2(n10084), .A(n9142), .B(n9141), .ZN(n9143)
         );
  NAND2_X1 U6052 ( .A1(n5591), .A2(n5057), .ZN(n5588) );
  INV_X1 U6053 ( .A(n5307), .ZN(n10547) );
  NAND2_X1 U6054 ( .A1(n5586), .A2(n5584), .ZN(n10550) );
  NOR2_X1 U6055 ( .A1(n9136), .A2(n5585), .ZN(n5584) );
  INV_X1 U6056 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n5306) );
  OAI21_X1 U6057 ( .B1(n5586), .B2(n10990), .A(n5582), .ZN(P1_U3519) );
  NAND2_X1 U6058 ( .A1(n5580), .A2(n5579), .ZN(n5582) );
  NAND2_X1 U6059 ( .A1(n5589), .A2(n10990), .ZN(n5579) );
  INV_X2 U6060 ( .A(n5722), .ZN(n5783) );
  AND2_X2 U6061 ( .A1(n7208), .A2(n7111), .ZN(n7104) );
  INV_X1 U6062 ( .A(n7467), .ZN(n5504) );
  NAND2_X1 U6063 ( .A1(n5685), .A2(n5684), .ZN(n5054) );
  NAND2_X1 U6064 ( .A1(n5243), .A2(n8721), .ZN(n10088) );
  NAND2_X1 U6065 ( .A1(n5597), .A2(n6440), .ZN(n7144) );
  INV_X1 U6066 ( .A(n7669), .ZN(n7679) );
  AND2_X1 U6067 ( .A1(n6449), .A2(n6575), .ZN(n7669) );
  OR2_X1 U6068 ( .A1(n10099), .A2(n9953), .ZN(n5055) );
  OAI21_X2 U6069 ( .B1(n7012), .B2(n5709), .A(n5708), .ZN(n10742) );
  AND2_X1 U6070 ( .A1(n8729), .A2(n5547), .ZN(n5056) );
  AND2_X1 U6071 ( .A1(n5590), .A2(n10879), .ZN(n5057) );
  NAND2_X1 U6072 ( .A1(n6078), .A2(n6077), .ZN(n9644) );
  AND2_X1 U6073 ( .A1(n5309), .A2(n5312), .ZN(n5058) );
  AND2_X1 U6074 ( .A1(n5097), .A2(n5170), .ZN(n5059) );
  INV_X1 U6075 ( .A(n9136), .ZN(n5581) );
  AND2_X1 U6076 ( .A1(n5602), .A2(n10936), .ZN(n5060) );
  AND2_X1 U6077 ( .A1(n5314), .A2(n5313), .ZN(n5061) );
  AND2_X1 U6078 ( .A1(n10912), .A2(n5310), .ZN(n5062) );
  INV_X1 U6079 ( .A(n9007), .ZN(n5572) );
  NAND2_X1 U6080 ( .A1(n8080), .A2(n5084), .ZN(n8100) );
  OR2_X1 U6081 ( .A1(n9664), .A2(n9052), .ZN(n6594) );
  INV_X1 U6082 ( .A(n9547), .ZN(n9573) );
  AND2_X1 U6083 ( .A1(n7526), .A2(n7528), .ZN(n8996) );
  OR2_X1 U6084 ( .A1(n10320), .A2(n10321), .ZN(n5063) );
  INV_X1 U6085 ( .A(n10288), .ZN(n5377) );
  OR2_X1 U6086 ( .A1(n5127), .A2(n10291), .ZN(n5064) );
  AND2_X1 U6087 ( .A1(n6675), .A2(n6674), .ZN(n6957) );
  NAND2_X2 U6088 ( .A1(n5703), .A2(n6789), .ZN(n5722) );
  NAND2_X1 U6089 ( .A1(n6412), .A2(n6411), .ZN(n9365) );
  AND3_X1 U6090 ( .A1(n5730), .A2(n5729), .A3(n5728), .ZN(n5065) );
  OR2_X1 U6091 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5066) );
  AND2_X1 U6092 ( .A1(n5055), .A2(n9116), .ZN(n5067) );
  AND2_X1 U6093 ( .A1(n6551), .A2(n6611), .ZN(n9447) );
  AND2_X1 U6094 ( .A1(n8892), .A2(n8891), .ZN(n9002) );
  AND2_X1 U6095 ( .A1(n5277), .A2(n9109), .ZN(n5068) );
  AND2_X1 U6096 ( .A1(n10105), .A2(n9971), .ZN(n5069) );
  AND2_X1 U6097 ( .A1(n7974), .A2(n8120), .ZN(n5070) );
  OR2_X1 U6098 ( .A1(n6817), .A2(n10568), .ZN(n6947) );
  INV_X1 U6099 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6928) );
  AND2_X1 U6100 ( .A1(n9743), .A2(n8535), .ZN(n5071) );
  INV_X1 U6101 ( .A(n9082), .ZN(n9372) );
  XNOR2_X1 U6102 ( .A(n9592), .B(n9393), .ZN(n9082) );
  INV_X1 U6103 ( .A(n9828), .ZN(n7313) );
  NOR2_X1 U6104 ( .A1(n7793), .A2(n5147), .ZN(n5072) );
  NAND2_X1 U6105 ( .A1(n7148), .A2(n10742), .ZN(n6438) );
  NAND2_X1 U6106 ( .A1(n6802), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6681) );
  AND2_X1 U6107 ( .A1(n9014), .A2(n9024), .ZN(n5073) );
  NAND2_X1 U6108 ( .A1(n6173), .A2(n6172), .ZN(n9624) );
  AND2_X1 U6109 ( .A1(n8768), .A2(n5982), .ZN(n5074) );
  AND2_X1 U6110 ( .A1(n6724), .A2(n6643), .ZN(n6690) );
  INV_X1 U6111 ( .A(n7466), .ZN(n5503) );
  INV_X1 U6112 ( .A(n9123), .ZN(n5328) );
  INV_X1 U6113 ( .A(n9006), .ZN(n5266) );
  OR2_X1 U6114 ( .A1(n8358), .A2(n9272), .ZN(n5075) );
  NOR2_X1 U6115 ( .A1(n8498), .A2(n8497), .ZN(n5076) );
  AND2_X1 U6116 ( .A1(n6618), .A2(n6617), .ZN(n9088) );
  NOR2_X1 U6117 ( .A1(n9623), .A2(n9076), .ZN(n5077) );
  AND2_X1 U6118 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n5078) );
  AND2_X1 U6119 ( .A1(n7774), .A2(n7772), .ZN(n5079) );
  NAND2_X1 U6120 ( .A1(n7475), .A2(n7476), .ZN(n5080) );
  NAND2_X1 U6121 ( .A1(n8654), .A2(n8653), .ZN(n10126) );
  INV_X1 U6122 ( .A(n10938), .ZN(n8358) );
  OR2_X1 U6123 ( .A1(n8358), .A2(n8767), .ZN(n5081) );
  INV_X1 U6124 ( .A(n5547), .ZN(n5544) );
  INV_X1 U6125 ( .A(n5317), .ZN(n9151) );
  NOR3_X1 U6126 ( .A1(n5318), .A2(n9933), .A3(n9922), .ZN(n5317) );
  AND2_X1 U6127 ( .A1(n5590), .A2(n5587), .ZN(n5082) );
  NAND2_X1 U6128 ( .A1(n8751), .A2(n8750), .ZN(n10083) );
  AND2_X1 U6129 ( .A1(n5604), .A2(n9089), .ZN(n5083) );
  AND2_X1 U6130 ( .A1(n8082), .A2(n8079), .ZN(n5084) );
  AND2_X1 U6131 ( .A1(n5459), .A2(n9435), .ZN(n5085) );
  INV_X1 U6132 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n10330) );
  NAND2_X1 U6133 ( .A1(n5243), .A2(n5241), .ZN(n9129) );
  NAND2_X1 U6134 ( .A1(n7334), .A2(n7335), .ZN(n5086) );
  AND2_X1 U6135 ( .A1(n6465), .A2(n6585), .ZN(n7779) );
  NAND2_X1 U6136 ( .A1(n6130), .A2(n6129), .ZN(n9634) );
  AND2_X1 U6137 ( .A1(n8915), .A2(n8917), .ZN(n8991) );
  AND2_X1 U6138 ( .A1(n8926), .A2(n8925), .ZN(n9009) );
  OR2_X1 U6139 ( .A1(n9028), .A2(n9016), .ZN(n5087) );
  AND2_X1 U6140 ( .A1(n8941), .A2(n9123), .ZN(n10012) );
  INV_X1 U6141 ( .A(n10012), .ZN(n5330) );
  NOR2_X1 U6142 ( .A1(n10541), .A2(n10978), .ZN(n5088) );
  NOR2_X1 U6143 ( .A1(n10872), .A2(n9821), .ZN(n5089) );
  NOR2_X1 U6144 ( .A1(n8511), .A2(n9818), .ZN(n5090) );
  AND2_X1 U6145 ( .A1(n6587), .A2(n6554), .ZN(n7948) );
  AND2_X1 U6146 ( .A1(n5538), .A2(n5534), .ZN(n5091) );
  AND2_X1 U6147 ( .A1(n10126), .A2(n10040), .ZN(n5092) );
  NAND2_X1 U6148 ( .A1(n6679), .A2(n6678), .ZN(n5093) );
  NOR2_X1 U6149 ( .A1(n9922), .A2(n9942), .ZN(n5094) );
  NOR2_X1 U6150 ( .A1(n10094), .A2(n9738), .ZN(n5095) );
  INV_X1 U6151 ( .A(n5596), .ZN(n5595) );
  NAND2_X1 U6152 ( .A1(n8931), .A2(n8465), .ZN(n5596) );
  AND2_X1 U6153 ( .A1(n9418), .A2(n9432), .ZN(n5096) );
  AND2_X1 U6154 ( .A1(n8820), .A2(n8913), .ZN(n9004) );
  NAND2_X1 U6155 ( .A1(n6616), .A2(n6532), .ZN(n9080) );
  INV_X1 U6156 ( .A(n9080), .ZN(n5143) );
  AND2_X1 U6157 ( .A1(n9072), .A2(n5640), .ZN(n5097) );
  INV_X1 U6158 ( .A(n5609), .ZN(n5607) );
  NAND2_X1 U6159 ( .A1(n9390), .A2(n9375), .ZN(n5609) );
  AND2_X1 U6160 ( .A1(n5512), .A2(n5510), .ZN(n5098) );
  NAND2_X1 U6161 ( .A1(n5457), .A2(n6614), .ZN(n5099) );
  AND2_X1 U6162 ( .A1(n5391), .A2(n9129), .ZN(n5100) );
  NAND2_X1 U6163 ( .A1(n5568), .A2(n9117), .ZN(n5101) );
  INV_X1 U6164 ( .A(n5511), .ZN(n5510) );
  NAND2_X1 U6165 ( .A1(n5513), .A2(n8635), .ZN(n5511) );
  INV_X1 U6166 ( .A(n10085), .ZN(n5585) );
  AND2_X1 U6167 ( .A1(n7526), .A2(n7525), .ZN(n5102) );
  AND2_X1 U6168 ( .A1(n5606), .A2(n9088), .ZN(n5103) );
  AND2_X1 U6169 ( .A1(n9062), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5104) );
  NAND2_X1 U6170 ( .A1(n8221), .A2(n8220), .ZN(n5105) );
  NAND2_X1 U6171 ( .A1(n5541), .A2(n9744), .ZN(n5106) );
  AND2_X1 U6172 ( .A1(n8135), .A2(n8132), .ZN(n5107) );
  AND2_X1 U6173 ( .A1(n5283), .A2(n10330), .ZN(n5108) );
  INV_X1 U6174 ( .A(n5543), .ZN(n5542) );
  NAND2_X1 U6175 ( .A1(n5546), .A2(n5544), .ZN(n5543) );
  NAND2_X1 U6176 ( .A1(n6038), .A2(n6037), .ZN(n9655) );
  AND2_X1 U6177 ( .A1(n5456), .A2(n5459), .ZN(n5109) );
  INV_X1 U6178 ( .A(n7509), .ZN(n8638) );
  BUF_X1 U6179 ( .A(n7183), .Z(n7509) );
  XNOR2_X1 U6180 ( .A(n6671), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8985) );
  INV_X1 U6181 ( .A(n8985), .ZN(n5509) );
  INV_X1 U6182 ( .A(n6682), .ZN(n5284) );
  AND2_X1 U6183 ( .A1(n5464), .A2(n6594), .ZN(n5110) );
  AND3_X1 U6184 ( .A1(n8534), .A2(n8544), .A3(n8535), .ZN(n5111) );
  NAND2_X1 U6185 ( .A1(n9110), .A2(n5068), .ZN(n10002) );
  AND2_X1 U6186 ( .A1(n10032), .A2(n8752), .ZN(n5112) );
  AND2_X1 U6187 ( .A1(n8101), .A2(n5303), .ZN(n5113) );
  BUF_X1 U6188 ( .A(n5697), .Z(n6369) );
  XNOR2_X1 U6189 ( .A(n6006), .B(SI_14_), .ZN(n6005) );
  NAND2_X1 U6190 ( .A1(n8290), .A2(n8241), .ZN(n8377) );
  NAND2_X1 U6191 ( .A1(n9542), .A2(n5625), .ZN(n5624) );
  INV_X1 U6192 ( .A(n5624), .ZN(n5620) );
  NAND2_X1 U6193 ( .A1(n8602), .A2(n8601), .ZN(n10109) );
  INV_X1 U6194 ( .A(n10109), .ZN(n5313) );
  NAND2_X1 U6195 ( .A1(n5280), .A2(n5570), .ZN(n8378) );
  NAND2_X1 U6196 ( .A1(n5512), .A2(n5513), .ZN(n5114) );
  NAND2_X1 U6197 ( .A1(n5477), .A2(n6158), .ZN(n9225) );
  NAND2_X1 U6198 ( .A1(n6160), .A2(SI_21_), .ZN(n5115) );
  AND2_X1 U6199 ( .A1(n9121), .A2(n9120), .ZN(n5116) );
  NAND2_X1 U6200 ( .A1(n9435), .A2(n5616), .ZN(n5615) );
  INV_X1 U6201 ( .A(n5615), .ZN(n5611) );
  AND2_X1 U6202 ( .A1(n6086), .A2(n6085), .ZN(n9539) );
  INV_X1 U6203 ( .A(n5216), .ZN(n5215) );
  NAND2_X1 U6204 ( .A1(n6027), .A2(n5217), .ZN(n5216) );
  AND2_X1 U6205 ( .A1(n6275), .A2(n6274), .ZN(n5117) );
  INV_X1 U6206 ( .A(n5614), .ZN(n9623) );
  NAND2_X1 U6207 ( .A1(n5617), .A2(n9443), .ZN(n5614) );
  INV_X1 U6208 ( .A(n5428), .ZN(n5427) );
  NAND2_X1 U6209 ( .A1(n6096), .A2(n5429), .ZN(n5428) );
  NAND2_X1 U6210 ( .A1(n6377), .A2(n6376), .ZN(n5118) );
  NAND2_X1 U6211 ( .A1(n6030), .A2(n6052), .ZN(n5119) );
  NAND2_X1 U6212 ( .A1(n5966), .A2(n5943), .ZN(n5944) );
  NAND2_X1 U6213 ( .A1(n7533), .A2(n10741), .ZN(n10022) );
  INV_X1 U6214 ( .A(n8557), .ZN(n5475) );
  INV_X1 U6215 ( .A(n9099), .ZN(n9248) );
  NAND2_X1 U6216 ( .A1(n8100), .A2(n8099), .ZN(n8357) );
  OAI21_X1 U6217 ( .B1(n7918), .B2(n5070), .A(n5273), .ZN(n8014) );
  NAND2_X1 U6218 ( .A1(n6013), .A2(n6012), .ZN(n9659) );
  INV_X1 U6219 ( .A(n9659), .ZN(n5304) );
  NAND2_X1 U6220 ( .A1(n8237), .A2(n8236), .ZN(n10928) );
  INV_X1 U6221 ( .A(n10928), .ZN(n5312) );
  OR2_X1 U6222 ( .A1(n10993), .A2(n5306), .ZN(n5120) );
  INV_X1 U6223 ( .A(n9742), .ZN(n5514) );
  INV_X1 U6224 ( .A(n5221), .ZN(n7479) );
  NAND2_X1 U6225 ( .A1(n8018), .A2(n8017), .ZN(n8170) );
  NAND2_X1 U6226 ( .A1(n5520), .A2(n5518), .ZN(n7964) );
  INV_X1 U6227 ( .A(n9744), .ZN(n5540) );
  AND2_X1 U6228 ( .A1(n10196), .A2(n10195), .ZN(n5121) );
  NAND2_X1 U6229 ( .A1(n6655), .A2(n6654), .ZN(n5122) );
  AND2_X1 U6230 ( .A1(n6383), .A2(n10153), .ZN(n5123) );
  AND2_X1 U6231 ( .A1(n7947), .A2(n6587), .ZN(n5124) );
  AND2_X1 U6232 ( .A1(n8080), .A2(n8079), .ZN(n5125) );
  AND2_X1 U6233 ( .A1(n7490), .A2(n7445), .ZN(n5126) );
  XNOR2_X1 U6234 ( .A(n6681), .B(n6803), .ZN(n6751) );
  NAND2_X1 U6235 ( .A1(n5903), .A2(n5902), .ZN(n8029) );
  INV_X1 U6236 ( .A(n8029), .ZN(n5299) );
  NAND2_X1 U6237 ( .A1(n7169), .A2(n10875), .ZN(n5587) );
  INV_X1 U6238 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5141) );
  NAND2_X1 U6239 ( .A1(n7921), .A2(n7920), .ZN(n10872) );
  INV_X1 U6240 ( .A(n10872), .ZN(n5310) );
  NAND4_X1 U6241 ( .A1(n5696), .A2(n5695), .A3(n5694), .A4(n5693), .ZN(n6436)
         );
  NAND2_X1 U6242 ( .A1(n5881), .A2(n5880), .ZN(n10863) );
  INV_X1 U6243 ( .A(n10863), .ZN(n5301) );
  AOI21_X1 U6244 ( .B1(n7773), .B2(n5079), .A(n5177), .ZN(n9570) );
  OR2_X1 U6245 ( .A1(n5377), .A2(n10284), .ZN(n5127) );
  NAND2_X1 U6246 ( .A1(n10283), .A2(n10282), .ZN(n5128) );
  NAND3_X1 U6247 ( .A1(n10297), .A2(n10296), .A3(n10295), .ZN(n5129) );
  INV_X1 U6248 ( .A(n9347), .ZN(n5153) );
  AND4_X1 U6249 ( .A1(n10329), .A2(n10328), .A3(n10327), .A4(n10326), .ZN(
        n5130) );
  XOR2_X1 U6250 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_242), .Z(n5131) );
  NAND2_X1 U6251 ( .A1(n10334), .A2(n10335), .ZN(n5132) );
  NAND2_X1 U6252 ( .A1(n10332), .A2(n10331), .ZN(n5133) );
  OR2_X1 U6253 ( .A1(keyinput_217), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n5134)
         );
  AND2_X1 U6254 ( .A1(n6629), .A2(n10800), .ZN(n5135) );
  NOR2_X1 U6255 ( .A1(n7664), .A2(n9538), .ZN(n5201) );
  INV_X1 U6256 ( .A(n7664), .ZN(n5200) );
  AOI21_X1 U6257 ( .B1(n5202), .B2(n10794), .A(n9095), .ZN(n9589) );
  NOR2_X4 U6258 ( .A1(n7665), .A2(n6635), .ZN(n6542) );
  NAND2_X1 U6259 ( .A1(n5142), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6288) );
  OAI21_X1 U6260 ( .B1(n5443), .B2(n5442), .A(n6618), .ZN(n6621) );
  NOR2_X2 U6261 ( .A1(n9371), .A2(n9372), .ZN(n9370) );
  NAND2_X1 U6262 ( .A1(n5149), .A2(n9357), .ZN(P2_U3264) );
  NAND2_X1 U6263 ( .A1(n5150), .A2(n10696), .ZN(n5149) );
  XNOR2_X1 U6264 ( .A(n5151), .B(n9346), .ZN(n5150) );
  NAND2_X1 U6265 ( .A1(n9340), .A2(n9341), .ZN(n9345) );
  AOI21_X1 U6266 ( .B1(n10720), .B2(n10721), .A(n5160), .ZN(n5159) );
  NOR2_X1 U6267 ( .A1(n10721), .A2(n10720), .ZN(n5160) );
  NAND2_X1 U6268 ( .A1(n5168), .A2(n5167), .ZN(n9672) );
  NAND3_X1 U6269 ( .A1(n5598), .A2(n7750), .A3(n5178), .ZN(n7773) );
  AND3_X2 U6270 ( .A1(n5725), .A2(n5724), .A3(n5726), .ZN(n10752) );
  OAI21_X2 U6271 ( .B1(n9536), .B2(n9542), .A(n6603), .ZN(n9526) );
  NAND2_X2 U6272 ( .A1(n5467), .A2(n5465), .ZN(n5464) );
  OR2_X2 U6273 ( .A1(n8092), .A2(n8098), .ZN(n5467) );
  NAND2_X1 U6274 ( .A1(n5186), .A2(n5184), .ZN(n5185) );
  OR2_X2 U6275 ( .A1(n9444), .A2(n5189), .ZN(n5186) );
  INV_X1 U6276 ( .A(n9434), .ZN(n5460) );
  NAND2_X1 U6277 ( .A1(n9694), .A2(n5104), .ZN(n5194) );
  NAND2_X1 U6278 ( .A1(n5197), .A2(n5195), .ZN(n5688) );
  NOR2_X1 U6279 ( .A1(n6055), .A2(n5673), .ZN(n5686) );
  NAND2_X1 U6280 ( .A1(n5743), .A2(n5744), .ZN(n5204) );
  NAND2_X1 U6281 ( .A1(n5717), .A2(n5716), .ZN(n5205) );
  NAND2_X1 U6282 ( .A1(n5823), .A2(n5822), .ZN(n5826) );
  NAND2_X1 U6283 ( .A1(n5331), .A2(n5207), .ZN(n5206) );
  NAND2_X1 U6284 ( .A1(n5759), .A2(n5333), .ZN(n5207) );
  NAND2_X1 U6285 ( .A1(n8110), .A2(n8109), .ZN(n8115) );
  NAND2_X2 U6286 ( .A1(n5208), .A2(n7965), .ZN(n8110) );
  NAND2_X1 U6287 ( .A1(n6009), .A2(n6008), .ZN(n5212) );
  NAND2_X1 U6288 ( .A1(n5222), .A2(n7468), .ZN(n5219) );
  NAND3_X1 U6289 ( .A1(n5220), .A2(n5219), .A3(n5080), .ZN(n7691) );
  INV_X1 U6290 ( .A(n8543), .ZN(n5224) );
  NAND2_X1 U6291 ( .A1(n8543), .A2(n8546), .ZN(n8534) );
  OAI211_X1 U6292 ( .C1(n5227), .C2(n5224), .A(n5225), .B(n5223), .ZN(n9786)
         );
  NAND3_X1 U6293 ( .A1(n8533), .A2(n8532), .A3(n5228), .ZN(n5223) );
  NAND2_X2 U6294 ( .A1(n8533), .A2(n8532), .ZN(n8544) );
  NAND2_X1 U6295 ( .A1(n6143), .A2(n5232), .ZN(n5231) );
  NAND2_X1 U6296 ( .A1(n5231), .A2(n5115), .ZN(n6162) );
  OAI21_X1 U6297 ( .B1(n6240), .B2(n5236), .A(n5233), .ZN(n6283) );
  INV_X1 U6298 ( .A(n5720), .ZN(n5680) );
  NAND2_X4 U6299 ( .A1(n5249), .A2(n5248), .ZN(n5720) );
  NAND3_X1 U6300 ( .A1(n5706), .A2(n5246), .A3(n5244), .ZN(n5718) );
  NAND2_X1 U6301 ( .A1(n5245), .A2(n5078), .ZN(n5244) );
  INV_X1 U6302 ( .A(n5248), .ZN(n5245) );
  NAND2_X1 U6303 ( .A1(n5247), .A2(n5078), .ZN(n5246) );
  INV_X1 U6304 ( .A(n5249), .ZN(n5247) );
  NAND3_X1 U6305 ( .A1(n5249), .A2(n5248), .A3(n5679), .ZN(n5706) );
  NAND3_X1 U6306 ( .A1(n8159), .A2(n5105), .A3(n8158), .ZN(n5251) );
  NAND3_X1 U6307 ( .A1(n5393), .A2(n9128), .A3(n9939), .ZN(n5256) );
  NAND2_X1 U6308 ( .A1(n7918), .A2(n5268), .ZN(n5267) );
  OAI21_X1 U6309 ( .B1(n7918), .B2(n5270), .A(n5268), .ZN(n8131) );
  AOI21_X1 U6310 ( .B1(n5268), .B2(n5270), .A(n5266), .ZN(n5265) );
  NAND2_X1 U6311 ( .A1(n5284), .A2(n5053), .ZN(n6930) );
  OAI211_X1 U6312 ( .C1(n10082), .C2(n10539), .A(n10080), .B(n10081), .ZN(
        n10549) );
  NAND2_X1 U6313 ( .A1(n9364), .A2(n5294), .ZN(n5291) );
  NAND3_X1 U6314 ( .A1(n5291), .A2(n5290), .A3(n5292), .ZN(n9578) );
  NAND3_X1 U6315 ( .A1(n5291), .A2(n5290), .A3(n5288), .ZN(n5295) );
  NAND2_X1 U6316 ( .A1(n9364), .A2(n9586), .ZN(n9582) );
  NAND2_X1 U6317 ( .A1(n5295), .A2(n9581), .ZN(n9669) );
  OAI21_X1 U6318 ( .B1(n5307), .B2(n10990), .A(n5120), .ZN(P1_U3522) );
  OAI21_X1 U6319 ( .B1(n10072), .B2(n10984), .A(n10075), .ZN(n5308) );
  NAND2_X1 U6320 ( .A1(n10038), .A2(n9122), .ZN(n10011) );
  NAND2_X1 U6321 ( .A1(n5759), .A2(n5758), .ZN(n5779) );
  NAND2_X1 U6322 ( .A1(n5355), .A2(n5356), .ZN(n10344) );
  NAND2_X1 U6323 ( .A1(n10323), .A2(n5357), .ZN(n5355) );
  NAND2_X1 U6324 ( .A1(n10285), .A2(n5371), .ZN(n5369) );
  NAND2_X1 U6325 ( .A1(n5369), .A2(n5370), .ZN(n10307) );
  NAND3_X1 U6326 ( .A1(n10292), .A2(n5134), .A3(n5376), .ZN(n5375) );
  AOI21_X1 U6327 ( .B1(n10344), .B2(n10343), .A(n10342), .ZN(n10346) );
  AOI21_X1 U6328 ( .B1(n10349), .B2(keyinput_255), .A(keyinput_127), .ZN(
        n10528) );
  OAI22_X1 U6329 ( .A1(n10207), .A2(n10206), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(keyinput_170), .ZN(n10208) );
  INV_X1 U6330 ( .A(n5443), .ZN(n9090) );
  NAND2_X1 U6331 ( .A1(n5917), .A2(n5411), .ZN(n5410) );
  INV_X1 U6332 ( .A(n9120), .ZN(n5397) );
  NAND2_X1 U6333 ( .A1(n5983), .A2(n5635), .ZN(n5985) );
  NAND2_X1 U6334 ( .A1(n9939), .A2(n9128), .ZN(n9913) );
  NAND2_X1 U6335 ( .A1(n5430), .A2(n6096), .ZN(n6118) );
  NAND2_X1 U6336 ( .A1(n5967), .A2(n5966), .ZN(n5983) );
  NAND2_X1 U6337 ( .A1(n8013), .A2(n8902), .ZN(n5389) );
  NAND2_X1 U6338 ( .A1(n7933), .A2(n8898), .ZN(n7935) );
  NAND2_X1 U6339 ( .A1(n8881), .A2(n7528), .ZN(n5395) );
  NAND3_X1 U6340 ( .A1(n5394), .A2(n8865), .A3(n8888), .ZN(n9020) );
  OR2_X1 U6341 ( .A1(n8139), .A2(n5401), .ZN(n5400) );
  NAND2_X1 U6342 ( .A1(n5400), .A2(n5398), .ZN(n8254) );
  INV_X1 U6343 ( .A(n7166), .ZN(n5403) );
  NAND2_X1 U6344 ( .A1(n8851), .A2(n7278), .ZN(n7163) );
  NAND3_X1 U6345 ( .A1(n5403), .A2(n8851), .A3(n7278), .ZN(n7279) );
  NAND2_X1 U6346 ( .A1(n7269), .A2(n9829), .ZN(n8851) );
  NAND2_X1 U6347 ( .A1(n5410), .A2(n5408), .ZN(n5967) );
  NAND2_X1 U6348 ( .A1(n5917), .A2(n5916), .ZN(n5939) );
  NAND2_X1 U6349 ( .A1(n6168), .A2(n6167), .ZN(n6190) );
  NAND4_X1 U6350 ( .A1(n5448), .A2(n5422), .A3(n5447), .A4(n5419), .ZN(n5446)
         );
  NAND3_X1 U6351 ( .A1(n5420), .A2(n8063), .A3(n6573), .ZN(n5419) );
  NAND2_X1 U6352 ( .A1(n6094), .A2(n6093), .ZN(n5430) );
  NAND2_X1 U6353 ( .A1(n6283), .A2(n5434), .ZN(n5433) );
  NAND2_X1 U6354 ( .A1(n6283), .A2(n6282), .ZN(n6315) );
  AND2_X1 U6355 ( .A1(n5648), .A2(n5647), .ZN(n5763) );
  AND2_X1 U6356 ( .A1(n5438), .A2(n5441), .ZN(n5650) );
  NOR2_X1 U6357 ( .A1(n5491), .A2(n5490), .ZN(n5438) );
  NAND4_X2 U6358 ( .A1(n5440), .A2(n5439), .A3(n5784), .A4(n5441), .ZN(n6055)
         );
  AND3_X2 U6359 ( .A1(n5648), .A2(n5647), .A3(n5649), .ZN(n5784) );
  AND2_X1 U6360 ( .A1(n5645), .A2(n5644), .ZN(n5441) );
  NAND2_X1 U6361 ( .A1(n8034), .A2(n8035), .ZN(n6591) );
  NAND3_X1 U6362 ( .A1(n7947), .A2(n6588), .A3(n6587), .ZN(n7985) );
  NAND2_X1 U6363 ( .A1(n5445), .A2(n6638), .ZN(P2_U3244) );
  NAND2_X1 U6364 ( .A1(n5446), .A2(n6633), .ZN(n5445) );
  NAND2_X1 U6365 ( .A1(n6632), .A2(n6631), .ZN(n5447) );
  NAND2_X1 U6366 ( .A1(n5449), .A2(n5135), .ZN(n5448) );
  INV_X1 U6367 ( .A(n6632), .ZN(n5449) );
  NAND3_X1 U6368 ( .A1(n5451), .A2(n6582), .A3(n5450), .ZN(n7803) );
  NAND3_X1 U6369 ( .A1(n7742), .A2(n6581), .A3(n5455), .ZN(n5451) );
  NAND2_X1 U6370 ( .A1(n7742), .A2(n6577), .ZN(n10788) );
  INV_X1 U6371 ( .A(n6615), .ZN(n5456) );
  INV_X1 U6372 ( .A(n6613), .ZN(n5459) );
  OAI21_X1 U6373 ( .B1(n5460), .B2(n6613), .A(n5458), .ZN(n5461) );
  INV_X1 U6374 ( .A(n5461), .ZN(n9419) );
  NAND2_X1 U6375 ( .A1(n5467), .A2(n5075), .ZN(n8363) );
  INV_X1 U6376 ( .A(n5464), .ZN(n8362) );
  INV_X1 U6377 ( .A(n5075), .ZN(n5466) );
  NAND2_X1 U6378 ( .A1(n8561), .A2(n5473), .ZN(n5469) );
  NAND2_X1 U6379 ( .A1(n5470), .A2(n5469), .ZN(n8759) );
  NAND2_X1 U6380 ( .A1(n9196), .A2(n5481), .ZN(n5479) );
  NAND2_X1 U6381 ( .A1(n7570), .A2(n5484), .ZN(n9217) );
  NAND2_X1 U6382 ( .A1(n5732), .A2(n7567), .ZN(n7570) );
  NAND2_X1 U6383 ( .A1(n8197), .A2(n5485), .ZN(n8406) );
  NAND2_X1 U6384 ( .A1(n8406), .A2(n6069), .ZN(n6087) );
  NAND2_X1 U6385 ( .A1(n7588), .A2(n5486), .ZN(n7643) );
  NAND2_X1 U6386 ( .A1(n7643), .A2(n5842), .ZN(n5867) );
  NAND2_X1 U6387 ( .A1(n7844), .A2(n5914), .ZN(n5489) );
  NAND3_X1 U6388 ( .A1(n5646), .A2(n5948), .A3(n5990), .ZN(n5490) );
  NAND3_X1 U6389 ( .A1(n5643), .A2(n5642), .A3(n5949), .ZN(n5491) );
  NAND2_X1 U6390 ( .A1(n6313), .A2(n5494), .ZN(n5492) );
  OAI211_X1 U6391 ( .C1(n6313), .C2(n5496), .A(n5492), .B(n5493), .ZN(P2_U3222) );
  NAND2_X1 U6392 ( .A1(n5501), .A2(n7124), .ZN(n8570) );
  NAND2_X1 U6393 ( .A1(n6963), .A2(n7122), .ZN(n5501) );
  OAI21_X1 U6394 ( .B1(n6963), .B2(n7122), .A(n5501), .ZN(n7081) );
  NAND2_X1 U6395 ( .A1(n5505), .A2(n7338), .ZN(n7468) );
  NAND3_X1 U6396 ( .A1(n7242), .A2(n7241), .A3(n5086), .ZN(n5505) );
  NAND2_X1 U6397 ( .A1(n7242), .A2(n7241), .ZN(n7339) );
  NAND2_X1 U6398 ( .A1(n8159), .A2(n8158), .ZN(n5507) );
  XNOR2_X1 U6399 ( .A(n5507), .B(n8164), .ZN(n8172) );
  INV_X1 U6400 ( .A(n8795), .ZN(n8716) );
  AND2_X4 U6401 ( .A1(n7415), .A2(n7208), .ZN(n8795) );
  NAND2_X1 U6402 ( .A1(n8110), .A2(n5515), .ZN(n8157) );
  NAND2_X1 U6403 ( .A1(n7691), .A2(n5521), .ZN(n5520) );
  NAND2_X1 U6404 ( .A1(n7691), .A2(n7690), .ZN(n7692) );
  INV_X1 U6405 ( .A(n5533), .ZN(n5529) );
  NAND2_X1 U6406 ( .A1(n8499), .A2(n5532), .ZN(n5530) );
  AND2_X1 U6407 ( .A1(n5532), .A2(n8516), .ZN(n5531) );
  OR2_X1 U6408 ( .A1(n8498), .A2(n8497), .ZN(n5532) );
  AND2_X1 U6409 ( .A1(n8498), .A2(n8497), .ZN(n5533) );
  AOI21_X1 U6410 ( .B1(n5545), .B2(n5548), .A(n5543), .ZN(n8808) );
  OR2_X2 U6411 ( .A1(n9803), .A2(n5106), .ZN(n5536) );
  INV_X1 U6412 ( .A(n8729), .ZN(n5546) );
  NOR2_X1 U6413 ( .A1(n8719), .A2(n8720), .ZN(n5547) );
  NAND3_X1 U6414 ( .A1(n9790), .A2(n9787), .A3(n5550), .ZN(n5549) );
  NAND2_X1 U6415 ( .A1(n5549), .A2(n5553), .ZN(n9778) );
  NAND3_X1 U6416 ( .A1(n9790), .A2(n9787), .A3(n9714), .ZN(n9713) );
  NAND3_X1 U6417 ( .A1(n7490), .A2(n7446), .A3(n7445), .ZN(n7552) );
  NAND2_X1 U6418 ( .A1(n8133), .A2(n5107), .ZN(n8233) );
  NAND2_X1 U6419 ( .A1(n8133), .A2(n8132), .ZN(n8134) );
  NAND2_X1 U6420 ( .A1(n5575), .A2(n5573), .ZN(n9110) );
  NAND2_X1 U6421 ( .A1(n10030), .A2(n9107), .ZN(n5575) );
  NAND2_X1 U6422 ( .A1(n7856), .A2(n5576), .ZN(n7884) );
  NAND2_X1 U6423 ( .A1(n5578), .A2(n5108), .ZN(n6677) );
  NAND3_X1 U6424 ( .A1(n5581), .A2(n5589), .A3(n10085), .ZN(n5580) );
  NAND3_X1 U6425 ( .A1(n7748), .A2(n7678), .A3(n7717), .ZN(n5598) );
  NAND2_X1 U6426 ( .A1(n5650), .A2(n5784), .ZN(n6035) );
  NAND2_X1 U6427 ( .A1(n9384), .A2(n5103), .ZN(n5599) );
  NAND3_X1 U6428 ( .A1(n5608), .A2(n9588), .A3(n9589), .ZN(n9671) );
  NAND3_X1 U6429 ( .A1(n5600), .A2(n5602), .A3(n5599), .ZN(n9590) );
  NAND3_X1 U6430 ( .A1(n5600), .A2(n5060), .A3(n5599), .ZN(n5608) );
  NAND2_X1 U6431 ( .A1(n9448), .A2(n5611), .ZN(n5610) );
  NAND2_X1 U6432 ( .A1(n10846), .A2(n5618), .ZN(n7982) );
  INV_X1 U6433 ( .A(n8423), .ZN(n5627) );
  AND2_X1 U6434 ( .A1(n9655), .A2(n9269), .ZN(n5628) );
  OAI21_X1 U6435 ( .B1(n7809), .B2(n5630), .A(n7808), .ZN(n10834) );
  AND4_X1 U6436 ( .A1(n7161), .A2(n7160), .A3(n7159), .A4(n7158), .ZN(n7280)
         );
  INV_X1 U6437 ( .A(n10568), .ZN(n6814) );
  NAND2_X1 U6438 ( .A1(n10568), .A2(n6817), .ZN(n6948) );
  NAND3_X1 U6439 ( .A1(n6693), .A2(n6644), .A3(n6690), .ZN(n6682) );
  NAND2_X1 U6440 ( .A1(n5686), .A2(n5684), .ZN(n5674) );
  NAND2_X1 U6441 ( .A1(n5052), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7102) );
  CLKBUF_X1 U6442 ( .A(n8782), .Z(n9216) );
  CLKBUF_X1 U6443 ( .A(n7602), .Z(n7645) );
  CLKBUF_X1 U6444 ( .A(n8759), .Z(n9056) );
  XNOR2_X1 U6445 ( .A(n9911), .B(n9914), .ZN(n10093) );
  AOI21_X1 U6446 ( .B1(n9705), .B2(n9703), .A(n9702), .ZN(n9755) );
  OR2_X1 U6447 ( .A1(n7113), .A2(n10676), .ZN(n5631) );
  OR2_X1 U6448 ( .A1(n7208), .A2(n10655), .ZN(n5632) );
  INV_X1 U6449 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6653) );
  OR2_X1 U6450 ( .A1(n9592), .A2(n5042), .ZN(n5633) );
  INV_X1 U6451 ( .A(n6573), .ZN(n5698) );
  AND2_X1 U6452 ( .A1(n6251), .A2(n6250), .ZN(n9437) );
  INV_X1 U6453 ( .A(n9437), .ZN(n9078) );
  AND2_X1 U6454 ( .A1(n5984), .A2(n5971), .ZN(n5635) );
  AND2_X1 U6455 ( .A1(n5916), .A2(n5899), .ZN(n5636) );
  NAND2_X1 U6456 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n5637) );
  INV_X1 U6457 ( .A(n9694), .ZN(n9695) );
  AND2_X1 U6458 ( .A1(n6959), .A2(n6958), .ZN(n5638) );
  INV_X1 U6459 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5709) );
  OR2_X1 U6460 ( .A1(n7012), .A2(n10709), .ZN(n5639) );
  NAND2_X1 U6461 ( .A1(n7659), .A2(n9549), .ZN(n10803) );
  OR2_X1 U6462 ( .A1(n7291), .A2(n7156), .ZN(n10945) );
  INV_X1 U6463 ( .A(n9002), .ZN(n7857) );
  INV_X1 U6464 ( .A(n9608), .ZN(n9418) );
  INV_X1 U6465 ( .A(n9624), .ZN(n9074) );
  INV_X1 U6466 ( .A(n8354), .ZN(n6633) );
  OR2_X1 U6467 ( .A1(n9132), .A2(n9131), .ZN(n5641) );
  OAI22_X1 U6468 ( .A1(n10172), .A2(keyinput_141), .B1(n10171), .B2(SI_19_), 
        .ZN(n10173) );
  INV_X1 U6469 ( .A(n10173), .ZN(n10174) );
  XNOR2_X1 U6470 ( .A(keyinput_161), .B(P2_RD_REG_SCAN_IN), .ZN(n10203) );
  OR2_X1 U6471 ( .A1(n10204), .A2(n10203), .ZN(n10205) );
  INV_X1 U6472 ( .A(keyinput_181), .ZN(n10222) );
  XNOR2_X1 U6473 ( .A(n10222), .B(P2_REG3_REG_9__SCAN_IN), .ZN(n10223) );
  OAI22_X1 U6474 ( .A1(n10228), .A2(keyinput_183), .B1(n10227), .B2(
        P2_REG3_REG_20__SCAN_IN), .ZN(n10229) );
  OAI22_X1 U6475 ( .A1(n10233), .A2(keyinput_185), .B1(n10232), .B2(
        P2_REG3_REG_22__SCAN_IN), .ZN(n10234) );
  INV_X1 U6476 ( .A(n10234), .ZN(n10235) );
  NAND2_X1 U6477 ( .A1(n10236), .A2(n10235), .ZN(n10242) );
  OAI22_X1 U6478 ( .A1(n10576), .A2(keyinput_198), .B1(n10255), .B2(
        P2_DATAO_REG_26__SCAN_IN), .ZN(n10256) );
  INV_X1 U6479 ( .A(n10256), .ZN(n10257) );
  NAND2_X1 U6480 ( .A1(n10258), .A2(n10257), .ZN(n10259) );
  XNOR2_X1 U6481 ( .A(keyinput_203), .B(P2_DATAO_REG_21__SCAN_IN), .ZN(n10267)
         );
  AOI21_X1 U6482 ( .B1(n10269), .B2(n10268), .A(n10267), .ZN(n10270) );
  INV_X1 U6483 ( .A(n10270), .ZN(n10276) );
  INV_X1 U6484 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6645) );
  OR2_X1 U6485 ( .A1(n9360), .A2(n8174), .ZN(n6619) );
  NAND2_X1 U6486 ( .A1(keyinput_251), .A2(P1_D_REG_0__SCAN_IN), .ZN(n10340) );
  INV_X1 U6487 ( .A(n7983), .ZN(n6588) );
  INV_X1 U6488 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5649) );
  NAND2_X1 U6489 ( .A1(n10341), .A2(n10340), .ZN(n10342) );
  INV_X1 U6490 ( .A(n8991), .ZN(n8239) );
  INV_X1 U6491 ( .A(n6624), .ZN(n6625) );
  NAND2_X1 U6492 ( .A1(n6014), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6040) );
  INV_X1 U6493 ( .A(n9485), .ZN(n9073) );
  INV_X1 U6494 ( .A(n8081), .ZN(n8082) );
  NAND2_X1 U6495 ( .A1(n6436), .A2(n7674), .ZN(n6440) );
  INV_X1 U6496 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5651) );
  NOR2_X1 U6497 ( .A1(n7925), .A2(n6815), .ZN(n6846) );
  INV_X1 U6498 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7517) );
  NOR2_X1 U6499 ( .A1(n8257), .A2(n8256), .ZN(n8255) );
  INV_X1 U6500 ( .A(n9004), .ZN(n8135) );
  INV_X1 U6501 ( .A(n8996), .ZN(n7446) );
  INV_X1 U6502 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6809) );
  INV_X1 U6503 ( .A(n5843), .ZN(n5844) );
  OR2_X1 U6504 ( .A1(n6196), .A2(n10141), .ZN(n6215) );
  INV_X1 U6505 ( .A(n9228), .ZN(n6187) );
  NAND2_X1 U6506 ( .A1(n8063), .A2(n9546), .ZN(n6354) );
  OR2_X1 U6507 ( .A1(n6288), .A2(n9165), .ZN(n6301) );
  INV_X1 U6508 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10140) );
  INV_X1 U6509 ( .A(n9510), .ZN(n9070) );
  INV_X1 U6510 ( .A(n10613), .ZN(n6346) );
  NAND2_X1 U6511 ( .A1(n9831), .A2(n5040), .ZN(n6962) );
  OR2_X1 U6512 ( .A1(n8472), .A2(n9792), .ZN(n8615) );
  AND2_X1 U6513 ( .A1(n8613), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n8666) );
  AND2_X1 U6514 ( .A1(n10972), .A2(n8930), .ZN(n10058) );
  INV_X1 U6515 ( .A(n8886), .ZN(n7448) );
  NAND2_X1 U6516 ( .A1(n6809), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6810) );
  NAND2_X1 U6517 ( .A1(n5897), .A2(n10144), .ZN(n5916) );
  NAND2_X1 U6518 ( .A1(n5850), .A2(n5849), .ZN(n5868) );
  INV_X1 U6519 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5761) );
  INV_X1 U6520 ( .A(n7592), .ZN(n5841) );
  INV_X1 U6521 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7650) );
  OR2_X1 U6522 ( .A1(n6215), .A2(n10219), .ZN(n6244) );
  NAND2_X1 U6523 ( .A1(n5882), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5904) );
  NAND2_X1 U6524 ( .A1(n5924), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5955) );
  OR2_X1 U6525 ( .A1(n6371), .A2(n7571), .ZN(n6379) );
  INV_X1 U6526 ( .A(n6217), .ZN(n6357) );
  OR2_X1 U6527 ( .A1(n9651), .A2(n9527), .ZN(n9067) );
  AND2_X1 U6528 ( .A1(n8416), .A2(n6597), .ZN(n8445) );
  AND2_X1 U6529 ( .A1(n7155), .A2(n7154), .ZN(n7290) );
  NAND2_X1 U6530 ( .A1(n7352), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7518) );
  INV_X1 U6531 ( .A(n9942), .ZN(n9738) );
  AND2_X1 U6532 ( .A1(n8732), .A2(n8711), .ZN(n9925) );
  OR2_X1 U6533 ( .A1(n6883), .A2(n6882), .ZN(n6920) );
  INV_X1 U6534 ( .A(n9134), .ZN(n9135) );
  NAND2_X1 U6535 ( .A1(n8959), .A2(n9128), .ZN(n9117) );
  INV_X1 U6536 ( .A(n9922), .ZN(n10094) );
  NAND2_X1 U6537 ( .A1(n6396), .A2(n6395), .ZN(n6400) );
  INV_X1 U6538 ( .A(SI_4_), .ZN(n10193) );
  INV_X1 U6539 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10563) );
  NAND2_X1 U6540 ( .A1(n9098), .A2(n10742), .ZN(n9180) );
  AND2_X1 U6541 ( .A1(n9257), .A2(n10791), .ZN(n9244) );
  NOR2_X1 U6542 ( .A1(n6379), .A2(n6356), .ZN(n9220) );
  AND2_X1 U6543 ( .A1(n6364), .A2(n6363), .ZN(n9374) );
  AND2_X1 U6544 ( .A1(n6138), .A2(n6137), .ZN(n9510) );
  AND2_X1 U6545 ( .A1(n7014), .A2(n7013), .ZN(n10726) );
  INV_X1 U6546 ( .A(n9559), .ZN(n10791) );
  AND2_X1 U6547 ( .A1(n9544), .A2(n10750), .ZN(n10904) );
  OR2_X1 U6548 ( .A1(n9700), .A2(n6336), .ZN(n10613) );
  AND2_X1 U6549 ( .A1(n5788), .A2(n5827), .ZN(n6999) );
  INV_X1 U6550 ( .A(n9794), .ZN(n9805) );
  AND3_X1 U6551 ( .A1(n8621), .A2(n8620), .A3(n8619), .ZN(n10014) );
  OR2_X1 U6552 ( .A1(n7613), .A2(n7612), .ZN(n7615) );
  INV_X1 U6553 ( .A(n9958), .ZN(n10021) );
  INV_X2 U6554 ( .A(n7185), .ZN(n8749) );
  NAND2_X1 U6555 ( .A1(n5641), .A2(n9135), .ZN(n9136) );
  OR2_X1 U6556 ( .A1(n10875), .A2(n6957), .ZN(n7074) );
  INV_X1 U6557 ( .A(n10873), .ZN(n10984) );
  AND2_X1 U6558 ( .A1(n10093), .A2(n10933), .ZN(n10098) );
  OR2_X1 U6559 ( .A1(n8972), .A2(n9037), .ZN(n10875) );
  AND2_X1 U6560 ( .A1(n6700), .A2(n6699), .ZN(n8128) );
  XNOR2_X1 U6561 ( .A(n5824), .B(n5805), .ZN(n5822) );
  AND2_X1 U6562 ( .A1(n6858), .A2(n6857), .ZN(n10718) );
  INV_X1 U6563 ( .A(n9246), .ZN(n9259) );
  INV_X1 U6564 ( .A(n9244), .ZN(n9229) );
  INV_X1 U6565 ( .A(n9197), .ZN(n9445) );
  INV_X1 U6566 ( .A(n6445), .ZN(n9280) );
  INV_X1 U6567 ( .A(n9365), .ZN(n9586) );
  AND3_X1 U6568 ( .A1(n10944), .A2(n10943), .A3(n10942), .ZN(n10949) );
  OR2_X1 U6569 ( .A1(n7291), .A2(n7656), .ZN(n10947) );
  INV_X1 U6570 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6907) );
  OR2_X1 U6571 ( .A1(n7080), .A2(n7079), .ZN(n9813) );
  AND2_X1 U6572 ( .A1(n7374), .A2(n7373), .ZN(n9133) );
  OR2_X1 U6573 ( .A1(n11006), .A2(n7420), .ZN(n10734) );
  INV_X1 U6574 ( .A(n10022), .ZN(n11006) );
  OR3_X1 U6575 ( .A1(n10738), .A2(n7506), .A3(n8724), .ZN(n10070) );
  OR2_X1 U6576 ( .A1(n7174), .A2(n7411), .ZN(n10987) );
  OR2_X1 U6577 ( .A1(n7174), .A2(n10562), .ZN(n10990) );
  CLKBUF_X1 U6578 ( .A(n10605), .Z(n10612) );
  INV_X1 U6579 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10279) );
  INV_X1 U6580 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6833) );
  NOR2_X1 U6581 ( .A1(n8334), .A2(n8333), .ZN(n10642) );
  NOR2_X1 U6582 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5645) );
  INV_X1 U6583 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5642) );
  INV_X1 U6584 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5646) );
  INV_X1 U6585 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5652) );
  NAND2_X1 U6586 ( .A1(n6076), .A2(n5652), .ZN(n5653) );
  NAND2_X1 U6587 ( .A1(n5653), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5660) );
  INV_X1 U6588 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5659) );
  NAND2_X1 U6589 ( .A1(n5660), .A2(n5659), .ZN(n5661) );
  XNOR2_X2 U6590 ( .A(n5654), .B(P2_IR_REG_20__SCAN_IN), .ZN(n5697) );
  INV_X1 U6591 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5655) );
  NAND2_X1 U6592 ( .A1(n5659), .A2(n5655), .ZN(n5668) );
  NOR2_X1 U6593 ( .A1(n5668), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U6594 ( .A1(n5657), .A2(n5656), .ZN(n5663) );
  INV_X1 U6595 ( .A(n5663), .ZN(n5658) );
  INV_X1 U6596 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5667) );
  NAND2_X1 U6597 ( .A1(n5658), .A2(n5667), .ZN(n6319) );
  INV_X1 U6598 ( .A(n6355), .ZN(n8371) );
  NAND2_X1 U6599 ( .A1(n5697), .A2(n8371), .ZN(n5665) );
  OR2_X1 U6600 ( .A1(n5660), .A2(n5659), .ZN(n5662) );
  NAND2_X1 U6601 ( .A1(n5663), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5664) );
  NAND3_X1 U6602 ( .A1(n5665), .A2(n9546), .A3(n6573), .ZN(n7143) );
  NAND2_X1 U6603 ( .A1(n7143), .A2(n8174), .ZN(n5666) );
  NAND2_X1 U6604 ( .A1(n6369), .A2(n6435), .ZN(n7147) );
  NAND2_X4 U6605 ( .A1(n5666), .A2(n7147), .ZN(n6310) );
  INV_X1 U6606 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6322) );
  INV_X1 U6607 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6325) );
  AND4_X1 U6608 ( .A1(n6322), .A2(n5667), .A3(n6325), .A4(n6327), .ZN(n5672)
         );
  NOR2_X1 U6609 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n5671) );
  INV_X1 U6610 ( .A(n5668), .ZN(n5670) );
  NOR2_X1 U6611 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5669) );
  NAND4_X1 U6612 ( .A1(n5672), .A2(n5671), .A3(n5670), .A4(n5669), .ZN(n5673)
         );
  INV_X1 U6613 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5684) );
  INV_X1 U6614 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5685) );
  INV_X1 U6615 ( .A(n5686), .ZN(n5676) );
  INV_X1 U6616 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6786) );
  OR2_X1 U6617 ( .A1(n5722), .A2(n6786), .ZN(n5683) );
  INV_X1 U6618 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5678) );
  AND2_X1 U6619 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5679) );
  INV_X1 U6620 ( .A(SI_1_), .ZN(n5681) );
  XNOR2_X1 U6621 ( .A(n5718), .B(n5681), .ZN(n5717) );
  MUX2_X1 U6622 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5720), .Z(n5716) );
  XNOR2_X1 U6623 ( .A(n5717), .B(n5716), .ZN(n7114) );
  XNOR2_X1 U6624 ( .A(n5046), .B(n7674), .ZN(n5713) );
  XNOR2_X2 U6625 ( .A(n5687), .B(P2_IR_REG_30__SCAN_IN), .ZN(n9694) );
  NAND2_X1 U6626 ( .A1(n5689), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5690) );
  NOR2_X2 U6627 ( .A1(n9694), .A2(n9062), .ZN(n5767) );
  NAND2_X1 U6628 ( .A1(n5767), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5696) );
  INV_X1 U6629 ( .A(n9062), .ZN(n5692) );
  AND2_X2 U6630 ( .A1(n9694), .A2(n5692), .ZN(n5737) );
  NAND2_X1 U6631 ( .A1(n5737), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5694) );
  NOR2_X2 U6632 ( .A1(n9694), .A2(n5692), .ZN(n5727) );
  NAND2_X1 U6633 ( .A1(n5727), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5693) );
  INV_X1 U6634 ( .A(n5697), .ZN(n8063) );
  INV_X1 U6635 ( .A(n6354), .ZN(n5699) );
  AND2_X4 U6636 ( .A1(n5699), .A2(n5698), .ZN(n6628) );
  NAND2_X1 U6637 ( .A1(n5737), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U6638 ( .A1(n5767), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5701) );
  NAND2_X1 U6639 ( .A1(n5727), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U6640 ( .A1(n5680), .A2(SI_0_), .ZN(n5705) );
  INV_X1 U6641 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5704) );
  NAND2_X1 U6642 ( .A1(n5705), .A2(n5704), .ZN(n5707) );
  AND2_X1 U6643 ( .A1(n5707), .A2(n5706), .ZN(n9701) );
  INV_X1 U6644 ( .A(n10742), .ZN(n9102) );
  NAND2_X1 U6645 ( .A1(n6310), .A2(n9102), .ZN(n9183) );
  OAI21_X1 U6646 ( .B1(n9180), .B2(n6628), .A(n9183), .ZN(n5710) );
  INV_X1 U6647 ( .A(n5710), .ZN(n5711) );
  NAND2_X1 U6648 ( .A1(n9179), .A2(n5711), .ZN(n7566) );
  INV_X1 U6649 ( .A(n5712), .ZN(n5714) );
  OR2_X1 U6650 ( .A1(n5714), .A2(n5713), .ZN(n5715) );
  NAND2_X1 U6651 ( .A1(n7566), .A2(n5715), .ZN(n5732) );
  NAND2_X1 U6652 ( .A1(n5718), .A2(SI_1_), .ZN(n5719) );
  MUX2_X1 U6653 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5720), .Z(n5745) );
  INV_X1 U6654 ( .A(SI_2_), .ZN(n5721) );
  XNOR2_X1 U6655 ( .A(n5745), .B(n5721), .ZN(n5744) );
  XNOR2_X1 U6656 ( .A(n5743), .B(n5744), .ZN(n7105) );
  OR2_X1 U6657 ( .A1(n5762), .A2(n7105), .ZN(n5726) );
  INV_X1 U6658 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6788) );
  OR2_X1 U6659 ( .A1(n5722), .A2(n6788), .ZN(n5725) );
  NAND2_X1 U6660 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5066), .ZN(n5723) );
  XNOR2_X1 U6661 ( .A(n5723), .B(P2_IR_REG_2__SCAN_IN), .ZN(n10723) );
  INV_X1 U6662 ( .A(n10723), .ZN(n6787) );
  OR2_X1 U6663 ( .A1(n7012), .A2(n6787), .ZN(n5724) );
  XNOR2_X1 U6664 ( .A(n6310), .B(n10752), .ZN(n5733) );
  NAND2_X1 U6665 ( .A1(n5727), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5731) );
  NAND2_X1 U6666 ( .A1(n5767), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5729) );
  NAND2_X1 U6667 ( .A1(n5737), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5728) );
  NAND2_X1 U6668 ( .A1(n9281), .A2(n9101), .ZN(n5734) );
  XNOR2_X1 U6669 ( .A(n5733), .B(n5734), .ZN(n7567) );
  INV_X1 U6670 ( .A(n5733), .ZN(n5735) );
  NAND2_X1 U6671 ( .A1(n5735), .A2(n5734), .ZN(n5736) );
  NAND2_X1 U6672 ( .A1(n5727), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5741) );
  NAND2_X1 U6673 ( .A1(n5767), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5740) );
  INV_X1 U6674 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7049) );
  NAND2_X1 U6675 ( .A1(n5737), .A2(n7049), .ZN(n5739) );
  NAND2_X1 U6676 ( .A1(n5768), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5738) );
  NOR2_X1 U6677 ( .A1(n6445), .A2(n6628), .ZN(n5750) );
  OAI21_X1 U6678 ( .B1(P2_IR_REG_2__SCAN_IN), .B2(n5066), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5742) );
  XNOR2_X1 U6679 ( .A(n5742), .B(P2_IR_REG_3__SCAN_IN), .ZN(n7003) );
  INV_X1 U6680 ( .A(n7003), .ZN(n7056) );
  NAND2_X1 U6681 ( .A1(n5745), .A2(SI_2_), .ZN(n5746) );
  MUX2_X1 U6682 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n6789), .Z(n5757) );
  INV_X1 U6683 ( .A(SI_3_), .ZN(n5747) );
  XNOR2_X1 U6684 ( .A(n5756), .B(n5755), .ZN(n7186) );
  OR2_X1 U6685 ( .A1(n7186), .A2(n5762), .ZN(n5749) );
  INV_X1 U6686 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6790) );
  XNOR2_X1 U6687 ( .A(n5047), .B(n10759), .ZN(n5751) );
  NAND2_X1 U6688 ( .A1(n5750), .A2(n5751), .ZN(n5773) );
  INV_X1 U6689 ( .A(n5750), .ZN(n5752) );
  INV_X1 U6690 ( .A(n5751), .ZN(n9212) );
  NAND2_X1 U6691 ( .A1(n5752), .A2(n9212), .ZN(n5753) );
  NAND2_X1 U6692 ( .A1(n5773), .A2(n5753), .ZN(n7733) );
  NAND2_X1 U6693 ( .A1(n5756), .A2(n5755), .ZN(n5759) );
  NAND2_X1 U6694 ( .A1(n5757), .A2(SI_3_), .ZN(n5758) );
  XNOR2_X1 U6695 ( .A(n5779), .B(n5778), .ZN(n7243) );
  OR2_X1 U6696 ( .A1(n7243), .A2(n5762), .ZN(n5766) );
  OR2_X1 U6697 ( .A1(n5763), .A2(n5651), .ZN(n5764) );
  XNOR2_X1 U6698 ( .A(n5764), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7001) );
  AOI22_X1 U6699 ( .A1(n5783), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n5041), .B2(
        n7001), .ZN(n5765) );
  XNOR2_X1 U6700 ( .A(n6310), .B(n10775), .ZN(n5775) );
  OAI21_X1 U6701 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n5791), .ZN(n7754) );
  INV_X1 U6702 ( .A(n7754), .ZN(n9215) );
  NAND2_X1 U6703 ( .A1(n5737), .A2(n9215), .ZN(n5772) );
  NAND2_X1 U6704 ( .A1(n6403), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5771) );
  NAND2_X1 U6705 ( .A1(n5727), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5770) );
  NAND2_X1 U6706 ( .A1(n5768), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U6707 ( .A1(n10790), .A2(n9101), .ZN(n5776) );
  XNOR2_X1 U6708 ( .A(n5775), .B(n5776), .ZN(n9218) );
  AND2_X1 U6709 ( .A1(n9218), .A2(n5773), .ZN(n5774) );
  NAND2_X1 U6710 ( .A1(n9217), .A2(n5774), .ZN(n8782) );
  INV_X1 U6711 ( .A(n5775), .ZN(n8780) );
  NAND2_X1 U6712 ( .A1(n8780), .A2(n5776), .ZN(n5777) );
  NAND2_X1 U6713 ( .A1(n8782), .A2(n5777), .ZN(n5797) );
  NAND2_X1 U6714 ( .A1(n5780), .A2(SI_4_), .ZN(n5781) );
  MUX2_X1 U6715 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n6789), .Z(n5803) );
  INV_X1 U6716 ( .A(SI_5_), .ZN(n5782) );
  XNOR2_X1 U6717 ( .A(n5802), .B(n5801), .ZN(n7340) );
  OR2_X1 U6718 ( .A1(n7340), .A2(n5762), .ZN(n5790) );
  NOR2_X1 U6719 ( .A1(n5784), .A2(n5651), .ZN(n5785) );
  MUX2_X1 U6720 ( .A(n5651), .B(n5785), .S(P2_IR_REG_5__SCAN_IN), .Z(n5786) );
  INV_X1 U6721 ( .A(n5786), .ZN(n5788) );
  INV_X1 U6722 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5787) );
  NAND2_X1 U6723 ( .A1(n5784), .A2(n5787), .ZN(n5827) );
  AOI22_X1 U6724 ( .A1(n5783), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n5041), .B2(
        n6999), .ZN(n5789) );
  NAND2_X1 U6725 ( .A1(n5790), .A2(n5789), .ZN(n10795) );
  XNOR2_X1 U6726 ( .A(n6214), .B(n10795), .ZN(n5798) );
  NAND2_X1 U6727 ( .A1(n5768), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5796) );
  NAND2_X1 U6728 ( .A1(n6403), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5795) );
  INV_X1 U6729 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7037) );
  NAND2_X1 U6730 ( .A1(n5791), .A2(n7037), .ZN(n5792) );
  AND2_X1 U6731 ( .A1(n5811), .A2(n5792), .ZN(n10797) );
  NAND2_X1 U6732 ( .A1(n5737), .A2(n10797), .ZN(n5794) );
  NAND2_X1 U6733 ( .A1(n6414), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5793) );
  OR2_X1 U6734 ( .A1(n9562), .A2(n6628), .ZN(n5799) );
  XNOR2_X1 U6735 ( .A(n5798), .B(n5799), .ZN(n8783) );
  NAND2_X1 U6736 ( .A1(n5797), .A2(n8783), .ZN(n8788) );
  INV_X1 U6737 ( .A(n5798), .ZN(n7582) );
  NAND2_X1 U6738 ( .A1(n5799), .A2(n7582), .ZN(n5800) );
  NAND2_X1 U6739 ( .A1(n8788), .A2(n5800), .ZN(n5817) );
  NAND2_X1 U6740 ( .A1(n5803), .A2(SI_5_), .ZN(n5804) );
  MUX2_X1 U6741 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6789), .Z(n5824) );
  INV_X1 U6742 ( .A(SI_6_), .ZN(n5805) );
  XNOR2_X1 U6743 ( .A(n5823), .B(n5822), .ZN(n7436) );
  OR2_X1 U6744 ( .A1(n7436), .A2(n5762), .ZN(n5808) );
  NAND2_X1 U6745 ( .A1(n5827), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5806) );
  XNOR2_X1 U6746 ( .A(n5806), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6998) );
  AOI22_X1 U6747 ( .A1(n5783), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5041), .B2(
        n6998), .ZN(n5807) );
  NAND2_X1 U6748 ( .A1(n5808), .A2(n5807), .ZN(n10821) );
  XNOR2_X1 U6749 ( .A(n10821), .B(n6214), .ZN(n5818) );
  NAND2_X1 U6750 ( .A1(n5768), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5816) );
  NAND2_X1 U6751 ( .A1(n6403), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5815) );
  INV_X1 U6752 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5810) );
  NAND2_X1 U6753 ( .A1(n5811), .A2(n5810), .ZN(n5812) );
  AND2_X1 U6754 ( .A1(n5831), .A2(n5812), .ZN(n9567) );
  NAND2_X1 U6755 ( .A1(n5737), .A2(n9567), .ZN(n5814) );
  NAND2_X1 U6756 ( .A1(n6414), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5813) );
  NAND4_X1 U6757 ( .A1(n5816), .A2(n5815), .A3(n5814), .A4(n5813), .ZN(n10792)
         );
  NAND2_X1 U6758 ( .A1(n10792), .A2(n9101), .ZN(n5819) );
  XNOR2_X1 U6759 ( .A(n5818), .B(n5819), .ZN(n7583) );
  NAND2_X1 U6760 ( .A1(n5817), .A2(n7583), .ZN(n7588) );
  INV_X1 U6761 ( .A(n5818), .ZN(n5820) );
  NAND2_X1 U6762 ( .A1(n5820), .A2(n5819), .ZN(n5821) );
  NAND2_X1 U6763 ( .A1(n5824), .A2(SI_6_), .ZN(n5825) );
  NAND2_X1 U6764 ( .A1(n5826), .A2(n5825), .ZN(n5845) );
  MUX2_X1 U6765 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5720), .Z(n5846) );
  XNOR2_X1 U6766 ( .A(n5845), .B(n5843), .ZN(n7512) );
  INV_X2 U6767 ( .A(n5762), .ZN(n6421) );
  NAND2_X1 U6768 ( .A1(n7512), .A2(n6421), .ZN(n5830) );
  NAND2_X1 U6769 ( .A1(n5853), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5828) );
  XNOR2_X1 U6770 ( .A(n5828), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7085) );
  AOI22_X1 U6771 ( .A1(n5783), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5041), .B2(
        n7085), .ZN(n5829) );
  NAND2_X1 U6772 ( .A1(n5830), .A2(n5829), .ZN(n7813) );
  XNOR2_X1 U6773 ( .A(n7813), .B(n6214), .ZN(n5837) );
  INV_X2 U6774 ( .A(n6109), .ZN(n6413) );
  NAND2_X1 U6775 ( .A1(n6413), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5836) );
  NAND2_X1 U6776 ( .A1(n6403), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5835) );
  INV_X1 U6777 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7589) );
  NAND2_X1 U6778 ( .A1(n5831), .A2(n7589), .ZN(n5832) );
  AND2_X1 U6779 ( .A1(n5857), .A2(n5832), .ZN(n7812) );
  NAND2_X1 U6780 ( .A1(n6217), .A2(n7812), .ZN(n5834) );
  NAND2_X1 U6781 ( .A1(n6414), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5833) );
  NOR2_X1 U6782 ( .A1(n9560), .A2(n6628), .ZN(n5838) );
  NAND2_X1 U6783 ( .A1(n5837), .A2(n5838), .ZN(n5842) );
  INV_X1 U6784 ( .A(n5837), .ZN(n7644) );
  INV_X1 U6785 ( .A(n5838), .ZN(n5839) );
  NAND2_X1 U6786 ( .A1(n7644), .A2(n5839), .ZN(n5840) );
  NAND2_X1 U6787 ( .A1(n5842), .A2(n5840), .ZN(n7592) );
  NAND2_X1 U6788 ( .A1(n5845), .A2(n5844), .ZN(n5848) );
  NAND2_X1 U6789 ( .A1(n5846), .A2(SI_7_), .ZN(n5847) );
  MUX2_X1 U6790 ( .A(n6831), .B(n6833), .S(n5720), .Z(n5850) );
  INV_X1 U6791 ( .A(SI_8_), .ZN(n5849) );
  INV_X1 U6792 ( .A(n5850), .ZN(n5851) );
  NAND2_X1 U6793 ( .A1(n5851), .A2(SI_8_), .ZN(n5852) );
  XNOR2_X1 U6794 ( .A(n5870), .B(n5869), .ZN(n7819) );
  NAND2_X1 U6795 ( .A1(n7819), .A2(n6421), .ZN(n5856) );
  NOR2_X1 U6796 ( .A1(n5853), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5879) );
  OR2_X1 U6797 ( .A1(n5879), .A2(n5651), .ZN(n5854) );
  XNOR2_X1 U6798 ( .A(n5854), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7221) );
  AOI22_X1 U6799 ( .A1(n5783), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5041), .B2(
        n7221), .ZN(n5855) );
  NAND2_X1 U6800 ( .A1(n5856), .A2(n5855), .ZN(n7943) );
  XNOR2_X1 U6801 ( .A(n7943), .B(n6214), .ZN(n7604) );
  NAND2_X1 U6802 ( .A1(n6413), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U6803 ( .A1(n6403), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5861) );
  NAND2_X1 U6804 ( .A1(n5857), .A2(n7650), .ZN(n5858) );
  AND2_X1 U6805 ( .A1(n5883), .A2(n5858), .ZN(n7768) );
  NAND2_X1 U6806 ( .A1(n6217), .A2(n7768), .ZN(n5860) );
  NAND2_X1 U6807 ( .A1(n6414), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5859) );
  NOR2_X1 U6808 ( .A1(n7603), .A2(n6628), .ZN(n5863) );
  NAND2_X1 U6809 ( .A1(n7604), .A2(n5863), .ZN(n5889) );
  INV_X1 U6810 ( .A(n7604), .ZN(n5865) );
  INV_X1 U6811 ( .A(n5863), .ZN(n5864) );
  NAND2_X1 U6812 ( .A1(n5865), .A2(n5864), .ZN(n5866) );
  AND2_X1 U6813 ( .A1(n5889), .A2(n5866), .ZN(n7641) );
  NAND2_X1 U6814 ( .A1(n5867), .A2(n7641), .ZN(n7602) );
  OAI21_X1 U6815 ( .B1(n5870), .B2(n5869), .A(n5868), .ZN(n5876) );
  INV_X1 U6816 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5871) );
  MUX2_X1 U6817 ( .A(n5871), .B(n6872), .S(n5720), .Z(n5872) );
  INV_X1 U6818 ( .A(SI_9_), .ZN(n10186) );
  INV_X1 U6819 ( .A(n5872), .ZN(n5873) );
  NAND2_X1 U6820 ( .A1(n5873), .A2(SI_9_), .ZN(n5874) );
  NAND2_X1 U6821 ( .A1(n5876), .A2(n5875), .ZN(n5896) );
  OR2_X1 U6822 ( .A1(n5876), .A2(n5875), .ZN(n5877) );
  NAND2_X1 U6823 ( .A1(n5896), .A2(n5877), .ZN(n7859) );
  NAND2_X1 U6824 ( .A1(n7859), .A2(n6421), .ZN(n5881) );
  INV_X1 U6825 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U6826 ( .A1(n5879), .A2(n5878), .ZN(n5951) );
  NAND2_X1 U6827 ( .A1(n5951), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5900) );
  XNOR2_X1 U6828 ( .A(n5900), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7377) );
  AOI22_X1 U6829 ( .A1(n5783), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5041), .B2(
        n7377), .ZN(n5880) );
  XNOR2_X1 U6830 ( .A(n10863), .B(n6310), .ZN(n5893) );
  NAND2_X1 U6831 ( .A1(n6403), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U6832 ( .A1(n6413), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5887) );
  INV_X1 U6833 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7226) );
  NAND2_X1 U6834 ( .A1(n5883), .A2(n7226), .ZN(n5884) );
  AND2_X1 U6835 ( .A1(n5904), .A2(n5884), .ZN(n7952) );
  NAND2_X1 U6836 ( .A1(n5737), .A2(n7952), .ZN(n5886) );
  NAND2_X1 U6837 ( .A1(n6414), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5885) );
  NOR2_X1 U6838 ( .A1(n7986), .A2(n6628), .ZN(n5891) );
  XNOR2_X1 U6839 ( .A(n5893), .B(n5891), .ZN(n7606) );
  AND2_X1 U6840 ( .A1(n7606), .A2(n5889), .ZN(n5890) );
  NAND2_X1 U6841 ( .A1(n7602), .A2(n5890), .ZN(n7611) );
  INV_X1 U6842 ( .A(n5891), .ZN(n5892) );
  NAND2_X1 U6843 ( .A1(n5893), .A2(n5892), .ZN(n5894) );
  NAND2_X1 U6844 ( .A1(n7611), .A2(n5894), .ZN(n7844) );
  NAND2_X1 U6845 ( .A1(n5896), .A2(n5895), .ZN(n5915) );
  MUX2_X1 U6846 ( .A(n6907), .B(n6908), .S(n5720), .Z(n5897) );
  INV_X1 U6847 ( .A(SI_10_), .ZN(n10144) );
  INV_X1 U6848 ( .A(n5897), .ZN(n5898) );
  NAND2_X1 U6849 ( .A1(n5898), .A2(SI_10_), .ZN(n5899) );
  XNOR2_X1 U6850 ( .A(n5915), .B(n5636), .ZN(n7919) );
  NAND2_X1 U6851 ( .A1(n7919), .A2(n6421), .ZN(n5903) );
  NAND2_X1 U6852 ( .A1(n5900), .A2(n5949), .ZN(n5901) );
  NAND2_X1 U6853 ( .A1(n5901), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5919) );
  XNOR2_X1 U6854 ( .A(n5919), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7794) );
  AOI22_X1 U6855 ( .A1(n5783), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7794), .B2(
        n5041), .ZN(n5902) );
  XNOR2_X1 U6856 ( .A(n8029), .B(n6214), .ZN(n5910) );
  NAND2_X1 U6857 ( .A1(n6403), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U6858 ( .A1(n6413), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U6859 ( .A1(n5904), .A2(n10140), .ZN(n5905) );
  AND2_X1 U6860 ( .A1(n5925), .A2(n5905), .ZN(n7990) );
  NAND2_X1 U6861 ( .A1(n6217), .A2(n7990), .ZN(n5907) );
  NAND2_X1 U6862 ( .A1(n6414), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5906) );
  NOR2_X1 U6863 ( .A1(n9239), .A2(n6628), .ZN(n5911) );
  NAND2_X1 U6864 ( .A1(n5910), .A2(n5911), .ZN(n5914) );
  INV_X1 U6865 ( .A(n5910), .ZN(n9238) );
  INV_X1 U6866 ( .A(n5911), .ZN(n5912) );
  NAND2_X1 U6867 ( .A1(n9238), .A2(n5912), .ZN(n5913) );
  NAND2_X1 U6868 ( .A1(n5914), .A2(n5913), .ZN(n7845) );
  NAND2_X1 U6869 ( .A1(n5915), .A2(n5636), .ZN(n5917) );
  MUX2_X1 U6870 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6789), .Z(n5936) );
  INV_X1 U6871 ( .A(SI_11_), .ZN(n5918) );
  XNOR2_X1 U6872 ( .A(n5939), .B(n5935), .ZN(n8015) );
  NAND2_X1 U6873 ( .A1(n8015), .A2(n6421), .ZN(n5923) );
  NAND2_X1 U6874 ( .A1(n5919), .A2(n5948), .ZN(n5920) );
  NAND2_X1 U6875 ( .A1(n5920), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5921) );
  XNOR2_X1 U6876 ( .A(n5921), .B(P2_IR_REG_11__SCAN_IN), .ZN(n9285) );
  AOI22_X1 U6877 ( .A1(n9285), .A2(n5041), .B1(n5783), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n5922) );
  NAND2_X1 U6878 ( .A1(n5923), .A2(n5922), .ZN(n10901) );
  XNOR2_X1 U6879 ( .A(n10901), .B(n6214), .ZN(n5931) );
  NAND2_X1 U6880 ( .A1(n6403), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5930) );
  NAND2_X1 U6881 ( .A1(n6413), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5929) );
  INV_X1 U6882 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10137) );
  NAND2_X1 U6883 ( .A1(n5925), .A2(n10137), .ZN(n5926) );
  AND2_X1 U6884 ( .A1(n5955), .A2(n5926), .ZN(n9245) );
  NAND2_X1 U6885 ( .A1(n6217), .A2(n9245), .ZN(n5928) );
  NAND2_X1 U6886 ( .A1(n6414), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5927) );
  NOR2_X1 U6887 ( .A1(n8075), .A2(n6628), .ZN(n5932) );
  NAND2_X1 U6888 ( .A1(n5931), .A2(n5932), .ZN(n5961) );
  INV_X1 U6889 ( .A(n5931), .ZN(n8000) );
  INV_X1 U6890 ( .A(n5932), .ZN(n5933) );
  NAND2_X1 U6891 ( .A1(n8000), .A2(n5933), .ZN(n5934) );
  AND2_X1 U6892 ( .A1(n5961), .A2(n5934), .ZN(n9235) );
  NAND2_X1 U6893 ( .A1(n5936), .A2(SI_11_), .ZN(n5937) );
  INV_X1 U6894 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5940) );
  MUX2_X1 U6895 ( .A(n5940), .B(n10279), .S(n5720), .Z(n5941) );
  INV_X1 U6896 ( .A(SI_12_), .ZN(n10146) );
  INV_X1 U6897 ( .A(n5941), .ZN(n5942) );
  NAND2_X1 U6898 ( .A1(n5942), .A2(SI_12_), .ZN(n5943) );
  NAND2_X1 U6899 ( .A1(n5945), .A2(n5944), .ZN(n5946) );
  NAND2_X1 U6900 ( .A1(n5967), .A2(n5946), .ZN(n8127) );
  NAND2_X1 U6901 ( .A1(n8127), .A2(n6421), .ZN(n5954) );
  INV_X1 U6902 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5947) );
  NAND3_X1 U6903 ( .A1(n5949), .A2(n5948), .A3(n5947), .ZN(n5950) );
  OR2_X1 U6904 ( .A1(n5951), .A2(n5950), .ZN(n5972) );
  NAND2_X1 U6905 ( .A1(n5972), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5952) );
  XNOR2_X1 U6906 ( .A(n5952), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7907) );
  AOI22_X1 U6907 ( .A1(n5783), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5041), .B2(
        n7907), .ZN(n5953) );
  NAND2_X1 U6908 ( .A1(n5954), .A2(n5953), .ZN(n8095) );
  XNOR2_X1 U6909 ( .A(n8095), .B(n6310), .ZN(n8558) );
  NAND2_X1 U6910 ( .A1(n6403), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U6911 ( .A1(n6414), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5959) );
  INV_X1 U6912 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7790) );
  NAND2_X1 U6913 ( .A1(n5955), .A2(n7790), .ZN(n5956) );
  AND2_X1 U6914 ( .A1(n5975), .A2(n5956), .ZN(n8085) );
  NAND2_X1 U6915 ( .A1(n5737), .A2(n8085), .ZN(n5958) );
  NAND2_X1 U6916 ( .A1(n6413), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5957) );
  NOR2_X1 U6917 ( .A1(n8559), .A2(n6628), .ZN(n5963) );
  XNOR2_X1 U6918 ( .A(n8558), .B(n5963), .ZN(n8012) );
  AND2_X1 U6919 ( .A1(n8012), .A2(n5961), .ZN(n5962) );
  INV_X1 U6920 ( .A(n5963), .ZN(n5964) );
  NAND2_X1 U6921 ( .A1(n8558), .A2(n5964), .ZN(n5965) );
  INV_X1 U6922 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7295) );
  INV_X1 U6923 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7296) );
  MUX2_X1 U6924 ( .A(n7295), .B(n7296), .S(n6789), .Z(n5969) );
  INV_X1 U6925 ( .A(SI_13_), .ZN(n5968) );
  NAND2_X1 U6926 ( .A1(n5969), .A2(n5968), .ZN(n5984) );
  INV_X1 U6927 ( .A(n5969), .ZN(n5970) );
  NAND2_X1 U6928 ( .A1(n5970), .A2(SI_13_), .ZN(n5971) );
  XNOR2_X1 U6929 ( .A(n5983), .B(n5635), .ZN(n8234) );
  NAND2_X1 U6930 ( .A1(n8234), .A2(n6421), .ZN(n5974) );
  OAI21_X1 U6931 ( .B1(n5972), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5988) );
  XNOR2_X1 U6932 ( .A(n5988), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8051) );
  AOI22_X1 U6933 ( .A1(n8051), .A2(n5041), .B1(n5783), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n5973) );
  XNOR2_X1 U6934 ( .A(n10938), .B(n6310), .ZN(n8768) );
  NAND2_X1 U6935 ( .A1(n6413), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5980) );
  NAND2_X1 U6936 ( .A1(n6403), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5979) );
  INV_X1 U6937 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10231) );
  NAND2_X1 U6938 ( .A1(n5975), .A2(n10231), .ZN(n5976) );
  AND2_X1 U6939 ( .A1(n5996), .A2(n5976), .ZN(n8564) );
  NAND2_X1 U6940 ( .A1(n5737), .A2(n8564), .ZN(n5978) );
  NAND2_X1 U6941 ( .A1(n6414), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5977) );
  NOR2_X1 U6942 ( .A1(n8767), .A2(n6628), .ZN(n5981) );
  XNOR2_X1 U6943 ( .A(n8768), .B(n5981), .ZN(n8557) );
  INV_X1 U6944 ( .A(n5981), .ZN(n5982) );
  INV_X1 U6945 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7333) );
  INV_X1 U6946 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5986) );
  MUX2_X1 U6947 ( .A(n7333), .B(n5986), .S(n5720), .Z(n6006) );
  XNOR2_X1 U6948 ( .A(n6009), .B(n6005), .ZN(n8242) );
  NAND2_X1 U6949 ( .A1(n8242), .A2(n6421), .ZN(n5994) );
  INV_X1 U6950 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U6951 ( .A1(n5988), .A2(n5987), .ZN(n5989) );
  NAND2_X1 U6952 ( .A1(n5989), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U6953 ( .A1(n5991), .A2(n5990), .ZN(n6010) );
  OR2_X1 U6954 ( .A1(n5991), .A2(n5990), .ZN(n5992) );
  AOI22_X1 U6955 ( .A1(n8199), .A2(n5041), .B1(n5783), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5993) );
  XNOR2_X1 U6956 ( .A(n9664), .B(n6310), .ZN(n9053) );
  NAND2_X1 U6957 ( .A1(n6413), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6001) );
  INV_X1 U6958 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U6959 ( .A1(n5996), .A2(n5995), .ZN(n5997) );
  AND2_X1 U6960 ( .A1(n6016), .A2(n5997), .ZN(n8760) );
  NAND2_X1 U6961 ( .A1(n6217), .A2(n8760), .ZN(n6000) );
  NAND2_X1 U6962 ( .A1(n6403), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5999) );
  NAND2_X1 U6963 ( .A1(n6414), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5998) );
  NOR2_X1 U6964 ( .A1(n9052), .A2(n6628), .ZN(n6002) );
  XNOR2_X1 U6965 ( .A(n9053), .B(n6002), .ZN(n8766) );
  INV_X1 U6966 ( .A(n6002), .ZN(n6003) );
  NAND2_X1 U6967 ( .A1(n9053), .A2(n6003), .ZN(n6004) );
  NAND2_X1 U6968 ( .A1(n8759), .A2(n6004), .ZN(n6022) );
  INV_X1 U6969 ( .A(n6006), .ZN(n6007) );
  NAND2_X1 U6970 ( .A1(n6007), .A2(SI_14_), .ZN(n6008) );
  MUX2_X1 U6971 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6789), .Z(n6029) );
  XNOR2_X1 U6972 ( .A(n6029), .B(SI_15_), .ZN(n6026) );
  XNOR2_X1 U6973 ( .A(n6028), .B(n6026), .ZN(n8372) );
  NAND2_X1 U6974 ( .A1(n8372), .A2(n6421), .ZN(n6013) );
  NAND2_X1 U6975 ( .A1(n6010), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6011) );
  XNOR2_X1 U6976 ( .A(n6011), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9302) );
  AOI22_X1 U6977 ( .A1(n9302), .A2(n5041), .B1(n5783), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6012) );
  XNOR2_X1 U6978 ( .A(n9659), .B(n6310), .ZN(n8192) );
  INV_X1 U6979 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U6980 ( .A1(n6016), .A2(n6015), .ZN(n6017) );
  NAND2_X1 U6981 ( .A1(n6040), .A2(n6017), .ZN(n8443) );
  OR2_X1 U6982 ( .A1(n6357), .A2(n8443), .ZN(n6021) );
  NAND2_X1 U6983 ( .A1(n6413), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6020) );
  NAND2_X1 U6984 ( .A1(n6403), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U6985 ( .A1(n6414), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6018) );
  NOR2_X1 U6986 ( .A1(n8422), .A2(n6628), .ZN(n6023) );
  XNOR2_X1 U6987 ( .A(n8192), .B(n6023), .ZN(n9051) );
  NAND2_X1 U6988 ( .A1(n6022), .A2(n9051), .ZN(n8190) );
  INV_X1 U6989 ( .A(n6023), .ZN(n6024) );
  NAND2_X1 U6990 ( .A1(n8192), .A2(n6024), .ZN(n6025) );
  NAND2_X1 U6991 ( .A1(n8190), .A2(n6025), .ZN(n6045) );
  NAND2_X1 U6992 ( .A1(n6029), .A2(SI_15_), .ZN(n6030) );
  INV_X1 U6993 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7542) );
  INV_X1 U6994 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7540) );
  MUX2_X1 U6995 ( .A(n7542), .B(n7540), .S(n5720), .Z(n6032) );
  INV_X1 U6996 ( .A(SI_16_), .ZN(n6031) );
  NAND2_X1 U6997 ( .A1(n6032), .A2(n6031), .ZN(n6053) );
  INV_X1 U6998 ( .A(n6032), .ZN(n6033) );
  NAND2_X1 U6999 ( .A1(n6033), .A2(SI_16_), .ZN(n6034) );
  NAND2_X1 U7000 ( .A1(n6053), .A2(n6034), .ZN(n6051) );
  XNOR2_X1 U7001 ( .A(n6050), .B(n6051), .ZN(n8461) );
  NAND2_X1 U7002 ( .A1(n8461), .A2(n6421), .ZN(n6038) );
  NAND2_X1 U7003 ( .A1(n6035), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6036) );
  XNOR2_X1 U7004 ( .A(n6036), .B(P2_IR_REG_16__SCAN_IN), .ZN(n9316) );
  AOI22_X1 U7005 ( .A1(n5783), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5041), .B2(
        n9316), .ZN(n6037) );
  XNOR2_X1 U7006 ( .A(n9655), .B(n6310), .ZN(n6048) );
  INV_X1 U7007 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U7008 ( .A1(n6040), .A2(n6039), .ZN(n6041) );
  AND2_X1 U7009 ( .A1(n6059), .A2(n6041), .ZN(n8187) );
  NAND2_X1 U7010 ( .A1(n8187), .A2(n6217), .ZN(n6044) );
  AOI22_X1 U7011 ( .A1(n6413), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n6403), .B2(
        P2_REG1_REG_16__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7012 ( .A1(n6414), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6042) );
  NOR2_X1 U7013 ( .A1(n9540), .A2(n6628), .ZN(n6046) );
  XNOR2_X1 U7014 ( .A(n6048), .B(n6046), .ZN(n8191) );
  NAND2_X1 U7015 ( .A1(n6045), .A2(n8191), .ZN(n8197) );
  INV_X1 U7016 ( .A(n6046), .ZN(n6047) );
  NAND2_X1 U7017 ( .A1(n6048), .A2(n6047), .ZN(n6049) );
  INV_X1 U7018 ( .A(n6051), .ZN(n6052) );
  INV_X1 U7019 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6054) );
  INV_X1 U7020 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7626) );
  MUX2_X1 U7021 ( .A(n6054), .B(n7626), .S(n6789), .Z(n6071) );
  XNOR2_X1 U7022 ( .A(n6071), .B(SI_17_), .ZN(n6070) );
  XNOR2_X1 U7023 ( .A(n6075), .B(n6070), .ZN(n8466) );
  NAND2_X1 U7024 ( .A1(n8466), .A2(n6421), .ZN(n6058) );
  NAND2_X1 U7025 ( .A1(n6055), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6056) );
  XNOR2_X1 U7026 ( .A(n6056), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9339) );
  AOI22_X1 U7027 ( .A1(n5783), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5041), .B2(
        n9339), .ZN(n6057) );
  XNOR2_X1 U7028 ( .A(n9651), .B(n6214), .ZN(n6064) );
  INV_X1 U7029 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9319) );
  NAND2_X1 U7030 ( .A1(n6059), .A2(n9319), .ZN(n6060) );
  NAND2_X1 U7031 ( .A1(n6079), .A2(n6060), .ZN(n9550) );
  OR2_X1 U7032 ( .A1(n9550), .A2(n6357), .ZN(n6063) );
  AOI22_X1 U7033 ( .A1(n6413), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n6403), .B2(
        P2_REG1_REG_17__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7034 ( .A1(n6414), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6061) );
  NOR2_X1 U7035 ( .A1(n9066), .A2(n6628), .ZN(n6065) );
  NAND2_X1 U7036 ( .A1(n6064), .A2(n6065), .ZN(n6069) );
  INV_X1 U7037 ( .A(n6064), .ZN(n8407) );
  INV_X1 U7038 ( .A(n6065), .ZN(n6066) );
  NAND2_X1 U7039 ( .A1(n8407), .A2(n6066), .ZN(n6067) );
  NAND2_X1 U7040 ( .A1(n6069), .A2(n6067), .ZN(n6664) );
  INV_X1 U7041 ( .A(n6664), .ZN(n6068) );
  INV_X1 U7042 ( .A(n6070), .ZN(n6074) );
  INV_X1 U7043 ( .A(n6071), .ZN(n6072) );
  NAND2_X1 U7044 ( .A1(n6072), .A2(SI_17_), .ZN(n6073) );
  MUX2_X1 U7045 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6789), .Z(n6095) );
  XNOR2_X1 U7046 ( .A(n6095), .B(SI_18_), .ZN(n6092) );
  XNOR2_X1 U7047 ( .A(n6094), .B(n6092), .ZN(n8636) );
  NAND2_X1 U7048 ( .A1(n8636), .A2(n6421), .ZN(n6078) );
  XNOR2_X1 U7049 ( .A(n6076), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9347) );
  AOI22_X1 U7050 ( .A1(n5783), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5041), .B2(
        n9347), .ZN(n6077) );
  XNOR2_X1 U7051 ( .A(n9644), .B(n6310), .ZN(n6088) );
  INV_X1 U7052 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8411) );
  NAND2_X1 U7053 ( .A1(n6079), .A2(n8411), .ZN(n6080) );
  AND2_X1 U7054 ( .A1(n6104), .A2(n6080), .ZN(n9522) );
  NAND2_X1 U7055 ( .A1(n9522), .A2(n6217), .ZN(n6086) );
  INV_X1 U7056 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n6083) );
  NAND2_X1 U7057 ( .A1(n6403), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6082) );
  NAND2_X1 U7058 ( .A1(n6414), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6081) );
  OAI211_X1 U7059 ( .C1(n6083), .C2(n6109), .A(n6082), .B(n6081), .ZN(n6084)
         );
  INV_X1 U7060 ( .A(n6084), .ZN(n6085) );
  NOR2_X1 U7061 ( .A1(n9539), .A2(n6628), .ZN(n6089) );
  XNOR2_X1 U7062 ( .A(n6088), .B(n6089), .ZN(n8404) );
  NAND2_X1 U7063 ( .A1(n6087), .A2(n8404), .ZN(n8408) );
  INV_X1 U7064 ( .A(n6088), .ZN(n6090) );
  NAND2_X1 U7065 ( .A1(n6090), .A2(n6089), .ZN(n6091) );
  NAND2_X1 U7066 ( .A1(n8408), .A2(n6091), .ZN(n8454) );
  INV_X1 U7067 ( .A(n6092), .ZN(n6093) );
  NAND2_X1 U7068 ( .A1(n6095), .A2(SI_18_), .ZN(n6096) );
  INV_X1 U7069 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7916) );
  INV_X1 U7070 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10272) );
  MUX2_X1 U7071 ( .A(n7916), .B(n10272), .S(n5720), .Z(n6097) );
  INV_X1 U7072 ( .A(SI_19_), .ZN(n10172) );
  NAND2_X1 U7073 ( .A1(n6097), .A2(n10172), .ZN(n6119) );
  INV_X1 U7074 ( .A(n6097), .ZN(n6098) );
  NAND2_X1 U7075 ( .A1(n6098), .A2(SI_19_), .ZN(n6099) );
  NAND2_X1 U7076 ( .A1(n6119), .A2(n6099), .ZN(n6117) );
  XNOR2_X1 U7077 ( .A(n6118), .B(n6117), .ZN(n8610) );
  NAND2_X1 U7078 ( .A1(n8610), .A2(n6421), .ZN(n6101) );
  INV_X1 U7079 ( .A(n9546), .ZN(n10800) );
  AOI22_X1 U7080 ( .A1(n5783), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n10800), 
        .B2(n5041), .ZN(n6100) );
  XNOR2_X1 U7081 ( .A(n9641), .B(n6214), .ZN(n6113) );
  INV_X1 U7082 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7083 ( .A1(n6104), .A2(n6103), .ZN(n6105) );
  NAND2_X1 U7084 ( .A1(n6131), .A2(n6105), .ZN(n9512) );
  OR2_X1 U7085 ( .A1(n9512), .A2(n6357), .ZN(n6112) );
  INV_X1 U7086 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U7087 ( .A1(n6414), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U7088 ( .A1(n6403), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6106) );
  OAI211_X1 U7089 ( .C1(n6109), .C2(n6108), .A(n6107), .B(n6106), .ZN(n6110)
         );
  INV_X1 U7090 ( .A(n6110), .ZN(n6111) );
  NOR2_X1 U7091 ( .A1(n9068), .A2(n6628), .ZN(n6114) );
  AND2_X1 U7092 ( .A1(n6113), .A2(n6114), .ZN(n8451) );
  INV_X1 U7093 ( .A(n6113), .ZN(n6116) );
  INV_X1 U7094 ( .A(n6114), .ZN(n6115) );
  NAND2_X1 U7095 ( .A1(n6116), .A2(n6115), .ZN(n8450) );
  OAI21_X2 U7096 ( .B1(n8454), .B2(n8451), .A(n8450), .ZN(n8487) );
  INV_X1 U7097 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8652) );
  INV_X1 U7098 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6128) );
  MUX2_X1 U7099 ( .A(n8652), .B(n6128), .S(n5680), .Z(n6120) );
  INV_X1 U7100 ( .A(SI_20_), .ZN(n10170) );
  NAND2_X1 U7101 ( .A1(n6120), .A2(n10170), .ZN(n6142) );
  INV_X1 U7102 ( .A(n6120), .ZN(n6121) );
  NAND2_X1 U7103 ( .A1(n6121), .A2(SI_20_), .ZN(n6122) );
  NAND2_X1 U7104 ( .A1(n6142), .A2(n6122), .ZN(n6124) );
  NAND2_X1 U7105 ( .A1(n6123), .A2(n6124), .ZN(n6127) );
  INV_X1 U7106 ( .A(n6124), .ZN(n6125) );
  NAND2_X1 U7107 ( .A1(n6126), .A2(n6125), .ZN(n6143) );
  NAND2_X1 U7108 ( .A1(n6127), .A2(n6143), .ZN(n8651) );
  NAND2_X1 U7109 ( .A1(n8651), .A2(n6421), .ZN(n6130) );
  OR2_X1 U7110 ( .A1(n5722), .A2(n6128), .ZN(n6129) );
  XNOR2_X1 U7111 ( .A(n9634), .B(n6214), .ZN(n6140) );
  INV_X1 U7112 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10228) );
  NAND2_X1 U7113 ( .A1(n6131), .A2(n10228), .ZN(n6132) );
  AND2_X1 U7114 ( .A1(n6147), .A2(n6132), .ZN(n8488) );
  NAND2_X1 U7115 ( .A1(n8488), .A2(n5737), .ZN(n6138) );
  INV_X1 U7116 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7117 ( .A1(n6413), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U7118 ( .A1(n6403), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6133) );
  OAI211_X1 U7119 ( .C1(n6135), .C2(n6360), .A(n6134), .B(n6133), .ZN(n6136)
         );
  INV_X1 U7120 ( .A(n6136), .ZN(n6137) );
  NOR2_X1 U7121 ( .A1(n9510), .A2(n6628), .ZN(n6139) );
  XNOR2_X1 U7122 ( .A(n6140), .B(n6139), .ZN(n8486) );
  NAND2_X1 U7123 ( .A1(n6140), .A2(n6139), .ZN(n6141) );
  OAI21_X1 U7124 ( .B1(n8487), .B2(n8486), .A(n6141), .ZN(n9190) );
  MUX2_X1 U7125 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n5680), .Z(n6160) );
  INV_X1 U7126 ( .A(SI_21_), .ZN(n6144) );
  XNOR2_X1 U7127 ( .A(n6160), .B(n6144), .ZN(n6159) );
  XNOR2_X1 U7128 ( .A(n6161), .B(n6159), .ZN(n8662) );
  NAND2_X1 U7129 ( .A1(n8662), .A2(n6421), .ZN(n6146) );
  INV_X1 U7130 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8175) );
  OR2_X1 U7131 ( .A1(n5722), .A2(n8175), .ZN(n6145) );
  XNOR2_X1 U7132 ( .A(n9629), .B(n5047), .ZN(n6155) );
  NAND2_X1 U7133 ( .A1(n6147), .A2(n5141), .ZN(n6148) );
  NAND2_X1 U7134 ( .A1(n6174), .A2(n6148), .ZN(n9479) );
  OR2_X1 U7135 ( .A1(n9479), .A2(n6357), .ZN(n6154) );
  INV_X1 U7136 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7137 ( .A1(n6403), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U7138 ( .A1(n6413), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6149) );
  OAI211_X1 U7139 ( .C1(n6151), .C2(n6360), .A(n6150), .B(n6149), .ZN(n6152)
         );
  INV_X1 U7140 ( .A(n6152), .ZN(n6153) );
  NOR2_X1 U7141 ( .A1(n9266), .A2(n6628), .ZN(n6156) );
  XNOR2_X1 U7142 ( .A(n6155), .B(n6156), .ZN(n9189) );
  INV_X1 U7143 ( .A(n6155), .ZN(n6157) );
  NAND2_X1 U7144 ( .A1(n6157), .A2(n6156), .ZN(n6158) );
  INV_X1 U7145 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10266) );
  INV_X1 U7146 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n6171) );
  MUX2_X1 U7147 ( .A(n10266), .B(n6171), .S(n5680), .Z(n6164) );
  INV_X1 U7148 ( .A(SI_22_), .ZN(n6163) );
  NAND2_X1 U7149 ( .A1(n6164), .A2(n6163), .ZN(n6189) );
  INV_X1 U7150 ( .A(n6164), .ZN(n6165) );
  NAND2_X1 U7151 ( .A1(n6165), .A2(SI_22_), .ZN(n6166) );
  NAND2_X1 U7152 ( .A1(n6189), .A2(n6166), .ZN(n6169) );
  INV_X1 U7153 ( .A(n6169), .ZN(n6167) );
  NAND2_X1 U7154 ( .A1(n6162), .A2(n6169), .ZN(n6170) );
  NAND2_X1 U7155 ( .A1(n6190), .A2(n6170), .ZN(n8679) );
  NAND2_X1 U7156 ( .A1(n8679), .A2(n6421), .ZN(n6173) );
  OR2_X1 U7157 ( .A1(n5722), .A2(n6171), .ZN(n6172) );
  XNOR2_X1 U7158 ( .A(n9624), .B(n6310), .ZN(n6182) );
  INV_X1 U7159 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10233) );
  NAND2_X1 U7160 ( .A1(n6174), .A2(n10233), .ZN(n6175) );
  NAND2_X1 U7161 ( .A1(n6196), .A2(n6175), .ZN(n9462) );
  OR2_X1 U7162 ( .A1(n9462), .A2(n6357), .ZN(n6181) );
  INV_X1 U7163 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n6178) );
  NAND2_X1 U7164 ( .A1(n6403), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U7165 ( .A1(n6413), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6176) );
  OAI211_X1 U7166 ( .C1(n6178), .C2(n6360), .A(n6177), .B(n6176), .ZN(n6179)
         );
  INV_X1 U7167 ( .A(n6179), .ZN(n6180) );
  NAND2_X1 U7168 ( .A1(n6181), .A2(n6180), .ZN(n9485) );
  NAND2_X1 U7169 ( .A1(n9485), .A2(n9101), .ZN(n6183) );
  NAND2_X1 U7170 ( .A1(n6182), .A2(n6183), .ZN(n6188) );
  INV_X1 U7171 ( .A(n6182), .ZN(n6185) );
  INV_X1 U7172 ( .A(n6183), .ZN(n6184) );
  NAND2_X1 U7173 ( .A1(n6185), .A2(n6184), .ZN(n6186) );
  NAND2_X1 U7174 ( .A1(n6188), .A2(n6186), .ZN(n9228) );
  NAND2_X1 U7175 ( .A1(n9226), .A2(n6188), .ZN(n6207) );
  INV_X1 U7176 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8600) );
  INV_X1 U7177 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8356) );
  MUX2_X1 U7178 ( .A(n8600), .B(n8356), .S(n5680), .Z(n6191) );
  INV_X1 U7179 ( .A(SI_23_), .ZN(n10161) );
  NAND2_X1 U7180 ( .A1(n6191), .A2(n10161), .ZN(n6211) );
  INV_X1 U7181 ( .A(n6191), .ZN(n6192) );
  NAND2_X1 U7182 ( .A1(n6192), .A2(SI_23_), .ZN(n6193) );
  AND2_X1 U7183 ( .A1(n6211), .A2(n6193), .ZN(n6209) );
  NAND2_X1 U7184 ( .A1(n8599), .A2(n6421), .ZN(n6195) );
  OR2_X1 U7185 ( .A1(n5722), .A2(n8356), .ZN(n6194) );
  XNOR2_X1 U7186 ( .A(n9618), .B(n6214), .ZN(n6205) );
  XNOR2_X1 U7187 ( .A(n6207), .B(n6205), .ZN(n9172) );
  INV_X1 U7188 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10141) );
  NAND2_X1 U7189 ( .A1(n6196), .A2(n10141), .ZN(n6197) );
  NAND2_X1 U7190 ( .A1(n6215), .A2(n6197), .ZN(n9451) );
  OR2_X1 U7191 ( .A1(n9451), .A2(n6357), .ZN(n6203) );
  INV_X1 U7192 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U7193 ( .A1(n6403), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6199) );
  NAND2_X1 U7194 ( .A1(n6413), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6198) );
  OAI211_X1 U7195 ( .C1(n6200), .C2(n6360), .A(n6199), .B(n6198), .ZN(n6201)
         );
  INV_X1 U7196 ( .A(n6201), .ZN(n6202) );
  NAND2_X1 U7197 ( .A1(n9468), .A2(n9101), .ZN(n6204) );
  NAND2_X1 U7198 ( .A1(n9172), .A2(n6204), .ZN(n9178) );
  INV_X1 U7199 ( .A(n6205), .ZN(n6206) );
  NAND2_X1 U7200 ( .A1(n6207), .A2(n6206), .ZN(n6208) );
  NAND2_X1 U7201 ( .A1(n9178), .A2(n6208), .ZN(n6226) );
  MUX2_X1 U7202 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n5680), .Z(n6230) );
  INV_X1 U7203 ( .A(SI_24_), .ZN(n6232) );
  XNOR2_X1 U7204 ( .A(n6230), .B(n6232), .ZN(n6229) );
  XNOR2_X1 U7205 ( .A(n6234), .B(n6229), .ZN(n8688) );
  NAND2_X1 U7206 ( .A1(n8688), .A2(n6421), .ZN(n6213) );
  INV_X1 U7207 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8401) );
  OR2_X1 U7208 ( .A1(n5722), .A2(n8401), .ZN(n6212) );
  XNOR2_X1 U7209 ( .A(n9612), .B(n6214), .ZN(n6224) );
  XNOR2_X1 U7210 ( .A(n6226), .B(n6224), .ZN(n9205) );
  INV_X1 U7211 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10219) );
  NAND2_X1 U7212 ( .A1(n6215), .A2(n10219), .ZN(n6216) );
  AND2_X1 U7213 ( .A1(n6244), .A2(n6216), .ZN(n9430) );
  NAND2_X1 U7214 ( .A1(n9430), .A2(n6217), .ZN(n6223) );
  INV_X1 U7215 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7216 ( .A1(n6413), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U7217 ( .A1(n6403), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6218) );
  OAI211_X1 U7218 ( .C1(n6220), .C2(n6360), .A(n6219), .B(n6218), .ZN(n6221)
         );
  INV_X1 U7219 ( .A(n6221), .ZN(n6222) );
  NOR2_X1 U7220 ( .A1(n9197), .A2(n6628), .ZN(n9204) );
  NAND2_X1 U7221 ( .A1(n9205), .A2(n9204), .ZN(n6228) );
  INV_X1 U7222 ( .A(n6224), .ZN(n6225) );
  OR2_X1 U7223 ( .A1(n6226), .A2(n6225), .ZN(n6227) );
  INV_X1 U7224 ( .A(n6229), .ZN(n6233) );
  INV_X1 U7225 ( .A(n6230), .ZN(n6231) );
  INV_X1 U7226 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10260) );
  INV_X1 U7227 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8439) );
  MUX2_X1 U7228 ( .A(n10260), .B(n8439), .S(n5680), .Z(n6236) );
  INV_X1 U7229 ( .A(SI_25_), .ZN(n6235) );
  NAND2_X1 U7230 ( .A1(n6236), .A2(n6235), .ZN(n6256) );
  INV_X1 U7231 ( .A(n6236), .ZN(n6237) );
  NAND2_X1 U7232 ( .A1(n6237), .A2(SI_25_), .ZN(n6238) );
  NAND2_X1 U7233 ( .A1(n6256), .A2(n6238), .ZN(n6239) );
  NAND2_X1 U7234 ( .A1(n6240), .A2(n6239), .ZN(n6241) );
  NAND2_X1 U7235 ( .A1(n6257), .A2(n6241), .ZN(n8586) );
  NAND2_X1 U7236 ( .A1(n8586), .A2(n6421), .ZN(n6243) );
  OR2_X1 U7237 ( .A1(n5722), .A2(n8439), .ZN(n6242) );
  XNOR2_X1 U7238 ( .A(n9608), .B(n5047), .ZN(n6252) );
  INV_X1 U7239 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10213) );
  NAND2_X1 U7240 ( .A1(n6244), .A2(n10213), .ZN(n6245) );
  NAND2_X1 U7241 ( .A1(n6265), .A2(n6245), .ZN(n9415) );
  INV_X1 U7242 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n6248) );
  NAND2_X1 U7243 ( .A1(n6403), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U7244 ( .A1(n6413), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6246) );
  OAI211_X1 U7245 ( .C1(n6360), .C2(n6248), .A(n6247), .B(n6246), .ZN(n6249)
         );
  INV_X1 U7246 ( .A(n6249), .ZN(n6250) );
  NOR2_X1 U7247 ( .A1(n9437), .A2(n6628), .ZN(n6253) );
  XNOR2_X1 U7248 ( .A(n6252), .B(n6253), .ZN(n9195) );
  INV_X1 U7249 ( .A(n6252), .ZN(n6254) );
  NAND2_X1 U7250 ( .A1(n6254), .A2(n6253), .ZN(n6255) );
  INV_X1 U7251 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10576) );
  INV_X1 U7252 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9699) );
  MUX2_X1 U7253 ( .A(n10576), .B(n9699), .S(n5680), .Z(n6259) );
  INV_X1 U7254 ( .A(SI_26_), .ZN(n6258) );
  NAND2_X1 U7255 ( .A1(n6259), .A2(n6258), .ZN(n6278) );
  INV_X1 U7256 ( .A(n6259), .ZN(n6260) );
  NAND2_X1 U7257 ( .A1(n6260), .A2(SI_26_), .ZN(n6261) );
  AND2_X1 U7258 ( .A1(n6278), .A2(n6261), .ZN(n6276) );
  NAND2_X1 U7259 ( .A1(n9697), .A2(n6421), .ZN(n6263) );
  OR2_X1 U7260 ( .A1(n5722), .A2(n9699), .ZN(n6262) );
  NAND2_X2 U7261 ( .A1(n6263), .A2(n6262), .ZN(n9603) );
  XNOR2_X1 U7262 ( .A(n9603), .B(n6310), .ZN(n6273) );
  INV_X1 U7263 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6264) );
  NAND2_X1 U7264 ( .A1(n6265), .A2(n6264), .ZN(n6266) );
  NAND2_X1 U7265 ( .A1(n6288), .A2(n6266), .ZN(n9408) );
  INV_X1 U7266 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U7267 ( .A1(n6413), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6268) );
  NAND2_X1 U7268 ( .A1(n6403), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6267) );
  OAI211_X1 U7269 ( .C1(n6269), .C2(n6360), .A(n6268), .B(n6267), .ZN(n6270)
         );
  INV_X1 U7270 ( .A(n6270), .ZN(n6271) );
  NOR2_X1 U7271 ( .A1(n9198), .A2(n6628), .ZN(n6274) );
  XNOR2_X1 U7272 ( .A(n6273), .B(n6274), .ZN(n9254) );
  INV_X1 U7273 ( .A(n6273), .ZN(n6275) );
  INV_X1 U7274 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10253) );
  INV_X1 U7275 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6285) );
  MUX2_X1 U7276 ( .A(n10253), .B(n6285), .S(n5680), .Z(n6279) );
  INV_X1 U7277 ( .A(SI_27_), .ZN(n10154) );
  NAND2_X1 U7278 ( .A1(n6279), .A2(n10154), .ZN(n6314) );
  INV_X1 U7279 ( .A(n6279), .ZN(n6280) );
  NAND2_X1 U7280 ( .A1(n6280), .A2(SI_27_), .ZN(n6281) );
  AND2_X1 U7281 ( .A1(n6314), .A2(n6281), .ZN(n6282) );
  OR2_X1 U7282 ( .A1(n5722), .A2(n6285), .ZN(n6286) );
  XNOR2_X1 U7283 ( .A(n9597), .B(n5047), .ZN(n6294) );
  INV_X1 U7284 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9165) );
  NAND2_X1 U7285 ( .A1(n6288), .A2(n9165), .ZN(n6289) );
  INV_X1 U7286 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6292) );
  NAND2_X1 U7287 ( .A1(n6413), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U7288 ( .A1(n6403), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6290) );
  OAI211_X1 U7289 ( .C1(n6292), .C2(n6360), .A(n6291), .B(n6290), .ZN(n6293)
         );
  AOI21_X1 U7290 ( .B1(n9388), .B2(n5737), .A(n6293), .ZN(n9375) );
  NOR2_X1 U7291 ( .A1(n9375), .A2(n6628), .ZN(n6295) );
  XNOR2_X1 U7292 ( .A(n6294), .B(n6295), .ZN(n9164) );
  NAND2_X1 U7293 ( .A1(n9163), .A2(n9164), .ZN(n6298) );
  INV_X1 U7294 ( .A(n6294), .ZN(n6296) );
  NAND2_X1 U7295 ( .A1(n6296), .A2(n6295), .ZN(n6297) );
  INV_X1 U7296 ( .A(n6301), .ZN(n6299) );
  NAND2_X1 U7297 ( .A1(n6299), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n9084) );
  INV_X1 U7298 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U7299 ( .A1(n6301), .A2(n6300), .ZN(n6302) );
  NAND2_X1 U7300 ( .A1(n9084), .A2(n6302), .ZN(n6368) );
  INV_X1 U7301 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6305) );
  NAND2_X1 U7302 ( .A1(n6413), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6304) );
  NAND2_X1 U7303 ( .A1(n6403), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6303) );
  OAI211_X1 U7304 ( .C1(n6305), .C2(n6360), .A(n6304), .B(n6303), .ZN(n6306)
         );
  INV_X1 U7305 ( .A(n6306), .ZN(n6307) );
  NAND3_X1 U7306 ( .A1(n9393), .A2(n9101), .A3(n6310), .ZN(n6309) );
  OAI21_X1 U7307 ( .B1(n6310), .B2(n9393), .A(n6309), .ZN(n6311) );
  INV_X1 U7308 ( .A(n6311), .ZN(n6312) );
  MUX2_X1 U7309 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n5680), .Z(n6382) );
  XNOR2_X1 U7310 ( .A(n6382), .B(n10153), .ZN(n6380) );
  NAND2_X1 U7311 ( .A1(n9144), .A2(n6421), .ZN(n6317) );
  INV_X1 U7312 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9146) );
  OR2_X1 U7313 ( .A1(n5722), .A2(n9146), .ZN(n6316) );
  INV_X1 U7314 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10615) );
  NAND3_X1 U7315 ( .A1(n6322), .A2(n6325), .A3(n6327), .ZN(n6318) );
  NOR2_X1 U7316 ( .A1(n6319), .A2(n6318), .ZN(n6329) );
  INV_X1 U7317 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6330) );
  NAND2_X1 U7318 ( .A1(n6329), .A2(n6330), .ZN(n6332) );
  NAND2_X1 U7319 ( .A1(n6332), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6321) );
  INV_X1 U7320 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6320) );
  XNOR2_X1 U7321 ( .A(n6321), .B(n6320), .ZN(n9700) );
  NAND2_X1 U7322 ( .A1(n6323), .A2(n6322), .ZN(n6324) );
  NAND2_X1 U7323 ( .A1(n6324), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6353) );
  NAND2_X1 U7324 ( .A1(n6353), .A2(n6325), .ZN(n6326) );
  NAND2_X1 U7325 ( .A1(n6326), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6328) );
  XNOR2_X1 U7326 ( .A(n6328), .B(n6327), .ZN(n8403) );
  INV_X1 U7327 ( .A(n8403), .ZN(n6352) );
  INV_X1 U7328 ( .A(P2_B_REG_SCAN_IN), .ZN(n6334) );
  OR2_X1 U7329 ( .A1(n6329), .A2(n5651), .ZN(n6331) );
  MUX2_X1 U7330 ( .A(n6331), .B(P2_IR_REG_31__SCAN_IN), .S(n6330), .Z(n6333)
         );
  NAND2_X1 U7331 ( .A1(n6333), .A2(n6332), .ZN(n8437) );
  OAI221_X1 U7332 ( .B1(P2_B_REG_SCAN_IN), .B2(n6352), .C1(n6334), .C2(n8403), 
        .A(n8437), .ZN(n6335) );
  INV_X1 U7333 ( .A(n6335), .ZN(n6336) );
  AND2_X1 U7334 ( .A1(n8437), .A2(n9700), .ZN(n10616) );
  AOI21_X1 U7335 ( .B1(n10615), .B2(n6346), .A(n10616), .ZN(n7657) );
  NOR4_X1 U7336 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6345) );
  OR4_X1 U7337 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6342) );
  NOR4_X1 U7338 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6340) );
  NOR4_X1 U7339 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6339) );
  NOR4_X1 U7340 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6338) );
  NOR4_X1 U7341 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6337) );
  NAND4_X1 U7342 ( .A1(n6340), .A2(n6339), .A3(n6338), .A4(n6337), .ZN(n6341)
         );
  NOR4_X1 U7343 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        n6342), .A4(n6341), .ZN(n6344) );
  NOR4_X1 U7344 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6343) );
  NAND3_X1 U7345 ( .A1(n6345), .A2(n6344), .A3(n6343), .ZN(n6347) );
  NAND2_X1 U7346 ( .A1(n6347), .A2(n6346), .ZN(n7155) );
  AND2_X1 U7347 ( .A1(n8403), .A2(n9700), .ZN(n10695) );
  INV_X1 U7348 ( .A(n10695), .ZN(n6349) );
  OR2_X1 U7349 ( .A1(n10613), .A2(P2_D_REG_0__SCAN_IN), .ZN(n6348) );
  AND2_X1 U7350 ( .A1(n7155), .A2(n7288), .ZN(n6350) );
  NAND2_X1 U7351 ( .A1(n7657), .A2(n6350), .ZN(n6371) );
  NOR2_X1 U7352 ( .A1(n9700), .A2(n8437), .ZN(n6351) );
  NAND2_X1 U7353 ( .A1(n6352), .A2(n6351), .ZN(n6660) );
  XNOR2_X1 U7354 ( .A(n6353), .B(P2_IR_REG_23__SCAN_IN), .ZN(n6661) );
  NOR2_X1 U7355 ( .A1(n6661), .A2(P2_U3152), .ZN(n10694) );
  INV_X1 U7356 ( .A(n10614), .ZN(n7571) );
  OR2_X1 U7357 ( .A1(n10939), .A2(n6855), .ZN(n6356) );
  OR2_X1 U7358 ( .A1(n9084), .A2(n6357), .ZN(n6364) );
  INV_X1 U7359 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6361) );
  NAND2_X1 U7360 ( .A1(n6413), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6359) );
  NAND2_X1 U7361 ( .A1(n6403), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6358) );
  OAI211_X1 U7362 ( .C1(n6361), .C2(n6360), .A(n6359), .B(n6358), .ZN(n6362)
         );
  INV_X1 U7363 ( .A(n6362), .ZN(n6363) );
  INV_X1 U7364 ( .A(n9374), .ZN(n9264) );
  NOR2_X1 U7365 ( .A1(n6379), .A2(n6354), .ZN(n9257) );
  INV_X1 U7366 ( .A(n6855), .ZN(n7141) );
  INV_X1 U7367 ( .A(n6366), .ZN(n6367) );
  INV_X1 U7368 ( .A(n6368), .ZN(n9378) );
  OR3_X1 U7369 ( .A1(n6369), .A2(n6635), .A3(n9546), .ZN(n10750) );
  NOR2_X1 U7370 ( .A1(n10750), .A2(n6435), .ZN(n7152) );
  INV_X1 U7371 ( .A(n7152), .ZN(n6370) );
  NAND2_X1 U7372 ( .A1(n6371), .A2(n6370), .ZN(n6372) );
  NAND2_X1 U7373 ( .A1(n6354), .A2(n6855), .ZN(n7153) );
  NAND2_X1 U7374 ( .A1(n6372), .A2(n7153), .ZN(n7572) );
  INV_X1 U7375 ( .A(n6661), .ZN(n6373) );
  NAND2_X1 U7376 ( .A1(n6660), .A2(n6373), .ZN(n6374) );
  OR2_X1 U7377 ( .A1(n7572), .A2(n6374), .ZN(n6375) );
  AOI22_X1 U7378 ( .A1(n9264), .A2(n9244), .B1(n9378), .B2(n9246), .ZN(n6377)
         );
  INV_X1 U7379 ( .A(n9375), .ZN(n9265) );
  AOI22_X1 U7380 ( .A1(n9265), .A2(n9247), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n6376) );
  AND2_X1 U7381 ( .A1(n5698), .A2(n6369), .ZN(n10796) );
  INV_X1 U7382 ( .A(n10796), .ZN(n6378) );
  NAND2_X1 U7383 ( .A1(n10614), .A2(n7152), .ZN(n9549) );
  OAI21_X1 U7384 ( .B1(n6379), .B2(n6378), .A(n9549), .ZN(n9261) );
  INV_X1 U7385 ( .A(n9261), .ZN(n9099) );
  INV_X1 U7386 ( .A(n6382), .ZN(n6383) );
  MUX2_X1 U7387 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n5680), .Z(n6391) );
  INV_X1 U7388 ( .A(SI_29_), .ZN(n6384) );
  XNOR2_X1 U7389 ( .A(n6391), .B(n6384), .ZN(n6419) );
  MUX2_X1 U7390 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n5680), .Z(n6387) );
  INV_X1 U7391 ( .A(n6387), .ZN(n6385) );
  INV_X1 U7392 ( .A(SI_30_), .ZN(n6386) );
  NAND2_X1 U7393 ( .A1(n6385), .A2(n6386), .ZN(n6392) );
  INV_X1 U7394 ( .A(n6392), .ZN(n6388) );
  XNOR2_X1 U7395 ( .A(n6387), .B(n6386), .ZN(n6409) );
  OR2_X1 U7396 ( .A1(n6388), .A2(n6409), .ZN(n6390) );
  AND2_X1 U7397 ( .A1(n6419), .A2(n6390), .ZN(n6389) );
  NAND2_X1 U7398 ( .A1(n6420), .A2(n6389), .ZN(n6396) );
  INV_X1 U7399 ( .A(n6390), .ZN(n6394) );
  OR2_X1 U7400 ( .A1(n6391), .A2(SI_29_), .ZN(n6407) );
  AND2_X1 U7401 ( .A1(n6407), .A2(n6392), .ZN(n6393) );
  OR2_X1 U7402 ( .A1(n6394), .A2(n6393), .ZN(n6395) );
  MUX2_X1 U7403 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n5680), .Z(n6398) );
  INV_X1 U7404 ( .A(SI_31_), .ZN(n6397) );
  XNOR2_X1 U7405 ( .A(n6398), .B(n6397), .ZN(n6399) );
  NAND2_X1 U7406 ( .A1(n9687), .A2(n6421), .ZN(n6402) );
  INV_X1 U7407 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9689) );
  OR2_X1 U7408 ( .A1(n5722), .A2(n9689), .ZN(n6401) );
  NAND2_X1 U7409 ( .A1(n6403), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6406) );
  NAND2_X1 U7410 ( .A1(n6413), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6405) );
  NAND2_X1 U7411 ( .A1(n6414), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6404) );
  NAND3_X1 U7412 ( .A1(n6406), .A2(n6405), .A3(n6404), .ZN(n9360) );
  INV_X1 U7413 ( .A(n9360), .ZN(n6543) );
  OR2_X1 U7414 ( .A1(n9580), .A2(n6543), .ZN(n6418) );
  NAND2_X1 U7415 ( .A1(n6420), .A2(n6419), .ZN(n6408) );
  NAND2_X1 U7416 ( .A1(n6408), .A2(n6407), .ZN(n6410) );
  NAND2_X1 U7417 ( .A1(n9693), .A2(n6421), .ZN(n6412) );
  INV_X1 U7418 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9696) );
  OR2_X1 U7419 ( .A1(n5722), .A2(n9696), .ZN(n6411) );
  NAND2_X1 U7420 ( .A1(n6413), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6417) );
  NAND2_X1 U7421 ( .A1(n6403), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6416) );
  NAND2_X1 U7422 ( .A1(n6414), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6415) );
  AND3_X1 U7423 ( .A1(n6417), .A2(n6416), .A3(n6415), .ZN(n9094) );
  NAND2_X1 U7424 ( .A1(n9365), .A2(n9094), .ZN(n6539) );
  NOR2_X1 U7425 ( .A1(n9365), .A2(n9094), .ZN(n6620) );
  INV_X1 U7426 ( .A(n6620), .ZN(n6540) );
  AND2_X1 U7427 ( .A1(n6624), .A2(n6540), .ZN(n6548) );
  OR2_X1 U7428 ( .A1(n8174), .A2(n9546), .ZN(n7665) );
  MUX2_X1 U7429 ( .A(n6626), .B(n6548), .S(n6531), .Z(n6547) );
  NAND2_X1 U7430 ( .A1(n9060), .A2(n6421), .ZN(n6423) );
  INV_X1 U7431 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9061) );
  OR2_X1 U7432 ( .A1(n5722), .A2(n9061), .ZN(n6422) );
  NAND2_X1 U7433 ( .A1(n9083), .A2(n9374), .ZN(n6617) );
  NAND2_X1 U7434 ( .A1(n6549), .A2(n9399), .ZN(n6615) );
  NAND2_X1 U7435 ( .A1(n9603), .A2(n9198), .ZN(n6614) );
  NAND2_X1 U7436 ( .A1(n9608), .A2(n9437), .ZN(n6521) );
  NAND2_X1 U7437 ( .A1(n6614), .A2(n6521), .ZN(n6424) );
  MUX2_X1 U7438 ( .A(n6615), .B(n6424), .S(n6542), .Z(n6425) );
  INV_X1 U7439 ( .A(n6425), .ZN(n6530) );
  NAND2_X1 U7440 ( .A1(n9612), .A2(n9197), .ZN(n6550) );
  NAND2_X1 U7441 ( .A1(n9618), .A2(n9436), .ZN(n6611) );
  NAND2_X1 U7442 ( .A1(n6550), .A2(n6611), .ZN(n6427) );
  NAND2_X1 U7443 ( .A1(n6612), .A2(n6551), .ZN(n6426) );
  MUX2_X1 U7444 ( .A(n6427), .B(n6426), .S(n6542), .Z(n6428) );
  INV_X1 U7445 ( .A(n6428), .ZN(n6520) );
  NAND2_X1 U7446 ( .A1(n9074), .A2(n9485), .ZN(n6610) );
  INV_X1 U7447 ( .A(n6610), .ZN(n6430) );
  OAI21_X1 U7448 ( .B1(n9074), .B2(n9485), .A(n6611), .ZN(n6429) );
  MUX2_X1 U7449 ( .A(n6430), .B(n6429), .S(n6542), .Z(n6431) );
  INV_X1 U7450 ( .A(n6431), .ZN(n6518) );
  NAND2_X1 U7451 ( .A1(n9629), .A2(n9266), .ZN(n6607) );
  NAND2_X1 U7452 ( .A1(n6609), .A2(n6607), .ZN(n9475) );
  INV_X1 U7453 ( .A(n9475), .ZN(n9483) );
  NAND2_X1 U7454 ( .A1(n9634), .A2(n9510), .ZN(n6432) );
  MUX2_X1 U7455 ( .A(n6604), .B(n6432), .S(n6542), .Z(n6512) );
  NAND2_X1 U7456 ( .A1(n6604), .A2(n6432), .ZN(n9495) );
  INV_X1 U7457 ( .A(n9495), .ZN(n6606) );
  NAND2_X1 U7458 ( .A1(n9651), .A2(n9066), .ZN(n6499) );
  NAND2_X1 U7459 ( .A1(n6603), .A2(n6499), .ZN(n9542) );
  INV_X1 U7460 ( .A(n9542), .ZN(n6498) );
  NAND2_X1 U7461 ( .A1(n9655), .A2(n9540), .ZN(n6596) );
  MUX2_X1 U7462 ( .A(n6596), .B(n6600), .S(n6542), .Z(n6497) );
  NAND2_X1 U7463 ( .A1(n9659), .A2(n8422), .ZN(n6597) );
  MUX2_X1 U7464 ( .A(n8416), .B(n6597), .S(n6542), .Z(n6495) );
  INV_X1 U7465 ( .A(n10790), .ZN(n8781) );
  NAND2_X1 U7466 ( .A1(n8781), .A2(n10775), .ZN(n7772) );
  NAND2_X1 U7467 ( .A1(n9098), .A2(n9102), .ZN(n6439) );
  AND2_X1 U7468 ( .A1(n6439), .A2(n6435), .ZN(n6437) );
  OAI21_X1 U7469 ( .B1(n6441), .B2(n6437), .A(n6440), .ZN(n6443) );
  NAND2_X1 U7470 ( .A1(n6438), .A2(n6439), .ZN(n10743) );
  OAI21_X1 U7471 ( .B1(n7144), .B2(n10743), .A(n7713), .ZN(n6442) );
  MUX2_X1 U7472 ( .A(n6443), .B(n6442), .S(n6542), .Z(n6444) );
  INV_X1 U7473 ( .A(n7714), .ZN(n7712) );
  NAND2_X1 U7474 ( .A1(n6444), .A2(n7712), .ZN(n6448) );
  NAND2_X1 U7475 ( .A1(n9281), .A2(n10752), .ZN(n6446) );
  INV_X1 U7476 ( .A(n9281), .ZN(n7677) );
  NAND2_X1 U7477 ( .A1(n7677), .A2(n7728), .ZN(n6574) );
  MUX2_X1 U7478 ( .A(n6446), .B(n6574), .S(n6542), .Z(n6447) );
  NAND3_X1 U7479 ( .A1(n6448), .A2(n7669), .A3(n6447), .ZN(n6451) );
  MUX2_X1 U7480 ( .A(n6449), .B(n6575), .S(n6531), .Z(n6450) );
  NAND2_X1 U7481 ( .A1(n6451), .A2(n6450), .ZN(n6456) );
  INV_X1 U7482 ( .A(n10775), .ZN(n9214) );
  NAND3_X1 U7483 ( .A1(n6456), .A2(n10790), .A3(n9214), .ZN(n6453) );
  MUX2_X1 U7484 ( .A(n10790), .B(n9214), .S(n6542), .Z(n6452) );
  NAND2_X1 U7485 ( .A1(n6453), .A2(n6452), .ZN(n6455) );
  NAND2_X1 U7486 ( .A1(n9562), .A2(n10795), .ZN(n6579) );
  INV_X1 U7487 ( .A(n10795), .ZN(n10808) );
  INV_X1 U7488 ( .A(n9562), .ZN(n9279) );
  INV_X1 U7489 ( .A(n10787), .ZN(n6454) );
  OAI211_X1 U7490 ( .C1(n7772), .C2(n6456), .A(n6455), .B(n6454), .ZN(n6458)
         );
  MUX2_X1 U7491 ( .A(n6578), .B(n6579), .S(n6531), .Z(n6457) );
  NAND2_X1 U7492 ( .A1(n6458), .A2(n6457), .ZN(n6460) );
  NAND2_X1 U7493 ( .A1(n10821), .A2(n10792), .ZN(n7777) );
  MUX2_X1 U7494 ( .A(n10821), .B(n10792), .S(n6542), .Z(n6459) );
  OAI21_X1 U7495 ( .B1(n6460), .B2(n7777), .A(n6459), .ZN(n6462) );
  INV_X1 U7496 ( .A(n10821), .ZN(n7766) );
  INV_X1 U7497 ( .A(n10792), .ZN(n8777) );
  NAND3_X1 U7498 ( .A1(n6460), .A2(n7766), .A3(n8777), .ZN(n6461) );
  NAND2_X1 U7499 ( .A1(n6462), .A2(n6461), .ZN(n6464) );
  OR2_X1 U7500 ( .A1(n7813), .A2(n9560), .ZN(n6467) );
  NAND2_X1 U7501 ( .A1(n7813), .A2(n9560), .ZN(n6583) );
  OR2_X1 U7502 ( .A1(n7943), .A2(n7603), .ZN(n6465) );
  NAND2_X1 U7503 ( .A1(n7943), .A2(n7603), .ZN(n6585) );
  OAI21_X1 U7504 ( .B1(n6542), .B2(n6583), .A(n7779), .ZN(n6463) );
  AOI21_X1 U7505 ( .B1(n6464), .B2(n7807), .A(n6463), .ZN(n6472) );
  MUX2_X1 U7506 ( .A(n6585), .B(n6465), .S(n6531), .Z(n6466) );
  OR2_X1 U7507 ( .A1(n10863), .A2(n7986), .ZN(n6587) );
  NAND2_X1 U7508 ( .A1(n6466), .A2(n6587), .ZN(n6471) );
  NAND2_X1 U7509 ( .A1(n8029), .A2(n9239), .ZN(n6589) );
  NAND2_X1 U7510 ( .A1(n10863), .A2(n7986), .ZN(n6554) );
  INV_X1 U7511 ( .A(n6554), .ZN(n6473) );
  OR2_X1 U7512 ( .A1(n8029), .A2(n9239), .ZN(n6553) );
  OAI211_X1 U7513 ( .C1(n6467), .C2(n6471), .A(n6553), .B(n6587), .ZN(n6468)
         );
  MUX2_X1 U7514 ( .A(n6473), .B(n6468), .S(n6542), .Z(n6469) );
  INV_X1 U7515 ( .A(n6469), .ZN(n6470) );
  OAI211_X1 U7516 ( .C1(n6472), .C2(n6471), .A(n6589), .B(n6470), .ZN(n6479)
         );
  OR2_X1 U7517 ( .A1(n8095), .A2(n8559), .ZN(n6481) );
  NAND2_X1 U7518 ( .A1(n8095), .A2(n8559), .ZN(n6592) );
  NAND2_X1 U7519 ( .A1(n10901), .A2(n8075), .ZN(n6590) );
  NAND2_X1 U7520 ( .A1(n6553), .A2(n6473), .ZN(n6474) );
  NAND3_X1 U7521 ( .A1(n6590), .A2(n6589), .A3(n6474), .ZN(n6476) );
  OR2_X1 U7522 ( .A1(n10901), .A2(n8075), .ZN(n6552) );
  NAND2_X1 U7523 ( .A1(n6552), .A2(n6553), .ZN(n6475) );
  MUX2_X1 U7524 ( .A(n6476), .B(n6475), .S(n6531), .Z(n6477) );
  INV_X1 U7525 ( .A(n6477), .ZN(n6478) );
  NAND3_X1 U7526 ( .A1(n6479), .A2(n8081), .A3(n6478), .ZN(n6486) );
  XNOR2_X1 U7527 ( .A(n10938), .B(n8767), .ZN(n8098) );
  INV_X1 U7528 ( .A(n8098), .ZN(n6559) );
  NAND2_X1 U7529 ( .A1(n6481), .A2(n6552), .ZN(n6480) );
  NAND2_X1 U7530 ( .A1(n6480), .A2(n6592), .ZN(n6484) );
  NAND2_X1 U7531 ( .A1(n6592), .A2(n6590), .ZN(n6482) );
  NAND2_X1 U7532 ( .A1(n6482), .A2(n6481), .ZN(n6483) );
  MUX2_X1 U7533 ( .A(n6484), .B(n6483), .S(n6531), .Z(n6485) );
  NAND3_X1 U7534 ( .A1(n6486), .A2(n6559), .A3(n6485), .ZN(n6490) );
  NAND2_X1 U7535 ( .A1(n9664), .A2(n9052), .ZN(n6491) );
  OR2_X1 U7536 ( .A1(n8767), .A2(n6542), .ZN(n6488) );
  NAND2_X1 U7537 ( .A1(n8767), .A2(n6542), .ZN(n6487) );
  MUX2_X1 U7538 ( .A(n6488), .B(n6487), .S(n10938), .Z(n6489) );
  NAND3_X1 U7539 ( .A1(n6490), .A2(n8360), .A3(n6489), .ZN(n6493) );
  MUX2_X1 U7540 ( .A(n6594), .B(n6491), .S(n6531), .Z(n6492) );
  NAND3_X1 U7541 ( .A1(n6493), .A2(n8445), .A3(n6492), .ZN(n6494) );
  NAND3_X1 U7542 ( .A1(n6495), .A2(n8424), .A3(n6494), .ZN(n6496) );
  NAND3_X1 U7543 ( .A1(n6498), .A2(n6497), .A3(n6496), .ZN(n6501) );
  MUX2_X1 U7544 ( .A(n6499), .B(n6603), .S(n6531), .Z(n6500) );
  NAND2_X1 U7545 ( .A1(n6501), .A2(n6500), .ZN(n6505) );
  XNOR2_X1 U7546 ( .A(n9644), .B(n9539), .ZN(n9525) );
  INV_X1 U7547 ( .A(n9539), .ZN(n9268) );
  NAND2_X1 U7548 ( .A1(n9268), .A2(n6542), .ZN(n6503) );
  NAND2_X1 U7549 ( .A1(n9539), .A2(n6531), .ZN(n6502) );
  MUX2_X1 U7550 ( .A(n6503), .B(n6502), .S(n9644), .Z(n6504) );
  OAI21_X1 U7551 ( .B1(n6505), .B2(n9525), .A(n6504), .ZN(n6509) );
  XNOR2_X1 U7552 ( .A(n9641), .B(n9068), .ZN(n9507) );
  INV_X1 U7553 ( .A(n9068), .ZN(n9528) );
  NAND2_X1 U7554 ( .A1(n9528), .A2(n6531), .ZN(n6507) );
  NAND2_X1 U7555 ( .A1(n9068), .A2(n6542), .ZN(n6506) );
  MUX2_X1 U7556 ( .A(n6507), .B(n6506), .S(n9641), .Z(n6508) );
  OAI21_X1 U7557 ( .B1(n6509), .B2(n9507), .A(n6508), .ZN(n6510) );
  NAND2_X1 U7558 ( .A1(n6606), .A2(n6510), .ZN(n6511) );
  NAND2_X1 U7559 ( .A1(n6512), .A2(n6511), .ZN(n6513) );
  NAND2_X1 U7560 ( .A1(n9483), .A2(n6513), .ZN(n6515) );
  MUX2_X1 U7561 ( .A(n6609), .B(n6607), .S(n6542), .Z(n6514) );
  NAND2_X1 U7562 ( .A1(n6515), .A2(n6514), .ZN(n6516) );
  NAND2_X1 U7563 ( .A1(n6516), .A2(n9466), .ZN(n6517) );
  NAND3_X1 U7564 ( .A1(n6518), .A2(n6551), .A3(n6517), .ZN(n6519) );
  NAND2_X1 U7565 ( .A1(n6520), .A2(n6519), .ZN(n6522) );
  INV_X1 U7566 ( .A(n9612), .ZN(n9432) );
  AOI21_X1 U7567 ( .B1(n6522), .B2(n9432), .A(n9420), .ZN(n6525) );
  AND2_X1 U7568 ( .A1(n6521), .A2(n6531), .ZN(n6524) );
  OAI211_X1 U7569 ( .C1(n9445), .C2(n6531), .A(n6522), .B(n6612), .ZN(n6523)
         );
  OAI21_X1 U7570 ( .B1(n6525), .B2(n6524), .A(n6523), .ZN(n6529) );
  INV_X1 U7571 ( .A(n6614), .ZN(n6527) );
  INV_X1 U7572 ( .A(n6549), .ZN(n6526) );
  MUX2_X1 U7573 ( .A(n6527), .B(n6526), .S(n6542), .Z(n6528) );
  AOI21_X1 U7574 ( .B1(n6530), .B2(n6529), .A(n6528), .ZN(n6534) );
  NAND2_X1 U7575 ( .A1(n9597), .A2(n9375), .ZN(n6532) );
  MUX2_X1 U7576 ( .A(n6616), .B(n6532), .S(n6531), .Z(n6533) );
  OAI211_X1 U7577 ( .C1(n6534), .C2(n9080), .A(n9082), .B(n6533), .ZN(n6537)
         );
  INV_X1 U7578 ( .A(n9393), .ZN(n9166) );
  OR3_X1 U7579 ( .A1(n9592), .A2(n9166), .A3(n6542), .ZN(n6536) );
  NAND3_X1 U7580 ( .A1(n9592), .A2(n9166), .A3(n6542), .ZN(n6535) );
  NAND4_X1 U7581 ( .A1(n9088), .A2(n6537), .A3(n6536), .A4(n6535), .ZN(n6541)
         );
  MUX2_X1 U7582 ( .A(n6617), .B(n6618), .S(n6542), .Z(n6538) );
  NAND4_X1 U7583 ( .A1(n6541), .A2(n6540), .A3(n6539), .A4(n6538), .ZN(n6546)
         );
  AOI21_X1 U7584 ( .B1(n9580), .B2(n9360), .A(n6544), .ZN(n6545) );
  INV_X1 U7585 ( .A(n6548), .ZN(n6569) );
  INV_X1 U7586 ( .A(n6626), .ZN(n6568) );
  NAND2_X1 U7587 ( .A1(n6552), .A2(n6590), .ZN(n8032) );
  INV_X1 U7588 ( .A(n8032), .ZN(n8034) );
  NAND2_X1 U7589 ( .A1(n6553), .A2(n6589), .ZN(n7983) );
  NOR2_X1 U7590 ( .A1(n7144), .A2(n8063), .ZN(n6555) );
  INV_X1 U7591 ( .A(n10743), .ZN(n7741) );
  NAND4_X1 U7592 ( .A1(n6555), .A2(n7669), .A3(n7741), .A4(n7712), .ZN(n6556)
         );
  NOR3_X1 U7593 ( .A1(n6556), .A2(n7750), .A3(n10787), .ZN(n6557) );
  XNOR2_X1 U7594 ( .A(n10821), .B(n10792), .ZN(n9571) );
  AND4_X1 U7595 ( .A1(n7948), .A2(n7807), .A3(n6557), .A4(n9571), .ZN(n6558)
         );
  AND4_X1 U7596 ( .A1(n8081), .A2(n6588), .A3(n7779), .A4(n6558), .ZN(n6560)
         );
  AND4_X1 U7597 ( .A1(n8360), .A2(n8034), .A3(n6560), .A4(n6559), .ZN(n6561)
         );
  NAND3_X1 U7598 ( .A1(n8424), .A2(n8445), .A3(n6561), .ZN(n6562) );
  NOR4_X1 U7599 ( .A1(n9495), .A2(n9525), .A3(n9542), .A4(n6562), .ZN(n6564)
         );
  INV_X1 U7600 ( .A(n9507), .ZN(n6563) );
  NAND4_X1 U7601 ( .A1(n9466), .A2(n9483), .A3(n6564), .A4(n6563), .ZN(n6565)
         );
  NOR4_X1 U7602 ( .A1(n9420), .A2(n9435), .A3(n9443), .A4(n6565), .ZN(n6566)
         );
  NAND4_X1 U7603 ( .A1(n9088), .A2(n5143), .A3(n9401), .A4(n6566), .ZN(n6567)
         );
  XNOR2_X1 U7604 ( .A(n6570), .B(n9546), .ZN(n6571) );
  NAND2_X1 U7605 ( .A1(n6635), .A2(n10800), .ZN(n7146) );
  INV_X1 U7606 ( .A(n6575), .ZN(n6576) );
  INV_X1 U7607 ( .A(n7750), .ZN(n7743) );
  NAND2_X1 U7608 ( .A1(n7744), .A2(n7743), .ZN(n7742) );
  NAND2_X1 U7609 ( .A1(n10790), .A2(n10775), .ZN(n6577) );
  INV_X1 U7610 ( .A(n6578), .ZN(n6580) );
  NAND2_X1 U7611 ( .A1(n7766), .A2(n10792), .ZN(n6581) );
  NAND2_X1 U7612 ( .A1(n10821), .A2(n8777), .ZN(n6582) );
  NAND2_X1 U7613 ( .A1(n7803), .A2(n7807), .ZN(n6584) );
  NAND2_X1 U7614 ( .A1(n6584), .A2(n6583), .ZN(n7763) );
  INV_X1 U7615 ( .A(n6585), .ZN(n6586) );
  NAND2_X1 U7616 ( .A1(n7949), .A2(n7948), .ZN(n7947) );
  NAND2_X1 U7617 ( .A1(n6591), .A2(n6590), .ZN(n8073) );
  INV_X1 U7618 ( .A(n6592), .ZN(n6593) );
  INV_X1 U7619 ( .A(n8767), .ZN(n9272) );
  INV_X1 U7620 ( .A(n8360), .ZN(n8364) );
  INV_X1 U7621 ( .A(n6594), .ZN(n6595) );
  INV_X1 U7622 ( .A(n6596), .ZN(n6599) );
  INV_X1 U7623 ( .A(n6597), .ZN(n6598) );
  INV_X1 U7624 ( .A(n6600), .ZN(n6601) );
  NOR2_X1 U7625 ( .A1(n6602), .A2(n6601), .ZN(n9536) );
  INV_X1 U7626 ( .A(n9525), .ZN(n9517) );
  INV_X1 U7627 ( .A(n9644), .ZN(n9524) );
  INV_X1 U7628 ( .A(n6604), .ZN(n6605) );
  INV_X1 U7629 ( .A(n6607), .ZN(n6608) );
  NAND2_X1 U7630 ( .A1(n9467), .A2(n9466), .ZN(n9465) );
  NAND2_X1 U7631 ( .A1(n9465), .A2(n6610), .ZN(n9444) );
  INV_X1 U7632 ( .A(n6612), .ZN(n6613) );
  INV_X1 U7633 ( .A(n6621), .ZN(n6623) );
  OAI21_X1 U7634 ( .B1(n6621), .B2(n6620), .A(n6619), .ZN(n6622) );
  OAI21_X1 U7635 ( .B1(n6623), .B2(n9365), .A(n6622), .ZN(n6627) );
  AOI21_X1 U7636 ( .B1(n6627), .B2(n6626), .A(n6625), .ZN(n6632) );
  INV_X1 U7637 ( .A(n7147), .ZN(n6629) );
  AOI21_X1 U7638 ( .B1(n6629), .B2(n9546), .A(n6628), .ZN(n6630) );
  INV_X1 U7639 ( .A(n6630), .ZN(n6631) );
  NAND2_X1 U7640 ( .A1(n6661), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8354) );
  NOR4_X1 U7641 ( .A1(n7571), .A2(n6354), .A3(n9091), .A4(n9561), .ZN(n6637)
         );
  OAI21_X1 U7642 ( .B1(n8354), .B2(n6635), .A(P2_B_REG_SCAN_IN), .ZN(n6636) );
  OR2_X1 U7643 ( .A1(n6637), .A2(n6636), .ZN(n6638) );
  NAND2_X1 U7644 ( .A1(n6677), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6647) );
  NAND2_X1 U7645 ( .A1(n6647), .A2(n6678), .ZN(n6650) );
  OR2_X1 U7646 ( .A1(n6647), .A2(n6678), .ZN(n6648) );
  NAND2_X1 U7647 ( .A1(n6650), .A2(n6648), .ZN(n8436) );
  NOR2_X1 U7648 ( .A1(n8436), .A2(n8400), .ZN(n6652) );
  INV_X1 U7649 ( .A(n6669), .ZN(n6655) );
  NAND2_X1 U7650 ( .A1(n5122), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6657) );
  XNOR2_X1 U7651 ( .A(n6657), .B(n6656), .ZN(n8351) );
  INV_X1 U7652 ( .A(n8351), .ZN(n6658) );
  NOR2_X1 U7653 ( .A1(n7208), .A2(n6658), .ZN(n6780) );
  AND2_X2 U7654 ( .A1(n6780), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  OR2_X1 U7655 ( .A1(n6660), .A2(P2_U3152), .ZN(n6989) );
  INV_X2 U7656 ( .A(n9267), .ZN(P2_U3966) );
  INV_X1 U7657 ( .A(n8406), .ZN(n6662) );
  AOI211_X1 U7658 ( .C1(n6664), .C2(n6663), .A(n5042), .B(n6662), .ZN(n6668)
         );
  INV_X1 U7659 ( .A(n9651), .ZN(n9548) );
  NOR2_X1 U7660 ( .A1(n9548), .A2(n9099), .ZN(n6667) );
  OAI22_X1 U7661 ( .A1(n9229), .A2(n9539), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9319), .ZN(n6666) );
  OAI22_X1 U7662 ( .A1(n9230), .A2(n9540), .B1(n9259), .B2(n9550), .ZN(n6665)
         );
  OR4_X1 U7663 ( .A1(n6668), .A2(n6667), .A3(n6666), .A4(n6665), .ZN(P2_U3230)
         );
  NAND2_X1 U7664 ( .A1(n6669), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6929) );
  NAND2_X1 U7665 ( .A1(n6929), .A2(n6928), .ZN(n6670) );
  NAND2_X1 U7666 ( .A1(n6670), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6673) );
  NAND2_X1 U7667 ( .A1(n6673), .A2(n6672), .ZN(n6675) );
  NAND2_X1 U7668 ( .A1(n6675), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6671) );
  OR2_X1 U7669 ( .A1(n6673), .A2(n6672), .ZN(n6674) );
  NAND2_X1 U7670 ( .A1(n7208), .A2(n7205), .ZN(n6676) );
  NAND2_X1 U7671 ( .A1(n6676), .A2(n8351), .ZN(n6752) );
  INV_X1 U7672 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6679) );
  NAND2_X1 U7673 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n6680) );
  INV_X1 U7674 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6803) );
  NAND2_X1 U7675 ( .A1(n6752), .A2(n7510), .ZN(n6777) );
  NAND2_X1 U7676 ( .A1(n6777), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  OR2_X1 U7677 ( .A1(n6682), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n6688) );
  NAND2_X1 U7678 ( .A1(n6688), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6683) );
  MUX2_X1 U7679 ( .A(n6683), .B(P1_IR_REG_31__SCAN_IN), .S(n10319), .Z(n6685)
         );
  INV_X1 U7680 ( .A(n6688), .ZN(n6684) );
  NAND2_X1 U7681 ( .A1(n6684), .A2(n10319), .ZN(n6749) );
  NAND2_X1 U7682 ( .A1(n6685), .A2(n6749), .ZN(n8183) );
  INV_X1 U7683 ( .A(n8183), .ZN(n8462) );
  NAND2_X1 U7684 ( .A1(n6682), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6687) );
  MUX2_X1 U7685 ( .A(n6687), .B(P1_IR_REG_31__SCAN_IN), .S(n6686), .Z(n6689)
         );
  NAND2_X1 U7686 ( .A1(n6689), .A2(n6688), .ZN(n8373) );
  NAND2_X1 U7687 ( .A1(n6690), .A2(n6691), .ZN(n6722) );
  NOR2_X1 U7688 ( .A1(n6722), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n6712) );
  NOR2_X1 U7689 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n6692) );
  NAND2_X1 U7690 ( .A1(n6712), .A2(n6692), .ZN(n6708) );
  INV_X1 U7691 ( .A(n6693), .ZN(n6694) );
  OAI21_X1 U7692 ( .B1(n6708), .B2(n6694), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6695) );
  MUX2_X1 U7693 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6695), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n6696) );
  AND2_X1 U7694 ( .A1(n6682), .A2(n6696), .ZN(n8243) );
  OAI21_X1 U7695 ( .B1(n6742), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6698) );
  INV_X1 U7696 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10310) );
  NAND2_X1 U7697 ( .A1(n6698), .A2(n10310), .ZN(n6699) );
  NAND2_X1 U7698 ( .A1(n6699), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6697) );
  XNOR2_X1 U7699 ( .A(n6697), .B(P1_IR_REG_13__SCAN_IN), .ZN(n8235) );
  NAND2_X1 U7700 ( .A1(n8235), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6746) );
  OR2_X1 U7701 ( .A1(n6698), .A2(n10310), .ZN(n6700) );
  NAND2_X1 U7702 ( .A1(n6706), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6701) );
  MUX2_X1 U7703 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6701), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n6702) );
  NAND2_X1 U7704 ( .A1(n6702), .A2(n6742), .ZN(n6910) );
  INV_X1 U7705 ( .A(n6910), .ZN(n10662) );
  NAND2_X1 U7706 ( .A1(n10662), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6741) );
  INV_X1 U7707 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6703) );
  MUX2_X1 U7708 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n6703), .S(n6910), .Z(n6704)
         );
  INV_X1 U7709 ( .A(n6704), .ZN(n10669) );
  NAND2_X1 U7710 ( .A1(n6710), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6705) );
  MUX2_X1 U7711 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6705), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n6707) );
  AND2_X1 U7712 ( .A1(n6707), .A2(n6706), .ZN(n7860) );
  INV_X1 U7713 ( .A(n7860), .ZN(n6924) );
  INV_X1 U7714 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6740) );
  NAND2_X1 U7715 ( .A1(n6708), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6709) );
  MUX2_X1 U7716 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6709), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n6711) );
  AND2_X1 U7717 ( .A1(n6711), .A2(n6710), .ZN(n7820) );
  INV_X1 U7718 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7892) );
  OR2_X1 U7719 ( .A1(n6712), .A2(n10563), .ZN(n6714) );
  INV_X1 U7720 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n10300) );
  NAND2_X1 U7721 ( .A1(n6714), .A2(n10300), .ZN(n6716) );
  NAND2_X1 U7722 ( .A1(n6716), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6713) );
  XNOR2_X1 U7723 ( .A(n6713), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7511) );
  NOR2_X1 U7724 ( .A1(n7511), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6739) );
  OR2_X1 U7725 ( .A1(n6714), .A2(n10300), .ZN(n6715) );
  NAND2_X1 U7726 ( .A1(n6842), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6738) );
  INV_X1 U7727 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6717) );
  INV_X1 U7728 ( .A(n6842), .ZN(n7440) );
  AOI22_X1 U7729 ( .A1(n6842), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n6717), .B2(
        n7440), .ZN(n6836) );
  NAND2_X1 U7730 ( .A1(n6722), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6719) );
  XNOR2_X1 U7731 ( .A(n6719), .B(n6718), .ZN(n7344) );
  INV_X1 U7732 ( .A(n7344), .ZN(n6899) );
  NOR2_X1 U7733 ( .A1(n6899), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6737) );
  NOR2_X1 U7734 ( .A1(n6690), .A2(n10563), .ZN(n6720) );
  MUX2_X1 U7735 ( .A(n10563), .B(n6720), .S(P1_IR_REG_4__SCAN_IN), .Z(n6721)
         );
  INV_X1 U7736 ( .A(n6721), .ZN(n6723) );
  NAND2_X1 U7737 ( .A1(n6723), .A2(n6722), .ZN(n7247) );
  INV_X1 U7738 ( .A(n7247), .ZN(n6969) );
  NOR2_X1 U7739 ( .A1(n6969), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6735) );
  INV_X1 U7740 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7417) );
  OR2_X1 U7741 ( .A1(n6724), .A2(n10563), .ZN(n6732) );
  INV_X1 U7742 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6731) );
  NAND2_X1 U7743 ( .A1(n6732), .A2(n6731), .ZN(n6725) );
  NAND2_X1 U7744 ( .A1(n6725), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6726) );
  INV_X1 U7745 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n10294) );
  XNOR2_X1 U7746 ( .A(n6726), .B(n10294), .ZN(n9850) );
  INV_X1 U7747 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6729) );
  INV_X1 U7748 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n6728) );
  NAND2_X1 U7749 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6727) );
  XNOR2_X1 U7750 ( .A(n6728), .B(n6727), .ZN(n10676) );
  MUX2_X1 U7751 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6729), .S(n10676), .Z(n6730)
         );
  INV_X1 U7752 ( .A(n6730), .ZN(n10682) );
  NAND3_X1 U7753 ( .A1(n10682), .A2(P1_REG2_REG_0__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n10680) );
  INV_X1 U7754 ( .A(n10676), .ZN(n6758) );
  NAND2_X1 U7755 ( .A1(n6758), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9838) );
  INV_X1 U7756 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7428) );
  XNOR2_X1 U7757 ( .A(n6732), .B(n6731), .ZN(n7109) );
  MUX2_X1 U7758 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n7428), .S(n7109), .Z(n9837)
         );
  AOI21_X1 U7759 ( .B1(n10680), .B2(n9838), .A(n9837), .ZN(n9853) );
  NOR2_X1 U7760 ( .A1(n7109), .A2(n7428), .ZN(n9852) );
  MUX2_X1 U7761 ( .A(n7417), .B(P1_REG2_REG_3__SCAN_IN), .S(n9850), .Z(n9854)
         );
  OAI21_X1 U7762 ( .B1(n9853), .B2(n9852), .A(n9854), .ZN(n9856) );
  OAI21_X1 U7763 ( .B1(n7417), .B2(n9850), .A(n9856), .ZN(n6968) );
  INV_X1 U7764 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6734) );
  INV_X1 U7765 ( .A(n6735), .ZN(n6733) );
  OAI21_X1 U7766 ( .B1(n6734), .B2(n7247), .A(n6733), .ZN(n6967) );
  NOR2_X1 U7767 ( .A1(n6968), .A2(n6967), .ZN(n6966) );
  NOR2_X1 U7768 ( .A1(n6735), .A2(n6966), .ZN(n6895) );
  INV_X1 U7769 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7551) );
  INV_X1 U7770 ( .A(n6737), .ZN(n6736) );
  OAI21_X1 U7771 ( .B1(n7551), .B2(n7344), .A(n6736), .ZN(n6896) );
  NOR2_X1 U7772 ( .A1(n6895), .A2(n6896), .ZN(n6894) );
  NOR2_X1 U7773 ( .A1(n6737), .A2(n6894), .ZN(n6835) );
  NAND2_X1 U7774 ( .A1(n6836), .A2(n6835), .ZN(n6834) );
  NAND2_X1 U7775 ( .A1(n6738), .A2(n6834), .ZN(n6861) );
  INV_X1 U7776 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7535) );
  INV_X1 U7777 ( .A(n7511), .ZN(n6863) );
  AOI22_X1 U7778 ( .A1(n7511), .A2(n7535), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n6863), .ZN(n6860) );
  NOR2_X1 U7779 ( .A1(n6861), .A2(n6860), .ZN(n6859) );
  NOR2_X1 U7780 ( .A1(n6739), .A2(n6859), .ZN(n6879) );
  MUX2_X1 U7781 ( .A(n7892), .B(P1_REG2_REG_8__SCAN_IN), .S(n7820), .Z(n6878)
         );
  OAI21_X1 U7782 ( .B1(n7820), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6876), .ZN(
        n6916) );
  MUX2_X1 U7783 ( .A(n6740), .B(P1_REG2_REG_9__SCAN_IN), .S(n7860), .Z(n6915)
         );
  OAI21_X1 U7784 ( .B1(n6924), .B2(n6740), .A(n6913), .ZN(n10670) );
  NAND2_X1 U7785 ( .A1(n10669), .A2(n10670), .ZN(n10668) );
  NAND2_X1 U7786 ( .A1(n6741), .A2(n10668), .ZN(n7308) );
  AND2_X1 U7787 ( .A1(n7308), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7302) );
  NAND2_X1 U7788 ( .A1(n6742), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6743) );
  XNOR2_X1 U7789 ( .A(n6743), .B(P1_IR_REG_11__SCAN_IN), .ZN(n8016) );
  OAI22_X1 U7790 ( .A1(n7302), .A2(n8016), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n7308), .ZN(n7406) );
  NAND2_X1 U7791 ( .A1(n8128), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6744) );
  OAI21_X1 U7792 ( .B1(n8128), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6744), .ZN(
        n7405) );
  NOR2_X1 U7793 ( .A1(n7406), .A2(n7405), .ZN(n7404) );
  AOI21_X1 U7794 ( .B1(n8128), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7404), .ZN(
        n7635) );
  OAI21_X1 U7795 ( .B1(n8235), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6746), .ZN(
        n7634) );
  NOR2_X1 U7796 ( .A1(n7635), .A2(n7634), .ZN(n7633) );
  INV_X1 U7797 ( .A(n7633), .ZN(n6745) );
  NAND2_X1 U7798 ( .A1(n6746), .A2(n6745), .ZN(n7613) );
  XNOR2_X1 U7799 ( .A(n8243), .B(P1_REG2_REG_14__SCAN_IN), .ZN(n7612) );
  OAI21_X1 U7800 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n8243), .A(n7615), .ZN(
        n6747) );
  NOR2_X1 U7801 ( .A1(n8373), .A2(n6747), .ZN(n6748) );
  INV_X1 U7802 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8067) );
  XNOR2_X1 U7803 ( .A(n6747), .B(n8373), .ZN(n8068) );
  NOR2_X1 U7804 ( .A1(n8067), .A2(n8068), .ZN(n8066) );
  NOR2_X1 U7805 ( .A1(n6748), .A2(n8066), .ZN(n8178) );
  XNOR2_X1 U7806 ( .A(n8462), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n8177) );
  NOR2_X1 U7807 ( .A1(n8178), .A2(n8177), .ZN(n8176) );
  AOI21_X1 U7808 ( .B1(n8462), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8176), .ZN(
        n6755) );
  NAND2_X1 U7809 ( .A1(n6749), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7850) );
  XNOR2_X1 U7810 ( .A(n7850), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9868) );
  NAND2_X1 U7811 ( .A1(n9868), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6750) );
  OAI21_X1 U7812 ( .B1(n9868), .B2(P1_REG2_REG_17__SCAN_IN), .A(n6750), .ZN(
        n6754) );
  NOR2_X1 U7813 ( .A1(n5050), .A2(P1_U3084), .ZN(n10570) );
  NAND2_X1 U7814 ( .A1(n6752), .A2(n10570), .ZN(n7298) );
  OR2_X1 U7815 ( .A1(n7298), .A2(n6753), .ZN(n9890) );
  NOR2_X1 U7816 ( .A1(n6755), .A2(n6754), .ZN(n9867) );
  AOI211_X1 U7817 ( .C1(n6755), .C2(n6754), .A(n9890), .B(n9867), .ZN(n6785)
         );
  INV_X1 U7818 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6756) );
  MUX2_X1 U7819 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n6756), .S(n8235), .Z(n7629)
         );
  NOR2_X1 U7820 ( .A1(n7511), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6764) );
  NAND2_X1 U7821 ( .A1(n6842), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6763) );
  INV_X1 U7822 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6757) );
  MUX2_X1 U7823 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6757), .S(n6842), .Z(n6838)
         );
  INV_X1 U7824 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6762) );
  MUX2_X1 U7825 ( .A(n6762), .B(P1_REG1_REG_5__SCAN_IN), .S(n7344), .Z(n6901)
         );
  INV_X1 U7826 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6761) );
  INV_X1 U7827 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6760) );
  XOR2_X1 U7828 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10676), .Z(n10687) );
  NAND2_X1 U7829 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n10686) );
  NOR2_X1 U7830 ( .A1(n10687), .A2(n10686), .ZN(n10685) );
  AOI21_X1 U7831 ( .B1(n6758), .B2(P1_REG1_REG_1__SCAN_IN), .A(n10685), .ZN(
        n9835) );
  INV_X1 U7832 ( .A(n9835), .ZN(n6759) );
  XNOR2_X1 U7833 ( .A(n7109), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9834) );
  INV_X1 U7834 ( .A(n7109), .ZN(n9833) );
  AOI22_X1 U7835 ( .A1(n6759), .A2(n9834), .B1(P1_REG1_REG_2__SCAN_IN), .B2(
        n9833), .ZN(n9848) );
  MUX2_X1 U7836 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6760), .S(n9850), .Z(n9847)
         );
  OR2_X1 U7837 ( .A1(n9848), .A2(n9847), .ZN(n9845) );
  OAI21_X1 U7838 ( .B1(n6760), .B2(n9850), .A(n9845), .ZN(n6974) );
  MUX2_X1 U7839 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6761), .S(n7247), .Z(n6973)
         );
  NOR2_X1 U7840 ( .A1(n6974), .A2(n6973), .ZN(n6972) );
  AOI21_X1 U7841 ( .B1(n7247), .B2(n6761), .A(n6972), .ZN(n6902) );
  NAND2_X1 U7842 ( .A1(n6901), .A2(n6902), .ZN(n6900) );
  OAI21_X1 U7843 ( .B1(n6762), .B2(n7344), .A(n6900), .ZN(n6839) );
  NAND2_X1 U7844 ( .A1(n6838), .A2(n6839), .ZN(n6837) );
  NAND2_X1 U7845 ( .A1(n6763), .A2(n6837), .ZN(n6866) );
  INV_X1 U7846 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7709) );
  AOI22_X1 U7847 ( .A1(n7511), .A2(n7709), .B1(P1_REG1_REG_7__SCAN_IN), .B2(
        n6863), .ZN(n6865) );
  NOR2_X1 U7848 ( .A1(n6866), .A2(n6865), .ZN(n6864) );
  NOR2_X1 U7849 ( .A1(n6764), .A2(n6864), .ZN(n6883) );
  INV_X1 U7850 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6765) );
  MUX2_X1 U7851 ( .A(n6765), .B(P1_REG1_REG_8__SCAN_IN), .S(n7820), .Z(n6882)
         );
  OR2_X1 U7852 ( .A1(n7820), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6918) );
  NAND2_X1 U7853 ( .A1(n6920), .A2(n6918), .ZN(n6766) );
  INV_X1 U7854 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10859) );
  MUX2_X1 U7855 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10859), .S(n7860), .Z(n6917)
         );
  NAND2_X1 U7856 ( .A1(n6766), .A2(n6917), .ZN(n6922) );
  NAND2_X1 U7857 ( .A1(n6924), .A2(n10859), .ZN(n6767) );
  NAND2_X1 U7858 ( .A1(n6922), .A2(n6767), .ZN(n10664) );
  INV_X1 U7859 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10880) );
  MUX2_X1 U7860 ( .A(n10880), .B(P1_REG1_REG_10__SCAN_IN), .S(n6910), .Z(
        n10665) );
  NAND2_X1 U7861 ( .A1(n10664), .A2(n10665), .ZN(n10663) );
  NAND2_X1 U7862 ( .A1(n6910), .A2(n10880), .ZN(n6768) );
  NAND2_X1 U7863 ( .A1(n10663), .A2(n6768), .ZN(n7303) );
  INV_X1 U7864 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10897) );
  NOR2_X1 U7865 ( .A1(n7303), .A2(n10897), .ZN(n6770) );
  INV_X1 U7866 ( .A(n7303), .ZN(n6769) );
  OAI22_X1 U7867 ( .A1(n6770), .A2(n8016), .B1(n6769), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7400) );
  INV_X1 U7868 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6771) );
  MUX2_X1 U7869 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6771), .S(n8128), .Z(n7401)
         );
  NAND2_X1 U7870 ( .A1(n7400), .A2(n7401), .ZN(n7399) );
  OAI21_X1 U7871 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n8128), .A(n7399), .ZN(
        n7630) );
  NAND2_X1 U7872 ( .A1(n7629), .A2(n7630), .ZN(n7628) );
  OAI21_X1 U7873 ( .B1(n8235), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7628), .ZN(
        n7617) );
  NOR2_X1 U7874 ( .A1(n8243), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6772) );
  AOI21_X1 U7875 ( .B1(n8243), .B2(P1_REG1_REG_14__SCAN_IN), .A(n6772), .ZN(
        n7618) );
  NAND2_X1 U7876 ( .A1(n7617), .A2(n7618), .ZN(n7616) );
  OAI21_X1 U7877 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n8243), .A(n7616), .ZN(
        n6773) );
  NOR2_X1 U7878 ( .A1(n8373), .A2(n6773), .ZN(n6774) );
  INV_X1 U7879 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10965) );
  XNOR2_X1 U7880 ( .A(n6773), .B(n8373), .ZN(n8065) );
  NOR2_X1 U7881 ( .A1(n10965), .A2(n8065), .ZN(n8064) );
  NOR2_X1 U7882 ( .A1(n6774), .A2(n8064), .ZN(n8181) );
  NAND2_X1 U7883 ( .A1(n8183), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6775) );
  OAI21_X1 U7884 ( .B1(n8183), .B2(P1_REG1_REG_16__SCAN_IN), .A(n6775), .ZN(
        n6776) );
  INV_X1 U7885 ( .A(n6776), .ZN(n8180) );
  NOR2_X1 U7886 ( .A1(n8181), .A2(n8180), .ZN(n8179) );
  AOI21_X1 U7887 ( .B1(n8462), .B2(P1_REG1_REG_16__SCAN_IN), .A(n8179), .ZN(
        n6779) );
  XNOR2_X1 U7888 ( .A(n9868), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n6778) );
  NOR2_X1 U7889 ( .A1(n6777), .A2(P1_U3084), .ZN(n10659) );
  AND2_X1 U7890 ( .A1(n10659), .A2(n5050), .ZN(n10666) );
  INV_X1 U7891 ( .A(n10666), .ZN(n10684) );
  NOR2_X1 U7892 ( .A1(n6779), .A2(n6778), .ZN(n9860) );
  AOI211_X1 U7893 ( .C1(n6779), .C2(n6778), .A(n10684), .B(n9860), .ZN(n6784)
         );
  OR2_X1 U7894 ( .A1(P1_U3083), .A2(n6780), .ZN(n6906) );
  INV_X1 U7895 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n6781) );
  NOR2_X1 U7896 ( .A1(n6906), .A2(n6781), .ZN(n6783) );
  INV_X1 U7897 ( .A(n6753), .ZN(n7135) );
  OR2_X1 U7898 ( .A1(n7298), .A2(n7135), .ZN(n10677) );
  INV_X1 U7899 ( .A(n9868), .ZN(n7627) );
  NAND2_X1 U7900 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9746) );
  OAI21_X1 U7901 ( .B1(n10677), .B2(n7627), .A(n9746), .ZN(n6782) );
  OR4_X1 U7902 ( .A1(n6785), .A2(n6784), .A3(n6783), .A4(n6782), .ZN(P1_U3258)
         );
  AND2_X1 U7903 ( .A1(n5720), .A2(P2_U3152), .ZN(n7761) );
  INV_X2 U7904 ( .A(n7761), .ZN(n9698) );
  AND2_X1 U7905 ( .A1(n5680), .A2(P2_U3152), .ZN(n8353) );
  OAI222_X1 U7906 ( .A1(n9698), .A2(n6786), .B1(n5043), .B2(n7114), .C1(
        P2_U3152), .C2(n10709), .ZN(P2_U3357) );
  OAI222_X1 U7907 ( .A1(n9698), .A2(n6788), .B1(n5043), .B2(n7105), .C1(
        P2_U3152), .C2(n6787), .ZN(P2_U3356) );
  NAND2_X1 U7908 ( .A1(n5680), .A2(P1_U3084), .ZN(n10575) );
  INV_X1 U7909 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7112) );
  AND2_X1 U7910 ( .A1(n6789), .A2(P1_U3084), .ZN(n8350) );
  OAI222_X1 U7911 ( .A1(n10575), .A2(n7112), .B1(n5044), .B2(n7114), .C1(
        n10676), .C2(P1_U3084), .ZN(P1_U3352) );
  INV_X1 U7912 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7184) );
  OAI222_X1 U7913 ( .A1(n10575), .A2(n7184), .B1(n5044), .B2(n7186), .C1(n9850), .C2(P1_U3084), .ZN(P1_U3350) );
  OAI222_X1 U7914 ( .A1(n9698), .A2(n6790), .B1(n5043), .B2(n7186), .C1(
        P2_U3152), .C2(n7056), .ZN(P2_U3355) );
  INV_X1 U7915 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7106) );
  OAI222_X1 U7916 ( .A1(n7109), .A2(P1_U3084), .B1(n5044), .B2(n7105), .C1(
        n7106), .C2(n10575), .ZN(P1_U3351) );
  INV_X1 U7917 ( .A(n7001), .ZN(n7031) );
  OAI222_X1 U7918 ( .A1(n9698), .A2(n5761), .B1(n5043), .B2(n7243), .C1(
        P2_U3152), .C2(n7031), .ZN(P2_U3354) );
  INV_X1 U7919 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7244) );
  OAI222_X1 U7920 ( .A1(n7247), .A2(P1_U3084), .B1(n5044), .B2(n7243), .C1(
        n7244), .C2(n10575), .ZN(P1_U3349) );
  NAND2_X1 U7921 ( .A1(n8436), .A2(P1_B_REG_SCAN_IN), .ZN(n6791) );
  INV_X1 U7922 ( .A(n8400), .ZN(n6943) );
  MUX2_X1 U7923 ( .A(n6791), .B(P1_B_REG_SCAN_IN), .S(n6943), .Z(n6792) );
  NAND2_X1 U7924 ( .A1(n6792), .A2(n10574), .ZN(n6944) );
  INV_X1 U7925 ( .A(n8436), .ZN(n6793) );
  OAI22_X1 U7926 ( .A1(n6944), .A2(P1_D_REG_1__SCAN_IN), .B1(n10574), .B2(
        n6793), .ZN(n7071) );
  AND2_X1 U7927 ( .A1(n8351), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6794) );
  NAND2_X1 U7928 ( .A1(n7208), .A2(n6794), .ZN(n10580) );
  NAND2_X1 U7929 ( .A1(n10580), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6795) );
  OAI21_X1 U7930 ( .B1(n7071), .B2(n10580), .A(n6795), .ZN(P1_U3441) );
  INV_X1 U7931 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6796) );
  INV_X1 U7932 ( .A(n6999), .ZN(n7043) );
  OAI222_X1 U7933 ( .A1(n9698), .A2(n6796), .B1(n5043), .B2(n7340), .C1(
        P2_U3152), .C2(n7043), .ZN(P2_U3353) );
  INV_X1 U7934 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7341) );
  INV_X1 U7935 ( .A(n10575), .ZN(n10571) );
  INV_X1 U7936 ( .A(n10571), .ZN(n8399) );
  OAI222_X1 U7937 ( .A1(n7344), .A2(P1_U3084), .B1(n5044), .B2(n7340), .C1(
        n7341), .C2(n8399), .ZN(P1_U3348) );
  INV_X1 U7938 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6797) );
  INV_X1 U7939 ( .A(n6998), .ZN(n7067) );
  OAI222_X1 U7940 ( .A1(n9698), .A2(n6797), .B1(n5043), .B2(n7436), .C1(
        P2_U3152), .C2(n7067), .ZN(P2_U3352) );
  INV_X1 U7941 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7437) );
  OAI222_X1 U7942 ( .A1(n7440), .A2(P1_U3084), .B1(n5044), .B2(n7436), .C1(
        n7437), .C2(n10575), .ZN(P1_U3347) );
  INV_X1 U7943 ( .A(n7512), .ZN(n6799) );
  INV_X1 U7944 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6798) );
  OAI222_X1 U7945 ( .A1(n6863), .A2(P1_U3084), .B1(n5044), .B2(n6799), .C1(
        n6798), .C2(n8399), .ZN(P1_U3346) );
  INV_X1 U7946 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6800) );
  INV_X1 U7947 ( .A(n7085), .ZN(n7091) );
  OAI222_X1 U7948 ( .A1(n9698), .A2(n6800), .B1(n5043), .B2(n6799), .C1(
        P2_U3152), .C2(n7091), .ZN(P2_U3351) );
  NAND2_X1 U7949 ( .A1(n9267), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6801) );
  OAI21_X1 U7950 ( .B1(n9267), .B2(n9094), .A(n6801), .ZN(P2_U3582) );
  INV_X1 U7951 ( .A(n6802), .ZN(n6806) );
  INV_X1 U7952 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6804) );
  AND3_X1 U7953 ( .A1(n6804), .A2(n6803), .A3(n6809), .ZN(n6805) );
  NAND2_X1 U7954 ( .A1(n6806), .A2(n6805), .ZN(n6813) );
  XNOR2_X2 U7955 ( .A(n6808), .B(n6807), .ZN(n10568) );
  NAND2_X1 U7956 ( .A1(n7351), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6821) );
  NAND2_X1 U7957 ( .A1(n6823), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7867) );
  INV_X1 U7958 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7866) );
  INV_X1 U7959 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7922) );
  INV_X1 U7960 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6815) );
  INV_X1 U7961 ( .A(n6846), .ZN(n8141) );
  NAND2_X1 U7962 ( .A1(n7925), .A2(n6815), .ZN(n6816) );
  AND2_X1 U7963 ( .A1(n8141), .A2(n6816), .ZN(n8223) );
  NAND2_X1 U7964 ( .A1(n7099), .A2(n8223), .ZN(n6820) );
  NAND2_X1 U7965 ( .A1(n5051), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6819) );
  NAND2_X1 U7966 ( .A1(n5038), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6818) );
  NAND4_X1 U7967 ( .A1(n6821), .A2(n6820), .A3(n6819), .A4(n6818), .ZN(n8284)
         );
  NAND2_X1 U7968 ( .A1(n8284), .A2(P1_U4006), .ZN(n6822) );
  OAI21_X1 U7969 ( .B1(n5940), .B2(P1_U4006), .A(n6822), .ZN(P1_U3567) );
  NAND2_X1 U7970 ( .A1(n7351), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6829) );
  INV_X1 U7971 ( .A(n6823), .ZN(n7520) );
  INV_X1 U7972 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6824) );
  NAND2_X1 U7973 ( .A1(n7520), .A2(n6824), .ZN(n6825) );
  AND2_X1 U7974 ( .A1(n7867), .A2(n6825), .ZN(n7977) );
  NAND2_X1 U7975 ( .A1(n7099), .A2(n7977), .ZN(n6828) );
  NAND2_X1 U7976 ( .A1(n5051), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6827) );
  NAND2_X1 U7977 ( .A1(n5038), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6826) );
  NAND4_X1 U7978 ( .A1(n6829), .A2(n6828), .A3(n6827), .A4(n6826), .ZN(n8120)
         );
  NAND2_X1 U7979 ( .A1(n8120), .A2(P1_U4006), .ZN(n6830) );
  OAI21_X1 U7980 ( .B1(P1_U4006), .B2(n5871), .A(n6830), .ZN(P1_U3564) );
  INV_X1 U7981 ( .A(n7819), .ZN(n6832) );
  INV_X1 U7982 ( .A(n7221), .ZN(n7228) );
  OAI222_X1 U7983 ( .A1(n9698), .A2(n6831), .B1(n5043), .B2(n6832), .C1(
        P2_U3152), .C2(n7228), .ZN(P2_U3350) );
  INV_X1 U7984 ( .A(n7820), .ZN(n6881) );
  OAI222_X1 U7985 ( .A1(n10575), .A2(n6833), .B1(n5044), .B2(n6832), .C1(n6881), .C2(P1_U3084), .ZN(P1_U3345) );
  OAI21_X1 U7986 ( .B1(n6836), .B2(n6835), .A(n6834), .ZN(n6845) );
  OAI211_X1 U7987 ( .C1(n6839), .C2(n6838), .A(n10666), .B(n6837), .ZN(n6840)
         );
  INV_X1 U7988 ( .A(n6840), .ZN(n6841) );
  AOI21_X1 U7989 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(n10679), .A(n6841), .ZN(
        n6844) );
  INV_X1 U7990 ( .A(n10677), .ZN(n10661) );
  INV_X1 U7991 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7353) );
  NOR2_X1 U7992 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7353), .ZN(n7483) );
  AOI21_X1 U7993 ( .B1(n10661), .B2(n6842), .A(n7483), .ZN(n6843) );
  OAI211_X1 U7994 ( .C1(n6845), .C2(n9890), .A(n6844), .B(n6843), .ZN(P1_U3247) );
  NAND2_X1 U7995 ( .A1(n6846), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8247) );
  INV_X1 U7996 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8246) );
  INV_X1 U7997 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8256) );
  NAND2_X1 U7998 ( .A1(n6847), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8472) );
  INV_X1 U7999 ( .A(n6847), .ZN(n8383) );
  INV_X1 U8000 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6848) );
  NAND2_X1 U8001 ( .A1(n8383), .A2(n6848), .ZN(n6849) );
  AND2_X1 U8002 ( .A1(n8472), .A2(n6849), .ZN(n9751) );
  NAND2_X1 U8003 ( .A1(n7099), .A2(n9751), .ZN(n6853) );
  NAND2_X1 U8004 ( .A1(n7351), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6852) );
  NAND2_X1 U8005 ( .A1(n5051), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6851) );
  NAND2_X1 U8006 ( .A1(n5039), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6850) );
  NAND4_X1 U8007 ( .A1(n6853), .A2(n6852), .A3(n6851), .A4(n6850), .ZN(n10978)
         );
  NAND2_X1 U8008 ( .A1(n10978), .A2(P1_U4006), .ZN(n6854) );
  OAI21_X1 U8009 ( .B1(n6054), .B2(P1_U4006), .A(n6854), .ZN(P1_U3572) );
  NAND2_X1 U8010 ( .A1(n10614), .A2(n6855), .ZN(n6856) );
  NAND2_X1 U8011 ( .A1(n6856), .A2(n7012), .ZN(n6858) );
  OR2_X1 U8012 ( .A1(n10614), .A2(n6633), .ZN(n6857) );
  NOR2_X1 U8013 ( .A1(n10718), .A2(P2_U3966), .ZN(P2_U3151) );
  AOI21_X1 U8014 ( .B1(n6861), .B2(n6860), .A(n6859), .ZN(n6871) );
  NAND2_X1 U8015 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3084), .ZN(n6862) );
  OAI21_X1 U8016 ( .B1(n10677), .B2(n6863), .A(n6862), .ZN(n6869) );
  AOI21_X1 U8017 ( .B1(n6866), .B2(n6865), .A(n6864), .ZN(n6867) );
  NOR2_X1 U8018 ( .A1(n10684), .A2(n6867), .ZN(n6868) );
  AOI211_X1 U8019 ( .C1(n10679), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n6869), .B(
        n6868), .ZN(n6870) );
  OAI21_X1 U8020 ( .B1(n6871), .B2(n9890), .A(n6870), .ZN(P1_U3248) );
  INV_X1 U8021 ( .A(n7377), .ZN(n7384) );
  INV_X1 U8022 ( .A(n7859), .ZN(n6873) );
  OAI222_X1 U8023 ( .A1(P2_U3152), .A2(n7384), .B1(n5043), .B2(n6873), .C1(
        n9698), .C2(n5871), .ZN(P2_U3349) );
  OAI222_X1 U8024 ( .A1(n6924), .A2(P1_U3084), .B1(n5044), .B2(n6873), .C1(
        n6872), .C2(n10575), .ZN(P1_U3344) );
  INV_X1 U8025 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6875) );
  NAND2_X1 U8026 ( .A1(P2_U3966), .A2(n9098), .ZN(n6874) );
  OAI21_X1 U8027 ( .B1(P2_U3966), .B2(n6875), .A(n6874), .ZN(P2_U3552) );
  INV_X1 U8028 ( .A(n6876), .ZN(n6877) );
  AOI21_X1 U8029 ( .B1(n6879), .B2(n6878), .A(n6877), .ZN(n6888) );
  NOR2_X1 U8030 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7517), .ZN(n7838) );
  INV_X1 U8031 ( .A(n7838), .ZN(n6880) );
  OAI21_X1 U8032 ( .B1(n10677), .B2(n6881), .A(n6880), .ZN(n6886) );
  NAND2_X1 U8033 ( .A1(n6883), .A2(n6882), .ZN(n6884) );
  AOI21_X1 U8034 ( .B1(n6920), .B2(n6884), .A(n10684), .ZN(n6885) );
  AOI211_X1 U8035 ( .C1(n10679), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n6886), .B(
        n6885), .ZN(n6887) );
  OAI21_X1 U8036 ( .B1(n6888), .B2(n9890), .A(n6887), .ZN(P1_U3249) );
  INV_X1 U8037 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9792) );
  INV_X1 U8038 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8614) );
  NOR2_X1 U8039 ( .A1(n8613), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6889) );
  OR2_X1 U8040 ( .A1(n8666), .A2(n6889), .ZN(n10025) );
  AOI22_X1 U8041 ( .A1(n5051), .A2(P1_REG0_REG_20__SCAN_IN), .B1(n5038), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n6891) );
  NAND2_X1 U8042 ( .A1(n7351), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6890) );
  OAI211_X1 U8043 ( .C1(n10025), .C2(n8618), .A(n6891), .B(n6890), .ZN(n10040)
         );
  NAND2_X1 U8044 ( .A1(n10040), .A2(P1_U4006), .ZN(n6892) );
  OAI21_X1 U8045 ( .B1(n6128), .B2(P1_U4006), .A(n6892), .ZN(P1_U3575) );
  INV_X1 U8046 ( .A(n8015), .ZN(n6912) );
  AOI22_X1 U8047 ( .A1(n9285), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n7761), .ZN(n6893) );
  OAI21_X1 U8048 ( .B1(n6912), .B2(n5043), .A(n6893), .ZN(P2_U3347) );
  INV_X1 U8049 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6905) );
  AND2_X1 U8050 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7361) );
  AOI21_X1 U8051 ( .B1(n6896), .B2(n6895), .A(n6894), .ZN(n6897) );
  NOR2_X1 U8052 ( .A1(n9890), .A2(n6897), .ZN(n6898) );
  AOI211_X1 U8053 ( .C1(n10661), .C2(n6899), .A(n7361), .B(n6898), .ZN(n6904)
         );
  OAI211_X1 U8054 ( .C1(n6902), .C2(n6901), .A(n10666), .B(n6900), .ZN(n6903)
         );
  OAI211_X1 U8055 ( .C1(n6906), .C2(n6905), .A(n6904), .B(n6903), .ZN(P1_U3246) );
  INV_X1 U8056 ( .A(n7919), .ZN(n6909) );
  INV_X1 U8057 ( .A(n7794), .ZN(n7785) );
  OAI222_X1 U8058 ( .A1(n9698), .A2(n6907), .B1(n5043), .B2(n6909), .C1(n7785), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  OAI222_X1 U8059 ( .A1(P1_U3084), .A2(n6910), .B1(n5044), .B2(n6909), .C1(
        n6908), .C2(n10575), .ZN(P1_U3343) );
  INV_X1 U8060 ( .A(n8016), .ZN(n7311) );
  INV_X1 U8061 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10287) );
  OAI222_X1 U8062 ( .A1(P1_U3084), .A2(n7311), .B1(n5044), .B2(n6912), .C1(
        n10287), .C2(n8399), .ZN(P1_U3342) );
  INV_X1 U8063 ( .A(n6913), .ZN(n6914) );
  AOI211_X1 U8064 ( .C1(n6916), .C2(n6915), .A(n9890), .B(n6914), .ZN(n6927)
         );
  INV_X1 U8065 ( .A(n6917), .ZN(n6919) );
  NAND3_X1 U8066 ( .A1(n6920), .A2(n6919), .A3(n6918), .ZN(n6921) );
  AOI21_X1 U8067 ( .B1(n6922), .B2(n6921), .A(n10684), .ZN(n6926) );
  NAND2_X1 U8068 ( .A1(n10679), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n6923) );
  NAND2_X1 U8069 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7971) );
  OAI211_X1 U8070 ( .C1(n10677), .C2(n6924), .A(n6923), .B(n7971), .ZN(n6925)
         );
  OR3_X1 U8071 ( .A1(n6927), .A2(n6926), .A3(n6925), .ZN(P1_U3250) );
  XNOR2_X1 U8072 ( .A(n6929), .B(n6928), .ZN(n8061) );
  AND2_X1 U8073 ( .A1(n8061), .A2(n9958), .ZN(n7207) );
  NOR2_X1 U8074 ( .A1(n7205), .A2(n7207), .ZN(n6932) );
  NOR2_X1 U8075 ( .A1(n10580), .A2(n6932), .ZN(n7412) );
  INV_X1 U8076 ( .A(n6944), .ZN(n10581) );
  NOR4_X1 U8077 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n6941) );
  NOR4_X1 U8078 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n6940) );
  INV_X1 U8079 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10583) );
  INV_X1 U8080 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10582) );
  INV_X1 U8081 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10611) );
  INV_X1 U8082 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10610) );
  NAND4_X1 U8083 ( .A1(n10583), .A2(n10582), .A3(n10611), .A4(n10610), .ZN(
        n6938) );
  NOR4_X1 U8084 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n6936) );
  NOR4_X1 U8085 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6935) );
  NOR4_X1 U8086 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n6934) );
  NOR4_X1 U8087 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6933) );
  NAND4_X1 U8088 ( .A1(n6936), .A2(n6935), .A3(n6934), .A4(n6933), .ZN(n6937)
         );
  NOR4_X1 U8089 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        n6938), .A4(n6937), .ZN(n6939) );
  NAND3_X1 U8090 ( .A1(n6941), .A2(n6940), .A3(n6939), .ZN(n6942) );
  NAND2_X1 U8091 ( .A1(n10581), .A2(n6942), .ZN(n7070) );
  INV_X1 U8092 ( .A(n8061), .ZN(n9037) );
  NAND4_X1 U8093 ( .A1(n7412), .A2(n7071), .A3(n7070), .A4(n7074), .ZN(n7174)
         );
  OAI22_X1 U8094 ( .A1(n6944), .A2(P1_D_REG_0__SCAN_IN), .B1(n10574), .B2(
        n6943), .ZN(n7411) );
  INV_X1 U8095 ( .A(n7411), .ZN(n10562) );
  INV_X2 U8096 ( .A(n10990), .ZN(n10993) );
  INV_X1 U8097 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6956) );
  NAND2_X1 U8098 ( .A1(n6789), .A2(SI_0_), .ZN(n6945) );
  XNOR2_X1 U8099 ( .A(n6945), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n10579) );
  MUX2_X1 U8100 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10579), .S(n7113), .Z(n7162)
         );
  INV_X1 U8101 ( .A(n7162), .ZN(n10732) );
  OR2_X1 U8102 ( .A1(n8985), .A2(n6957), .ZN(n7419) );
  INV_X1 U8103 ( .A(n7205), .ZN(n7506) );
  AND2_X1 U8104 ( .A1(n6753), .A2(n7506), .ZN(n10977) );
  NAND2_X1 U8105 ( .A1(n5051), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n7159) );
  INV_X1 U8106 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6946) );
  OR2_X1 U8107 ( .A1(n6948), .A2(n6946), .ZN(n7160) );
  NAND2_X1 U8108 ( .A1(n5039), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7158) );
  NAND2_X1 U8109 ( .A1(n7099), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n7161) );
  NAND2_X1 U8110 ( .A1(n5038), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6952) );
  NAND2_X1 U8111 ( .A1(n7099), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6951) );
  NAND4_X2 U8112 ( .A1(n6952), .A2(n6951), .A3(n6950), .A4(n6949), .ZN(n9831)
         );
  INV_X1 U8113 ( .A(n9831), .ZN(n6953) );
  NAND2_X1 U8114 ( .A1(n6953), .A2(n7162), .ZN(n7166) );
  NAND2_X1 U8115 ( .A1(n9831), .A2(n10732), .ZN(n8850) );
  AND2_X1 U8116 ( .A1(n7166), .A2(n8850), .ZN(n8994) );
  INV_X1 U8117 ( .A(n7419), .ZN(n7073) );
  NOR3_X1 U8118 ( .A1(n8994), .A2(n7506), .A3(n7073), .ZN(n6954) );
  AOI21_X1 U8119 ( .B1(n10977), .B2(n9829), .A(n6954), .ZN(n10735) );
  OAI21_X1 U8120 ( .B1(n10732), .B2(n7419), .A(n10735), .ZN(n10546) );
  NAND2_X1 U8121 ( .A1(n10546), .A2(n10993), .ZN(n6955) );
  OAI21_X1 U8122 ( .B1(n10993), .B2(n6956), .A(n6955), .ZN(P1_U3454) );
  INV_X1 U8123 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10656) );
  NAND2_X1 U8124 ( .A1(n7162), .A2(n5040), .ZN(n6959) );
  OR2_X1 U8125 ( .A1(n7208), .A2(n10656), .ZN(n6958) );
  AND2_X1 U8126 ( .A1(n6960), .A2(n5638), .ZN(n6963) );
  NAND2_X1 U8127 ( .A1(n7162), .A2(n8795), .ZN(n6961) );
  INV_X1 U8128 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10655) );
  NAND3_X1 U8129 ( .A1(n6962), .A2(n6961), .A3(n5632), .ZN(n7122) );
  MUX2_X1 U8130 ( .A(n10656), .B(n7081), .S(n5050), .Z(n6965) );
  OAI21_X1 U8131 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n5050), .A(n7135), .ZN(
        n10654) );
  NAND2_X1 U8132 ( .A1(n10654), .A2(n10656), .ZN(n6964) );
  OAI211_X1 U8133 ( .C1(n6965), .C2(n10654), .A(P1_U4006), .B(n6964), .ZN(
        n9844) );
  AOI21_X1 U8134 ( .B1(n6968), .B2(n6967), .A(n6966), .ZN(n6971) );
  AND2_X1 U8135 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7264) );
  AOI21_X1 U8136 ( .B1(n10661), .B2(n6969), .A(n7264), .ZN(n6970) );
  OAI21_X1 U8137 ( .B1(n6971), .B2(n9890), .A(n6970), .ZN(n6977) );
  AOI21_X1 U8138 ( .B1(n6974), .B2(n6973), .A(n6972), .ZN(n6975) );
  NOR2_X1 U8139 ( .A1(n10684), .A2(n6975), .ZN(n6976) );
  AOI211_X1 U8140 ( .C1(n10679), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n6977), .B(
        n6976), .ZN(n6978) );
  NAND2_X1 U8141 ( .A1(n9844), .A2(n6978), .ZN(P1_U3245) );
  INV_X1 U8142 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6979) );
  INV_X1 U8143 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6980) );
  MUX2_X1 U8144 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6980), .S(n10709), .Z(n10704) );
  NOR3_X1 U8145 ( .A1(n5709), .A2(n6979), .A3(n10704), .ZN(n10705) );
  NOR2_X1 U8146 ( .A1(n10709), .A2(n6980), .ZN(n6981) );
  NOR2_X1 U8147 ( .A1(n10705), .A2(n6981), .ZN(n10721) );
  NAND2_X1 U8148 ( .A1(n10723), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6982) );
  OAI21_X1 U8149 ( .B1(n10723), .B2(P2_REG2_REG_2__SCAN_IN), .A(n6982), .ZN(
        n10720) );
  NAND2_X1 U8150 ( .A1(n7003), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6983) );
  OAI21_X1 U8151 ( .B1(n7003), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6983), .ZN(
        n7047) );
  NOR2_X1 U8152 ( .A1(n7048), .A2(n7047), .ZN(n7046) );
  AOI21_X1 U8153 ( .B1(n7003), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7046), .ZN(
        n7023) );
  NAND2_X1 U8154 ( .A1(n7001), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6984) );
  OAI21_X1 U8155 ( .B1(n7001), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6984), .ZN(
        n7022) );
  NOR2_X1 U8156 ( .A1(n7023), .A2(n7022), .ZN(n7021) );
  AOI21_X1 U8157 ( .B1(n7001), .B2(P2_REG2_REG_4__SCAN_IN), .A(n7021), .ZN(
        n7036) );
  NAND2_X1 U8158 ( .A1(n6999), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6985) );
  OAI21_X1 U8159 ( .B1(n6999), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6985), .ZN(
        n7035) );
  NOR2_X1 U8160 ( .A1(n7036), .A2(n7035), .ZN(n7034) );
  AOI21_X1 U8161 ( .B1(n6999), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7034), .ZN(
        n7061) );
  INV_X1 U8162 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6986) );
  MUX2_X1 U8163 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6986), .S(n6998), .Z(n6987)
         );
  INV_X1 U8164 ( .A(n6987), .ZN(n7060) );
  NAND2_X1 U8165 ( .A1(n7085), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6988) );
  OAI21_X1 U8166 ( .B1(n7085), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6988), .ZN(
        n6994) );
  NAND2_X1 U8167 ( .A1(n10614), .A2(n7141), .ZN(n6991) );
  AND2_X1 U8168 ( .A1(n6989), .A2(n8354), .ZN(n6990) );
  NAND2_X1 U8169 ( .A1(n6991), .A2(n6990), .ZN(n7014) );
  NAND2_X1 U8170 ( .A1(n7014), .A2(n7012), .ZN(n6992) );
  NAND2_X1 U8171 ( .A1(n9267), .A2(n6992), .ZN(n6996) );
  NOR2_X1 U8172 ( .A1(n6366), .A2(n9091), .ZN(n6993) );
  NAND2_X1 U8173 ( .A1(n6996), .A2(n6993), .ZN(n10719) );
  AOI211_X1 U8174 ( .C1(n6995), .C2(n6994), .A(n7084), .B(n10719), .ZN(n7020)
         );
  NAND2_X1 U8175 ( .A1(n6996), .A2(n6366), .ZN(n10710) );
  NOR2_X1 U8176 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7589), .ZN(n6997) );
  AOI21_X1 U8177 ( .B1(n10718), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6997), .ZN(
        n7018) );
  INV_X1 U8178 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10827) );
  MUX2_X1 U8179 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10827), .S(n6998), .Z(n7063)
         );
  NAND2_X1 U8180 ( .A1(n6999), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7010) );
  INV_X1 U8181 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7000) );
  MUX2_X1 U8182 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n7000), .S(n6999), .Z(n7039)
         );
  NAND2_X1 U8183 ( .A1(n7001), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7009) );
  INV_X1 U8184 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7002) );
  MUX2_X1 U8185 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n7002), .S(n7001), .Z(n7027)
         );
  NAND2_X1 U8186 ( .A1(n7003), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7008) );
  INV_X1 U8187 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7004) );
  MUX2_X1 U8188 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n7004), .S(n7003), .Z(n7052)
         );
  NAND2_X1 U8189 ( .A1(n10723), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7007) );
  INV_X1 U8190 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7005) );
  MUX2_X1 U8191 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n7005), .S(n10723), .Z(n10727) );
  INV_X1 U8192 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7006) );
  MUX2_X1 U8193 ( .A(n7006), .B(P2_REG1_REG_1__SCAN_IN), .S(n10709), .Z(n10713) );
  NAND3_X1 U8194 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n10713), .ZN(n10712) );
  OAI21_X1 U8195 ( .B1(n10709), .B2(n7006), .A(n10712), .ZN(n10728) );
  NAND2_X1 U8196 ( .A1(n10727), .A2(n10728), .ZN(n10725) );
  NAND2_X1 U8197 ( .A1(n7007), .A2(n10725), .ZN(n7053) );
  NAND2_X1 U8198 ( .A1(n7052), .A2(n7053), .ZN(n7051) );
  NAND2_X1 U8199 ( .A1(n7008), .A2(n7051), .ZN(n7028) );
  NAND2_X1 U8200 ( .A1(n7027), .A2(n7028), .ZN(n7026) );
  NAND2_X1 U8201 ( .A1(n7009), .A2(n7026), .ZN(n7040) );
  NAND2_X1 U8202 ( .A1(n7039), .A2(n7040), .ZN(n7038) );
  NAND2_X1 U8203 ( .A1(n7010), .A2(n7038), .ZN(n7064) );
  NAND2_X1 U8204 ( .A1(n7063), .A2(n7064), .ZN(n7062) );
  OAI21_X1 U8205 ( .B1(n7067), .B2(n10827), .A(n7062), .ZN(n7016) );
  INV_X1 U8206 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7011) );
  MUX2_X1 U8207 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n7011), .S(n7085), .Z(n7015)
         );
  AND2_X1 U8208 ( .A1(n7012), .A2(n9091), .ZN(n7013) );
  NAND2_X1 U8209 ( .A1(n7015), .A2(n7016), .ZN(n7090) );
  OAI211_X1 U8210 ( .C1(n7016), .C2(n7015), .A(n10726), .B(n7090), .ZN(n7017)
         );
  OAI211_X1 U8211 ( .C1(n10710), .C2(n7091), .A(n7018), .B(n7017), .ZN(n7019)
         );
  OR2_X1 U8212 ( .A1(n7020), .A2(n7019), .ZN(P2_U3252) );
  AOI211_X1 U8213 ( .C1(n7023), .C2(n7022), .A(n7021), .B(n10719), .ZN(n7033)
         );
  INV_X1 U8214 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7024) );
  NOR2_X1 U8215 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7024), .ZN(n7025) );
  AOI21_X1 U8216 ( .B1(n10718), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n7025), .ZN(
        n7030) );
  OAI211_X1 U8217 ( .C1(n7028), .C2(n7027), .A(n10726), .B(n7026), .ZN(n7029)
         );
  OAI211_X1 U8218 ( .C1(n10710), .C2(n7031), .A(n7030), .B(n7029), .ZN(n7032)
         );
  OR2_X1 U8219 ( .A1(n7033), .A2(n7032), .ZN(P2_U3249) );
  AOI211_X1 U8220 ( .C1(n7036), .C2(n7035), .A(n7034), .B(n10719), .ZN(n7045)
         );
  NOR2_X1 U8221 ( .A1(n7037), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8774) );
  AOI21_X1 U8222 ( .B1(n10718), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8774), .ZN(
        n7042) );
  OAI211_X1 U8223 ( .C1(n7040), .C2(n7039), .A(n10726), .B(n7038), .ZN(n7041)
         );
  OAI211_X1 U8224 ( .C1(n10710), .C2(n7043), .A(n7042), .B(n7041), .ZN(n7044)
         );
  OR2_X1 U8225 ( .A1(n7045), .A2(n7044), .ZN(P2_U3250) );
  AOI211_X1 U8226 ( .C1(n7048), .C2(n7047), .A(n7046), .B(n10719), .ZN(n7058)
         );
  NOR2_X1 U8227 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7049), .ZN(n7050) );
  AOI21_X1 U8228 ( .B1(n10718), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n7050), .ZN(
        n7055) );
  OAI211_X1 U8229 ( .C1(n7053), .C2(n7052), .A(n10726), .B(n7051), .ZN(n7054)
         );
  OAI211_X1 U8230 ( .C1(n10710), .C2(n7056), .A(n7055), .B(n7054), .ZN(n7057)
         );
  OR2_X1 U8231 ( .A1(n7058), .A2(n7057), .ZN(P2_U3248) );
  AOI211_X1 U8232 ( .C1(n7061), .C2(n7060), .A(n7059), .B(n10719), .ZN(n7069)
         );
  NOR2_X1 U8233 ( .A1(n5810), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7577) );
  AOI21_X1 U8234 ( .B1(n10718), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n7577), .ZN(
        n7066) );
  OAI211_X1 U8235 ( .C1(n7064), .C2(n7063), .A(n10726), .B(n7062), .ZN(n7065)
         );
  OAI211_X1 U8236 ( .C1(n10710), .C2(n7067), .A(n7066), .B(n7065), .ZN(n7068)
         );
  OR2_X1 U8237 ( .A1(n7069), .A2(n7068), .ZN(P2_U3251) );
  INV_X1 U8238 ( .A(n7070), .ZN(n7072) );
  NOR2_X1 U8239 ( .A1(n7072), .A2(n7071), .ZN(n7414) );
  NAND2_X1 U8240 ( .A1(n7414), .A2(n10562), .ZN(n7136) );
  OR2_X1 U8241 ( .A1(n7136), .A2(n10580), .ZN(n7080) );
  NAND2_X1 U8242 ( .A1(n7073), .A2(n9037), .ZN(n7420) );
  OR2_X1 U8243 ( .A1(n7080), .A2(n7420), .ZN(n7075) );
  NAND2_X1 U8244 ( .A1(n7075), .A2(n10741), .ZN(n9811) );
  INV_X1 U8245 ( .A(n9811), .ZN(n9801) );
  NAND2_X1 U8246 ( .A1(n10977), .A2(n7207), .ZN(n7076) );
  INV_X1 U8247 ( .A(n9808), .ZN(n9798) );
  AND2_X1 U8248 ( .A1(n7420), .A2(n7205), .ZN(n7077) );
  NOR2_X1 U8249 ( .A1(n10580), .A2(n7077), .ZN(n7078) );
  NAND2_X1 U8250 ( .A1(n7136), .A2(n7078), .ZN(n7211) );
  NOR2_X2 U8251 ( .A1(n7419), .A2(n7207), .ZN(n10873) );
  NAND2_X1 U8252 ( .A1(n7136), .A2(n10984), .ZN(n7206) );
  NAND3_X1 U8253 ( .A1(n7211), .A2(n7206), .A3(n7412), .ZN(n8574) );
  AOI22_X1 U8254 ( .A1(n9798), .A2(n9829), .B1(n8574), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n7083) );
  OR2_X1 U8255 ( .A1(n10873), .A2(n7506), .ZN(n7079) );
  INV_X1 U8256 ( .A(n9813), .ZN(n9744) );
  NAND2_X1 U8257 ( .A1(n7081), .A2(n9744), .ZN(n7082) );
  OAI211_X1 U8258 ( .C1(n9801), .C2(n10732), .A(n7083), .B(n7082), .ZN(
        P1_U3230) );
  NAND2_X1 U8259 ( .A1(n7221), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7086) );
  OAI21_X1 U8260 ( .B1(n7221), .B2(P2_REG2_REG_8__SCAN_IN), .A(n7086), .ZN(
        n7087) );
  NOR2_X1 U8261 ( .A1(n7088), .A2(n7087), .ZN(n7220) );
  AOI211_X1 U8262 ( .C1(n7088), .C2(n7087), .A(n7220), .B(n10719), .ZN(n7098)
         );
  NOR2_X1 U8263 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7650), .ZN(n7089) );
  AOI21_X1 U8264 ( .B1(n10718), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7089), .ZN(
        n7096) );
  OAI21_X1 U8265 ( .B1(n7091), .B2(n7011), .A(n7090), .ZN(n7094) );
  INV_X1 U8266 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7092) );
  MUX2_X1 U8267 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7092), .S(n7221), .Z(n7093)
         );
  NAND2_X1 U8268 ( .A1(n7093), .A2(n7094), .ZN(n7227) );
  OAI211_X1 U8269 ( .C1(n7094), .C2(n7093), .A(n10726), .B(n7227), .ZN(n7095)
         );
  OAI211_X1 U8270 ( .C1(n10710), .C2(n7228), .A(n7096), .B(n7095), .ZN(n7097)
         );
  OR2_X1 U8271 ( .A1(n7098), .A2(n7097), .ZN(P2_U3253) );
  NAND2_X1 U8272 ( .A1(n7099), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n7103) );
  NAND2_X1 U8273 ( .A1(n5038), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7100) );
  NAND2_X1 U8274 ( .A1(n7113), .A2(n5720), .ZN(n7185) );
  OR2_X1 U8275 ( .A1(n7185), .A2(n7105), .ZN(n7108) );
  NAND2_X1 U8276 ( .A1(n7113), .A2(n5680), .ZN(n7183) );
  OR2_X1 U8277 ( .A1(n7183), .A2(n7106), .ZN(n7107) );
  NAND2_X1 U8278 ( .A1(n7272), .A2(n8795), .ZN(n7110) );
  OAI211_X1 U8279 ( .C1(n8985), .C2(n7111), .A(n9958), .B(n7205), .ZN(n7169)
         );
  AOI22_X1 U8280 ( .A1(n9828), .A2(n8790), .B1(n5040), .B2(n7272), .ZN(n7195)
         );
  XNOR2_X1 U8281 ( .A(n7194), .B(n7195), .ZN(n7192) );
  NAND2_X1 U8282 ( .A1(n9829), .A2(n5040), .ZN(n7118) );
  OR2_X1 U8283 ( .A1(n7183), .A2(n7112), .ZN(n7116) );
  NAND3_X2 U8284 ( .A1(n7116), .A2(n5631), .A3(n7115), .ZN(n8582) );
  NAND2_X1 U8285 ( .A1(n8582), .A2(n8795), .ZN(n7117) );
  NAND2_X1 U8286 ( .A1(n9829), .A2(n8790), .ZN(n7121) );
  NAND2_X1 U8287 ( .A1(n8582), .A2(n5040), .ZN(n7120) );
  NAND2_X1 U8288 ( .A1(n7121), .A2(n7120), .ZN(n7127) );
  NAND2_X1 U8289 ( .A1(n7126), .A2(n7127), .ZN(n7125) );
  INV_X1 U8290 ( .A(n7122), .ZN(n7123) );
  NAND2_X1 U8291 ( .A1(n7123), .A2(n8793), .ZN(n7124) );
  NAND2_X1 U8292 ( .A1(n7125), .A2(n8570), .ZN(n7129) );
  INV_X1 U8293 ( .A(n7127), .ZN(n8571) );
  NAND2_X1 U8294 ( .A1(n8573), .A2(n8571), .ZN(n7128) );
  NAND2_X1 U8295 ( .A1(n7129), .A2(n7128), .ZN(n7193) );
  XOR2_X1 U8296 ( .A(n7192), .B(n7130), .Z(n7139) );
  NAND2_X1 U8297 ( .A1(n7351), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7134) );
  INV_X1 U8298 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7200) );
  NAND2_X1 U8299 ( .A1(n7099), .A2(n7200), .ZN(n7133) );
  NAND2_X1 U8300 ( .A1(n5051), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n7132) );
  NAND2_X1 U8301 ( .A1(n7412), .A2(n10975), .ZN(n9043) );
  OR2_X1 U8302 ( .A1(n7136), .A2(n9043), .ZN(n9794) );
  AOI22_X1 U8303 ( .A1(n9798), .A2(n9827), .B1(n9805), .B2(n9829), .ZN(n7138)
         );
  AOI22_X1 U8304 ( .A1(n9811), .A2(n7272), .B1(n8574), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7137) );
  OAI211_X1 U8305 ( .C1(n7139), .C2(n9813), .A(n7138), .B(n7137), .ZN(P1_U3235) );
  INV_X1 U8306 ( .A(n8128), .ZN(n7403) );
  INV_X1 U8307 ( .A(n8127), .ZN(n7140) );
  OAI222_X1 U8308 ( .A1(n7403), .A2(P1_U3084), .B1(n5044), .B2(n7140), .C1(
        n10279), .C2(n8399), .ZN(P1_U3341) );
  INV_X1 U8309 ( .A(n7907), .ZN(n7903) );
  OAI222_X1 U8310 ( .A1(P2_U3152), .A2(n7903), .B1(n5043), .B2(n7140), .C1(
        n9698), .C2(n5940), .ZN(P2_U3346) );
  NOR2_X1 U8311 ( .A1(n7141), .A2(n6369), .ZN(n7142) );
  OR2_X1 U8312 ( .A1(n7143), .A2(n7142), .ZN(n9544) );
  INV_X1 U8313 ( .A(n10904), .ZN(n10936) );
  OAI21_X1 U8314 ( .B1(n7144), .B2(n9180), .A(n7676), .ZN(n7666) );
  NAND2_X1 U8315 ( .A1(n6433), .A2(n10742), .ZN(n7145) );
  NAND2_X1 U8316 ( .A1(n7711), .A2(n7145), .ZN(n7660) );
  AND2_X1 U8317 ( .A1(n5698), .A2(n8063), .ZN(n10940) );
  INV_X1 U8318 ( .A(n10940), .ZN(n10921) );
  INV_X1 U8319 ( .A(n10939), .ZN(n10919) );
  OAI22_X1 U8320 ( .A1(n7660), .A2(n10921), .B1(n10919), .B2(n7674), .ZN(n7151) );
  XOR2_X1 U8321 ( .A(n6438), .B(n7144), .Z(n7150) );
  NAND2_X1 U8322 ( .A1(n7147), .A2(n7146), .ZN(n10794) );
  INV_X1 U8323 ( .A(n10794), .ZN(n9538) );
  OAI22_X1 U8324 ( .A1(n7148), .A2(n9561), .B1(n7677), .B2(n9559), .ZN(n9184)
         );
  INV_X1 U8325 ( .A(n9184), .ZN(n7149) );
  OAI21_X1 U8326 ( .B1(n7150), .B2(n9538), .A(n7149), .ZN(n7663) );
  AOI211_X1 U8327 ( .C1(n10936), .C2(n7666), .A(n7151), .B(n7663), .ZN(n7292)
         );
  OR2_X1 U8328 ( .A1(n7657), .A2(n7152), .ZN(n7291) );
  AND2_X1 U8329 ( .A1(n10614), .A2(n7153), .ZN(n7154) );
  NAND2_X1 U8330 ( .A1(n7290), .A2(n7288), .ZN(n7156) );
  NAND2_X1 U8331 ( .A1(n10945), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7157) );
  OAI21_X1 U8332 ( .B1(n7292), .B2(n10945), .A(n7157), .ZN(P2_U3521) );
  INV_X1 U8333 ( .A(n10875), .ZN(n10933) );
  NAND2_X1 U8334 ( .A1(n7280), .A2(n8582), .ZN(n7278) );
  NAND2_X1 U8335 ( .A1(n9831), .A2(n7162), .ZN(n7164) );
  OAI21_X1 U8336 ( .B1(n7163), .B2(n7164), .A(n7271), .ZN(n8583) );
  NOR2_X2 U8337 ( .A1(n7419), .A2(n9037), .ZN(n10981) );
  NAND2_X1 U8338 ( .A1(n7269), .A2(n10732), .ZN(n7275) );
  OAI211_X1 U8339 ( .C1(n7269), .C2(n10732), .A(n10981), .B(n7275), .ZN(n8578)
         );
  OAI21_X1 U8340 ( .B1(n7269), .B2(n10984), .A(n8578), .ZN(n7173) );
  INV_X1 U8341 ( .A(n7279), .ZN(n7165) );
  AOI21_X1 U8342 ( .B1(n7163), .B2(n7166), .A(n7165), .ZN(n7172) );
  NAND2_X1 U8343 ( .A1(n8985), .A2(n10021), .ZN(n7168) );
  NAND2_X1 U8344 ( .A1(n6957), .A2(n9037), .ZN(n7167) );
  NAND2_X1 U8345 ( .A1(n7168), .A2(n7167), .ZN(n10980) );
  INV_X1 U8346 ( .A(n10980), .ZN(n9131) );
  AOI22_X1 U8347 ( .A1(n10975), .A2(n9831), .B1(n9828), .B2(n10977), .ZN(n7171) );
  INV_X1 U8348 ( .A(n7169), .ZN(n10879) );
  NAND2_X1 U8349 ( .A1(n8583), .A2(n10879), .ZN(n7170) );
  OAI211_X1 U8350 ( .C1(n7172), .C2(n9131), .A(n7171), .B(n7170), .ZN(n8580)
         );
  AOI211_X1 U8351 ( .C1(n10933), .C2(n8583), .A(n7173), .B(n8580), .ZN(n7217)
         );
  NAND2_X1 U8352 ( .A1(n10987), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7175) );
  OAI21_X1 U8353 ( .B1(n7217), .B2(n10987), .A(n7175), .ZN(P1_U3524) );
  NAND2_X1 U8354 ( .A1(n5052), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n7181) );
  INV_X1 U8355 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n7177) );
  NAND2_X1 U8356 ( .A1(n8666), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8667) );
  INV_X1 U8357 ( .A(n8667), .ZN(n7176) );
  NAND2_X1 U8358 ( .A1(n7176), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8603) );
  AOI21_X1 U8359 ( .B1(n7177), .B2(n8667), .A(n7367), .ZN(n9981) );
  NAND2_X1 U8360 ( .A1(n7099), .A2(n9981), .ZN(n7180) );
  NAND2_X1 U8361 ( .A1(n5051), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n7179) );
  NAND2_X1 U8362 ( .A1(n5039), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n7178) );
  NAND4_X1 U8363 ( .A1(n7181), .A2(n7180), .A3(n7179), .A4(n7178), .ZN(n9997)
         );
  NAND2_X1 U8364 ( .A1(n9997), .A2(P1_U4006), .ZN(n7182) );
  OAI21_X1 U8365 ( .B1(n6171), .B2(P1_U4006), .A(n7182), .ZN(P1_U3577) );
  NAND2_X1 U8366 ( .A1(n9827), .A2(n5040), .ZN(n7190) );
  OR2_X1 U8367 ( .A1(n7185), .A2(n7186), .ZN(n7187) );
  NAND2_X1 U8368 ( .A1(n7199), .A2(n8795), .ZN(n7189) );
  NAND2_X1 U8369 ( .A1(n7190), .A2(n7189), .ZN(n7191) );
  AOI22_X1 U8370 ( .A1(n9827), .A2(n8790), .B1(n5040), .B2(n7199), .ZN(n7239)
         );
  NAND2_X1 U8371 ( .A1(n7193), .A2(n7192), .ZN(n7198) );
  INV_X1 U8372 ( .A(n7194), .ZN(n7196) );
  NAND2_X1 U8373 ( .A1(n7196), .A2(n7195), .ZN(n7197) );
  NAND2_X1 U8374 ( .A1(n7198), .A2(n7197), .ZN(n7237) );
  XOR2_X1 U8375 ( .A(n7236), .B(n7237), .Z(n7216) );
  NAND2_X1 U8376 ( .A1(n7351), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7204) );
  XNOR2_X1 U8377 ( .A(n7200), .B(P1_REG3_REG_4__SCAN_IN), .ZN(n7499) );
  NAND2_X1 U8378 ( .A1(n7099), .A2(n7499), .ZN(n7203) );
  NAND2_X1 U8379 ( .A1(n5051), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n7202) );
  NAND2_X1 U8380 ( .A1(n5038), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7201) );
  NAND4_X1 U8381 ( .A1(n7204), .A2(n7203), .A3(n7202), .A4(n7201), .ZN(n9826)
         );
  INV_X1 U8382 ( .A(n9826), .ZN(n7444) );
  OAI22_X1 U8383 ( .A1(n9808), .A2(n7444), .B1(n7313), .B2(n9794), .ZN(n7214)
         );
  MUX2_X1 U8384 ( .A(n7207), .B(n7206), .S(n7205), .Z(n7209) );
  NAND3_X1 U8385 ( .A1(n7209), .A2(n7208), .A3(n8351), .ZN(n7210) );
  NAND2_X1 U8386 ( .A1(n7210), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7212) );
  NAND2_X1 U8387 ( .A1(n7212), .A2(n7211), .ZN(n9804) );
  MUX2_X1 U8388 ( .A(n9804), .B(P1_U3084), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n7213) );
  AOI211_X1 U8389 ( .C1(n7199), .C2(n9811), .A(n7214), .B(n7213), .ZN(n7215)
         );
  OAI21_X1 U8390 ( .B1(n7216), .B2(n9813), .A(n7215), .ZN(P1_U3216) );
  INV_X1 U8391 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7219) );
  OR2_X1 U8392 ( .A1(n7217), .A2(n10990), .ZN(n7218) );
  OAI21_X1 U8393 ( .B1(n10993), .B2(n7219), .A(n7218), .ZN(P1_U3457) );
  AOI21_X1 U8394 ( .B1(n7221), .B2(P2_REG2_REG_8__SCAN_IN), .A(n7220), .ZN(
        n7225) );
  INV_X1 U8395 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7222) );
  MUX2_X1 U8396 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7222), .S(n7377), .Z(n7223)
         );
  INV_X1 U8397 ( .A(n7223), .ZN(n7224) );
  NOR2_X1 U8398 ( .A1(n7225), .A2(n7224), .ZN(n7376) );
  AOI211_X1 U8399 ( .C1(n7225), .C2(n7224), .A(n7376), .B(n10719), .ZN(n7235)
         );
  NOR2_X1 U8400 ( .A1(n7226), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7597) );
  AOI21_X1 U8401 ( .B1(n10718), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7597), .ZN(
        n7233) );
  OAI21_X1 U8402 ( .B1(n7228), .B2(n7092), .A(n7227), .ZN(n7231) );
  INV_X1 U8403 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7229) );
  MUX2_X1 U8404 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n7229), .S(n7377), .Z(n7230)
         );
  NAND2_X1 U8405 ( .A1(n7230), .A2(n7231), .ZN(n7383) );
  OAI211_X1 U8406 ( .C1(n7231), .C2(n7230), .A(n10726), .B(n7383), .ZN(n7232)
         );
  OAI211_X1 U8407 ( .C1(n10710), .C2(n7384), .A(n7233), .B(n7232), .ZN(n7234)
         );
  OR2_X1 U8408 ( .A1(n7235), .A2(n7234), .ZN(P2_U3254) );
  NAND2_X1 U8409 ( .A1(n7237), .A2(n7236), .ZN(n7242) );
  INV_X1 U8410 ( .A(n7238), .ZN(n7240) );
  NAND2_X1 U8411 ( .A1(n7240), .A2(n7239), .ZN(n7241) );
  NAND2_X1 U8412 ( .A1(n9826), .A2(n5040), .ZN(n7249) );
  OR2_X1 U8413 ( .A1(n7185), .A2(n7243), .ZN(n7246) );
  OR2_X1 U8414 ( .A1(n7509), .A2(n7244), .ZN(n7245) );
  OAI211_X1 U8415 ( .C1(n7510), .C2(n7247), .A(n7246), .B(n7245), .ZN(n7500)
         );
  NAND2_X1 U8416 ( .A1(n7500), .A2(n8795), .ZN(n7248) );
  NAND2_X1 U8417 ( .A1(n7249), .A2(n7248), .ZN(n7251) );
  XNOR2_X1 U8418 ( .A(n7251), .B(n8724), .ZN(n7334) );
  NAND2_X1 U8419 ( .A1(n9826), .A2(n8790), .ZN(n7253) );
  NAND2_X1 U8420 ( .A1(n7500), .A2(n5040), .ZN(n7252) );
  AND2_X1 U8421 ( .A1(n7253), .A2(n7252), .ZN(n7335) );
  XNOR2_X1 U8422 ( .A(n7334), .B(n7335), .ZN(n7254) );
  XNOR2_X1 U8423 ( .A(n7339), .B(n7254), .ZN(n7268) );
  INV_X1 U8424 ( .A(n7500), .ZN(n10767) );
  NAND2_X1 U8425 ( .A1(n7351), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7262) );
  INV_X1 U8426 ( .A(n7255), .ZN(n7354) );
  INV_X1 U8427 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7257) );
  NAND2_X1 U8428 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7256) );
  NAND2_X1 U8429 ( .A1(n7257), .A2(n7256), .ZN(n7258) );
  AND2_X1 U8430 ( .A1(n7354), .A2(n7258), .ZN(n7549) );
  NAND2_X1 U8431 ( .A1(n7099), .A2(n7549), .ZN(n7261) );
  NAND2_X1 U8432 ( .A1(n5051), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n7260) );
  NAND2_X1 U8433 ( .A1(n5039), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7259) );
  NAND4_X1 U8434 ( .A1(n7262), .A2(n7261), .A3(n7260), .A4(n7259), .ZN(n9825)
         );
  INV_X1 U8435 ( .A(n9827), .ZN(n7493) );
  NOR2_X1 U8436 ( .A1(n9794), .A2(n7493), .ZN(n7263) );
  AOI211_X1 U8437 ( .C1(n9798), .C2(n9825), .A(n7264), .B(n7263), .ZN(n7265)
         );
  OAI21_X1 U8438 ( .B1(n10767), .B2(n9801), .A(n7265), .ZN(n7266) );
  AOI21_X1 U8439 ( .B1(n7499), .B2(n9804), .A(n7266), .ZN(n7267) );
  OAI21_X1 U8440 ( .B1(n7268), .B2(n9813), .A(n7267), .ZN(P1_U3228) );
  NAND2_X1 U8441 ( .A1(n7280), .A2(n7269), .ZN(n7270) );
  NAND2_X1 U8442 ( .A1(n7271), .A2(n7270), .ZN(n7273) );
  NAND2_X1 U8443 ( .A1(n9828), .A2(n7274), .ZN(n8854) );
  NAND2_X1 U8444 ( .A1(n8852), .A2(n8854), .ZN(n7277) );
  NAND2_X1 U8445 ( .A1(n7273), .A2(n7277), .ZN(n7315) );
  OAI21_X1 U8446 ( .B1(n7273), .B2(n7277), .A(n7315), .ZN(n7285) );
  INV_X1 U8447 ( .A(n7275), .ZN(n7276) );
  OAI21_X1 U8448 ( .B1(n7276), .B2(n7274), .A(n7326), .ZN(n7427) );
  INV_X1 U8449 ( .A(n10981), .ZN(n10960) );
  OAI22_X1 U8450 ( .A1(n7427), .A2(n10960), .B1(n7274), .B2(n10984), .ZN(n7284) );
  INV_X1 U8451 ( .A(n7285), .ZN(n7433) );
  INV_X1 U8452 ( .A(n7277), .ZN(n8995) );
  NAND2_X1 U8453 ( .A1(n8856), .A2(n8995), .ZN(n7318) );
  OAI21_X1 U8454 ( .B1(n8995), .B2(n8856), .A(n7318), .ZN(n7282) );
  INV_X1 U8455 ( .A(n10975), .ZN(n10013) );
  INV_X1 U8456 ( .A(n10977), .ZN(n10015) );
  OAI22_X1 U8457 ( .A1(n7280), .A2(n10013), .B1(n7493), .B2(n10015), .ZN(n7281) );
  AOI21_X1 U8458 ( .B1(n7282), .B2(n10980), .A(n7281), .ZN(n7283) );
  OAI21_X1 U8459 ( .B1(n7433), .B2(n7169), .A(n7283), .ZN(n7426) );
  AOI211_X1 U8460 ( .C1(n10933), .C2(n7285), .A(n7284), .B(n7426), .ZN(n10749)
         );
  NAND2_X1 U8461 ( .A1(n10987), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7286) );
  OAI21_X1 U8462 ( .B1(n10749), .B2(n10987), .A(n7286), .ZN(P1_U3525) );
  INV_X1 U8463 ( .A(n8242), .ZN(n7332) );
  AOI22_X1 U8464 ( .A1(n8243), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n10571), .ZN(n7287) );
  OAI21_X1 U8465 ( .B1(n7332), .B2(n5044), .A(n7287), .ZN(P1_U3339) );
  INV_X1 U8466 ( .A(n7288), .ZN(n7289) );
  NAND2_X1 U8467 ( .A1(n7290), .A2(n7289), .ZN(n7656) );
  INV_X2 U8468 ( .A(n10947), .ZN(n10950) );
  INV_X1 U8469 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7294) );
  OR2_X1 U8470 ( .A1(n7292), .A2(n10947), .ZN(n7293) );
  OAI21_X1 U8471 ( .B1(n10950), .B2(n7294), .A(n7293), .ZN(P2_U3454) );
  INV_X1 U8472 ( .A(n8234), .ZN(n7297) );
  INV_X1 U8473 ( .A(n8051), .ZN(n8046) );
  OAI222_X1 U8474 ( .A1(n9698), .A2(n7295), .B1(n5043), .B2(n7297), .C1(n8046), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8475 ( .A(n8235), .ZN(n7632) );
  OAI222_X1 U8476 ( .A1(P1_U3084), .A2(n7632), .B1(n5044), .B2(n7297), .C1(
        n7296), .C2(n8399), .ZN(P1_U3340) );
  INV_X1 U8477 ( .A(n7298), .ZN(n7301) );
  NAND2_X1 U8478 ( .A1(n10666), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7299) );
  OAI21_X1 U8479 ( .B1(n7303), .B2(n7299), .A(n10677), .ZN(n7300) );
  AOI21_X1 U8480 ( .B1(n7302), .B2(n7301), .A(n7300), .ZN(n7312) );
  AND2_X1 U8481 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8166) );
  NAND3_X1 U8482 ( .A1(n7303), .A2(n10897), .A3(n7311), .ZN(n7304) );
  AND3_X1 U8483 ( .A1(n7400), .A2(n10666), .A3(n7304), .ZN(n7305) );
  AOI211_X1 U8484 ( .C1(n10679), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n8166), .B(
        n7305), .ZN(n7310) );
  INV_X1 U8485 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7306) );
  NAND2_X1 U8486 ( .A1(n7311), .A2(n7306), .ZN(n7307) );
  INV_X1 U8487 ( .A(n9890), .ZN(n10681) );
  OAI211_X1 U8488 ( .C1(n7308), .C2(n7307), .A(n7406), .B(n10681), .ZN(n7309)
         );
  OAI211_X1 U8489 ( .C1(n7312), .C2(n7311), .A(n7310), .B(n7309), .ZN(P1_U3252) );
  INV_X2 U8490 ( .A(n10987), .ZN(n10989) );
  NAND2_X1 U8491 ( .A1(n7313), .A2(n7274), .ZN(n7314) );
  NAND2_X1 U8492 ( .A1(n7315), .A2(n7314), .ZN(n7316) );
  NAND2_X1 U8493 ( .A1(n9827), .A2(n7441), .ZN(n8859) );
  NAND2_X1 U8494 ( .A1(n7316), .A2(n8992), .ZN(n7443) );
  OR2_X1 U8495 ( .A1(n7316), .A2(n8992), .ZN(n7317) );
  NAND2_X1 U8496 ( .A1(n7443), .A2(n7317), .ZN(n7322) );
  INV_X1 U8497 ( .A(n7322), .ZN(n7425) );
  INV_X1 U8498 ( .A(n8992), .ZN(n7320) );
  NAND2_X1 U8499 ( .A1(n7318), .A2(n8852), .ZN(n7319) );
  NAND2_X1 U8500 ( .A1(n7319), .A2(n7320), .ZN(n7434) );
  OAI21_X1 U8501 ( .B1(n7320), .B2(n7319), .A(n7434), .ZN(n7321) );
  NAND2_X1 U8502 ( .A1(n7321), .A2(n10980), .ZN(n7325) );
  NAND2_X1 U8503 ( .A1(n7322), .A2(n10879), .ZN(n7324) );
  AOI22_X1 U8504 ( .A1(n10975), .A2(n9828), .B1(n9826), .B2(n10977), .ZN(n7323) );
  AND3_X1 U8505 ( .A1(n7325), .A2(n7324), .A3(n7323), .ZN(n7416) );
  AOI21_X1 U8506 ( .B1(n7199), .B2(n7326), .A(n7497), .ZN(n7422) );
  AOI22_X1 U8507 ( .A1(n7422), .A2(n10981), .B1(n10873), .B2(n7199), .ZN(n7327) );
  OAI211_X1 U8508 ( .C1(n7425), .C2(n10875), .A(n7416), .B(n7327), .ZN(n7329)
         );
  NAND2_X1 U8509 ( .A1(n7329), .A2(n10989), .ZN(n7328) );
  OAI21_X1 U8510 ( .B1(n10989), .B2(n6760), .A(n7328), .ZN(P1_U3526) );
  INV_X1 U8511 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7331) );
  NAND2_X1 U8512 ( .A1(n7329), .A2(n10993), .ZN(n7330) );
  OAI21_X1 U8513 ( .B1(n10993), .B2(n7331), .A(n7330), .ZN(P1_U3463) );
  INV_X1 U8514 ( .A(n8199), .ZN(n8207) );
  OAI222_X1 U8515 ( .A1(n9698), .A2(n7333), .B1(n5043), .B2(n7332), .C1(n8207), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8516 ( .A(n7334), .ZN(n7337) );
  INV_X1 U8517 ( .A(n7335), .ZN(n7336) );
  NAND2_X1 U8518 ( .A1(n7337), .A2(n7336), .ZN(n7338) );
  NAND2_X1 U8519 ( .A1(n9825), .A2(n8790), .ZN(n7346) );
  OR2_X1 U8520 ( .A1(n7185), .A2(n7340), .ZN(n7343) );
  OR2_X1 U8521 ( .A1(n7509), .A2(n7341), .ZN(n7342) );
  OAI211_X1 U8522 ( .C1(n7510), .C2(n7344), .A(n7343), .B(n7342), .ZN(n7558)
         );
  NAND2_X1 U8523 ( .A1(n7558), .A2(n5040), .ZN(n7345) );
  NAND2_X1 U8524 ( .A1(n7346), .A2(n7345), .ZN(n7466) );
  NAND2_X1 U8525 ( .A1(n9825), .A2(n5040), .ZN(n7348) );
  NAND2_X1 U8526 ( .A1(n7558), .A2(n8795), .ZN(n7347) );
  NAND2_X1 U8527 ( .A1(n7348), .A2(n7347), .ZN(n7349) );
  XNOR2_X1 U8528 ( .A(n7349), .B(n8793), .ZN(n7467) );
  XOR2_X1 U8529 ( .A(n7466), .B(n7467), .Z(n7350) );
  XNOR2_X1 U8530 ( .A(n7468), .B(n7350), .ZN(n7366) );
  INV_X1 U8531 ( .A(n7558), .ZN(n7363) );
  NAND2_X1 U8532 ( .A1(n7351), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7359) );
  INV_X1 U8533 ( .A(n7352), .ZN(n7451) );
  NAND2_X1 U8534 ( .A1(n7354), .A2(n7353), .ZN(n7355) );
  AND2_X1 U8535 ( .A1(n7451), .A2(n7355), .ZN(n7486) );
  NAND2_X1 U8536 ( .A1(n7099), .A2(n7486), .ZN(n7358) );
  NAND2_X1 U8537 ( .A1(n5051), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n7357) );
  NAND2_X1 U8538 ( .A1(n5039), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7356) );
  NAND4_X1 U8539 ( .A1(n7359), .A2(n7358), .A3(n7357), .A4(n7356), .ZN(n9824)
         );
  NOR2_X1 U8540 ( .A1(n9794), .A2(n7444), .ZN(n7360) );
  AOI211_X1 U8541 ( .C1(n9798), .C2(n9824), .A(n7361), .B(n7360), .ZN(n7362)
         );
  OAI21_X1 U8542 ( .B1(n7363), .B2(n9801), .A(n7362), .ZN(n7364) );
  AOI21_X1 U8543 ( .B1(n7549), .B2(n9804), .A(n7364), .ZN(n7365) );
  OAI21_X1 U8544 ( .B1(n7366), .B2(n9813), .A(n7365), .ZN(P1_U3225) );
  AOI22_X1 U8545 ( .A1(n5052), .A2(P1_REG1_REG_29__SCAN_IN), .B1(n5051), .B2(
        P1_REG0_REG_29__SCAN_IN), .ZN(n7374) );
  NAND2_X1 U8546 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(n7367), .ZN(n8692) );
  INV_X1 U8547 ( .A(n8692), .ZN(n7368) );
  NAND2_X1 U8548 ( .A1(n7368), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8694) );
  INV_X1 U8549 ( .A(n8694), .ZN(n7369) );
  NAND2_X1 U8550 ( .A1(n7369), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8710) );
  INV_X1 U8551 ( .A(n8710), .ZN(n7370) );
  NAND2_X1 U8552 ( .A1(n7370), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8732) );
  INV_X1 U8553 ( .A(n8732), .ZN(n7372) );
  AND2_X1 U8554 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n7371) );
  NAND2_X1 U8555 ( .A1(n7372), .A2(n7371), .ZN(n8734) );
  INV_X1 U8556 ( .A(n8734), .ZN(n9152) );
  AOI22_X1 U8557 ( .A1(n7099), .A2(n9152), .B1(n5039), .B2(
        P1_REG2_REG_29__SCAN_IN), .ZN(n7373) );
  INV_X1 U8558 ( .A(P1_U4006), .ZN(n9830) );
  NAND2_X1 U8559 ( .A1(n9830), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7375) );
  OAI21_X1 U8560 ( .B1(n9133), .B2(n9830), .A(n7375), .ZN(P1_U3584) );
  INV_X1 U8561 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7378) );
  MUX2_X1 U8562 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7378), .S(n7794), .Z(n7379)
         );
  INV_X1 U8563 ( .A(n7379), .ZN(n7380) );
  AOI211_X1 U8564 ( .C1(n7381), .C2(n7380), .A(n7793), .B(n10719), .ZN(n7391)
         );
  NOR2_X1 U8565 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10140), .ZN(n7382) );
  AOI21_X1 U8566 ( .B1(n10718), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7382), .ZN(
        n7389) );
  OAI21_X1 U8567 ( .B1(n7384), .B2(n7229), .A(n7383), .ZN(n7387) );
  INV_X1 U8568 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7385) );
  MUX2_X1 U8569 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7385), .S(n7794), .Z(n7386)
         );
  NAND2_X1 U8570 ( .A1(n7386), .A2(n7387), .ZN(n7784) );
  OAI211_X1 U8571 ( .C1(n7387), .C2(n7386), .A(n10726), .B(n7784), .ZN(n7388)
         );
  OAI211_X1 U8572 ( .C1(n10710), .C2(n7785), .A(n7389), .B(n7388), .ZN(n7390)
         );
  OR2_X1 U8573 ( .A1(n7391), .A2(n7390), .ZN(P2_U3255) );
  NAND2_X1 U8574 ( .A1(n5052), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n7395) );
  XNOR2_X1 U8575 ( .A(n8732), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9906) );
  NAND2_X1 U8576 ( .A1(n7099), .A2(n9906), .ZN(n7394) );
  NAND2_X1 U8577 ( .A1(n5051), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n7393) );
  NAND2_X1 U8578 ( .A1(n5039), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n7392) );
  NAND4_X1 U8579 ( .A1(n7395), .A2(n7394), .A3(n7393), .A4(n7392), .ZN(n9915)
         );
  NAND2_X1 U8580 ( .A1(n9915), .A2(P1_U4006), .ZN(n7396) );
  OAI21_X1 U8581 ( .B1(n6285), .B2(P1_U4006), .A(n7396), .ZN(P1_U3582) );
  INV_X1 U8582 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7397) );
  INV_X1 U8583 ( .A(n8372), .ZN(n7398) );
  INV_X1 U8584 ( .A(n9302), .ZN(n9295) );
  OAI222_X1 U8585 ( .A1(n9698), .A2(n7397), .B1(n5043), .B2(n7398), .C1(
        P2_U3152), .C2(n9295), .ZN(P2_U3343) );
  INV_X1 U8586 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10280) );
  OAI222_X1 U8587 ( .A1(n8373), .A2(P1_U3084), .B1(n5044), .B2(n7398), .C1(
        n10280), .C2(n8399), .ZN(P1_U3338) );
  OAI21_X1 U8588 ( .B1(n7401), .B2(n7400), .A(n7399), .ZN(n7409) );
  NAND2_X1 U8589 ( .A1(n10679), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n7402) );
  NAND2_X1 U8590 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8224) );
  OAI211_X1 U8591 ( .C1(n10677), .C2(n7403), .A(n7402), .B(n8224), .ZN(n7408)
         );
  AOI211_X1 U8592 ( .C1(n7406), .C2(n7405), .A(n9890), .B(n7404), .ZN(n7407)
         );
  AOI211_X1 U8593 ( .C1(n10666), .C2(n7409), .A(n7408), .B(n7407), .ZN(n7410)
         );
  INV_X1 U8594 ( .A(n7410), .ZN(P1_U3253) );
  AND2_X1 U8595 ( .A1(n7412), .A2(n7411), .ZN(n7413) );
  NAND2_X1 U8596 ( .A1(n7414), .A2(n7413), .ZN(n7533) );
  INV_X2 U8597 ( .A(n10022), .ZN(n10738) );
  OR3_X1 U8598 ( .A1(n10738), .A2(n7415), .A3(n9958), .ZN(n10029) );
  MUX2_X1 U8599 ( .A(n7417), .B(n7416), .S(n10022), .Z(n7424) );
  OR3_X1 U8600 ( .A1(n10738), .A2(n7419), .A3(n7418), .ZN(n10733) );
  OAI22_X1 U8601 ( .A1(n10734), .A2(n7441), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10741), .ZN(n7421) );
  AOI21_X1 U8602 ( .B1(n7422), .B2(n10068), .A(n7421), .ZN(n7423) );
  OAI211_X1 U8603 ( .C1(n7425), .C2(n10029), .A(n7424), .B(n7423), .ZN(
        P1_U3288) );
  NAND2_X1 U8604 ( .A1(n7426), .A2(n10022), .ZN(n7432) );
  NOR2_X1 U8605 ( .A1(n10733), .A2(n7427), .ZN(n7430) );
  INV_X1 U8606 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9832) );
  OAI22_X1 U8607 ( .A1(n10022), .A2(n7428), .B1(n9832), .B2(n10741), .ZN(n7429) );
  AOI211_X1 U8608 ( .C1(n10996), .C2(n7272), .A(n7430), .B(n7429), .ZN(n7431)
         );
  OAI211_X1 U8609 ( .C1(n7433), .C2(n10029), .A(n7432), .B(n7431), .ZN(
        P1_U3289) );
  NAND2_X1 U8610 ( .A1(n7434), .A2(n8857), .ZN(n7489) );
  NAND2_X1 U8611 ( .A1(n9826), .A2(n10767), .ZN(n8860) );
  NAND2_X1 U8612 ( .A1(n7444), .A2(n7500), .ZN(n7525) );
  NAND2_X1 U8613 ( .A1(n7527), .A2(n7525), .ZN(n7546) );
  INV_X1 U8614 ( .A(n9825), .ZN(n7492) );
  OR2_X1 U8615 ( .A1(n7492), .A2(n7558), .ZN(n7528) );
  NAND2_X1 U8616 ( .A1(n7546), .A2(n7528), .ZN(n7435) );
  NAND2_X1 U8617 ( .A1(n7492), .A2(n7558), .ZN(n7526) );
  NAND2_X1 U8618 ( .A1(n7435), .A2(n7526), .ZN(n8880) );
  INV_X1 U8619 ( .A(n9824), .ZN(n7530) );
  OR2_X1 U8620 ( .A1(n7185), .A2(n7436), .ZN(n7439) );
  OR2_X1 U8621 ( .A1(n7509), .A2(n7437), .ZN(n7438) );
  OAI211_X1 U8622 ( .C1(n7510), .C2(n7440), .A(n7439), .B(n7438), .ZN(n7472)
         );
  NAND2_X1 U8623 ( .A1(n7530), .A2(n7472), .ZN(n8882) );
  INV_X1 U8624 ( .A(n7472), .ZN(n10814) );
  NAND2_X1 U8625 ( .A1(n9824), .A2(n10814), .ZN(n8881) );
  AND2_X1 U8626 ( .A1(n8882), .A2(n8881), .ZN(n8886) );
  XNOR2_X1 U8627 ( .A(n8880), .B(n7448), .ZN(n7459) );
  NAND2_X1 U8628 ( .A1(n7493), .A2(n7441), .ZN(n7442) );
  NAND2_X1 U8629 ( .A1(n7443), .A2(n7442), .ZN(n7491) );
  NAND2_X1 U8630 ( .A1(n7525), .A2(n8860), .ZN(n8993) );
  NAND2_X1 U8631 ( .A1(n7444), .A2(n10767), .ZN(n7445) );
  NAND2_X1 U8632 ( .A1(n9825), .A2(n7558), .ZN(n7447) );
  OAI21_X1 U8633 ( .B1(n7449), .B2(n7448), .A(n7508), .ZN(n10818) );
  INV_X1 U8634 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7450) );
  NAND2_X1 U8635 ( .A1(n7451), .A2(n7450), .ZN(n7452) );
  AND2_X1 U8636 ( .A1(n7518), .A2(n7452), .ZN(n7534) );
  NAND2_X1 U8637 ( .A1(n7099), .A2(n7534), .ZN(n7456) );
  NAND2_X1 U8638 ( .A1(n7351), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7455) );
  NAND2_X1 U8639 ( .A1(n5051), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n7454) );
  NAND2_X1 U8640 ( .A1(n5038), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7453) );
  NAND4_X1 U8641 ( .A1(n7456), .A2(n7455), .A3(n7454), .A4(n7453), .ZN(n9823)
         );
  INV_X1 U8642 ( .A(n9823), .ZN(n7888) );
  OAI22_X1 U8643 ( .A1(n7492), .A2(n10013), .B1(n7888), .B2(n10015), .ZN(n7457) );
  AOI21_X1 U8644 ( .B1(n10818), .B2(n10879), .A(n7457), .ZN(n7458) );
  OAI21_X1 U8645 ( .B1(n9131), .B2(n7459), .A(n7458), .ZN(n10816) );
  INV_X1 U8646 ( .A(n10816), .ZN(n7465) );
  INV_X1 U8647 ( .A(n10029), .ZN(n9929) );
  NAND2_X1 U8648 ( .A1(n7497), .A2(n10767), .ZN(n7545) );
  AND2_X1 U8649 ( .A1(n7543), .A2(n7472), .ZN(n7460) );
  OR2_X1 U8650 ( .A1(n7460), .A2(n7531), .ZN(n10815) );
  INV_X1 U8651 ( .A(n10741), .ZN(n10994) );
  AOI22_X1 U8652 ( .A1(n10738), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7486), .B2(
        n10994), .ZN(n7462) );
  NAND2_X1 U8653 ( .A1(n10996), .A2(n7472), .ZN(n7461) );
  OAI211_X1 U8654 ( .C1(n10815), .C2(n10733), .A(n7462), .B(n7461), .ZN(n7463)
         );
  AOI21_X1 U8655 ( .B1(n10818), .B2(n9929), .A(n7463), .ZN(n7464) );
  OAI21_X1 U8656 ( .B1(n7465), .B2(n10738), .A(n7464), .ZN(P1_U3285) );
  NAND2_X1 U8657 ( .A1(n9824), .A2(n7104), .ZN(n7470) );
  NAND2_X1 U8658 ( .A1(n7472), .A2(n8795), .ZN(n7469) );
  NAND2_X1 U8659 ( .A1(n7470), .A2(n7469), .ZN(n7471) );
  XNOR2_X1 U8660 ( .A(n7471), .B(n8793), .ZN(n7475) );
  NAND2_X1 U8661 ( .A1(n9824), .A2(n8790), .ZN(n7474) );
  NAND2_X1 U8662 ( .A1(n7472), .A2(n5040), .ZN(n7473) );
  NAND2_X1 U8663 ( .A1(n7474), .A2(n7473), .ZN(n7476) );
  INV_X1 U8664 ( .A(n7691), .ZN(n7481) );
  INV_X1 U8665 ( .A(n7475), .ZN(n7478) );
  INV_X1 U8666 ( .A(n7476), .ZN(n7477) );
  NAND2_X1 U8667 ( .A1(n7478), .A2(n7477), .ZN(n7690) );
  NAND2_X1 U8668 ( .A1(n5080), .A2(n7690), .ZN(n7480) );
  AOI22_X1 U8669 ( .A1(n7481), .A2(n7690), .B1(n7479), .B2(n7480), .ZN(n7488)
         );
  NOR2_X1 U8670 ( .A1(n9794), .A2(n7492), .ZN(n7482) );
  AOI211_X1 U8671 ( .C1(n9798), .C2(n9823), .A(n7483), .B(n7482), .ZN(n7484)
         );
  OAI21_X1 U8672 ( .B1(n10814), .B2(n9801), .A(n7484), .ZN(n7485) );
  AOI21_X1 U8673 ( .B1(n7486), .B2(n9804), .A(n7485), .ZN(n7487) );
  OAI21_X1 U8674 ( .B1(n7488), .B2(n9813), .A(n7487), .ZN(P1_U3237) );
  XNOR2_X1 U8675 ( .A(n7489), .B(n8993), .ZN(n7496) );
  OAI21_X1 U8676 ( .B1(n7491), .B2(n8993), .A(n7490), .ZN(n10771) );
  OAI22_X1 U8677 ( .A1(n7493), .A2(n10013), .B1(n7492), .B2(n10015), .ZN(n7494) );
  AOI21_X1 U8678 ( .B1(n10771), .B2(n10879), .A(n7494), .ZN(n7495) );
  OAI21_X1 U8679 ( .B1(n9131), .B2(n7496), .A(n7495), .ZN(n10769) );
  INV_X1 U8680 ( .A(n10769), .ZN(n7505) );
  OR2_X1 U8681 ( .A1(n7497), .A2(n10767), .ZN(n7498) );
  NAND2_X1 U8682 ( .A1(n7545), .A2(n7498), .ZN(n10768) );
  AOI22_X1 U8683 ( .A1(n10738), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7499), .B2(
        n10994), .ZN(n7502) );
  NAND2_X1 U8684 ( .A1(n10996), .A2(n7500), .ZN(n7501) );
  OAI211_X1 U8685 ( .C1(n10768), .C2(n10733), .A(n7502), .B(n7501), .ZN(n7503)
         );
  AOI21_X1 U8686 ( .B1(n10771), .B2(n9929), .A(n7503), .ZN(n7504) );
  OAI21_X1 U8687 ( .B1(n7505), .B2(n10738), .A(n7504), .ZN(P1_U3287) );
  NAND2_X1 U8688 ( .A1(n7530), .A2(n10814), .ZN(n7507) );
  AOI22_X1 U8689 ( .A1(n8638), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8637), .B2(
        n7511), .ZN(n7514) );
  NAND2_X1 U8690 ( .A1(n7512), .A2(n8749), .ZN(n7513) );
  NAND2_X1 U8691 ( .A1(n7514), .A2(n7513), .ZN(n7702) );
  NAND2_X1 U8692 ( .A1(n7888), .A2(n7702), .ZN(n8889) );
  INV_X1 U8693 ( .A(n7702), .ZN(n7854) );
  NAND2_X1 U8694 ( .A1(n9823), .A2(n7854), .ZN(n8888) );
  NAND2_X1 U8695 ( .A1(n8889), .A2(n8888), .ZN(n8999) );
  OAI21_X1 U8696 ( .B1(n7515), .B2(n8999), .A(n7856), .ZN(n7516) );
  INV_X1 U8697 ( .A(n7516), .ZN(n7704) );
  NAND2_X1 U8698 ( .A1(n7351), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7524) );
  NAND2_X1 U8699 ( .A1(n7518), .A2(n7517), .ZN(n7519) );
  AND2_X1 U8700 ( .A1(n7520), .A2(n7519), .ZN(n7836) );
  NAND2_X1 U8701 ( .A1(n7099), .A2(n7836), .ZN(n7523) );
  NAND2_X1 U8702 ( .A1(n5051), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7522) );
  NAND2_X1 U8703 ( .A1(n5039), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7521) );
  NAND4_X1 U8704 ( .A1(n7524), .A2(n7523), .A3(n7522), .A4(n7521), .ZN(n9822)
         );
  INV_X1 U8705 ( .A(n9822), .ZN(n7873) );
  XOR2_X1 U8706 ( .A(n8999), .B(n7863), .Z(n7529) );
  OAI222_X1 U8707 ( .A1(n10015), .A2(n7873), .B1(n10013), .B2(n7530), .C1(
        n9131), .C2(n7529), .ZN(n7700) );
  NAND2_X1 U8708 ( .A1(n7700), .A2(n10022), .ZN(n7539) );
  INV_X1 U8709 ( .A(n7531), .ZN(n7532) );
  AOI211_X1 U8710 ( .C1(n7702), .C2(n7532), .A(n10960), .B(n7893), .ZN(n7701)
         );
  NOR2_X1 U8711 ( .A1(n7533), .A2(n10021), .ZN(n10999) );
  NOR2_X1 U8712 ( .A1(n10734), .A2(n7854), .ZN(n7537) );
  INV_X1 U8713 ( .A(n7534), .ZN(n7699) );
  OAI22_X1 U8714 ( .A1(n10022), .A2(n7535), .B1(n7699), .B2(n10741), .ZN(n7536) );
  AOI211_X1 U8715 ( .C1(n7701), .C2(n10999), .A(n7537), .B(n7536), .ZN(n7538)
         );
  OAI211_X1 U8716 ( .C1(n10070), .C2(n7704), .A(n7539), .B(n7538), .ZN(
        P1_U3284) );
  INV_X1 U8717 ( .A(n8461), .ZN(n7541) );
  OAI222_X1 U8718 ( .A1(n8183), .A2(P1_U3084), .B1(n5044), .B2(n7541), .C1(
        n7540), .C2(n8399), .ZN(P1_U3337) );
  INV_X1 U8719 ( .A(n9316), .ZN(n9323) );
  OAI222_X1 U8720 ( .A1(n9698), .A2(n7542), .B1(n5043), .B2(n7541), .C1(
        P2_U3152), .C2(n9323), .ZN(P2_U3342) );
  INV_X1 U8721 ( .A(n7543), .ZN(n7544) );
  AOI211_X1 U8722 ( .C1(n7558), .C2(n7545), .A(n10960), .B(n7544), .ZN(n7557)
         );
  XNOR2_X1 U8723 ( .A(n7546), .B(n8996), .ZN(n7547) );
  AOI222_X1 U8724 ( .A1(n10980), .A2(n7547), .B1(n9824), .B2(n10977), .C1(
        n9826), .C2(n10975), .ZN(n7560) );
  INV_X1 U8725 ( .A(n7560), .ZN(n7548) );
  AOI21_X1 U8726 ( .B1(n7557), .B2(n9958), .A(n7548), .ZN(n7556) );
  INV_X1 U8727 ( .A(n7549), .ZN(n7550) );
  OAI22_X1 U8728 ( .A1(n10022), .A2(n7551), .B1(n7550), .B2(n10741), .ZN(n7554) );
  OAI21_X1 U8729 ( .B1(n5126), .B2(n7446), .A(n7552), .ZN(n7561) );
  NOR2_X1 U8730 ( .A1(n7561), .A2(n10070), .ZN(n7553) );
  AOI211_X1 U8731 ( .C1(n10996), .C2(n7558), .A(n7554), .B(n7553), .ZN(n7555)
         );
  OAI21_X1 U8732 ( .B1(n7556), .B2(n10738), .A(n7555), .ZN(P1_U3286) );
  INV_X1 U8733 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7563) );
  AND2_X1 U8734 ( .A1(n7169), .A2(n10875), .ZN(n10539) );
  AOI21_X1 U8735 ( .B1(n10873), .B2(n7558), .A(n7557), .ZN(n7559) );
  OAI211_X1 U8736 ( .C1(n10539), .C2(n7561), .A(n7560), .B(n7559), .ZN(n7564)
         );
  NAND2_X1 U8737 ( .A1(n7564), .A2(n10993), .ZN(n7562) );
  OAI21_X1 U8738 ( .B1(n10993), .B2(n7563), .A(n7562), .ZN(P1_U3469) );
  NAND2_X1 U8739 ( .A1(n7564), .A2(n10989), .ZN(n7565) );
  OAI21_X1 U8740 ( .B1(n10989), .B2(n6762), .A(n7565), .ZN(P1_U3528) );
  AND2_X1 U8741 ( .A1(n9220), .A2(n9101), .ZN(n9203) );
  AOI22_X1 U8742 ( .A1(n9203), .A2(n6436), .B1(n9220), .B2(n5713), .ZN(n7569)
         );
  INV_X1 U8743 ( .A(n9182), .ZN(n7568) );
  NOR3_X1 U8744 ( .A1(n7569), .A2(n7568), .A3(n7567), .ZN(n7576) );
  OAI22_X1 U8745 ( .A1(n9229), .A2(n6445), .B1(n5042), .B2(n7570), .ZN(n7575)
         );
  OR2_X1 U8746 ( .A1(n7572), .A2(n7571), .ZN(n9181) );
  AOI22_X1 U8747 ( .A1(n9248), .A2(n7728), .B1(n9181), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n7573) );
  OAI21_X1 U8748 ( .B1(n9230), .B2(n6434), .A(n7573), .ZN(n7574) );
  OR3_X1 U8749 ( .A1(n7576), .A2(n7575), .A3(n7574), .ZN(P2_U3239) );
  NAND2_X1 U8750 ( .A1(n9248), .A2(n10821), .ZN(n7579) );
  INV_X1 U8751 ( .A(n7577), .ZN(n7578) );
  NAND2_X1 U8752 ( .A1(n7579), .A2(n7578), .ZN(n7581) );
  OAI22_X1 U8753 ( .A1(n9562), .A2(n9230), .B1(n9229), .B2(n9560), .ZN(n7580)
         );
  AOI211_X1 U8754 ( .C1(n9567), .C2(n9246), .A(n7581), .B(n7580), .ZN(n7587)
         );
  INV_X1 U8755 ( .A(n9203), .ZN(n9240) );
  OAI22_X1 U8756 ( .A1(n9240), .A2(n9562), .B1(n5042), .B2(n7582), .ZN(n7585)
         );
  INV_X1 U8757 ( .A(n7583), .ZN(n7584) );
  NAND3_X1 U8758 ( .A1(n7585), .A2(n8788), .A3(n7584), .ZN(n7586) );
  OAI211_X1 U8759 ( .C1(n5042), .C2(n7588), .A(n7587), .B(n7586), .ZN(P2_U3241) );
  INV_X1 U8760 ( .A(n7813), .ZN(n10830) );
  OAI22_X1 U8761 ( .A1(n9099), .A2(n10830), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7589), .ZN(n7591) );
  OAI22_X1 U8762 ( .A1(n7603), .A2(n9229), .B1(n9230), .B2(n8777), .ZN(n7590)
         );
  AOI211_X1 U8763 ( .C1(n7812), .C2(n9246), .A(n7591), .B(n7590), .ZN(n7596)
         );
  AOI21_X1 U8764 ( .B1(n7593), .B2(n7592), .A(n5042), .ZN(n7594) );
  NAND2_X1 U8765 ( .A1(n7594), .A2(n7643), .ZN(n7595) );
  NAND2_X1 U8766 ( .A1(n7596), .A2(n7595), .ZN(P2_U3215) );
  NAND2_X1 U8767 ( .A1(n9248), .A2(n10863), .ZN(n7599) );
  INV_X1 U8768 ( .A(n7597), .ZN(n7598) );
  NAND2_X1 U8769 ( .A1(n7599), .A2(n7598), .ZN(n7601) );
  OAI22_X1 U8770 ( .A1(n7603), .A2(n9230), .B1(n9229), .B2(n9239), .ZN(n7600)
         );
  AOI211_X1 U8771 ( .C1(n7952), .C2(n9246), .A(n7601), .B(n7600), .ZN(n7610)
         );
  INV_X1 U8772 ( .A(n7603), .ZN(n9277) );
  NAND3_X1 U8773 ( .A1(n9203), .A2(n7604), .A3(n9277), .ZN(n7605) );
  OAI21_X1 U8774 ( .B1(n7645), .B2(n5042), .A(n7605), .ZN(n7608) );
  INV_X1 U8775 ( .A(n7606), .ZN(n7607) );
  NAND2_X1 U8776 ( .A1(n7608), .A2(n7607), .ZN(n7609) );
  OAI211_X1 U8777 ( .C1(n5042), .C2(n7611), .A(n7610), .B(n7609), .ZN(P2_U3233) );
  NAND2_X1 U8778 ( .A1(n7613), .A2(n7612), .ZN(n7614) );
  AND2_X1 U8779 ( .A1(n7615), .A2(n7614), .ZN(n7625) );
  OAI21_X1 U8780 ( .B1(n7618), .B2(n7617), .A(n7616), .ZN(n7619) );
  AOI22_X1 U8781 ( .A1(n10666), .A2(n7619), .B1(n10679), .B2(
        P1_ADDR_REG_14__SCAN_IN), .ZN(n7624) );
  INV_X1 U8782 ( .A(n8243), .ZN(n7621) );
  NAND2_X1 U8783 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3084), .ZN(n7620) );
  OAI21_X1 U8784 ( .B1(n10677), .B2(n7621), .A(n7620), .ZN(n7622) );
  INV_X1 U8785 ( .A(n7622), .ZN(n7623) );
  OAI211_X1 U8786 ( .C1(n7625), .C2(n9890), .A(n7624), .B(n7623), .ZN(P1_U3255) );
  INV_X1 U8787 ( .A(n8466), .ZN(n7640) );
  OAI222_X1 U8788 ( .A1(P1_U3084), .A2(n7627), .B1(n5044), .B2(n7640), .C1(
        n7626), .C2(n8399), .ZN(P1_U3336) );
  OAI21_X1 U8789 ( .B1(n7630), .B2(n7629), .A(n7628), .ZN(n7638) );
  NAND2_X1 U8790 ( .A1(n10679), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n7631) );
  NAND2_X1 U8791 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8282) );
  OAI211_X1 U8792 ( .C1(n10677), .C2(n7632), .A(n7631), .B(n8282), .ZN(n7637)
         );
  AOI211_X1 U8793 ( .C1(n7635), .C2(n7634), .A(n7633), .B(n9890), .ZN(n7636)
         );
  AOI211_X1 U8794 ( .C1(n10666), .C2(n7638), .A(n7637), .B(n7636), .ZN(n7639)
         );
  INV_X1 U8795 ( .A(n7639), .ZN(P1_U3254) );
  INV_X1 U8796 ( .A(n9339), .ZN(n9331) );
  OAI222_X1 U8797 ( .A1(P2_U3152), .A2(n9331), .B1(n9698), .B2(n6054), .C1(
        n7640), .C2(n5043), .ZN(P2_U3341) );
  INV_X1 U8798 ( .A(n7768), .ZN(n7655) );
  INV_X1 U8799 ( .A(n7641), .ZN(n7642) );
  AOI21_X1 U8800 ( .B1(n7643), .B2(n7642), .A(n5042), .ZN(n7647) );
  NOR3_X1 U8801 ( .A1(n9240), .A2(n9560), .A3(n7644), .ZN(n7646) );
  OAI21_X1 U8802 ( .B1(n7647), .B2(n7646), .A(n7645), .ZN(n7654) );
  INV_X1 U8803 ( .A(n9257), .ZN(n7651) );
  OR2_X1 U8804 ( .A1(n7986), .A2(n9559), .ZN(n7649) );
  OR2_X1 U8805 ( .A1(n9560), .A2(n9561), .ZN(n7648) );
  AND2_X1 U8806 ( .A1(n7649), .A2(n7648), .ZN(n7764) );
  OAI22_X1 U8807 ( .A1(n7651), .A2(n7764), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7650), .ZN(n7652) );
  AOI21_X1 U8808 ( .B1(n7943), .B2(n9261), .A(n7652), .ZN(n7653) );
  OAI211_X1 U8809 ( .C1(n9259), .C2(n7655), .A(n7654), .B(n7653), .ZN(P2_U3223) );
  INV_X1 U8810 ( .A(n7656), .ZN(n7658) );
  NAND2_X1 U8811 ( .A1(n7658), .A2(n7657), .ZN(n7659) );
  NOR2_X1 U8812 ( .A1(n10803), .A2(n6980), .ZN(n7662) );
  OR2_X1 U8813 ( .A1(n7659), .A2(n9101), .ZN(n9363) );
  INV_X1 U8814 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10210) );
  OAI22_X1 U8815 ( .A1(n9363), .A2(n7660), .B1(n10210), .B2(n9549), .ZN(n7661)
         );
  AOI211_X1 U8816 ( .C1(n10803), .C2(n7663), .A(n7662), .B(n7661), .ZN(n7668)
         );
  OR2_X1 U8817 ( .A1(n7665), .A2(n5697), .ZN(n7727) );
  NAND2_X1 U8818 ( .A1(n9544), .A2(n7727), .ZN(n10802) );
  NAND2_X1 U8819 ( .A1(n10803), .A2(n10802), .ZN(n9533) );
  INV_X1 U8820 ( .A(n9533), .ZN(n9572) );
  NAND2_X1 U8821 ( .A1(n10803), .A2(n10796), .ZN(n9547) );
  AOI22_X1 U8822 ( .A1(n9572), .A2(n7666), .B1(n9573), .B2(n6433), .ZN(n7667)
         );
  NAND2_X1 U8823 ( .A1(n7668), .A2(n7667), .ZN(P2_U3295) );
  XNOR2_X1 U8824 ( .A(n7670), .B(n7669), .ZN(n7671) );
  NAND2_X1 U8825 ( .A1(n7671), .A2(n10794), .ZN(n7673) );
  AOI22_X1 U8826 ( .A1(n10791), .A2(n10790), .B1(n9281), .B2(n10789), .ZN(
        n7672) );
  AND2_X1 U8827 ( .A1(n7673), .A2(n7672), .ZN(n10761) );
  NAND2_X1 U8828 ( .A1(n6434), .A2(n7674), .ZN(n7675) );
  NAND2_X1 U8829 ( .A1(n7676), .A2(n7675), .ZN(n7715) );
  NAND2_X1 U8830 ( .A1(n7715), .A2(n7714), .ZN(n7717) );
  NAND2_X1 U8831 ( .A1(n7677), .A2(n10752), .ZN(n7678) );
  OAI21_X1 U8832 ( .B1(n7680), .B2(n7679), .A(n7749), .ZN(n10764) );
  AOI22_X1 U8833 ( .A1(n9572), .A2(n10764), .B1(n9573), .B2(n7681), .ZN(n7684)
         );
  OAI21_X1 U8834 ( .B1(n7710), .B2(n10759), .A(n7752), .ZN(n10760) );
  OAI22_X1 U8835 ( .A1(n9363), .A2(n10760), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9549), .ZN(n7682) );
  AOI21_X1 U8836 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n7664), .A(n7682), .ZN(
        n7683) );
  OAI211_X1 U8837 ( .C1(n7664), .C2(n10761), .A(n7684), .B(n7683), .ZN(
        P2_U3293) );
  INV_X1 U8838 ( .A(n9804), .ZN(n9795) );
  NAND2_X1 U8839 ( .A1(n9823), .A2(n7104), .ZN(n7686) );
  NAND2_X1 U8840 ( .A1(n7702), .A2(n8795), .ZN(n7685) );
  NAND2_X1 U8841 ( .A1(n7686), .A2(n7685), .ZN(n7687) );
  XNOR2_X1 U8842 ( .A(n7687), .B(n8724), .ZN(n7827) );
  NAND2_X1 U8843 ( .A1(n9823), .A2(n8790), .ZN(n7689) );
  NAND2_X1 U8844 ( .A1(n7702), .A2(n5040), .ZN(n7688) );
  NAND2_X1 U8845 ( .A1(n7689), .A2(n7688), .ZN(n7825) );
  XNOR2_X1 U8846 ( .A(n7827), .B(n7825), .ZN(n7693) );
  OAI21_X1 U8847 ( .B1(n7693), .B2(n7692), .A(n7834), .ZN(n7694) );
  NAND2_X1 U8848 ( .A1(n7694), .A2(n9744), .ZN(n7698) );
  AOI22_X1 U8849 ( .A1(n9805), .A2(n9824), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3084), .ZN(n7695) );
  OAI21_X1 U8850 ( .B1(n7873), .B2(n9808), .A(n7695), .ZN(n7696) );
  AOI21_X1 U8851 ( .B1(n7702), .B2(n9811), .A(n7696), .ZN(n7697) );
  OAI211_X1 U8852 ( .C1(n9795), .C2(n7699), .A(n7698), .B(n7697), .ZN(P1_U3211) );
  INV_X1 U8853 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7706) );
  AOI211_X1 U8854 ( .C1(n10873), .C2(n7702), .A(n7701), .B(n7700), .ZN(n7703)
         );
  OAI21_X1 U8855 ( .B1(n10539), .B2(n7704), .A(n7703), .ZN(n7707) );
  NAND2_X1 U8856 ( .A1(n7707), .A2(n10993), .ZN(n7705) );
  OAI21_X1 U8857 ( .B1(n10993), .B2(n7706), .A(n7705), .ZN(P1_U3475) );
  NAND2_X1 U8858 ( .A1(n7707), .A2(n10989), .ZN(n7708) );
  OAI21_X1 U8859 ( .B1(n10989), .B2(n7709), .A(n7708), .ZN(P1_U3530) );
  AOI21_X1 U8860 ( .B1(n7728), .B2(n7711), .A(n7710), .ZN(n10751) );
  INV_X1 U8861 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10238) );
  NOR2_X1 U8862 ( .A1(n10238), .A2(n9549), .ZN(n7726) );
  INV_X1 U8863 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7724) );
  XNOR2_X1 U8864 ( .A(n7713), .B(n7712), .ZN(n7722) );
  OR2_X1 U8865 ( .A1(n7715), .A2(n7714), .ZN(n7716) );
  NAND2_X1 U8866 ( .A1(n7717), .A2(n7716), .ZN(n10756) );
  INV_X1 U8867 ( .A(n9544), .ZN(n7718) );
  NAND2_X1 U8868 ( .A1(n10756), .A2(n7718), .ZN(n7721) );
  OAI22_X1 U8869 ( .A1(n6434), .A2(n9561), .B1(n6445), .B2(n9559), .ZN(n7719)
         );
  INV_X1 U8870 ( .A(n7719), .ZN(n7720) );
  OAI211_X1 U8871 ( .C1(n9538), .C2(n7722), .A(n7721), .B(n7720), .ZN(n10754)
         );
  NAND2_X1 U8872 ( .A1(n10803), .A2(n10754), .ZN(n7723) );
  OAI21_X1 U8873 ( .B1(n10803), .B2(n7724), .A(n7723), .ZN(n7725) );
  AOI211_X1 U8874 ( .C1(n9568), .C2(n10751), .A(n7726), .B(n7725), .ZN(n7730)
         );
  NOR2_X1 U8875 ( .A1(n7664), .A2(n7727), .ZN(n9554) );
  AOI22_X1 U8876 ( .A1(n9554), .A2(n10756), .B1(n9573), .B2(n7728), .ZN(n7729)
         );
  NAND2_X1 U8877 ( .A1(n7730), .A2(n7729), .ZN(P2_U3294) );
  OAI22_X1 U8878 ( .A1(n9229), .A2(n8781), .B1(n10759), .B2(n9099), .ZN(n7735)
         );
  INV_X1 U8879 ( .A(n9217), .ZN(n7731) );
  AOI211_X1 U8880 ( .C1(n7733), .C2(n7732), .A(n7731), .B(n5042), .ZN(n7734)
         );
  AOI211_X1 U8881 ( .C1(n9247), .C2(n9281), .A(n7735), .B(n7734), .ZN(n7737)
         );
  MUX2_X1 U8882 ( .A(n9259), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n7736) );
  NAND2_X1 U8883 ( .A1(n7737), .A2(n7736), .ZN(P2_U3220) );
  AOI22_X1 U8884 ( .A1(n10743), .A2(n10794), .B1(n10791), .B2(n6436), .ZN(
        n10745) );
  INV_X1 U8885 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10225) );
  OAI22_X1 U8886 ( .A1(n7664), .A2(n10745), .B1(n10225), .B2(n9549), .ZN(n7738) );
  AOI21_X1 U8887 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n7664), .A(n7738), .ZN(
        n7740) );
  OAI21_X1 U8888 ( .B1(n9573), .B2(n9568), .A(n10742), .ZN(n7739) );
  OAI211_X1 U8889 ( .C1(n7741), .C2(n9533), .A(n7740), .B(n7739), .ZN(P2_U3296) );
  OAI211_X1 U8890 ( .C1(n7744), .C2(n7743), .A(n7742), .B(n10794), .ZN(n7747)
         );
  OAI22_X1 U8891 ( .A1(n9562), .A2(n9559), .B1(n6445), .B2(n9561), .ZN(n7745)
         );
  INV_X1 U8892 ( .A(n7745), .ZN(n7746) );
  NAND2_X1 U8893 ( .A1(n7747), .A2(n7746), .ZN(n10777) );
  INV_X1 U8894 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7758) );
  NAND2_X1 U8895 ( .A1(n6445), .A2(n10759), .ZN(n7748) );
  OAI21_X1 U8896 ( .B1(n7751), .B2(n7750), .A(n7773), .ZN(n10779) );
  AOI22_X1 U8897 ( .A1(n9572), .A2(n10779), .B1(n9573), .B2(n9214), .ZN(n7757)
         );
  NAND2_X1 U8898 ( .A1(n7752), .A2(n9214), .ZN(n7753) );
  AND2_X1 U8899 ( .A1(n10783), .A2(n7753), .ZN(n10774) );
  NOR2_X1 U8900 ( .A1(n7754), .A2(n9549), .ZN(n7755) );
  AOI21_X1 U8901 ( .B1(n9568), .B2(n10774), .A(n7755), .ZN(n7756) );
  OAI211_X1 U8902 ( .C1(n7758), .C2(n10803), .A(n7757), .B(n7756), .ZN(n7759)
         );
  AOI21_X1 U8903 ( .B1(n10803), .B2(n10777), .A(n7759), .ZN(n7760) );
  INV_X1 U8904 ( .A(n7760), .ZN(P2_U3292) );
  INV_X1 U8905 ( .A(n8636), .ZN(n7853) );
  AOI22_X1 U8906 ( .A1(n9347), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n7761), .ZN(n7762) );
  OAI21_X1 U8907 ( .B1(n7853), .B2(n5043), .A(n7762), .ZN(P2_U3340) );
  XOR2_X1 U8908 ( .A(n7763), .B(n7779), .Z(n7765) );
  OAI21_X1 U8909 ( .B1(n7765), .B2(n9538), .A(n7764), .ZN(n10851) );
  INV_X1 U8910 ( .A(n10851), .ZN(n7783) );
  AND2_X1 U8911 ( .A1(n10803), .A2(n9546), .ZN(n9426) );
  AND2_X1 U8912 ( .A1(n10786), .A2(n7766), .ZN(n9565) );
  INV_X1 U8913 ( .A(n7811), .ZN(n7767) );
  INV_X1 U8914 ( .A(n7943), .ZN(n10849) );
  OAI211_X1 U8915 ( .C1(n7767), .C2(n10849), .A(n10940), .B(n7992), .ZN(n10847) );
  INV_X1 U8916 ( .A(n10847), .ZN(n7771) );
  INV_X1 U8917 ( .A(n9549), .ZN(n10798) );
  AOI22_X1 U8918 ( .A1(n7664), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n7768), .B2(
        n10798), .ZN(n7769) );
  OAI21_X1 U8919 ( .B1(n10849), .B2(n9547), .A(n7769), .ZN(n7770) );
  AOI21_X1 U8920 ( .B1(n9426), .B2(n7771), .A(n7770), .ZN(n7782) );
  NAND2_X1 U8921 ( .A1(n9562), .A2(n10808), .ZN(n7774) );
  INV_X1 U8922 ( .A(n9570), .ZN(n7776) );
  INV_X1 U8923 ( .A(n9571), .ZN(n7775) );
  NAND2_X1 U8924 ( .A1(n7776), .A2(n7775), .ZN(n9569) );
  INV_X1 U8925 ( .A(n9560), .ZN(n9278) );
  OR2_X1 U8926 ( .A1(n7813), .A2(n9278), .ZN(n7778) );
  NAND2_X1 U8927 ( .A1(n7780), .A2(n7779), .ZN(n10845) );
  NAND3_X1 U8928 ( .A1(n10846), .A2(n10845), .A3(n9572), .ZN(n7781) );
  OAI211_X1 U8929 ( .C1(n7783), .C2(n7664), .A(n7782), .B(n7781), .ZN(P2_U3288) );
  INV_X1 U8930 ( .A(n10710), .ZN(n10724) );
  INV_X1 U8931 ( .A(n10726), .ZN(n9355) );
  INV_X1 U8932 ( .A(n9285), .ZN(n7786) );
  INV_X1 U8933 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10907) );
  MUX2_X1 U8934 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10907), .S(n9285), .Z(n9288) );
  OAI21_X1 U8935 ( .B1(n7785), .B2(n7385), .A(n7784), .ZN(n9289) );
  NAND2_X1 U8936 ( .A1(n9288), .A2(n9289), .ZN(n9287) );
  OAI21_X1 U8937 ( .B1(n7786), .B2(n10907), .A(n9287), .ZN(n7789) );
  INV_X1 U8938 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7787) );
  MUX2_X1 U8939 ( .A(n7787), .B(P2_REG1_REG_12__SCAN_IN), .S(n7907), .Z(n7788)
         );
  NOR2_X1 U8940 ( .A1(n7788), .A2(n7789), .ZN(n7902) );
  AOI21_X1 U8941 ( .B1(n7789), .B2(n7788), .A(n7902), .ZN(n7792) );
  NOR2_X1 U8942 ( .A1(n7790), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8003) );
  AOI21_X1 U8943 ( .B1(n10718), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8003), .ZN(
        n7791) );
  OAI21_X1 U8944 ( .B1(n9355), .B2(n7792), .A(n7791), .ZN(n7801) );
  INV_X1 U8945 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7795) );
  MUX2_X1 U8946 ( .A(n7795), .B(P2_REG2_REG_11__SCAN_IN), .S(n9285), .Z(n7796)
         );
  INV_X1 U8947 ( .A(n7796), .ZN(n9283) );
  OAI21_X1 U8948 ( .B1(n9285), .B2(P2_REG2_REG_11__SCAN_IN), .A(n9282), .ZN(
        n7799) );
  INV_X1 U8949 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7797) );
  MUX2_X1 U8950 ( .A(n7797), .B(P2_REG2_REG_12__SCAN_IN), .S(n7907), .Z(n7798)
         );
  NOR2_X1 U8951 ( .A1(n7798), .A2(n7799), .ZN(n7906) );
  AOI211_X1 U8952 ( .C1(n7799), .C2(n7798), .A(n7906), .B(n10719), .ZN(n7800)
         );
  AOI211_X1 U8953 ( .C1(n10724), .C2(n7907), .A(n7801), .B(n7800), .ZN(n7802)
         );
  INV_X1 U8954 ( .A(n7802), .ZN(P2_U3257) );
  XNOR2_X1 U8955 ( .A(n7803), .B(n7807), .ZN(n7804) );
  NAND2_X1 U8956 ( .A1(n7804), .A2(n10794), .ZN(n7806) );
  AOI22_X1 U8957 ( .A1(n9277), .A2(n10791), .B1(n10789), .B2(n10792), .ZN(
        n7805) );
  NAND2_X1 U8958 ( .A1(n7806), .A2(n7805), .ZN(n10832) );
  INV_X1 U8959 ( .A(n10832), .ZN(n7818) );
  INV_X1 U8960 ( .A(n7807), .ZN(n7809) );
  OR2_X1 U8961 ( .A1(n9565), .A2(n10830), .ZN(n7810) );
  NAND2_X1 U8962 ( .A1(n7811), .A2(n7810), .ZN(n10831) );
  AOI22_X1 U8963 ( .A1(n7664), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n7812), .B2(
        n10798), .ZN(n7815) );
  NAND2_X1 U8964 ( .A1(n9573), .A2(n7813), .ZN(n7814) );
  OAI211_X1 U8965 ( .C1(n10831), .C2(n9363), .A(n7815), .B(n7814), .ZN(n7816)
         );
  AOI21_X1 U8966 ( .B1(n10834), .B2(n9572), .A(n7816), .ZN(n7817) );
  OAI21_X1 U8967 ( .B1(n7664), .B2(n7818), .A(n7817), .ZN(P2_U3289) );
  NAND2_X1 U8968 ( .A1(n7819), .A2(n8749), .ZN(n7822) );
  AOI22_X1 U8969 ( .A1(n8638), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8637), .B2(
        n7820), .ZN(n7821) );
  NAND2_X1 U8970 ( .A1(n9822), .A2(n7104), .ZN(n7823) );
  OAI21_X1 U8971 ( .B1(n7898), .B2(n8716), .A(n7823), .ZN(n7824) );
  XNOR2_X1 U8972 ( .A(n7824), .B(n8793), .ZN(n7963) );
  INV_X1 U8973 ( .A(n7825), .ZN(n7826) );
  NAND2_X1 U8974 ( .A1(n7827), .A2(n7826), .ZN(n7832) );
  OR2_X1 U8975 ( .A1(n7898), .A2(n7961), .ZN(n7829) );
  NAND2_X1 U8976 ( .A1(n9822), .A2(n8790), .ZN(n7828) );
  AND2_X1 U8977 ( .A1(n7829), .A2(n7828), .ZN(n7830) );
  INV_X1 U8978 ( .A(n7830), .ZN(n7831) );
  AND2_X1 U8979 ( .A1(n7832), .A2(n7831), .ZN(n7833) );
  NAND2_X1 U8980 ( .A1(n7834), .A2(n7833), .ZN(n7965) );
  NAND2_X1 U8981 ( .A1(n7964), .A2(n7965), .ZN(n7835) );
  XOR2_X1 U8982 ( .A(n7963), .B(n7835), .Z(n7842) );
  INV_X1 U8983 ( .A(n7898), .ZN(n10837) );
  INV_X1 U8984 ( .A(n7836), .ZN(n7897) );
  NOR2_X1 U8985 ( .A1(n9794), .A2(n7888), .ZN(n7837) );
  AOI211_X1 U8986 ( .C1(n9798), .C2(n8120), .A(n7838), .B(n7837), .ZN(n7839)
         );
  OAI21_X1 U8987 ( .B1(n9795), .B2(n7897), .A(n7839), .ZN(n7840) );
  AOI21_X1 U8988 ( .B1(n10837), .B2(n9811), .A(n7840), .ZN(n7841) );
  OAI21_X1 U8989 ( .B1(n7842), .B2(n9813), .A(n7841), .ZN(P1_U3219) );
  INV_X1 U8990 ( .A(n9237), .ZN(n7843) );
  AOI211_X1 U8991 ( .C1(n7845), .C2(n7844), .A(n5042), .B(n7843), .ZN(n7849)
         );
  INV_X1 U8992 ( .A(n8075), .ZN(n9274) );
  AOI22_X1 U8993 ( .A1(n9244), .A2(n9274), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3152), .ZN(n7847) );
  INV_X1 U8994 ( .A(n7986), .ZN(n9276) );
  AOI22_X1 U8995 ( .A1(n9247), .A2(n9276), .B1(n9246), .B2(n7990), .ZN(n7846)
         );
  OAI211_X1 U8996 ( .C1(n5299), .C2(n9099), .A(n7847), .B(n7846), .ZN(n7848)
         );
  OR2_X1 U8997 ( .A1(n7849), .A2(n7848), .ZN(P2_U3219) );
  NAND2_X1 U8998 ( .A1(n7850), .A2(n10318), .ZN(n7851) );
  NAND2_X1 U8999 ( .A1(n7851), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7852) );
  XNOR2_X1 U9000 ( .A(n7852), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9882) );
  INV_X1 U9001 ( .A(n9882), .ZN(n9866) );
  INV_X1 U9002 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10274) );
  OAI222_X1 U9003 ( .A1(n9866), .A2(P1_U3084), .B1(n5044), .B2(n7853), .C1(
        n10274), .C2(n8399), .ZN(P1_U3335) );
  NAND2_X1 U9004 ( .A1(n7888), .A2(n7854), .ZN(n7855) );
  NAND2_X1 U9005 ( .A1(n7898), .A2(n9822), .ZN(n8892) );
  NAND2_X1 U9006 ( .A1(n7873), .A2(n10837), .ZN(n8891) );
  NAND2_X1 U9007 ( .A1(n10837), .A2(n9822), .ZN(n7858) );
  NAND2_X1 U9008 ( .A1(n7859), .A2(n8749), .ZN(n7862) );
  AOI22_X1 U9009 ( .A1(n8638), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8637), .B2(
        n7860), .ZN(n7861) );
  INV_X1 U9010 ( .A(n8120), .ZN(n7937) );
  OR2_X1 U9011 ( .A1(n7974), .A2(n7937), .ZN(n8898) );
  NAND2_X1 U9012 ( .A1(n7974), .A2(n7937), .ZN(n8897) );
  NAND2_X1 U9013 ( .A1(n8898), .A2(n8897), .ZN(n8998) );
  XNOR2_X1 U9014 ( .A(n7918), .B(n8998), .ZN(n7877) );
  NAND2_X1 U9015 ( .A1(n9020), .A2(n8889), .ZN(n7864) );
  NAND2_X1 U9016 ( .A1(n7864), .A2(n9002), .ZN(n7932) );
  NAND2_X1 U9017 ( .A1(n7932), .A2(n8891), .ZN(n7865) );
  INV_X1 U9018 ( .A(n8998), .ZN(n8894) );
  XNOR2_X1 U9019 ( .A(n7865), .B(n8894), .ZN(n7875) );
  NAND2_X1 U9020 ( .A1(n7351), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7872) );
  NAND2_X1 U9021 ( .A1(n7867), .A2(n7866), .ZN(n7868) );
  AND2_X1 U9022 ( .A1(n7923), .A2(n7868), .ZN(n8118) );
  NAND2_X1 U9023 ( .A1(n7099), .A2(n8118), .ZN(n7871) );
  NAND2_X1 U9024 ( .A1(n5051), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7870) );
  NAND2_X1 U9025 ( .A1(n5039), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7869) );
  NAND4_X1 U9026 ( .A1(n7872), .A2(n7871), .A3(n7870), .A4(n7869), .ZN(n9821)
         );
  INV_X1 U9027 ( .A(n9821), .ZN(n7973) );
  OAI22_X1 U9028 ( .A1(n7873), .A2(n10013), .B1(n7973), .B2(n10015), .ZN(n7874) );
  AOI21_X1 U9029 ( .B1(n7875), .B2(n10980), .A(n7874), .ZN(n7876) );
  OAI21_X1 U9030 ( .B1(n7877), .B2(n7169), .A(n7876), .ZN(n10856) );
  INV_X1 U9031 ( .A(n10856), .ZN(n7883) );
  INV_X1 U9032 ( .A(n7877), .ZN(n10858) );
  NAND2_X1 U9033 ( .A1(n7893), .A2(n7898), .ZN(n7894) );
  NAND2_X1 U9034 ( .A1(n7894), .A2(n7974), .ZN(n7878) );
  NAND2_X1 U9035 ( .A1(n7938), .A2(n7878), .ZN(n10855) );
  AOI22_X1 U9036 ( .A1(n10738), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7977), .B2(
        n10994), .ZN(n7880) );
  NAND2_X1 U9037 ( .A1(n10996), .A2(n7974), .ZN(n7879) );
  OAI211_X1 U9038 ( .C1(n10855), .C2(n10733), .A(n7880), .B(n7879), .ZN(n7881)
         );
  AOI21_X1 U9039 ( .B1(n10858), .B2(n9929), .A(n7881), .ZN(n7882) );
  OAI21_X1 U9040 ( .B1(n7883), .B2(n10738), .A(n7882), .ZN(P1_U3282) );
  INV_X1 U9041 ( .A(n7884), .ZN(n7885) );
  AOI21_X1 U9042 ( .B1(n9002), .B2(n7886), .A(n7885), .ZN(n7891) );
  INV_X1 U9043 ( .A(n7891), .ZN(n10841) );
  NAND3_X1 U9044 ( .A1(n9020), .A2(n7857), .A3(n8889), .ZN(n7887) );
  AOI21_X1 U9045 ( .B1(n7932), .B2(n7887), .A(n9131), .ZN(n7890) );
  OAI22_X1 U9046 ( .A1(n7888), .A2(n10013), .B1(n7937), .B2(n10015), .ZN(n7889) );
  AOI211_X1 U9047 ( .C1(n7891), .C2(n10879), .A(n7890), .B(n7889), .ZN(n10840)
         );
  MUX2_X1 U9048 ( .A(n7892), .B(n10840), .S(n10022), .Z(n7901) );
  INV_X1 U9049 ( .A(n7893), .ZN(n7896) );
  INV_X1 U9050 ( .A(n7894), .ZN(n7895) );
  AOI21_X1 U9051 ( .B1(n10837), .B2(n7896), .A(n7895), .ZN(n10838) );
  OAI22_X1 U9052 ( .A1(n10734), .A2(n7898), .B1(n7897), .B2(n10741), .ZN(n7899) );
  AOI21_X1 U9053 ( .B1(n10838), .B2(n10068), .A(n7899), .ZN(n7900) );
  OAI211_X1 U9054 ( .C1(n10841), .C2(n10029), .A(n7901), .B(n7900), .ZN(
        P1_U3283) );
  AOI21_X1 U9055 ( .B1(n7903), .B2(n7787), .A(n7902), .ZN(n7905) );
  INV_X1 U9056 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10946) );
  AOI22_X1 U9057 ( .A1(n8051), .A2(n10946), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n8046), .ZN(n7904) );
  NOR2_X1 U9058 ( .A1(n7905), .A2(n7904), .ZN(n8045) );
  AOI21_X1 U9059 ( .B1(n7905), .B2(n7904), .A(n8045), .ZN(n7915) );
  NOR2_X1 U9060 ( .A1(n8051), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7908) );
  AOI21_X1 U9061 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n8051), .A(n7908), .ZN(
        n7909) );
  OAI21_X1 U9062 ( .B1(n7910), .B2(n7909), .A(n8050), .ZN(n7911) );
  INV_X1 U9063 ( .A(n10719), .ZN(n10696) );
  NAND2_X1 U9064 ( .A1(n7911), .A2(n10696), .ZN(n7914) );
  INV_X1 U9065 ( .A(n10718), .ZN(n8056) );
  INV_X1 U9066 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8335) );
  NAND2_X1 U9067 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3152), .ZN(n8562) );
  OAI21_X1 U9068 ( .B1(n8056), .B2(n8335), .A(n8562), .ZN(n7912) );
  AOI21_X1 U9069 ( .B1(n8051), .B2(n10724), .A(n7912), .ZN(n7913) );
  OAI211_X1 U9070 ( .C1(n7915), .C2(n9355), .A(n7914), .B(n7913), .ZN(P2_U3258) );
  INV_X1 U9071 ( .A(n8610), .ZN(n7917) );
  OAI222_X1 U9072 ( .A1(n9698), .A2(n7916), .B1(n5043), .B2(n7917), .C1(n9546), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI222_X1 U9073 ( .A1(P1_U3084), .A2(n9958), .B1(n5044), .B2(n7917), .C1(
        n10272), .C2(n8399), .ZN(P1_U3334) );
  NAND2_X1 U9074 ( .A1(n7919), .A2(n8749), .ZN(n7921) );
  AOI22_X1 U9075 ( .A1(n8638), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n8637), .B2(
        n10662), .ZN(n7920) );
  OR2_X1 U9076 ( .A1(n10872), .A2(n7973), .ZN(n8901) );
  NAND2_X1 U9077 ( .A1(n10872), .A2(n7973), .ZN(n8902) );
  NAND2_X1 U9078 ( .A1(n8901), .A2(n8902), .ZN(n8013) );
  INV_X1 U9079 ( .A(n8013), .ZN(n9003) );
  XNOR2_X1 U9080 ( .A(n8014), .B(n9003), .ZN(n10876) );
  NAND2_X1 U9081 ( .A1(n7923), .A2(n7922), .ZN(n7924) );
  AND2_X1 U9082 ( .A1(n7925), .A2(n7924), .ZN(n8165) );
  NAND2_X1 U9083 ( .A1(n7099), .A2(n8165), .ZN(n7929) );
  NAND2_X1 U9084 ( .A1(n7351), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7928) );
  NAND2_X1 U9085 ( .A1(n5051), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7927) );
  NAND2_X1 U9086 ( .A1(n5039), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7926) );
  NAND4_X1 U9087 ( .A1(n7929), .A2(n7928), .A3(n7927), .A4(n7926), .ZN(n9820)
         );
  INV_X1 U9088 ( .A(n9820), .ZN(n8147) );
  INV_X1 U9089 ( .A(n8891), .ZN(n7930) );
  NOR2_X1 U9090 ( .A1(n8998), .A2(n7930), .ZN(n7931) );
  NAND2_X1 U9091 ( .A1(n7932), .A2(n7931), .ZN(n7933) );
  INV_X1 U9092 ( .A(n8019), .ZN(n7934) );
  AOI21_X1 U9093 ( .B1(n8013), .B2(n7935), .A(n7934), .ZN(n7936) );
  OAI222_X1 U9094 ( .A1(n10015), .A2(n8147), .B1(n10013), .B2(n7937), .C1(
        n9131), .C2(n7936), .ZN(n10870) );
  AOI211_X1 U9095 ( .C1(n10872), .C2(n7938), .A(n10960), .B(n8023), .ZN(n10871) );
  NAND2_X1 U9096 ( .A1(n10871), .A2(n10999), .ZN(n7940) );
  AOI22_X1 U9097 ( .A1(n11006), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n8118), .B2(
        n10994), .ZN(n7939) );
  OAI211_X1 U9098 ( .C1(n5310), .C2(n10734), .A(n7940), .B(n7939), .ZN(n7941)
         );
  AOI21_X1 U9099 ( .B1(n10870), .B2(n10022), .A(n7941), .ZN(n7942) );
  OAI21_X1 U9100 ( .B1(n10070), .B2(n10876), .A(n7942), .ZN(P1_U3281) );
  NAND2_X1 U9101 ( .A1(n7943), .A2(n9277), .ZN(n7944) );
  INV_X1 U9102 ( .A(n7982), .ZN(n7945) );
  AOI21_X1 U9103 ( .B1(n7948), .B2(n7946), .A(n7945), .ZN(n10862) );
  INV_X1 U9104 ( .A(n9554), .ZN(n7999) );
  INV_X1 U9105 ( .A(n9239), .ZN(n9275) );
  AOI22_X1 U9106 ( .A1(n10789), .A2(n9277), .B1(n9275), .B2(n10791), .ZN(n7951) );
  OAI211_X1 U9107 ( .C1(n7949), .C2(n7948), .A(n7947), .B(n10794), .ZN(n7950)
         );
  OAI211_X1 U9108 ( .C1(n10862), .C2(n9544), .A(n7951), .B(n7950), .ZN(n10865)
         );
  NAND2_X1 U9109 ( .A1(n10865), .A2(n10803), .ZN(n7957) );
  XNOR2_X1 U9110 ( .A(n7992), .B(n10863), .ZN(n10864) );
  NOR2_X1 U9111 ( .A1(n9363), .A2(n10864), .ZN(n7955) );
  INV_X1 U9112 ( .A(n7952), .ZN(n7953) );
  OAI22_X1 U9113 ( .A1(n10803), .A2(n7222), .B1(n7953), .B2(n9549), .ZN(n7954)
         );
  AOI211_X1 U9114 ( .C1(n9573), .C2(n10863), .A(n7955), .B(n7954), .ZN(n7956)
         );
  OAI211_X1 U9115 ( .C1(n10862), .C2(n7999), .A(n7957), .B(n7956), .ZN(
        P2_U3287) );
  NAND2_X1 U9116 ( .A1(n7974), .A2(n8795), .ZN(n7959) );
  NAND2_X1 U9117 ( .A1(n8120), .A2(n7104), .ZN(n7958) );
  NAND2_X1 U9118 ( .A1(n7959), .A2(n7958), .ZN(n7960) );
  XNOR2_X1 U9119 ( .A(n7960), .B(n8724), .ZN(n8108) );
  INV_X1 U9120 ( .A(n7961), .ZN(n8676) );
  AND2_X1 U9121 ( .A1(n8120), .A2(n8790), .ZN(n7962) );
  AOI21_X1 U9122 ( .B1(n7974), .B2(n8676), .A(n7962), .ZN(n8107) );
  XNOR2_X1 U9123 ( .A(n8108), .B(n8107), .ZN(n7970) );
  NAND2_X1 U9124 ( .A1(n7964), .A2(n7963), .ZN(n7966) );
  INV_X1 U9125 ( .A(n7970), .ZN(n7967) );
  INV_X1 U9126 ( .A(n8110), .ZN(n7968) );
  AOI21_X1 U9127 ( .B1(n7970), .B2(n7969), .A(n7968), .ZN(n7979) );
  NAND2_X1 U9128 ( .A1(n9805), .A2(n9822), .ZN(n7972) );
  OAI211_X1 U9129 ( .C1(n9808), .C2(n7973), .A(n7972), .B(n7971), .ZN(n7976)
         );
  INV_X1 U9130 ( .A(n7974), .ZN(n10854) );
  NOR2_X1 U9131 ( .A1(n9801), .A2(n10854), .ZN(n7975) );
  AOI211_X1 U9132 ( .C1(n7977), .C2(n9804), .A(n7976), .B(n7975), .ZN(n7978)
         );
  OAI21_X1 U9133 ( .B1(n7979), .B2(n9813), .A(n7978), .ZN(P1_U3229) );
  OR2_X1 U9134 ( .A1(n10863), .A2(n9276), .ZN(n7980) );
  AND2_X1 U9135 ( .A1(n7982), .A2(n7980), .ZN(n7984) );
  AND2_X1 U9136 ( .A1(n7983), .A2(n7980), .ZN(n7981) );
  NAND2_X1 U9137 ( .A1(n7982), .A2(n7981), .ZN(n8031) );
  OAI21_X1 U9138 ( .B1(n7984), .B2(n7983), .A(n8031), .ZN(n10883) );
  OAI21_X1 U9139 ( .B1(n5124), .B2(n6588), .A(n7985), .ZN(n7988) );
  OAI22_X1 U9140 ( .A1(n8075), .A2(n9559), .B1(n7986), .B2(n9561), .ZN(n7987)
         );
  AOI21_X1 U9141 ( .B1(n7988), .B2(n10794), .A(n7987), .ZN(n7989) );
  OAI21_X1 U9142 ( .B1(n10883), .B2(n9544), .A(n7989), .ZN(n10885) );
  NAND2_X1 U9143 ( .A1(n10885), .A2(n10803), .ZN(n7998) );
  INV_X1 U9144 ( .A(n7990), .ZN(n7991) );
  OAI22_X1 U9145 ( .A1(n10803), .A2(n7378), .B1(n7991), .B2(n9549), .ZN(n7996)
         );
  AND2_X1 U9146 ( .A1(n7993), .A2(n8029), .ZN(n7994) );
  OR2_X1 U9147 ( .A1(n7994), .A2(n8039), .ZN(n10884) );
  NOR2_X1 U9148 ( .A1(n10884), .A2(n9363), .ZN(n7995) );
  AOI211_X1 U9149 ( .C1(n9573), .C2(n8029), .A(n7996), .B(n7995), .ZN(n7997)
         );
  OAI211_X1 U9150 ( .C1(n10883), .C2(n7999), .A(n7998), .B(n7997), .ZN(
        P2_U3286) );
  INV_X1 U9151 ( .A(n9241), .ZN(n8002) );
  NOR3_X1 U9152 ( .A1(n9240), .A2(n8075), .A3(n8000), .ZN(n8001) );
  AOI21_X1 U9153 ( .B1(n8002), .B2(n9220), .A(n8001), .ZN(n8011) );
  INV_X1 U9154 ( .A(n8561), .ZN(n8009) );
  AOI22_X1 U9155 ( .A1(n9244), .A2(n9272), .B1(n9246), .B2(n8085), .ZN(n8007)
         );
  INV_X1 U9156 ( .A(n8003), .ZN(n8006) );
  NAND2_X1 U9157 ( .A1(n9248), .A2(n8095), .ZN(n8005) );
  NAND2_X1 U9158 ( .A1(n9247), .A2(n9274), .ZN(n8004) );
  NAND4_X1 U9159 ( .A1(n8007), .A2(n8006), .A3(n8005), .A4(n8004), .ZN(n8008)
         );
  AOI21_X1 U9160 ( .B1(n8009), .B2(n9220), .A(n8008), .ZN(n8010) );
  OAI21_X1 U9161 ( .B1(n8012), .B2(n8011), .A(n8010), .ZN(P2_U3226) );
  NAND2_X1 U9162 ( .A1(n8015), .A2(n8749), .ZN(n8018) );
  AOI22_X1 U9163 ( .A1(n8638), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8637), .B2(
        n8016), .ZN(n8017) );
  OR2_X1 U9164 ( .A1(n8170), .A2(n8147), .ZN(n8905) );
  NAND2_X1 U9165 ( .A1(n8170), .A2(n8147), .ZN(n8906) );
  NAND2_X1 U9166 ( .A1(n8905), .A2(n8906), .ZN(n9006) );
  XNOR2_X1 U9167 ( .A(n8131), .B(n9006), .ZN(n10894) );
  XNOR2_X1 U9168 ( .A(n8137), .B(n9006), .ZN(n8021) );
  AOI22_X1 U9169 ( .A1(n10975), .A2(n9821), .B1(n8284), .B2(n10977), .ZN(n8020) );
  OAI21_X1 U9170 ( .B1(n8021), .B2(n9131), .A(n8020), .ZN(n8022) );
  AOI21_X1 U9171 ( .B1(n10894), .B2(n10879), .A(n8022), .ZN(n10896) );
  INV_X1 U9172 ( .A(n8170), .ZN(n10891) );
  NOR2_X1 U9173 ( .A1(n8023), .A2(n10891), .ZN(n8024) );
  OR2_X1 U9174 ( .A1(n8150), .A2(n8024), .ZN(n10892) );
  AOI22_X1 U9175 ( .A1(n10738), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8165), .B2(
        n10994), .ZN(n8026) );
  NAND2_X1 U9176 ( .A1(n8170), .A2(n10996), .ZN(n8025) );
  OAI211_X1 U9177 ( .C1(n10892), .C2(n10733), .A(n8026), .B(n8025), .ZN(n8027)
         );
  AOI21_X1 U9178 ( .B1(n10894), .B2(n9929), .A(n8027), .ZN(n8028) );
  OAI21_X1 U9179 ( .B1(n10896), .B2(n11006), .A(n8028), .ZN(P1_U3280) );
  NAND2_X1 U9180 ( .A1(n8029), .A2(n9275), .ZN(n8030) );
  NAND2_X1 U9181 ( .A1(n8031), .A2(n8030), .ZN(n8033) );
  OAI21_X1 U9182 ( .B1(n8033), .B2(n8032), .A(n8080), .ZN(n10905) );
  XNOR2_X1 U9183 ( .A(n8035), .B(n8034), .ZN(n8037) );
  OAI22_X1 U9184 ( .A1(n8559), .A2(n9559), .B1(n9239), .B2(n9561), .ZN(n8036)
         );
  AOI21_X1 U9185 ( .B1(n8037), .B2(n10794), .A(n8036), .ZN(n10903) );
  INV_X1 U9186 ( .A(n8039), .ZN(n8040) );
  INV_X1 U9187 ( .A(n10901), .ZN(n8038) );
  AOI211_X1 U9188 ( .C1(n10901), .C2(n8040), .A(n10921), .B(n8083), .ZN(n10900) );
  AOI22_X1 U9189 ( .A1(n10900), .A2(n9546), .B1(n10798), .B2(n9245), .ZN(n8041) );
  AOI21_X1 U9190 ( .B1(n10903), .B2(n8041), .A(n7664), .ZN(n8042) );
  INV_X1 U9191 ( .A(n8042), .ZN(n8044) );
  AOI22_X1 U9192 ( .A1(n9573), .A2(n10901), .B1(n7664), .B2(
        P2_REG2_REG_11__SCAN_IN), .ZN(n8043) );
  OAI211_X1 U9193 ( .C1(n9533), .C2(n10905), .A(n8044), .B(n8043), .ZN(
        P2_U3285) );
  AOI21_X1 U9194 ( .B1(n8046), .B2(n10946), .A(n8045), .ZN(n8048) );
  INV_X1 U9195 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8206) );
  AOI22_X1 U9196 ( .A1(n8199), .A2(n8206), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n8207), .ZN(n8047) );
  NOR2_X1 U9197 ( .A1(n8048), .A2(n8047), .ZN(n8205) );
  AOI21_X1 U9198 ( .B1(n8048), .B2(n8047), .A(n8205), .ZN(n8060) );
  NOR2_X1 U9199 ( .A1(n8199), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8049) );
  AOI21_X1 U9200 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8199), .A(n8049), .ZN(
        n8053) );
  OAI21_X1 U9201 ( .B1(n8053), .B2(n8052), .A(n8198), .ZN(n8054) );
  NAND2_X1 U9202 ( .A1(n8054), .A2(n10696), .ZN(n8059) );
  INV_X1 U9203 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8055) );
  NAND2_X1 U9204 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8762) );
  OAI21_X1 U9205 ( .B1(n8056), .B2(n8055), .A(n8762), .ZN(n8057) );
  AOI21_X1 U9206 ( .B1(n8199), .B2(n10724), .A(n8057), .ZN(n8058) );
  OAI211_X1 U9207 ( .C1(n8060), .C2(n9355), .A(n8059), .B(n8058), .ZN(P2_U3259) );
  INV_X1 U9208 ( .A(n8651), .ZN(n8062) );
  OAI222_X1 U9209 ( .A1(P1_U3084), .A2(n8061), .B1(n5044), .B2(n8062), .C1(
        n8652), .C2(n8399), .ZN(P1_U3333) );
  OAI222_X1 U9210 ( .A1(P2_U3152), .A2(n8063), .B1(n5043), .B2(n8062), .C1(
        n9698), .C2(n6128), .ZN(P2_U3338) );
  AOI211_X1 U9211 ( .C1(n10965), .C2(n8065), .A(n8064), .B(n10684), .ZN(n8072)
         );
  AOI211_X1 U9212 ( .C1(n8068), .C2(n8067), .A(n8066), .B(n9890), .ZN(n8071)
         );
  NAND2_X1 U9213 ( .A1(n10679), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n8069) );
  NAND2_X1 U9214 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8548) );
  OAI211_X1 U9215 ( .C1(n10677), .C2(n8373), .A(n8069), .B(n8548), .ZN(n8070)
         );
  OR3_X1 U9216 ( .A1(n8072), .A2(n8071), .A3(n8070), .ZN(P1_U3256) );
  XNOR2_X1 U9217 ( .A(n8073), .B(n8081), .ZN(n8074) );
  NAND2_X1 U9218 ( .A1(n8074), .A2(n10794), .ZN(n8078) );
  OAI22_X1 U9219 ( .A1(n8767), .A2(n9559), .B1(n8075), .B2(n9561), .ZN(n8076)
         );
  INV_X1 U9220 ( .A(n8076), .ZN(n8077) );
  NAND2_X1 U9221 ( .A1(n8078), .A2(n8077), .ZN(n10924) );
  INV_X1 U9222 ( .A(n10924), .ZN(n8091) );
  NAND2_X1 U9223 ( .A1(n10901), .A2(n9274), .ZN(n8079) );
  OAI21_X1 U9224 ( .B1(n5125), .B2(n8082), .A(n8100), .ZN(n10925) );
  INV_X1 U9225 ( .A(n8095), .ZN(n10920) );
  NOR2_X1 U9226 ( .A1(n8083), .A2(n10920), .ZN(n8084) );
  OR2_X1 U9227 ( .A1(n8101), .A2(n8084), .ZN(n10922) );
  INV_X1 U9228 ( .A(n8085), .ZN(n8086) );
  OAI22_X1 U9229 ( .A1(n10803), .A2(n7797), .B1(n8086), .B2(n9549), .ZN(n8087)
         );
  AOI21_X1 U9230 ( .B1(n9573), .B2(n8095), .A(n8087), .ZN(n8088) );
  OAI21_X1 U9231 ( .B1(n10922), .B2(n9363), .A(n8088), .ZN(n8089) );
  AOI21_X1 U9232 ( .B1(n10925), .B2(n9572), .A(n8089), .ZN(n8090) );
  OAI21_X1 U9233 ( .B1(n7664), .B2(n8091), .A(n8090), .ZN(P2_U3284) );
  XNOR2_X1 U9234 ( .A(n8092), .B(n8098), .ZN(n8094) );
  OAI22_X1 U9235 ( .A1(n9052), .A2(n9559), .B1(n8559), .B2(n9561), .ZN(n8093)
         );
  AOI21_X1 U9236 ( .B1(n8094), .B2(n10794), .A(n8093), .ZN(n10943) );
  INV_X1 U9237 ( .A(n8559), .ZN(n9273) );
  OR2_X1 U9238 ( .A1(n8095), .A2(n9273), .ZN(n8097) );
  AND2_X1 U9239 ( .A1(n8100), .A2(n8097), .ZN(n8096) );
  OR2_X1 U9240 ( .A1(n8096), .A2(n8098), .ZN(n10937) );
  AND2_X1 U9241 ( .A1(n8098), .A2(n8097), .ZN(n8099) );
  NAND3_X1 U9242 ( .A1(n10937), .A2(n9572), .A3(n8357), .ZN(n8106) );
  OR2_X1 U9243 ( .A1(n8101), .A2(n8358), .ZN(n8102) );
  AND2_X1 U9244 ( .A1(n8102), .A2(n8429), .ZN(n10941) );
  AOI22_X1 U9245 ( .A1(n7664), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8564), .B2(
        n10798), .ZN(n8103) );
  OAI21_X1 U9246 ( .B1(n8358), .B2(n9547), .A(n8103), .ZN(n8104) );
  AOI21_X1 U9247 ( .B1(n10941), .B2(n9568), .A(n8104), .ZN(n8105) );
  OAI211_X1 U9248 ( .C1(n7664), .C2(n10943), .A(n8106), .B(n8105), .ZN(
        P2_U3283) );
  NAND2_X1 U9249 ( .A1(n8108), .A2(n8107), .ZN(n8109) );
  NAND2_X1 U9250 ( .A1(n10872), .A2(n8795), .ZN(n8112) );
  NAND2_X1 U9251 ( .A1(n9821), .A2(n8676), .ZN(n8111) );
  NAND2_X1 U9252 ( .A1(n8112), .A2(n8111), .ZN(n8113) );
  XNOR2_X1 U9253 ( .A(n8113), .B(n8724), .ZN(n8114) );
  NAND2_X1 U9254 ( .A1(n8115), .A2(n8114), .ZN(n8158) );
  NAND2_X1 U9255 ( .A1(n8157), .A2(n8158), .ZN(n8117) );
  AND2_X1 U9256 ( .A1(n9821), .A2(n8790), .ZN(n8116) );
  AOI21_X1 U9257 ( .B1(n10872), .B2(n8676), .A(n8116), .ZN(n8156) );
  XNOR2_X1 U9258 ( .A(n8117), .B(n8156), .ZN(n8125) );
  NAND2_X1 U9259 ( .A1(n9804), .A2(n8118), .ZN(n8122) );
  NAND2_X1 U9260 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10673) );
  INV_X1 U9261 ( .A(n10673), .ZN(n8119) );
  AOI21_X1 U9262 ( .B1(n9805), .B2(n8120), .A(n8119), .ZN(n8121) );
  OAI211_X1 U9263 ( .C1(n8147), .C2(n9808), .A(n8122), .B(n8121), .ZN(n8123)
         );
  AOI21_X1 U9264 ( .B1(n10872), .B2(n9811), .A(n8123), .ZN(n8124) );
  OAI21_X1 U9265 ( .B1(n8125), .B2(n9813), .A(n8124), .ZN(P1_U3215) );
  INV_X1 U9266 ( .A(n6957), .ZN(n8126) );
  INV_X1 U9267 ( .A(n8662), .ZN(n8173) );
  INV_X1 U9268 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8663) );
  OAI222_X1 U9269 ( .A1(n8126), .A2(P1_U3084), .B1(n5044), .B2(n8173), .C1(
        n8663), .C2(n8399), .ZN(P1_U3332) );
  NAND2_X1 U9270 ( .A1(n8127), .A2(n8749), .ZN(n8130) );
  AOI22_X1 U9271 ( .A1(n8638), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n8637), .B2(
        n8128), .ZN(n8129) );
  INV_X1 U9272 ( .A(n8284), .ZN(n8295) );
  NAND2_X1 U9273 ( .A1(n8231), .A2(n8295), .ZN(n8913) );
  OR2_X1 U9274 ( .A1(n8170), .A2(n9820), .ZN(n8132) );
  INV_X1 U9275 ( .A(n8233), .ZN(n8136) );
  AOI21_X1 U9276 ( .B1(n9004), .B2(n8134), .A(n8136), .ZN(n10916) );
  INV_X1 U9277 ( .A(n10916), .ZN(n10913) );
  NAND2_X1 U9278 ( .A1(n8138), .A2(n8906), .ZN(n8139) );
  AOI21_X1 U9279 ( .B1(n8139), .B2(n8135), .A(n9131), .ZN(n8149) );
  INV_X1 U9280 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8140) );
  NAND2_X1 U9281 ( .A1(n8141), .A2(n8140), .ZN(n8142) );
  AND2_X1 U9282 ( .A1(n8247), .A2(n8142), .ZN(n8303) );
  NAND2_X1 U9283 ( .A1(n7099), .A2(n8303), .ZN(n8146) );
  NAND2_X1 U9284 ( .A1(n5052), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8145) );
  NAND2_X1 U9285 ( .A1(n5051), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8144) );
  NAND2_X1 U9286 ( .A1(n5038), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8143) );
  NAND4_X1 U9287 ( .A1(n8146), .A2(n8145), .A3(n8144), .A4(n8143), .ZN(n9819)
         );
  INV_X1 U9288 ( .A(n9819), .ZN(n8238) );
  OAI22_X1 U9289 ( .A1(n8147), .A2(n10013), .B1(n8238), .B2(n10015), .ZN(n8148) );
  AOI21_X1 U9290 ( .B1(n8149), .B2(n8253), .A(n8148), .ZN(n10911) );
  INV_X1 U9291 ( .A(n10911), .ZN(n8154) );
  INV_X1 U9292 ( .A(n8231), .ZN(n10912) );
  OAI211_X1 U9293 ( .C1(n8150), .C2(n10912), .A(n10981), .B(n8300), .ZN(n10910) );
  INV_X1 U9294 ( .A(n10999), .ZN(n8268) );
  AOI22_X1 U9295 ( .A1(n11006), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8223), .B2(
        n10994), .ZN(n8152) );
  NAND2_X1 U9296 ( .A1(n8231), .A2(n10996), .ZN(n8151) );
  OAI211_X1 U9297 ( .C1(n10910), .C2(n8268), .A(n8152), .B(n8151), .ZN(n8153)
         );
  AOI21_X1 U9298 ( .B1(n8154), .B2(n10022), .A(n8153), .ZN(n8155) );
  OAI21_X1 U9299 ( .B1(n10913), .B2(n10070), .A(n8155), .ZN(P1_U3279) );
  NAND2_X1 U9300 ( .A1(n8157), .A2(n8156), .ZN(n8159) );
  NAND2_X1 U9301 ( .A1(n8170), .A2(n8795), .ZN(n8161) );
  NAND2_X1 U9302 ( .A1(n9820), .A2(n8676), .ZN(n8160) );
  NAND2_X1 U9303 ( .A1(n8161), .A2(n8160), .ZN(n8162) );
  XNOR2_X1 U9304 ( .A(n8162), .B(n8724), .ZN(n8221) );
  AND2_X1 U9305 ( .A1(n9820), .A2(n8790), .ZN(n8163) );
  AOI21_X1 U9306 ( .B1(n8170), .B2(n8676), .A(n8163), .ZN(n8220) );
  XNOR2_X1 U9307 ( .A(n8221), .B(n8220), .ZN(n8164) );
  NAND2_X1 U9308 ( .A1(n9804), .A2(n8165), .ZN(n8168) );
  AOI21_X1 U9309 ( .B1(n9805), .B2(n9821), .A(n8166), .ZN(n8167) );
  OAI211_X1 U9310 ( .C1(n8295), .C2(n9808), .A(n8168), .B(n8167), .ZN(n8169)
         );
  AOI21_X1 U9311 ( .B1(n8170), .B2(n9811), .A(n8169), .ZN(n8171) );
  OAI21_X1 U9312 ( .B1(n8172), .B2(n9813), .A(n8171), .ZN(P1_U3234) );
  OAI222_X1 U9313 ( .A1(n9698), .A2(n8175), .B1(P2_U3152), .B2(n8174), .C1(
        n5043), .C2(n8173), .ZN(P2_U3337) );
  AOI211_X1 U9314 ( .C1(n8178), .C2(n8177), .A(n9890), .B(n8176), .ZN(n8186)
         );
  AOI211_X1 U9315 ( .C1(n8181), .C2(n8180), .A(n10684), .B(n8179), .ZN(n8185)
         );
  NAND2_X1 U9316 ( .A1(n10679), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n8182) );
  NAND2_X1 U9317 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8537) );
  OAI211_X1 U9318 ( .C1(n10677), .C2(n8183), .A(n8182), .B(n8537), .ZN(n8184)
         );
  OR3_X1 U9319 ( .A1(n8186), .A2(n8185), .A3(n8184), .ZN(P1_U3257) );
  INV_X1 U9320 ( .A(n8187), .ZN(n8426) );
  OAI22_X1 U9321 ( .A1(n9066), .A2(n9559), .B1(n8422), .B2(n9561), .ZN(n8418)
         );
  AOI22_X1 U9322 ( .A1(n9257), .A2(n8418), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3152), .ZN(n8188) );
  OAI21_X1 U9323 ( .B1(n9259), .B2(n8426), .A(n8188), .ZN(n8189) );
  AOI21_X1 U9324 ( .B1(n9655), .B2(n9261), .A(n8189), .ZN(n8196) );
  INV_X1 U9325 ( .A(n8191), .ZN(n8194) );
  OAI22_X1 U9326 ( .A1(n8192), .A2(n5042), .B1(n8422), .B2(n9240), .ZN(n8193)
         );
  NAND3_X1 U9327 ( .A1(n9059), .A2(n8194), .A3(n8193), .ZN(n8195) );
  OAI211_X1 U9328 ( .C1(n8197), .C2(n5042), .A(n8196), .B(n8195), .ZN(P2_U3228) );
  OAI21_X1 U9329 ( .B1(n8199), .B2(P2_REG2_REG_14__SCAN_IN), .A(n8198), .ZN(
        n9294) );
  XNOR2_X1 U9330 ( .A(n9294), .B(n9302), .ZN(n8201) );
  INV_X1 U9331 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8200) );
  OAI21_X1 U9332 ( .B1(n8201), .B2(n8200), .A(n9296), .ZN(n8202) );
  INV_X1 U9333 ( .A(n8202), .ZN(n8211) );
  NAND2_X1 U9334 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n9048) );
  INV_X1 U9335 ( .A(n9048), .ZN(n8204) );
  NOR2_X1 U9336 ( .A1(n10710), .A2(n9295), .ZN(n8203) );
  AOI211_X1 U9337 ( .C1(n10718), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n8204), .B(
        n8203), .ZN(n8210) );
  AOI21_X1 U9338 ( .B1(n8207), .B2(n8206), .A(n8205), .ZN(n9301) );
  XNOR2_X1 U9339 ( .A(n9301), .B(n9295), .ZN(n8208) );
  NAND2_X1 U9340 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8208), .ZN(n9303) );
  OAI211_X1 U9341 ( .C1(n8208), .C2(P2_REG1_REG_15__SCAN_IN), .A(n10726), .B(
        n9303), .ZN(n8209) );
  OAI211_X1 U9342 ( .C1(n8211), .C2(n10719), .A(n8210), .B(n8209), .ZN(
        P2_U3260) );
  NAND2_X1 U9343 ( .A1(n8231), .A2(n8795), .ZN(n8213) );
  NAND2_X1 U9344 ( .A1(n8284), .A2(n8676), .ZN(n8212) );
  NAND2_X1 U9345 ( .A1(n8213), .A2(n8212), .ZN(n8214) );
  XNOR2_X1 U9346 ( .A(n8214), .B(n8724), .ZN(n8219) );
  INV_X1 U9347 ( .A(n8219), .ZN(n8217) );
  AND2_X1 U9348 ( .A1(n8284), .A2(n8790), .ZN(n8215) );
  AOI21_X1 U9349 ( .B1(n8231), .B2(n8676), .A(n8215), .ZN(n8218) );
  INV_X1 U9350 ( .A(n8218), .ZN(n8216) );
  NAND2_X1 U9351 ( .A1(n8217), .A2(n8216), .ZN(n8274) );
  NAND2_X1 U9352 ( .A1(n8219), .A2(n8218), .ZN(n8272) );
  NAND2_X1 U9353 ( .A1(n8274), .A2(n8272), .ZN(n8222) );
  XOR2_X1 U9354 ( .A(n8222), .B(n8273), .Z(n8230) );
  NAND2_X1 U9355 ( .A1(n9804), .A2(n8223), .ZN(n8227) );
  INV_X1 U9356 ( .A(n8224), .ZN(n8225) );
  AOI21_X1 U9357 ( .B1(n9805), .B2(n9820), .A(n8225), .ZN(n8226) );
  OAI211_X1 U9358 ( .C1(n8238), .C2(n9808), .A(n8227), .B(n8226), .ZN(n8228)
         );
  AOI21_X1 U9359 ( .B1(n8231), .B2(n9811), .A(n8228), .ZN(n8229) );
  OAI21_X1 U9360 ( .B1(n8230), .B2(n9813), .A(n8229), .ZN(P1_U3222) );
  NAND2_X1 U9361 ( .A1(n8231), .A2(n8284), .ZN(n8232) );
  INV_X1 U9362 ( .A(n8292), .ZN(n8240) );
  NAND2_X1 U9363 ( .A1(n8234), .A2(n8749), .ZN(n8237) );
  AOI22_X1 U9364 ( .A1(n8638), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n8637), .B2(
        n8235), .ZN(n8236) );
  OR2_X1 U9365 ( .A1(n10928), .A2(n8238), .ZN(n8915) );
  NAND2_X1 U9366 ( .A1(n10928), .A2(n8238), .ZN(n8917) );
  OR2_X1 U9367 ( .A1(n10928), .A2(n9819), .ZN(n8241) );
  NAND2_X1 U9368 ( .A1(n8242), .A2(n8749), .ZN(n8245) );
  AOI22_X1 U9369 ( .A1(n8638), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n8637), .B2(
        n8243), .ZN(n8244) );
  NAND2_X1 U9370 ( .A1(n7351), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8252) );
  NAND2_X1 U9371 ( .A1(n8247), .A2(n8246), .ZN(n8248) );
  AND2_X1 U9372 ( .A1(n8257), .A2(n8248), .ZN(n8493) );
  NAND2_X1 U9373 ( .A1(n7099), .A2(n8493), .ZN(n8251) );
  NAND2_X1 U9374 ( .A1(n5051), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n8250) );
  NAND2_X1 U9375 ( .A1(n5038), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8249) );
  NAND4_X1 U9376 ( .A1(n8252), .A2(n8251), .A3(n8250), .A4(n8249), .ZN(n9818)
         );
  INV_X1 U9377 ( .A(n9818), .ZN(n8390) );
  NAND2_X1 U9378 ( .A1(n8511), .A2(n8390), .ZN(n8921) );
  NAND2_X1 U9379 ( .A1(n8922), .A2(n8921), .ZN(n9007) );
  XNOR2_X1 U9380 ( .A(n8377), .B(n9007), .ZN(n10955) );
  INV_X1 U9381 ( .A(n10955), .ZN(n8271) );
  OAI211_X1 U9382 ( .C1(n8254), .C2(n5572), .A(n8388), .B(n10980), .ZN(n8264)
         );
  NAND2_X1 U9383 ( .A1(n5052), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n8262) );
  INV_X1 U9384 ( .A(n8255), .ZN(n8381) );
  NAND2_X1 U9385 ( .A1(n8257), .A2(n8256), .ZN(n8258) );
  AND2_X1 U9386 ( .A1(n8381), .A2(n8258), .ZN(n8547) );
  NAND2_X1 U9387 ( .A1(n7099), .A2(n8547), .ZN(n8261) );
  NAND2_X1 U9388 ( .A1(n5051), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8260) );
  NAND2_X1 U9389 ( .A1(n5038), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n8259) );
  NAND4_X1 U9390 ( .A1(n8262), .A2(n8261), .A3(n8260), .A4(n8259), .ZN(n10976)
         );
  AOI22_X1 U9391 ( .A1(n10975), .A2(n9819), .B1(n10976), .B2(n10977), .ZN(
        n8263) );
  NAND2_X1 U9392 ( .A1(n8264), .A2(n8263), .ZN(n10954) );
  INV_X1 U9393 ( .A(n8302), .ZN(n8265) );
  INV_X1 U9394 ( .A(n8511), .ZN(n10952) );
  OAI211_X1 U9395 ( .C1(n8265), .C2(n10952), .A(n10981), .B(n8391), .ZN(n10951) );
  AOI22_X1 U9396 ( .A1(n10738), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8493), .B2(
        n10994), .ZN(n8267) );
  NAND2_X1 U9397 ( .A1(n8511), .A2(n10996), .ZN(n8266) );
  OAI211_X1 U9398 ( .C1(n10951), .C2(n8268), .A(n8267), .B(n8266), .ZN(n8269)
         );
  AOI21_X1 U9399 ( .B1(n10954), .B2(n10022), .A(n8269), .ZN(n8270) );
  OAI21_X1 U9400 ( .B1(n8271), .B2(n10070), .A(n8270), .ZN(P1_U3277) );
  NAND2_X1 U9401 ( .A1(n10928), .A2(n8676), .ZN(n8277) );
  NAND2_X1 U9402 ( .A1(n9819), .A2(n8790), .ZN(n8276) );
  NAND2_X1 U9403 ( .A1(n8277), .A2(n8276), .ZN(n8497) );
  NAND2_X1 U9404 ( .A1(n10928), .A2(n8795), .ZN(n8279) );
  NAND2_X1 U9405 ( .A1(n9819), .A2(n8676), .ZN(n8278) );
  NAND2_X1 U9406 ( .A1(n8279), .A2(n8278), .ZN(n8280) );
  XNOR2_X1 U9407 ( .A(n8280), .B(n8793), .ZN(n8498) );
  XOR2_X1 U9408 ( .A(n8497), .B(n8498), .Z(n8281) );
  XNOR2_X1 U9409 ( .A(n8499), .B(n8281), .ZN(n8289) );
  NAND2_X1 U9410 ( .A1(n9804), .A2(n8303), .ZN(n8286) );
  INV_X1 U9411 ( .A(n8282), .ZN(n8283) );
  AOI21_X1 U9412 ( .B1(n9805), .B2(n8284), .A(n8283), .ZN(n8285) );
  OAI211_X1 U9413 ( .C1(n8390), .C2(n9808), .A(n8286), .B(n8285), .ZN(n8287)
         );
  AOI21_X1 U9414 ( .B1(n10928), .B2(n9811), .A(n8287), .ZN(n8288) );
  OAI21_X1 U9415 ( .B1(n8289), .B2(n9813), .A(n8288), .ZN(P1_U3232) );
  INV_X1 U9416 ( .A(n8679), .ZN(n8370) );
  OAI222_X1 U9417 ( .A1(P1_U3084), .A2(n5509), .B1(n5044), .B2(n8370), .C1(
        n10266), .C2(n8399), .ZN(P1_U3331) );
  INV_X1 U9418 ( .A(n8290), .ZN(n8291) );
  AOI21_X1 U9419 ( .B1(n8991), .B2(n8292), .A(n8291), .ZN(n8299) );
  OAI21_X1 U9420 ( .B1(n8991), .B2(n8294), .A(n8293), .ZN(n8297) );
  OAI22_X1 U9421 ( .A1(n8295), .A2(n10013), .B1(n8390), .B2(n10015), .ZN(n8296) );
  AOI21_X1 U9422 ( .B1(n8297), .B2(n10980), .A(n8296), .ZN(n8298) );
  OAI21_X1 U9423 ( .B1(n8299), .B2(n7169), .A(n8298), .ZN(n10930) );
  INV_X1 U9424 ( .A(n10930), .ZN(n8308) );
  INV_X1 U9425 ( .A(n8299), .ZN(n10932) );
  NAND2_X1 U9426 ( .A1(n8300), .A2(n10928), .ZN(n8301) );
  NAND2_X1 U9427 ( .A1(n8302), .A2(n8301), .ZN(n10929) );
  AOI22_X1 U9428 ( .A1(n10738), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8303), .B2(
        n10994), .ZN(n8305) );
  NAND2_X1 U9429 ( .A1(n10928), .A2(n10996), .ZN(n8304) );
  OAI211_X1 U9430 ( .C1(n10929), .C2(n10733), .A(n8305), .B(n8304), .ZN(n8306)
         );
  AOI21_X1 U9431 ( .B1(n10932), .B2(n9929), .A(n8306), .ZN(n8307) );
  OAI21_X1 U9432 ( .B1(n8308), .B2(n10738), .A(n8307), .ZN(P1_U3278) );
  NOR2_X1 U9433 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n8345) );
  NOR2_X1 U9434 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n8343) );
  NOR2_X1 U9435 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n8341) );
  NOR2_X1 U9436 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n8339) );
  NOR2_X1 U9437 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n8337) );
  NOR2_X1 U9438 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n8334) );
  NAND2_X1 U9439 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n8332) );
  XOR2_X1 U9440 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n10638) );
  NAND2_X1 U9441 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n8330) );
  XOR2_X1 U9442 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n10636) );
  NOR2_X1 U9443 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n8314) );
  XNOR2_X1 U9444 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10627) );
  NAND2_X1 U9445 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n8312) );
  XOR2_X1 U9446 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(P1_ADDR_REG_3__SCAN_IN), .Z(
        n10625) );
  NAND2_X1 U9447 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n8310) );
  XOR2_X1 U9448 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10623) );
  AOI21_X1 U9449 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10617) );
  INV_X1 U9450 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10621) );
  NAND3_X1 U9451 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10619) );
  OAI21_X1 U9452 ( .B1(n10617), .B2(n10621), .A(n10619), .ZN(n10622) );
  NAND2_X1 U9453 ( .A1(n10623), .A2(n10622), .ZN(n8309) );
  NAND2_X1 U9454 ( .A1(n8310), .A2(n8309), .ZN(n10624) );
  NAND2_X1 U9455 ( .A1(n10625), .A2(n10624), .ZN(n8311) );
  NAND2_X1 U9456 ( .A1(n8312), .A2(n8311), .ZN(n10626) );
  NOR2_X1 U9457 ( .A1(n10627), .A2(n10626), .ZN(n8313) );
  NOR2_X1 U9458 ( .A1(n8314), .A2(n8313), .ZN(n8315) );
  NOR2_X1 U9459 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n8315), .ZN(n10629) );
  AND2_X1 U9460 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n8315), .ZN(n10628) );
  NOR2_X1 U9461 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10628), .ZN(n8316) );
  NOR2_X1 U9462 ( .A1(n10629), .A2(n8316), .ZN(n8317) );
  NAND2_X1 U9463 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n8317), .ZN(n8319) );
  XOR2_X1 U9464 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n8317), .Z(n10631) );
  NAND2_X1 U9465 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10631), .ZN(n8318) );
  NAND2_X1 U9466 ( .A1(n8319), .A2(n8318), .ZN(n8320) );
  NAND2_X1 U9467 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n8320), .ZN(n8322) );
  XOR2_X1 U9468 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n8320), .Z(n10632) );
  NAND2_X1 U9469 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10632), .ZN(n8321) );
  NAND2_X1 U9470 ( .A1(n8322), .A2(n8321), .ZN(n8323) );
  NAND2_X1 U9471 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n8323), .ZN(n8325) );
  XOR2_X1 U9472 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n8323), .Z(n10633) );
  NAND2_X1 U9473 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10633), .ZN(n8324) );
  NAND2_X1 U9474 ( .A1(n8325), .A2(n8324), .ZN(n8326) );
  NAND2_X1 U9475 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n8326), .ZN(n8328) );
  XOR2_X1 U9476 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n8326), .Z(n10634) );
  NAND2_X1 U9477 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10634), .ZN(n8327) );
  NAND2_X1 U9478 ( .A1(n8328), .A2(n8327), .ZN(n10635) );
  NAND2_X1 U9479 ( .A1(n10636), .A2(n10635), .ZN(n8329) );
  NAND2_X1 U9480 ( .A1(n8330), .A2(n8329), .ZN(n10637) );
  NAND2_X1 U9481 ( .A1(n10638), .A2(n10637), .ZN(n8331) );
  NAND2_X1 U9482 ( .A1(n8332), .A2(n8331), .ZN(n10640) );
  XNOR2_X1 U9483 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10639) );
  NOR2_X1 U9484 ( .A1(n10640), .A2(n10639), .ZN(n8333) );
  XOR2_X1 U9485 ( .A(n8335), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n10641) );
  NOR2_X1 U9486 ( .A1(n10642), .A2(n10641), .ZN(n8336) );
  NOR2_X1 U9487 ( .A1(n8337), .A2(n8336), .ZN(n10644) );
  XNOR2_X1 U9488 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10643) );
  NOR2_X1 U9489 ( .A1(n10644), .A2(n10643), .ZN(n8338) );
  NOR2_X1 U9490 ( .A1(n8339), .A2(n8338), .ZN(n10646) );
  XNOR2_X1 U9491 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10645) );
  NOR2_X1 U9492 ( .A1(n10646), .A2(n10645), .ZN(n8340) );
  NOR2_X1 U9493 ( .A1(n8341), .A2(n8340), .ZN(n10648) );
  XNOR2_X1 U9494 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10647) );
  NOR2_X1 U9495 ( .A1(n10648), .A2(n10647), .ZN(n8342) );
  NOR2_X1 U9496 ( .A1(n8343), .A2(n8342), .ZN(n10650) );
  XNOR2_X1 U9497 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10649) );
  NOR2_X1 U9498 ( .A1(n10650), .A2(n10649), .ZN(n8344) );
  NOR2_X1 U9499 ( .A1(n8345), .A2(n8344), .ZN(n8346) );
  AND2_X1 U9500 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n8346), .ZN(n10651) );
  NOR2_X1 U9501 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10651), .ZN(n8347) );
  NOR2_X1 U9502 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n8346), .ZN(n10652) );
  NOR2_X1 U9503 ( .A1(n8347), .A2(n10652), .ZN(n8349) );
  XNOR2_X1 U9504 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n8348) );
  XNOR2_X1 U9505 ( .A(n8349), .B(n8348), .ZN(ADD_1071_U4) );
  NAND2_X1 U9506 ( .A1(n8599), .A2(n8350), .ZN(n8352) );
  NOR2_X1 U9507 ( .A1(n8351), .A2(P1_U3084), .ZN(n9041) );
  INV_X1 U9508 ( .A(n9041), .ZN(n9045) );
  OAI211_X1 U9509 ( .C1(n8600), .C2(n10575), .A(n8352), .B(n9045), .ZN(
        P1_U3330) );
  NAND2_X1 U9510 ( .A1(n8599), .A2(n8353), .ZN(n8355) );
  OAI211_X1 U9511 ( .C1(n8356), .C2(n9698), .A(n8355), .B(n8354), .ZN(P2_U3335) );
  AOI21_X1 U9512 ( .B1(n8360), .B2(n8359), .A(n8420), .ZN(n9668) );
  INV_X1 U9513 ( .A(n9664), .ZN(n8421) );
  XNOR2_X1 U9514 ( .A(n8421), .B(n8429), .ZN(n9665) );
  AOI22_X1 U9515 ( .A1(n7664), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8760), .B2(
        n10798), .ZN(n8361) );
  OAI21_X1 U9516 ( .B1(n8421), .B2(n9547), .A(n8361), .ZN(n8368) );
  AOI211_X1 U9517 ( .C1(n8364), .C2(n8363), .A(n9538), .B(n8362), .ZN(n8366)
         );
  OAI22_X1 U9518 ( .A1(n8422), .A2(n9559), .B1(n8767), .B2(n9561), .ZN(n8365)
         );
  NOR2_X1 U9519 ( .A1(n8366), .A2(n8365), .ZN(n9667) );
  NOR2_X1 U9520 ( .A1(n9667), .A2(n7664), .ZN(n8367) );
  AOI211_X1 U9521 ( .C1(n9665), .C2(n9568), .A(n8368), .B(n8367), .ZN(n8369)
         );
  OAI21_X1 U9522 ( .B1(n9668), .B2(n9533), .A(n8369), .ZN(P2_U3282) );
  OAI222_X1 U9523 ( .A1(P2_U3152), .A2(n8371), .B1(n5043), .B2(n8370), .C1(
        n9698), .C2(n6171), .ZN(P2_U3336) );
  NAND2_X1 U9524 ( .A1(n8372), .A2(n8749), .ZN(n8376) );
  INV_X1 U9525 ( .A(n8373), .ZN(n8374) );
  AOI22_X1 U9526 ( .A1(n8638), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8637), .B2(
        n8374), .ZN(n8375) );
  INV_X1 U9527 ( .A(n10976), .ZN(n8496) );
  NAND2_X1 U9528 ( .A1(n8554), .A2(n8496), .ZN(n8925) );
  INV_X1 U9529 ( .A(n8460), .ZN(n8379) );
  AOI21_X1 U9530 ( .B1(n9009), .B2(n8378), .A(n8379), .ZN(n10964) );
  INV_X1 U9531 ( .A(n10964), .ZN(n8398) );
  NAND2_X1 U9532 ( .A1(n5052), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8387) );
  INV_X1 U9533 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8380) );
  NAND2_X1 U9534 ( .A1(n8381), .A2(n8380), .ZN(n8382) );
  AND2_X1 U9535 ( .A1(n8383), .A2(n8382), .ZN(n10995) );
  NAND2_X1 U9536 ( .A1(n7099), .A2(n10995), .ZN(n8386) );
  NAND2_X1 U9537 ( .A1(n5051), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8385) );
  NAND2_X1 U9538 ( .A1(n5039), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8384) );
  NAND4_X1 U9539 ( .A1(n8387), .A2(n8386), .A3(n8385), .A4(n8384), .ZN(n9817)
         );
  INV_X1 U9540 ( .A(n9817), .ZN(n8552) );
  XNOR2_X1 U9541 ( .A(n8471), .B(n9009), .ZN(n8389) );
  OAI222_X1 U9542 ( .A1(n10015), .A2(n8552), .B1(n10013), .B2(n8390), .C1(
        n9131), .C2(n8389), .ZN(n10963) );
  INV_X1 U9543 ( .A(n8554), .ZN(n10959) );
  INV_X1 U9544 ( .A(n8391), .ZN(n8393) );
  INV_X1 U9545 ( .A(n10983), .ZN(n8392) );
  OAI21_X1 U9546 ( .B1(n10959), .B2(n8393), .A(n8392), .ZN(n10961) );
  AOI22_X1 U9547 ( .A1(n10738), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8547), .B2(
        n10994), .ZN(n8395) );
  NAND2_X1 U9548 ( .A1(n8554), .A2(n10996), .ZN(n8394) );
  OAI211_X1 U9549 ( .C1(n10961), .C2(n10733), .A(n8395), .B(n8394), .ZN(n8396)
         );
  AOI21_X1 U9550 ( .B1(n10963), .B2(n10022), .A(n8396), .ZN(n8397) );
  OAI21_X1 U9551 ( .B1(n8398), .B2(n10070), .A(n8397), .ZN(P1_U3276) );
  INV_X1 U9552 ( .A(n8688), .ZN(n8402) );
  INV_X1 U9553 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10264) );
  OAI222_X1 U9554 ( .A1(n8400), .A2(P1_U3084), .B1(n5044), .B2(n8402), .C1(
        n10264), .C2(n8399), .ZN(P1_U3329) );
  OAI222_X1 U9555 ( .A1(P2_U3152), .A2(n8403), .B1(n5043), .B2(n8402), .C1(
        n8401), .C2(n9698), .ZN(P2_U3334) );
  INV_X1 U9556 ( .A(n8404), .ZN(n8405) );
  AOI21_X1 U9557 ( .B1(n8406), .B2(n8405), .A(n5042), .ZN(n8410) );
  NOR3_X1 U9558 ( .A1(n8407), .A2(n9066), .A3(n9240), .ZN(n8409) );
  OAI21_X1 U9559 ( .B1(n8410), .B2(n8409), .A(n8408), .ZN(n8415) );
  NOR2_X1 U9560 ( .A1(n8411), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9335) );
  INV_X1 U9561 ( .A(n9522), .ZN(n8412) );
  OAI22_X1 U9562 ( .A1(n9230), .A2(n9066), .B1(n9259), .B2(n8412), .ZN(n8413)
         );
  AOI211_X1 U9563 ( .C1(n9244), .C2(n9528), .A(n9335), .B(n8413), .ZN(n8414)
         );
  OAI211_X1 U9564 ( .C1(n9524), .C2(n9099), .A(n8415), .B(n8414), .ZN(P2_U3240) );
  INV_X1 U9565 ( .A(n8445), .ZN(n8440) );
  OAI21_X1 U9566 ( .B1(n5110), .B2(n8440), .A(n8416), .ZN(n8417) );
  XOR2_X1 U9567 ( .A(n8424), .B(n8417), .Z(n8419) );
  AOI21_X1 U9568 ( .B1(n8419), .B2(n10794), .A(n8418), .ZN(n9657) );
  INV_X1 U9569 ( .A(n8422), .ZN(n9270) );
  AOI21_X1 U9570 ( .B1(n8424), .B2(n8423), .A(n9065), .ZN(n8425) );
  INV_X1 U9571 ( .A(n8425), .ZN(n9658) );
  INV_X1 U9572 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8427) );
  OAI22_X1 U9573 ( .A1(n10803), .A2(n8427), .B1(n8426), .B2(n9549), .ZN(n8428)
         );
  AOI21_X1 U9574 ( .B1(n9655), .B2(n9573), .A(n8428), .ZN(n8433) );
  INV_X1 U9575 ( .A(n9655), .ZN(n8430) );
  OAI21_X1 U9576 ( .B1(n8430), .B2(n5113), .A(n10940), .ZN(n8431) );
  NOR2_X1 U9577 ( .A1(n8431), .A2(n9534), .ZN(n9654) );
  NAND2_X1 U9578 ( .A1(n9654), .A2(n9426), .ZN(n8432) );
  OAI211_X1 U9579 ( .C1(n9658), .C2(n9533), .A(n8433), .B(n8432), .ZN(n8434)
         );
  INV_X1 U9580 ( .A(n8434), .ZN(n8435) );
  OAI21_X1 U9581 ( .B1(n7664), .B2(n9657), .A(n8435), .ZN(P2_U3280) );
  INV_X1 U9582 ( .A(n8586), .ZN(n8438) );
  OAI222_X1 U9583 ( .A1(P1_U3084), .A2(n8436), .B1(n5044), .B2(n8438), .C1(
        n10260), .C2(n10575), .ZN(P1_U3328) );
  OAI222_X1 U9584 ( .A1(n9698), .A2(n8439), .B1(n5043), .B2(n8438), .C1(
        P2_U3152), .C2(n8437), .ZN(P2_U3333) );
  XNOR2_X1 U9585 ( .A(n8441), .B(n8440), .ZN(n9663) );
  AOI21_X1 U9586 ( .B1(n9659), .B2(n8442), .A(n5113), .ZN(n9660) );
  INV_X1 U9587 ( .A(n8443), .ZN(n9047) );
  AOI22_X1 U9588 ( .A1(n7664), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n9047), .B2(
        n10798), .ZN(n8444) );
  OAI21_X1 U9589 ( .B1(n5304), .B2(n9547), .A(n8444), .ZN(n8448) );
  XNOR2_X1 U9590 ( .A(n5110), .B(n8445), .ZN(n8446) );
  INV_X1 U9591 ( .A(n9540), .ZN(n9269) );
  INV_X1 U9592 ( .A(n9052), .ZN(n9271) );
  AOI222_X1 U9593 ( .A1(n10794), .A2(n8446), .B1(n9269), .B2(n10791), .C1(
        n9271), .C2(n10789), .ZN(n9662) );
  NOR2_X1 U9594 ( .A1(n9662), .A2(n7664), .ZN(n8447) );
  AOI211_X1 U9595 ( .C1(n9660), .C2(n9568), .A(n8448), .B(n8447), .ZN(n8449)
         );
  OAI21_X1 U9596 ( .B1(n9663), .B2(n9533), .A(n8449), .ZN(P2_U3281) );
  INV_X1 U9597 ( .A(n8450), .ZN(n8452) );
  NOR2_X1 U9598 ( .A1(n8452), .A2(n8451), .ZN(n8453) );
  XNOR2_X1 U9599 ( .A(n8454), .B(n8453), .ZN(n8458) );
  NAND2_X1 U9600 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9353) );
  OAI21_X1 U9601 ( .B1(n9230), .B2(n9539), .A(n9353), .ZN(n8456) );
  OAI22_X1 U9602 ( .A1(n9229), .A2(n9510), .B1(n9259), .B2(n9512), .ZN(n8455)
         );
  AOI211_X1 U9603 ( .C1(n9641), .C2(n9261), .A(n8456), .B(n8455), .ZN(n8457)
         );
  OAI21_X1 U9604 ( .B1(n8458), .B2(n5042), .A(n8457), .ZN(P2_U3221) );
  NAND2_X1 U9605 ( .A1(n8554), .A2(n10976), .ZN(n8459) );
  NAND2_X1 U9606 ( .A1(n8460), .A2(n8459), .ZN(n10970) );
  NAND2_X1 U9607 ( .A1(n8461), .A2(n8749), .ZN(n8464) );
  AOI22_X1 U9608 ( .A1(n8638), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8637), .B2(
        n8462), .ZN(n8463) );
  OR2_X1 U9609 ( .A1(n10997), .A2(n8552), .ZN(n8929) );
  NAND2_X1 U9610 ( .A1(n10997), .A2(n8552), .ZN(n8930) );
  NAND2_X1 U9611 ( .A1(n8929), .A2(n8930), .ZN(n10969) );
  NAND2_X1 U9612 ( .A1(n10997), .A2(n9817), .ZN(n8465) );
  NAND2_X1 U9613 ( .A1(n8466), .A2(n8749), .ZN(n8468) );
  AOI22_X1 U9614 ( .A1(n8638), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8637), .B2(
        n9868), .ZN(n8467) );
  INV_X1 U9615 ( .A(n10978), .ZN(n9793) );
  NAND2_X1 U9616 ( .A1(n10541), .A2(n9793), .ZN(n10057) );
  INV_X1 U9617 ( .A(n10054), .ZN(n8931) );
  OAI21_X1 U9618 ( .B1(n8469), .B2(n8931), .A(n9106), .ZN(n10540) );
  INV_X1 U9619 ( .A(n8926), .ZN(n8470) );
  INV_X1 U9620 ( .A(n10969), .ZN(n10974) );
  XNOR2_X1 U9621 ( .A(n10058), .B(n10054), .ZN(n8479) );
  NAND2_X1 U9622 ( .A1(n8472), .A2(n9792), .ZN(n8473) );
  NAND2_X1 U9623 ( .A1(n8615), .A2(n8473), .ZN(n10049) );
  INV_X1 U9624 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8474) );
  OAI22_X1 U9625 ( .A1(n10049), .A2(n8618), .B1(n6947), .B2(n8474), .ZN(n8477)
         );
  INV_X1 U9626 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9861) );
  INV_X1 U9627 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n8475) );
  OAI22_X1 U9628 ( .A1(n6948), .A2(n9861), .B1(n5037), .B2(n8475), .ZN(n8476)
         );
  OR2_X1 U9629 ( .A1(n8477), .A2(n8476), .ZN(n10041) );
  AOI22_X1 U9630 ( .A1(n10977), .A2(n10041), .B1(n9817), .B2(n10975), .ZN(
        n8478) );
  OAI21_X1 U9631 ( .B1(n8479), .B2(n9131), .A(n8478), .ZN(n8480) );
  AOI21_X1 U9632 ( .B1(n10540), .B2(n10879), .A(n8480), .ZN(n10544) );
  INV_X1 U9633 ( .A(n10541), .ZN(n9754) );
  INV_X1 U9634 ( .A(n10997), .ZN(n10985) );
  NAND2_X1 U9635 ( .A1(n10983), .A2(n10985), .ZN(n10982) );
  INV_X1 U9636 ( .A(n10048), .ZN(n8481) );
  AOI21_X1 U9637 ( .B1(n10541), .B2(n10982), .A(n8481), .ZN(n10542) );
  NAND2_X1 U9638 ( .A1(n10542), .A2(n10068), .ZN(n8483) );
  AOI22_X1 U9639 ( .A1(n10738), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9751), .B2(
        n10994), .ZN(n8482) );
  OAI211_X1 U9640 ( .C1(n9754), .C2(n10734), .A(n8483), .B(n8482), .ZN(n8484)
         );
  AOI21_X1 U9641 ( .B1(n10540), .B2(n9929), .A(n8484), .ZN(n8485) );
  OAI21_X1 U9642 ( .B1(n10544), .B2(n10738), .A(n8485), .ZN(P1_U3274) );
  XNOR2_X1 U9643 ( .A(n8487), .B(n8486), .ZN(n8492) );
  OAI22_X1 U9644 ( .A1(n9229), .A2(n9266), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10228), .ZN(n8490) );
  INV_X1 U9645 ( .A(n8488), .ZN(n9493) );
  OAI22_X1 U9646 ( .A1(n9230), .A2(n9068), .B1(n9259), .B2(n9493), .ZN(n8489)
         );
  AOI211_X1 U9647 ( .C1(n9634), .C2(n9248), .A(n8490), .B(n8489), .ZN(n8491)
         );
  OAI21_X1 U9648 ( .B1(n8492), .B2(n5042), .A(n8491), .ZN(P2_U3235) );
  NAND2_X1 U9649 ( .A1(n9804), .A2(n8493), .ZN(n8495) );
  AOI22_X1 U9650 ( .A1(n9805), .A2(n9819), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3084), .ZN(n8494) );
  OAI211_X1 U9651 ( .C1(n8496), .C2(n9808), .A(n8495), .B(n8494), .ZN(n8510)
         );
  NAND2_X1 U9652 ( .A1(n8511), .A2(n8795), .ZN(n8501) );
  NAND2_X1 U9653 ( .A1(n9818), .A2(n8676), .ZN(n8500) );
  NAND2_X1 U9654 ( .A1(n8501), .A2(n8500), .ZN(n8502) );
  XNOR2_X1 U9655 ( .A(n8502), .B(n8793), .ZN(n8516) );
  XOR2_X1 U9656 ( .A(n8517), .B(n8516), .Z(n8505) );
  NAND2_X1 U9657 ( .A1(n8511), .A2(n8676), .ZN(n8504) );
  NAND2_X1 U9658 ( .A1(n9818), .A2(n8790), .ZN(n8503) );
  NAND2_X1 U9659 ( .A1(n8504), .A2(n8503), .ZN(n8506) );
  OAI21_X1 U9660 ( .B1(n8505), .B2(n8506), .A(n8530), .ZN(n8508) );
  NAND3_X1 U9661 ( .A1(n8517), .A2(n8516), .A3(n8506), .ZN(n8507) );
  AOI21_X1 U9662 ( .B1(n8508), .B2(n8507), .A(n9813), .ZN(n8509) );
  AOI211_X1 U9663 ( .C1(n8511), .C2(n9811), .A(n8510), .B(n8509), .ZN(n8512)
         );
  INV_X1 U9664 ( .A(n8512), .ZN(P1_U3213) );
  NAND2_X1 U9665 ( .A1(n8554), .A2(n8795), .ZN(n8514) );
  NAND2_X1 U9666 ( .A1(n10976), .A2(n8676), .ZN(n8513) );
  NAND2_X1 U9667 ( .A1(n8514), .A2(n8513), .ZN(n8515) );
  XNOR2_X1 U9668 ( .A(n8515), .B(n8724), .ZN(n8531) );
  NAND3_X1 U9669 ( .A1(n8530), .A2(n8531), .A3(n8529), .ZN(n8543) );
  NAND2_X1 U9670 ( .A1(n8554), .A2(n8676), .ZN(n8519) );
  NAND2_X1 U9671 ( .A1(n10976), .A2(n8790), .ZN(n8518) );
  NAND2_X1 U9672 ( .A1(n8519), .A2(n8518), .ZN(n8546) );
  NAND2_X1 U9673 ( .A1(n10997), .A2(n8795), .ZN(n8521) );
  NAND2_X1 U9674 ( .A1(n9817), .A2(n8676), .ZN(n8520) );
  NAND2_X1 U9675 ( .A1(n8521), .A2(n8520), .ZN(n8522) );
  XNOR2_X1 U9676 ( .A(n8522), .B(n8724), .ZN(n8524) );
  AND2_X1 U9677 ( .A1(n9817), .A2(n8790), .ZN(n8523) );
  AOI21_X1 U9678 ( .B1(n10997), .B2(n8676), .A(n8523), .ZN(n8525) );
  NAND2_X1 U9679 ( .A1(n8524), .A2(n8525), .ZN(n9742) );
  INV_X1 U9680 ( .A(n8524), .ZN(n8527) );
  INV_X1 U9681 ( .A(n8525), .ZN(n8526) );
  NAND2_X1 U9682 ( .A1(n8527), .A2(n8526), .ZN(n8528) );
  AND2_X1 U9683 ( .A1(n9742), .A2(n8528), .ZN(n8535) );
  INV_X1 U9684 ( .A(n8531), .ZN(n8532) );
  AOI21_X1 U9685 ( .B1(n8534), .B2(n8544), .A(n8535), .ZN(n8536) );
  OAI21_X1 U9686 ( .B1(n5111), .B2(n8536), .A(n9744), .ZN(n8542) );
  INV_X1 U9687 ( .A(n8537), .ZN(n8538) );
  AOI21_X1 U9688 ( .B1(n9805), .B2(n10976), .A(n8538), .ZN(n8539) );
  OAI21_X1 U9689 ( .B1(n9793), .B2(n9808), .A(n8539), .ZN(n8540) );
  AOI21_X1 U9690 ( .B1(n9804), .B2(n10995), .A(n8540), .ZN(n8541) );
  OAI211_X1 U9691 ( .C1(n10985), .C2(n9801), .A(n8542), .B(n8541), .ZN(
        P1_U3224) );
  NAND2_X1 U9692 ( .A1(n8544), .A2(n8543), .ZN(n8545) );
  XOR2_X1 U9693 ( .A(n8546), .B(n8545), .Z(n8556) );
  NAND2_X1 U9694 ( .A1(n9804), .A2(n8547), .ZN(n8551) );
  INV_X1 U9695 ( .A(n8548), .ZN(n8549) );
  AOI21_X1 U9696 ( .B1(n9805), .B2(n9818), .A(n8549), .ZN(n8550) );
  OAI211_X1 U9697 ( .C1(n8552), .C2(n9808), .A(n8551), .B(n8550), .ZN(n8553)
         );
  AOI21_X1 U9698 ( .B1(n8554), .B2(n9811), .A(n8553), .ZN(n8555) );
  OAI21_X1 U9699 ( .B1(n8556), .B2(n9813), .A(n8555), .ZN(P1_U3239) );
  OAI22_X1 U9700 ( .A1(n9240), .A2(n8559), .B1(n8558), .B2(n5042), .ZN(n8560)
         );
  NAND3_X1 U9701 ( .A1(n8561), .A2(n5475), .A3(n8560), .ZN(n8568) );
  INV_X1 U9702 ( .A(n8562), .ZN(n8563) );
  AOI21_X1 U9703 ( .B1(n9247), .B2(n9273), .A(n8563), .ZN(n8567) );
  AOI22_X1 U9704 ( .A1(n9244), .A2(n9271), .B1(n9246), .B2(n8564), .ZN(n8566)
         );
  NAND2_X1 U9705 ( .A1(n10938), .A2(n9261), .ZN(n8565) );
  AND4_X1 U9706 ( .A1(n8568), .A2(n8567), .A3(n8566), .A4(n8565), .ZN(n8569)
         );
  OAI21_X1 U9707 ( .B1(n8771), .B2(n5042), .A(n8569), .ZN(P2_U3236) );
  XNOR2_X1 U9708 ( .A(n8570), .B(n8571), .ZN(n8572) );
  XNOR2_X1 U9709 ( .A(n8573), .B(n8572), .ZN(n8577) );
  AOI22_X1 U9710 ( .A1(n9798), .A2(n9828), .B1(n9805), .B2(n9831), .ZN(n8576)
         );
  AOI22_X1 U9711 ( .A1(n9811), .A2(n8582), .B1(n8574), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n8575) );
  OAI211_X1 U9712 ( .C1(n8577), .C2(n9813), .A(n8576), .B(n8575), .ZN(P1_U3220) );
  INV_X1 U9713 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10675) );
  OAI22_X1 U9714 ( .A1(n8578), .A2(n10021), .B1(n10675), .B2(n10741), .ZN(
        n8579) );
  NOR2_X1 U9715 ( .A1(n8580), .A2(n8579), .ZN(n8581) );
  MUX2_X1 U9716 ( .A(n6729), .B(n8581), .S(n10022), .Z(n8585) );
  AOI22_X1 U9717 ( .A1(n8583), .A2(n9929), .B1(n10996), .B2(n8582), .ZN(n8584)
         );
  NAND2_X1 U9718 ( .A1(n8585), .A2(n8584), .ZN(P1_U3290) );
  NAND2_X1 U9719 ( .A1(n8586), .A2(n8749), .ZN(n8588) );
  OR2_X1 U9720 ( .A1(n7183), .A2(n10260), .ZN(n8587) );
  NAND2_X1 U9721 ( .A1(n10099), .A2(n8795), .ZN(n8596) );
  NAND2_X1 U9722 ( .A1(n5052), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8594) );
  INV_X1 U9723 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8589) );
  NAND2_X1 U9724 ( .A1(n8694), .A2(n8589), .ZN(n8590) );
  AND2_X1 U9725 ( .A1(n8710), .A2(n8590), .ZN(n9936) );
  NAND2_X1 U9726 ( .A1(n7099), .A2(n9936), .ZN(n8593) );
  NAND2_X1 U9727 ( .A1(n5051), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8592) );
  NAND2_X1 U9728 ( .A1(n5038), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8591) );
  NAND4_X1 U9729 ( .A1(n8594), .A2(n8593), .A3(n8592), .A4(n8591), .ZN(n9953)
         );
  NAND2_X1 U9730 ( .A1(n9953), .A2(n7104), .ZN(n8595) );
  NAND2_X1 U9731 ( .A1(n8596), .A2(n8595), .ZN(n8597) );
  XNOR2_X1 U9732 ( .A(n8597), .B(n8724), .ZN(n9733) );
  INV_X1 U9733 ( .A(n9733), .ZN(n8706) );
  AND2_X1 U9734 ( .A1(n9953), .A2(n8790), .ZN(n8598) );
  AOI21_X1 U9735 ( .B1(n10099), .B2(n8676), .A(n8598), .ZN(n9732) );
  INV_X1 U9736 ( .A(n9732), .ZN(n8705) );
  NAND2_X1 U9737 ( .A1(n8599), .A2(n8749), .ZN(n8602) );
  OR2_X1 U9738 ( .A1(n7183), .A2(n8600), .ZN(n8601) );
  INV_X1 U9739 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8604) );
  NAND2_X1 U9740 ( .A1(n8604), .A2(n8603), .ZN(n8605) );
  AND2_X1 U9741 ( .A1(n8605), .A2(n8692), .ZN(n9966) );
  NAND2_X1 U9742 ( .A1(n7099), .A2(n9966), .ZN(n8609) );
  NAND2_X1 U9743 ( .A1(n7351), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8608) );
  NAND2_X1 U9744 ( .A1(n5051), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8607) );
  NAND2_X1 U9745 ( .A1(n5039), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8606) );
  NAND4_X1 U9746 ( .A1(n8609), .A2(n8608), .A3(n8607), .A4(n8606), .ZN(n9988)
         );
  AOI22_X1 U9747 ( .A1(n10109), .A2(n5040), .B1(n8790), .B2(n9988), .ZN(n9705)
         );
  NAND2_X1 U9748 ( .A1(n8610), .A2(n8749), .ZN(n8612) );
  AOI22_X1 U9749 ( .A1(n8638), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10021), 
        .B2(n8637), .ZN(n8611) );
  NAND2_X1 U9750 ( .A1(n10130), .A2(n8795), .ZN(n8623) );
  INV_X1 U9751 ( .A(n8613), .ZN(n8617) );
  NAND2_X1 U9752 ( .A1(n8615), .A2(n8614), .ZN(n8616) );
  NAND2_X1 U9753 ( .A1(n8617), .A2(n8616), .ZN(n10034) );
  INV_X1 U9754 ( .A(n7099), .ZN(n8618) );
  OR2_X1 U9755 ( .A1(n10034), .A2(n8618), .ZN(n8621) );
  AOI22_X1 U9756 ( .A1(n5051), .A2(P1_REG0_REG_19__SCAN_IN), .B1(n5039), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n8620) );
  NAND2_X1 U9757 ( .A1(n5052), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n8619) );
  OR2_X1 U9758 ( .A1(n10014), .A2(n7961), .ZN(n8622) );
  NAND2_X1 U9759 ( .A1(n8623), .A2(n8622), .ZN(n8624) );
  XNOR2_X1 U9760 ( .A(n8624), .B(n8793), .ZN(n8650) );
  INV_X1 U9761 ( .A(n8790), .ZN(n8699) );
  NOR2_X1 U9762 ( .A1(n10014), .A2(n8699), .ZN(n8625) );
  AOI21_X1 U9763 ( .B1(n10130), .B2(n8676), .A(n8625), .ZN(n8646) );
  INV_X1 U9764 ( .A(n8646), .ZN(n8649) );
  NAND2_X1 U9765 ( .A1(n10541), .A2(n8795), .ZN(n8627) );
  NAND2_X1 U9766 ( .A1(n10978), .A2(n8676), .ZN(n8626) );
  NAND2_X1 U9767 ( .A1(n8627), .A2(n8626), .ZN(n8628) );
  XNOR2_X1 U9768 ( .A(n8628), .B(n8724), .ZN(n8630) );
  AND2_X1 U9769 ( .A1(n10978), .A2(n8790), .ZN(n8629) );
  AOI21_X1 U9770 ( .B1(n10541), .B2(n8676), .A(n8629), .ZN(n8631) );
  NAND2_X1 U9771 ( .A1(n8630), .A2(n8631), .ZN(n8635) );
  INV_X1 U9772 ( .A(n8630), .ZN(n8633) );
  INV_X1 U9773 ( .A(n8631), .ZN(n8632) );
  NAND2_X1 U9774 ( .A1(n8633), .A2(n8632), .ZN(n8634) );
  AND2_X1 U9775 ( .A1(n8635), .A2(n8634), .ZN(n9743) );
  NAND2_X1 U9776 ( .A1(n8636), .A2(n8749), .ZN(n8640) );
  AOI22_X1 U9777 ( .A1(n8638), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8637), .B2(
        n9882), .ZN(n8639) );
  NAND2_X1 U9778 ( .A1(n10534), .A2(n8795), .ZN(n8642) );
  NAND2_X1 U9779 ( .A1(n10041), .A2(n8676), .ZN(n8641) );
  NAND2_X1 U9780 ( .A1(n8642), .A2(n8641), .ZN(n8643) );
  XNOR2_X1 U9781 ( .A(n8643), .B(n8724), .ZN(n8647) );
  NAND2_X1 U9782 ( .A1(n10534), .A2(n8676), .ZN(n8645) );
  NAND2_X1 U9783 ( .A1(n10041), .A2(n8790), .ZN(n8644) );
  NAND2_X1 U9784 ( .A1(n8645), .A2(n8644), .ZN(n9785) );
  NAND2_X1 U9785 ( .A1(n9786), .A2(n9785), .ZN(n9790) );
  XNOR2_X1 U9786 ( .A(n8650), .B(n8646), .ZN(n9714) );
  INV_X1 U9787 ( .A(n8647), .ZN(n8648) );
  NAND2_X2 U9788 ( .A1(n5098), .A2(n8648), .ZN(n9787) );
  NAND2_X1 U9789 ( .A1(n8651), .A2(n8749), .ZN(n8654) );
  OR2_X1 U9790 ( .A1(n7509), .A2(n8652), .ZN(n8653) );
  NAND2_X1 U9791 ( .A1(n10126), .A2(n8795), .ZN(n8656) );
  NAND2_X1 U9792 ( .A1(n10040), .A2(n8676), .ZN(n8655) );
  NAND2_X1 U9793 ( .A1(n8656), .A2(n8655), .ZN(n8657) );
  XNOR2_X1 U9794 ( .A(n8657), .B(n8793), .ZN(n8661) );
  NAND2_X1 U9795 ( .A1(n10126), .A2(n8676), .ZN(n8659) );
  NAND2_X1 U9796 ( .A1(n10040), .A2(n8790), .ZN(n8658) );
  NAND2_X1 U9797 ( .A1(n8659), .A2(n8658), .ZN(n8660) );
  NOR2_X1 U9798 ( .A1(n8661), .A2(n8660), .ZN(n9763) );
  NAND2_X1 U9799 ( .A1(n8661), .A2(n8660), .ZN(n9764) );
  NAND2_X1 U9800 ( .A1(n8662), .A2(n8749), .ZN(n8665) );
  OR2_X1 U9801 ( .A1(n7509), .A2(n8663), .ZN(n8664) );
  NAND2_X1 U9802 ( .A1(n10120), .A2(n8795), .ZN(n8673) );
  OR2_X1 U9803 ( .A1(n8666), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8668) );
  AND2_X1 U9804 ( .A1(n8668), .A2(n8667), .ZN(n10001) );
  NAND2_X1 U9805 ( .A1(n10001), .A2(n7099), .ZN(n8671) );
  AOI22_X1 U9806 ( .A1(n7351), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n5051), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n8670) );
  NAND2_X1 U9807 ( .A1(n5039), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8669) );
  AND3_X1 U9808 ( .A1(n8671), .A2(n8670), .A3(n8669), .ZN(n10016) );
  OR2_X1 U9809 ( .A1(n10016), .A2(n7961), .ZN(n8672) );
  NAND2_X1 U9810 ( .A1(n8673), .A2(n8672), .ZN(n8674) );
  XNOR2_X1 U9811 ( .A(n8674), .B(n8724), .ZN(n8678) );
  NOR2_X1 U9812 ( .A1(n10016), .A2(n8699), .ZN(n8675) );
  AOI21_X1 U9813 ( .B1(n10120), .B2(n8676), .A(n8675), .ZN(n8677) );
  NOR2_X1 U9814 ( .A1(n8678), .A2(n8677), .ZN(n9723) );
  NAND2_X1 U9815 ( .A1(n8678), .A2(n8677), .ZN(n9721) );
  NAND2_X1 U9816 ( .A1(n8679), .A2(n8749), .ZN(n8681) );
  OR2_X1 U9817 ( .A1(n7183), .A2(n10266), .ZN(n8680) );
  INV_X1 U9818 ( .A(n9997), .ZN(n9728) );
  OAI22_X1 U9819 ( .A1(n9983), .A2(n8716), .B1(n9728), .B2(n7961), .ZN(n8682)
         );
  XNOR2_X1 U9820 ( .A(n8682), .B(n8793), .ZN(n8684) );
  OAI22_X1 U9821 ( .A1(n9983), .A2(n7961), .B1(n9728), .B2(n8699), .ZN(n8683)
         );
  NAND2_X1 U9822 ( .A1(n8684), .A2(n8683), .ZN(n9775) );
  NOR2_X1 U9823 ( .A1(n8684), .A2(n8683), .ZN(n9774) );
  AOI21_X2 U9824 ( .B1(n9778), .B2(n9775), .A(n9774), .ZN(n8687) );
  AOI22_X1 U9825 ( .A1(n10109), .A2(n8795), .B1(n5040), .B2(n9988), .ZN(n8685)
         );
  XNOR2_X1 U9826 ( .A(n8685), .B(n8724), .ZN(n8686) );
  NAND2_X1 U9827 ( .A1(n8687), .A2(n8686), .ZN(n9703) );
  NAND2_X1 U9828 ( .A1(n8688), .A2(n8749), .ZN(n8690) );
  OR2_X1 U9829 ( .A1(n7183), .A2(n10264), .ZN(n8689) );
  INV_X1 U9830 ( .A(n10105), .ZN(n9949) );
  NAND2_X1 U9831 ( .A1(n7351), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8698) );
  INV_X1 U9832 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8691) );
  NAND2_X1 U9833 ( .A1(n8692), .A2(n8691), .ZN(n8693) );
  AND2_X1 U9834 ( .A1(n8694), .A2(n8693), .ZN(n9957) );
  NAND2_X1 U9835 ( .A1(n7099), .A2(n9957), .ZN(n8697) );
  NAND2_X1 U9836 ( .A1(n5051), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8696) );
  NAND2_X1 U9837 ( .A1(n5038), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8695) );
  NAND4_X1 U9838 ( .A1(n8698), .A2(n8697), .A3(n8696), .A4(n8695), .ZN(n9971)
         );
  INV_X1 U9839 ( .A(n9971), .ZN(n9709) );
  OAI22_X1 U9840 ( .A1(n9949), .A2(n7961), .B1(n9709), .B2(n8699), .ZN(n8704)
         );
  NAND2_X1 U9841 ( .A1(n10105), .A2(n8795), .ZN(n8701) );
  NAND2_X1 U9842 ( .A1(n9971), .A2(n5040), .ZN(n8700) );
  NAND2_X1 U9843 ( .A1(n8701), .A2(n8700), .ZN(n8702) );
  XNOR2_X1 U9844 ( .A(n8702), .B(n8724), .ZN(n8703) );
  XOR2_X1 U9845 ( .A(n8704), .B(n8703), .Z(n9756) );
  OR2_X1 U9846 ( .A1(n7183), .A2(n10576), .ZN(n8707) );
  NAND2_X1 U9847 ( .A1(n7351), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8715) );
  INV_X1 U9848 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8709) );
  NAND2_X1 U9849 ( .A1(n8710), .A2(n8709), .ZN(n8711) );
  NAND2_X1 U9850 ( .A1(n7099), .A2(n9925), .ZN(n8714) );
  NAND2_X1 U9851 ( .A1(n5051), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8713) );
  NAND2_X1 U9852 ( .A1(n5038), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8712) );
  NAND4_X1 U9853 ( .A1(n8715), .A2(n8714), .A3(n8713), .A4(n8712), .ZN(n9942)
         );
  OAI22_X1 U9854 ( .A1(n10094), .A2(n8716), .B1(n9738), .B2(n7961), .ZN(n8717)
         );
  XNOR2_X1 U9855 ( .A(n8717), .B(n8724), .ZN(n8719) );
  AND2_X1 U9856 ( .A1(n9942), .A2(n8790), .ZN(n8718) );
  AOI21_X1 U9857 ( .B1(n9922), .B2(n5040), .A(n8718), .ZN(n8720) );
  XNOR2_X1 U9858 ( .A(n8719), .B(n8720), .ZN(n9802) );
  OR2_X1 U9859 ( .A1(n7183), .A2(n10253), .ZN(n8721) );
  NAND2_X1 U9860 ( .A1(n10088), .A2(n8795), .ZN(n8723) );
  NAND2_X1 U9861 ( .A1(n9915), .A2(n7104), .ZN(n8722) );
  NAND2_X1 U9862 ( .A1(n8723), .A2(n8722), .ZN(n8725) );
  XNOR2_X1 U9863 ( .A(n8725), .B(n8724), .ZN(n8728) );
  AND2_X1 U9864 ( .A1(n9915), .A2(n8790), .ZN(n8726) );
  AOI21_X1 U9865 ( .B1(n10088), .B2(n5040), .A(n8726), .ZN(n8727) );
  NAND2_X1 U9866 ( .A1(n8728), .A2(n8727), .ZN(n8801) );
  OAI21_X1 U9867 ( .B1(n8728), .B2(n8727), .A(n8801), .ZN(n8729) );
  INV_X1 U9868 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8731) );
  OAI22_X1 U9869 ( .A1(n9794), .A2(n9738), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8731), .ZN(n8740) );
  NAND2_X1 U9870 ( .A1(n5052), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8738) );
  INV_X1 U9871 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8730) );
  OAI21_X1 U9872 ( .B1(n8732), .B2(n8731), .A(n8730), .ZN(n8733) );
  NAND2_X1 U9873 ( .A1(n7099), .A2(n9138), .ZN(n8737) );
  NAND2_X1 U9874 ( .A1(n5051), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8736) );
  NAND2_X1 U9875 ( .A1(n5038), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8735) );
  NAND4_X1 U9876 ( .A1(n8738), .A2(n8737), .A3(n8736), .A4(n8735), .ZN(n9905)
         );
  INV_X1 U9877 ( .A(n9905), .ZN(n8841) );
  NOR2_X1 U9878 ( .A1(n9808), .A2(n8841), .ZN(n8739) );
  AOI211_X1 U9879 ( .C1(n9804), .C2(n9906), .A(n8740), .B(n8739), .ZN(n8742)
         );
  NAND2_X1 U9880 ( .A1(n10088), .A2(n9811), .ZN(n8741) );
  INV_X1 U9881 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n8743) );
  NOR2_X1 U9882 ( .A1(n7183), .A2(n8743), .ZN(n8744) );
  NAND2_X1 U9883 ( .A1(n9693), .A2(n8749), .ZN(n8746) );
  INV_X1 U9884 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10567) );
  OR2_X1 U9885 ( .A1(n7183), .A2(n10567), .ZN(n8745) );
  NAND2_X1 U9886 ( .A1(n9060), .A2(n8749), .ZN(n8748) );
  INV_X1 U9887 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10246) );
  OR2_X1 U9888 ( .A1(n7183), .A2(n10246), .ZN(n8747) );
  NAND2_X1 U9889 ( .A1(n9144), .A2(n8749), .ZN(n8751) );
  INV_X1 U9890 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9145) );
  OR2_X1 U9891 ( .A1(n7183), .A2(n9145), .ZN(n8750) );
  INV_X1 U9892 ( .A(n10083), .ZN(n9140) );
  INV_X1 U9893 ( .A(n10099), .ZN(n9938) );
  INV_X1 U9894 ( .A(n10130), .ZN(n10037) );
  INV_X1 U9895 ( .A(n10126), .ZN(n8752) );
  AND2_X2 U9896 ( .A1(n9965), .A2(n9949), .ZN(n9955) );
  INV_X1 U9897 ( .A(n10088), .ZN(n9902) );
  NAND2_X1 U9898 ( .A1(n10077), .A2(n9892), .ZN(n10073) );
  NAND2_X1 U9899 ( .A1(n10071), .A2(n10068), .ZN(n8758) );
  NAND2_X1 U9900 ( .A1(n5052), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U9901 ( .A1(n5039), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8754) );
  NAND2_X1 U9902 ( .A1(n5051), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8753) );
  NAND3_X1 U9903 ( .A1(n8755), .A2(n8754), .A3(n8753), .ZN(n9815) );
  INV_X1 U9904 ( .A(P1_B_REG_SCAN_IN), .ZN(n9040) );
  OR2_X1 U9905 ( .A1(n5050), .A2(n9040), .ZN(n8756) );
  AND2_X1 U9906 ( .A1(n10977), .A2(n8756), .ZN(n9160) );
  NAND2_X1 U9907 ( .A1(n9815), .A2(n9160), .ZN(n10075) );
  NOR2_X1 U9908 ( .A1(n10738), .A2(n10075), .ZN(n9895) );
  AOI21_X1 U9909 ( .B1(n11006), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9895), .ZN(
        n8757) );
  OAI211_X1 U9910 ( .C1(n10072), .C2(n10734), .A(n8758), .B(n8757), .ZN(
        P1_U3261) );
  NAND2_X1 U9911 ( .A1(n9244), .A2(n9270), .ZN(n8764) );
  NAND2_X1 U9912 ( .A1(n9247), .A2(n9272), .ZN(n8763) );
  NAND2_X1 U9913 ( .A1(n9246), .A2(n8760), .ZN(n8761) );
  NAND4_X1 U9914 ( .A1(n8764), .A2(n8763), .A3(n8762), .A4(n8761), .ZN(n8765)
         );
  AOI21_X1 U9915 ( .B1(n9664), .B2(n9261), .A(n8765), .ZN(n8773) );
  INV_X1 U9916 ( .A(n8766), .ZN(n8770) );
  OAI22_X1 U9917 ( .A1(n8768), .A2(n5042), .B1(n8767), .B2(n9240), .ZN(n8769)
         );
  NAND3_X1 U9918 ( .A1(n8771), .A2(n8770), .A3(n8769), .ZN(n8772) );
  OAI211_X1 U9919 ( .C1(n9056), .C2(n5042), .A(n8773), .B(n8772), .ZN(P2_U3217) );
  NAND2_X1 U9920 ( .A1(n9248), .A2(n10795), .ZN(n8776) );
  INV_X1 U9921 ( .A(n8774), .ZN(n8775) );
  NAND2_X1 U9922 ( .A1(n8776), .A2(n8775), .ZN(n8779) );
  OAI22_X1 U9923 ( .A1(n8781), .A2(n9230), .B1(n9229), .B2(n8777), .ZN(n8778)
         );
  AOI211_X1 U9924 ( .C1(n10797), .C2(n9246), .A(n8779), .B(n8778), .ZN(n8787)
         );
  OAI22_X1 U9925 ( .A1(n9240), .A2(n8781), .B1(n5042), .B2(n8780), .ZN(n8785)
         );
  INV_X1 U9926 ( .A(n8783), .ZN(n8784) );
  NAND3_X1 U9927 ( .A1(n8785), .A2(n9216), .A3(n8784), .ZN(n8786) );
  OAI211_X1 U9928 ( .C1(n5042), .C2(n8788), .A(n8787), .B(n8786), .ZN(P2_U3229) );
  INV_X1 U9929 ( .A(n8789), .ZN(n10573) );
  OAI222_X1 U9930 ( .A1(P2_U3152), .A2(n9091), .B1(n5043), .B2(n10573), .C1(
        n9698), .C2(n6285), .ZN(P2_U3331) );
  NAND2_X1 U9931 ( .A1(n10083), .A2(n7104), .ZN(n8792) );
  NAND2_X1 U9932 ( .A1(n9905), .A2(n8790), .ZN(n8791) );
  NAND2_X1 U9933 ( .A1(n8792), .A2(n8791), .ZN(n8794) );
  XNOR2_X1 U9934 ( .A(n8794), .B(n8793), .ZN(n8797) );
  AOI22_X1 U9935 ( .A1(n10083), .A2(n8795), .B1(n5040), .B2(n9905), .ZN(n8796)
         );
  XNOR2_X1 U9936 ( .A(n8797), .B(n8796), .ZN(n8798) );
  INV_X1 U9937 ( .A(n8798), .ZN(n8802) );
  NAND3_X1 U9938 ( .A1(n8802), .A2(n9744), .A3(n8801), .ZN(n8807) );
  NAND3_X1 U9939 ( .A1(n8808), .A2(n9744), .A3(n8798), .ZN(n8806) );
  NAND2_X1 U9940 ( .A1(n9804), .A2(n9138), .ZN(n8800) );
  AOI22_X1 U9941 ( .A1(n9805), .A2(n9915), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8799) );
  OAI211_X1 U9942 ( .C1(n9133), .C2(n9808), .A(n8800), .B(n8799), .ZN(n8804)
         );
  NOR3_X1 U9943 ( .A1(n8802), .A2(n9813), .A3(n8801), .ZN(n8803) );
  AOI211_X1 U9944 ( .C1(n10083), .C2(n9811), .A(n8804), .B(n8803), .ZN(n8805)
         );
  OAI211_X1 U9945 ( .C1(n8808), .C2(n8807), .A(n8806), .B(n8805), .ZN(P1_U3218) );
  INV_X1 U9946 ( .A(n10072), .ZN(n8876) );
  INV_X1 U9947 ( .A(n9815), .ZN(n8981) );
  NAND2_X1 U9948 ( .A1(n8876), .A2(n8981), .ZN(n8984) );
  NAND2_X1 U9949 ( .A1(n7351), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8811) );
  NAND2_X1 U9950 ( .A1(n5038), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8810) );
  NAND2_X1 U9951 ( .A1(n5051), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8809) );
  NAND3_X1 U9952 ( .A1(n8811), .A2(n8810), .A3(n8809), .ZN(n9816) );
  INV_X1 U9953 ( .A(n9816), .ZN(n8869) );
  OR2_X1 U9954 ( .A1(n9893), .A2(n8869), .ZN(n8982) );
  NAND2_X1 U9955 ( .A1(n8984), .A2(n8982), .ZN(n9017) );
  INV_X1 U9956 ( .A(n9017), .ZN(n8872) );
  NAND2_X1 U9957 ( .A1(n9014), .A2(n9155), .ZN(n9026) );
  INV_X1 U9958 ( .A(n9026), .ZN(n8967) );
  INV_X1 U9959 ( .A(n9915), .ZN(n9809) );
  INV_X1 U9960 ( .A(n9953), .ZN(n9759) );
  OR2_X1 U9961 ( .A1(n10099), .A2(n9759), .ZN(n8959) );
  NAND3_X1 U9962 ( .A1(n9129), .A2(n8879), .A3(n8959), .ZN(n8849) );
  OR2_X1 U9963 ( .A1(n10105), .A2(n9709), .ZN(n8956) );
  INV_X1 U9964 ( .A(n9988), .ZN(n9781) );
  OR2_X1 U9965 ( .A1(n10109), .A2(n9781), .ZN(n8953) );
  AND2_X1 U9966 ( .A1(n8956), .A2(n8953), .ZN(n8847) );
  OR2_X1 U9967 ( .A1(n10120), .A2(n10016), .ZN(n8940) );
  INV_X1 U9968 ( .A(n10040), .ZN(n8815) );
  NAND2_X1 U9969 ( .A1(n10126), .A2(n8815), .ZN(n9123) );
  NAND2_X1 U9970 ( .A1(n8940), .A2(n5328), .ZN(n8812) );
  NAND2_X1 U9971 ( .A1(n10120), .A2(n10016), .ZN(n9124) );
  AND2_X1 U9972 ( .A1(n8812), .A2(n9124), .ZN(n8946) );
  NAND2_X1 U9973 ( .A1(n10130), .A2(n10014), .ZN(n9122) );
  NAND2_X1 U9974 ( .A1(n10114), .A2(n9728), .ZN(n9125) );
  NAND3_X1 U9975 ( .A1(n8946), .A2(n9122), .A3(n9125), .ZN(n8836) );
  INV_X1 U9976 ( .A(n10041), .ZN(n9749) );
  NAND2_X1 U9977 ( .A1(n10534), .A2(n9749), .ZN(n8935) );
  INV_X1 U9978 ( .A(n10059), .ZN(n10053) );
  NAND2_X1 U9979 ( .A1(n8935), .A2(n10053), .ZN(n8813) );
  OR2_X1 U9980 ( .A1(n10534), .A2(n9749), .ZN(n8936) );
  OR2_X1 U9981 ( .A1(n10130), .A2(n10014), .ZN(n8942) );
  AND2_X1 U9982 ( .A1(n9120), .A2(n8942), .ZN(n8814) );
  OR2_X1 U9983 ( .A1(n8836), .A2(n8814), .ZN(n8818) );
  OR2_X1 U9984 ( .A1(n10126), .A2(n8815), .ZN(n8941) );
  NAND2_X1 U9985 ( .A1(n8940), .A2(n8941), .ZN(n8948) );
  NAND3_X1 U9986 ( .A1(n8946), .A2(n9125), .A3(n8948), .ZN(n8816) );
  NAND2_X1 U9987 ( .A1(n9983), .A2(n9997), .ZN(n8947) );
  AND2_X1 U9988 ( .A1(n8816), .A2(n8947), .ZN(n8817) );
  NAND2_X1 U9989 ( .A1(n8818), .A2(n8817), .ZN(n8844) );
  AND2_X1 U9990 ( .A1(n10057), .A2(n8930), .ZN(n8819) );
  AND2_X1 U9991 ( .A1(n8935), .A2(n8819), .ZN(n9119) );
  NAND2_X1 U9992 ( .A1(n8925), .A2(n8921), .ZN(n8832) );
  NAND2_X1 U9993 ( .A1(n8915), .A2(n8820), .ZN(n8910) );
  INV_X1 U9994 ( .A(n8897), .ZN(n8821) );
  NAND2_X1 U9995 ( .A1(n8901), .A2(n8821), .ZN(n8822) );
  NAND4_X1 U9996 ( .A1(n8913), .A2(n8906), .A3(n8902), .A4(n8822), .ZN(n8829)
         );
  AND3_X1 U9997 ( .A1(n8901), .A2(n8892), .A3(n8898), .ZN(n8824) );
  INV_X1 U9998 ( .A(n8913), .ZN(n8823) );
  OAI22_X1 U9999 ( .A1(n8829), .A2(n8824), .B1(n8823), .B2(n8905), .ZN(n8825)
         );
  OAI21_X1 U10000 ( .B1(n8910), .B2(n8825), .A(n8917), .ZN(n8826) );
  AND2_X1 U10001 ( .A1(n8826), .A2(n8922), .ZN(n8827) );
  OAI211_X1 U10002 ( .C1(n8832), .C2(n8827), .A(n8929), .B(n8926), .ZN(n8828)
         );
  NAND2_X1 U10003 ( .A1(n9119), .A2(n8828), .ZN(n8845) );
  INV_X1 U10004 ( .A(n8829), .ZN(n8830) );
  NAND4_X1 U10005 ( .A1(n8917), .A2(n8830), .A3(n8891), .A4(n8889), .ZN(n8831)
         );
  NOR2_X1 U10006 ( .A1(n8832), .A2(n8831), .ZN(n8833) );
  NAND2_X1 U10007 ( .A1(n9119), .A2(n8833), .ZN(n8834) );
  AND2_X1 U10008 ( .A1(n8845), .A2(n8834), .ZN(n8835) );
  NOR2_X1 U10009 ( .A1(n8836), .A2(n8835), .ZN(n8837) );
  NAND2_X1 U10010 ( .A1(n10109), .A2(n9781), .ZN(n9126) );
  OAI21_X1 U10011 ( .B1(n8844), .B2(n8837), .A(n9126), .ZN(n8838) );
  NAND2_X1 U10012 ( .A1(n8847), .A2(n8838), .ZN(n8839) );
  NAND2_X1 U10013 ( .A1(n10099), .A2(n9759), .ZN(n9128) );
  NAND2_X1 U10014 ( .A1(n10105), .A2(n9709), .ZN(n9127) );
  AND3_X1 U10015 ( .A1(n8839), .A2(n9128), .A3(n9127), .ZN(n8843) );
  NAND2_X1 U10016 ( .A1(n9922), .A2(n9738), .ZN(n9903) );
  INV_X1 U10017 ( .A(n9903), .ZN(n8878) );
  NAND2_X1 U10018 ( .A1(n9129), .A2(n8878), .ZN(n8840) );
  NAND2_X1 U10019 ( .A1(n10088), .A2(n9809), .ZN(n8963) );
  AND2_X1 U10020 ( .A1(n8840), .A2(n8963), .ZN(n8842) );
  NAND2_X1 U10021 ( .A1(n10083), .A2(n8841), .ZN(n9157) );
  OAI211_X1 U10022 ( .C1(n8849), .C2(n8843), .A(n8842), .B(n9157), .ZN(n9021)
         );
  INV_X1 U10023 ( .A(n9021), .ZN(n8867) );
  INV_X1 U10024 ( .A(n8844), .ZN(n8846) );
  NAND3_X1 U10025 ( .A1(n8847), .A2(n8846), .A3(n8845), .ZN(n8848) );
  NOR2_X1 U10026 ( .A1(n8849), .A2(n8848), .ZN(n9022) );
  NAND3_X1 U10027 ( .A1(n8851), .A2(n8850), .A3(n6957), .ZN(n8853) );
  NAND2_X1 U10028 ( .A1(n8853), .A2(n8852), .ZN(n8855) );
  OAI21_X1 U10029 ( .B1(n8856), .B2(n8855), .A(n8854), .ZN(n8858) );
  NAND2_X1 U10030 ( .A1(n8858), .A2(n8857), .ZN(n8861) );
  NAND3_X1 U10031 ( .A1(n8861), .A2(n8860), .A3(n8859), .ZN(n8863) );
  NAND2_X1 U10032 ( .A1(n8863), .A2(n8862), .ZN(n8864) );
  NAND4_X1 U10033 ( .A1(n9022), .A2(n8888), .A3(n8865), .A4(n8864), .ZN(n8866)
         );
  NAND2_X1 U10034 ( .A1(n8867), .A2(n8866), .ZN(n8868) );
  NAND2_X1 U10035 ( .A1(n8967), .A2(n8868), .ZN(n8870) );
  AND2_X1 U10036 ( .A1(n9893), .A2(n8869), .ZN(n9016) );
  INV_X1 U10037 ( .A(n9016), .ZN(n8874) );
  NAND3_X1 U10038 ( .A1(n8870), .A2(n8874), .A3(n9024), .ZN(n8871) );
  AND2_X1 U10039 ( .A1(n10072), .A2(n9815), .ZN(n9028) );
  AOI21_X1 U10040 ( .B1(n8872), .B2(n8871), .A(n9028), .ZN(n8873) );
  XNOR2_X1 U10041 ( .A(n8873), .B(n9958), .ZN(n9039) );
  NAND3_X1 U10042 ( .A1(n8982), .A2(n8874), .A3(n9815), .ZN(n8875) );
  OAI21_X1 U10043 ( .B1(n8876), .B2(n9893), .A(n8875), .ZN(n8970) );
  INV_X1 U10044 ( .A(n8879), .ZN(n8877) );
  MUX2_X1 U10045 ( .A(n8878), .B(n8877), .S(n8972), .Z(n8966) );
  INV_X1 U10046 ( .A(n8972), .ZN(n8977) );
  XNOR2_X1 U10047 ( .A(n8880), .B(n8972), .ZN(n8887) );
  NAND2_X1 U10048 ( .A1(n8888), .A2(n8881), .ZN(n8884) );
  NAND2_X1 U10049 ( .A1(n8889), .A2(n8882), .ZN(n8883) );
  MUX2_X1 U10050 ( .A(n8884), .B(n8883), .S(n8972), .Z(n8885) );
  AOI21_X1 U10051 ( .B1(n8887), .B2(n8886), .A(n8885), .ZN(n8896) );
  MUX2_X1 U10052 ( .A(n8889), .B(n8888), .S(n8972), .Z(n8890) );
  NAND2_X1 U10053 ( .A1(n8890), .A2(n9002), .ZN(n8895) );
  MUX2_X1 U10054 ( .A(n8892), .B(n8891), .S(n8972), .Z(n8893) );
  OAI211_X1 U10055 ( .C1(n8896), .C2(n8895), .A(n8894), .B(n8893), .ZN(n8900)
         );
  MUX2_X1 U10056 ( .A(n8898), .B(n8897), .S(n8977), .Z(n8899) );
  NAND3_X1 U10057 ( .A1(n8900), .A2(n9003), .A3(n8899), .ZN(n8904) );
  MUX2_X1 U10058 ( .A(n8902), .B(n8901), .S(n8977), .Z(n8903) );
  NAND3_X1 U10059 ( .A1(n8904), .A2(n5266), .A3(n8903), .ZN(n8909) );
  MUX2_X1 U10060 ( .A(n8906), .B(n8905), .S(n8972), .Z(n8907) );
  AND2_X1 U10061 ( .A1(n9004), .A2(n8907), .ZN(n8908) );
  NAND2_X1 U10062 ( .A1(n8909), .A2(n8908), .ZN(n8914) );
  INV_X1 U10063 ( .A(n8910), .ZN(n8912) );
  INV_X1 U10064 ( .A(n8917), .ZN(n8911) );
  AOI21_X1 U10065 ( .B1(n8914), .B2(n8912), .A(n8911), .ZN(n8920) );
  NAND2_X1 U10066 ( .A1(n8914), .A2(n8913), .ZN(n8916) );
  NAND2_X1 U10067 ( .A1(n8916), .A2(n8915), .ZN(n8918) );
  NAND2_X1 U10068 ( .A1(n8918), .A2(n8917), .ZN(n8919) );
  MUX2_X1 U10069 ( .A(n8920), .B(n8919), .S(n8972), .Z(n8924) );
  MUX2_X1 U10070 ( .A(n8922), .B(n8921), .S(n8977), .Z(n8923) );
  OAI211_X1 U10071 ( .C1(n8924), .C2(n9007), .A(n9009), .B(n8923), .ZN(n8928)
         );
  MUX2_X1 U10072 ( .A(n8926), .B(n8925), .S(n8972), .Z(n8927) );
  NAND3_X1 U10073 ( .A1(n8928), .A2(n10974), .A3(n8927), .ZN(n8933) );
  MUX2_X1 U10074 ( .A(n8930), .B(n8929), .S(n8972), .Z(n8932) );
  AOI21_X1 U10075 ( .B1(n8933), .B2(n8932), .A(n8931), .ZN(n8939) );
  MUX2_X1 U10076 ( .A(n10057), .B(n10059), .S(n8972), .Z(n8934) );
  NAND2_X1 U10077 ( .A1(n10060), .A2(n8934), .ZN(n8938) );
  INV_X1 U10078 ( .A(n10031), .ZN(n10039) );
  MUX2_X1 U10079 ( .A(n8936), .B(n8935), .S(n8972), .Z(n8937) );
  OAI211_X1 U10080 ( .C1(n8939), .C2(n8938), .A(n10039), .B(n8937), .ZN(n8944)
         );
  MUX2_X1 U10081 ( .A(n8942), .B(n9122), .S(n8977), .Z(n8943) );
  NAND4_X1 U10082 ( .A1(n8944), .A2(n10003), .A3(n10012), .A4(n8943), .ZN(
        n8945) );
  NAND2_X1 U10083 ( .A1(n8947), .A2(n9125), .ZN(n9977) );
  INV_X1 U10084 ( .A(n9977), .ZN(n9986) );
  OAI211_X1 U10085 ( .C1(n8977), .C2(n8946), .A(n8945), .B(n9986), .ZN(n8950)
         );
  NAND2_X1 U10086 ( .A1(n8950), .A2(n8947), .ZN(n8952) );
  AND2_X1 U10087 ( .A1(n8948), .A2(n9124), .ZN(n8949) );
  OAI21_X1 U10088 ( .B1(n8950), .B2(n8949), .A(n9125), .ZN(n8951) );
  MUX2_X1 U10089 ( .A(n8952), .B(n8951), .S(n8977), .Z(n8955) );
  INV_X1 U10090 ( .A(n9970), .ZN(n9964) );
  MUX2_X1 U10091 ( .A(n8953), .B(n9126), .S(n8972), .Z(n8954) );
  OAI211_X1 U10092 ( .C1(n8955), .C2(n9964), .A(n9952), .B(n8954), .ZN(n8958)
         );
  MUX2_X1 U10093 ( .A(n9127), .B(n8956), .S(n8972), .Z(n8957) );
  NAND3_X1 U10094 ( .A1(n8958), .A2(n9941), .A3(n8957), .ZN(n8961) );
  MUX2_X1 U10095 ( .A(n8959), .B(n9128), .S(n8972), .Z(n8960) );
  NAND3_X1 U10096 ( .A1(n9914), .A2(n8961), .A3(n8960), .ZN(n8962) );
  NAND2_X1 U10097 ( .A1(n9904), .A2(n8962), .ZN(n8965) );
  MUX2_X1 U10098 ( .A(n9129), .B(n8963), .S(n8972), .Z(n8964) );
  OAI211_X1 U10099 ( .C1(n8966), .C2(n8965), .A(n9130), .B(n8964), .ZN(n8976)
         );
  NAND2_X1 U10100 ( .A1(n8967), .A2(n8976), .ZN(n8968) );
  NAND3_X1 U10101 ( .A1(n8968), .A2(n8972), .A3(n9024), .ZN(n8969) );
  NAND2_X1 U10102 ( .A1(n8970), .A2(n8969), .ZN(n8975) );
  NAND2_X1 U10103 ( .A1(n9815), .A2(n9816), .ZN(n8971) );
  NAND2_X1 U10104 ( .A1(n9893), .A2(n8971), .ZN(n9025) );
  INV_X1 U10105 ( .A(n9025), .ZN(n8973) );
  NAND3_X1 U10106 ( .A1(n8984), .A2(n8973), .A3(n8972), .ZN(n8974) );
  NAND2_X1 U10107 ( .A1(n8975), .A2(n8974), .ZN(n8980) );
  NAND3_X1 U10108 ( .A1(n8976), .A2(n9157), .A3(n9024), .ZN(n8978) );
  NAND3_X1 U10109 ( .A1(n8978), .A2(n8977), .A3(n9014), .ZN(n8979) );
  NAND2_X1 U10110 ( .A1(n8980), .A2(n8979), .ZN(n8990) );
  OR2_X1 U10111 ( .A1(n8982), .A2(n8981), .ZN(n8983) );
  AND2_X1 U10112 ( .A1(n8984), .A2(n8983), .ZN(n9030) );
  INV_X1 U10113 ( .A(n9030), .ZN(n8986) );
  OAI21_X1 U10114 ( .B1(n8986), .B2(n8985), .A(n10021), .ZN(n8989) );
  INV_X1 U10115 ( .A(n9028), .ZN(n8987) );
  NAND2_X1 U10116 ( .A1(n8987), .A2(n6957), .ZN(n8988) );
  AOI21_X1 U10117 ( .B1(n8990), .B2(n8989), .A(n8988), .ZN(n9036) );
  OR2_X1 U10118 ( .A1(n8990), .A2(n5509), .ZN(n9035) );
  INV_X1 U10119 ( .A(n9904), .ZN(n9013) );
  INV_X1 U10120 ( .A(n9952), .ZN(n9948) );
  INV_X1 U10121 ( .A(n10060), .ZN(n10055) );
  NOR3_X1 U10122 ( .A1(n8993), .A2(n8992), .A3(n7163), .ZN(n8997) );
  NAND4_X1 U10123 ( .A1(n8997), .A2(n8996), .A3(n8995), .A4(n8994), .ZN(n9000)
         );
  NOR4_X1 U10124 ( .A1(n9000), .A2(n8999), .A3(n7448), .A4(n8998), .ZN(n9001)
         );
  NAND4_X1 U10125 ( .A1(n9004), .A2(n9003), .A3(n9002), .A4(n9001), .ZN(n9005)
         );
  NOR4_X1 U10126 ( .A1(n9007), .A2(n8239), .A3(n9006), .A4(n9005), .ZN(n9008)
         );
  NAND4_X1 U10127 ( .A1(n10054), .A2(n10974), .A3(n9009), .A4(n9008), .ZN(
        n9010) );
  NOR4_X1 U10128 ( .A1(n5330), .A2(n10055), .A3(n10031), .A4(n9010), .ZN(n9011) );
  NAND4_X1 U10129 ( .A1(n9970), .A2(n9986), .A3(n10003), .A4(n9011), .ZN(n9012) );
  NOR4_X1 U10130 ( .A1(n9013), .A2(n9948), .A3(n9117), .A4(n9012), .ZN(n9015)
         );
  NAND4_X1 U10131 ( .A1(n9015), .A2(n5073), .A3(n9130), .A4(n9914), .ZN(n9018)
         );
  NOR3_X1 U10132 ( .A1(n9018), .A2(n9017), .A3(n5087), .ZN(n9019) );
  XNOR2_X1 U10133 ( .A(n9019), .B(n9958), .ZN(n9033) );
  INV_X1 U10134 ( .A(n9020), .ZN(n9023) );
  AOI21_X1 U10135 ( .B1(n9023), .B2(n9022), .A(n9021), .ZN(n9027) );
  OAI211_X1 U10136 ( .C1(n9027), .C2(n9026), .A(n9025), .B(n9024), .ZN(n9029)
         );
  AOI21_X1 U10137 ( .B1(n9030), .B2(n9029), .A(n9028), .ZN(n9031) );
  NOR2_X1 U10138 ( .A1(n9031), .A2(n10021), .ZN(n9032) );
  MUX2_X1 U10139 ( .A(n9033), .B(n9032), .S(n6957), .Z(n9034) );
  AOI21_X1 U10140 ( .B1(n9036), .B2(n9035), .A(n9034), .ZN(n9038) );
  AOI21_X1 U10141 ( .B1(n5509), .B2(n9041), .A(n9040), .ZN(n9042) );
  OAI21_X1 U10142 ( .B1(n9043), .B2(n5050), .A(n9042), .ZN(n9044) );
  OAI21_X1 U10143 ( .B1(n9046), .B2(n9045), .A(n9044), .ZN(P1_U3240) );
  AOI22_X1 U10144 ( .A1(n9244), .A2(n9269), .B1(n9246), .B2(n9047), .ZN(n9049)
         );
  OAI211_X1 U10145 ( .C1(n9230), .C2(n9052), .A(n9049), .B(n9048), .ZN(n9050)
         );
  AOI21_X1 U10146 ( .B1(n9659), .B2(n9261), .A(n9050), .ZN(n9058) );
  INV_X1 U10147 ( .A(n9051), .ZN(n9055) );
  OAI22_X1 U10148 ( .A1(n9053), .A2(n5042), .B1(n9052), .B2(n9240), .ZN(n9054)
         );
  NAND3_X1 U10149 ( .A1(n9056), .A2(n9055), .A3(n9054), .ZN(n9057) );
  OAI211_X1 U10150 ( .C1(n9059), .C2(n5042), .A(n9058), .B(n9057), .ZN(
        P2_U3243) );
  INV_X1 U10151 ( .A(n9060), .ZN(n9064) );
  OAI222_X1 U10152 ( .A1(n5043), .A2(n9064), .B1(P2_U3152), .B2(n9062), .C1(
        n9061), .C2(n9698), .ZN(P2_U3329) );
  OAI222_X1 U10153 ( .A1(n5044), .A2(n9064), .B1(n9063), .B2(P1_U3084), .C1(
        n10246), .C2(n10575), .ZN(P1_U3324) );
  INV_X1 U10154 ( .A(n9066), .ZN(n9527) );
  NAND2_X1 U10155 ( .A1(n9506), .A2(n9507), .ZN(n9505) );
  INV_X1 U10156 ( .A(n9641), .ZN(n9069) );
  NAND2_X1 U10157 ( .A1(n9505), .A2(n5634), .ZN(n9496) );
  INV_X1 U10158 ( .A(n9634), .ZN(n9497) );
  NAND2_X1 U10159 ( .A1(n9634), .A2(n9070), .ZN(n9071) );
  INV_X1 U10160 ( .A(n9629), .ZN(n9482) );
  INV_X1 U10161 ( .A(n9466), .ZN(n9072) );
  NAND2_X1 U10162 ( .A1(n9074), .A2(n9073), .ZN(n9075) );
  NAND2_X1 U10163 ( .A1(n9458), .A2(n9075), .ZN(n9448) );
  INV_X1 U10164 ( .A(n9597), .ZN(n9390) );
  INV_X1 U10165 ( .A(n9618), .ZN(n9454) );
  NAND2_X1 U10166 ( .A1(n9548), .A2(n9534), .ZN(n9521) );
  NAND2_X1 U10167 ( .A1(n9497), .A2(n9511), .ZN(n9498) );
  NAND2_X1 U10168 ( .A1(n9405), .A2(n9390), .ZN(n9385) );
  AOI21_X1 U10169 ( .B1(n9083), .B2(n9376), .A(n9364), .ZN(n9587) );
  INV_X1 U10170 ( .A(n9083), .ZN(n9087) );
  INV_X1 U10171 ( .A(n9084), .ZN(n9085) );
  AOI22_X1 U10172 ( .A1(n9085), .A2(n10798), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n7664), .ZN(n9086) );
  OAI21_X1 U10173 ( .B1(n9087), .B2(n9547), .A(n9086), .ZN(n9096) );
  INV_X1 U10174 ( .A(n9088), .ZN(n9089) );
  INV_X1 U10175 ( .A(n9091), .ZN(n9092) );
  AND2_X1 U10176 ( .A1(n9092), .A2(P2_B_REG_SCAN_IN), .ZN(n9093) );
  OR2_X1 U10177 ( .A1(n9559), .A2(n9093), .ZN(n9358) );
  OAI22_X1 U10178 ( .A1(n9166), .A2(n9561), .B1(n9094), .B2(n9358), .ZN(n9095)
         );
  OAI21_X1 U10179 ( .B1(n9590), .B2(n9533), .A(n9097), .ZN(P2_U3267) );
  NAND2_X1 U10180 ( .A1(n9203), .A2(n9098), .ZN(n9100) );
  MUX2_X1 U10181 ( .A(n9100), .B(n9099), .S(n10742), .Z(n9105) );
  OAI21_X1 U10182 ( .B1(n9102), .B2(n9101), .A(n6438), .ZN(n9103) );
  AOI22_X1 U10183 ( .A1(n9220), .A2(n9103), .B1(n9181), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n9104) );
  OAI211_X1 U10184 ( .C1(n6434), .C2(n9229), .A(n9105), .B(n9104), .ZN(
        P2_U3234) );
  INV_X1 U10185 ( .A(n10534), .ZN(n10052) );
  OAI22_X1 U10186 ( .A1(n10046), .A2(n10060), .B1(n9749), .B2(n10052), .ZN(
        n10030) );
  INV_X1 U10187 ( .A(n10014), .ZN(n10064) );
  OR2_X1 U10188 ( .A1(n10130), .A2(n10064), .ZN(n9107) );
  NAND2_X1 U10189 ( .A1(n10130), .A2(n10064), .ZN(n9108) );
  OR2_X1 U10190 ( .A1(n10126), .A2(n10040), .ZN(n9109) );
  INV_X1 U10191 ( .A(n10016), .ZN(n9987) );
  NAND2_X1 U10192 ( .A1(n10120), .A2(n9987), .ZN(n9111) );
  NAND2_X1 U10193 ( .A1(n10114), .A2(n9997), .ZN(n9112) );
  NAND2_X1 U10194 ( .A1(n9976), .A2(n9112), .ZN(n9963) );
  OR2_X1 U10195 ( .A1(n10109), .A2(n9988), .ZN(n9113) );
  NAND2_X1 U10196 ( .A1(n9963), .A2(n9113), .ZN(n9115) );
  NAND2_X1 U10197 ( .A1(n10109), .A2(n9988), .ZN(n9114) );
  NAND2_X1 U10198 ( .A1(n10972), .A2(n9119), .ZN(n9121) );
  NAND2_X1 U10199 ( .A1(n9996), .A2(n10003), .ZN(n9995) );
  NAND2_X1 U10200 ( .A1(n9995), .A2(n9124), .ZN(n9985) );
  NAND2_X1 U10201 ( .A1(n9985), .A2(n9986), .ZN(n9984) );
  NAND2_X1 U10202 ( .A1(n9984), .A2(n9125), .ZN(n9969) );
  NAND2_X1 U10203 ( .A1(n9969), .A2(n9970), .ZN(n9968) );
  NAND2_X1 U10204 ( .A1(n9968), .A2(n9126), .ZN(n9951) );
  NAND2_X1 U10205 ( .A1(n9951), .A2(n9952), .ZN(n9950) );
  NAND2_X1 U10206 ( .A1(n9950), .A2(n9127), .ZN(n9940) );
  NAND2_X1 U10207 ( .A1(n9940), .A2(n9941), .ZN(n9939) );
  XNOR2_X1 U10208 ( .A(n9158), .B(n9130), .ZN(n9132) );
  OAI22_X1 U10209 ( .A1(n9133), .A2(n10015), .B1(n9809), .B2(n10013), .ZN(
        n9134) );
  INV_X1 U10210 ( .A(n9899), .ZN(n9137) );
  AOI21_X1 U10211 ( .B1(n10083), .B2(n9137), .A(n5317), .ZN(n10084) );
  AOI22_X1 U10212 ( .A1(n10738), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9138), 
        .B2(n10994), .ZN(n9139) );
  OAI21_X1 U10213 ( .B1(n9140), .B2(n10734), .A(n9139), .ZN(n9142) );
  NOR2_X1 U10214 ( .A1(n10087), .A2(n10029), .ZN(n9141) );
  OAI21_X1 U10215 ( .B1(n10086), .B2(n10738), .A(n9143), .ZN(P1_U3263) );
  INV_X1 U10216 ( .A(n9144), .ZN(n9147) );
  OAI222_X1 U10217 ( .A1(n5043), .A2(n9147), .B1(P2_U3152), .B2(n6366), .C1(
        n9146), .C2(n9698), .ZN(P2_U3330) );
  AOI21_X1 U10218 ( .B1(n10078), .B2(n9151), .A(n9892), .ZN(n10079) );
  INV_X1 U10219 ( .A(n10078), .ZN(n9154) );
  AOI22_X1 U10220 ( .A1(n10738), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9152), 
        .B2(n10994), .ZN(n9153) );
  OAI21_X1 U10221 ( .B1(n9154), .B2(n10734), .A(n9153), .ZN(n9161) );
  INV_X1 U10222 ( .A(n9155), .ZN(n9156) );
  OAI21_X1 U10223 ( .B1(n10082), .B2(n10070), .A(n9162), .ZN(P1_U3355) );
  XNOR2_X1 U10224 ( .A(n9163), .B(n9164), .ZN(n9171) );
  OAI22_X1 U10225 ( .A1(n9166), .A2(n9229), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9165), .ZN(n9169) );
  INV_X1 U10226 ( .A(n9388), .ZN(n9167) );
  OAI22_X1 U10227 ( .A1(n9167), .A2(n9259), .B1(n9198), .B2(n9230), .ZN(n9168)
         );
  AOI211_X1 U10228 ( .C1(n9597), .C2(n9261), .A(n9169), .B(n9168), .ZN(n9170)
         );
  OAI21_X1 U10229 ( .B1(n9171), .B2(n5042), .A(n9170), .ZN(P2_U3216) );
  INV_X1 U10230 ( .A(n9172), .ZN(n9173) );
  NAND3_X1 U10231 ( .A1(n9173), .A2(n9203), .A3(n9468), .ZN(n9177) );
  OAI22_X1 U10232 ( .A1(n9229), .A2(n9197), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10141), .ZN(n9175) );
  OAI22_X1 U10233 ( .A1(n9230), .A2(n9073), .B1(n9259), .B2(n9451), .ZN(n9174)
         );
  AOI211_X1 U10234 ( .C1(n9618), .C2(n9248), .A(n9175), .B(n9174), .ZN(n9176)
         );
  OAI211_X1 U10235 ( .C1(n9178), .C2(n5042), .A(n9177), .B(n9176), .ZN(
        P2_U3218) );
  OR3_X1 U10236 ( .A1(n9240), .A2(n9179), .A3(n9180), .ZN(n9188) );
  AOI22_X1 U10237 ( .A1(n9248), .A2(n6433), .B1(n9181), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n9187) );
  OAI21_X1 U10238 ( .B1(n9179), .B2(n9183), .A(n9182), .ZN(n9185) );
  AOI22_X1 U10239 ( .A1(n9220), .A2(n9185), .B1(n9257), .B2(n9184), .ZN(n9186)
         );
  NAND3_X1 U10240 ( .A1(n9188), .A2(n9187), .A3(n9186), .ZN(P2_U3224) );
  XNOR2_X1 U10241 ( .A(n9190), .B(n9189), .ZN(n9194) );
  OAI22_X1 U10242 ( .A1(n9229), .A2(n9073), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5141), .ZN(n9192) );
  OAI22_X1 U10243 ( .A1(n9230), .A2(n9510), .B1(n9259), .B2(n9479), .ZN(n9191)
         );
  AOI211_X1 U10244 ( .C1(n9629), .C2(n9261), .A(n9192), .B(n9191), .ZN(n9193)
         );
  OAI21_X1 U10245 ( .B1(n9194), .B2(n5042), .A(n9193), .ZN(P2_U3225) );
  XNOR2_X1 U10246 ( .A(n9196), .B(n9195), .ZN(n9202) );
  OAI22_X1 U10247 ( .A1(n9198), .A2(n9559), .B1(n9197), .B2(n9561), .ZN(n9422)
         );
  AOI22_X1 U10248 ( .A1(n9422), .A2(n9257), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n9199) );
  OAI21_X1 U10249 ( .B1(n9415), .B2(n9259), .A(n9199), .ZN(n9200) );
  AOI21_X1 U10250 ( .B1(n9608), .B2(n9261), .A(n9200), .ZN(n9201) );
  OAI21_X1 U10251 ( .B1(n9202), .B2(n5042), .A(n9201), .ZN(P2_U3227) );
  NAND2_X1 U10252 ( .A1(n9445), .A2(n9203), .ZN(n9207) );
  OR2_X1 U10253 ( .A1(n9204), .A2(n5042), .ZN(n9206) );
  MUX2_X1 U10254 ( .A(n9207), .B(n9206), .S(n9205), .Z(n9211) );
  AOI22_X1 U10255 ( .A1(n9247), .A2(n9468), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n9210) );
  AOI22_X1 U10256 ( .A1(n9078), .A2(n9244), .B1(n9246), .B2(n9430), .ZN(n9209)
         );
  NAND2_X1 U10257 ( .A1(n9612), .A2(n9248), .ZN(n9208) );
  NAND4_X1 U10258 ( .A1(n9211), .A2(n9210), .A3(n9209), .A4(n9208), .ZN(
        P2_U3231) );
  NOR3_X1 U10259 ( .A1(n9240), .A2(n9218), .A3(n9212), .ZN(n9213) );
  OAI21_X1 U10260 ( .B1(n9213), .B2(n9247), .A(n9280), .ZN(n9224) );
  AOI22_X1 U10261 ( .A1(n9248), .A2(n9214), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n9223) );
  AOI22_X1 U10262 ( .A1(n9244), .A2(n9279), .B1(n9246), .B2(n9215), .ZN(n9222)
         );
  OAI21_X1 U10263 ( .B1(n9218), .B2(n9217), .A(n9216), .ZN(n9219) );
  NAND2_X1 U10264 ( .A1(n9220), .A2(n9219), .ZN(n9221) );
  NAND4_X1 U10265 ( .A1(n9224), .A2(n9223), .A3(n9222), .A4(n9221), .ZN(
        P2_U3232) );
  INV_X1 U10266 ( .A(n9226), .ZN(n9227) );
  AOI21_X1 U10267 ( .B1(n9225), .B2(n9228), .A(n9227), .ZN(n9234) );
  OAI22_X1 U10268 ( .A1(n9229), .A2(n9436), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10233), .ZN(n9232) );
  OAI22_X1 U10269 ( .A1(n9230), .A2(n9266), .B1(n9259), .B2(n9462), .ZN(n9231)
         );
  AOI211_X1 U10270 ( .C1(n9624), .C2(n9248), .A(n9232), .B(n9231), .ZN(n9233)
         );
  OAI21_X1 U10271 ( .B1(n9234), .B2(n5042), .A(n9233), .ZN(P2_U3237) );
  INV_X1 U10272 ( .A(n9235), .ZN(n9236) );
  AOI21_X1 U10273 ( .B1(n9237), .B2(n9236), .A(n5042), .ZN(n9243) );
  NOR3_X1 U10274 ( .A1(n9240), .A2(n9239), .A3(n9238), .ZN(n9242) );
  OAI21_X1 U10275 ( .B1(n9243), .B2(n9242), .A(n9241), .ZN(n9252) );
  AOI22_X1 U10276 ( .A1(n9244), .A2(n9273), .B1(P2_REG3_REG_11__SCAN_IN), .B2(
        P2_U3152), .ZN(n9251) );
  AOI22_X1 U10277 ( .A1(n9247), .A2(n9275), .B1(n9246), .B2(n9245), .ZN(n9250)
         );
  NAND2_X1 U10278 ( .A1(n9248), .A2(n10901), .ZN(n9249) );
  NAND4_X1 U10279 ( .A1(n9252), .A2(n9251), .A3(n9250), .A4(n9249), .ZN(
        P2_U3238) );
  XNOR2_X1 U10280 ( .A(n9253), .B(n9254), .ZN(n9263) );
  OR2_X1 U10281 ( .A1(n9375), .A2(n9559), .ZN(n9256) );
  NAND2_X1 U10282 ( .A1(n9078), .A2(n10789), .ZN(n9255) );
  NAND2_X1 U10283 ( .A1(n9256), .A2(n9255), .ZN(n9403) );
  AOI22_X1 U10284 ( .A1(n9403), .A2(n9257), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n9258) );
  OAI21_X1 U10285 ( .B1(n9408), .B2(n9259), .A(n9258), .ZN(n9260) );
  AOI21_X1 U10286 ( .B1(n9603), .B2(n9261), .A(n9260), .ZN(n9262) );
  OAI21_X1 U10287 ( .B1(n9263), .B2(n5042), .A(n9262), .ZN(P2_U3242) );
  MUX2_X1 U10288 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n9360), .S(P2_U3966), .Z(
        P2_U3583) );
  MUX2_X1 U10289 ( .A(n9264), .B(P2_DATAO_REG_29__SCAN_IN), .S(n9267), .Z(
        P2_U3581) );
  MUX2_X1 U10290 ( .A(n9393), .B(P2_DATAO_REG_28__SCAN_IN), .S(n9267), .Z(
        P2_U3580) );
  MUX2_X1 U10291 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n9265), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U10292 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n9392), .S(P2_U3966), .Z(
        P2_U3578) );
  MUX2_X1 U10293 ( .A(n9078), .B(P2_DATAO_REG_25__SCAN_IN), .S(n9267), .Z(
        P2_U3577) );
  MUX2_X1 U10294 ( .A(n9445), .B(P2_DATAO_REG_24__SCAN_IN), .S(n9267), .Z(
        P2_U3576) );
  MUX2_X1 U10295 ( .A(n9468), .B(P2_DATAO_REG_23__SCAN_IN), .S(n9267), .Z(
        P2_U3575) );
  MUX2_X1 U10296 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9485), .S(P2_U3966), .Z(
        P2_U3574) );
  INV_X1 U10297 ( .A(n9266), .ZN(n9491) );
  MUX2_X1 U10298 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9491), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U10299 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9070), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U10300 ( .A(n9528), .B(P2_DATAO_REG_19__SCAN_IN), .S(n9267), .Z(
        P2_U3571) );
  MUX2_X1 U10301 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9268), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U10302 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9527), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U10303 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9269), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10304 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9270), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10305 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n9271), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U10306 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n9272), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U10307 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n9273), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U10308 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n9274), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U10309 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n9275), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U10310 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n9276), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U10311 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n9277), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U10312 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n9278), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U10313 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n10792), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U10314 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n9279), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U10315 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n10790), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U10316 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n9280), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U10317 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n9281), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U10318 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6436), .S(P2_U3966), .Z(
        P2_U3553) );
  OAI21_X1 U10319 ( .B1(n9283), .B2(n5072), .A(n9282), .ZN(n9284) );
  NAND2_X1 U10320 ( .A1(n10696), .A2(n9284), .ZN(n9293) );
  NAND2_X1 U10321 ( .A1(n10724), .A2(n9285), .ZN(n9292) );
  NOR2_X1 U10322 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10137), .ZN(n9286) );
  AOI21_X1 U10323 ( .B1(n10718), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n9286), .ZN(
        n9291) );
  OAI211_X1 U10324 ( .C1(n9289), .C2(n9288), .A(n10726), .B(n9287), .ZN(n9290)
         );
  NAND4_X1 U10325 ( .A1(n9293), .A2(n9292), .A3(n9291), .A4(n9290), .ZN(
        P2_U3256) );
  NAND2_X1 U10326 ( .A1(n9295), .A2(n9294), .ZN(n9297) );
  NAND2_X1 U10327 ( .A1(n9316), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n9298) );
  OAI21_X1 U10328 ( .B1(n9316), .B2(P2_REG2_REG_16__SCAN_IN), .A(n9298), .ZN(
        n9299) );
  AOI211_X1 U10329 ( .C1(n9300), .C2(n9299), .A(n9315), .B(n10719), .ZN(n9312)
         );
  NAND2_X1 U10330 ( .A1(n9302), .A2(n9301), .ZN(n9304) );
  NAND2_X1 U10331 ( .A1(n9304), .A2(n9303), .ZN(n9306) );
  XNOR2_X1 U10332 ( .A(n9316), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n9305) );
  NOR2_X1 U10333 ( .A1(n9306), .A2(n9305), .ZN(n9321) );
  AOI21_X1 U10334 ( .B1(n9306), .B2(n9305), .A(n9321), .ZN(n9307) );
  NOR2_X1 U10335 ( .A1(n9307), .A2(n9355), .ZN(n9311) );
  AND2_X1 U10336 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9308) );
  AOI21_X1 U10337 ( .B1(n10718), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n9308), .ZN(
        n9309) );
  OAI21_X1 U10338 ( .B1(n10710), .B2(n9323), .A(n9309), .ZN(n9310) );
  OR3_X1 U10339 ( .A1(n9312), .A2(n9311), .A3(n9310), .ZN(P2_U3261) );
  INV_X1 U10340 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9551) );
  OR2_X1 U10341 ( .A1(n9339), .A2(n9551), .ZN(n9314) );
  NAND2_X1 U10342 ( .A1(n9339), .A2(n9551), .ZN(n9313) );
  AND2_X1 U10343 ( .A1(n9314), .A2(n9313), .ZN(n9318) );
  NOR2_X1 U10344 ( .A1(n9317), .A2(n9318), .ZN(n9338) );
  AOI211_X1 U10345 ( .C1(n9318), .C2(n9317), .A(n9338), .B(n10719), .ZN(n9329)
         );
  NOR2_X1 U10346 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9319), .ZN(n9320) );
  AOI21_X1 U10347 ( .B1(n10718), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n9320), .ZN(
        n9327) );
  XNOR2_X1 U10348 ( .A(n9331), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n9325) );
  INV_X1 U10349 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9322) );
  AOI21_X1 U10350 ( .B1(n9323), .B2(n9322), .A(n9321), .ZN(n9324) );
  NAND2_X1 U10351 ( .A1(n9325), .A2(n9324), .ZN(n9330) );
  OAI211_X1 U10352 ( .C1(n9325), .C2(n9324), .A(n10726), .B(n9330), .ZN(n9326)
         );
  OAI211_X1 U10353 ( .C1(n10710), .C2(n9331), .A(n9327), .B(n9326), .ZN(n9328)
         );
  OR2_X1 U10354 ( .A1(n9329), .A2(n9328), .ZN(P2_U3262) );
  INV_X1 U10355 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9332) );
  OAI21_X1 U10356 ( .B1(n9332), .B2(n9331), .A(n9330), .ZN(n9348) );
  XNOR2_X1 U10357 ( .A(n9347), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n9349) );
  XOR2_X1 U10358 ( .A(n9348), .B(n9349), .Z(n9333) );
  NOR2_X1 U10359 ( .A1(n9355), .A2(n9333), .ZN(n9334) );
  AOI211_X1 U10360 ( .C1(n10718), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n9335), .B(
        n9334), .ZN(n9344) );
  OR2_X1 U10361 ( .A1(n9347), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9337) );
  NAND2_X1 U10362 ( .A1(n9347), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9336) );
  AND2_X1 U10363 ( .A1(n9337), .A2(n9336), .ZN(n9341) );
  AOI21_X1 U10364 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n9339), .A(n9338), .ZN(
        n9340) );
  OAI21_X1 U10365 ( .B1(n9341), .B2(n9340), .A(n9345), .ZN(n9342) );
  NAND2_X1 U10366 ( .A1(n10696), .A2(n9342), .ZN(n9343) );
  OAI211_X1 U10367 ( .C1(n10710), .C2(n5153), .A(n9344), .B(n9343), .ZN(
        P2_U3263) );
  MUX2_X1 U10368 ( .A(n6108), .B(P2_REG2_REG_19__SCAN_IN), .S(n9546), .Z(n9346) );
  OAI22_X1 U10369 ( .A1(n9349), .A2(n9348), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n9347), .ZN(n9351) );
  XNOR2_X1 U10370 ( .A(n10800), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n9350) );
  XNOR2_X1 U10371 ( .A(n9351), .B(n9350), .ZN(n9354) );
  NAND2_X1 U10372 ( .A1(n10718), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n9352) );
  OAI211_X1 U10373 ( .C1(n9355), .C2(n9354), .A(n9353), .B(n9352), .ZN(n9356)
         );
  AOI21_X1 U10374 ( .B1(n10800), .B2(n10724), .A(n9356), .ZN(n9357) );
  INV_X1 U10375 ( .A(n9358), .ZN(n9359) );
  AND2_X1 U10376 ( .A1(n9360), .A2(n9359), .ZN(n9579) );
  INV_X1 U10377 ( .A(n9579), .ZN(n9584) );
  NOR2_X1 U10378 ( .A1(n7664), .A2(n9584), .ZN(n9367) );
  AOI211_X1 U10379 ( .C1(n7664), .C2(P2_REG2_REG_31__SCAN_IN), .A(n9367), .B(
        n9361), .ZN(n9362) );
  OAI21_X1 U10380 ( .B1(n9363), .B2(n9578), .A(n9362), .ZN(P2_U3265) );
  INV_X1 U10381 ( .A(n9364), .ZN(n9366) );
  NAND2_X1 U10382 ( .A1(n9366), .A2(n9365), .ZN(n9583) );
  NAND3_X1 U10383 ( .A1(n9583), .A2(n9568), .A3(n9582), .ZN(n9369) );
  AOI21_X1 U10384 ( .B1(n7664), .B2(P2_REG2_REG_30__SCAN_IN), .A(n9367), .ZN(
        n9368) );
  OAI211_X1 U10385 ( .C1(n9586), .C2(n9547), .A(n9369), .B(n9368), .ZN(
        P2_U3266) );
  AOI21_X1 U10386 ( .B1(n9372), .B2(n9371), .A(n9370), .ZN(n9373) );
  OAI222_X1 U10387 ( .A1(n9561), .A2(n9375), .B1(n9559), .B2(n9374), .C1(n9538), .C2(n9373), .ZN(n9591) );
  INV_X1 U10388 ( .A(n9592), .ZN(n9381) );
  INV_X1 U10389 ( .A(n9376), .ZN(n9377) );
  AOI21_X1 U10390 ( .B1(n9592), .B2(n9385), .A(n9377), .ZN(n9593) );
  NAND2_X1 U10391 ( .A1(n9593), .A2(n9568), .ZN(n9380) );
  AOI22_X1 U10392 ( .A1(n9378), .A2(n10798), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n7664), .ZN(n9379) );
  OAI211_X1 U10393 ( .C1(n9381), .C2(n9547), .A(n9380), .B(n9379), .ZN(n9382)
         );
  AOI21_X1 U10394 ( .B1(n9591), .B2(n10803), .A(n9382), .ZN(n9383) );
  OAI21_X1 U10395 ( .B1(n9596), .B2(n9533), .A(n9383), .ZN(P2_U3268) );
  XNOR2_X1 U10396 ( .A(n9384), .B(n5143), .ZN(n9601) );
  INV_X1 U10397 ( .A(n9405), .ZN(n9387) );
  INV_X1 U10398 ( .A(n9385), .ZN(n9386) );
  AOI21_X1 U10399 ( .B1(n9597), .B2(n9387), .A(n9386), .ZN(n9598) );
  AOI22_X1 U10400 ( .A1(n9388), .A2(n10798), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n7664), .ZN(n9389) );
  OAI21_X1 U10401 ( .B1(n9390), .B2(n9547), .A(n9389), .ZN(n9396) );
  XNOR2_X1 U10402 ( .A(n9391), .B(n5143), .ZN(n9394) );
  AOI222_X1 U10403 ( .A1(n10794), .A2(n9394), .B1(n9393), .B2(n10791), .C1(
        n9392), .C2(n10789), .ZN(n9600) );
  NOR2_X1 U10404 ( .A1(n9600), .A2(n7664), .ZN(n9395) );
  AOI211_X1 U10405 ( .C1(n9568), .C2(n9598), .A(n9396), .B(n9395), .ZN(n9397)
         );
  OAI21_X1 U10406 ( .B1(n9601), .B2(n9533), .A(n9397), .ZN(P2_U3269) );
  XOR2_X1 U10407 ( .A(n9401), .B(n9398), .Z(n9606) );
  AOI22_X1 U10408 ( .A1(n9603), .A2(n9573), .B1(n7664), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n9411) );
  INV_X1 U10409 ( .A(n9399), .ZN(n9400) );
  NOR2_X1 U10410 ( .A1(n9419), .A2(n9400), .ZN(n9402) );
  XNOR2_X1 U10411 ( .A(n9402), .B(n9401), .ZN(n9404) );
  AOI21_X1 U10412 ( .B1(n9404), .B2(n10794), .A(n9403), .ZN(n9605) );
  INV_X1 U10413 ( .A(n9413), .ZN(n9406) );
  AOI211_X1 U10414 ( .C1(n9603), .C2(n9406), .A(n10921), .B(n9405), .ZN(n9602)
         );
  NAND2_X1 U10415 ( .A1(n9602), .A2(n9546), .ZN(n9407) );
  OAI211_X1 U10416 ( .C1(n9549), .C2(n9408), .A(n9605), .B(n9407), .ZN(n9409)
         );
  NAND2_X1 U10417 ( .A1(n9409), .A2(n10803), .ZN(n9410) );
  OAI211_X1 U10418 ( .C1(n9606), .C2(n9533), .A(n9411), .B(n9410), .ZN(
        P2_U3270) );
  XOR2_X1 U10419 ( .A(n9420), .B(n9412), .Z(n9611) );
  AOI21_X1 U10420 ( .B1(n9432), .B2(n9449), .A(n9418), .ZN(n9414) );
  NOR3_X1 U10421 ( .A1(n9414), .A2(n9413), .A3(n10921), .ZN(n9607) );
  INV_X1 U10422 ( .A(n9415), .ZN(n9416) );
  AOI22_X1 U10423 ( .A1(n9416), .A2(n10798), .B1(n7664), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n9417) );
  OAI21_X1 U10424 ( .B1(n9418), .B2(n9547), .A(n9417), .ZN(n9425) );
  AOI211_X1 U10425 ( .C1(n9421), .C2(n9420), .A(n9538), .B(n9419), .ZN(n9423)
         );
  NOR2_X1 U10426 ( .A1(n9423), .A2(n9422), .ZN(n9610) );
  NOR2_X1 U10427 ( .A1(n9610), .A2(n7664), .ZN(n9424) );
  AOI211_X1 U10428 ( .C1(n9607), .C2(n9426), .A(n9425), .B(n9424), .ZN(n9427)
         );
  OAI21_X1 U10429 ( .B1(n9611), .B2(n9533), .A(n9427), .ZN(P2_U3271) );
  OAI21_X1 U10430 ( .B1(n5077), .B2(n9435), .A(n9428), .ZN(n9429) );
  INV_X1 U10431 ( .A(n9429), .ZN(n9616) );
  XNOR2_X1 U10432 ( .A(n9449), .B(n9612), .ZN(n9613) );
  AOI22_X1 U10433 ( .A1(n7664), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n9430), .B2(
        n10798), .ZN(n9431) );
  OAI21_X1 U10434 ( .B1(n9432), .B2(n9547), .A(n9431), .ZN(n9441) );
  AOI211_X1 U10435 ( .C1(n9435), .C2(n9434), .A(n9538), .B(n9433), .ZN(n9439)
         );
  OAI22_X1 U10436 ( .A1(n9437), .A2(n9559), .B1(n9436), .B2(n9561), .ZN(n9438)
         );
  NOR2_X1 U10437 ( .A1(n9439), .A2(n9438), .ZN(n9615) );
  NOR2_X1 U10438 ( .A1(n9615), .A2(n7664), .ZN(n9440) );
  AOI211_X1 U10439 ( .C1(n9613), .C2(n9568), .A(n9441), .B(n9440), .ZN(n9442)
         );
  OAI21_X1 U10440 ( .B1(n9616), .B2(n9533), .A(n9442), .ZN(P2_U3272) );
  XNOR2_X1 U10441 ( .A(n9444), .B(n9443), .ZN(n9446) );
  AOI222_X1 U10442 ( .A1(n10794), .A2(n9446), .B1(n9485), .B2(n10789), .C1(
        n9445), .C2(n10791), .ZN(n9621) );
  NAND2_X1 U10443 ( .A1(n9448), .A2(n9447), .ZN(n9617) );
  NAND3_X1 U10444 ( .A1(n5614), .A2(n9572), .A3(n9617), .ZN(n9457) );
  INV_X1 U10445 ( .A(n9461), .ZN(n9450) );
  AOI21_X1 U10446 ( .B1(n9618), .B2(n9450), .A(n9449), .ZN(n9619) );
  INV_X1 U10447 ( .A(n9451), .ZN(n9452) );
  AOI22_X1 U10448 ( .A1(n7664), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n9452), .B2(
        n10798), .ZN(n9453) );
  OAI21_X1 U10449 ( .B1(n9454), .B2(n9547), .A(n9453), .ZN(n9455) );
  AOI21_X1 U10450 ( .B1(n9619), .B2(n9568), .A(n9455), .ZN(n9456) );
  OAI211_X1 U10451 ( .C1(n7664), .C2(n9621), .A(n9457), .B(n9456), .ZN(
        P2_U3273) );
  INV_X1 U10452 ( .A(n9458), .ZN(n9459) );
  AOI21_X1 U10453 ( .B1(n9466), .B2(n9460), .A(n9459), .ZN(n9628) );
  AOI21_X1 U10454 ( .B1(n9624), .B2(n9477), .A(n9461), .ZN(n9625) );
  INV_X1 U10455 ( .A(n9462), .ZN(n9463) );
  AOI22_X1 U10456 ( .A1(n7664), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9463), .B2(
        n10798), .ZN(n9464) );
  OAI21_X1 U10457 ( .B1(n9074), .B2(n9547), .A(n9464), .ZN(n9472) );
  OAI211_X1 U10458 ( .C1(n9467), .C2(n9466), .A(n9465), .B(n10794), .ZN(n9470)
         );
  AOI22_X1 U10459 ( .A1(n9468), .A2(n10791), .B1(n10789), .B2(n9491), .ZN(
        n9469) );
  AND2_X1 U10460 ( .A1(n9470), .A2(n9469), .ZN(n9627) );
  NOR2_X1 U10461 ( .A1(n9627), .A2(n7664), .ZN(n9471) );
  AOI211_X1 U10462 ( .C1(n9625), .C2(n9568), .A(n9472), .B(n9471), .ZN(n9473)
         );
  OAI21_X1 U10463 ( .B1(n9628), .B2(n9533), .A(n9473), .ZN(P2_U3274) );
  OAI21_X1 U10464 ( .B1(n9476), .B2(n9475), .A(n9474), .ZN(n9633) );
  INV_X1 U10465 ( .A(n9477), .ZN(n9478) );
  AOI21_X1 U10466 ( .B1(n9629), .B2(n9498), .A(n9478), .ZN(n9630) );
  INV_X1 U10467 ( .A(n9479), .ZN(n9480) );
  AOI22_X1 U10468 ( .A1(n7664), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9480), .B2(
        n10798), .ZN(n9481) );
  OAI21_X1 U10469 ( .B1(n9482), .B2(n9547), .A(n9481), .ZN(n9488) );
  XNOR2_X1 U10470 ( .A(n9484), .B(n9483), .ZN(n9486) );
  AOI222_X1 U10471 ( .A1(n10794), .A2(n9486), .B1(n9485), .B2(n10791), .C1(
        n9070), .C2(n10789), .ZN(n9632) );
  NOR2_X1 U10472 ( .A1(n9632), .A2(n7664), .ZN(n9487) );
  AOI211_X1 U10473 ( .C1(n9630), .C2(n9568), .A(n9488), .B(n9487), .ZN(n9489)
         );
  OAI21_X1 U10474 ( .B1(n9533), .B2(n9633), .A(n9489), .ZN(P2_U3275) );
  XNOR2_X1 U10475 ( .A(n9490), .B(n9495), .ZN(n9492) );
  AOI222_X1 U10476 ( .A1(n10794), .A2(n9492), .B1(n9491), .B2(n10791), .C1(
        n9528), .C2(n10789), .ZN(n9637) );
  OAI21_X1 U10477 ( .B1(n9493), .B2(n9549), .A(n9637), .ZN(n9503) );
  OAI21_X1 U10478 ( .B1(n9496), .B2(n9495), .A(n9494), .ZN(n9638) );
  AOI22_X1 U10479 ( .A1(n9634), .A2(n9573), .B1(n7664), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n9501) );
  OR2_X1 U10480 ( .A1(n9497), .A2(n9511), .ZN(n9499) );
  AND2_X1 U10481 ( .A1(n9499), .A2(n9498), .ZN(n9635) );
  NAND2_X1 U10482 ( .A1(n9635), .A2(n9568), .ZN(n9500) );
  OAI211_X1 U10483 ( .C1(n9638), .C2(n9533), .A(n9501), .B(n9500), .ZN(n9502)
         );
  AOI21_X1 U10484 ( .B1(n10803), .B2(n9503), .A(n9502), .ZN(n9504) );
  INV_X1 U10485 ( .A(n9504), .ZN(P2_U3276) );
  OAI21_X1 U10486 ( .B1(n9506), .B2(n9507), .A(n9505), .ZN(n9643) );
  AOI22_X1 U10487 ( .A1(n9641), .A2(n9573), .B1(P2_REG2_REG_19__SCAN_IN), .B2(
        n7664), .ZN(n9516) );
  XNOR2_X1 U10488 ( .A(n9508), .B(n9507), .ZN(n9509) );
  OAI222_X1 U10489 ( .A1(n9559), .A2(n9510), .B1(n9561), .B2(n9539), .C1(n9509), .C2(n9538), .ZN(n9639) );
  AOI211_X1 U10490 ( .C1(n9641), .C2(n9519), .A(n10921), .B(n9511), .ZN(n9640)
         );
  INV_X1 U10491 ( .A(n9640), .ZN(n9513) );
  OAI22_X1 U10492 ( .A1(n9513), .A2(n10800), .B1(n9549), .B2(n9512), .ZN(n9514) );
  OAI21_X1 U10493 ( .B1(n9639), .B2(n9514), .A(n10803), .ZN(n9515) );
  OAI211_X1 U10494 ( .C1(n9643), .C2(n9533), .A(n9516), .B(n9515), .ZN(
        P2_U3277) );
  XNOR2_X1 U10495 ( .A(n9518), .B(n9517), .ZN(n9648) );
  INV_X1 U10496 ( .A(n9519), .ZN(n9520) );
  AOI21_X1 U10497 ( .B1(n9644), .B2(n9521), .A(n9520), .ZN(n9645) );
  AOI22_X1 U10498 ( .A1(n7664), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9522), .B2(
        n10798), .ZN(n9523) );
  OAI21_X1 U10499 ( .B1(n9524), .B2(n9547), .A(n9523), .ZN(n9531) );
  XNOR2_X1 U10500 ( .A(n9526), .B(n9525), .ZN(n9529) );
  AOI222_X1 U10501 ( .A1(n10794), .A2(n9529), .B1(n9528), .B2(n10791), .C1(
        n9527), .C2(n10789), .ZN(n9647) );
  NOR2_X1 U10502 ( .A1(n9647), .A2(n7664), .ZN(n9530) );
  AOI211_X1 U10503 ( .C1(n9645), .C2(n9568), .A(n9531), .B(n9530), .ZN(n9532)
         );
  OAI21_X1 U10504 ( .B1(n9533), .B2(n9648), .A(n9532), .ZN(P2_U3278) );
  XNOR2_X1 U10505 ( .A(n9548), .B(n9534), .ZN(n9535) );
  NOR2_X1 U10506 ( .A1(n9535), .A2(n10921), .ZN(n9650) );
  XNOR2_X1 U10507 ( .A(n9536), .B(n9542), .ZN(n9537) );
  OAI222_X1 U10508 ( .A1(n9561), .A2(n9540), .B1(n9559), .B2(n9539), .C1(n9538), .C2(n9537), .ZN(n9649) );
  OAI21_X1 U10509 ( .B1(n9543), .B2(n9542), .A(n9541), .ZN(n9555) );
  INV_X1 U10510 ( .A(n9555), .ZN(n9653) );
  NOR2_X1 U10511 ( .A1(n9653), .A2(n9544), .ZN(n9545) );
  AOI211_X1 U10512 ( .C1(n9650), .C2(n9546), .A(n9649), .B(n9545), .ZN(n9557)
         );
  NOR2_X1 U10513 ( .A1(n9548), .A2(n9547), .ZN(n9553) );
  OAI22_X1 U10514 ( .A1(n10803), .A2(n9551), .B1(n9550), .B2(n9549), .ZN(n9552) );
  AOI211_X1 U10515 ( .C1(n9555), .C2(n9554), .A(n9553), .B(n9552), .ZN(n9556)
         );
  OAI21_X1 U10516 ( .B1(n9557), .B2(n7664), .A(n9556), .ZN(P2_U3279) );
  XNOR2_X1 U10517 ( .A(n9558), .B(n9571), .ZN(n9564) );
  OAI22_X1 U10518 ( .A1(n9562), .A2(n9561), .B1(n9560), .B2(n9559), .ZN(n9563)
         );
  AOI21_X1 U10519 ( .B1(n9564), .B2(n10794), .A(n9563), .ZN(n10826) );
  MUX2_X1 U10520 ( .A(n6986), .B(n10826), .S(n10803), .Z(n9577) );
  INV_X1 U10521 ( .A(n10786), .ZN(n9566) );
  AOI21_X1 U10522 ( .B1(n10821), .B2(n9566), .A(n9565), .ZN(n10822) );
  AOI22_X1 U10523 ( .A1(n9568), .A2(n10822), .B1(n9567), .B2(n10798), .ZN(
        n9576) );
  NAND2_X1 U10524 ( .A1(n9570), .A2(n9571), .ZN(n10823) );
  NAND3_X1 U10525 ( .A1(n9569), .A2(n10823), .A3(n9572), .ZN(n9575) );
  NAND2_X1 U10526 ( .A1(n9573), .A2(n10821), .ZN(n9574) );
  NAND4_X1 U10527 ( .A1(n9577), .A2(n9576), .A3(n9575), .A4(n9574), .ZN(
        P2_U3290) );
  AOI21_X1 U10528 ( .B1(n9580), .B2(n10939), .A(n9579), .ZN(n9581) );
  INV_X2 U10529 ( .A(n10945), .ZN(n10811) );
  MUX2_X1 U10530 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9669), .S(n10811), .Z(
        P2_U3551) );
  NAND3_X1 U10531 ( .A1(n9583), .A2(n10940), .A3(n9582), .ZN(n9585) );
  OAI211_X1 U10532 ( .C1(n9586), .C2(n10919), .A(n9585), .B(n9584), .ZN(n9670)
         );
  MUX2_X1 U10533 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9670), .S(n10811), .Z(
        P2_U3550) );
  AOI22_X1 U10534 ( .A1(n9587), .A2(n10940), .B1(n10939), .B2(n9083), .ZN(
        n9588) );
  MUX2_X1 U10535 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9671), .S(n10811), .Z(
        P2_U3549) );
  INV_X1 U10536 ( .A(n9591), .ZN(n9595) );
  AOI22_X1 U10537 ( .A1(n9593), .A2(n10940), .B1(n10939), .B2(n9592), .ZN(
        n9594) );
  MUX2_X1 U10538 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9672), .S(n10811), .Z(
        P2_U3548) );
  AOI22_X1 U10539 ( .A1(n9598), .A2(n10940), .B1(n10939), .B2(n9597), .ZN(
        n9599) );
  OAI211_X1 U10540 ( .C1(n9601), .C2(n10904), .A(n9600), .B(n9599), .ZN(n9673)
         );
  MUX2_X1 U10541 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9673), .S(n10811), .Z(
        P2_U3547) );
  AOI21_X1 U10542 ( .B1(n10939), .B2(n9603), .A(n9602), .ZN(n9604) );
  OAI211_X1 U10543 ( .C1(n9606), .C2(n10904), .A(n9605), .B(n9604), .ZN(n9674)
         );
  MUX2_X1 U10544 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9674), .S(n10811), .Z(
        P2_U3546) );
  AOI21_X1 U10545 ( .B1(n10939), .B2(n9608), .A(n9607), .ZN(n9609) );
  OAI211_X1 U10546 ( .C1(n9611), .C2(n10904), .A(n9610), .B(n9609), .ZN(n9675)
         );
  MUX2_X1 U10547 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9675), .S(n10811), .Z(
        P2_U3545) );
  AOI22_X1 U10548 ( .A1(n9613), .A2(n10940), .B1(n10939), .B2(n9612), .ZN(
        n9614) );
  OAI211_X1 U10549 ( .C1(n9616), .C2(n10904), .A(n9615), .B(n9614), .ZN(n9676)
         );
  MUX2_X1 U10550 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9676), .S(n10811), .Z(
        P2_U3544) );
  NAND2_X1 U10551 ( .A1(n9617), .A2(n10936), .ZN(n9622) );
  AOI22_X1 U10552 ( .A1(n9619), .A2(n10940), .B1(n10939), .B2(n9618), .ZN(
        n9620) );
  OAI211_X1 U10553 ( .C1(n9623), .C2(n9622), .A(n9621), .B(n9620), .ZN(n9677)
         );
  MUX2_X1 U10554 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9677), .S(n10811), .Z(
        P2_U3543) );
  AOI22_X1 U10555 ( .A1(n9625), .A2(n10940), .B1(n10939), .B2(n9624), .ZN(
        n9626) );
  OAI211_X1 U10556 ( .C1(n9628), .C2(n10904), .A(n9627), .B(n9626), .ZN(n9678)
         );
  MUX2_X1 U10557 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9678), .S(n10811), .Z(
        P2_U3542) );
  AOI22_X1 U10558 ( .A1(n9630), .A2(n10940), .B1(n10939), .B2(n9629), .ZN(
        n9631) );
  OAI211_X1 U10559 ( .C1(n9633), .C2(n10904), .A(n9632), .B(n9631), .ZN(n9679)
         );
  MUX2_X1 U10560 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9679), .S(n10811), .Z(
        P2_U3541) );
  AOI22_X1 U10561 ( .A1(n9635), .A2(n10940), .B1(n10939), .B2(n9634), .ZN(
        n9636) );
  OAI211_X1 U10562 ( .C1(n9638), .C2(n10904), .A(n9637), .B(n9636), .ZN(n9680)
         );
  MUX2_X1 U10563 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9680), .S(n10811), .Z(
        P2_U3540) );
  AOI211_X1 U10564 ( .C1(n10939), .C2(n9641), .A(n9640), .B(n9639), .ZN(n9642)
         );
  OAI21_X1 U10565 ( .B1(n9643), .B2(n10904), .A(n9642), .ZN(n9681) );
  MUX2_X1 U10566 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9681), .S(n10811), .Z(
        P2_U3539) );
  AOI22_X1 U10567 ( .A1(n9645), .A2(n10940), .B1(n10939), .B2(n9644), .ZN(
        n9646) );
  OAI211_X1 U10568 ( .C1(n9648), .C2(n10904), .A(n9647), .B(n9646), .ZN(n9682)
         );
  MUX2_X1 U10569 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9682), .S(n10811), .Z(
        P2_U3538) );
  AOI211_X1 U10570 ( .C1(n10939), .C2(n9651), .A(n9650), .B(n9649), .ZN(n9652)
         );
  OAI21_X1 U10571 ( .B1(n9653), .B2(n10904), .A(n9652), .ZN(n9683) );
  MUX2_X1 U10572 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9683), .S(n10811), .Z(
        P2_U3537) );
  AOI21_X1 U10573 ( .B1(n10939), .B2(n9655), .A(n9654), .ZN(n9656) );
  OAI211_X1 U10574 ( .C1(n9658), .C2(n10904), .A(n9657), .B(n9656), .ZN(n9684)
         );
  MUX2_X1 U10575 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9684), .S(n10811), .Z(
        P2_U3536) );
  AOI22_X1 U10576 ( .A1(n9660), .A2(n10940), .B1(n10939), .B2(n9659), .ZN(
        n9661) );
  OAI211_X1 U10577 ( .C1(n9663), .C2(n10904), .A(n9662), .B(n9661), .ZN(n9685)
         );
  MUX2_X1 U10578 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9685), .S(n10811), .Z(
        P2_U3535) );
  AOI22_X1 U10579 ( .A1(n9665), .A2(n10940), .B1(n10939), .B2(n9664), .ZN(
        n9666) );
  OAI211_X1 U10580 ( .C1(n9668), .C2(n10904), .A(n9667), .B(n9666), .ZN(n9686)
         );
  MUX2_X1 U10581 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n9686), .S(n10811), .Z(
        P2_U3534) );
  MUX2_X1 U10582 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9669), .S(n10950), .Z(
        P2_U3519) );
  MUX2_X1 U10583 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9670), .S(n10950), .Z(
        P2_U3518) );
  MUX2_X1 U10584 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9671), .S(n10950), .Z(
        P2_U3517) );
  MUX2_X1 U10585 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9672), .S(n10950), .Z(
        P2_U3516) );
  MUX2_X1 U10586 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9673), .S(n10950), .Z(
        P2_U3515) );
  MUX2_X1 U10587 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9674), .S(n10950), .Z(
        P2_U3514) );
  MUX2_X1 U10588 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9675), .S(n10950), .Z(
        P2_U3513) );
  MUX2_X1 U10589 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9676), .S(n10950), .Z(
        P2_U3512) );
  MUX2_X1 U10590 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9677), .S(n10950), .Z(
        P2_U3511) );
  MUX2_X1 U10591 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9678), .S(n10950), .Z(
        P2_U3510) );
  MUX2_X1 U10592 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9679), .S(n10950), .Z(
        P2_U3509) );
  MUX2_X1 U10593 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9680), .S(n10950), .Z(
        P2_U3508) );
  MUX2_X1 U10594 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9681), .S(n10950), .Z(
        P2_U3507) );
  MUX2_X1 U10595 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9682), .S(n10950), .Z(
        P2_U3505) );
  MUX2_X1 U10596 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9683), .S(n10950), .Z(
        P2_U3502) );
  MUX2_X1 U10597 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9684), .S(n10950), .Z(
        P2_U3499) );
  MUX2_X1 U10598 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9685), .S(n10950), .Z(
        P2_U3496) );
  MUX2_X1 U10599 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n9686), .S(n10950), .Z(
        P2_U3493) );
  INV_X1 U10600 ( .A(n9687), .ZN(n10566) );
  INV_X1 U10601 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9688) );
  NAND3_X1 U10602 ( .A1(n9688), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n9690) );
  OAI22_X1 U10603 ( .A1(n5688), .A2(n9690), .B1(n9689), .B2(n9698), .ZN(n9691)
         );
  INV_X1 U10604 ( .A(n9691), .ZN(n9692) );
  OAI21_X1 U10605 ( .B1(n10566), .B2(n5043), .A(n9692), .ZN(P2_U3327) );
  INV_X1 U10606 ( .A(n9693), .ZN(n10569) );
  OAI222_X1 U10607 ( .A1(n5043), .A2(n10569), .B1(P2_U3152), .B2(n9695), .C1(
        n9696), .C2(n9698), .ZN(P2_U3328) );
  INV_X1 U10608 ( .A(n9697), .ZN(n10577) );
  OAI222_X1 U10609 ( .A1(P2_U3152), .A2(n9700), .B1(n5043), .B2(n10577), .C1(
        n9699), .C2(n9698), .ZN(P2_U3332) );
  MUX2_X1 U10610 ( .A(n9701), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10611 ( .A(n9702), .ZN(n9704) );
  NAND2_X1 U10612 ( .A1(n9704), .A2(n9703), .ZN(n9706) );
  XNOR2_X1 U10613 ( .A(n9706), .B(n9705), .ZN(n9712) );
  NAND2_X1 U10614 ( .A1(n9804), .A2(n9966), .ZN(n9708) );
  AOI22_X1 U10615 ( .A1(n9805), .A2(n9997), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9707) );
  OAI211_X1 U10616 ( .C1(n9709), .C2(n9808), .A(n9708), .B(n9707), .ZN(n9710)
         );
  AOI21_X1 U10617 ( .B1(n10109), .B2(n9811), .A(n9710), .ZN(n9711) );
  OAI21_X1 U10618 ( .B1(n9712), .B2(n9813), .A(n9711), .ZN(P1_U3214) );
  INV_X1 U10619 ( .A(n9713), .ZN(n9716) );
  AOI21_X1 U10620 ( .B1(n9790), .B2(n9787), .A(n9714), .ZN(n9715) );
  OAI21_X1 U10621 ( .B1(n9716), .B2(n9715), .A(n9744), .ZN(n9720) );
  NAND2_X1 U10622 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9886) );
  OAI21_X1 U10623 ( .B1(n9794), .B2(n9749), .A(n9886), .ZN(n9718) );
  NOR2_X1 U10624 ( .A1(n9795), .A2(n10034), .ZN(n9717) );
  AOI211_X1 U10625 ( .C1(n9798), .C2(n10040), .A(n9718), .B(n9717), .ZN(n9719)
         );
  OAI211_X1 U10626 ( .C1(n10037), .C2(n9801), .A(n9720), .B(n9719), .ZN(
        P1_U3217) );
  INV_X1 U10627 ( .A(n9721), .ZN(n9722) );
  NOR2_X1 U10628 ( .A1(n9723), .A2(n9722), .ZN(n9724) );
  XNOR2_X1 U10629 ( .A(n9725), .B(n9724), .ZN(n9731) );
  NAND2_X1 U10630 ( .A1(n9804), .A2(n10001), .ZN(n9727) );
  AOI22_X1 U10631 ( .A1(n10040), .A2(n9805), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9726) );
  OAI211_X1 U10632 ( .C1(n9728), .C2(n9808), .A(n9727), .B(n9726), .ZN(n9729)
         );
  AOI21_X1 U10633 ( .B1(n10120), .B2(n9811), .A(n9729), .ZN(n9730) );
  OAI21_X1 U10634 ( .B1(n9731), .B2(n9813), .A(n9730), .ZN(P1_U3221) );
  XNOR2_X1 U10635 ( .A(n9733), .B(n9732), .ZN(n9734) );
  XNOR2_X1 U10636 ( .A(n9735), .B(n9734), .ZN(n9741) );
  NAND2_X1 U10637 ( .A1(n9804), .A2(n9936), .ZN(n9737) );
  AOI22_X1 U10638 ( .A1(n9805), .A2(n9971), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9736) );
  OAI211_X1 U10639 ( .C1(n9738), .C2(n9808), .A(n9737), .B(n9736), .ZN(n9739)
         );
  AOI21_X1 U10640 ( .B1(n10099), .B2(n9811), .A(n9739), .ZN(n9740) );
  OAI21_X1 U10641 ( .B1(n9741), .B2(n9813), .A(n9740), .ZN(P1_U3223) );
  NOR3_X1 U10642 ( .A1(n5111), .A2(n5514), .A3(n9743), .ZN(n9745) );
  OAI21_X1 U10643 ( .B1(n9745), .B2(n5114), .A(n9744), .ZN(n9753) );
  INV_X1 U10644 ( .A(n9746), .ZN(n9747) );
  AOI21_X1 U10645 ( .B1(n9805), .B2(n9817), .A(n9747), .ZN(n9748) );
  OAI21_X1 U10646 ( .B1(n9749), .B2(n9808), .A(n9748), .ZN(n9750) );
  AOI21_X1 U10647 ( .B1(n9804), .B2(n9751), .A(n9750), .ZN(n9752) );
  OAI211_X1 U10648 ( .C1(n9754), .C2(n9801), .A(n9753), .B(n9752), .ZN(
        P1_U3226) );
  XOR2_X1 U10649 ( .A(n9756), .B(n9755), .Z(n9762) );
  NAND2_X1 U10650 ( .A1(n9804), .A2(n9957), .ZN(n9758) );
  AOI22_X1 U10651 ( .A1(n9805), .A2(n9988), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9757) );
  OAI211_X1 U10652 ( .C1(n9759), .C2(n9808), .A(n9758), .B(n9757), .ZN(n9760)
         );
  AOI21_X1 U10653 ( .B1(n10105), .B2(n9811), .A(n9760), .ZN(n9761) );
  OAI21_X1 U10654 ( .B1(n9762), .B2(n9813), .A(n9761), .ZN(P1_U3227) );
  INV_X1 U10655 ( .A(n9763), .ZN(n9765) );
  NAND2_X1 U10656 ( .A1(n9765), .A2(n9764), .ZN(n9766) );
  XNOR2_X1 U10657 ( .A(n9767), .B(n9766), .ZN(n9773) );
  INV_X1 U10658 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9768) );
  OAI22_X1 U10659 ( .A1(n10014), .A2(n9794), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9768), .ZN(n9769) );
  AOI21_X1 U10660 ( .B1(n9987), .B2(n9798), .A(n9769), .ZN(n9770) );
  OAI21_X1 U10661 ( .B1(n9795), .B2(n10025), .A(n9770), .ZN(n9771) );
  AOI21_X1 U10662 ( .B1(n10126), .B2(n9811), .A(n9771), .ZN(n9772) );
  OAI21_X1 U10663 ( .B1(n9773), .B2(n9813), .A(n9772), .ZN(P1_U3231) );
  INV_X1 U10664 ( .A(n9774), .ZN(n9776) );
  NAND2_X1 U10665 ( .A1(n9776), .A2(n9775), .ZN(n9777) );
  XNOR2_X1 U10666 ( .A(n9778), .B(n9777), .ZN(n9784) );
  AOI22_X1 U10667 ( .A1(n9987), .A2(n9805), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9780) );
  NAND2_X1 U10668 ( .A1(n9804), .A2(n9981), .ZN(n9779) );
  OAI211_X1 U10669 ( .C1(n9781), .C2(n9808), .A(n9780), .B(n9779), .ZN(n9782)
         );
  AOI21_X1 U10670 ( .B1(n10114), .B2(n9811), .A(n9782), .ZN(n9783) );
  OAI21_X1 U10671 ( .B1(n9784), .B2(n9813), .A(n9783), .ZN(P1_U3233) );
  INV_X1 U10672 ( .A(n9787), .ZN(n9791) );
  AOI21_X1 U10673 ( .B1(n9787), .B2(n9786), .A(n9785), .ZN(n9788) );
  NOR2_X1 U10674 ( .A1(n9788), .A2(n9813), .ZN(n9789) );
  OAI21_X1 U10675 ( .B1(n9791), .B2(n9790), .A(n9789), .ZN(n9800) );
  OAI22_X1 U10676 ( .A1(n9794), .A2(n9793), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9792), .ZN(n9797) );
  NOR2_X1 U10677 ( .A1(n9795), .A2(n10049), .ZN(n9796) );
  AOI211_X1 U10678 ( .C1(n9798), .C2(n10064), .A(n9797), .B(n9796), .ZN(n9799)
         );
  OAI211_X1 U10679 ( .C1(n10052), .C2(n9801), .A(n9800), .B(n9799), .ZN(
        P1_U3236) );
  XNOR2_X1 U10680 ( .A(n9803), .B(n9802), .ZN(n9814) );
  NAND2_X1 U10681 ( .A1(n9804), .A2(n9925), .ZN(n9807) );
  AOI22_X1 U10682 ( .A1(n9805), .A2(n9953), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9806) );
  OAI211_X1 U10683 ( .C1(n9809), .C2(n9808), .A(n9807), .B(n9806), .ZN(n9810)
         );
  AOI21_X1 U10684 ( .B1(n9922), .B2(n9811), .A(n9810), .ZN(n9812) );
  OAI21_X1 U10685 ( .B1(n9814), .B2(n9813), .A(n9812), .ZN(P1_U3238) );
  MUX2_X1 U10686 ( .A(n9815), .B(P1_DATAO_REG_31__SCAN_IN), .S(n9830), .Z(
        P1_U3586) );
  MUX2_X1 U10687 ( .A(n9816), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9830), .Z(
        P1_U3585) );
  MUX2_X1 U10688 ( .A(n9905), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9830), .Z(
        P1_U3583) );
  MUX2_X1 U10689 ( .A(n9942), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9830), .Z(
        P1_U3581) );
  MUX2_X1 U10690 ( .A(n9953), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9830), .Z(
        P1_U3580) );
  MUX2_X1 U10691 ( .A(n9971), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9830), .Z(
        P1_U3579) );
  MUX2_X1 U10692 ( .A(n9988), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9830), .Z(
        P1_U3578) );
  MUX2_X1 U10693 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9987), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10694 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n10064), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10695 ( .A(n10041), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9830), .Z(
        P1_U3573) );
  MUX2_X1 U10696 ( .A(n9817), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9830), .Z(
        P1_U3571) );
  MUX2_X1 U10697 ( .A(n10976), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9830), .Z(
        P1_U3570) );
  MUX2_X1 U10698 ( .A(n9818), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9830), .Z(
        P1_U3569) );
  MUX2_X1 U10699 ( .A(n9819), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9830), .Z(
        P1_U3568) );
  MUX2_X1 U10700 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9820), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10701 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9821), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10702 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9822), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10703 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9823), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10704 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9824), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10705 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9825), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10706 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9826), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10707 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9827), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10708 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9828), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10709 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9829), .S(P1_U4006), .Z(
        P1_U3556) );
  MUX2_X1 U10710 ( .A(n9831), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9830), .Z(
        P1_U3555) );
  AOI22_X1 U10711 ( .A1(n10661), .A2(n9833), .B1(P1_U3084), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n9843) );
  XNOR2_X1 U10712 ( .A(n9835), .B(n9834), .ZN(n9836) );
  AOI22_X1 U10713 ( .A1(n10666), .A2(n9836), .B1(n10679), .B2(
        P1_ADDR_REG_2__SCAN_IN), .ZN(n9842) );
  INV_X1 U10714 ( .A(n9853), .ZN(n9840) );
  NAND3_X1 U10715 ( .A1(n10680), .A2(n9838), .A3(n9837), .ZN(n9839) );
  NAND3_X1 U10716 ( .A1(n10681), .A2(n9840), .A3(n9839), .ZN(n9841) );
  NAND4_X1 U10717 ( .A1(n9844), .A2(n9843), .A3(n9842), .A4(n9841), .ZN(
        P1_U3243) );
  INV_X1 U10718 ( .A(n9845), .ZN(n9846) );
  AOI211_X1 U10719 ( .C1(n9848), .C2(n9847), .A(n9846), .B(n10684), .ZN(n9849)
         );
  AOI21_X1 U10720 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(n10679), .A(n9849), .ZN(
        n9859) );
  INV_X1 U10721 ( .A(n9850), .ZN(n9851) );
  AOI22_X1 U10722 ( .A1(n10661), .A2(n9851), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        P1_U3084), .ZN(n9858) );
  OR3_X1 U10723 ( .A1(n9854), .A2(n9853), .A3(n9852), .ZN(n9855) );
  NAND3_X1 U10724 ( .A1(n10681), .A2(n9856), .A3(n9855), .ZN(n9857) );
  NAND3_X1 U10725 ( .A1(n9859), .A2(n9858), .A3(n9857), .ZN(P1_U3244) );
  AOI21_X1 U10726 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9868), .A(n9860), .ZN(
        n9863) );
  XNOR2_X1 U10727 ( .A(n9882), .B(n9861), .ZN(n9862) );
  NAND2_X1 U10728 ( .A1(n9863), .A2(n9862), .ZN(n9881) );
  OAI21_X1 U10729 ( .B1(n9863), .B2(n9862), .A(n9881), .ZN(n9874) );
  NAND2_X1 U10730 ( .A1(n10679), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n9865) );
  NAND2_X1 U10731 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3084), .ZN(n9864) );
  OAI211_X1 U10732 ( .C1(n9866), .C2(n10677), .A(n9865), .B(n9864), .ZN(n9873)
         );
  AOI21_X1 U10733 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n9868), .A(n9867), .ZN(
        n9871) );
  NAND2_X1 U10734 ( .A1(n9882), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9869) );
  OAI21_X1 U10735 ( .B1(n9882), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9869), .ZN(
        n9870) );
  NOR2_X1 U10736 ( .A1(n9871), .A2(n9870), .ZN(n9877) );
  AOI211_X1 U10737 ( .C1(n9871), .C2(n9870), .A(n9877), .B(n9890), .ZN(n9872)
         );
  AOI211_X1 U10738 ( .C1(n10666), .C2(n9874), .A(n9873), .B(n9872), .ZN(n9875)
         );
  INV_X1 U10739 ( .A(n9875), .ZN(P1_U3259) );
  INV_X1 U10740 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9876) );
  MUX2_X1 U10741 ( .A(n9876), .B(P1_REG2_REG_19__SCAN_IN), .S(n9958), .Z(n9879) );
  AOI21_X1 U10742 ( .B1(n9882), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9877), .ZN(
        n9878) );
  XOR2_X1 U10743 ( .A(n9879), .B(n9878), .Z(n9891) );
  INV_X1 U10744 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9880) );
  MUX2_X1 U10745 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9880), .S(n9958), .Z(n9884) );
  OAI21_X1 U10746 ( .B1(n9882), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9881), .ZN(
        n9883) );
  XOR2_X1 U10747 ( .A(n9884), .B(n9883), .Z(n9885) );
  AOI22_X1 U10748 ( .A1(n10666), .A2(n9885), .B1(n10679), .B2(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n9889) );
  INV_X1 U10749 ( .A(n9886), .ZN(n9887) );
  AOI21_X1 U10750 ( .B1(n10661), .B2(n10021), .A(n9887), .ZN(n9888) );
  OAI211_X1 U10751 ( .C1(n9891), .C2(n9890), .A(n9889), .B(n9888), .ZN(
        P1_U3260) );
  INV_X1 U10752 ( .A(n9892), .ZN(n9894) );
  NAND2_X1 U10753 ( .A1(n9894), .A2(n9893), .ZN(n10074) );
  NAND3_X1 U10754 ( .A1(n10074), .A2(n10068), .A3(n10073), .ZN(n9897) );
  AOI21_X1 U10755 ( .B1(n11006), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9895), .ZN(
        n9896) );
  OAI211_X1 U10756 ( .C1(n10077), .C2(n10734), .A(n9897), .B(n9896), .ZN(
        P1_U3262) );
  XOR2_X1 U10757 ( .A(n9904), .B(n9898), .Z(n10092) );
  NOR2_X1 U10758 ( .A1(n9902), .A2(n9924), .ZN(n9900) );
  NOR2_X1 U10759 ( .A1(n9900), .A2(n9899), .ZN(n10089) );
  INV_X1 U10760 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9901) );
  OAI22_X1 U10761 ( .A1(n9902), .A2(n10734), .B1(n9901), .B2(n10022), .ZN(
        n9909) );
  NAND2_X1 U10762 ( .A1(n10994), .A2(n9906), .ZN(n9907) );
  AOI21_X1 U10763 ( .B1(n10091), .B2(n9907), .A(n10738), .ZN(n9908) );
  AOI211_X1 U10764 ( .C1(n10068), .C2(n10089), .A(n9909), .B(n9908), .ZN(n9910) );
  OAI21_X1 U10765 ( .B1(n10092), .B2(n10070), .A(n9910), .ZN(P1_U3264) );
  NAND2_X1 U10766 ( .A1(n10093), .A2(n10879), .ZN(n9921) );
  OAI21_X1 U10767 ( .B1(n9914), .B2(n9913), .A(n9912), .ZN(n9919) );
  NAND2_X1 U10768 ( .A1(n9953), .A2(n10975), .ZN(n9917) );
  NAND2_X1 U10769 ( .A1(n9915), .A2(n10977), .ZN(n9916) );
  NAND2_X1 U10770 ( .A1(n9917), .A2(n9916), .ZN(n9918) );
  AOI21_X1 U10771 ( .B1(n9919), .B2(n10980), .A(n9918), .ZN(n9920) );
  NAND2_X1 U10772 ( .A1(n9921), .A2(n9920), .ZN(n10097) );
  INV_X1 U10773 ( .A(n10097), .ZN(n9931) );
  AND2_X1 U10774 ( .A1(n9922), .A2(n9933), .ZN(n9923) );
  NOR2_X1 U10775 ( .A1(n10095), .A2(n10733), .ZN(n9928) );
  AOI22_X1 U10776 ( .A1(n10738), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9925), 
        .B2(n10994), .ZN(n9926) );
  OAI21_X1 U10777 ( .B1(n10094), .B2(n10734), .A(n9926), .ZN(n9927) );
  AOI211_X1 U10778 ( .C1(n10093), .C2(n9929), .A(n9928), .B(n9927), .ZN(n9930)
         );
  OAI21_X1 U10779 ( .B1(n9931), .B2(n11006), .A(n9930), .ZN(P1_U3265) );
  XNOR2_X1 U10780 ( .A(n9932), .B(n9941), .ZN(n10103) );
  INV_X1 U10781 ( .A(n9955), .ZN(n9935) );
  INV_X1 U10782 ( .A(n9933), .ZN(n9934) );
  AOI21_X1 U10783 ( .B1(n10099), .B2(n9935), .A(n9934), .ZN(n10100) );
  AOI22_X1 U10784 ( .A1(n10738), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9936), 
        .B2(n10994), .ZN(n9937) );
  OAI21_X1 U10785 ( .B1(n9938), .B2(n10734), .A(n9937), .ZN(n9945) );
  OAI21_X1 U10786 ( .B1(n9941), .B2(n9940), .A(n9939), .ZN(n9943) );
  AOI222_X1 U10787 ( .A1(n9943), .A2(n10980), .B1(n9942), .B2(n10977), .C1(
        n9971), .C2(n10975), .ZN(n10102) );
  NOR2_X1 U10788 ( .A1(n10102), .A2(n10738), .ZN(n9944) );
  AOI211_X1 U10789 ( .C1(n10100), .C2(n10068), .A(n9945), .B(n9944), .ZN(n9946) );
  OAI21_X1 U10790 ( .B1(n10103), .B2(n10070), .A(n9946), .ZN(P1_U3266) );
  XNOR2_X1 U10791 ( .A(n9947), .B(n9948), .ZN(n10108) );
  NOR2_X1 U10792 ( .A1(n9949), .A2(n10734), .ZN(n9961) );
  OAI21_X1 U10793 ( .B1(n9952), .B2(n9951), .A(n9950), .ZN(n9954) );
  AOI222_X1 U10794 ( .A1(n9954), .A2(n10980), .B1(n9953), .B2(n10977), .C1(
        n9988), .C2(n10975), .ZN(n10107) );
  INV_X1 U10795 ( .A(n9965), .ZN(n9956) );
  AOI211_X1 U10796 ( .C1(n10105), .C2(n9956), .A(n10960), .B(n9955), .ZN(
        n10104) );
  AOI22_X1 U10797 ( .A1(n10104), .A2(n9958), .B1(n10994), .B2(n9957), .ZN(
        n9959) );
  AOI21_X1 U10798 ( .B1(n10107), .B2(n9959), .A(n10738), .ZN(n9960) );
  AOI211_X1 U10799 ( .C1(n11006), .C2(P1_REG2_REG_24__SCAN_IN), .A(n9961), .B(
        n9960), .ZN(n9962) );
  OAI21_X1 U10800 ( .B1(n10070), .B2(n10108), .A(n9962), .ZN(P1_U3267) );
  XNOR2_X1 U10801 ( .A(n9963), .B(n9964), .ZN(n10113) );
  AOI21_X1 U10802 ( .B1(n10109), .B2(n9979), .A(n9965), .ZN(n10110) );
  AOI22_X1 U10803 ( .A1(n10738), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9966), 
        .B2(n10994), .ZN(n9967) );
  OAI21_X1 U10804 ( .B1(n5313), .B2(n10734), .A(n9967), .ZN(n9974) );
  OAI21_X1 U10805 ( .B1(n9970), .B2(n9969), .A(n9968), .ZN(n9972) );
  AOI222_X1 U10806 ( .A1(n9972), .A2(n10980), .B1(n9971), .B2(n10977), .C1(
        n9997), .C2(n10975), .ZN(n10112) );
  NOR2_X1 U10807 ( .A1(n10112), .A2(n11006), .ZN(n9973) );
  AOI211_X1 U10808 ( .C1(n10110), .C2(n10068), .A(n9974), .B(n9973), .ZN(n9975) );
  OAI21_X1 U10809 ( .B1(n10070), .B2(n10113), .A(n9975), .ZN(P1_U3268) );
  OAI21_X1 U10810 ( .B1(n9978), .B2(n9977), .A(n9976), .ZN(n10118) );
  INV_X1 U10811 ( .A(n9979), .ZN(n9980) );
  AOI21_X1 U10812 ( .B1(n10114), .B2(n9993), .A(n9980), .ZN(n10115) );
  AOI22_X1 U10813 ( .A1(n10738), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9981), 
        .B2(n10994), .ZN(n9982) );
  OAI21_X1 U10814 ( .B1(n9983), .B2(n10734), .A(n9982), .ZN(n9991) );
  OAI21_X1 U10815 ( .B1(n9986), .B2(n9985), .A(n9984), .ZN(n9989) );
  AOI222_X1 U10816 ( .A1(n9989), .A2(n10980), .B1(n9988), .B2(n10977), .C1(
        n9987), .C2(n10975), .ZN(n10117) );
  NOR2_X1 U10817 ( .A1(n10117), .A2(n10738), .ZN(n9990) );
  AOI211_X1 U10818 ( .C1(n10115), .C2(n10068), .A(n9991), .B(n9990), .ZN(n9992) );
  OAI21_X1 U10819 ( .B1(n10070), .B2(n10118), .A(n9992), .ZN(P1_U3269) );
  INV_X1 U10820 ( .A(n10120), .ZN(n9994) );
  OAI211_X1 U10821 ( .C1(n5112), .C2(n9994), .A(n10981), .B(n9993), .ZN(n10121) );
  NOR2_X1 U10822 ( .A1(n10121), .A2(n10021), .ZN(n10000) );
  OAI21_X1 U10823 ( .B1(n10003), .B2(n9996), .A(n9995), .ZN(n9998) );
  AOI222_X1 U10824 ( .A1(n9998), .A2(n10980), .B1(n9997), .B2(n10977), .C1(
        n10040), .C2(n10975), .ZN(n10123) );
  INV_X1 U10825 ( .A(n10123), .ZN(n9999) );
  AOI211_X1 U10826 ( .C1(n10994), .C2(n10001), .A(n10000), .B(n9999), .ZN(
        n10007) );
  AOI22_X1 U10827 ( .A1(n10120), .A2(n10996), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n10738), .ZN(n10006) );
  NAND2_X1 U10828 ( .A1(n10004), .A2(n10003), .ZN(n10119) );
  INV_X1 U10829 ( .A(n10070), .ZN(n11001) );
  NAND3_X1 U10830 ( .A1(n10002), .A2(n10119), .A3(n11001), .ZN(n10005) );
  OAI211_X1 U10831 ( .C1(n10007), .C2(n10738), .A(n10006), .B(n10005), .ZN(
        P1_U3270) );
  XNOR2_X1 U10832 ( .A(n10008), .B(n5330), .ZN(n10129) );
  INV_X1 U10833 ( .A(n10032), .ZN(n10009) );
  AOI211_X1 U10834 ( .C1(n10009), .C2(n10126), .A(n10960), .B(n5112), .ZN(
        n10125) );
  INV_X1 U10835 ( .A(n10125), .ZN(n10020) );
  OAI21_X1 U10836 ( .B1(n10012), .B2(n10011), .A(n10010), .ZN(n10019) );
  OAI22_X1 U10837 ( .A1(n10016), .A2(n10015), .B1(n10014), .B2(n10013), .ZN(
        n10018) );
  NOR2_X1 U10838 ( .A1(n10129), .A2(n7169), .ZN(n10017) );
  AOI211_X1 U10839 ( .C1(n10980), .C2(n10019), .A(n10018), .B(n10017), .ZN(
        n10128) );
  OAI21_X1 U10840 ( .B1(n10021), .B2(n10020), .A(n10128), .ZN(n10023) );
  NAND2_X1 U10841 ( .A1(n10023), .A2(n10022), .ZN(n10028) );
  NAND2_X1 U10842 ( .A1(n10738), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n10024) );
  OAI21_X1 U10843 ( .B1(n10741), .B2(n10025), .A(n10024), .ZN(n10026) );
  AOI21_X1 U10844 ( .B1(n10126), .B2(n10996), .A(n10026), .ZN(n10027) );
  OAI211_X1 U10845 ( .C1(n10129), .C2(n10029), .A(n10028), .B(n10027), .ZN(
        P1_U3271) );
  XNOR2_X1 U10846 ( .A(n10030), .B(n10031), .ZN(n10134) );
  INV_X1 U10847 ( .A(n10047), .ZN(n10033) );
  AOI21_X1 U10848 ( .B1(n10130), .B2(n10033), .A(n10032), .ZN(n10131) );
  INV_X1 U10849 ( .A(n10034), .ZN(n10035) );
  AOI22_X1 U10850 ( .A1(n10738), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n10035), 
        .B2(n10994), .ZN(n10036) );
  OAI21_X1 U10851 ( .B1(n10037), .B2(n10734), .A(n10036), .ZN(n10044) );
  OAI21_X1 U10852 ( .B1(n5116), .B2(n10039), .A(n10038), .ZN(n10042) );
  AOI222_X1 U10853 ( .A1(n10042), .A2(n10980), .B1(n10041), .B2(n10975), .C1(
        n10040), .C2(n10977), .ZN(n10133) );
  NOR2_X1 U10854 ( .A1(n10133), .A2(n10738), .ZN(n10043) );
  AOI211_X1 U10855 ( .C1(n10068), .C2(n10131), .A(n10044), .B(n10043), .ZN(
        n10045) );
  OAI21_X1 U10856 ( .B1(n10134), .B2(n10070), .A(n10045), .ZN(P1_U3272) );
  XNOR2_X1 U10857 ( .A(n10046), .B(n10060), .ZN(n10538) );
  AOI21_X1 U10858 ( .B1(n10534), .B2(n10048), .A(n10047), .ZN(n10535) );
  INV_X1 U10859 ( .A(n10049), .ZN(n10050) );
  AOI22_X1 U10860 ( .A1(n10738), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n10050), 
        .B2(n10994), .ZN(n10051) );
  OAI21_X1 U10861 ( .B1(n10052), .B2(n10734), .A(n10051), .ZN(n10067) );
  AOI21_X1 U10862 ( .B1(n10058), .B2(n10054), .A(n10053), .ZN(n10056) );
  MUX2_X1 U10863 ( .A(n10057), .B(n10056), .S(n10055), .Z(n10063) );
  INV_X1 U10864 ( .A(n10058), .ZN(n10061) );
  NAND3_X1 U10865 ( .A1(n10061), .A2(n10060), .A3(n10059), .ZN(n10062) );
  NAND2_X1 U10866 ( .A1(n10063), .A2(n10062), .ZN(n10065) );
  AOI222_X1 U10867 ( .A1(n10980), .A2(n10065), .B1(n10978), .B2(n10975), .C1(
        n10064), .C2(n10977), .ZN(n10537) );
  NOR2_X1 U10868 ( .A1(n10537), .A2(n11006), .ZN(n10066) );
  AOI211_X1 U10869 ( .C1(n10535), .C2(n10068), .A(n10067), .B(n10066), .ZN(
        n10069) );
  OAI21_X1 U10870 ( .B1(n10538), .B2(n10070), .A(n10069), .ZN(P1_U3273) );
  MUX2_X1 U10871 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10547), .S(n10989), .Z(
        P1_U3554) );
  NAND3_X1 U10872 ( .A1(n10074), .A2(n10981), .A3(n10073), .ZN(n10076) );
  OAI211_X1 U10873 ( .C1(n10077), .C2(n10984), .A(n10076), .B(n10075), .ZN(
        n10548) );
  MUX2_X1 U10874 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10548), .S(n10989), .Z(
        P1_U3553) );
  AOI22_X1 U10875 ( .A1(n10079), .A2(n10981), .B1(n10873), .B2(n10078), .ZN(
        n10080) );
  MUX2_X1 U10876 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10549), .S(n10989), .Z(
        P1_U3552) );
  AOI22_X1 U10877 ( .A1(n10084), .A2(n10981), .B1(n10873), .B2(n10083), .ZN(
        n10085) );
  MUX2_X1 U10878 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10550), .S(n10989), .Z(
        P1_U3551) );
  AOI22_X1 U10879 ( .A1(n10089), .A2(n10981), .B1(n10873), .B2(n10088), .ZN(
        n10090) );
  OAI211_X1 U10880 ( .C1(n10092), .C2(n10539), .A(n10091), .B(n10090), .ZN(
        n10551) );
  MUX2_X1 U10881 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10551), .S(n10989), .Z(
        P1_U3550) );
  OAI22_X1 U10882 ( .A1(n10095), .A2(n10960), .B1(n10094), .B2(n10984), .ZN(
        n10096) );
  MUX2_X1 U10883 ( .A(n10552), .B(P1_REG1_REG_26__SCAN_IN), .S(n10987), .Z(
        P1_U3549) );
  AOI22_X1 U10884 ( .A1(n10100), .A2(n10981), .B1(n10873), .B2(n10099), .ZN(
        n10101) );
  OAI211_X1 U10885 ( .C1(n10103), .C2(n10539), .A(n10102), .B(n10101), .ZN(
        n10553) );
  MUX2_X1 U10886 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10553), .S(n10989), .Z(
        P1_U3548) );
  AOI21_X1 U10887 ( .B1(n10873), .B2(n10105), .A(n10104), .ZN(n10106) );
  OAI211_X1 U10888 ( .C1(n10108), .C2(n10539), .A(n10107), .B(n10106), .ZN(
        n10554) );
  MUX2_X1 U10889 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10554), .S(n10989), .Z(
        P1_U3547) );
  AOI22_X1 U10890 ( .A1(n10110), .A2(n10981), .B1(n10873), .B2(n10109), .ZN(
        n10111) );
  OAI211_X1 U10891 ( .C1(n10113), .C2(n10539), .A(n10112), .B(n10111), .ZN(
        n10555) );
  MUX2_X1 U10892 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10555), .S(n10989), .Z(
        P1_U3546) );
  AOI22_X1 U10893 ( .A1(n10115), .A2(n10981), .B1(n10873), .B2(n10114), .ZN(
        n10116) );
  OAI211_X1 U10894 ( .C1(n10118), .C2(n10539), .A(n10117), .B(n10116), .ZN(
        n10556) );
  MUX2_X1 U10895 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10556), .S(n10989), .Z(
        P1_U3545) );
  NAND3_X1 U10896 ( .A1(n10002), .A2(n5587), .A3(n10119), .ZN(n10124) );
  NAND2_X1 U10897 ( .A1(n10120), .A2(n10873), .ZN(n10122) );
  NAND4_X1 U10898 ( .A1(n10124), .A2(n10123), .A3(n10122), .A4(n10121), .ZN(
        n10557) );
  MUX2_X1 U10899 ( .A(n10557), .B(P1_REG1_REG_21__SCAN_IN), .S(n10987), .Z(
        P1_U3544) );
  AOI21_X1 U10900 ( .B1(n10873), .B2(n10126), .A(n10125), .ZN(n10127) );
  OAI211_X1 U10901 ( .C1(n10875), .C2(n10129), .A(n10128), .B(n10127), .ZN(
        n10558) );
  MUX2_X1 U10902 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10558), .S(n10989), .Z(
        P1_U3543) );
  AOI22_X1 U10903 ( .A1(n10131), .A2(n10981), .B1(n10873), .B2(n10130), .ZN(
        n10132) );
  OAI211_X1 U10904 ( .C1(n10134), .C2(n10539), .A(n10133), .B(n10132), .ZN(
        n10559) );
  MUX2_X1 U10905 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10559), .S(n10989), .Z(
        n10533) );
  INV_X1 U10906 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10531) );
  INV_X1 U10907 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10136) );
  AOI22_X1 U10908 ( .A1(n10136), .A2(keyinput_252), .B1(n10582), .B2(
        keyinput_253), .ZN(n10135) );
  OAI221_X1 U10909 ( .B1(n10136), .B2(keyinput_252), .C1(n10582), .C2(
        keyinput_253), .A(n10135), .ZN(n10347) );
  INV_X1 U10910 ( .A(keyinput_200), .ZN(n10263) );
  INV_X1 U10911 ( .A(keyinput_199), .ZN(n10261) );
  INV_X1 U10912 ( .A(keyinput_197), .ZN(n10254) );
  XOR2_X1 U10913 ( .A(n10137), .B(keyinput_186), .Z(n10243) );
  INV_X1 U10914 ( .A(keyinput_184), .ZN(n10230) );
  INV_X1 U10915 ( .A(keyinput_182), .ZN(n10226) );
  OAI22_X1 U10916 ( .A1(n7650), .A2(keyinput_171), .B1(keyinput_169), .B2(
        P2_REG3_REG_19__SCAN_IN), .ZN(n10138) );
  AOI221_X1 U10917 ( .B1(n7650), .B2(keyinput_171), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput_169), .A(n10138), .ZN(n10209)
         );
  AOI22_X1 U10918 ( .A1(n10141), .A2(keyinput_166), .B1(n10140), .B2(
        keyinput_167), .ZN(n10139) );
  OAI221_X1 U10919 ( .B1(n10141), .B2(keyinput_166), .C1(n10140), .C2(
        keyinput_167), .A(n10139), .ZN(n10207) );
  INV_X1 U10920 ( .A(SI_7_), .ZN(n10143) );
  OAI22_X1 U10921 ( .A1(n10143), .A2(keyinput_153), .B1(keyinput_154), .B2(
        SI_6_), .ZN(n10142) );
  AOI221_X1 U10922 ( .B1(n10143), .B2(keyinput_153), .C1(SI_6_), .C2(
        keyinput_154), .A(n10142), .ZN(n10191) );
  XNOR2_X1 U10923 ( .A(n10144), .B(keyinput_150), .ZN(n10189) );
  AOI22_X1 U10924 ( .A1(SI_13_), .A2(keyinput_147), .B1(n10146), .B2(
        keyinput_148), .ZN(n10145) );
  OAI221_X1 U10925 ( .B1(SI_13_), .B2(keyinput_147), .C1(n10146), .C2(
        keyinput_148), .A(n10145), .ZN(n10184) );
  XNOR2_X1 U10926 ( .A(SI_18_), .B(keyinput_142), .ZN(n10183) );
  INV_X1 U10927 ( .A(keyinput_140), .ZN(n10169) );
  OAI22_X1 U10928 ( .A1(SI_25_), .A2(keyinput_135), .B1(keyinput_136), .B2(
        SI_24_), .ZN(n10147) );
  AOI221_X1 U10929 ( .B1(SI_25_), .B2(keyinput_135), .C1(SI_24_), .C2(
        keyinput_136), .A(n10147), .ZN(n10160) );
  OAI221_X1 U10930 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_128), .C1(SI_31_), 
        .C2(keyinput_129), .A(n10148), .ZN(n10151) );
  INV_X1 U10931 ( .A(keyinput_130), .ZN(n10149) );
  MUX2_X1 U10932 ( .A(keyinput_130), .B(n10149), .S(SI_30_), .Z(n10150) );
  NAND2_X1 U10933 ( .A1(n10151), .A2(n10150), .ZN(n10158) );
  INV_X1 U10934 ( .A(keyinput_131), .ZN(n10152) );
  MUX2_X1 U10935 ( .A(keyinput_131), .B(n10152), .S(SI_29_), .Z(n10157) );
  XNOR2_X1 U10936 ( .A(n10153), .B(keyinput_132), .ZN(n10156) );
  XNOR2_X1 U10937 ( .A(n10154), .B(keyinput_133), .ZN(n10155) );
  AOI211_X1 U10938 ( .C1(n10158), .C2(n10157), .A(n10156), .B(n10155), .ZN(
        n10159) );
  INV_X1 U10939 ( .A(keyinput_138), .ZN(n10162) );
  MUX2_X1 U10940 ( .A(n10162), .B(keyinput_138), .S(SI_22_), .Z(n10163) );
  NAND2_X1 U10941 ( .A1(n10164), .A2(n10163), .ZN(n10167) );
  INV_X1 U10942 ( .A(keyinput_139), .ZN(n10165) );
  MUX2_X1 U10943 ( .A(n10165), .B(keyinput_139), .S(SI_21_), .Z(n10166) );
  NAND2_X1 U10944 ( .A1(n10167), .A2(n10166), .ZN(n10168) );
  OAI221_X1 U10945 ( .B1(SI_20_), .B2(keyinput_140), .C1(n10170), .C2(n10169), 
        .A(n10168), .ZN(n10175) );
  INV_X1 U10946 ( .A(keyinput_141), .ZN(n10171) );
  INV_X1 U10947 ( .A(SI_15_), .ZN(n10178) );
  INV_X1 U10948 ( .A(SI_17_), .ZN(n10177) );
  AOI22_X1 U10949 ( .A1(n10178), .A2(keyinput_145), .B1(n10177), .B2(
        keyinput_143), .ZN(n10176) );
  OAI221_X1 U10950 ( .B1(n10178), .B2(keyinput_145), .C1(n10177), .C2(
        keyinput_143), .A(n10176), .ZN(n10182) );
  INV_X1 U10951 ( .A(SI_14_), .ZN(n10180) );
  AOI22_X1 U10952 ( .A1(SI_16_), .A2(keyinput_144), .B1(n10180), .B2(
        keyinput_146), .ZN(n10179) );
  OAI221_X1 U10953 ( .B1(SI_16_), .B2(keyinput_144), .C1(n10180), .C2(
        keyinput_146), .A(n10179), .ZN(n10181) );
  OAI22_X1 U10954 ( .A1(n10186), .A2(keyinput_151), .B1(SI_8_), .B2(
        keyinput_152), .ZN(n10185) );
  AOI221_X1 U10955 ( .B1(n10186), .B2(keyinput_151), .C1(keyinput_152), .C2(
        SI_8_), .A(n10185), .ZN(n10187) );
  OAI21_X1 U10956 ( .B1(n10189), .B2(n10188), .A(n10187), .ZN(n10190) );
  AOI22_X1 U10957 ( .A1(SI_3_), .A2(keyinput_157), .B1(n10193), .B2(
        keyinput_156), .ZN(n10192) );
  OAI221_X1 U10958 ( .B1(SI_3_), .B2(keyinput_157), .C1(n10193), .C2(
        keyinput_156), .A(n10192), .ZN(n10194) );
  XNOR2_X1 U10959 ( .A(SI_1_), .B(keyinput_159), .ZN(n10196) );
  XNOR2_X1 U10960 ( .A(SI_2_), .B(keyinput_158), .ZN(n10195) );
  OAI22_X1 U10961 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput_163), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_164), .ZN(n10197) );
  AOI221_X1 U10962 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_163), .C1(
        keyinput_164), .C2(P2_REG3_REG_27__SCAN_IN), .A(n10197), .ZN(n10201)
         );
  INV_X1 U10963 ( .A(SI_0_), .ZN(n10199) );
  OAI22_X1 U10964 ( .A1(n10199), .A2(keyinput_160), .B1(keyinput_168), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n10198) );
  AOI221_X1 U10965 ( .B1(n10199), .B2(keyinput_160), .C1(
        P2_REG3_REG_3__SCAN_IN), .C2(keyinput_168), .A(n10198), .ZN(n10200) );
  AOI22_X1 U10966 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_165), .B1(
        P2_U3152), .B2(keyinput_162), .ZN(n10202) );
  OAI221_X1 U10967 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_165), .C1(
        P2_U3152), .C2(keyinput_162), .A(n10202), .ZN(n10204) );
  AOI22_X1 U10968 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_173), .B1(
        P2_REG3_REG_12__SCAN_IN), .B2(keyinput_174), .ZN(n10211) );
  OAI221_X1 U10969 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_173), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_174), .A(n10211), .ZN(n10217)
         );
  OAI22_X1 U10970 ( .A1(n10213), .A2(keyinput_175), .B1(keyinput_178), .B2(
        P2_REG3_REG_17__SCAN_IN), .ZN(n10212) );
  AOI221_X1 U10971 ( .B1(n10213), .B2(keyinput_175), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput_178), .A(n10212), .ZN(n10216)
         );
  OAI22_X1 U10972 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_177), .B1(
        keyinput_176), .B2(P2_REG3_REG_16__SCAN_IN), .ZN(n10214) );
  AOI221_X1 U10973 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_177), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput_176), .A(n10214), .ZN(n10215)
         );
  OAI22_X1 U10974 ( .A1(n10219), .A2(keyinput_179), .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_180), .ZN(n10218) );
  AOI221_X1 U10975 ( .B1(n10219), .B2(keyinput_179), .C1(keyinput_180), .C2(
        P2_REG3_REG_4__SCAN_IN), .A(n10218), .ZN(n10220) );
  NAND2_X1 U10976 ( .A1(n10221), .A2(n10220), .ZN(n10224) );
  INV_X1 U10977 ( .A(keyinput_183), .ZN(n10227) );
  INV_X1 U10978 ( .A(keyinput_185), .ZN(n10232) );
  AOI22_X1 U10979 ( .A1(n5810), .A2(keyinput_189), .B1(keyinput_187), .B2(
        n10238), .ZN(n10237) );
  OAI221_X1 U10980 ( .B1(n5810), .B2(keyinput_189), .C1(n10238), .C2(
        keyinput_187), .A(n10237), .ZN(n10241) );
  AOI22_X1 U10981 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_190), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_188), .ZN(n10239) );
  OAI221_X1 U10982 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_190), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput_188), .A(n10239), .ZN(n10240)
         );
  AOI211_X1 U10983 ( .C1(n10243), .C2(n10242), .A(n10241), .B(n10240), .ZN(
        n10251) );
  AOI22_X1 U10984 ( .A1(P2_B_REG_SCAN_IN), .A2(keyinput_192), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput_191), .ZN(n10244) );
  OAI221_X1 U10985 ( .B1(P2_B_REG_SCAN_IN), .B2(keyinput_192), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput_191), .A(n10244), .ZN(n10250)
         );
  OAI22_X1 U10986 ( .A1(n10246), .A2(keyinput_195), .B1(keyinput_194), .B2(
        P2_DATAO_REG_30__SCAN_IN), .ZN(n10245) );
  AOI221_X1 U10987 ( .B1(n10246), .B2(keyinput_195), .C1(
        P2_DATAO_REG_30__SCAN_IN), .C2(keyinput_194), .A(n10245), .ZN(n10249)
         );
  OAI22_X1 U10988 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(keyinput_196), .B1(
        keyinput_193), .B2(P2_DATAO_REG_31__SCAN_IN), .ZN(n10247) );
  AOI221_X1 U10989 ( .B1(P2_DATAO_REG_28__SCAN_IN), .B2(keyinput_196), .C1(
        P2_DATAO_REG_31__SCAN_IN), .C2(keyinput_193), .A(n10247), .ZN(n10248)
         );
  OAI211_X1 U10990 ( .C1(n10251), .C2(n10250), .A(n10249), .B(n10248), .ZN(
        n10252) );
  OAI221_X1 U10991 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(n10254), .C1(n10253), 
        .C2(keyinput_197), .A(n10252), .ZN(n10258) );
  INV_X1 U10992 ( .A(keyinput_198), .ZN(n10255) );
  OAI221_X1 U10993 ( .B1(P2_DATAO_REG_25__SCAN_IN), .B2(n10261), .C1(n10260), 
        .C2(keyinput_199), .A(n10259), .ZN(n10262) );
  OAI221_X1 U10994 ( .B1(P2_DATAO_REG_24__SCAN_IN), .B2(keyinput_200), .C1(
        n10264), .C2(n10263), .A(n10262), .ZN(n10269) );
  OAI22_X1 U10995 ( .A1(n10266), .A2(keyinput_202), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(keyinput_201), .ZN(n10265) );
  AOI221_X1 U10996 ( .B1(n10266), .B2(keyinput_202), .C1(keyinput_201), .C2(
        P2_DATAO_REG_23__SCAN_IN), .A(n10265), .ZN(n10268) );
  OAI22_X1 U10997 ( .A1(n10272), .A2(keyinput_205), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_204), .ZN(n10271) );
  AOI221_X1 U10998 ( .B1(n10272), .B2(keyinput_205), .C1(keyinput_204), .C2(
        P2_DATAO_REG_20__SCAN_IN), .A(n10271), .ZN(n10275) );
  NOR2_X1 U10999 ( .A1(n10274), .A2(keyinput_206), .ZN(n10273) );
  AOI22_X1 U11000 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput_208), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_207), .ZN(n10277) );
  OAI221_X1 U11001 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput_208), .C1(
        P2_DATAO_REG_17__SCAN_IN), .C2(keyinput_207), .A(n10277), .ZN(n10284)
         );
  OAI22_X1 U11002 ( .A1(n10280), .A2(keyinput_209), .B1(n10279), .B2(
        keyinput_212), .ZN(n10278) );
  AOI221_X1 U11003 ( .B1(n10280), .B2(keyinput_209), .C1(keyinput_212), .C2(
        n10279), .A(n10278), .ZN(n10283) );
  OAI22_X1 U11004 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(keyinput_210), .B1(
        keyinput_211), .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n10281) );
  AOI221_X1 U11005 ( .B1(P2_DATAO_REG_14__SCAN_IN), .B2(keyinput_210), .C1(
        P2_DATAO_REG_13__SCAN_IN), .C2(keyinput_211), .A(n10281), .ZN(n10282)
         );
  OAI22_X1 U11006 ( .A1(n10287), .A2(keyinput_213), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_214), .ZN(n10286) );
  AOI221_X1 U11007 ( .B1(n10287), .B2(keyinput_213), .C1(keyinput_214), .C2(
        P2_DATAO_REG_10__SCAN_IN), .A(n10286), .ZN(n10288) );
  OAI22_X1 U11008 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput_215), .B1(
        keyinput_216), .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n10289) );
  AOI221_X1 U11009 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_215), .C1(
        P2_DATAO_REG_8__SCAN_IN), .C2(keyinput_216), .A(n10289), .ZN(n10292)
         );
  AOI22_X1 U11010 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(keyinput_218), .B1(
        n10656), .B2(keyinput_219), .ZN(n10290) );
  OAI221_X1 U11011 ( .B1(P2_DATAO_REG_6__SCAN_IN), .B2(keyinput_218), .C1(
        n10656), .C2(keyinput_219), .A(n10290), .ZN(n10291) );
  INV_X1 U11012 ( .A(keyinput_220), .ZN(n10293) );
  MUX2_X1 U11013 ( .A(n10293), .B(keyinput_220), .S(P1_IR_REG_1__SCAN_IN), .Z(
        n10298) );
  XNOR2_X1 U11014 ( .A(n10294), .B(keyinput_222), .ZN(n10297) );
  XNOR2_X1 U11015 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_221), .ZN(n10296) );
  XNOR2_X1 U11016 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_223), .ZN(n10295) );
  INV_X1 U11017 ( .A(keyinput_224), .ZN(n10299) );
  MUX2_X1 U11018 ( .A(n10299), .B(keyinput_224), .S(P1_IR_REG_5__SCAN_IN), .Z(
        n10306) );
  XNOR2_X1 U11019 ( .A(n10300), .B(keyinput_225), .ZN(n10304) );
  XNOR2_X1 U11020 ( .A(n10301), .B(keyinput_226), .ZN(n10303) );
  XNOR2_X1 U11021 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_227), .ZN(n10302) );
  NAND3_X1 U11022 ( .A1(n10304), .A2(n10303), .A3(n10302), .ZN(n10305) );
  AOI21_X1 U11023 ( .B1(n10307), .B2(n10306), .A(n10305), .ZN(n10314) );
  INV_X1 U11024 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n10309) );
  AOI22_X1 U11025 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput_228), .B1(n10309), 
        .B2(keyinput_229), .ZN(n10308) );
  OAI221_X1 U11026 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput_228), .C1(n10309), 
        .C2(keyinput_229), .A(n10308), .ZN(n10313) );
  XNOR2_X1 U11027 ( .A(n10310), .B(keyinput_231), .ZN(n10312) );
  XNOR2_X1 U11028 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_230), .ZN(n10311)
         );
  XOR2_X1 U11029 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_233), .Z(n10317) );
  XNOR2_X1 U11030 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_234), .ZN(n10316)
         );
  XNOR2_X1 U11031 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_232), .ZN(n10315)
         );
  NOR3_X1 U11032 ( .A1(n10317), .A2(n10316), .A3(n10315), .ZN(n10322) );
  XNOR2_X1 U11033 ( .A(n10318), .B(keyinput_236), .ZN(n10321) );
  XNOR2_X1 U11034 ( .A(n10319), .B(keyinput_235), .ZN(n10320) );
  OAI22_X1 U11035 ( .A1(n10325), .A2(keyinput_237), .B1(P1_IR_REG_19__SCAN_IN), 
        .B2(keyinput_238), .ZN(n10324) );
  AOI221_X1 U11036 ( .B1(n10325), .B2(keyinput_237), .C1(keyinput_238), .C2(
        P1_IR_REG_19__SCAN_IN), .A(n10324), .ZN(n10329) );
  XNOR2_X1 U11037 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_239), .ZN(n10328)
         );
  XNOR2_X1 U11038 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_241), .ZN(n10327)
         );
  XNOR2_X1 U11039 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_240), .ZN(n10326)
         );
  XNOR2_X1 U11040 ( .A(n10330), .B(keyinput_243), .ZN(n10332) );
  XNOR2_X1 U11041 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_244), .ZN(n10331)
         );
  XNOR2_X1 U11042 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_246), .ZN(n10335)
         );
  OAI22_X1 U11043 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(keyinput_245), .B1(
        P1_IR_REG_28__SCAN_IN), .B2(keyinput_247), .ZN(n10333) );
  AOI221_X1 U11044 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(keyinput_245), .C1(
        keyinput_247), .C2(P1_IR_REG_28__SCAN_IN), .A(n10333), .ZN(n10334) );
  INV_X1 U11045 ( .A(keyinput_248), .ZN(n10336) );
  MUX2_X1 U11046 ( .A(keyinput_248), .B(n10336), .S(P1_IR_REG_29__SCAN_IN), 
        .Z(n10343) );
  XOR2_X1 U11047 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_250), .Z(n10338) );
  XNOR2_X1 U11048 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_249), .ZN(n10337)
         );
  OAI211_X1 U11049 ( .C1(P1_D_REG_0__SCAN_IN), .C2(keyinput_251), .A(n10338), 
        .B(n10337), .ZN(n10339) );
  INV_X1 U11050 ( .A(n10339), .ZN(n10341) );
  NAND2_X1 U11051 ( .A1(n10583), .A2(keyinput_254), .ZN(n10345) );
  INV_X1 U11052 ( .A(n10349), .ZN(n10348) );
  OAI21_X1 U11053 ( .B1(n10348), .B2(keyinput_255), .A(keyinput_127), .ZN(
        n10530) );
  XOR2_X1 U11054 ( .A(SI_29_), .B(keyinput_3), .Z(n10356) );
  XNOR2_X1 U11055 ( .A(SI_31_), .B(keyinput_1), .ZN(n10352) );
  XNOR2_X1 U11056 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_0), .ZN(n10351) );
  XOR2_X1 U11057 ( .A(SI_30_), .B(keyinput_2), .Z(n10350) );
  OAI21_X1 U11058 ( .B1(n10352), .B2(n10351), .A(n10350), .ZN(n10355) );
  XNOR2_X1 U11059 ( .A(SI_27_), .B(keyinput_5), .ZN(n10354) );
  XOR2_X1 U11060 ( .A(SI_28_), .B(keyinput_4), .Z(n10353) );
  AOI211_X1 U11061 ( .C1(n10356), .C2(n10355), .A(n10354), .B(n10353), .ZN(
        n10360) );
  XOR2_X1 U11062 ( .A(SI_26_), .B(keyinput_6), .Z(n10359) );
  XOR2_X1 U11063 ( .A(SI_25_), .B(keyinput_7), .Z(n10358) );
  XNOR2_X1 U11064 ( .A(SI_24_), .B(keyinput_8), .ZN(n10357) );
  OAI211_X1 U11065 ( .C1(n10360), .C2(n10359), .A(n10358), .B(n10357), .ZN(
        n10363) );
  XOR2_X1 U11066 ( .A(SI_23_), .B(keyinput_9), .Z(n10362) );
  XNOR2_X1 U11067 ( .A(SI_22_), .B(keyinput_10), .ZN(n10361) );
  AOI21_X1 U11068 ( .B1(n10363), .B2(n10362), .A(n10361), .ZN(n10366) );
  XNOR2_X1 U11069 ( .A(SI_21_), .B(keyinput_11), .ZN(n10365) );
  XOR2_X1 U11070 ( .A(SI_20_), .B(keyinput_12), .Z(n10364) );
  OAI21_X1 U11071 ( .B1(n10366), .B2(n10365), .A(n10364), .ZN(n10369) );
  XNOR2_X1 U11072 ( .A(SI_19_), .B(keyinput_13), .ZN(n10368) );
  XNOR2_X1 U11073 ( .A(SI_18_), .B(keyinput_14), .ZN(n10367) );
  AOI21_X1 U11074 ( .B1(n10369), .B2(n10368), .A(n10367), .ZN(n10377) );
  XOR2_X1 U11075 ( .A(SI_17_), .B(keyinput_15), .Z(n10373) );
  XOR2_X1 U11076 ( .A(SI_16_), .B(keyinput_16), .Z(n10372) );
  XNOR2_X1 U11077 ( .A(SI_14_), .B(keyinput_18), .ZN(n10371) );
  XNOR2_X1 U11078 ( .A(SI_15_), .B(keyinput_17), .ZN(n10370) );
  NAND4_X1 U11079 ( .A1(n10373), .A2(n10372), .A3(n10371), .A4(n10370), .ZN(
        n10376) );
  XOR2_X1 U11080 ( .A(SI_12_), .B(keyinput_20), .Z(n10375) );
  XNOR2_X1 U11081 ( .A(SI_13_), .B(keyinput_19), .ZN(n10374) );
  OAI211_X1 U11082 ( .C1(n10377), .C2(n10376), .A(n10375), .B(n10374), .ZN(
        n10380) );
  XOR2_X1 U11083 ( .A(SI_11_), .B(keyinput_21), .Z(n10379) );
  XOR2_X1 U11084 ( .A(SI_10_), .B(keyinput_22), .Z(n10378) );
  AOI21_X1 U11085 ( .B1(n10380), .B2(n10379), .A(n10378), .ZN(n10383) );
  XOR2_X1 U11086 ( .A(SI_9_), .B(keyinput_23), .Z(n10382) );
  XNOR2_X1 U11087 ( .A(SI_8_), .B(keyinput_24), .ZN(n10381) );
  NOR3_X1 U11088 ( .A1(n10383), .A2(n10382), .A3(n10381), .ZN(n10386) );
  XNOR2_X1 U11089 ( .A(SI_7_), .B(keyinput_25), .ZN(n10385) );
  XNOR2_X1 U11090 ( .A(SI_6_), .B(keyinput_26), .ZN(n10384) );
  NOR3_X1 U11091 ( .A1(n10386), .A2(n10385), .A3(n10384), .ZN(n10390) );
  XOR2_X1 U11092 ( .A(SI_5_), .B(keyinput_27), .Z(n10389) );
  XOR2_X1 U11093 ( .A(SI_4_), .B(keyinput_28), .Z(n10388) );
  XOR2_X1 U11094 ( .A(SI_3_), .B(keyinput_29), .Z(n10387) );
  OAI211_X1 U11095 ( .C1(n10390), .C2(n10389), .A(n10388), .B(n10387), .ZN(
        n10393) );
  XNOR2_X1 U11096 ( .A(SI_1_), .B(keyinput_31), .ZN(n10392) );
  XNOR2_X1 U11097 ( .A(SI_2_), .B(keyinput_30), .ZN(n10391) );
  NAND3_X1 U11098 ( .A1(n10393), .A2(n10392), .A3(n10391), .ZN(n10410) );
  XOR2_X1 U11099 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput_34), .Z(n10396) );
  XNOR2_X1 U11100 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_37), .ZN(n10395)
         );
  XNOR2_X1 U11101 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_35), .ZN(n10394)
         );
  NAND3_X1 U11102 ( .A1(n10396), .A2(n10395), .A3(n10394), .ZN(n10404) );
  XNOR2_X1 U11103 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_40), .ZN(n10400)
         );
  XNOR2_X1 U11104 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_36), .ZN(n10399)
         );
  XNOR2_X1 U11105 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_39), .ZN(n10398)
         );
  XNOR2_X1 U11106 ( .A(SI_0_), .B(keyinput_32), .ZN(n10397) );
  NAND4_X1 U11107 ( .A1(n10400), .A2(n10399), .A3(n10398), .A4(n10397), .ZN(
        n10403) );
  XNOR2_X1 U11108 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_38), .ZN(n10402)
         );
  XNOR2_X1 U11109 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_33), .ZN(n10401) );
  NOR4_X1 U11110 ( .A1(n10404), .A2(n10403), .A3(n10402), .A4(n10401), .ZN(
        n10409) );
  XOR2_X1 U11111 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_43), .Z(n10407) );
  XOR2_X1 U11112 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_42), .Z(n10406) );
  XNOR2_X1 U11113 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput_41), .ZN(n10405)
         );
  NAND3_X1 U11114 ( .A1(n10407), .A2(n10406), .A3(n10405), .ZN(n10408) );
  AOI21_X1 U11115 ( .B1(n10410), .B2(n10409), .A(n10408), .ZN(n10414) );
  XOR2_X1 U11116 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_46), .Z(n10413) );
  XNOR2_X1 U11117 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_44), .ZN(n10412)
         );
  XNOR2_X1 U11118 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_45), .ZN(n10411)
         );
  NOR4_X1 U11119 ( .A1(n10414), .A2(n10413), .A3(n10412), .A4(n10411), .ZN(
        n10422) );
  XOR2_X1 U11120 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput_47), .Z(n10418) );
  XOR2_X1 U11121 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_48), .Z(n10417) );
  XNOR2_X1 U11122 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_50), .ZN(n10416)
         );
  XNOR2_X1 U11123 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput_49), .ZN(n10415)
         );
  NAND4_X1 U11124 ( .A1(n10418), .A2(n10417), .A3(n10416), .A4(n10415), .ZN(
        n10421) );
  XOR2_X1 U11125 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput_51), .Z(n10420) );
  XOR2_X1 U11126 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_52), .Z(n10419) );
  OAI211_X1 U11127 ( .C1(n10422), .C2(n10421), .A(n10420), .B(n10419), .ZN(
        n10425) );
  XNOR2_X1 U11128 ( .A(P2_REG3_REG_9__SCAN_IN), .B(keyinput_53), .ZN(n10424)
         );
  XNOR2_X1 U11129 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_54), .ZN(n10423)
         );
  AOI21_X1 U11130 ( .B1(n10425), .B2(n10424), .A(n10423), .ZN(n10428) );
  XNOR2_X1 U11131 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_55), .ZN(n10427)
         );
  XNOR2_X1 U11132 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput_56), .ZN(n10426)
         );
  OAI21_X1 U11133 ( .B1(n10428), .B2(n10427), .A(n10426), .ZN(n10431) );
  XNOR2_X1 U11134 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_57), .ZN(n10430)
         );
  XOR2_X1 U11135 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_58), .Z(n10429) );
  AOI21_X1 U11136 ( .B1(n10431), .B2(n10430), .A(n10429), .ZN(n10439) );
  XOR2_X1 U11137 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_62), .Z(n10435) );
  XOR2_X1 U11138 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_59), .Z(n10434) );
  XOR2_X1 U11139 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_61), .Z(n10433) );
  XNOR2_X1 U11140 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_60), .ZN(n10432)
         );
  NAND4_X1 U11141 ( .A1(n10435), .A2(n10434), .A3(n10433), .A4(n10432), .ZN(
        n10438) );
  XOR2_X1 U11142 ( .A(P2_REG3_REG_15__SCAN_IN), .B(keyinput_63), .Z(n10437) );
  XNOR2_X1 U11143 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_64), .ZN(n10436) );
  OAI211_X1 U11144 ( .C1(n10439), .C2(n10438), .A(n10437), .B(n10436), .ZN(
        n10446) );
  XOR2_X1 U11145 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_66), .Z(n10443)
         );
  XOR2_X1 U11146 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_65), .Z(n10442)
         );
  XOR2_X1 U11147 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_67), .Z(n10441)
         );
  XOR2_X1 U11148 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_68), .Z(n10440)
         );
  NOR4_X1 U11149 ( .A1(n10443), .A2(n10442), .A3(n10441), .A4(n10440), .ZN(
        n10445) );
  XNOR2_X1 U11150 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput_69), .ZN(n10444)
         );
  AOI21_X1 U11151 ( .B1(n10446), .B2(n10445), .A(n10444), .ZN(n10449) );
  XOR2_X1 U11152 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput_70), .Z(n10448)
         );
  XNOR2_X1 U11153 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_71), .ZN(n10447)
         );
  OAI21_X1 U11154 ( .B1(n10449), .B2(n10448), .A(n10447), .ZN(n10453) );
  XOR2_X1 U11155 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_72), .Z(n10452)
         );
  XOR2_X1 U11156 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_73), .Z(n10451)
         );
  XNOR2_X1 U11157 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_74), .ZN(n10450)
         );
  AOI211_X1 U11158 ( .C1(n10453), .C2(n10452), .A(n10451), .B(n10450), .ZN(
        n10457) );
  XNOR2_X1 U11159 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .ZN(n10456)
         );
  XOR2_X1 U11160 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .Z(n10455)
         );
  XNOR2_X1 U11161 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput_76), .ZN(n10454)
         );
  OAI211_X1 U11162 ( .C1(n10457), .C2(n10456), .A(n10455), .B(n10454), .ZN(
        n10461) );
  XOR2_X1 U11163 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .Z(n10460)
         );
  XOR2_X1 U11164 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_79), .Z(n10459)
         );
  XNOR2_X1 U11165 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput_80), .ZN(n10458)
         );
  AOI211_X1 U11166 ( .C1(n10461), .C2(n10460), .A(n10459), .B(n10458), .ZN(
        n10469) );
  XOR2_X1 U11167 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_83), .Z(n10465)
         );
  XOR2_X1 U11168 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_81), .Z(n10464)
         );
  XOR2_X1 U11169 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_82), .Z(n10463)
         );
  XNOR2_X1 U11170 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_84), .ZN(n10462)
         );
  NAND4_X1 U11171 ( .A1(n10465), .A2(n10464), .A3(n10463), .A4(n10462), .ZN(
        n10468) );
  XOR2_X1 U11172 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_86), .Z(n10467)
         );
  XNOR2_X1 U11173 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_85), .ZN(n10466)
         );
  OAI211_X1 U11174 ( .C1(n10469), .C2(n10468), .A(n10467), .B(n10466), .ZN(
        n10473) );
  XOR2_X1 U11175 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_88), .Z(n10472) );
  XOR2_X1 U11176 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .Z(n10471) );
  XOR2_X1 U11177 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_87), .Z(n10470) );
  NAND4_X1 U11178 ( .A1(n10473), .A2(n10472), .A3(n10471), .A4(n10470), .ZN(
        n10476) );
  XOR2_X1 U11179 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_91), .Z(n10475) );
  XNOR2_X1 U11180 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput_90), .ZN(n10474)
         );
  NAND3_X1 U11181 ( .A1(n10476), .A2(n10475), .A3(n10474), .ZN(n10482) );
  XOR2_X1 U11182 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_92), .Z(n10481) );
  XNOR2_X1 U11183 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_93), .ZN(n10480) );
  XNOR2_X1 U11184 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_95), .ZN(n10478) );
  XNOR2_X1 U11185 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_94), .ZN(n10477) );
  NAND2_X1 U11186 ( .A1(n10478), .A2(n10477), .ZN(n10479) );
  AOI211_X1 U11187 ( .C1(n10482), .C2(n10481), .A(n10480), .B(n10479), .ZN(
        n10484) );
  XNOR2_X1 U11188 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_96), .ZN(n10483) );
  NOR2_X1 U11189 ( .A1(n10484), .A2(n10483), .ZN(n10488) );
  XOR2_X1 U11190 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_98), .Z(n10487) );
  XNOR2_X1 U11191 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_97), .ZN(n10486) );
  XNOR2_X1 U11192 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_99), .ZN(n10485) );
  NOR4_X1 U11193 ( .A1(n10488), .A2(n10487), .A3(n10486), .A4(n10485), .ZN(
        n10491) );
  XOR2_X1 U11194 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_101), .Z(n10490) );
  XOR2_X1 U11195 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_100), .Z(n10489) );
  NOR3_X1 U11196 ( .A1(n10491), .A2(n10490), .A3(n10489), .ZN(n10494) );
  XOR2_X1 U11197 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_103), .Z(n10493) );
  XNOR2_X1 U11198 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_102), .ZN(n10492)
         );
  NOR3_X1 U11199 ( .A1(n10494), .A2(n10493), .A3(n10492), .ZN(n10498) );
  XOR2_X1 U11200 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_106), .Z(n10497) );
  XOR2_X1 U11201 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_105), .Z(n10496) );
  XOR2_X1 U11202 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_104), .Z(n10495) );
  NOR4_X1 U11203 ( .A1(n10498), .A2(n10497), .A3(n10496), .A4(n10495), .ZN(
        n10501) );
  XOR2_X1 U11204 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_108), .Z(n10500) );
  XNOR2_X1 U11205 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_107), .ZN(n10499)
         );
  NOR3_X1 U11206 ( .A1(n10501), .A2(n10500), .A3(n10499), .ZN(n10508) );
  XNOR2_X1 U11207 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_109), .ZN(n10507)
         );
  XNOR2_X1 U11208 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_112), .ZN(n10506)
         );
  XOR2_X1 U11209 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_111), .Z(n10504) );
  XOR2_X1 U11210 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_110), .Z(n10503) );
  XNOR2_X1 U11211 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_113), .ZN(n10502)
         );
  NAND3_X1 U11212 ( .A1(n10504), .A2(n10503), .A3(n10502), .ZN(n10505) );
  NOR4_X1 U11213 ( .A1(n10508), .A2(n10507), .A3(n10506), .A4(n10505), .ZN(
        n10512) );
  XNOR2_X1 U11214 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_114), .ZN(n10511)
         );
  XOR2_X1 U11215 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_116), .Z(n10510) );
  XNOR2_X1 U11216 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_115), .ZN(n10509)
         );
  OAI211_X1 U11217 ( .C1(n10512), .C2(n10511), .A(n10510), .B(n10509), .ZN(
        n10516) );
  XOR2_X1 U11218 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_119), .Z(n10515) );
  XOR2_X1 U11219 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_117), .Z(n10514) );
  XNOR2_X1 U11220 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_118), .ZN(n10513)
         );
  NAND4_X1 U11221 ( .A1(n10516), .A2(n10515), .A3(n10514), .A4(n10513), .ZN(
        n10522) );
  XOR2_X1 U11222 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_120), .Z(n10521) );
  XOR2_X1 U11223 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_122), .Z(n10519) );
  XNOR2_X1 U11224 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_121), .ZN(n10518)
         );
  XNOR2_X1 U11225 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_123), .ZN(n10517) );
  NAND3_X1 U11226 ( .A1(n10519), .A2(n10518), .A3(n10517), .ZN(n10520) );
  AOI21_X1 U11227 ( .B1(n10522), .B2(n10521), .A(n10520), .ZN(n10525) );
  XNOR2_X1 U11228 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_124), .ZN(n10524) );
  XNOR2_X1 U11229 ( .A(P1_D_REG_2__SCAN_IN), .B(keyinput_125), .ZN(n10523) );
  NOR3_X1 U11230 ( .A1(n10525), .A2(n10524), .A3(n10523), .ZN(n10527) );
  XOR2_X1 U11231 ( .A(keyinput_126), .B(P1_D_REG_3__SCAN_IN), .Z(n10526) );
  OAI22_X1 U11232 ( .A1(n10528), .A2(n10531), .B1(n10527), .B2(n10526), .ZN(
        n10529) );
  AOI21_X1 U11233 ( .B1(n10531), .B2(n10530), .A(n10529), .ZN(n10532) );
  XOR2_X1 U11234 ( .A(n10533), .B(n10532), .Z(P1_U3542) );
  AOI22_X1 U11235 ( .A1(n10535), .A2(n10981), .B1(n10873), .B2(n10534), .ZN(
        n10536) );
  OAI211_X1 U11236 ( .C1(n10539), .C2(n10538), .A(n10537), .B(n10536), .ZN(
        n10560) );
  MUX2_X1 U11237 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10560), .S(n10989), .Z(
        P1_U3541) );
  INV_X1 U11238 ( .A(n10540), .ZN(n10545) );
  AOI22_X1 U11239 ( .A1(n10542), .A2(n10981), .B1(n10873), .B2(n10541), .ZN(
        n10543) );
  OAI211_X1 U11240 ( .C1(n10545), .C2(n10875), .A(n10544), .B(n10543), .ZN(
        n10561) );
  MUX2_X1 U11241 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10561), .S(n10989), .Z(
        P1_U3540) );
  MUX2_X1 U11242 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n10546), .S(n10989), .Z(
        P1_U3523) );
  MUX2_X1 U11243 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10548), .S(n10993), .Z(
        P1_U3521) );
  MUX2_X1 U11244 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10549), .S(n10993), .Z(
        P1_U3520) );
  MUX2_X1 U11245 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10551), .S(n10993), .Z(
        P1_U3518) );
  MUX2_X1 U11246 ( .A(n10552), .B(P1_REG0_REG_26__SCAN_IN), .S(n10990), .Z(
        P1_U3517) );
  MUX2_X1 U11247 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10553), .S(n10993), .Z(
        P1_U3516) );
  MUX2_X1 U11248 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10554), .S(n10993), .Z(
        P1_U3515) );
  MUX2_X1 U11249 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10555), .S(n10993), .Z(
        P1_U3514) );
  MUX2_X1 U11250 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10556), .S(n10993), .Z(
        P1_U3513) );
  MUX2_X1 U11251 ( .A(n10557), .B(P1_REG0_REG_21__SCAN_IN), .S(n10990), .Z(
        P1_U3512) );
  MUX2_X1 U11252 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10558), .S(n10993), .Z(
        P1_U3511) );
  MUX2_X1 U11253 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10559), .S(n10993), .Z(
        P1_U3510) );
  MUX2_X1 U11254 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10560), .S(n10993), .Z(
        P1_U3508) );
  MUX2_X1 U11255 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10561), .S(n10993), .Z(
        P1_U3505) );
  MUX2_X1 U11256 ( .A(n10562), .B(P1_D_REG_0__SCAN_IN), .S(n10580), .Z(
        P1_U3440) );
  NOR4_X1 U11257 ( .A1(n6813), .A2(P1_IR_REG_30__SCAN_IN), .A3(n10563), .A4(
        P1_U3084), .ZN(n10564) );
  AOI21_X1 U11258 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n10571), .A(n10564), 
        .ZN(n10565) );
  OAI21_X1 U11259 ( .B1(n10566), .B2(n5044), .A(n10565), .ZN(P1_U3322) );
  OAI222_X1 U11260 ( .A1(n5044), .A2(n10569), .B1(n10568), .B2(P1_U3084), .C1(
        n10567), .C2(n10575), .ZN(P1_U3323) );
  AOI21_X1 U11261 ( .B1(n10571), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n10570), 
        .ZN(n10572) );
  OAI21_X1 U11262 ( .B1(n10573), .B2(n5044), .A(n10572), .ZN(P1_U3326) );
  INV_X1 U11263 ( .A(n10574), .ZN(n10578) );
  OAI222_X1 U11264 ( .A1(n10578), .A2(P1_U3084), .B1(n5044), .B2(n10577), .C1(
        n10576), .C2(n10575), .ZN(P1_U3327) );
  MUX2_X1 U11265 ( .A(n10579), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NOR2_X1 U11266 ( .A1(n10581), .A2(n10580), .ZN(n10605) );
  NOR2_X1 U11267 ( .A1(n10612), .A2(n10582), .ZN(P1_U3321) );
  NOR2_X1 U11268 ( .A1(n10612), .A2(n10583), .ZN(P1_U3320) );
  NOR2_X1 U11269 ( .A1(n10612), .A2(n10531), .ZN(P1_U3319) );
  INV_X1 U11270 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10584) );
  NOR2_X1 U11271 ( .A1(n10612), .A2(n10584), .ZN(P1_U3318) );
  INV_X1 U11272 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10585) );
  NOR2_X1 U11273 ( .A1(n10612), .A2(n10585), .ZN(P1_U3317) );
  INV_X1 U11274 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10586) );
  NOR2_X1 U11275 ( .A1(n10612), .A2(n10586), .ZN(P1_U3316) );
  INV_X1 U11276 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10587) );
  NOR2_X1 U11277 ( .A1(n10612), .A2(n10587), .ZN(P1_U3315) );
  INV_X1 U11278 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10588) );
  NOR2_X1 U11279 ( .A1(n10612), .A2(n10588), .ZN(P1_U3314) );
  INV_X1 U11280 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10589) );
  NOR2_X1 U11281 ( .A1(n10612), .A2(n10589), .ZN(P1_U3313) );
  INV_X1 U11282 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10590) );
  NOR2_X1 U11283 ( .A1(n10612), .A2(n10590), .ZN(P1_U3312) );
  INV_X1 U11284 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10591) );
  NOR2_X1 U11285 ( .A1(n10612), .A2(n10591), .ZN(P1_U3311) );
  INV_X1 U11286 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10592) );
  NOR2_X1 U11287 ( .A1(n10605), .A2(n10592), .ZN(P1_U3310) );
  INV_X1 U11288 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10593) );
  NOR2_X1 U11289 ( .A1(n10605), .A2(n10593), .ZN(P1_U3309) );
  INV_X1 U11290 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10594) );
  NOR2_X1 U11291 ( .A1(n10605), .A2(n10594), .ZN(P1_U3308) );
  INV_X1 U11292 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10595) );
  NOR2_X1 U11293 ( .A1(n10605), .A2(n10595), .ZN(P1_U3307) );
  INV_X1 U11294 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10596) );
  NOR2_X1 U11295 ( .A1(n10605), .A2(n10596), .ZN(P1_U3306) );
  INV_X1 U11296 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10597) );
  NOR2_X1 U11297 ( .A1(n10605), .A2(n10597), .ZN(P1_U3305) );
  INV_X1 U11298 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10598) );
  NOR2_X1 U11299 ( .A1(n10605), .A2(n10598), .ZN(P1_U3304) );
  INV_X1 U11300 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10599) );
  NOR2_X1 U11301 ( .A1(n10612), .A2(n10599), .ZN(P1_U3303) );
  INV_X1 U11302 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10600) );
  NOR2_X1 U11303 ( .A1(n10612), .A2(n10600), .ZN(P1_U3302) );
  INV_X1 U11304 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10601) );
  NOR2_X1 U11305 ( .A1(n10605), .A2(n10601), .ZN(P1_U3301) );
  INV_X1 U11306 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10602) );
  NOR2_X1 U11307 ( .A1(n10605), .A2(n10602), .ZN(P1_U3300) );
  INV_X1 U11308 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10603) );
  NOR2_X1 U11309 ( .A1(n10605), .A2(n10603), .ZN(P1_U3299) );
  INV_X1 U11310 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10604) );
  NOR2_X1 U11311 ( .A1(n10605), .A2(n10604), .ZN(P1_U3298) );
  INV_X1 U11312 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10606) );
  NOR2_X1 U11313 ( .A1(n10612), .A2(n10606), .ZN(P1_U3297) );
  INV_X1 U11314 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10607) );
  NOR2_X1 U11315 ( .A1(n10612), .A2(n10607), .ZN(P1_U3296) );
  INV_X1 U11316 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10608) );
  NOR2_X1 U11317 ( .A1(n10612), .A2(n10608), .ZN(P1_U3295) );
  INV_X1 U11318 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10609) );
  NOR2_X1 U11319 ( .A1(n10612), .A2(n10609), .ZN(P1_U3294) );
  NOR2_X1 U11320 ( .A1(n10612), .A2(n10610), .ZN(P1_U3293) );
  NOR2_X1 U11321 ( .A1(n10612), .A2(n10611), .ZN(P1_U3292) );
  NAND2_X1 U11322 ( .A1(n10614), .A2(n10613), .ZN(n10692) );
  AOI22_X1 U11323 ( .A1(n10616), .A2(n10694), .B1(n10615), .B2(n10692), .ZN(
        P2_U3438) );
  AND2_X1 U11324 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10692), .ZN(P2_U3326) );
  AND2_X1 U11325 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10692), .ZN(P2_U3325) );
  AND2_X1 U11326 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10692), .ZN(P2_U3324) );
  AND2_X1 U11327 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10692), .ZN(P2_U3323) );
  AND2_X1 U11328 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10692), .ZN(P2_U3322) );
  AND2_X1 U11329 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10692), .ZN(P2_U3321) );
  AND2_X1 U11330 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10692), .ZN(P2_U3320) );
  AND2_X1 U11331 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10692), .ZN(P2_U3319) );
  AND2_X1 U11332 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10692), .ZN(P2_U3318) );
  AND2_X1 U11333 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10692), .ZN(P2_U3317) );
  AND2_X1 U11334 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10692), .ZN(P2_U3316) );
  AND2_X1 U11335 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10692), .ZN(P2_U3315) );
  AND2_X1 U11336 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10692), .ZN(P2_U3314) );
  AND2_X1 U11337 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10692), .ZN(P2_U3313) );
  AND2_X1 U11338 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10692), .ZN(P2_U3312) );
  AND2_X1 U11339 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10692), .ZN(P2_U3311) );
  AND2_X1 U11340 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10692), .ZN(P2_U3310) );
  AND2_X1 U11341 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10692), .ZN(P2_U3309) );
  AND2_X1 U11342 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10692), .ZN(P2_U3308) );
  AND2_X1 U11343 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10692), .ZN(P2_U3307) );
  AND2_X1 U11344 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10692), .ZN(P2_U3306) );
  AND2_X1 U11345 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10692), .ZN(P2_U3305) );
  AND2_X1 U11346 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10692), .ZN(P2_U3304) );
  AND2_X1 U11347 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10692), .ZN(P2_U3303) );
  AND2_X1 U11348 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10692), .ZN(P2_U3302) );
  AND2_X1 U11349 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10692), .ZN(P2_U3301) );
  AND2_X1 U11350 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10692), .ZN(P2_U3300) );
  AND2_X1 U11351 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10692), .ZN(P2_U3299) );
  AND2_X1 U11352 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10692), .ZN(P2_U3298) );
  AND2_X1 U11353 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10692), .ZN(P2_U3297) );
  XOR2_X1 U11354 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  INV_X1 U11355 ( .A(n10617), .ZN(n10618) );
  NAND2_X1 U11356 ( .A1(n10619), .A2(n10618), .ZN(n10620) );
  XOR2_X1 U11357 ( .A(n10621), .B(n10620), .Z(ADD_1071_U5) );
  XOR2_X1 U11358 ( .A(n10623), .B(n10622), .Z(ADD_1071_U54) );
  XOR2_X1 U11359 ( .A(n10625), .B(n10624), .Z(ADD_1071_U53) );
  XNOR2_X1 U11360 ( .A(n10627), .B(n10626), .ZN(ADD_1071_U52) );
  NOR2_X1 U11361 ( .A1(n10629), .A2(n10628), .ZN(n10630) );
  XOR2_X1 U11362 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n10630), .Z(ADD_1071_U51) );
  XOR2_X1 U11363 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10631), .Z(ADD_1071_U50) );
  XOR2_X1 U11364 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10632), .Z(ADD_1071_U49) );
  XOR2_X1 U11365 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10633), .Z(ADD_1071_U48) );
  XOR2_X1 U11366 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n10634), .Z(ADD_1071_U47) );
  XOR2_X1 U11367 ( .A(n10636), .B(n10635), .Z(ADD_1071_U63) );
  XOR2_X1 U11368 ( .A(n10638), .B(n10637), .Z(ADD_1071_U62) );
  XNOR2_X1 U11369 ( .A(n10640), .B(n10639), .ZN(ADD_1071_U61) );
  XNOR2_X1 U11370 ( .A(n10642), .B(n10641), .ZN(ADD_1071_U60) );
  XNOR2_X1 U11371 ( .A(n10644), .B(n10643), .ZN(ADD_1071_U59) );
  XNOR2_X1 U11372 ( .A(n10646), .B(n10645), .ZN(ADD_1071_U58) );
  XNOR2_X1 U11373 ( .A(n10648), .B(n10647), .ZN(ADD_1071_U57) );
  XNOR2_X1 U11374 ( .A(n10650), .B(n10649), .ZN(ADD_1071_U56) );
  NOR2_X1 U11375 ( .A1(n10652), .A2(n10651), .ZN(n10653) );
  XOR2_X1 U11376 ( .A(P1_ADDR_REG_18__SCAN_IN), .B(n10653), .Z(ADD_1071_U55)
         );
  INV_X1 U11377 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10740) );
  AOI21_X1 U11378 ( .B1(n5050), .B2(n10655), .A(n10654), .ZN(n10657) );
  XNOR2_X1 U11379 ( .A(n10657), .B(n10656), .ZN(n10658) );
  AOI22_X1 U11380 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n10679), .B1(n10659), 
        .B2(n10658), .ZN(n10660) );
  OAI21_X1 U11381 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n10740), .A(n10660), .ZN(
        P1_U3241) );
  AOI22_X1 U11382 ( .A1(n10679), .A2(P1_ADDR_REG_10__SCAN_IN), .B1(n10662), 
        .B2(n10661), .ZN(n10674) );
  OAI21_X1 U11383 ( .B1(n10665), .B2(n10664), .A(n10663), .ZN(n10667) );
  NAND2_X1 U11384 ( .A1(n10667), .A2(n10666), .ZN(n10672) );
  OAI211_X1 U11385 ( .C1(n10670), .C2(n10669), .A(n10681), .B(n10668), .ZN(
        n10671) );
  NAND4_X1 U11386 ( .A1(n10674), .A2(n10673), .A3(n10672), .A4(n10671), .ZN(
        P1_U3251) );
  OAI22_X1 U11387 ( .A1(n10677), .A2(n10676), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10675), .ZN(n10678) );
  AOI21_X1 U11388 ( .B1(n10679), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n10678), .ZN(
        n10691) );
  AND2_X1 U11389 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10683) );
  OAI211_X1 U11390 ( .C1(n10683), .C2(n10682), .A(n10681), .B(n10680), .ZN(
        n10690) );
  AOI211_X1 U11391 ( .C1(n10687), .C2(n10686), .A(n10685), .B(n10684), .ZN(
        n10688) );
  INV_X1 U11392 ( .A(n10688), .ZN(n10689) );
  NAND3_X1 U11393 ( .A1(n10691), .A2(n10690), .A3(n10689), .ZN(P1_U3242) );
  INV_X1 U11394 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10693) );
  AOI22_X1 U11395 ( .A1(n10695), .A2(n10694), .B1(n10693), .B2(n10692), .ZN(
        P2_U3437) );
  AOI22_X1 U11396 ( .A1(n10696), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10726), .ZN(n10702) );
  INV_X1 U11397 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10697) );
  NAND2_X1 U11398 ( .A1(n10726), .A2(n10697), .ZN(n10698) );
  OAI211_X1 U11399 ( .C1(n10719), .C2(P2_REG2_REG_0__SCAN_IN), .A(n10698), .B(
        n10710), .ZN(n10699) );
  INV_X1 U11400 ( .A(n10699), .ZN(n10701) );
  AOI22_X1 U11401 ( .A1(n10718), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10700) );
  OAI221_X1 U11402 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n10702), .C1(n5709), .C2(
        n10701), .A(n10700), .ZN(P2_U3245) );
  NAND2_X1 U11403 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10703) );
  AND2_X1 U11404 ( .A1(n10704), .A2(n10703), .ZN(n10706) );
  OR3_X1 U11405 ( .A1(n10719), .A2(n10706), .A3(n10705), .ZN(n10708) );
  AOI22_X1 U11406 ( .A1(n10718), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n10707) );
  OAI211_X1 U11407 ( .C1(n10710), .C2(n10709), .A(n10708), .B(n10707), .ZN(
        n10711) );
  INV_X1 U11408 ( .A(n10711), .ZN(n10716) );
  NOR2_X1 U11409 ( .A1(n5709), .A2(n10697), .ZN(n10714) );
  OAI211_X1 U11410 ( .C1(n10714), .C2(n10713), .A(n10726), .B(n10712), .ZN(
        n10715) );
  NAND2_X1 U11411 ( .A1(n10716), .A2(n10715), .ZN(P2_U3246) );
  AOI22_X1 U11412 ( .A1(n10718), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n10731) );
  AOI21_X1 U11413 ( .B1(n10724), .B2(n10723), .A(n10722), .ZN(n10730) );
  OAI211_X1 U11414 ( .C1(n10728), .C2(n10727), .A(n10726), .B(n10725), .ZN(
        n10729) );
  NAND3_X1 U11415 ( .A1(n10731), .A2(n10730), .A3(n10729), .ZN(P2_U3247) );
  XNOR2_X1 U11416 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  AOI21_X1 U11417 ( .B1(n10734), .B2(n10733), .A(n10732), .ZN(n10737) );
  NOR2_X1 U11418 ( .A1(n10735), .A2(n11006), .ZN(n10736) );
  AOI211_X1 U11419 ( .C1(n10738), .C2(P1_REG2_REG_0__SCAN_IN), .A(n10737), .B(
        n10736), .ZN(n10739) );
  OAI21_X1 U11420 ( .B1(n10741), .B2(n10740), .A(n10739), .ZN(P1_U3291) );
  AOI22_X1 U11421 ( .A1(n10743), .A2(n10936), .B1(n5698), .B2(n10742), .ZN(
        n10744) );
  AND2_X1 U11422 ( .A1(n10745), .A2(n10744), .ZN(n10747) );
  AOI22_X1 U11423 ( .A1(n10811), .A2(n10747), .B1(n10697), .B2(n10945), .ZN(
        P2_U3520) );
  INV_X1 U11424 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10746) );
  AOI22_X1 U11425 ( .A1(n10950), .A2(n10747), .B1(n10746), .B2(n10947), .ZN(
        P2_U3451) );
  INV_X1 U11426 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10748) );
  AOI22_X1 U11427 ( .A1(n10993), .A2(n10749), .B1(n10748), .B2(n10990), .ZN(
        P1_U3460) );
  INV_X1 U11428 ( .A(n10750), .ZN(n10888) );
  INV_X1 U11429 ( .A(n10751), .ZN(n10753) );
  OAI22_X1 U11430 ( .A1(n10753), .A2(n10921), .B1(n10752), .B2(n10919), .ZN(
        n10755) );
  AOI211_X1 U11431 ( .C1(n10888), .C2(n10756), .A(n10755), .B(n10754), .ZN(
        n10758) );
  AOI22_X1 U11432 ( .A1(n10811), .A2(n10758), .B1(n7005), .B2(n10945), .ZN(
        P2_U3522) );
  INV_X1 U11433 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10757) );
  AOI22_X1 U11434 ( .A1(n10950), .A2(n10758), .B1(n10757), .B2(n10947), .ZN(
        P2_U3457) );
  OAI22_X1 U11435 ( .A1(n10760), .A2(n10921), .B1(n10759), .B2(n10919), .ZN(
        n10763) );
  INV_X1 U11436 ( .A(n10761), .ZN(n10762) );
  AOI211_X1 U11437 ( .C1(n10936), .C2(n10764), .A(n10763), .B(n10762), .ZN(
        n10766) );
  AOI22_X1 U11438 ( .A1(n10811), .A2(n10766), .B1(n7004), .B2(n10945), .ZN(
        P2_U3523) );
  INV_X1 U11439 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10765) );
  AOI22_X1 U11440 ( .A1(n10950), .A2(n10766), .B1(n10765), .B2(n10947), .ZN(
        P2_U3460) );
  OAI22_X1 U11441 ( .A1(n10768), .A2(n10960), .B1(n10767), .B2(n10984), .ZN(
        n10770) );
  AOI211_X1 U11442 ( .C1(n10933), .C2(n10771), .A(n10770), .B(n10769), .ZN(
        n10773) );
  AOI22_X1 U11443 ( .A1(n10989), .A2(n10773), .B1(n6761), .B2(n10987), .ZN(
        P1_U3527) );
  INV_X1 U11444 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U11445 ( .A1(n10993), .A2(n10773), .B1(n10772), .B2(n10990), .ZN(
        P1_U3466) );
  INV_X1 U11446 ( .A(n10774), .ZN(n10776) );
  OAI22_X1 U11447 ( .A1(n10776), .A2(n10921), .B1(n10775), .B2(n10919), .ZN(
        n10778) );
  AOI211_X1 U11448 ( .C1(n10936), .C2(n10779), .A(n10778), .B(n10777), .ZN(
        n10781) );
  AOI22_X1 U11449 ( .A1(n10811), .A2(n10781), .B1(n7002), .B2(n10945), .ZN(
        P2_U3524) );
  INV_X1 U11450 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10780) );
  AOI22_X1 U11451 ( .A1(n10950), .A2(n10781), .B1(n10780), .B2(n10947), .ZN(
        P2_U3463) );
  INV_X1 U11452 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10805) );
  XNOR2_X1 U11453 ( .A(n10782), .B(n10787), .ZN(n10810) );
  NAND2_X1 U11454 ( .A1(n10783), .A2(n10795), .ZN(n10784) );
  NAND2_X1 U11455 ( .A1(n10784), .A2(n10940), .ZN(n10785) );
  OR2_X1 U11456 ( .A1(n10786), .A2(n10785), .ZN(n10806) );
  XNOR2_X1 U11457 ( .A(n10788), .B(n10787), .ZN(n10793) );
  AOI222_X1 U11458 ( .A1(n10794), .A2(n10793), .B1(n10792), .B2(n10791), .C1(
        n10790), .C2(n10789), .ZN(n10807) );
  AOI22_X1 U11459 ( .A1(n10798), .A2(n10797), .B1(n10796), .B2(n10795), .ZN(
        n10799) );
  OAI211_X1 U11460 ( .C1(n10800), .C2(n10806), .A(n10807), .B(n10799), .ZN(
        n10801) );
  AOI21_X1 U11461 ( .B1(n10802), .B2(n10810), .A(n10801), .ZN(n10804) );
  AOI22_X1 U11462 ( .A1(n7664), .A2(n10805), .B1(n10804), .B2(n10803), .ZN(
        P2_U3291) );
  OAI211_X1 U11463 ( .C1(n10808), .C2(n10919), .A(n10807), .B(n10806), .ZN(
        n10809) );
  AOI21_X1 U11464 ( .B1(n10936), .B2(n10810), .A(n10809), .ZN(n10813) );
  AOI22_X1 U11465 ( .A1(n10811), .A2(n10813), .B1(n7000), .B2(n10945), .ZN(
        P2_U3525) );
  INV_X1 U11466 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10812) );
  AOI22_X1 U11467 ( .A1(n10950), .A2(n10813), .B1(n10812), .B2(n10947), .ZN(
        P2_U3466) );
  OAI22_X1 U11468 ( .A1(n10815), .A2(n10960), .B1(n10814), .B2(n10984), .ZN(
        n10817) );
  AOI211_X1 U11469 ( .C1(n10933), .C2(n10818), .A(n10817), .B(n10816), .ZN(
        n10820) );
  AOI22_X1 U11470 ( .A1(n10989), .A2(n10820), .B1(n6757), .B2(n10987), .ZN(
        P1_U3529) );
  INV_X1 U11471 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10819) );
  AOI22_X1 U11472 ( .A1(n10993), .A2(n10820), .B1(n10819), .B2(n10990), .ZN(
        P1_U3472) );
  AOI22_X1 U11473 ( .A1(n10822), .A2(n10940), .B1(n10939), .B2(n10821), .ZN(
        n10825) );
  NAND3_X1 U11474 ( .A1(n9569), .A2(n10823), .A3(n10936), .ZN(n10824) );
  AND3_X1 U11475 ( .A1(n10826), .A2(n10825), .A3(n10824), .ZN(n10829) );
  AOI22_X1 U11476 ( .A1(n10811), .A2(n10829), .B1(n10827), .B2(n10945), .ZN(
        P2_U3526) );
  INV_X1 U11477 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10828) );
  AOI22_X1 U11478 ( .A1(n10950), .A2(n10829), .B1(n10828), .B2(n10947), .ZN(
        P2_U3469) );
  OAI22_X1 U11479 ( .A1(n10831), .A2(n10921), .B1(n10830), .B2(n10919), .ZN(
        n10833) );
  AOI211_X1 U11480 ( .C1(n10936), .C2(n10834), .A(n10833), .B(n10832), .ZN(
        n10836) );
  AOI22_X1 U11481 ( .A1(n10811), .A2(n10836), .B1(n7011), .B2(n10945), .ZN(
        P2_U3527) );
  INV_X1 U11482 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10835) );
  AOI22_X1 U11483 ( .A1(n10950), .A2(n10836), .B1(n10835), .B2(n10947), .ZN(
        P2_U3472) );
  AOI22_X1 U11484 ( .A1(n10838), .A2(n10981), .B1(n10873), .B2(n10837), .ZN(
        n10839) );
  OAI211_X1 U11485 ( .C1(n10875), .C2(n10841), .A(n10840), .B(n10839), .ZN(
        n10842) );
  INV_X1 U11486 ( .A(n10842), .ZN(n10844) );
  AOI22_X1 U11487 ( .A1(n10989), .A2(n10844), .B1(n6765), .B2(n10987), .ZN(
        P1_U3531) );
  INV_X1 U11488 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10843) );
  AOI22_X1 U11489 ( .A1(n10993), .A2(n10844), .B1(n10843), .B2(n10990), .ZN(
        P1_U3478) );
  NAND3_X1 U11490 ( .A1(n10846), .A2(n10845), .A3(n10936), .ZN(n10848) );
  OAI211_X1 U11491 ( .C1(n10849), .C2(n10919), .A(n10848), .B(n10847), .ZN(
        n10850) );
  NOR2_X1 U11492 ( .A1(n10851), .A2(n10850), .ZN(n10853) );
  AOI22_X1 U11493 ( .A1(n10811), .A2(n10853), .B1(n7092), .B2(n10945), .ZN(
        P2_U3528) );
  INV_X1 U11494 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10852) );
  AOI22_X1 U11495 ( .A1(n10950), .A2(n10853), .B1(n10852), .B2(n10947), .ZN(
        P2_U3475) );
  OAI22_X1 U11496 ( .A1(n10855), .A2(n10960), .B1(n10854), .B2(n10984), .ZN(
        n10857) );
  AOI211_X1 U11497 ( .C1(n10933), .C2(n10858), .A(n10857), .B(n10856), .ZN(
        n10861) );
  AOI22_X1 U11498 ( .A1(n10989), .A2(n10861), .B1(n10859), .B2(n10987), .ZN(
        P1_U3532) );
  INV_X1 U11499 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10860) );
  AOI22_X1 U11500 ( .A1(n10993), .A2(n10861), .B1(n10860), .B2(n10990), .ZN(
        P1_U3481) );
  INV_X1 U11501 ( .A(n10862), .ZN(n10867) );
  OAI22_X1 U11502 ( .A1(n10864), .A2(n10921), .B1(n5301), .B2(n10919), .ZN(
        n10866) );
  AOI211_X1 U11503 ( .C1(n10888), .C2(n10867), .A(n10866), .B(n10865), .ZN(
        n10869) );
  AOI22_X1 U11504 ( .A1(n10811), .A2(n10869), .B1(n7229), .B2(n10945), .ZN(
        P2_U3529) );
  INV_X1 U11505 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10868) );
  AOI22_X1 U11506 ( .A1(n10950), .A2(n10869), .B1(n10868), .B2(n10947), .ZN(
        P2_U3478) );
  INV_X1 U11507 ( .A(n10876), .ZN(n10878) );
  AOI211_X1 U11508 ( .C1(n10873), .C2(n10872), .A(n10871), .B(n10870), .ZN(
        n10874) );
  OAI21_X1 U11509 ( .B1(n10876), .B2(n10875), .A(n10874), .ZN(n10877) );
  AOI21_X1 U11510 ( .B1(n10879), .B2(n10878), .A(n10877), .ZN(n10882) );
  AOI22_X1 U11511 ( .A1(n10989), .A2(n10882), .B1(n10880), .B2(n10987), .ZN(
        P1_U3533) );
  INV_X1 U11512 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10881) );
  AOI22_X1 U11513 ( .A1(n10993), .A2(n10882), .B1(n10881), .B2(n10990), .ZN(
        P1_U3484) );
  INV_X1 U11514 ( .A(n10883), .ZN(n10887) );
  OAI22_X1 U11515 ( .A1(n10884), .A2(n10921), .B1(n5299), .B2(n10919), .ZN(
        n10886) );
  AOI211_X1 U11516 ( .C1(n10888), .C2(n10887), .A(n10886), .B(n10885), .ZN(
        n10890) );
  AOI22_X1 U11517 ( .A1(n10811), .A2(n10890), .B1(n7385), .B2(n10945), .ZN(
        P2_U3530) );
  INV_X1 U11518 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10889) );
  AOI22_X1 U11519 ( .A1(n10950), .A2(n10890), .B1(n10889), .B2(n10947), .ZN(
        P2_U3481) );
  OAI22_X1 U11520 ( .A1(n10892), .A2(n10960), .B1(n10891), .B2(n10984), .ZN(
        n10893) );
  AOI21_X1 U11521 ( .B1(n10894), .B2(n10933), .A(n10893), .ZN(n10895) );
  AND2_X1 U11522 ( .A1(n10896), .A2(n10895), .ZN(n10899) );
  AOI22_X1 U11523 ( .A1(n10989), .A2(n10899), .B1(n10897), .B2(n10987), .ZN(
        P1_U3534) );
  INV_X1 U11524 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10898) );
  AOI22_X1 U11525 ( .A1(n10993), .A2(n10899), .B1(n10898), .B2(n10990), .ZN(
        P1_U3487) );
  AOI21_X1 U11526 ( .B1(n10939), .B2(n10901), .A(n10900), .ZN(n10902) );
  OAI211_X1 U11527 ( .C1(n10905), .C2(n10904), .A(n10903), .B(n10902), .ZN(
        n10906) );
  INV_X1 U11528 ( .A(n10906), .ZN(n10909) );
  AOI22_X1 U11529 ( .A1(n10811), .A2(n10909), .B1(n10907), .B2(n10945), .ZN(
        P2_U3531) );
  INV_X1 U11530 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10908) );
  AOI22_X1 U11531 ( .A1(n10950), .A2(n10909), .B1(n10908), .B2(n10947), .ZN(
        P2_U3484) );
  OAI211_X1 U11532 ( .C1(n10912), .C2(n10984), .A(n10911), .B(n10910), .ZN(
        n10915) );
  NOR2_X1 U11533 ( .A1(n10913), .A2(n7169), .ZN(n10914) );
  AOI211_X1 U11534 ( .C1(n10916), .C2(n10933), .A(n10915), .B(n10914), .ZN(
        n10918) );
  AOI22_X1 U11535 ( .A1(n10989), .A2(n10918), .B1(n6771), .B2(n10987), .ZN(
        P1_U3535) );
  INV_X1 U11536 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U11537 ( .A1(n10993), .A2(n10918), .B1(n10917), .B2(n10990), .ZN(
        P1_U3490) );
  OAI22_X1 U11538 ( .A1(n10922), .A2(n10921), .B1(n10920), .B2(n10919), .ZN(
        n10923) );
  AOI211_X1 U11539 ( .C1(n10925), .C2(n10936), .A(n10924), .B(n10923), .ZN(
        n10927) );
  AOI22_X1 U11540 ( .A1(n10811), .A2(n10927), .B1(n7787), .B2(n10945), .ZN(
        P2_U3532) );
  INV_X1 U11541 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10926) );
  AOI22_X1 U11542 ( .A1(n10950), .A2(n10927), .B1(n10926), .B2(n10947), .ZN(
        P2_U3487) );
  OAI22_X1 U11543 ( .A1(n10929), .A2(n10960), .B1(n5312), .B2(n10984), .ZN(
        n10931) );
  AOI211_X1 U11544 ( .C1(n10933), .C2(n10932), .A(n10931), .B(n10930), .ZN(
        n10935) );
  AOI22_X1 U11545 ( .A1(n10989), .A2(n10935), .B1(n6756), .B2(n10987), .ZN(
        P1_U3536) );
  INV_X1 U11546 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10934) );
  AOI22_X1 U11547 ( .A1(n10993), .A2(n10935), .B1(n10934), .B2(n10990), .ZN(
        P1_U3493) );
  NAND3_X1 U11548 ( .A1(n10937), .A2(n10936), .A3(n8357), .ZN(n10944) );
  AOI22_X1 U11549 ( .A1(n10941), .A2(n10940), .B1(n10939), .B2(n10938), .ZN(
        n10942) );
  AOI22_X1 U11550 ( .A1(n10811), .A2(n10949), .B1(n10946), .B2(n10945), .ZN(
        P2_U3533) );
  INV_X1 U11551 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10948) );
  AOI22_X1 U11552 ( .A1(n10950), .A2(n10949), .B1(n10948), .B2(n10947), .ZN(
        P2_U3490) );
  OAI21_X1 U11553 ( .B1(n10952), .B2(n10984), .A(n10951), .ZN(n10953) );
  AOI211_X1 U11554 ( .C1(n10955), .C2(n5587), .A(n10954), .B(n10953), .ZN(
        n10958) );
  INV_X1 U11555 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10956) );
  AOI22_X1 U11556 ( .A1(n10989), .A2(n10958), .B1(n10956), .B2(n10987), .ZN(
        P1_U3537) );
  INV_X1 U11557 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10957) );
  AOI22_X1 U11558 ( .A1(n10993), .A2(n10958), .B1(n10957), .B2(n10990), .ZN(
        P1_U3496) );
  OAI22_X1 U11559 ( .A1(n10961), .A2(n10960), .B1(n10959), .B2(n10984), .ZN(
        n10962) );
  AOI211_X1 U11560 ( .C1(n10964), .C2(n5587), .A(n10963), .B(n10962), .ZN(
        n10967) );
  AOI22_X1 U11561 ( .A1(n10989), .A2(n10967), .B1(n10965), .B2(n10987), .ZN(
        P1_U3538) );
  INV_X1 U11562 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10966) );
  AOI22_X1 U11563 ( .A1(n10993), .A2(n10967), .B1(n10966), .B2(n10990), .ZN(
        P1_U3499) );
  OAI21_X1 U11564 ( .B1(n10970), .B2(n10969), .A(n10968), .ZN(n10971) );
  INV_X1 U11565 ( .A(n10971), .ZN(n11002) );
  OAI21_X1 U11566 ( .B1(n10974), .B2(n10973), .A(n10972), .ZN(n10979) );
  AOI222_X1 U11567 ( .A1(n10980), .A2(n10979), .B1(n10978), .B2(n10977), .C1(
        n10976), .C2(n10975), .ZN(n11005) );
  OAI211_X1 U11568 ( .C1(n10983), .C2(n10985), .A(n10982), .B(n10981), .ZN(
        n10998) );
  OAI211_X1 U11569 ( .C1(n10985), .C2(n10984), .A(n11005), .B(n10998), .ZN(
        n10986) );
  AOI21_X1 U11570 ( .B1(n11002), .B2(n5587), .A(n10986), .ZN(n10992) );
  INV_X1 U11571 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10988) );
  AOI22_X1 U11572 ( .A1(n10989), .A2(n10992), .B1(n10988), .B2(n10987), .ZN(
        P1_U3539) );
  INV_X1 U11573 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10991) );
  AOI22_X1 U11574 ( .A1(n10993), .A2(n10992), .B1(n10991), .B2(n10990), .ZN(
        P1_U3502) );
  AOI222_X1 U11575 ( .A1(n10997), .A2(n10996), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(n10738), .C1(n10995), .C2(n10994), .ZN(n11004) );
  INV_X1 U11576 ( .A(n10998), .ZN(n11000) );
  AOI22_X1 U11577 ( .A1(n11002), .A2(n11001), .B1(n11000), .B2(n10999), .ZN(
        n11003) );
  OAI211_X1 U11578 ( .C1(n11006), .C2(n11005), .A(n11004), .B(n11003), .ZN(
        P1_U3275) );
  XNOR2_X1 U11579 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U5143 ( .A(n7681), .ZN(n10759) );
  CLKBUF_X2 U5190 ( .A(n5703), .Z(n7012) );
  CLKBUF_X1 U5335 ( .A(n7113), .Z(n7510) );
endmodule

