

module b20_C_gen_AntiSAT_k_256_5 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, 
        keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, 
        keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, 
        keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, 
        keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, 
        keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, 
        keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, 
        keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, 
        keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104, 
        keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108, 
        keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112, 
        keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116, 
        keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120, 
        keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124, 
        keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, 
        keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, 
        keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, 
        keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, 
        keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, 
        keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, 
        keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, 
        keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562;

  AOI21_X2 U5013 ( .B1(n8094), .B2(n8093), .A(n8092), .ZN(n9143) );
  AOI21_X1 U5014 ( .B1(n9051), .B2(n8090), .A(n8087), .ZN(n9141) );
  INV_X1 U5015 ( .A(n9418), .ZN(n9658) );
  NAND2_X1 U5016 ( .A1(n5629), .A2(n5628), .ZN(n9612) );
  INV_X2 U5017 ( .A(n8356), .ZN(n6915) );
  CLKBUF_X2 U5018 ( .A(n5909), .Z(n7094) );
  OR2_X1 U5019 ( .A1(n5315), .A2(n5282), .ZN(n5334) );
  INV_X1 U5020 ( .A(n5850), .ZN(n9007) );
  NOR2_X1 U5021 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5701) );
  CLKBUF_X2 U5022 ( .A(n5287), .Z(n4513) );
  BUF_X2 U5023 ( .A(n5287), .Z(n4514) );
  NOR2_X1 U5024 ( .A1(n5833), .A2(n5832), .ZN(n4823) );
  INV_X1 U5025 ( .A(n8358), .ZN(n8120) );
  OAI21_X1 U5026 ( .B1(n7979), .B2(n4880), .A(n4878), .ZN(n6139) );
  AND2_X1 U5027 ( .A1(n5727), .A2(n6514), .ZN(n7729) );
  OR2_X1 U5028 ( .A1(n5883), .A2(n9888), .ZN(n5852) );
  OAI21_X1 U5029 ( .B1(n8728), .B2(n6105), .A(n6106), .ZN(n7977) );
  INV_X1 U5030 ( .A(n8353), .ZN(n8129) );
  NAND2_X1 U5032 ( .A1(n6492), .A2(n6317), .ZN(n9385) );
  INV_X1 U5033 ( .A(n5391), .ZN(n5594) );
  OAI21_X1 U5034 ( .B1(n5609), .B2(n10288), .A(n5248), .ZN(n5250) );
  NAND2_X2 U5035 ( .A1(n8144), .A2(n9007), .ZN(n5898) );
  NOR2_X1 U5036 ( .A1(n9935), .A2(n9936), .ZN(n9934) );
  INV_X1 U5037 ( .A(n8326), .ZN(n8336) );
  BUF_X1 U5038 ( .A(n5869), .Z(n6229) );
  AOI21_X1 U5039 ( .B1(n4812), .B2(n4818), .A(n8160), .ZN(n4810) );
  NAND2_X1 U5040 ( .A1(n4824), .A2(n4825), .ZN(n7821) );
  INV_X2 U5041 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9002) );
  INV_X2 U5042 ( .A(n5171), .ZN(n5382) );
  AND2_X1 U5043 ( .A1(n5170), .A2(n5166), .ZN(n5327) );
  NAND2_X2 U5044 ( .A1(n7973), .A2(n9684), .ZN(n6709) );
  INV_X1 U5045 ( .A(n7253), .ZN(n9809) );
  NAND4_X2 U5046 ( .A1(n5877), .A2(n5876), .A3(n5875), .A4(n5874), .ZN(n8207)
         );
  INV_X1 U5047 ( .A(n6020), .ZN(n8148) );
  NAND2_X1 U5048 ( .A1(n6243), .A2(n8272), .ZN(n8750) );
  NAND2_X1 U5049 ( .A1(n5484), .A2(n5483), .ZN(n8011) );
  XNOR2_X1 U5050 ( .A(n5008), .B(n6344), .ZN(n9001) );
  NAND2_X1 U5051 ( .A1(n5388), .A2(n5387), .ZN(n5390) );
  OAI21_X1 U5052 ( .B1(n5297), .B2(n5296), .A(n4991), .ZN(n5313) );
  NAND2_X1 U5053 ( .A1(n6272), .A2(n6271), .ZN(n9017) );
  AOI21_X1 U5054 ( .B1(n9001), .B2(n6347), .A(n6346), .ZN(n9579) );
  XNOR2_X1 U5055 ( .A(n5334), .B(n5333), .ZN(n6753) );
  NAND2_X2 U5056 ( .A1(n7631), .A2(n7630), .ZN(n7629) );
  CLKBUF_X2 U5057 ( .A(n8825), .Z(n4507) );
  NAND4_X1 U5058 ( .A1(n5887), .A2(n5886), .A3(n5885), .A4(n5884), .ZN(n8825)
         );
  AND2_X2 U5059 ( .A1(n4815), .A2(n4813), .ZN(n4812) );
  NAND2_X2 U5060 ( .A1(n5114), .A2(n5112), .ZN(n7996) );
  OAI222_X1 U5061 ( .A1(n9018), .A2(n7819), .B1(P2_U3151), .B2(n6276), .C1(
        n7808), .C2(n9015), .ZN(P2_U3271) );
  NAND2_X2 U5062 ( .A1(n4736), .A2(n4737), .ZN(n9051) );
  OAI21_X2 U5063 ( .B1(n5590), .B2(n5589), .A(n5247), .ZN(n5609) );
  OAI21_X2 U5064 ( .B1(n5572), .B2(n5241), .A(n5243), .ZN(n5590) );
  OAI21_X2 U5065 ( .B1(n7821), .B2(n8173), .A(n8250), .ZN(n7838) );
  OAI21_X2 U5066 ( .B1(n7386), .B2(n5720), .A(n4930), .ZN(n4929) );
  OR3_X4 U5067 ( .A1(n9139), .A2(n9143), .A3(n9035), .ZN(n9104) );
  AOI21_X2 U5068 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n7547), .A(n7546), .ZN(
        n7550) );
  OAI21_X2 U5069 ( .B1(n9409), .B2(n6461), .A(n6458), .ZN(n9396) );
  NAND2_X2 U5070 ( .A1(n9427), .A2(n6455), .ZN(n9409) );
  XNOR2_X2 U5071 ( .A(n5592), .B(P1_IR_REG_19__SCAN_IN), .ZN(n6542) );
  NAND2_X1 U5072 ( .A1(n8144), .A2(n5850), .ZN(n5909) );
  XNOR2_X2 U5073 ( .A(n5846), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5850) );
  AOI21_X2 U5074 ( .B1(n5095), .B2(n4555), .A(n5091), .ZN(n8373) );
  XNOR2_X1 U5075 ( .A(n5858), .B(n5840), .ZN(n4508) );
  INV_X8 U5076 ( .A(n8346), .ZN(n9876) );
  AOI21_X2 U5077 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n7867), .A(n7866), .ZN(
        n7868) );
  OAI222_X1 U5078 ( .A1(P1_U3086), .A2(n6756), .B1(n9687), .B2(n5295), .C1(
        n6688), .C2(n9689), .ZN(P1_U3354) );
  OR2_X1 U5079 ( .A1(n6488), .A2(n5711), .ZN(n4600) );
  INV_X1 U5080 ( .A(n8368), .ZN(n4510) );
  NAND2_X1 U5081 ( .A1(n5691), .A2(n5690), .ZN(n8368) );
  OR2_X1 U5082 ( .A1(n6461), .A2(n6464), .ZN(n9413) );
  NAND2_X1 U5083 ( .A1(n5277), .A2(n5276), .ZN(n5688) );
  NAND2_X1 U5084 ( .A1(n5642), .A2(n5641), .ZN(n9608) );
  NAND2_X1 U5085 ( .A1(n5620), .A2(n5619), .ZN(n9478) );
  NAND2_X1 U5086 ( .A1(n5541), .A2(n5540), .ZN(n9548) );
  NAND2_X2 U5087 ( .A1(n6425), .A2(n6510), .ZN(n7618) );
  INV_X1 U5088 ( .A(n7663), .ZN(n10053) );
  OR2_X1 U5089 ( .A1(n5463), .A2(n5462), .ZN(n5039) );
  INV_X4 U5090 ( .A(n6590), .ZN(n7997) );
  NAND2_X1 U5091 ( .A1(n6571), .A2(n6570), .ZN(n6582) );
  INV_X1 U5092 ( .A(n6991), .ZN(n9796) );
  NAND2_X2 U5093 ( .A1(n6237), .A2(n8199), .ZN(n7055) );
  NOR2_X1 U5094 ( .A1(n9218), .A2(n7228), .ZN(n7222) );
  XNOR2_X1 U5095 ( .A(n6859), .B(n9783), .ZN(n5713) );
  NAND4_X1 U5096 ( .A1(n5919), .A2(n5918), .A3(n5917), .A4(n5916), .ZN(n8527)
         );
  NAND4_X2 U5097 ( .A1(n5855), .A2(n5854), .A3(n5853), .A4(n5852), .ZN(n6572)
         );
  INV_X2 U5098 ( .A(n5898), .ZN(n5952) );
  BUF_X4 U5099 ( .A(n5988), .Z(n4509) );
  XNOR2_X1 U5100 ( .A(n5858), .B(n5840), .ZN(n6227) );
  NAND3_X1 U5101 ( .A1(n4660), .A2(n4823), .A3(n5890), .ZN(n4661) );
  NAND2_X1 U5102 ( .A1(n5879), .A2(n4968), .ZN(n6966) );
  AND2_X1 U5103 ( .A1(n5129), .A2(n4547), .ZN(n5127) );
  NOR2_X2 U5104 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5315) );
  INV_X1 U5105 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5776) );
  NAND2_X1 U5106 ( .A1(n4806), .A2(n4804), .ZN(n8611) );
  OR2_X1 U5107 ( .A1(n9364), .A2(n9365), .ZN(n5808) );
  AND2_X1 U5108 ( .A1(n4804), .A2(n10101), .ZN(n4803) );
  OAI21_X1 U5109 ( .B1(n6489), .B2(n9344), .A(n6883), .ZN(n4599) );
  OR2_X1 U5110 ( .A1(n6484), .A2(n4719), .ZN(n4718) );
  NOR2_X1 U5111 ( .A1(n8330), .A2(n4765), .ZN(n8337) );
  NOR2_X1 U5112 ( .A1(n4895), .A2(n6474), .ZN(n4894) );
  NOR2_X1 U5113 ( .A1(n4654), .A2(n4653), .ZN(n8333) );
  OR2_X1 U5114 ( .A1(n6549), .A2(n6485), .ZN(n4724) );
  AOI21_X1 U5115 ( .B1(n4902), .B2(n4908), .A(n4901), .ZN(n4900) );
  AND2_X1 U5116 ( .A1(n6348), .A2(n6481), .ZN(n6549) );
  INV_X1 U5117 ( .A(n9357), .ZN(n9649) );
  NAND2_X1 U5118 ( .A1(n8060), .A2(n8059), .ZN(n9156) );
  NAND2_X1 U5119 ( .A1(n5676), .A2(n5675), .ZN(n9401) );
  OAI21_X1 U5120 ( .B1(n6342), .B2(n6341), .A(n6340), .ZN(n5008) );
  XNOR2_X1 U5121 ( .A(n6342), .B(n6341), .ZN(n8146) );
  OR2_X1 U5122 ( .A1(n10019), .A2(n8538), .ZN(n4700) );
  OAI21_X1 U5123 ( .B1(n5733), .B2(n4941), .A(n4939), .ZN(n5735) );
  AND2_X1 U5124 ( .A1(n6252), .A2(n8315), .ZN(n4807) );
  NAND2_X1 U5125 ( .A1(n9021), .A2(n5066), .ZN(n5065) );
  NAND2_X1 U5126 ( .A1(n6189), .A2(n6188), .ZN(n8919) );
  NAND2_X1 U5127 ( .A1(n5289), .A2(n5288), .ZN(n9390) );
  OAI21_X1 U5128 ( .B1(n9454), .B2(n5637), .A(n5638), .ZN(n9441) );
  XNOR2_X1 U5129 ( .A(n6326), .B(n6324), .ZN(n6323) );
  AOI21_X1 U5130 ( .B1(n8587), .B2(n8586), .A(n8585), .ZN(n8593) );
  INV_X1 U5131 ( .A(n4940), .ZN(n4939) );
  XNOR2_X1 U5132 ( .A(n5688), .B(n5687), .ZN(n7991) );
  OAI21_X1 U5133 ( .B1(n5588), .B2(n4650), .A(n4648), .ZN(n9470) );
  AND2_X1 U5134 ( .A1(n5141), .A2(n6149), .ZN(n4884) );
  NAND2_X1 U5135 ( .A1(n6170), .A2(n6169), .ZN(n8931) );
  OR2_X1 U5136 ( .A1(n9984), .A2(n9983), .ZN(n4973) );
  NAND2_X1 U5137 ( .A1(n5655), .A2(n5654), .ZN(n9601) );
  OAI21_X1 U5138 ( .B1(n8750), .B2(n8752), .A(n8273), .ZN(n8740) );
  NAND2_X1 U5139 ( .A1(n6130), .A2(n6129), .ZN(n8953) );
  OAI21_X1 U5140 ( .B1(n5618), .B2(n5253), .A(n5252), .ZN(n5627) );
  NAND2_X1 U5141 ( .A1(n5611), .A2(n5610), .ZN(n9623) );
  NAND2_X1 U5142 ( .A1(n9961), .A2(n8553), .ZN(n9978) );
  OR2_X1 U5143 ( .A1(n7957), .A2(n7918), .ZN(n4701) );
  AND2_X1 U5144 ( .A1(n6520), .A2(n6417), .ZN(n9562) );
  NAND2_X1 U5145 ( .A1(n6591), .A2(n7453), .ZN(n7457) );
  XNOR2_X1 U5146 ( .A(n5537), .B(n5536), .ZN(n7075) );
  NAND2_X1 U5147 ( .A1(n5015), .A2(n5012), .ZN(n5537) );
  OR2_X1 U5148 ( .A1(n6741), .A2(n5341), .ZN(n5484) );
  NAND2_X1 U5149 ( .A1(n4865), .A2(n5950), .ZN(n7640) );
  NAND2_X1 U5150 ( .A1(n5494), .A2(n5493), .ZN(n9137) );
  OR2_X1 U5151 ( .A1(n9732), .A2(n7789), .ZN(n7617) );
  AOI21_X1 U5152 ( .B1(n8236), .B2(n4835), .A(n4834), .ZN(n4833) );
  NAND2_X1 U5153 ( .A1(n5455), .A2(n5454), .ZN(n9704) );
  OAI21_X1 U5154 ( .B1(n5506), .B2(SI_14_), .A(n5504), .ZN(n5231) );
  NAND2_X1 U5155 ( .A1(n5984), .A2(n5983), .ZN(n10071) );
  OR2_X1 U5156 ( .A1(n7751), .A2(n7752), .ZN(n4688) );
  NAND2_X1 U5157 ( .A1(n5467), .A2(n5466), .ZN(n9732) );
  AND2_X1 U5158 ( .A1(n8237), .A2(n8233), .ZN(n4835) );
  NAND2_X1 U5159 ( .A1(n7423), .A2(n5925), .ZN(n5927) );
  OR2_X1 U5160 ( .A1(n10065), .A2(n7676), .ZN(n8240) );
  NAND2_X1 U5161 ( .A1(n4986), .A2(n4985), .ZN(n4984) );
  NAND2_X1 U5162 ( .A1(n5973), .A2(n5972), .ZN(n10065) );
  OAI211_X1 U5163 ( .C1(n6229), .C2(n7475), .A(n5949), .B(n5948), .ZN(n7663)
         );
  OAI21_X1 U5164 ( .B1(n5402), .B2(n5401), .A(n5403), .ZN(n6699) );
  INV_X2 U5165 ( .A(n6582), .ZN(n6590) );
  NOR2_X1 U5166 ( .A1(P2_U3150), .A2(n6958), .ZN(n10007) );
  NOR2_X1 U5167 ( .A1(n7179), .A2(n7178), .ZN(n7474) );
  AND2_X1 U5168 ( .A1(n8223), .A2(n8216), .ZN(n8165) );
  BUF_X2 U5169 ( .A(n6981), .Z(n8358) );
  AOI21_X1 U5170 ( .B1(n6792), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6791), .ZN(
        n6817) );
  NOR2_X1 U5171 ( .A1(n9934), .A2(n4605), .ZN(n7031) );
  BUF_X4 U5172 ( .A(n6915), .Z(n8130) );
  NAND2_X1 U5173 ( .A1(n6843), .A2(n6842), .ZN(n6846) );
  AND4_X1 U5174 ( .A1(n5351), .A2(n5350), .A3(n5349), .A4(n5348), .ZN(n7263)
         );
  AND4_X1 U5175 ( .A1(n5386), .A2(n5385), .A3(n5384), .A4(n5383), .ZN(n7345)
         );
  AND4_X1 U5176 ( .A1(n5369), .A2(n5368), .A3(n5367), .A4(n5366), .ZN(n7260)
         );
  OAI211_X1 U5177 ( .C1(n6966), .C2(n6229), .A(n4889), .B(n4886), .ZN(n6578)
         );
  NAND2_X2 U5178 ( .A1(n6841), .A2(n6875), .ZN(n8356) );
  INV_X1 U5179 ( .A(n6572), .ZN(n5863) );
  NAND4_X1 U5180 ( .A1(n5307), .A2(n5306), .A3(n5305), .A4(n5304), .ZN(n9218)
         );
  INV_X1 U5181 ( .A(n5035), .ZN(n5034) );
  AOI21_X1 U5182 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n9266), .A(n6747), .ZN(
        n6750) );
  AOI21_X1 U5183 ( .B1(n5035), .B2(n5037), .A(n5490), .ZN(n5033) );
  NAND2_X1 U5184 ( .A1(n5780), .A2(n5043), .ZN(n6875) );
  INV_X1 U5185 ( .A(n7096), .ZN(n6231) );
  INV_X2 U5186 ( .A(n6542), .ZN(n5711) );
  NAND2_X1 U5187 ( .A1(n6266), .A2(n6265), .ZN(n6276) );
  AND3_X2 U5188 ( .A1(n5302), .A2(n5301), .A3(n5300), .ZN(n9783) );
  INV_X2 U5189 ( .A(n5341), .ZN(n6347) );
  XNOR2_X1 U5190 ( .A(n5777), .B(n5776), .ZN(n6842) );
  AND2_X1 U5191 ( .A1(n5170), .A2(n9682), .ZN(n5320) );
  OR2_X1 U5192 ( .A1(n6264), .A2(n6263), .ZN(n6265) );
  BUF_X2 U5193 ( .A(n5327), .Z(n4596) );
  AND2_X1 U5194 ( .A1(n5211), .A2(n5210), .ZN(n5401) );
  NAND2_X1 U5195 ( .A1(n5869), .A2(n4513), .ZN(n6020) );
  NAND2_X4 U5196 ( .A1(n6709), .A2(n4513), .ZN(n5391) );
  XNOR2_X1 U5197 ( .A(n5705), .B(n5704), .ZN(n6840) );
  AND2_X1 U5198 ( .A1(n5165), .A2(n9677), .ZN(n5166) );
  XNOR2_X1 U5199 ( .A(n6108), .B(n5835), .ZN(n8596) );
  INV_X1 U5200 ( .A(n6227), .ZN(n8346) );
  XNOR2_X1 U5201 ( .A(n5708), .B(n5707), .ZN(n7557) );
  OR2_X1 U5202 ( .A1(n5180), .A2(SI_1_), .ZN(n5181) );
  MUX2_X1 U5203 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5163), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5165) );
  XNOR2_X1 U5204 ( .A(n6224), .B(n5837), .ZN(n8343) );
  OR2_X1 U5205 ( .A1(n6270), .A2(n9002), .ZN(n5858) );
  NAND2_X1 U5206 ( .A1(n9003), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5846) );
  NAND2_X1 U5207 ( .A1(n4658), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5284) );
  INV_X2 U5208 ( .A(n9005), .ZN(n9015) );
  NOR2_X1 U5209 ( .A1(n4661), .A2(n4659), .ZN(n6270) );
  OR2_X1 U5210 ( .A1(n5072), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n4521) );
  AND2_X1 U5211 ( .A1(n4616), .A2(n4615), .ZN(n4617) );
  AND4_X1 U5212 ( .A1(n5149), .A2(n5148), .A3(n5147), .A4(n10494), .ZN(n5150)
         );
  AND2_X1 U5213 ( .A1(n5834), .A2(n5130), .ZN(n5129) );
  NOR2_X1 U5214 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5829) );
  NOR2_X1 U5215 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5828) );
  NOR2_X1 U5216 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5827) );
  INV_X4 U5217 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X4 U5218 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5219 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5921) );
  INV_X1 U5220 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4615) );
  INV_X1 U5221 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4616) );
  INV_X1 U5222 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6003) );
  INV_X1 U5223 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6007) );
  INV_X1 U5224 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n10235) );
  NOR2_X1 U5225 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n5159) );
  INV_X1 U5226 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5158) );
  INV_X1 U5227 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5704) );
  INV_X1 U5228 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5707) );
  INV_X1 U5229 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n10519) );
  INV_X1 U5231 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n10494) );
  NOR3_X1 U5232 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .A3(
        P2_IR_REG_24__SCAN_IN), .ZN(n5839) );
  INV_X1 U5233 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5130) );
  INV_X1 U5234 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5834) );
  NOR2_X1 U5235 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5148) );
  AOI21_X2 U5236 ( .B1(n8780), .B2(n8267), .A(n8269), .ZN(n8763) );
  AND2_X4 U5237 ( .A1(n5878), .A2(n5826), .ZN(n5890) );
  NAND2_X2 U5238 ( .A1(n5863), .A2(n5870), .ZN(n6237) );
  OAI22_X2 U5239 ( .A1(n8633), .A2(n8634), .B1(n8622), .B2(n8919), .ZN(n8618)
         );
  OAI21_X2 U5240 ( .B1(n6219), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6291) );
  OAI21_X2 U5241 ( .B1(n7270), .B2(n5896), .A(n5895), .ZN(n7281) );
  OAI21_X2 U5242 ( .B1(n7640), .B2(n8524), .A(n5966), .ZN(n7810) );
  BUF_X8 U5243 ( .A(n5859), .Z(n4511) );
  INV_X2 U5244 ( .A(n5287), .ZN(n5859) );
  AND2_X1 U5245 ( .A1(n5170), .A2(n9682), .ZN(n4512) );
  XNOR2_X2 U5246 ( .A(n5161), .B(n5160), .ZN(n8140) );
  AOI21_X2 U5247 ( .B1(n6273), .B2(n7881), .A(n9017), .ZN(n6275) );
  XNOR2_X2 U5248 ( .A(n5299), .B(n5298), .ZN(n6756) );
  NAND2_X1 U5249 ( .A1(n5178), .A2(n5179), .ZN(n5287) );
  AND2_X2 U5250 ( .A1(n5861), .A2(n4971), .ZN(n5878) );
  NOR2_X4 U5251 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5861) );
  NAND2_X1 U5252 ( .A1(n5848), .A2(n5850), .ZN(n5988) );
  NOR2_X2 U5253 ( .A1(n8470), .A2(n8402), .ZN(n5095) );
  NOR2_X2 U5254 ( .A1(n7928), .A2(n7929), .ZN(n8470) );
  NAND2_X1 U5255 ( .A1(n4630), .A2(n4629), .ZN(n8292) );
  NAND2_X1 U5256 ( .A1(n8288), .A2(n8326), .ZN(n4629) );
  OAI21_X1 U5257 ( .B1(n4632), .B2(n4627), .A(n4625), .ZN(n4630) );
  OR2_X1 U5258 ( .A1(n8324), .A2(n8623), .ZN(n8328) );
  OR2_X1 U5259 ( .A1(n5811), .A2(n7077), .ZN(n6476) );
  AOI21_X1 U5260 ( .B1(n5028), .B2(n5027), .A(n5026), .ZN(n5025) );
  NAND2_X1 U5261 ( .A1(n8285), .A2(n8274), .ZN(n4779) );
  AOI21_X1 U5262 ( .B1(n4781), .B2(n8273), .A(n8741), .ZN(n4780) );
  OR2_X1 U5263 ( .A1(n8295), .A2(n8326), .ZN(n4777) );
  NOR2_X1 U5264 ( .A1(n8322), .A2(n8323), .ZN(n4653) );
  AOI21_X1 U5265 ( .B1(n8317), .B2(n4656), .A(n4655), .ZN(n4654) );
  NAND2_X1 U5266 ( .A1(n5001), .A2(n5000), .ZN(n6326) );
  AOI21_X1 U5267 ( .B1(n5003), .B2(n5005), .A(n4588), .ZN(n5000) );
  NAND2_X1 U5268 ( .A1(n5688), .A2(n5003), .ZN(n5001) );
  NAND2_X1 U5269 ( .A1(n7515), .A2(n7514), .ZN(n4986) );
  NAND2_X1 U5270 ( .A1(n4701), .A2(n7919), .ZN(n4965) );
  INV_X1 U5271 ( .A(n7072), .ZN(n5870) );
  OR2_X1 U5272 ( .A1(n8953), .A2(n8691), .ZN(n8193) );
  OR2_X1 U5273 ( .A1(n4723), .A2(n6842), .ZN(n4719) );
  NAND2_X1 U5274 ( .A1(n5290), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5291) );
  OR2_X1 U5275 ( .A1(n9628), .A2(n5731), .ZN(n6433) );
  AND2_X1 U5276 ( .A1(n5276), .A2(n5275), .ZN(n5677) );
  AOI21_X1 U5277 ( .B1(n5663), .B2(n4998), .A(n4997), .ZN(n4996) );
  INV_X1 U5278 ( .A(n5267), .ZN(n4998) );
  INV_X1 U5279 ( .A(n5272), .ZN(n4997) );
  INV_X1 U5280 ( .A(n5663), .ZN(n4999) );
  INV_X1 U5281 ( .A(n8469), .ZN(n5088) );
  NOR2_X1 U5282 ( .A1(n8342), .A2(n4677), .ZN(n4676) );
  NAND2_X1 U5284 ( .A1(n7190), .A2(n7191), .ZN(n7466) );
  NAND2_X1 U5285 ( .A1(n7194), .A2(n7192), .ZN(n7190) );
  XNOR2_X1 U5286 ( .A(n4984), .B(n4983), .ZN(n7751) );
  XNOR2_X1 U5287 ( .A(n4966), .B(n7917), .ZN(n7958) );
  OR2_X1 U5288 ( .A1(n6160), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6171) );
  INV_X1 U5289 ( .A(n4879), .ZN(n4878) );
  INV_X1 U5290 ( .A(n7979), .ZN(n4882) );
  NAND2_X1 U5291 ( .A1(n6093), .A2(n6092), .ZN(n8728) );
  AOI21_X1 U5292 ( .B1(n4828), .B2(n4827), .A(n4826), .ZN(n4825) );
  INV_X1 U5293 ( .A(n8240), .ZN(n4826) );
  XNOR2_X1 U5294 ( .A(n8913), .B(n8636), .ZN(n8620) );
  OR2_X1 U5295 ( .A1(n8937), .A2(n8682), .ZN(n6167) );
  OR2_X1 U5296 ( .A1(n8943), .A2(n8692), .ZN(n8665) );
  NAND2_X1 U5297 ( .A1(n7979), .A2(n4883), .ZN(n8715) );
  OR2_X1 U5298 ( .A1(n8391), .A2(n8729), .ZN(n8711) );
  INV_X1 U5299 ( .A(n8261), .ZN(n4816) );
  NAND2_X1 U5300 ( .A1(n6709), .A2(n4633), .ZN(n4635) );
  AND2_X1 U5301 ( .A1(n4514), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4633) );
  NAND2_X1 U5302 ( .A1(n5065), .A2(n4517), .ZN(n4756) );
  NOR2_X1 U5303 ( .A1(n4724), .A2(n4535), .ZN(n4723) );
  AND2_X1 U5304 ( .A1(n4715), .A2(n4714), .ZN(n4722) );
  NAND2_X1 U5305 ( .A1(n4535), .A2(n9357), .ZN(n4714) );
  NAND2_X1 U5306 ( .A1(n4724), .A2(n4559), .ZN(n4715) );
  OAI211_X1 U5307 ( .C1(n6472), .C2(n6471), .A(n4566), .B(n4725), .ZN(n6475)
         );
  INV_X1 U5308 ( .A(n6483), .ZN(n6554) );
  OR2_X1 U5309 ( .A1(n5811), .A2(n5806), .ZN(n9356) );
  NOR2_X1 U5310 ( .A1(n5605), .A2(n4652), .ZN(n4651) );
  INV_X1 U5311 ( .A(n5587), .ZN(n4652) );
  NAND2_X1 U5312 ( .A1(n4957), .A2(n4956), .ZN(n5588) );
  AND2_X1 U5313 ( .A1(n5144), .A2(n5570), .ZN(n4956) );
  INV_X1 U5314 ( .A(n6416), .ZN(n4915) );
  INV_X1 U5315 ( .A(n9504), .ZN(n9756) );
  AND2_X1 U5316 ( .A1(n6875), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5781) );
  AND2_X1 U5317 ( .A1(n5392), .A2(n5156), .ZN(n4657) );
  NOR2_X1 U5318 ( .A1(n5626), .A2(n5031), .ZN(n5030) );
  INV_X1 U5319 ( .A(n5252), .ZN(n5031) );
  AND2_X1 U5320 ( .A1(n5262), .A2(n5261), .ZN(n5639) );
  INV_X1 U5321 ( .A(n6229), .ZN(n6682) );
  OR2_X1 U5322 ( .A1(n6613), .A2(n8754), .ZN(n6614) );
  NAND2_X1 U5323 ( .A1(n6623), .A2(n6622), .ZN(n8443) );
  INV_X1 U5324 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5856) );
  AND2_X1 U5325 ( .A1(n4938), .A2(n4516), .ZN(n5787) );
  NOR2_X1 U5326 ( .A1(n4667), .A2(n8246), .ZN(n4666) );
  NAND2_X1 U5327 ( .A1(n4665), .A2(n4668), .ZN(n4669) );
  NOR2_X1 U5328 ( .A1(n8246), .A2(n8326), .ZN(n4668) );
  NAND2_X1 U5329 ( .A1(n8252), .A2(n8254), .ZN(n4785) );
  NAND2_X1 U5330 ( .A1(n4618), .A2(n8764), .ZN(n8276) );
  INV_X1 U5331 ( .A(n8271), .ZN(n4619) );
  NAND2_X1 U5332 ( .A1(n4702), .A2(n6408), .ZN(n6422) );
  OAI21_X1 U5333 ( .B1(n6400), .B2(n6550), .A(n4703), .ZN(n4702) );
  OAI21_X1 U5334 ( .B1(n6418), .B2(n6493), .A(n6520), .ZN(n4713) );
  NOR2_X1 U5335 ( .A1(n6420), .A2(n6550), .ZN(n4711) );
  AOI21_X1 U5336 ( .B1(n4662), .B2(n4775), .A(n8304), .ZN(n8312) );
  INV_X1 U5337 ( .A(n6449), .ZN(n4709) );
  AND2_X1 U5338 ( .A1(n4537), .A2(n6627), .ZN(n5110) );
  NOR2_X1 U5339 ( .A1(n4873), .A2(n4871), .ZN(n4870) );
  INV_X1 U5340 ( .A(n6187), .ZN(n4871) );
  NAND2_X1 U5341 ( .A1(n6211), .A2(n6255), .ZN(n4873) );
  NAND2_X1 U5342 ( .A1(n6409), .A2(n7404), .ZN(n6405) );
  NOR2_X1 U5343 ( .A1(n9548), .A2(n9573), .ZN(n4856) );
  AND2_X1 U5344 ( .A1(n5110), .A2(n4545), .ZN(n5104) );
  INV_X1 U5345 ( .A(n8444), .ZN(n5102) );
  AOI22_X1 U5346 ( .A1(n5109), .A2(n4537), .B1(n5110), .B2(n8394), .ZN(n5108)
         );
  INV_X1 U5347 ( .A(n8461), .ZN(n5109) );
  OAI22_X1 U5348 ( .A1(n9892), .A2(n6946), .B1(n4972), .B2(n9878), .ZN(n9889)
         );
  NAND2_X1 U5349 ( .A1(n4792), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9891) );
  INV_X1 U5350 ( .A(n9889), .ZN(n4792) );
  OR2_X1 U5351 ( .A1(n9892), .A2(n6964), .ZN(n4692) );
  NOR2_X1 U5352 ( .A1(n7215), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6964) );
  NAND2_X1 U5353 ( .A1(n9904), .A2(n6967), .ZN(n6969) );
  NAND2_X1 U5354 ( .A1(n7037), .A2(n7036), .ZN(n7038) );
  NAND2_X1 U5355 ( .A1(n4961), .A2(n4960), .ZN(n4689) );
  INV_X1 U5356 ( .A(n7038), .ZN(n4961) );
  NAND2_X1 U5357 ( .A1(n8569), .A2(n4791), .ZN(n8572) );
  OR2_X1 U5358 ( .A1(n8570), .A2(n8899), .ZN(n4791) );
  NOR2_X1 U5359 ( .A1(n9966), .A2(n4974), .ZN(n8535) );
  NOR2_X1 U5360 ( .A1(n9957), .A2(n8784), .ZN(n4974) );
  OR2_X1 U5361 ( .A1(n8318), .A2(n8158), .ZN(n8313) );
  OR2_X1 U5362 ( .A1(n8937), .A2(n8414), .ZN(n8305) );
  AND2_X1 U5363 ( .A1(n8716), .A2(n6119), .ZN(n4883) );
  OR2_X1 U5364 ( .A1(n8968), .A2(n8756), .ZN(n8281) );
  OR2_X1 U5365 ( .A1(n8978), .A2(n8754), .ZN(n8272) );
  AND2_X1 U5366 ( .A1(n7204), .A2(n7068), .ZN(n6658) );
  NOR2_X1 U5367 ( .A1(n5132), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n4891) );
  NOR2_X1 U5368 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n5133) );
  NAND2_X1 U5369 ( .A1(n5127), .A2(n5837), .ZN(n5126) );
  INV_X1 U5370 ( .A(n9103), .ZN(n5085) );
  NOR2_X1 U5371 ( .A1(n9080), .A2(n5069), .ZN(n5066) );
  NAND2_X1 U5372 ( .A1(n4904), .A2(n4520), .ZN(n4726) );
  INV_X1 U5373 ( .A(n4719), .ZN(n4721) );
  INV_X1 U5374 ( .A(n4722), .ZN(n4717) );
  NOR2_X1 U5375 ( .A1(n9418), .A2(n9402), .ZN(n4845) );
  INV_X1 U5376 ( .A(n6443), .ZN(n4941) );
  NOR2_X1 U5377 ( .A1(n4548), .A2(n4944), .ZN(n4943) );
  INV_X1 U5378 ( .A(n5606), .ZN(n4944) );
  INV_X1 U5379 ( .A(n4651), .ZN(n4649) );
  INV_X1 U5380 ( .A(n6386), .ZN(n4942) );
  AND2_X1 U5381 ( .A1(n4856), .A2(n4855), .ZN(n4854) );
  AOI21_X1 U5382 ( .B1(n4927), .B2(n4923), .A(n4922), .ZN(n4921) );
  NAND2_X1 U5383 ( .A1(n4920), .A2(n4925), .ZN(n4919) );
  INV_X1 U5384 ( .A(n4921), .ZN(n4920) );
  OR2_X1 U5385 ( .A1(n9137), .A2(n8018), .ZN(n6514) );
  NOR2_X1 U5386 ( .A1(n6360), .A2(n4638), .ZN(n4637) );
  INV_X1 U5387 ( .A(n4641), .ZN(n4638) );
  NAND2_X1 U5388 ( .A1(n7238), .A2(n6396), .ZN(n7386) );
  NAND2_X1 U5389 ( .A1(n9215), .A2(n9789), .ZN(n6497) );
  NAND2_X1 U5390 ( .A1(n6328), .A2(n6327), .ZN(n6342) );
  OR2_X1 U5391 ( .A1(n6326), .A2(n6325), .ZN(n6327) );
  NAND2_X1 U5392 ( .A1(n5573), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5577) );
  AOI21_X1 U5393 ( .B1(n5013), .B2(n5011), .A(n4584), .ZN(n5010) );
  AOI21_X1 U5394 ( .B1(n4567), .B2(n4771), .A(n4528), .ZN(n4768) );
  INV_X1 U5395 ( .A(SI_9_), .ZN(n5215) );
  NOR2_X1 U5396 ( .A1(n8468), .A2(n4587), .ZN(n5087) );
  NAND2_X1 U5397 ( .A1(n7848), .A2(n6605), .ZN(n6606) );
  OR2_X1 U5398 ( .A1(n6615), .A2(n8509), .ZN(n6616) );
  INV_X1 U5399 ( .A(n5094), .ZN(n5093) );
  OAI21_X1 U5400 ( .B1(n8402), .B2(n5097), .A(n5099), .ZN(n5094) );
  OR2_X1 U5401 ( .A1(n6608), .A2(n8453), .ZN(n5099) );
  INV_X1 U5402 ( .A(n6607), .ZN(n5097) );
  XNOR2_X1 U5403 ( .A(n6578), .B(n6590), .ZN(n6580) );
  INV_X1 U5404 ( .A(n5121), .ZN(n5120) );
  OAI21_X1 U5405 ( .B1(n4533), .B2(n8486), .A(n8485), .ZN(n5121) );
  AND4_X1 U5406 ( .A1(n7101), .A2(n6217), .A3(n6216), .A4(n6215), .ZN(n8623)
         );
  AND3_X1 U5407 ( .A1(n6147), .A2(n6146), .A3(n6145), .ZN(n6148) );
  OAI22_X1 U5408 ( .A1(n7215), .A2(n5909), .B1(n5883), .B2(n9878), .ZN(n5865)
         );
  NAND2_X1 U5409 ( .A1(n4607), .A2(n4606), .ZN(n4605) );
  INV_X1 U5410 ( .A(n6941), .ZN(n4606) );
  INV_X1 U5411 ( .A(n6940), .ZN(n4607) );
  NAND2_X1 U5412 ( .A1(n7466), .A2(n4696), .ZN(n4698) );
  NOR2_X1 U5413 ( .A1(n7475), .A2(n4697), .ZN(n4696) );
  NAND2_X1 U5414 ( .A1(n7466), .A2(n7465), .ZN(n4694) );
  NOR2_X1 U5415 ( .A1(n7474), .A2(n7473), .ZN(n7477) );
  NOR2_X1 U5416 ( .A1(n7477), .A2(n7476), .ZN(n7497) );
  NAND2_X1 U5417 ( .A1(n7750), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4985) );
  NOR2_X1 U5418 ( .A1(n7959), .A2(n7960), .ZN(n7961) );
  INV_X1 U5419 ( .A(n4966), .ZN(n7916) );
  INV_X1 U5420 ( .A(n4965), .ZN(n8530) );
  NAND2_X1 U5421 ( .A1(n7955), .A2(n7907), .ZN(n7908) );
  NAND2_X1 U5422 ( .A1(n7908), .A2(n7909), .ZN(n8569) );
  XNOR2_X1 U5423 ( .A(n8572), .B(n9942), .ZN(n9947) );
  NOR2_X1 U5424 ( .A1(n9968), .A2(n9967), .ZN(n9966) );
  NAND2_X1 U5425 ( .A1(n5890), .A2(n4823), .ZN(n6069) );
  NAND2_X1 U5426 ( .A1(n8599), .A2(n8598), .ZN(n4799) );
  NAND2_X1 U5427 ( .A1(n8602), .A2(n10016), .ZN(n4795) );
  INV_X1 U5428 ( .A(n8601), .ZN(n4794) );
  AND2_X1 U5429 ( .A1(n6182), .A2(n10488), .ZN(n6190) );
  AND3_X1 U5430 ( .A1(n6137), .A2(n6136), .A3(n6135), .ZN(n8691) );
  INV_X1 U5431 ( .A(n6119), .ZN(n4881) );
  INV_X1 U5432 ( .A(n8243), .ZN(n4834) );
  NAND2_X1 U5433 ( .A1(n4861), .A2(n4860), .ZN(n4863) );
  AND2_X1 U5434 ( .A1(n8233), .A2(n8243), .ZN(n8170) );
  NAND2_X1 U5435 ( .A1(n5881), .A2(n5880), .ZN(n7270) );
  OAI21_X1 U5436 ( .B1(n7055), .B2(n7048), .A(n6237), .ZN(n4809) );
  INV_X1 U5437 ( .A(n8204), .ZN(n8822) );
  NAND2_X1 U5438 ( .A1(n7052), .A2(n8196), .ZN(n7053) );
  INV_X1 U5439 ( .A(n4805), .ZN(n4804) );
  NAND2_X1 U5440 ( .A1(n6213), .A2(n6212), .ZN(n8324) );
  NAND2_X1 U5441 ( .A1(n8925), .A2(n8658), .ZN(n4876) );
  AND2_X1 U5442 ( .A1(n6255), .A2(n6254), .ZN(n8634) );
  AND2_X1 U5443 ( .A1(n6178), .A2(n6177), .ZN(n8647) );
  OR2_X1 U5444 ( .A1(n8931), .A2(n8647), .ZN(n8315) );
  INV_X1 U5445 ( .A(n8313), .ZN(n8643) );
  NAND2_X1 U5446 ( .A1(n8688), .A2(n8693), .ZN(n4885) );
  INV_X1 U5447 ( .A(n8180), .ZN(n6117) );
  NAND2_X1 U5448 ( .A1(n6098), .A2(n6097), .ZN(n8483) );
  INV_X1 U5449 ( .A(n8757), .ZN(n8824) );
  NOR2_X1 U5450 ( .A1(n7070), .A2(n6297), .ZN(n6648) );
  INV_X1 U5451 ( .A(n8831), .ZN(n8808) );
  INV_X1 U5452 ( .A(n7881), .ZN(n6290) );
  INV_X1 U5453 ( .A(n6275), .ZN(n6731) );
  NAND2_X1 U5454 ( .A1(n6262), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6264) );
  INV_X1 U5455 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6263) );
  NAND2_X1 U5456 ( .A1(n6264), .A2(n6263), .ZN(n6266) );
  AND2_X1 U5457 ( .A1(n9002), .A2(n4971), .ZN(n4969) );
  OAI211_X1 U5458 ( .C1(n7164), .C2(n4732), .A(n7339), .B(n4730), .ZN(n7342)
         );
  NAND2_X1 U5459 ( .A1(n4731), .A2(n4538), .ZN(n4730) );
  NOR2_X1 U5460 ( .A1(n5077), .A2(n5084), .ZN(n5076) );
  INV_X1 U5461 ( .A(n5086), .ZN(n5077) );
  INV_X1 U5462 ( .A(n9215), .ZN(n6990) );
  AOI21_X1 U5463 ( .B1(n9218), .B2(n6915), .A(n6850), .ZN(n6855) );
  INV_X1 U5464 ( .A(n8068), .ZN(n4741) );
  INV_X1 U5465 ( .A(n9116), .ZN(n4738) );
  INV_X1 U5466 ( .A(n9042), .ZN(n4739) );
  NAND2_X1 U5467 ( .A1(n5064), .A2(n5067), .ZN(n5063) );
  INV_X1 U5468 ( .A(n9080), .ZN(n5064) );
  INV_X1 U5469 ( .A(n8030), .ZN(n5068) );
  OR2_X1 U5470 ( .A1(n5065), .A2(n5068), .ZN(n4757) );
  XNOR2_X1 U5471 ( .A(n6982), .B(n8354), .ZN(n7160) );
  OAI22_X1 U5472 ( .A1(n8358), .A2(n9796), .B1(n7087), .B2(n8356), .ZN(n6982)
         );
  NOR2_X1 U5473 ( .A1(n5438), .A2(n6799), .ZN(n5456) );
  INV_X1 U5474 ( .A(n9059), .ZN(n5055) );
  NOR2_X1 U5475 ( .A1(n5056), .A2(n5053), .ZN(n5052) );
  INV_X1 U5476 ( .A(n9131), .ZN(n5056) );
  OR2_X1 U5477 ( .A1(n8091), .A2(n8089), .ZN(n8087) );
  NAND2_X1 U5478 ( .A1(n9086), .A2(n4525), .ZN(n9154) );
  INV_X1 U5479 ( .A(n8054), .ZN(n5050) );
  NOR2_X1 U5480 ( .A1(n9356), .A2(n9357), .ZN(n9360) );
  NAND2_X1 U5481 ( .A1(n5795), .A2(n5794), .ZN(n5811) );
  NAND2_X1 U5482 ( .A1(n9385), .A2(n6317), .ZN(n4906) );
  OR2_X1 U5483 ( .A1(n6470), .A2(n4901), .ZN(n6374) );
  NAND2_X1 U5484 ( .A1(n9432), .A2(n4842), .ZN(n5806) );
  AND2_X1 U5485 ( .A1(n4843), .A2(n4510), .ZN(n4842) );
  NAND2_X1 U5486 ( .A1(n9401), .A2(n6371), .ZN(n4681) );
  OAI21_X1 U5487 ( .B1(n9470), .B2(n5625), .A(n4950), .ZN(n9454) );
  OR2_X1 U5488 ( .A1(n9478), .A2(n9198), .ZN(n4950) );
  NAND2_X1 U5489 ( .A1(n5733), .A2(n4534), .ZN(n9471) );
  OR2_X1 U5490 ( .A1(n9623), .A2(n5732), .ZN(n6386) );
  AND2_X1 U5491 ( .A1(n6386), .A2(n6387), .ZN(n9487) );
  NOR2_X1 U5492 ( .A1(n4561), .A2(n4645), .ZN(n4644) );
  INV_X1 U5493 ( .A(n5550), .ZN(n4645) );
  OAI21_X1 U5494 ( .B1(n9563), .B2(n5533), .A(n5532), .ZN(n9542) );
  OR2_X1 U5495 ( .A1(n7728), .A2(n4916), .ZN(n4909) );
  NAND2_X1 U5496 ( .A1(n4912), .A2(n4910), .ZN(n9543) );
  AND2_X1 U5497 ( .A1(n4647), .A2(n4911), .ZN(n4910) );
  NOR2_X1 U5498 ( .A1(n7407), .A2(n4642), .ZN(n4641) );
  INV_X1 U5499 ( .A(n7429), .ZN(n4642) );
  NOR2_X1 U5500 ( .A1(n4949), .A2(n4947), .ZN(n4946) );
  INV_X1 U5501 ( .A(n5416), .ZN(n4947) );
  AND2_X1 U5502 ( .A1(n6409), .A2(n6421), .ZN(n7407) );
  NAND2_X1 U5503 ( .A1(n7384), .A2(n7387), .ZN(n4948) );
  NAND2_X1 U5504 ( .A1(n4589), .A2(n9809), .ZN(n9748) );
  NAND2_X1 U5505 ( .A1(n7223), .A2(n7222), .ZN(n7221) );
  AND2_X1 U5506 ( .A1(n6884), .A2(n7557), .ZN(n9765) );
  NAND2_X1 U5507 ( .A1(n5596), .A2(n5595), .ZN(n9628) );
  INV_X1 U5508 ( .A(n9765), .ZN(n9850) );
  OR2_X1 U5509 ( .A1(n5391), .A2(n5295), .ZN(n5302) );
  AND2_X1 U5510 ( .A1(n5738), .A2(n6552), .ZN(n9504) );
  OR2_X1 U5511 ( .A1(n5752), .A2(n4521), .ZN(n5162) );
  AOI21_X1 U5512 ( .B1(n4996), .B2(n4999), .A(n4994), .ZN(n4993) );
  AND2_X1 U5513 ( .A1(n5689), .A2(n5281), .ZN(n5687) );
  INV_X1 U5514 ( .A(n5074), .ZN(n4859) );
  INV_X1 U5515 ( .A(n5257), .ZN(n5029) );
  NAND2_X1 U5516 ( .A1(n5703), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5777) );
  NAND2_X1 U5517 ( .A1(n5032), .A2(n5035), .ZN(n5491) );
  NAND2_X1 U5518 ( .A1(n5463), .A2(n5038), .ZN(n5032) );
  NAND2_X1 U5519 ( .A1(n5375), .A2(n5202), .ZN(n5388) );
  NAND2_X1 U5520 ( .A1(n4990), .A2(SI_0_), .ZN(n5296) );
  AOI21_X1 U5521 ( .B1(n4539), .B2(n5117), .A(n5113), .ZN(n5112) );
  INV_X1 U5522 ( .A(n8495), .ZN(n5113) );
  XNOR2_X1 U5523 ( .A(n7993), .B(n8622), .ZN(n7995) );
  AND4_X1 U5524 ( .A1(n6127), .A2(n6126), .A3(n6125), .A4(n6124), .ZN(n8398)
         );
  INV_X1 U5525 ( .A(n8527), .ZN(n8218) );
  NAND2_X1 U5526 ( .A1(n6141), .A2(n6140), .ZN(n8695) );
  AND4_X1 U5527 ( .A1(n6116), .A2(n6115), .A3(n6114), .A4(n6113), .ZN(n8729)
         );
  AND2_X1 U5528 ( .A1(n6611), .A2(n6612), .ZN(n4595) );
  INV_X1 U5529 ( .A(n8596), .ZN(n8344) );
  NAND2_X1 U5530 ( .A1(n6197), .A2(n6196), .ZN(n8645) );
  INV_X1 U5531 ( .A(n6666), .ZN(n8658) );
  NAND2_X1 U5532 ( .A1(n6166), .A2(n6165), .ZN(n8682) );
  INV_X1 U5533 ( .A(n6148), .ZN(n8704) );
  INV_X1 U5534 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9884) );
  OAI211_X1 U5535 ( .C1(n9876), .C2(n7215), .A(P2_IR_REG_0__SCAN_IN), .B(n4594), .ZN(n9900) );
  NAND2_X1 U5536 ( .A1(n9876), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4594) );
  NAND2_X1 U5537 ( .A1(n7941), .A2(n7942), .ZN(n7940) );
  NAND2_X1 U5538 ( .A1(n6121), .A2(n6120), .ZN(n8874) );
  NAND2_X1 U5539 ( .A1(n8610), .A2(n8823), .ZN(n4806) );
  NAND2_X1 U5540 ( .A1(n6200), .A2(n6199), .ZN(n8913) );
  NAND2_X1 U5541 ( .A1(n6151), .A2(n6150), .ZN(n8943) );
  OR2_X1 U5542 ( .A1(n6741), .A2(n6020), .ZN(n6023) );
  OR2_X1 U5543 ( .A1(n5869), .A2(n9892), .ZN(n5125) );
  NAND2_X1 U5544 ( .A1(n5869), .A2(n4519), .ZN(n5124) );
  NAND2_X1 U5545 ( .A1(n5869), .A2(n4836), .ZN(n5123) );
  NOR2_X1 U5546 ( .A1(n7883), .A2(n7820), .ZN(n5043) );
  NAND2_X1 U5547 ( .A1(n5318), .A2(n5317), .ZN(n7126) );
  AND2_X1 U5548 ( .A1(n4635), .A2(n4634), .ZN(n5317) );
  OR2_X1 U5549 ( .A1(n4723), .A2(n6484), .ZN(n4720) );
  NAND2_X1 U5550 ( .A1(n4600), .A2(n4598), .ZN(n6548) );
  INV_X1 U5551 ( .A(n4599), .ZN(n4598) );
  NOR2_X1 U5552 ( .A1(n6546), .A2(n6545), .ZN(n6547) );
  NOR2_X1 U5553 ( .A1(n6543), .A2(n6555), .ZN(n6546) );
  INV_X1 U5554 ( .A(n6544), .ZN(n6545) );
  INV_X1 U5555 ( .A(n5811), .ZN(n9369) );
  AOI21_X1 U5556 ( .B1(n4536), .B2(n4933), .A(n4527), .ZN(n4932) );
  NAND2_X1 U5557 ( .A1(n4536), .A2(n4518), .ZN(n4935) );
  NOR2_X1 U5558 ( .A1(n9369), .A2(n9645), .ZN(n5821) );
  INV_X1 U5559 ( .A(n9378), .ZN(n5750) );
  NAND2_X1 U5560 ( .A1(n4670), .A2(n4669), .ZN(n4673) );
  NAND2_X1 U5561 ( .A1(n4672), .A2(n8336), .ZN(n4671) );
  NOR2_X1 U5562 ( .A1(n8259), .A2(n4783), .ZN(n4782) );
  INV_X1 U5563 ( .A(n8262), .ZN(n4783) );
  NAND2_X1 U5564 ( .A1(n8275), .A2(n8326), .ZN(n4778) );
  AND2_X1 U5565 ( .A1(n8711), .A2(n8286), .ZN(n4631) );
  INV_X1 U5566 ( .A(n4704), .ZN(n4703) );
  OAI21_X1 U5567 ( .B1(n6401), .B2(n6468), .A(n6404), .ZN(n4704) );
  NAND2_X1 U5568 ( .A1(n4632), .A2(n4778), .ZN(n8287) );
  INV_X1 U5569 ( .A(n4631), .ZN(n4627) );
  AOI21_X1 U5570 ( .B1(n4631), .B2(n4626), .A(n8326), .ZN(n4625) );
  INV_X1 U5571 ( .A(n4778), .ZN(n4626) );
  OAI21_X1 U5572 ( .B1(n6422), .B2(n6410), .A(n6409), .ZN(n6411) );
  INV_X1 U5573 ( .A(n8297), .ZN(n4776) );
  NOR2_X1 U5574 ( .A1(n8693), .A2(n4552), .ZN(n4775) );
  OAI21_X1 U5575 ( .B1(n4712), .B2(n6468), .A(n4710), .ZN(n6431) );
  NOR2_X1 U5576 ( .A1(n4549), .A2(n4711), .ZN(n4710) );
  AOI21_X1 U5577 ( .B1(n4713), .B2(n6522), .A(n6419), .ZN(n4712) );
  NAND2_X1 U5578 ( .A1(n8321), .A2(n8320), .ZN(n4655) );
  AND2_X1 U5579 ( .A1(n8643), .A2(n8316), .ZN(n4656) );
  INV_X1 U5580 ( .A(n5689), .ZN(n5005) );
  INV_X1 U5581 ( .A(n5004), .ZN(n5003) );
  OAI21_X1 U5582 ( .B1(n5687), .B2(n5005), .A(n5788), .ZN(n5004) );
  INV_X1 U5583 ( .A(n5417), .ZN(n4770) );
  AND2_X1 U5584 ( .A1(n10012), .A2(n8556), .ZN(n8560) );
  NAND2_X1 U5585 ( .A1(n4532), .A2(n6454), .ZN(n4707) );
  INV_X1 U5586 ( .A(n5030), .ZN(n5027) );
  INV_X1 U5587 ( .A(n5639), .ZN(n5026) );
  INV_X1 U5588 ( .A(n5616), .ZN(n5251) );
  INV_X1 U5589 ( .A(SI_18_), .ZN(n10460) );
  INV_X1 U5590 ( .A(n4580), .ZN(n5011) );
  NAND2_X1 U5591 ( .A1(n5227), .A2(SI_13_), .ZN(n5228) );
  NAND2_X1 U5592 ( .A1(n8839), .A2(n8907), .ZN(n8153) );
  NAND2_X1 U5593 ( .A1(n4767), .A2(n4766), .ZN(n4765) );
  INV_X1 U5594 ( .A(n8333), .ZN(n8330) );
  NAND2_X1 U5595 ( .A1(n9891), .A2(n6947), .ZN(n9909) );
  NOR2_X1 U5596 ( .A1(n7761), .A2(n7760), .ZN(n7889) );
  OR2_X1 U5597 ( .A1(n7937), .A2(n4967), .ZN(n4966) );
  NOR2_X1 U5598 ( .A1(n7949), .A2(n7914), .ZN(n4967) );
  AND2_X1 U5599 ( .A1(n4965), .A2(n4964), .ZN(n8532) );
  NAND2_X1 U5600 ( .A1(n8531), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4964) );
  NAND2_X1 U5601 ( .A1(n9958), .A2(n4790), .ZN(n8575) );
  NAND2_X1 U5602 ( .A1(n8568), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4790) );
  NAND2_X1 U5603 ( .A1(n9991), .A2(n4786), .ZN(n8578) );
  NAND2_X1 U5604 ( .A1(n8567), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4786) );
  INV_X1 U5605 ( .A(n6128), .ZN(n4880) );
  OAI21_X1 U5606 ( .B1(n4883), .B2(n4880), .A(n8703), .ZN(n4879) );
  NAND2_X1 U5607 ( .A1(n4833), .A2(n4830), .ZN(n4829) );
  INV_X1 U5608 ( .A(n8172), .ZN(n4830) );
  INV_X1 U5609 ( .A(n4835), .ZN(n4827) );
  OR3_X1 U5610 ( .A1(n5951), .A2(n4867), .A3(n4862), .ZN(n4861) );
  NAND2_X1 U5611 ( .A1(n5927), .A2(n4546), .ZN(n4864) );
  NOR2_X1 U5612 ( .A1(n8526), .A2(n10047), .ZN(n4867) );
  AOI21_X1 U5613 ( .B1(n6211), .B2(n4875), .A(n4554), .ZN(n4872) );
  AND2_X1 U5614 ( .A1(n8308), .A2(n8666), .ZN(n6249) );
  AND2_X1 U5615 ( .A1(n6250), .A2(n8305), .ZN(n8309) );
  OR2_X1 U5616 ( .A1(n8306), .A2(n8665), .ZN(n6250) );
  OR2_X1 U5617 ( .A1(n8695), .A2(n6148), .ZN(n8300) );
  INV_X1 U5618 ( .A(n8343), .ZN(n6293) );
  OR2_X1 U5619 ( .A1(n8483), .A2(n6620), .ZN(n8286) );
  AND2_X1 U5620 ( .A1(n8159), .A2(n8267), .ZN(n8266) );
  OR2_X1 U5621 ( .A1(n6731), .A2(n6288), .ZN(n7068) );
  INV_X1 U5622 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6292) );
  AND2_X1 U5623 ( .A1(n5968), .A2(n5967), .ZN(n5970) );
  NOR2_X1 U5624 ( .A1(n5049), .A2(n4729), .ZN(n4728) );
  INV_X1 U5625 ( .A(n9717), .ZN(n4729) );
  INV_X1 U5626 ( .A(n7578), .ZN(n5044) );
  NAND2_X1 U5627 ( .A1(n6844), .A2(n7557), .ZN(n6847) );
  NOR2_X1 U5628 ( .A1(n5071), .A2(n5070), .ZN(n5069) );
  INV_X1 U5629 ( .A(n9176), .ZN(n5071) );
  NOR2_X1 U5630 ( .A1(n9165), .A2(n9166), .ZN(n5086) );
  NOR2_X1 U5631 ( .A1(n9390), .A2(n4844), .ZN(n4843) );
  INV_X1 U5632 ( .A(n4845), .ZN(n4844) );
  OR2_X1 U5633 ( .A1(n9601), .A2(n9071), .ZN(n6455) );
  NOR2_X1 U5634 ( .A1(n5543), .A2(n5542), .ZN(n9093) );
  NAND2_X1 U5635 ( .A1(n4848), .A2(n4522), .ZN(n7616) );
  AND2_X1 U5636 ( .A1(n7806), .A2(n4847), .ZN(n4849) );
  INV_X1 U5637 ( .A(n4850), .ZN(n4847) );
  INV_X1 U5638 ( .A(n7441), .ZN(n4848) );
  NAND2_X1 U5639 ( .A1(n7593), .A2(n4851), .ZN(n4850) );
  NAND2_X1 U5640 ( .A1(n6402), .A2(n7385), .ZN(n4931) );
  NAND2_X1 U5641 ( .A1(n7126), .A2(n6990), .ZN(n5715) );
  NAND2_X1 U5642 ( .A1(n9491), .A2(n5747), .ZN(n9492) );
  NAND2_X1 U5643 ( .A1(n9569), .A2(n4856), .ZN(n9549) );
  NAND2_X1 U5644 ( .A1(n9569), .A2(n9709), .ZN(n9568) );
  INV_X1 U5645 ( .A(n5677), .ZN(n4994) );
  NAND2_X1 U5646 ( .A1(n5159), .A2(n5158), .ZN(n5074) );
  AND2_X1 U5647 ( .A1(n5272), .A2(n5271), .ZN(n5663) );
  INV_X1 U5648 ( .A(SI_20_), .ZN(n10288) );
  INV_X1 U5649 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5555) );
  NOR2_X1 U5650 ( .A1(n5517), .A2(SI_15_), .ZN(n5014) );
  NAND2_X1 U5651 ( .A1(n5016), .A2(n4580), .ZN(n5015) );
  INV_X1 U5652 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n10406) );
  AOI21_X1 U5653 ( .B1(n5462), .B2(n5038), .A(n5036), .ZN(n5035) );
  INV_X1 U5654 ( .A(n5226), .ZN(n5036) );
  OR2_X1 U5655 ( .A1(n5449), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5450) );
  OR2_X1 U5656 ( .A1(n5434), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5449) );
  INV_X1 U5657 ( .A(n5401), .ZN(n4774) );
  INV_X1 U5658 ( .A(n5207), .ZN(n4773) );
  INV_X1 U5659 ( .A(n5211), .ZN(n4772) );
  AND2_X1 U5660 ( .A1(n5186), .A2(n5192), .ZN(n4988) );
  OAI21_X1 U5661 ( .B1(n4511), .B2(n4611), .A(n4610), .ZN(n5193) );
  NAND2_X1 U5662 ( .A1(n5859), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4610) );
  OR2_X1 U5663 ( .A1(n8411), .A2(n5117), .ZN(n5116) );
  INV_X1 U5664 ( .A(n6640), .ZN(n5117) );
  OR2_X1 U5665 ( .A1(n5986), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6013) );
  XNOR2_X1 U5666 ( .A(n6582), .B(n7072), .ZN(n6573) );
  INV_X1 U5667 ( .A(n5104), .ZN(n5103) );
  AND2_X1 U5668 ( .A1(n5108), .A2(n5101), .ZN(n5100) );
  NAND2_X1 U5669 ( .A1(n5104), .A2(n5102), .ZN(n5101) );
  NAND2_X1 U5670 ( .A1(n7671), .A2(n4557), .ZN(n7848) );
  NAND2_X1 U5671 ( .A1(n5975), .A2(n5974), .ZN(n5986) );
  INV_X1 U5672 ( .A(n8786), .ZN(n8453) );
  NAND2_X1 U5673 ( .A1(n5088), .A2(n5089), .ZN(n5098) );
  NOR2_X1 U5674 ( .A1(n5098), .A2(n8470), .ZN(n8467) );
  AND2_X1 U5675 ( .A1(n8190), .A2(n8338), .ZN(n8191) );
  NOR2_X1 U5676 ( .A1(n4677), .A2(n5020), .ZN(n5019) );
  INV_X1 U5677 ( .A(n5021), .ZN(n5020) );
  AOI21_X1 U5678 ( .B1(n8837), .B2(n8334), .A(n8343), .ZN(n5021) );
  OAI21_X1 U5679 ( .B1(n8339), .B2(n8636), .A(n4763), .ZN(n4762) );
  NOR2_X1 U5680 ( .A1(n8337), .A2(n4764), .ZN(n4763) );
  NAND2_X1 U5681 ( .A1(n4562), .A2(n8338), .ZN(n4764) );
  INV_X1 U5682 ( .A(n4761), .ZN(n4760) );
  OAI21_X1 U5683 ( .B1(n8341), .B2(n8154), .A(n8340), .ZN(n4761) );
  AND4_X1 U5684 ( .A1(n6080), .A2(n6079), .A3(n6078), .A4(n6077), .ZN(n8509)
         );
  AND4_X1 U5685 ( .A1(n6018), .A2(n6017), .A3(n6016), .A4(n6015), .ZN(n8403)
         );
  NAND2_X1 U5686 ( .A1(n6231), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5919) );
  NOR2_X1 U5687 ( .A1(n4691), .A2(n5849), .ZN(n4690) );
  INV_X1 U5688 ( .A(n6965), .ZN(n4691) );
  NAND2_X1 U5689 ( .A1(n4692), .A2(n6965), .ZN(n4693) );
  NAND2_X1 U5690 ( .A1(n4963), .A2(n4962), .ZN(n4687) );
  INV_X1 U5691 ( .A(n6969), .ZN(n4963) );
  NAND2_X1 U5692 ( .A1(n6969), .A2(n6968), .ZN(n6972) );
  NAND2_X1 U5693 ( .A1(n6971), .A2(n6970), .ZN(n7037) );
  NAND2_X1 U5694 ( .A1(n9923), .A2(n6972), .ZN(n6970) );
  AND2_X1 U5695 ( .A1(n4689), .A2(n7192), .ZN(n7039) );
  NAND2_X1 U5696 ( .A1(n7038), .A2(n7182), .ZN(n7192) );
  NAND3_X1 U5697 ( .A1(n4689), .A2(n7192), .A3(P2_REG2_REG_5__SCAN_IN), .ZN(
        n7194) );
  INV_X1 U5698 ( .A(n4986), .ZN(n7749) );
  INV_X1 U5699 ( .A(n4688), .ZN(n7913) );
  NOR2_X1 U5700 ( .A1(n7890), .A2(n7889), .ZN(n7944) );
  NAND2_X1 U5701 ( .A1(n7940), .A2(n4787), .ZN(n7906) );
  OR2_X1 U5702 ( .A1(n7949), .A2(n5985), .ZN(n4787) );
  AOI21_X1 U5703 ( .B1(n8550), .B2(n8549), .A(n8548), .ZN(n9945) );
  XNOR2_X1 U5704 ( .A(n8532), .B(n9942), .ZN(n9951) );
  NAND2_X1 U5705 ( .A1(n9946), .A2(n8573), .ZN(n9959) );
  NAND2_X1 U5706 ( .A1(n9962), .A2(n9963), .ZN(n9961) );
  NAND2_X1 U5707 ( .A1(n9959), .A2(n9960), .ZN(n9958) );
  XNOR2_X1 U5708 ( .A(n8575), .B(n9974), .ZN(n9976) );
  AND2_X1 U5709 ( .A1(n4973), .A2(n4544), .ZN(n10001) );
  NOR2_X1 U5710 ( .A1(n10001), .A2(n10000), .ZN(n9999) );
  NAND2_X1 U5711 ( .A1(n9992), .A2(n9993), .ZN(n9991) );
  NAND2_X1 U5712 ( .A1(n10013), .A2(n10014), .ZN(n10012) );
  XNOR2_X1 U5713 ( .A(n8578), .B(n10009), .ZN(n10011) );
  NAND2_X1 U5714 ( .A1(n10011), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n10010) );
  AOI21_X1 U5715 ( .B1(n8540), .B2(n4980), .A(n4979), .ZN(n4978) );
  NAND2_X1 U5716 ( .A1(n8597), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n4798) );
  NAND2_X1 U5717 ( .A1(n6143), .A2(n6142), .ZN(n6152) );
  NOR2_X1 U5718 ( .A1(n4822), .A2(n4820), .ZN(n4819) );
  INV_X1 U5719 ( .A(n8296), .ZN(n4820) );
  AND2_X1 U5720 ( .A1(n6133), .A2(n10491), .ZN(n6143) );
  NOR2_X1 U5721 ( .A1(n6122), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6133) );
  INV_X1 U5722 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10491) );
  INV_X1 U5723 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10450) );
  NAND2_X1 U5724 ( .A1(n6099), .A2(n10450), .ZN(n6111) );
  AND2_X1 U5725 ( .A1(n6086), .A2(n8429), .ZN(n6099) );
  AND4_X1 U5726 ( .A1(n6066), .A2(n6065), .A3(n6064), .A4(n6063), .ZN(n8754)
         );
  AND4_X1 U5727 ( .A1(n6091), .A2(n6090), .A3(n6089), .A4(n6088), .ZN(n8756)
         );
  INV_X1 U5728 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10462) );
  INV_X1 U5729 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10509) );
  OR2_X1 U5730 ( .A1(n6013), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6024) );
  NOR2_X1 U5731 ( .A1(n6024), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6036) );
  AND2_X1 U5732 ( .A1(n5954), .A2(n7518), .ZN(n5975) );
  NAND2_X1 U5733 ( .A1(n4868), .A2(n4866), .ZN(n7656) );
  INV_X1 U5734 ( .A(n4867), .ZN(n4866) );
  OR2_X1 U5735 ( .A1(n5929), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U5736 ( .A1(n5927), .A2(n5926), .ZN(n7487) );
  NAND2_X1 U5737 ( .A1(n4800), .A2(n8219), .ZN(n7425) );
  AND3_X1 U5738 ( .A1(n7208), .A2(n10078), .A3(n6259), .ZN(n8823) );
  AND2_X1 U5739 ( .A1(n8605), .A2(n8604), .ZN(n8905) );
  AND2_X1 U5740 ( .A1(n6181), .A2(n6180), .ZN(n6641) );
  AND2_X1 U5741 ( .A1(n8290), .A2(n8711), .ZN(n8180) );
  INV_X1 U5742 ( .A(n8270), .ZN(n8764) );
  INV_X1 U5743 ( .A(n8266), .ZN(n8781) );
  NOR2_X1 U5744 ( .A1(n6688), .A2(n4511), .ZN(n4836) );
  NAND2_X1 U5745 ( .A1(n6658), .A2(n7067), .ZN(n6661) );
  NAND2_X1 U5746 ( .A1(n6290), .A2(n6289), .ZN(n6679) );
  NOR2_X1 U5747 ( .A1(n5126), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4890) );
  INV_X1 U5748 ( .A(n5839), .ZN(n5131) );
  XNOR2_X1 U5749 ( .A(n6291), .B(n6292), .ZN(n6680) );
  OR2_X1 U5750 ( .A1(n5935), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5947) );
  INV_X1 U5751 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5920) );
  INV_X1 U5752 ( .A(n4748), .ZN(n4747) );
  AOI21_X1 U5753 ( .B1(n4750), .B2(n4749), .A(n4753), .ZN(n4748) );
  INV_X1 U5754 ( .A(n5076), .ZN(n4749) );
  INV_X1 U5755 ( .A(n4751), .ZN(n4746) );
  NAND2_X1 U5756 ( .A1(n9214), .A2(n8129), .ZN(n6984) );
  NAND2_X1 U5757 ( .A1(n9152), .A2(n9156), .ZN(n9041) );
  NOR2_X1 U5758 ( .A1(n4752), .A2(n8133), .ZN(n4751) );
  OR2_X1 U5759 ( .A1(n5409), .A2(n5408), .ZN(n5424) );
  INV_X1 U5760 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5423) );
  XNOR2_X1 U5761 ( .A(n4742), .B(n8354), .ZN(n6860) );
  OAI21_X1 U5762 ( .B1(n6981), .B2(n9783), .A(n6858), .ZN(n4742) );
  INV_X1 U5763 ( .A(n9069), .ZN(n5080) );
  NAND2_X1 U5764 ( .A1(n9102), .A2(n8111), .ZN(n5082) );
  NAND2_X1 U5765 ( .A1(n9104), .A2(n5083), .ZN(n5081) );
  INV_X1 U5766 ( .A(n5069), .ZN(n5062) );
  NOR2_X1 U5767 ( .A1(n9176), .A2(n9177), .ZN(n5067) );
  OR2_X1 U5768 ( .A1(n5424), .A2(n5423), .ZN(n5438) );
  OR2_X1 U5769 ( .A1(n5599), .A2(n5598), .ZN(n5612) );
  OR2_X1 U5770 ( .A1(n5612), .A2(n9120), .ZN(n5621) );
  NAND2_X1 U5771 ( .A1(n9041), .A2(n9042), .ZN(n9040) );
  NAND2_X1 U5772 ( .A1(n5057), .A2(n9059), .ZN(n9132) );
  NAND2_X1 U5773 ( .A1(n7799), .A2(n9058), .ZN(n5057) );
  NOR2_X1 U5774 ( .A1(n5621), .A2(n9053), .ZN(n5630) );
  CLKBUF_X1 U5775 ( .A(n8005), .Z(n7799) );
  NOR2_X1 U5776 ( .A1(n5049), .A2(n5048), .ZN(n5047) );
  INV_X1 U5777 ( .A(n4550), .ZN(n5048) );
  CLKBUF_X1 U5778 ( .A(n7796), .Z(n7785) );
  NAND2_X1 U5779 ( .A1(n5086), .A2(n5079), .ZN(n5075) );
  NAND2_X1 U5780 ( .A1(n4718), .A2(n4716), .ZN(n6487) );
  AOI21_X1 U5781 ( .B1(n4721), .B2(n4717), .A(n6840), .ZN(n4716) );
  AND2_X1 U5782 ( .A1(n6542), .A2(n7557), .ZN(n6845) );
  AND4_X1 U5783 ( .A1(n5686), .A2(n5685), .A3(n5684), .A4(n5683), .ZN(n9072)
         );
  AND4_X1 U5784 ( .A1(n5502), .A2(n5501), .A3(n5500), .A4(n5499), .ZN(n8018)
         );
  AND4_X1 U5785 ( .A1(n5488), .A2(n5487), .A3(n5486), .A4(n5485), .ZN(n8009)
         );
  AND4_X1 U5786 ( .A1(n5474), .A2(n5473), .A3(n5472), .A4(n5471), .ZN(n7789)
         );
  AND4_X1 U5787 ( .A1(n5461), .A2(n5460), .A3(n5459), .A4(n5458), .ZN(n7780)
         );
  AND4_X1 U5788 ( .A1(n5442), .A2(n5441), .A3(n5440), .A4(n5439), .ZN(n7574)
         );
  OR2_X1 U5789 ( .A1(n5602), .A2(n5328), .ZN(n5329) );
  AOI21_X1 U5790 ( .B1(n6795), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6808), .ZN(
        n6796) );
  AOI21_X1 U5791 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9292), .A(n9291), .ZN(
        n9315) );
  AND2_X1 U5792 ( .A1(n6872), .A2(n9232), .ZN(n9181) );
  OAI21_X1 U5793 ( .B1(n6474), .B2(n4900), .A(n4897), .ZN(n4896) );
  NAND2_X1 U5794 ( .A1(n4900), .A2(n4898), .ZN(n4897) );
  NAND2_X1 U5795 ( .A1(n4903), .A2(n4899), .ZN(n4898) );
  NAND2_X1 U5796 ( .A1(n4937), .A2(n4516), .ZN(n4936) );
  NAND2_X1 U5797 ( .A1(n4516), .A2(n4934), .ZN(n4933) );
  NAND2_X1 U5798 ( .A1(n4518), .A2(n9400), .ZN(n4934) );
  NAND2_X1 U5799 ( .A1(n4681), .A2(n4543), .ZN(n4938) );
  NAND2_X1 U5800 ( .A1(n9432), .A2(n4843), .ZN(n9387) );
  NOR2_X1 U5801 ( .A1(n5682), .A2(n9172), .ZN(n5681) );
  NAND2_X1 U5802 ( .A1(n9432), .A2(n9658), .ZN(n9415) );
  NOR2_X1 U5803 ( .A1(n9608), .A2(n9455), .ZN(n9446) );
  AND2_X1 U5804 ( .A1(n9436), .A2(n9446), .ZN(n9432) );
  NAND2_X1 U5805 ( .A1(n6455), .A2(n6456), .ZN(n9429) );
  OAI21_X1 U5806 ( .B1(n4534), .B2(n4941), .A(n9462), .ZN(n4940) );
  AND2_X1 U5807 ( .A1(n6450), .A2(n6451), .ZN(n9443) );
  AOI21_X1 U5808 ( .B1(n4943), .B2(n4649), .A(n4542), .ZN(n4648) );
  INV_X1 U5809 ( .A(n4943), .ZN(n4650) );
  NAND2_X1 U5810 ( .A1(n9569), .A2(n4524), .ZN(n9514) );
  INV_X1 U5811 ( .A(n4854), .ZN(n4853) );
  AOI22_X1 U5812 ( .A1(n4921), .A2(n4928), .B1(n4924), .B2(n4926), .ZN(n4917)
         );
  OR2_X1 U5813 ( .A1(n7616), .A2(n9137), .ZN(n7737) );
  NOR2_X2 U5814 ( .A1(n7737), .A2(n7740), .ZN(n9569) );
  AND2_X1 U5815 ( .A1(n6515), .A2(n6416), .ZN(n7730) );
  NOR2_X1 U5816 ( .A1(n5495), .A2(n5167), .ZN(n5510) );
  INV_X1 U5817 ( .A(n5724), .ZN(n4955) );
  NAND2_X1 U5818 ( .A1(n7709), .A2(n7708), .ZN(n7707) );
  AOI21_X1 U5819 ( .B1(n7530), .B2(n4640), .A(n4560), .ZN(n4639) );
  INV_X1 U5820 ( .A(n5443), .ZN(n4640) );
  NAND2_X1 U5821 ( .A1(n7528), .A2(n6360), .ZN(n7690) );
  INV_X1 U5822 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5468) );
  NAND2_X1 U5823 ( .A1(n4848), .A2(n4849), .ZN(n7685) );
  INV_X1 U5824 ( .A(n7690), .ZN(n7529) );
  NOR2_X1 U5825 ( .A1(n7441), .A2(n7576), .ZN(n7534) );
  NAND2_X1 U5826 ( .A1(n7395), .A2(n9823), .ZN(n7440) );
  NOR2_X1 U5827 ( .A1(n9748), .A2(n7381), .ZN(n7395) );
  INV_X1 U5828 ( .A(n9766), .ZN(n4841) );
  NAND2_X1 U5829 ( .A1(n9765), .A2(n9344), .ZN(n6886) );
  NAND2_X1 U5830 ( .A1(n6845), .A2(n6844), .ZN(n7220) );
  NOR2_X1 U5831 ( .A1(n7227), .A2(n7126), .ZN(n9767) );
  NAND2_X1 U5832 ( .A1(n7221), .A2(n5714), .ZN(n7117) );
  INV_X1 U5833 ( .A(n9168), .ZN(n9180) );
  INV_X1 U5834 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4838) );
  INV_X1 U5835 ( .A(n9691), .ZN(n4837) );
  INV_X1 U5836 ( .A(n6709), .ZN(n5593) );
  NAND2_X1 U5837 ( .A1(n5680), .A2(n5679), .ZN(n9402) );
  INV_X1 U5838 ( .A(n7126), .ZN(n9789) );
  INV_X1 U5839 ( .A(n9845), .ZN(n9805) );
  XNOR2_X1 U5840 ( .A(n6323), .B(n5793), .ZN(n8142) );
  XNOR2_X1 U5841 ( .A(n5757), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U5842 ( .A1(n5756), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5757) );
  XNOR2_X1 U5843 ( .A(n5678), .B(n5677), .ZN(n9014) );
  OAI21_X1 U5844 ( .B1(n5268), .B2(n4999), .A(n4996), .ZN(n5678) );
  NAND2_X1 U5845 ( .A1(n5755), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5759) );
  INV_X1 U5846 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U5847 ( .A1(n5591), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5592) );
  CLKBUF_X1 U5848 ( .A(n5577), .Z(n5574) );
  INV_X1 U5849 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5147) );
  NAND2_X1 U5850 ( .A1(n5444), .A2(n5222), .ZN(n5448) );
  AND2_X1 U5851 ( .A1(n5396), .A2(n5404), .ZN(n6792) );
  NAND2_X1 U5852 ( .A1(n5188), .A2(SI_3_), .ZN(n5192) );
  CLKBUF_X1 U5853 ( .A(n5354), .Z(n5355) );
  NAND2_X1 U5854 ( .A1(n5187), .A2(n5186), .ZN(n5338) );
  OAI21_X1 U5855 ( .B1(P1_RD_REG_SCAN_IN), .B2(P1_ADDR_REG_19__SCAN_IN), .A(
        n5176), .ZN(n5179) );
  INV_X1 U5856 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5176) );
  OAI21_X1 U5857 ( .B1(n5093), .B2(n4587), .A(n5092), .ZN(n5091) );
  INV_X1 U5858 ( .A(n8450), .ZN(n5092) );
  XNOR2_X1 U5859 ( .A(n6606), .B(n8522), .ZN(n7928) );
  AOI21_X1 U5860 ( .B1(n5120), .B2(n8486), .A(n4583), .ZN(n5119) );
  OR2_X1 U5861 ( .A1(n7993), .A2(n8622), .ZN(n7994) );
  INV_X1 U5862 ( .A(n8523), .ZN(n7676) );
  AND2_X1 U5863 ( .A1(n5105), .A2(n4545), .ZN(n8395) );
  NAND2_X1 U5864 ( .A1(n8443), .A2(n8444), .ZN(n5105) );
  INV_X1 U5865 ( .A(n8682), .ZN(n8414) );
  XNOR2_X1 U5866 ( .A(n6635), .B(n8682), .ZN(n8437) );
  AND2_X1 U5867 ( .A1(n7298), .A2(n6587), .ZN(n7308) );
  NAND2_X1 U5868 ( .A1(n7671), .A2(n6601), .ZN(n7850) );
  AND2_X1 U5869 ( .A1(n7132), .A2(n8351), .ZN(n8511) );
  NAND2_X1 U5870 ( .A1(n5090), .A2(n5093), .ZN(n8452) );
  NAND2_X1 U5871 ( .A1(n5095), .A2(n5096), .ZN(n5090) );
  INV_X1 U5872 ( .A(n5098), .ZN(n5096) );
  NAND2_X1 U5873 ( .A1(n5111), .A2(n6627), .ZN(n8460) );
  NAND2_X1 U5874 ( .A1(n5107), .A2(n5106), .ZN(n5111) );
  INV_X1 U5875 ( .A(n8394), .ZN(n5106) );
  INV_X1 U5876 ( .A(n8395), .ZN(n5107) );
  OAI21_X1 U5877 ( .B1(n8418), .B2(n8486), .A(n5120), .ZN(n8484) );
  INV_X1 U5878 ( .A(n8511), .ZN(n8497) );
  NAND2_X1 U5879 ( .A1(n7457), .A2(n6593), .ZN(n7606) );
  NAND2_X1 U5880 ( .A1(n6649), .A2(n8819), .ZN(n8501) );
  OR2_X1 U5881 ( .A1(n6665), .A2(n6662), .ZN(n8510) );
  NAND2_X1 U5882 ( .A1(n5115), .A2(n6640), .ZN(n8493) );
  NAND2_X1 U5883 ( .A1(n8410), .A2(n8411), .ZN(n5115) );
  INV_X1 U5884 ( .A(n8503), .ZN(n8505) );
  INV_X1 U5885 ( .A(n8476), .ZN(n8514) );
  XNOR2_X1 U5886 ( .A(n6220), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8348) );
  INV_X1 U5887 ( .A(n8647), .ZN(n8671) );
  INV_X1 U5888 ( .A(n8509), .ZN(n8766) );
  INV_X1 U5889 ( .A(n8754), .ZN(n8774) );
  NOR2_X1 U5890 ( .A1(n4509), .A2(n7210), .ZN(n5864) );
  NAND2_X1 U5891 ( .A1(n4789), .A2(n9884), .ZN(n4788) );
  NAND2_X1 U5892 ( .A1(n9876), .A2(n9878), .ZN(n4789) );
  OAI22_X1 U5893 ( .A1(n7175), .A2(n7174), .B1(n4960), .B2(n7173), .ZN(n7179)
         );
  AND2_X1 U5894 ( .A1(n7511), .A2(n4698), .ZN(n7467) );
  NOR2_X1 U5895 ( .A1(n7497), .A2(n4608), .ZN(n7504) );
  AND2_X1 U5896 ( .A1(n7498), .A2(n4959), .ZN(n4608) );
  AND2_X1 U5897 ( .A1(n4688), .A2(n4569), .ZN(n7939) );
  INV_X1 U5898 ( .A(n4984), .ZN(n7911) );
  NOR2_X1 U5899 ( .A1(n7939), .A2(n7938), .ZN(n7937) );
  NAND2_X1 U5900 ( .A1(n7904), .A2(n7905), .ZN(n7941) );
  XNOR2_X1 U5901 ( .A(n7906), .B(n7965), .ZN(n7956) );
  NOR2_X1 U5902 ( .A1(n7897), .A2(n7961), .ZN(n8550) );
  INV_X1 U5903 ( .A(n4701), .ZN(n7921) );
  INV_X1 U5904 ( .A(n4973), .ZN(n9982) );
  NAND2_X1 U5905 ( .A1(n6960), .A2(n6959), .ZN(n10008) );
  OR2_X1 U5906 ( .A1(n8540), .A2(n8591), .ZN(n4982) );
  INV_X1 U5907 ( .A(n4700), .ZN(n8539) );
  AND2_X1 U5908 ( .A1(n4978), .A2(n4981), .ZN(n4976) );
  XNOR2_X1 U5909 ( .A(n4797), .B(n8600), .ZN(n4796) );
  NAND2_X1 U5910 ( .A1(n4795), .A2(n4794), .ZN(n4793) );
  NAND2_X1 U5911 ( .A1(n4799), .A2(n4798), .ZN(n4797) );
  AND2_X1 U5912 ( .A1(n8606), .A2(n6204), .ZN(n8629) );
  OR2_X1 U5913 ( .A1(n6190), .A2(n6183), .ZN(n8651) );
  NOR2_X1 U5914 ( .A1(n4882), .A2(n4881), .ZN(n8717) );
  NAND2_X1 U5915 ( .A1(n6072), .A2(n6071), .ZN(n8887) );
  AND2_X1 U5916 ( .A1(n5999), .A2(n5998), .ZN(n7834) );
  NAND2_X1 U5917 ( .A1(n4831), .A2(n4833), .ZN(n7809) );
  NAND2_X1 U5918 ( .A1(n7655), .A2(n4835), .ZN(n4831) );
  NAND2_X1 U5919 ( .A1(n4832), .A2(n8237), .ZN(n7639) );
  OR2_X1 U5920 ( .A1(n7655), .A2(n8236), .ZN(n4832) );
  INV_X1 U5921 ( .A(n8819), .ZN(n8769) );
  INV_X1 U5922 ( .A(n8733), .ZN(n8813) );
  NAND2_X1 U5923 ( .A1(n7053), .A2(n6237), .ZN(n8818) );
  NAND2_X1 U5924 ( .A1(n7067), .A2(n7069), .ZN(n8819) );
  INV_X1 U5925 ( .A(n6575), .ZN(n7218) );
  OR2_X1 U5926 ( .A1(n7214), .A2(n8820), .ZN(n8733) );
  NOR2_X1 U5927 ( .A1(n8625), .A2(n8624), .ZN(n8626) );
  NOR2_X1 U5928 ( .A1(n8622), .A2(n8755), .ZN(n8625) );
  AOI21_X1 U5929 ( .B1(n9001), .B2(n8148), .A(n5006), .ZN(n8907) );
  NOR2_X1 U5930 ( .A1(n5905), .A2(n5007), .ZN(n5006) );
  INV_X1 U5931 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5007) );
  AOI21_X1 U5932 ( .B1(n8146), .B2(n8148), .A(n8145), .ZN(n8910) );
  AND2_X1 U5933 ( .A1(n4877), .A2(n4876), .ZN(n8635) );
  INV_X1 U5934 ( .A(n6641), .ZN(n8925) );
  NAND2_X1 U5935 ( .A1(n4808), .A2(n8315), .ZN(n8642) );
  NAND2_X1 U5936 ( .A1(n6159), .A2(n6158), .ZN(n8937) );
  NAND2_X1 U5937 ( .A1(n4885), .A2(n6149), .ZN(n8681) );
  NAND2_X1 U5938 ( .A1(n8715), .A2(n6128), .ZN(n8702) );
  NAND2_X1 U5939 ( .A1(n4821), .A2(n8296), .ZN(n8701) );
  NAND2_X1 U5940 ( .A1(n6110), .A2(n6109), .ZN(n8391) );
  INV_X1 U5941 ( .A(n8483), .ZN(n8965) );
  NAND2_X1 U5942 ( .A1(n6085), .A2(n6084), .ZN(n8968) );
  NAND2_X1 U5943 ( .A1(n6062), .A2(n6061), .ZN(n8978) );
  NAND2_X1 U5944 ( .A1(n6050), .A2(n6049), .ZN(n8984) );
  NAND2_X1 U5945 ( .A1(n6035), .A2(n6034), .ZN(n8990) );
  NAND2_X1 U5946 ( .A1(n4814), .A2(n4815), .ZN(n8794) );
  OR2_X1 U5947 ( .A1(n7838), .A2(n4818), .ZN(n4814) );
  OAI22_X1 U5948 ( .A1(n6731), .A2(P2_D_REG_1__SCAN_IN), .B1(n6274), .B2(n6290), .ZN(n7062) );
  AND2_X1 U5949 ( .A1(n6680), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7131) );
  NAND2_X1 U5950 ( .A1(n6731), .A2(n7067), .ZN(n6735) );
  XNOR2_X1 U5951 ( .A(n6268), .B(n6267), .ZN(n7881) );
  NAND2_X1 U5952 ( .A1(n6266), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6268) );
  INV_X1 U5953 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7718) );
  INV_X1 U5954 ( .A(n8348), .ZN(n7717) );
  INV_X1 U5955 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7598) );
  INV_X1 U5956 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7420) );
  INV_X1 U5957 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7236) );
  OR2_X1 U5958 ( .A1(n6010), .A2(n6009), .ZN(n7917) );
  INV_X1 U5959 ( .A(n7519), .ZN(n7750) );
  AOI21_X1 U5960 ( .B1(n4972), .B2(n4970), .A(n4969), .ZN(n4968) );
  NOR2_X1 U5961 ( .A1(n9002), .A2(n4971), .ZN(n4970) );
  NAND2_X1 U5962 ( .A1(n5862), .A2(n4972), .ZN(n9892) );
  NAND2_X1 U5963 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5860) );
  XNOR2_X1 U5964 ( .A(n5779), .B(n10519), .ZN(n6876) );
  CLKBUF_X1 U5965 ( .A(n7342), .Z(n7341) );
  CLKBUF_X1 U5966 ( .A(n7561), .Z(n7343) );
  AOI21_X1 U5967 ( .B1(n4747), .B2(n4746), .A(n9699), .ZN(n4744) );
  NAND2_X1 U5968 ( .A1(n4750), .A2(n4746), .ZN(n4745) );
  AOI21_X1 U5969 ( .B1(n4740), .B2(n4739), .A(n4738), .ZN(n4737) );
  NAND2_X1 U5970 ( .A1(n5081), .A2(n5082), .ZN(n9070) );
  NAND2_X1 U5971 ( .A1(n4757), .A2(n5063), .ZN(n8045) );
  INV_X1 U5972 ( .A(n5059), .ZN(n9079) );
  OAI21_X1 U5973 ( .B1(n5068), .B2(n5061), .A(n5060), .ZN(n5059) );
  INV_X1 U5974 ( .A(n5067), .ZN(n5060) );
  NAND2_X1 U5975 ( .A1(n9021), .A2(n5062), .ZN(n5061) );
  NAND2_X1 U5976 ( .A1(n4757), .A2(n4517), .ZN(n9087) );
  AOI21_X1 U5977 ( .B1(n9104), .B2(n9103), .A(n9102), .ZN(n9106) );
  NAND2_X1 U5978 ( .A1(n7164), .A2(n7163), .ZN(n7259) );
  NAND2_X1 U5979 ( .A1(n5055), .A2(n9131), .ZN(n5054) );
  NAND2_X1 U5980 ( .A1(n6922), .A2(n6923), .ZN(n6989) );
  INV_X1 U5981 ( .A(n9722), .ZN(n9703) );
  INV_X1 U5982 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9184) );
  INV_X1 U5983 ( .A(n9727), .ZN(n9187) );
  AND4_X1 U5984 ( .A1(n5744), .A2(n5743), .A3(n5742), .A4(n5741), .ZN(n7077)
         );
  AND2_X1 U5985 ( .A1(n5322), .A2(n5323), .ZN(n4597) );
  AOI21_X1 U5986 ( .B1(n7019), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7015), .ZN(
        n7018) );
  CLKBUF_X1 U5987 ( .A(n6542), .Z(n9344) );
  NOR2_X1 U5988 ( .A1(n4839), .A2(n9850), .ZN(n9352) );
  OR2_X1 U5989 ( .A1(n9360), .A2(n9359), .ZN(n9581) );
  NAND2_X1 U5990 ( .A1(n4905), .A2(n4906), .ZN(n5797) );
  NAND2_X1 U5991 ( .A1(n4679), .A2(n4938), .ZN(n9586) );
  NAND2_X1 U5992 ( .A1(n4680), .A2(n4937), .ZN(n4679) );
  NAND2_X1 U5993 ( .A1(n4681), .A2(n4518), .ZN(n4680) );
  NAND2_X1 U5994 ( .A1(n9471), .A2(n6443), .ZN(n9463) );
  NAND2_X1 U5995 ( .A1(n5733), .A2(n6386), .ZN(n9473) );
  NAND2_X1 U5996 ( .A1(n4945), .A2(n5606), .ZN(n9486) );
  NAND2_X1 U5997 ( .A1(n5588), .A2(n4651), .ZN(n4945) );
  NAND2_X1 U5998 ( .A1(n5588), .A2(n5587), .ZN(n9500) );
  NAND2_X1 U5999 ( .A1(n4957), .A2(n5570), .ZN(n9513) );
  NAND2_X1 U6000 ( .A1(n4646), .A2(n5550), .ZN(n9527) );
  NAND2_X1 U6001 ( .A1(n4909), .A2(n4913), .ZN(n9544) );
  INV_X1 U6002 ( .A(n9565), .ZN(n9759) );
  INV_X1 U6003 ( .A(n9452), .ZN(n9730) );
  NAND2_X1 U6004 ( .A1(n7527), .A2(n7530), .ZN(n7526) );
  NAND2_X1 U6005 ( .A1(n4643), .A2(n5443), .ZN(n7527) );
  NAND2_X1 U6006 ( .A1(n5431), .A2(n4641), .ZN(n4643) );
  NAND2_X1 U6007 ( .A1(n5431), .A2(n7429), .ZN(n7403) );
  NAND2_X1 U6008 ( .A1(n4948), .A2(n5416), .ZN(n7430) );
  OR2_X1 U6009 ( .A1(n6886), .A2(n9775), .ZN(n9565) );
  INV_X1 U6010 ( .A(n9556), .ZN(n9770) );
  OR2_X1 U6011 ( .A1(n9773), .A2(n9344), .ZN(n9570) );
  INV_X1 U6012 ( .A(n7228), .ZN(n7005) );
  INV_X1 U6013 ( .A(n9761), .ZN(n9731) );
  INV_X1 U6014 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n4684) );
  NOR2_X1 U6015 ( .A1(n9369), .A2(n9675), .ZN(n5812) );
  INV_X1 U6016 ( .A(n9402), .ZN(n9654) );
  INV_X1 U6017 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5160) );
  NAND2_X1 U6018 ( .A1(n5002), .A2(n5689), .ZN(n5789) );
  MUX2_X1 U6019 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5285), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n5286) );
  XNOR2_X1 U6020 ( .A(n5759), .B(n5758), .ZN(n7883) );
  NAND2_X1 U6021 ( .A1(n5754), .A2(n5755), .ZN(n7820) );
  NAND2_X1 U6022 ( .A1(n5024), .A2(n5028), .ZN(n5640) );
  NAND2_X1 U6023 ( .A1(n5618), .A2(n5030), .ZN(n5024) );
  INV_X1 U6024 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10446) );
  INV_X1 U6025 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7612) );
  INV_X1 U6026 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7422) );
  NAND2_X1 U6027 ( .A1(n5039), .A2(n5038), .ZN(n5478) );
  NAND2_X1 U6028 ( .A1(n5402), .A2(n5401), .ZN(n5403) );
  INV_X1 U6029 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n10542) );
  INV_X2 U6030 ( .A(n8528), .ZN(P2_U3893) );
  NOR2_X1 U6031 ( .A1(n9877), .A2(n4788), .ZN(n9880) );
  XNOR2_X1 U6032 ( .A(n4700), .B(n8540), .ZN(n4699) );
  OAI21_X1 U6033 ( .B1(n4802), .B2(n5143), .A(n8845), .ZN(n8846) );
  NAND2_X1 U6034 ( .A1(n10098), .A2(n8844), .ZN(n8845) );
  NOR2_X1 U6035 ( .A1(n5138), .A2(n6303), .ZN(n6304) );
  NOR2_X1 U6036 ( .A1(n5143), .A2(n8611), .ZN(n8843) );
  INV_X1 U6037 ( .A(n6562), .ZN(n6563) );
  OAI21_X1 U6038 ( .B1(n6561), .B2(n6560), .A(n6559), .ZN(n6562) );
  NOR2_X1 U6039 ( .A1(n5821), .A2(n5823), .ZN(n5824) );
  AOI21_X1 U6040 ( .B1(n8368), .B2(n7701), .A(n4603), .ZN(n4602) );
  NOR2_X1 U6041 ( .A1(n9875), .A2(n9585), .ZN(n4603) );
  INV_X1 U6042 ( .A(n4683), .ZN(n4682) );
  NAND2_X1 U6043 ( .A1(n9650), .A2(n9875), .ZN(n4685) );
  INV_X1 U6044 ( .A(n4612), .ZN(P1_U3517) );
  AOI21_X1 U6045 ( .B1(n9650), .B2(n9858), .A(n4613), .ZN(n4612) );
  OAI21_X1 U6046 ( .B1(n5748), .B2(n9675), .A(n4614), .ZN(n4613) );
  NAND2_X1 U6047 ( .A1(n5809), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n4614) );
  INV_X1 U6048 ( .A(n5327), .ZN(n5650) );
  AND2_X1 U6049 ( .A1(n8286), .A2(n8285), .ZN(n4515) );
  OR2_X1 U6050 ( .A1(n9390), .A2(n9193), .ZN(n4516) );
  AND2_X1 U6051 ( .A1(n5063), .A2(n8046), .ZN(n4517) );
  INV_X1 U6052 ( .A(n8332), .ZN(n4767) );
  NAND3_X1 U6053 ( .A1(n5073), .A2(n5058), .A3(n4657), .ZN(n4658) );
  INV_X1 U6054 ( .A(n7708), .ZN(n4923) );
  NAND2_X1 U6055 ( .A1(n6476), .A2(n6477), .ZN(n6474) );
  INV_X1 U6056 ( .A(n6474), .ZN(n4899) );
  NAND2_X1 U6057 ( .A1(n9402), .A2(n9194), .ZN(n4518) );
  AND2_X1 U6058 ( .A1(n4511), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4519) );
  AND2_X1 U6059 ( .A1(n6492), .A2(n6468), .ZN(n4520) );
  INV_X1 U6060 ( .A(n6318), .ZN(n4901) );
  INV_X1 U6061 ( .A(n8468), .ZN(n5089) );
  AND2_X1 U6062 ( .A1(n4852), .A2(n4849), .ZN(n4522) );
  NAND2_X1 U6063 ( .A1(n9608), .A2(n9145), .ZN(n4523) );
  NOR2_X1 U6064 ( .A1(n4853), .A2(n9632), .ZN(n4524) );
  NOR2_X1 U6065 ( .A1(n8059), .A2(n5050), .ZN(n4525) );
  INV_X1 U6066 ( .A(n4875), .ZN(n4874) );
  OAI21_X1 U6067 ( .B1(n8323), .B2(n4876), .A(n6254), .ZN(n4875) );
  INV_X1 U6068 ( .A(n9390), .ZN(n5748) );
  AND2_X1 U6069 ( .A1(n7307), .A2(n6587), .ZN(n4526) );
  AND2_X1 U6070 ( .A1(n4510), .A2(n8357), .ZN(n4527) );
  AND2_X1 U6071 ( .A1(n5214), .A2(n5213), .ZN(n4528) );
  AND2_X1 U6072 ( .A1(n6594), .A2(n6593), .ZN(n4529) );
  INV_X1 U6073 ( .A(n7182), .ZN(n4960) );
  NAND2_X2 U6074 ( .A1(n6709), .A2(n4511), .ZN(n5341) );
  NAND2_X1 U6075 ( .A1(n6221), .A2(n5838), .ZN(n6219) );
  NAND2_X1 U6076 ( .A1(n5157), .A2(n5156), .ZN(n5752) );
  INV_X1 U6077 ( .A(n5320), .ZN(n5171) );
  AND2_X1 U6078 ( .A1(n5081), .A2(n5078), .ZN(n4530) );
  INV_X1 U6079 ( .A(n6968), .ZN(n4962) );
  OR2_X1 U6080 ( .A1(n4510), .A2(n8357), .ZN(n4531) );
  AND2_X1 U6081 ( .A1(n6452), .A2(n6453), .ZN(n4532) );
  NOR2_X1 U6082 ( .A1(n8428), .A2(n5122), .ZN(n4533) );
  NOR2_X1 U6083 ( .A1(n9474), .A2(n4942), .ZN(n4534) );
  NAND2_X1 U6084 ( .A1(n4906), .A2(n4904), .ZN(n4903) );
  NOR2_X1 U6085 ( .A1(n6483), .A2(n6482), .ZN(n4535) );
  AND2_X1 U6086 ( .A1(n4936), .A2(n4531), .ZN(n4536) );
  INV_X1 U6087 ( .A(n7465), .ZN(n4697) );
  NOR2_X1 U6088 ( .A1(n8919), .A2(n8645), .ZN(n8323) );
  XNOR2_X1 U6089 ( .A(n8525), .B(n10053), .ZN(n8236) );
  INV_X1 U6090 ( .A(n8236), .ZN(n4665) );
  OR2_X1 U6091 ( .A1(n6629), .A2(n8704), .ZN(n4537) );
  NOR2_X1 U6092 ( .A1(n7331), .A2(n7330), .ZN(n4538) );
  NAND2_X1 U6093 ( .A1(n9040), .A2(n8068), .ZN(n9114) );
  AND2_X1 U6094 ( .A1(n5116), .A2(n8494), .ZN(n4539) );
  INV_X1 U6095 ( .A(n8263), .ZN(n4813) );
  NAND2_X1 U6096 ( .A1(n8526), .A2(n10047), .ZN(n4540) );
  AND2_X1 U6097 ( .A1(n6470), .A2(n6550), .ZN(n4541) );
  AND2_X1 U6098 ( .A1(n9623), .A2(n9199), .ZN(n4542) );
  XNOR2_X1 U6099 ( .A(n5789), .B(n5788), .ZN(n6198) );
  NOR3_X1 U6100 ( .A1(n5752), .A2(n4521), .A3(P1_IR_REG_29__SCAN_IN), .ZN(
        n5164) );
  INV_X1 U6101 ( .A(n6417), .ZN(n4914) );
  INV_X1 U6102 ( .A(n8340), .ZN(n4677) );
  AND2_X1 U6103 ( .A1(n9385), .A2(n4518), .ZN(n4543) );
  OR2_X1 U6104 ( .A1(n9974), .A2(n8535), .ZN(n4544) );
  OR2_X1 U6105 ( .A1(n6625), .A2(n8705), .ZN(n4545) );
  AND3_X1 U6106 ( .A1(n4540), .A2(n5926), .A3(n5950), .ZN(n4546) );
  AND2_X1 U6107 ( .A1(n5836), .A2(n5835), .ZN(n4547) );
  INV_X1 U6108 ( .A(n5038), .ZN(n5037) );
  NOR2_X1 U6109 ( .A1(n5476), .A2(n5041), .ZN(n5038) );
  NAND2_X1 U6110 ( .A1(n6333), .A2(n6332), .ZN(n9357) );
  INV_X1 U6111 ( .A(n8331), .ZN(n4766) );
  NAND2_X1 U6112 ( .A1(n5129), .A2(n5128), .ZN(n6094) );
  NOR2_X1 U6113 ( .A1(n9623), .A2(n9199), .ZN(n4548) );
  NOR2_X1 U6114 ( .A1(n6430), .A2(n6429), .ZN(n4549) );
  NAND2_X1 U6115 ( .A1(n5666), .A2(n5665), .ZN(n9418) );
  AND2_X1 U6116 ( .A1(n5509), .A2(n5508), .ZN(n9849) );
  INV_X1 U6117 ( .A(n9849), .ZN(n7740) );
  INV_X1 U6118 ( .A(n4925), .ZN(n4924) );
  XOR2_X1 U6119 ( .A(n7779), .B(n8128), .Z(n4550) );
  AND2_X1 U6120 ( .A1(n4754), .A2(n4751), .ZN(n4551) );
  AND2_X1 U6121 ( .A1(n8299), .A2(n8326), .ZN(n4552) );
  NOR2_X1 U6122 ( .A1(n9608), .A2(n9145), .ZN(n4553) );
  AND2_X1 U6123 ( .A1(n8913), .A2(n8636), .ZN(n4554) );
  AND2_X1 U6124 ( .A1(n5088), .A2(n5087), .ZN(n4555) );
  NAND2_X1 U6125 ( .A1(n9432), .A2(n4845), .ZN(n4846) );
  AND4_X1 U6126 ( .A1(n5175), .A2(n5174), .A3(n5173), .A4(n5172), .ZN(n9169)
         );
  NAND2_X1 U6127 ( .A1(n8126), .A2(n8125), .ZN(n4556) );
  INV_X1 U6128 ( .A(n8133), .ZN(n4753) );
  AND2_X1 U6129 ( .A1(n6602), .A2(n6601), .ZN(n4557) );
  INV_X1 U6130 ( .A(n4908), .ZN(n4907) );
  NAND2_X1 U6131 ( .A1(n6317), .A2(n6466), .ZN(n4908) );
  INV_X1 U6132 ( .A(n4928), .ZN(n4927) );
  NAND2_X1 U6133 ( .A1(n5503), .A2(n7740), .ZN(n4928) );
  AND2_X1 U6134 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n7750), .ZN(n4558) );
  OR2_X1 U6135 ( .A1(n6549), .A2(n9649), .ZN(n4559) );
  INV_X1 U6136 ( .A(n8259), .ZN(n8793) );
  NOR2_X1 U6137 ( .A1(n9704), .A2(n9207), .ZN(n4560) );
  INV_X1 U6138 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5837) );
  INV_X1 U6139 ( .A(n5079), .ZN(n5078) );
  NAND2_X1 U6140 ( .A1(n5080), .A2(n5082), .ZN(n5079) );
  AND2_X1 U6141 ( .A1(n9536), .A2(n9202), .ZN(n4561) );
  INV_X1 U6142 ( .A(n5041), .ZN(n5040) );
  NOR2_X1 U6143 ( .A1(n5224), .A2(SI_11_), .ZN(n5041) );
  AND2_X1 U6144 ( .A1(n8335), .A2(n8152), .ZN(n4562) );
  AND2_X1 U6145 ( .A1(n4754), .A2(n5075), .ZN(n4563) );
  AND4_X1 U6146 ( .A1(n5332), .A2(n5330), .A3(n5331), .A4(n5329), .ZN(n7087)
         );
  NAND2_X1 U6147 ( .A1(n5127), .A2(n5128), .ZN(n4564) );
  INV_X1 U6148 ( .A(n5084), .ZN(n5083) );
  OR2_X1 U6149 ( .A1(n8112), .A2(n5085), .ZN(n5084) );
  INV_X1 U6150 ( .A(n5861), .ZN(n4972) );
  INV_X1 U6151 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5838) );
  INV_X1 U6152 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5283) );
  OR3_X1 U6153 ( .A1(n6219), .A2(P2_IR_REG_22__SCAN_IN), .A3(n5131), .ZN(n4565) );
  OR2_X1 U6154 ( .A1(n6469), .A2(n4726), .ZN(n4566) );
  AND2_X1 U6155 ( .A1(n4510), .A2(n9192), .ZN(n6470) );
  INV_X1 U6156 ( .A(n6470), .ZN(n4904) );
  AND2_X1 U6157 ( .A1(n4774), .A2(n4770), .ZN(n4567) );
  INV_X1 U6158 ( .A(n4752), .ZN(n4750) );
  NAND2_X1 U6159 ( .A1(n5075), .A2(n4556), .ZN(n4752) );
  NOR2_X1 U6160 ( .A1(n5074), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n5073) );
  AND2_X1 U6161 ( .A1(n4771), .A2(n4770), .ZN(n4568) );
  OR2_X1 U6162 ( .A1(n7912), .A2(n7911), .ZN(n4569) );
  AND2_X1 U6163 ( .A1(n5156), .A2(n4859), .ZN(n4570) );
  NAND2_X1 U6164 ( .A1(n5580), .A2(n5579), .ZN(n9632) );
  AND2_X1 U6165 ( .A1(n8254), .A2(n8255), .ZN(n8176) );
  INV_X1 U6166 ( .A(n8176), .ZN(n4817) );
  NOR2_X1 U6167 ( .A1(n5951), .A2(n4867), .ZN(n4571) );
  AND2_X1 U6168 ( .A1(n4747), .A2(n5076), .ZN(n4572) );
  NOR2_X1 U6169 ( .A1(n5014), .A2(n5233), .ZN(n5013) );
  INV_X1 U6170 ( .A(n6364), .ZN(n4647) );
  NOR2_X1 U6171 ( .A1(n9115), .A2(n4741), .ZN(n4740) );
  AND2_X1 U6172 ( .A1(n4817), .A2(n5998), .ZN(n4573) );
  AND2_X1 U6173 ( .A1(n8265), .A2(n8266), .ZN(n4574) );
  AND2_X1 U6174 ( .A1(n5054), .A2(n9129), .ZN(n4575) );
  AND2_X1 U6175 ( .A1(n4540), .A2(n5926), .ZN(n4576) );
  INV_X1 U6176 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4971) );
  AND2_X1 U6177 ( .A1(n4720), .A2(n4722), .ZN(n4577) );
  OR2_X1 U6178 ( .A1(n4903), .A2(n4899), .ZN(n4578) );
  AND3_X1 U6179 ( .A1(n4975), .A2(n4977), .A3(n4593), .ZN(P2_U3201) );
  INV_X1 U6180 ( .A(n8524), .ZN(n4862) );
  OR2_X1 U6181 ( .A1(n5232), .A2(n5017), .ZN(n4580) );
  INV_X1 U6182 ( .A(n9385), .ZN(n4937) );
  INV_X1 U6183 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5836) );
  INV_X1 U6184 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4611) );
  AND2_X1 U6185 ( .A1(n5971), .A2(n5981), .ZN(n7912) );
  INV_X1 U6186 ( .A(n7912), .ZN(n4983) );
  INV_X1 U6187 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5835) );
  AND2_X1 U6188 ( .A1(n5392), .A2(n5150), .ZN(n5480) );
  OR2_X1 U6189 ( .A1(n6069), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n4581) );
  AND2_X1 U6190 ( .A1(n8418), .A2(n4533), .ZN(n4582) );
  AND2_X1 U6191 ( .A1(n6619), .A2(n6620), .ZN(n4583) );
  NOR2_X1 U6192 ( .A1(n9514), .A2(n9628), .ZN(n9491) );
  NAND2_X1 U6193 ( .A1(n9569), .A2(n4854), .ZN(n4857) );
  INV_X1 U6194 ( .A(n8357), .ZN(n9192) );
  AND4_X1 U6195 ( .A1(n5699), .A2(n5698), .A3(n5697), .A4(n5696), .ZN(n8357)
         );
  AND2_X1 U6196 ( .A1(n5535), .A2(SI_16_), .ZN(n4584) );
  NAND2_X1 U6197 ( .A1(n5746), .A2(n5745), .ZN(n4585) );
  NOR2_X1 U6198 ( .A1(n8467), .A2(n6607), .ZN(n4586) );
  AOI21_X1 U6199 ( .B1(n5030), .B2(n5253), .A(n5029), .ZN(n5028) );
  INV_X1 U6200 ( .A(n5157), .ZN(n5553) );
  NAND2_X1 U6201 ( .A1(n5564), .A2(n5563), .ZN(n9536) );
  INV_X1 U6202 ( .A(n9536), .ZN(n4855) );
  INV_X1 U6203 ( .A(n8011), .ZN(n4852) );
  AND4_X1 U6204 ( .A1(n5516), .A2(n5515), .A3(n5514), .A4(n5513), .ZN(n8025)
         );
  INV_X1 U6205 ( .A(n8025), .ZN(n4922) );
  NAND2_X1 U6206 ( .A1(n7259), .A2(n7258), .ZN(n7340) );
  NAND2_X1 U6207 ( .A1(n6277), .A2(n6732), .ZN(n6565) );
  INV_X1 U6208 ( .A(n9058), .ZN(n5053) );
  AND2_X1 U6209 ( .A1(n6610), .A2(n6609), .ZN(n4587) );
  NAND2_X1 U6210 ( .A1(n6240), .A2(n10044), .ZN(n7483) );
  INV_X1 U6211 ( .A(n4929), .ZN(n7528) );
  AND2_X1 U6212 ( .A1(n5792), .A2(n5791), .ZN(n4588) );
  NAND2_X1 U6213 ( .A1(n9715), .A2(n9717), .ZN(n7567) );
  INV_X1 U6214 ( .A(n7576), .ZN(n4851) );
  AND2_X1 U6215 ( .A1(n4841), .A2(n4840), .ZN(n4589) );
  AND2_X1 U6216 ( .A1(n6882), .A2(n6873), .ZN(n9724) );
  INV_X1 U6217 ( .A(n9724), .ZN(n9699) );
  INV_X1 U6218 ( .A(n5905), .ZN(n8147) );
  AND2_X1 U6219 ( .A1(n6577), .A2(n6574), .ZN(n7137) );
  AND2_X1 U6220 ( .A1(n8597), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n4590) );
  AND2_X1 U6221 ( .A1(n4982), .A2(n4978), .ZN(n4591) );
  INV_X1 U6222 ( .A(n4981), .ZN(n4980) );
  OR2_X1 U6223 ( .A1(n8588), .A2(n4590), .ZN(n4981) );
  AND3_X1 U6224 ( .A1(n5125), .A2(n5124), .A3(n5123), .ZN(n7072) );
  INV_X1 U6225 ( .A(n5166), .ZN(n9682) );
  INV_X1 U6226 ( .A(n6840), .ZN(n6844) );
  INV_X1 U6227 ( .A(n8161), .ZN(n8195) );
  NAND2_X1 U6228 ( .A1(n6219), .A2(n6223), .ZN(n8161) );
  AND2_X1 U6229 ( .A1(n4687), .A2(n6972), .ZN(n4592) );
  AND2_X1 U6230 ( .A1(n6662), .A2(n8336), .ZN(n8827) );
  NOR2_X1 U6231 ( .A1(n8799), .A2(n8336), .ZN(n4784) );
  NAND2_X1 U6232 ( .A1(n4694), .A2(n7475), .ZN(n7511) );
  AOI21_X1 U6233 ( .B1(n4697), .B2(n7475), .A(n7661), .ZN(n4695) );
  INV_X1 U6234 ( .A(n7475), .ZN(n4959) );
  XNOR2_X1 U6235 ( .A(n8535), .B(n9974), .ZN(n9984) );
  NOR2_X1 U6236 ( .A1(n7958), .A2(n7884), .ZN(n7957) );
  NAND2_X1 U6237 ( .A1(n9994), .A2(n8555), .ZN(n10013) );
  NAND3_X1 U6238 ( .A1(n8603), .A2(n4700), .A3(n4591), .ZN(n4593) );
  AOI21_X2 U6239 ( .B1(n5433), .B2(n5432), .A(n5217), .ZN(n5444) );
  OAI21_X2 U6240 ( .B1(n9502), .B2(n9501), .A(n6433), .ZN(n9488) );
  MUX2_X2 U6241 ( .A(n5783), .B(n9584), .S(n9858), .Z(n5786) );
  OAI21_X1 U6242 ( .B1(n4699), .B2(n10023), .A(n8583), .ZN(P2_U3200) );
  INV_X1 U6243 ( .A(n7406), .ZN(n6398) );
  AND2_X2 U6244 ( .A1(n5150), .A2(n5151), .ZN(n5058) );
  NAND2_X1 U6245 ( .A1(n4913), .A2(n4916), .ZN(n4911) );
  NAND2_X1 U6246 ( .A1(n5229), .A2(n5228), .ZN(n5506) );
  AOI21_X2 U6247 ( .B1(n5739), .B2(n9756), .A(n4585), .ZN(n5139) );
  AOI21_X2 U6248 ( .B1(n8373), .B2(n8372), .A(n4595), .ZN(n8508) );
  NAND2_X2 U6249 ( .A1(n8420), .A2(n8419), .ZN(n8418) );
  INV_X1 U6250 ( .A(n4903), .ZN(n4902) );
  NAND2_X1 U6251 ( .A1(n9542), .A2(n6364), .ZN(n4646) );
  INV_X1 U6252 ( .A(n4900), .ZN(n4895) );
  NAND2_X1 U6253 ( .A1(n4918), .A2(n4917), .ZN(n9563) );
  NAND2_X1 U6254 ( .A1(n5263), .A2(n5262), .ZN(n5653) );
  NAND2_X1 U6255 ( .A1(n4987), .A2(n5240), .ZN(n5572) );
  NAND2_X1 U6256 ( .A1(n4636), .A2(n4639), .ZN(n7683) );
  INV_X1 U6257 ( .A(n9441), .ZN(n5651) );
  NAND3_X1 U6258 ( .A1(n5321), .A2(n5324), .A3(n4597), .ZN(n9215) );
  NAND2_X1 U6259 ( .A1(n5009), .A2(n5010), .ZN(n5552) );
  NAND2_X1 U6260 ( .A1(n4995), .A2(n4993), .ZN(n5277) );
  NAND2_X1 U6261 ( .A1(n5239), .A2(n5238), .ZN(n4987) );
  INV_X1 U6262 ( .A(n5519), .ZN(n5016) );
  NAND2_X1 U6263 ( .A1(n7776), .A2(n5047), .ZN(n7795) );
  AND2_X1 U6264 ( .A1(n7166), .A2(n7258), .ZN(n4731) );
  OAI21_X1 U6265 ( .B1(n8627), .B2(n8831), .A(n8626), .ZN(n8848) );
  NAND2_X1 U6266 ( .A1(n8821), .A2(n8204), .ZN(n5881) );
  OAI21_X1 U6267 ( .B1(n4877), .B2(n8323), .A(n4874), .ZN(n8619) );
  INV_X1 U6268 ( .A(n7977), .ZN(n6118) );
  OAI21_X2 U6269 ( .B1(n8669), .B2(n6168), .A(n6167), .ZN(n8657) );
  NAND2_X1 U6270 ( .A1(n4868), .A2(n4571), .ZN(n4865) );
  NAND2_X1 U6271 ( .A1(n5999), .A2(n4573), .ZN(n7833) );
  NAND2_X2 U6272 ( .A1(n6118), .A2(n6117), .ZN(n7979) );
  XNOR2_X2 U6273 ( .A(n8207), .B(n4601), .ZN(n8204) );
  INV_X1 U6274 ( .A(n6578), .ZN(n4601) );
  NAND2_X1 U6275 ( .A1(n6248), .A2(n8300), .ZN(n8679) );
  INV_X1 U6276 ( .A(n4829), .ZN(n4828) );
  OAI21_X1 U6277 ( .B1(n5022), .B2(n8191), .A(n5019), .ZN(n5018) );
  NAND2_X1 U6278 ( .A1(n4604), .A2(n4602), .ZN(P1_U3550) );
  OR2_X1 U6279 ( .A1(n9584), .A2(n5819), .ZN(n4604) );
  OR2_X1 U6280 ( .A1(n5164), .A2(n5282), .ZN(n5161) );
  INV_X1 U6281 ( .A(n5073), .ZN(n5072) );
  INV_X1 U6282 ( .A(n4958), .ZN(n9753) );
  XNOR2_X1 U6283 ( .A(n6630), .B(n6631), .ZN(n8379) );
  NAND2_X1 U6284 ( .A1(n5839), .A2(n5133), .ZN(n5132) );
  NAND3_X1 U6285 ( .A1(n8603), .A2(n4976), .A3(n8539), .ZN(n4975) );
  XNOR2_X2 U6286 ( .A(n9328), .B(n9327), .ZN(n9340) );
  OAI211_X1 U6287 ( .C1(n5337), .C2(n4989), .A(n4609), .B(n5142), .ZN(n5198)
         );
  NAND2_X1 U6288 ( .A1(n5187), .A2(n4988), .ZN(n4609) );
  NAND2_X2 U6289 ( .A1(n5448), .A2(n5223), .ZN(n5463) );
  NAND2_X1 U6290 ( .A1(n8655), .A2(n8314), .ZN(n4808) );
  NOR2_X2 U6291 ( .A1(n8798), .A2(n8799), .ZN(n6242) );
  NAND2_X1 U6292 ( .A1(n5039), .A2(n5040), .ZN(n5477) );
  OAI21_X1 U6293 ( .B1(n5859), .B2(n6687), .A(n4992), .ZN(n5180) );
  NAND2_X1 U6294 ( .A1(n4769), .A2(n4768), .ZN(n5433) );
  NAND2_X1 U6295 ( .A1(n5177), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5178) );
  NAND2_X1 U6296 ( .A1(n4811), .A2(n4810), .ZN(n8780) );
  AOI21_X1 U6297 ( .B1(n8156), .B2(n8157), .A(n8161), .ZN(n5022) );
  OR2_X2 U6298 ( .A1(n9425), .A2(n9429), .ZN(n9427) );
  AND2_X1 U6299 ( .A1(n9588), .A2(n9587), .ZN(n4686) );
  OR2_X2 U6300 ( .A1(n9529), .A2(n9528), .ZN(n9531) );
  NAND2_X2 U6301 ( .A1(n7729), .A2(n7730), .ZN(n7728) );
  AND2_X1 U6302 ( .A1(n6407), .A2(n7431), .ZN(n7406) );
  NAND2_X2 U6303 ( .A1(n9396), .A2(n9400), .ZN(n9395) );
  NAND2_X1 U6304 ( .A1(n6505), .A2(n6353), .ZN(n4930) );
  NAND3_X1 U6305 ( .A1(n4617), .A2(n5315), .A3(n5146), .ZN(n5354) );
  NAND2_X1 U6306 ( .A1(n4617), .A2(n5315), .ZN(n5352) );
  NAND2_X1 U6307 ( .A1(n4620), .A2(n4619), .ZN(n4618) );
  NAND2_X1 U6308 ( .A1(n4621), .A2(n4574), .ZN(n4620) );
  NAND2_X1 U6309 ( .A1(n4622), .A2(n4782), .ZN(n4621) );
  NAND3_X1 U6310 ( .A1(n4624), .A2(n8803), .A3(n4623), .ZN(n4622) );
  NAND2_X1 U6311 ( .A1(n8258), .A2(n8336), .ZN(n4623) );
  NAND2_X1 U6312 ( .A1(n4785), .A2(n4784), .ZN(n4624) );
  OR2_X1 U6313 ( .A1(n4780), .A2(n4779), .ZN(n4628) );
  NAND2_X1 U6314 ( .A1(n4628), .A2(n8336), .ZN(n4632) );
  NAND3_X1 U6315 ( .A1(n7973), .A2(n9684), .A3(n9239), .ZN(n4634) );
  NAND2_X1 U6316 ( .A1(n5431), .A2(n4637), .ZN(n4636) );
  NAND2_X1 U6317 ( .A1(n4646), .A2(n4644), .ZN(n4957) );
  AND2_X2 U6318 ( .A1(n5058), .A2(n5392), .ZN(n5157) );
  INV_X1 U6319 ( .A(n4891), .ZN(n4659) );
  INV_X1 U6320 ( .A(n5126), .ZN(n4660) );
  INV_X1 U6321 ( .A(n4661), .ZN(n6221) );
  NAND2_X1 U6322 ( .A1(n4663), .A2(n4776), .ZN(n4662) );
  NAND2_X1 U6323 ( .A1(n4664), .A2(n8298), .ZN(n4663) );
  NAND2_X1 U6324 ( .A1(n8294), .A2(n4777), .ZN(n4664) );
  NAND2_X1 U6325 ( .A1(n8232), .A2(n8231), .ZN(n4672) );
  NAND2_X1 U6326 ( .A1(n4665), .A2(n8229), .ZN(n4667) );
  NAND2_X1 U6327 ( .A1(n8222), .A2(n4666), .ZN(n4670) );
  AOI21_X1 U6328 ( .B1(n4673), .B2(n4671), .A(n8249), .ZN(n8257) );
  NAND3_X1 U6329 ( .A1(n5018), .A2(n4675), .A3(n4674), .ZN(n8345) );
  NAND3_X1 U6330 ( .A1(n4676), .A2(n8343), .A3(n4678), .ZN(n4674) );
  NAND3_X1 U6331 ( .A1(n4762), .A2(n8343), .A3(n4760), .ZN(n4675) );
  OR2_X1 U6332 ( .A1(n8339), .A2(n8913), .ZN(n4678) );
  INV_X1 U6333 ( .A(n7048), .ZN(n8196) );
  NAND2_X1 U6334 ( .A1(n7135), .A2(n6575), .ZN(n7048) );
  NAND2_X1 U6335 ( .A1(n4685), .A2(n4682), .ZN(P1_U3549) );
  OAI22_X1 U6336 ( .A1(n5748), .A2(n9645), .B1(n9875), .B2(n4684), .ZN(n4683)
         );
  NAND2_X1 U6337 ( .A1(n9589), .A2(n4686), .ZN(n9650) );
  NAND3_X1 U6338 ( .A1(n4687), .A2(P2_REG2_REG_3__SCAN_IN), .A3(n6972), .ZN(
        n9923) );
  NAND2_X1 U6339 ( .A1(n4690), .A2(n4692), .ZN(n9887) );
  NAND2_X1 U6340 ( .A1(n4693), .A2(n5849), .ZN(n9886) );
  OAI211_X1 U6341 ( .C1(n7466), .C2(n4959), .A(n4698), .B(n4695), .ZN(n7512)
         );
  XNOR2_X2 U6342 ( .A(n5284), .B(n5283), .ZN(n7973) );
  NAND4_X1 U6343 ( .A1(n4707), .A2(n4706), .A3(n4705), .A4(n6457), .ZN(n6465)
         );
  NAND3_X1 U6344 ( .A1(n6447), .A2(n4532), .A3(n4708), .ZN(n4705) );
  NAND3_X1 U6345 ( .A1(n6445), .A2(n4709), .A3(n4532), .ZN(n4706) );
  AND2_X1 U6346 ( .A1(n4709), .A2(n6446), .ZN(n4708) );
  NOR2_X1 U6347 ( .A1(n6473), .A2(n4541), .ZN(n4725) );
  AOI21_X1 U6348 ( .B1(n9716), .B2(n4728), .A(n4550), .ZN(n4727) );
  NAND2_X1 U6349 ( .A1(n5045), .A2(n4727), .ZN(n5046) );
  NAND2_X1 U6350 ( .A1(n7567), .A2(n7578), .ZN(n7776) );
  NAND2_X1 U6351 ( .A1(n4538), .A2(n7258), .ZN(n4732) );
  NAND2_X1 U6352 ( .A1(n7342), .A2(n7344), .ZN(n7561) );
  NAND3_X1 U6353 ( .A1(n4734), .A2(n7161), .A3(n4733), .ZN(n7162) );
  NAND2_X1 U6354 ( .A1(n7156), .A2(n4735), .ZN(n4733) );
  NAND3_X1 U6355 ( .A1(n7156), .A2(n6922), .A3(n6923), .ZN(n4734) );
  INV_X1 U6356 ( .A(n6988), .ZN(n4735) );
  NAND2_X1 U6357 ( .A1(n6989), .A2(n6988), .ZN(n7157) );
  NAND3_X1 U6358 ( .A1(n9152), .A2(n4740), .A3(n9156), .ZN(n4736) );
  AND2_X2 U6359 ( .A1(n8353), .A2(n7152), .ZN(n6981) );
  NAND2_X1 U6360 ( .A1(n9104), .A2(n4572), .ZN(n4743) );
  NAND2_X1 U6361 ( .A1(n9104), .A2(n5076), .ZN(n4754) );
  OAI211_X1 U6362 ( .C1(n9104), .C2(n4745), .A(n4743), .B(n4744), .ZN(n8139)
         );
  NAND2_X1 U6363 ( .A1(n5068), .A2(n4517), .ZN(n4755) );
  NAND3_X1 U6364 ( .A1(n4756), .A2(n9088), .A3(n4755), .ZN(n9086) );
  NAND2_X1 U6365 ( .A1(n4758), .A2(n5158), .ZN(n5755) );
  INV_X1 U6366 ( .A(n5752), .ZN(n4758) );
  NAND2_X1 U6367 ( .A1(n4759), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5177) );
  INV_X2 U6368 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4759) );
  MUX2_X1 U6369 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n4514), .Z(n5188) );
  NAND2_X1 U6370 ( .A1(n5390), .A2(n4568), .ZN(n4769) );
  OAI21_X1 U6371 ( .B1(n5390), .B2(n4774), .A(n4771), .ZN(n5418) );
  NAND2_X1 U6372 ( .A1(n5390), .A2(n5207), .ZN(n5402) );
  AOI21_X2 U6373 ( .B1(n5401), .B2(n4773), .A(n4772), .ZN(n4771) );
  NAND3_X1 U6374 ( .A1(n8276), .A2(n8278), .A3(n8272), .ZN(n4781) );
  MUX2_X1 U6375 ( .A(n9019), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  MUX2_X1 U6376 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9019), .S(n6229), .Z(n6575) );
  AOI21_X2 U6377 ( .B1(n4796), .B2(n10017), .A(n4793), .ZN(n8603) );
  NAND2_X1 U6378 ( .A1(n7285), .A2(n8162), .ZN(n4800) );
  NAND2_X1 U6379 ( .A1(n4801), .A2(n8223), .ZN(n7285) );
  NAND2_X1 U6380 ( .A1(n7274), .A2(n8165), .ZN(n4801) );
  NAND2_X1 U6381 ( .A1(n4806), .A2(n4803), .ZN(n4802) );
  OAI21_X1 U6382 ( .B1(n6261), .B2(n8831), .A(n6260), .ZN(n4805) );
  NAND2_X1 U6383 ( .A1(n4808), .A2(n4807), .ZN(n6253) );
  INV_X1 U6384 ( .A(n7055), .ZN(n7052) );
  NAND2_X1 U6385 ( .A1(n4809), .A2(n8822), .ZN(n8817) );
  INV_X1 U6386 ( .A(n6578), .ZN(n10028) );
  NAND3_X1 U6387 ( .A1(n7484), .A2(n7483), .A3(n8231), .ZN(n6241) );
  NAND2_X1 U6388 ( .A1(n7838), .A2(n4812), .ZN(n4811) );
  AOI21_X1 U6389 ( .B1(n6242), .B2(n4817), .A(n4816), .ZN(n4815) );
  INV_X1 U6390 ( .A(n6242), .ZN(n4818) );
  NAND2_X1 U6391 ( .A1(n7837), .A2(n6242), .ZN(n8801) );
  NAND2_X1 U6392 ( .A1(n7838), .A2(n8176), .ZN(n7837) );
  NAND2_X1 U6393 ( .A1(n4821), .A2(n4819), .ZN(n6247) );
  NAND2_X1 U6394 ( .A1(n8712), .A2(n8289), .ZN(n4821) );
  INV_X1 U6395 ( .A(n8298), .ZN(n4822) );
  OR2_X1 U6396 ( .A1(n7655), .A2(n4829), .ZN(n4824) );
  NAND2_X2 U6397 ( .A1(n4508), .A2(n6226), .ZN(n5869) );
  MUX2_X1 U6398 ( .A(n4838), .B(n4837), .S(n6709), .Z(n7228) );
  NAND2_X2 U6399 ( .A1(n5286), .A2(n4658), .ZN(n9684) );
  NOR2_X1 U6400 ( .A1(n9352), .A2(n9353), .ZN(n9576) );
  XNOR2_X1 U6401 ( .A(n9360), .B(n9579), .ZN(n4839) );
  INV_X1 U6402 ( .A(n9800), .ZN(n4840) );
  INV_X1 U6403 ( .A(n4846), .ZN(n9386) );
  NOR2_X1 U6404 ( .A1(n7441), .A2(n4850), .ZN(n7684) );
  INV_X1 U6405 ( .A(n4857), .ZN(n9535) );
  NAND2_X1 U6406 ( .A1(n5157), .A2(n4570), .ZN(n4858) );
  NAND2_X1 U6407 ( .A1(n4858), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5285) );
  OR2_X1 U6408 ( .A1(n5950), .A2(n4862), .ZN(n4860) );
  NAND2_X1 U6409 ( .A1(n5927), .A2(n4576), .ZN(n4868) );
  NAND2_X1 U6410 ( .A1(n4864), .A2(n4863), .ZN(n5965) );
  NAND2_X1 U6411 ( .A1(n8644), .A2(n6187), .ZN(n4877) );
  NAND2_X1 U6412 ( .A1(n4869), .A2(n4872), .ZN(n6218) );
  NAND2_X1 U6413 ( .A1(n8644), .A2(n4870), .ZN(n4869) );
  OAI21_X2 U6414 ( .B1(n8773), .B2(n6057), .A(n6058), .ZN(n8765) );
  OAI22_X2 U6415 ( .A1(n8785), .A2(n6042), .B1(n8806), .B2(n8990), .ZN(n8773)
         );
  NAND2_X2 U6416 ( .A1(n6031), .A2(n6030), .ZN(n8785) );
  NAND2_X1 U6417 ( .A1(n7833), .A2(n6019), .ZN(n8804) );
  NAND2_X1 U6418 ( .A1(n4885), .A2(n4884), .ZN(n6157) );
  NAND2_X1 U6419 ( .A1(n4888), .A2(n4887), .ZN(n4886) );
  INV_X1 U6420 ( .A(n6690), .ZN(n4887) );
  INV_X1 U6421 ( .A(n6020), .ZN(n4888) );
  OR2_X1 U6422 ( .A1(n5905), .A2(n6691), .ZN(n4889) );
  AND3_X2 U6423 ( .A1(n4891), .A2(n4890), .A3(n5128), .ZN(n5845) );
  NAND2_X1 U6424 ( .A1(n4892), .A2(n5717), .ZN(n9763) );
  NAND3_X1 U6425 ( .A1(n6500), .A2(n6499), .A3(n4892), .ZN(n6501) );
  NAND2_X1 U6426 ( .A1(n9214), .A2(n9796), .ZN(n4892) );
  NAND2_X1 U6427 ( .A1(n9395), .A2(n4894), .ZN(n4893) );
  OAI211_X1 U6428 ( .C1(n9395), .C2(n4578), .A(n4896), .B(n4893), .ZN(n5805)
         );
  NAND2_X1 U6429 ( .A1(n9395), .A2(n4907), .ZN(n4905) );
  NAND2_X1 U6430 ( .A1(n9395), .A2(n6466), .ZN(n9381) );
  NAND2_X1 U6431 ( .A1(n7728), .A2(n4913), .ZN(n4912) );
  NAND2_X1 U6432 ( .A1(n7728), .A2(n6416), .ZN(n9558) );
  AOI21_X2 U6433 ( .B1(n9562), .B2(n4915), .A(n4914), .ZN(n4913) );
  INV_X1 U6434 ( .A(n9562), .ZN(n4916) );
  NAND2_X1 U6435 ( .A1(n7709), .A2(n4919), .ZN(n4918) );
  OAI21_X1 U6436 ( .B1(n7708), .B2(n4926), .A(n9849), .ZN(n4925) );
  INV_X1 U6437 ( .A(n5503), .ZN(n4926) );
  NAND2_X1 U6438 ( .A1(n7707), .A2(n5503), .ZN(n7727) );
  OR2_X1 U6439 ( .A1(n6405), .A2(n4931), .ZN(n6353) );
  NAND2_X2 U6440 ( .A1(n5719), .A2(n6500), .ZN(n7238) );
  OAI21_X1 U6441 ( .B1(n9401), .B2(n4935), .A(n4932), .ZN(n5796) );
  NAND2_X1 U6442 ( .A1(n4948), .A2(n4946), .ZN(n5431) );
  INV_X1 U6443 ( .A(n5136), .ZN(n4949) );
  NAND3_X1 U6444 ( .A1(n4953), .A2(n4951), .A3(n4952), .ZN(n5727) );
  NAND2_X1 U6445 ( .A1(n5726), .A2(n4955), .ZN(n4952) );
  NAND2_X1 U6446 ( .A1(n7529), .A2(n5726), .ZN(n4953) );
  NOR2_X1 U6447 ( .A1(n4954), .A2(n7708), .ZN(n4951) );
  NAND3_X1 U6448 ( .A1(n4953), .A2(n4952), .A3(n6510), .ZN(n7704) );
  NAND2_X1 U6449 ( .A1(n7690), .A2(n5724), .ZN(n7691) );
  INV_X1 U6450 ( .A(n6510), .ZN(n4954) );
  OAI21_X2 U6451 ( .B1(n7117), .B2(n5716), .A(n6497), .ZN(n4958) );
  OAI21_X2 U6452 ( .B1(n9520), .B2(n9519), .A(n6441), .ZN(n9502) );
  NAND2_X2 U6453 ( .A1(n9531), .A2(n6351), .ZN(n9520) );
  NAND2_X1 U6454 ( .A1(n8603), .A2(n10023), .ZN(n4977) );
  AND2_X1 U6455 ( .A1(n8588), .A2(n4590), .ZN(n4979) );
  INV_X1 U6456 ( .A(n5192), .ZN(n4989) );
  NAND2_X1 U6457 ( .A1(n5340), .A2(n5192), .ZN(n5358) );
  NAND2_X1 U6458 ( .A1(n5338), .A2(n5337), .ZN(n5340) );
  MUX2_X1 U6459 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(P1_DATAO_REG_0__SCAN_IN), 
        .S(n4513), .Z(n4990) );
  NAND2_X1 U6460 ( .A1(n5181), .A2(n4991), .ZN(n5297) );
  NAND2_X1 U6461 ( .A1(n5180), .A2(SI_1_), .ZN(n4991) );
  NAND2_X1 U6462 ( .A1(n5859), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4992) );
  NAND2_X1 U6463 ( .A1(n5268), .A2(n4996), .ZN(n4995) );
  NAND2_X1 U6464 ( .A1(n5268), .A2(n5267), .ZN(n5664) );
  NAND2_X1 U6465 ( .A1(n5688), .A2(n5687), .ZN(n5002) );
  NAND2_X1 U6466 ( .A1(n5519), .A2(n5013), .ZN(n5009) );
  INV_X1 U6467 ( .A(n5014), .ZN(n5012) );
  INV_X1 U6468 ( .A(SI_15_), .ZN(n5017) );
  NAND2_X1 U6469 ( .A1(n5250), .A2(n5249), .ZN(n5618) );
  NAND2_X1 U6470 ( .A1(n5023), .A2(n5025), .ZN(n5263) );
  NAND3_X1 U6471 ( .A1(n5250), .A2(n5028), .A3(n5249), .ZN(n5023) );
  OAI21_X1 U6472 ( .B1(n5463), .B2(n5034), .A(n5033), .ZN(n5229) );
  NAND2_X4 U6473 ( .A1(n6846), .A2(n5042), .ZN(n8353) );
  AND2_X2 U6474 ( .A1(n7220), .A2(n6875), .ZN(n5042) );
  NAND2_X1 U6475 ( .A1(n5044), .A2(n7775), .ZN(n5045) );
  NAND2_X1 U6476 ( .A1(n7795), .A2(n5046), .ZN(n9697) );
  INV_X1 U6477 ( .A(n7775), .ZN(n5049) );
  NAND2_X1 U6478 ( .A1(n9086), .A2(n8054), .ZN(n8060) );
  NAND2_X1 U6479 ( .A1(n8005), .A2(n5052), .ZN(n5051) );
  NAND2_X1 U6480 ( .A1(n5051), .A2(n4575), .ZN(n9134) );
  NAND3_X1 U6481 ( .A1(n5058), .A2(n5558), .A3(n5393), .ZN(n5560) );
  NAND2_X1 U6482 ( .A1(n9021), .A2(n8030), .ZN(n9179) );
  INV_X1 U6483 ( .A(n9177), .ZN(n5070) );
  OAI21_X2 U6484 ( .B1(n8443), .B2(n5103), .A(n5100), .ZN(n6630) );
  NAND2_X1 U6485 ( .A1(n8410), .A2(n4539), .ZN(n5114) );
  NAND2_X1 U6486 ( .A1(n8418), .A2(n5120), .ZN(n5118) );
  NAND2_X1 U6487 ( .A1(n5118), .A2(n5119), .ZN(n8385) );
  NAND2_X1 U6488 ( .A1(n8418), .A2(n6616), .ZN(n8427) );
  INV_X1 U6489 ( .A(n6616), .ZN(n5122) );
  NAND2_X2 U6490 ( .A1(n5869), .A2(n4511), .ZN(n5905) );
  AND2_X2 U6491 ( .A1(n7604), .A2(n6596), .ZN(n7631) );
  NAND2_X1 U6492 ( .A1(n7457), .A2(n4529), .ZN(n7604) );
  NAND2_X2 U6493 ( .A1(n6599), .A2(n7668), .ZN(n7671) );
  INV_X2 U6494 ( .A(n6069), .ZN(n5128) );
  NAND2_X1 U6495 ( .A1(n7298), .A2(n4526), .ZN(n7306) );
  NAND2_X1 U6496 ( .A1(n6584), .A2(n6583), .ZN(n7298) );
  NAND2_X1 U6497 ( .A1(n7306), .A2(n7454), .ZN(n6591) );
  NAND2_X1 U6498 ( .A1(n6548), .A2(n6547), .ZN(n6564) );
  NAND2_X1 U6499 ( .A1(n6475), .A2(n4899), .ZN(n6479) );
  XNOR2_X1 U6500 ( .A(n8621), .B(n8620), .ZN(n8627) );
  INV_X1 U6501 ( .A(n5319), .ZN(n5602) );
  INV_X1 U6502 ( .A(n8619), .ZN(n8621) );
  INV_X1 U6503 ( .A(n7162), .ZN(n7164) );
  OR2_X1 U6504 ( .A1(n5597), .A2(n5303), .ZN(n5307) );
  NAND2_X1 U6505 ( .A1(n5706), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5708) );
  OAI21_X2 U6506 ( .B1(n5706), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5705) );
  AOI21_X2 U6507 ( .B1(n8657), .B2(n8656), .A(n6179), .ZN(n8644) );
  NAND2_X1 U6508 ( .A1(n5139), .A2(n5750), .ZN(n5751) );
  NAND2_X2 U6509 ( .A1(n6637), .A2(n6636), .ZN(n8410) );
  NAND2_X1 U6510 ( .A1(n6245), .A2(n4515), .ZN(n6246) );
  NAND2_X1 U6511 ( .A1(n6572), .A2(n7072), .ZN(n8199) );
  CLKBUF_X1 U6512 ( .A(n6572), .Z(n8826) );
  XNOR2_X1 U6513 ( .A(n8150), .B(n8188), .ZN(n8610) );
  INV_X1 U6514 ( .A(n8140), .ZN(n5170) );
  AND2_X1 U6515 ( .A1(n6670), .A2(n6669), .ZN(n5134) );
  OR3_X1 U6516 ( .A1(n6472), .A2(n6492), .A3(n6468), .ZN(n5135) );
  INV_X1 U6517 ( .A(n10101), .ZN(n10098) );
  INV_X2 U6518 ( .A(n10086), .ZN(n10084) );
  NAND2_X1 U6519 ( .A1(n7214), .A2(n8819), .ZN(n8835) );
  INV_X1 U6520 ( .A(n8835), .ZN(n8812) );
  OR2_X1 U6521 ( .A1(n7566), .A2(n9209), .ZN(n5136) );
  AND2_X1 U6522 ( .A1(n6024), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5137) );
  INV_X1 U6523 ( .A(n8744), .ZN(n6620) );
  AND2_X2 U6524 ( .A1(n7003), .A2(n9565), .ZN(n9773) );
  NAND2_X1 U6525 ( .A1(n9858), .A2(n9801), .ZN(n9675) );
  AND2_X2 U6526 ( .A1(n5818), .A2(n5782), .ZN(n9858) );
  INV_X1 U6527 ( .A(n9858), .ZN(n5809) );
  AND2_X1 U6528 ( .A1(n8324), .A2(n6301), .ZN(n5138) );
  INV_X1 U6529 ( .A(n8913), .ZN(n6210) );
  NOR2_X1 U6530 ( .A1(n5581), .A2(n5565), .ZN(n5140) );
  OR2_X1 U6531 ( .A1(n8943), .A2(n8672), .ZN(n5141) );
  NOR2_X1 U6532 ( .A1(n5557), .A2(n5556), .ZN(n5558) );
  INV_X1 U6533 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8429) );
  AND2_X1 U6534 ( .A1(n5196), .A2(n5197), .ZN(n5142) );
  AND2_X1 U6535 ( .A1(n8610), .A2(n10076), .ZN(n5143) );
  AND2_X1 U6536 ( .A1(n4513), .A2(P2_U3151), .ZN(n9010) );
  INV_X1 U6537 ( .A(n8324), .ZN(n8847) );
  INV_X1 U6538 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5974) );
  OR2_X1 U6539 ( .A1(n9632), .A2(n9201), .ZN(n5144) );
  AND2_X1 U6540 ( .A1(n5438), .A2(n6799), .ZN(n5145) );
  INV_X1 U6541 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5831) );
  INV_X1 U6542 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5554) );
  INV_X1 U6543 ( .A(n8338), .ZN(n8154) );
  NAND2_X1 U6544 ( .A1(n8153), .A2(n4562), .ZN(n8155) );
  INV_X1 U6545 ( .A(n8636), .ZN(n6209) );
  INV_X1 U6546 ( .A(n9698), .ZN(n7783) );
  NOR2_X1 U6547 ( .A1(n8155), .A2(n8154), .ZN(n8156) );
  INV_X1 U6548 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5826) );
  INV_X1 U6549 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5363) );
  INV_X1 U6550 ( .A(n7607), .ZN(n6594) );
  INV_X1 U6551 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5912) );
  AND2_X1 U6552 ( .A1(n9093), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5581) );
  INV_X1 U6553 ( .A(n9623), .ZN(n5747) );
  INV_X1 U6554 ( .A(n6842), .ZN(n6551) );
  INV_X1 U6555 ( .A(SI_28_), .ZN(n5791) );
  INV_X1 U6556 ( .A(SI_26_), .ZN(n10239) );
  INV_X1 U6557 ( .A(SI_22_), .ZN(n10517) );
  INV_X1 U6558 ( .A(SI_19_), .ZN(n10253) );
  INV_X1 U6559 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5151) );
  INV_X1 U6560 ( .A(SI_7_), .ZN(n10449) );
  INV_X1 U6561 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5146) );
  INV_X1 U6562 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7518) );
  INV_X1 U6563 ( .A(n8806), .ZN(n6609) );
  INV_X1 U6564 ( .A(n4509), .ZN(n5911) );
  INV_X1 U6565 ( .A(n7917), .ZN(n7965) );
  NOR2_X1 U6566 ( .A1(n6171), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6182) );
  OR2_X1 U6567 ( .A1(n6111), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6122) );
  OR2_X1 U6568 ( .A1(n6051), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6075) );
  NOR2_X1 U6569 ( .A1(n5940), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5954) );
  INV_X1 U6570 ( .A(n8964), .ZN(n6301) );
  INV_X1 U6571 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5408) );
  INV_X1 U6572 ( .A(n7166), .ZN(n7163) );
  NAND2_X1 U6573 ( .A1(n9134), .A2(n8023), .ZN(n8029) );
  AND2_X1 U6574 ( .A1(n5643), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U6575 ( .A1(n5581), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5599) );
  AND2_X1 U6576 ( .A1(n5695), .A2(n5740), .ZN(n9375) );
  AND2_X1 U6577 ( .A1(n6551), .A2(n6844), .ZN(n6872) );
  INV_X1 U6578 ( .A(n9491), .ZN(n9506) );
  OR2_X1 U6579 ( .A1(n7440), .A2(n7566), .ZN(n7441) );
  NAND2_X1 U6580 ( .A1(n5225), .A2(SI_12_), .ZN(n5226) );
  NOR2_X1 U6581 ( .A1(n6075), .A2(n6074), .ZN(n6086) );
  OR2_X1 U6582 ( .A1(n6566), .A2(n6294), .ZN(n6655) );
  INV_X1 U6583 ( .A(n6226), .ZN(n6939) );
  OR2_X1 U6584 ( .A1(n6152), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6160) );
  INV_X1 U6585 ( .A(n8827), .ZN(n8755) );
  OR2_X1 U6586 ( .A1(n10057), .A2(n8524), .ZN(n8243) );
  NAND2_X1 U6587 ( .A1(n6664), .A2(n8336), .ZN(n8757) );
  OR2_X1 U6588 ( .A1(n6565), .A2(n7063), .ZN(n7064) );
  INV_X1 U6589 ( .A(n8645), .ZN(n8622) );
  NAND2_X1 U6590 ( .A1(n8953), .A2(n8691), .ZN(n8298) );
  AND2_X1 U6591 ( .A1(n6294), .A2(n6225), .ZN(n8831) );
  AND2_X1 U6592 ( .A1(n6644), .A2(n8820), .ZN(n6651) );
  INV_X1 U6593 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5842) );
  OR2_X1 U6594 ( .A1(n5526), .A2(n9184), .ZN(n5543) );
  AND2_X1 U6595 ( .A1(n5630), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5643) );
  INV_X1 U6596 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6799) );
  INV_X1 U6597 ( .A(n7557), .ZN(n6883) );
  INV_X1 U6598 ( .A(n6371), .ZN(n9400) );
  OR2_X1 U6599 ( .A1(n5469), .A2(n5468), .ZN(n5495) );
  OR2_X1 U6600 ( .A1(n6349), .A2(n9232), .ZN(n9168) );
  AND2_X1 U6601 ( .A1(n6872), .A2(n6555), .ZN(n6878) );
  INV_X1 U6602 ( .A(n9573), .ZN(n9709) );
  AND2_X1 U6604 ( .A1(n5267), .A2(n5266), .ZN(n5652) );
  OAI21_X1 U6605 ( .B1(n5227), .B2(SI_13_), .A(n5228), .ZN(n5490) );
  AND2_X1 U6606 ( .A1(n5207), .A2(n5206), .ZN(n5387) );
  INV_X1 U6607 ( .A(n8510), .ZN(n8480) );
  OR2_X1 U6608 ( .A1(n6661), .A2(n6655), .ZN(n6647) );
  OR2_X1 U6609 ( .A1(n4509), .A2(n8606), .ZN(n7101) );
  OR2_X1 U6610 ( .A1(n6679), .A2(n6678), .ZN(n6934) );
  INV_X1 U6611 ( .A(n9928), .ZN(n10017) );
  OR2_X1 U6612 ( .A1(n8823), .A2(n8833), .ZN(n7276) );
  OR2_X1 U6613 ( .A1(n10078), .A2(n6296), .ZN(n8820) );
  INV_X1 U6614 ( .A(n8882), .ZN(n8900) );
  OR2_X1 U6615 ( .A1(n7062), .A2(n6565), .ZN(n7070) );
  NAND2_X1 U6616 ( .A1(n7717), .A2(n8161), .ZN(n10078) );
  INV_X1 U6617 ( .A(n10078), .ZN(n10063) );
  AND2_X1 U6618 ( .A1(n7717), .A2(n6296), .ZN(n10076) );
  OR2_X1 U6619 ( .A1(n8823), .A2(n10076), .ZN(n10083) );
  INV_X1 U6620 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6267) );
  AND2_X1 U6621 ( .A1(n6059), .A2(n6048), .ZN(n9957) );
  INV_X1 U6622 ( .A(n9694), .ZN(n9719) );
  OR2_X1 U6623 ( .A1(n6885), .A2(n7004), .ZN(n6887) );
  AND4_X1 U6624 ( .A1(n5549), .A2(n5548), .A3(n5547), .A4(n5546), .ZN(n9092)
         );
  OR2_X1 U6625 ( .A1(n6752), .A2(n6748), .ZN(n9341) );
  OR2_X1 U6626 ( .A1(n6713), .A2(n6712), .ZN(n6752) );
  INV_X1 U6627 ( .A(n9341), .ZN(n9319) );
  INV_X1 U6628 ( .A(n9570), .ZN(n9769) );
  INV_X1 U6629 ( .A(n5713), .ZN(n7223) );
  INV_X1 U6630 ( .A(n9875), .ZN(n5819) );
  AND2_X1 U6631 ( .A1(n6842), .A2(n6840), .ZN(n6884) );
  INV_X1 U6632 ( .A(n9675), .ZN(n5784) );
  AND2_X1 U6633 ( .A1(n6884), .A2(n6555), .ZN(n9801) );
  NAND2_X1 U6634 ( .A1(n7688), .A2(n7681), .ZN(n9845) );
  NAND2_X1 U6635 ( .A1(n6876), .A2(n5781), .ZN(n9775) );
  AND2_X1 U6636 ( .A1(n5538), .A2(n5523), .ZN(n7860) );
  AND2_X1 U6637 ( .A1(n5453), .A2(n5464), .ZN(n7019) );
  NAND2_X1 U6638 ( .A1(n5373), .A2(n5372), .ZN(n5375) );
  INV_X1 U6639 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10118) );
  AND2_X1 U6640 ( .A1(n5964), .A2(n5963), .ZN(n10057) );
  AND2_X1 U6641 ( .A1(n6647), .A2(n6646), .ZN(n8503) );
  INV_X1 U6642 ( .A(n8501), .ZN(n8517) );
  NAND4_X1 U6643 ( .A1(n6208), .A2(n6207), .A3(n6206), .A4(n6205), .ZN(n8636)
         );
  INV_X1 U6644 ( .A(n8398), .ZN(n8705) );
  INV_X1 U6645 ( .A(n8403), .ZN(n8805) );
  OR2_X1 U6646 ( .A1(n6934), .A2(P2_U3151), .ZN(n8528) );
  INV_X1 U6647 ( .A(n10007), .ZN(n9941) );
  INV_X1 U6648 ( .A(n10016), .ZN(n9937) );
  NAND2_X1 U6649 ( .A1(n9881), .A2(n8346), .ZN(n10023) );
  INV_X1 U6650 ( .A(n8812), .ZN(n8810) );
  NAND2_X1 U6651 ( .A1(n8835), .A2(n7276), .ZN(n8816) );
  NAND2_X1 U6652 ( .A1(n10101), .A2(n10083), .ZN(n8903) );
  AND3_X2 U6653 ( .A1(n7205), .A2(n7071), .A3(n7070), .ZN(n10101) );
  OR2_X1 U6654 ( .A1(n10086), .A2(n10078), .ZN(n8964) );
  OR2_X1 U6655 ( .A1(n10086), .A2(n10058), .ZN(n8999) );
  AND2_X1 U6656 ( .A1(n10052), .A2(n10051), .ZN(n10092) );
  AND2_X1 U6657 ( .A1(n6300), .A2(n6299), .ZN(n10086) );
  AND2_X1 U6658 ( .A1(n6679), .A2(n7131), .ZN(n7067) );
  INV_X1 U6659 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7725) );
  INV_X1 U6660 ( .A(n9957), .ZN(n8568) );
  NAND2_X1 U6661 ( .A1(n9094), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9727) );
  OR2_X1 U6662 ( .A1(n6885), .A2(n6555), .ZN(n9694) );
  AND2_X1 U6663 ( .A1(n6887), .A2(n9565), .ZN(n9722) );
  OR2_X1 U6664 ( .A1(n5604), .A2(n5603), .ZN(n9200) );
  OR2_X1 U6665 ( .A1(n6752), .A2(n6751), .ZN(n9339) );
  OR2_X1 U6666 ( .A1(n9773), .A2(n7004), .ZN(n9761) );
  OR2_X1 U6667 ( .A1(n9773), .A2(n7084), .ZN(n9556) );
  NAND2_X1 U6668 ( .A1(n9875), .A2(n9801), .ZN(n9645) );
  AND2_X2 U6669 ( .A1(n5818), .A2(n5817), .ZN(n9875) );
  OR2_X1 U6670 ( .A1(n9775), .A2(n9774), .ZN(n9776) );
  INV_X1 U6671 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n10278) );
  INV_X1 U6672 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10447) );
  OR2_X1 U6673 ( .A1(n5482), .A2(n5157), .ZN(n7116) );
  INV_X1 U6674 ( .A(n7720), .ZN(n9686) );
  OAI21_X1 U6675 ( .B1(n8843), .B2(n10086), .A(n6304), .ZN(P2_U3456) );
  AND2_X2 U6676 ( .A1(n6876), .A2(n6677), .ZN(P1_U3973) );
  NAND2_X1 U6677 ( .A1(n6564), .A2(n6563), .ZN(P1_U3242) );
  INV_X1 U6678 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n5783) );
  NOR2_X2 U6679 ( .A1(n5354), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5392) );
  NOR2_X1 U6680 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5149) );
  NOR2_X1 U6681 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5153) );
  NOR2_X1 U6682 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5152) );
  NAND4_X1 U6683 ( .A1(n5701), .A2(n5153), .A3(n5152), .A4(n10519), .ZN(n5155)
         );
  NAND4_X1 U6684 ( .A1(n5707), .A2(n5704), .A3(n5776), .A4(n10235), .ZN(n5154)
         );
  NOR2_X2 U6685 ( .A1(n5155), .A2(n5154), .ZN(n5156) );
  NAND2_X1 U6686 ( .A1(n5162), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5163) );
  INV_X1 U6687 ( .A(n5164), .ZN(n9677) );
  NAND2_X2 U6688 ( .A1(n8140), .A2(n5166), .ZN(n5597) );
  INV_X4 U6689 ( .A(n5597), .ZN(n6334) );
  NAND2_X1 U6690 ( .A1(n6334), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5175) );
  AND2_X2 U6691 ( .A1(n8140), .A2(n9682), .ZN(n5319) );
  NAND2_X1 U6692 ( .A1(n5319), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5174) );
  NAND2_X1 U6693 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5364) );
  NOR2_X1 U6694 ( .A1(n5364), .A2(n5363), .ZN(n5380) );
  NAND2_X1 U6695 ( .A1(n5380), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5409) );
  NAND2_X1 U6696 ( .A1(n5456), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U6697 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n5167) );
  NAND2_X1 U6698 ( .A1(n5510), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5526) );
  INV_X1 U6699 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5542) );
  INV_X1 U6700 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5598) );
  INV_X1 U6701 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9120) );
  INV_X1 U6702 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9053) );
  NAND2_X1 U6703 ( .A1(n5656), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5668) );
  INV_X1 U6704 ( .A(n5668), .ZN(n5168) );
  NAND2_X1 U6705 ( .A1(n5168), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5682) );
  INV_X1 U6706 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9172) );
  NAND2_X1 U6707 ( .A1(n5681), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5693) );
  OAI21_X1 U6708 ( .B1(P1_REG3_REG_27__SCAN_IN), .B2(n5681), .A(n5693), .ZN(
        n5169) );
  INV_X1 U6709 ( .A(n5169), .ZN(n9389) );
  NAND2_X1 U6710 ( .A1(n4596), .A2(n9389), .ZN(n5173) );
  NAND2_X1 U6711 ( .A1(n5382), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5172) );
  MUX2_X1 U6712 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n4514), .Z(n5182) );
  NAND2_X1 U6713 ( .A1(n5182), .A2(SI_2_), .ZN(n5186) );
  INV_X1 U6714 ( .A(n5182), .ZN(n5184) );
  INV_X1 U6715 ( .A(SI_2_), .ZN(n5183) );
  NAND2_X1 U6716 ( .A1(n5184), .A2(n5183), .ZN(n5185) );
  AND2_X1 U6717 ( .A1(n5186), .A2(n5185), .ZN(n5314) );
  NAND2_X1 U6718 ( .A1(n5313), .A2(n5314), .ZN(n5187) );
  INV_X1 U6719 ( .A(n5188), .ZN(n5190) );
  INV_X1 U6720 ( .A(SI_3_), .ZN(n5189) );
  NAND2_X1 U6721 ( .A1(n5190), .A2(n5189), .ZN(n5191) );
  AND2_X1 U6722 ( .A1(n5192), .A2(n5191), .ZN(n5337) );
  NAND2_X1 U6723 ( .A1(n5193), .A2(SI_4_), .ZN(n5197) );
  INV_X1 U6724 ( .A(n5193), .ZN(n5195) );
  INV_X1 U6725 ( .A(SI_4_), .ZN(n5194) );
  NAND2_X1 U6726 ( .A1(n5195), .A2(n5194), .ZN(n5196) );
  NAND2_X1 U6727 ( .A1(n5198), .A2(n5197), .ZN(n5373) );
  MUX2_X1 U6728 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n4511), .Z(n5199) );
  NAND2_X1 U6729 ( .A1(n5199), .A2(SI_5_), .ZN(n5202) );
  INV_X1 U6730 ( .A(n5199), .ZN(n5200) );
  INV_X1 U6731 ( .A(SI_5_), .ZN(n10330) );
  NAND2_X1 U6732 ( .A1(n5200), .A2(n10330), .ZN(n5201) );
  AND2_X1 U6733 ( .A1(n5202), .A2(n5201), .ZN(n5372) );
  MUX2_X1 U6734 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n4511), .Z(n5203) );
  NAND2_X1 U6735 ( .A1(n5203), .A2(SI_6_), .ZN(n5207) );
  INV_X1 U6736 ( .A(n5203), .ZN(n5205) );
  INV_X1 U6737 ( .A(SI_6_), .ZN(n5204) );
  NAND2_X1 U6738 ( .A1(n5205), .A2(n5204), .ZN(n5206) );
  MUX2_X1 U6739 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4511), .Z(n5208) );
  NAND2_X1 U6740 ( .A1(n5208), .A2(SI_7_), .ZN(n5211) );
  INV_X1 U6741 ( .A(n5208), .ZN(n5209) );
  NAND2_X1 U6742 ( .A1(n5209), .A2(n10449), .ZN(n5210) );
  MUX2_X1 U6743 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n4511), .Z(n5212) );
  XNOR2_X1 U6744 ( .A(n5212), .B(SI_8_), .ZN(n5417) );
  INV_X1 U6745 ( .A(n5212), .ZN(n5214) );
  INV_X1 U6746 ( .A(SI_8_), .ZN(n5213) );
  MUX2_X1 U6747 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n4511), .Z(n5216) );
  XNOR2_X1 U6748 ( .A(n5216), .B(n5215), .ZN(n5432) );
  NOR2_X1 U6749 ( .A1(n5216), .A2(SI_9_), .ZN(n5217) );
  MUX2_X1 U6750 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n4511), .Z(n5218) );
  NAND2_X1 U6751 ( .A1(n5218), .A2(SI_10_), .ZN(n5223) );
  INV_X1 U6752 ( .A(n5218), .ZN(n5220) );
  INV_X1 U6753 ( .A(SI_10_), .ZN(n5219) );
  NAND2_X1 U6754 ( .A1(n5220), .A2(n5219), .ZN(n5221) );
  NAND2_X1 U6755 ( .A1(n5223), .A2(n5221), .ZN(n5445) );
  INV_X1 U6756 ( .A(n5445), .ZN(n5222) );
  MUX2_X1 U6757 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n4511), .Z(n5224) );
  XNOR2_X1 U6758 ( .A(n5224), .B(SI_11_), .ZN(n5462) );
  MUX2_X1 U6759 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n4511), .Z(n5225) );
  OAI21_X1 U6760 ( .B1(n5225), .B2(SI_12_), .A(n5226), .ZN(n5476) );
  MUX2_X1 U6761 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n4511), .Z(n5227) );
  MUX2_X1 U6762 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4511), .Z(n5504) );
  NAND2_X1 U6763 ( .A1(n5506), .A2(SI_14_), .ZN(n5230) );
  NAND2_X1 U6764 ( .A1(n5231), .A2(n5230), .ZN(n5519) );
  MUX2_X1 U6765 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n4511), .Z(n5517) );
  INV_X1 U6766 ( .A(n5517), .ZN(n5232) );
  MUX2_X1 U6767 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n4511), .Z(n5535) );
  NOR2_X1 U6768 ( .A1(n5535), .A2(SI_16_), .ZN(n5233) );
  INV_X1 U6769 ( .A(n5552), .ZN(n5239) );
  MUX2_X1 U6770 ( .A(n7236), .B(n10447), .S(n4511), .Z(n5235) );
  INV_X1 U6771 ( .A(SI_17_), .ZN(n5234) );
  NAND2_X1 U6772 ( .A1(n5235), .A2(n5234), .ZN(n5240) );
  INV_X1 U6773 ( .A(n5235), .ZN(n5236) );
  NAND2_X1 U6774 ( .A1(n5236), .A2(SI_17_), .ZN(n5237) );
  NAND2_X1 U6775 ( .A1(n5240), .A2(n5237), .ZN(n5551) );
  INV_X1 U6776 ( .A(n5551), .ZN(n5238) );
  MUX2_X1 U6777 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4511), .Z(n5242) );
  XNOR2_X1 U6778 ( .A(n5242), .B(n10460), .ZN(n5571) );
  INV_X1 U6779 ( .A(n5571), .ZN(n5241) );
  NAND2_X1 U6780 ( .A1(n5242), .A2(SI_18_), .ZN(n5243) );
  MUX2_X1 U6781 ( .A(n7420), .B(n7422), .S(n4511), .Z(n5244) );
  NAND2_X1 U6782 ( .A1(n5244), .A2(n10253), .ZN(n5247) );
  INV_X1 U6783 ( .A(n5244), .ZN(n5245) );
  NAND2_X1 U6784 ( .A1(n5245), .A2(SI_19_), .ZN(n5246) );
  NAND2_X1 U6785 ( .A1(n5247), .A2(n5246), .ZN(n5589) );
  MUX2_X1 U6786 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n4511), .Z(n5607) );
  INV_X1 U6787 ( .A(n5607), .ZN(n5248) );
  NAND2_X1 U6788 ( .A1(n5609), .A2(n10288), .ZN(n5249) );
  MUX2_X1 U6789 ( .A(n7598), .B(n7612), .S(n4511), .Z(n5616) );
  NOR2_X1 U6790 ( .A1(n5251), .A2(SI_21_), .ZN(n5253) );
  NAND2_X1 U6791 ( .A1(n5251), .A2(SI_21_), .ZN(n5252) );
  MUX2_X1 U6792 ( .A(n7718), .B(n10446), .S(n4511), .Z(n5254) );
  NAND2_X1 U6793 ( .A1(n5254), .A2(n10517), .ZN(n5257) );
  INV_X1 U6794 ( .A(n5254), .ZN(n5255) );
  NAND2_X1 U6795 ( .A1(n5255), .A2(SI_22_), .ZN(n5256) );
  NAND2_X1 U6796 ( .A1(n5257), .A2(n5256), .ZN(n5626) );
  MUX2_X1 U6797 ( .A(n7725), .B(n10278), .S(n4511), .Z(n5259) );
  INV_X1 U6798 ( .A(SI_23_), .ZN(n5258) );
  NAND2_X1 U6799 ( .A1(n5259), .A2(n5258), .ZN(n5262) );
  INV_X1 U6800 ( .A(n5259), .ZN(n5260) );
  NAND2_X1 U6801 ( .A1(n5260), .A2(SI_23_), .ZN(n5261) );
  INV_X1 U6802 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7808) );
  INV_X1 U6803 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7818) );
  MUX2_X1 U6804 ( .A(n7808), .B(n7818), .S(n4511), .Z(n5264) );
  INV_X1 U6805 ( .A(SI_24_), .ZN(n10506) );
  NAND2_X1 U6806 ( .A1(n5264), .A2(n10506), .ZN(n5267) );
  INV_X1 U6807 ( .A(n5264), .ZN(n5265) );
  NAND2_X1 U6808 ( .A1(n5265), .A2(SI_24_), .ZN(n5266) );
  NAND2_X1 U6809 ( .A1(n5653), .A2(n5652), .ZN(n5268) );
  INV_X1 U6810 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7880) );
  INV_X1 U6811 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10477) );
  MUX2_X1 U6812 ( .A(n7880), .B(n10477), .S(n4511), .Z(n5269) );
  INV_X1 U6813 ( .A(SI_25_), .ZN(n10291) );
  NAND2_X1 U6814 ( .A1(n5269), .A2(n10291), .ZN(n5272) );
  INV_X1 U6815 ( .A(n5269), .ZN(n5270) );
  NAND2_X1 U6816 ( .A1(n5270), .A2(SI_25_), .ZN(n5271) );
  INV_X1 U6817 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9016) );
  INV_X1 U6818 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10490) );
  MUX2_X1 U6819 ( .A(n9016), .B(n10490), .S(n4511), .Z(n5273) );
  NAND2_X1 U6820 ( .A1(n5273), .A2(n10239), .ZN(n5276) );
  INV_X1 U6821 ( .A(n5273), .ZN(n5274) );
  NAND2_X1 U6822 ( .A1(n5274), .A2(SI_26_), .ZN(n5275) );
  INV_X1 U6823 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7992) );
  INV_X1 U6824 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10317) );
  MUX2_X1 U6825 ( .A(n7992), .B(n10317), .S(n4511), .Z(n5279) );
  INV_X1 U6826 ( .A(SI_27_), .ZN(n5278) );
  NAND2_X1 U6827 ( .A1(n5279), .A2(n5278), .ZN(n5689) );
  INV_X1 U6828 ( .A(n5279), .ZN(n5280) );
  NAND2_X1 U6829 ( .A1(n5280), .A2(SI_27_), .ZN(n5281) );
  INV_X1 U6830 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5282) );
  NAND2_X1 U6831 ( .A1(n7991), .A2(n6347), .ZN(n5289) );
  OR2_X1 U6832 ( .A1(n5391), .A2(n10317), .ZN(n5288) );
  NAND2_X1 U6833 ( .A1(n5319), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5294) );
  NAND2_X1 U6834 ( .A1(n5327), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6835 ( .A1(n4512), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5292) );
  INV_X1 U6836 ( .A(n5597), .ZN(n5290) );
  NAND4_X1 U6837 ( .A1(n5294), .A2(n5293), .A3(n5292), .A4(n5291), .ZN(n6859)
         );
  INV_X1 U6838 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5295) );
  XNOR2_X1 U6839 ( .A(n5297), .B(n5296), .ZN(n6688) );
  OR2_X1 U6840 ( .A1(n5341), .A2(n6688), .ZN(n5301) );
  INV_X1 U6841 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5299) );
  NAND2_X1 U6842 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5298) );
  OR2_X1 U6843 ( .A1(n6709), .A2(n6756), .ZN(n5300) );
  INV_X1 U6844 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U6845 ( .A1(n5319), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U6846 ( .A1(n5320), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5305) );
  NAND2_X1 U6847 ( .A1(n5327), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5304) );
  INV_X1 U6848 ( .A(SI_0_), .ZN(n5308) );
  NOR2_X1 U6849 ( .A1(n4514), .A2(n5308), .ZN(n5310) );
  INV_X1 U6850 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5309) );
  XNOR2_X1 U6851 ( .A(n5310), .B(n5309), .ZN(n9691) );
  NAND2_X1 U6852 ( .A1(n9218), .A2(n7005), .ZN(n7219) );
  NAND2_X1 U6853 ( .A1(n5713), .A2(n7219), .ZN(n5312) );
  INV_X1 U6854 ( .A(n6859), .ZN(n6494) );
  NAND2_X1 U6855 ( .A1(n6494), .A2(n9783), .ZN(n5311) );
  NAND2_X1 U6856 ( .A1(n5312), .A2(n5311), .ZN(n7120) );
  XNOR2_X1 U6857 ( .A(n5313), .B(n5314), .ZN(n6690) );
  OR2_X1 U6858 ( .A1(n5341), .A2(n6690), .ZN(n5318) );
  INV_X1 U6859 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5316) );
  INV_X1 U6860 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U6861 ( .A1(n5290), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5324) );
  NAND2_X1 U6862 ( .A1(n5319), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U6863 ( .A1(n5320), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U6864 ( .A1(n5327), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5321) );
  NAND2_X1 U6865 ( .A1(n5715), .A2(n6497), .ZN(n7121) );
  NAND2_X1 U6866 ( .A1(n7120), .A2(n7121), .ZN(n5326) );
  NAND2_X1 U6867 ( .A1(n6990), .A2(n9789), .ZN(n5325) );
  NAND2_X1 U6868 ( .A1(n5326), .A2(n5325), .ZN(n9764) );
  INV_X1 U6869 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9758) );
  NAND2_X1 U6870 ( .A1(n5327), .A2(n9758), .ZN(n5332) );
  NAND2_X1 U6871 ( .A1(n6334), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5331) );
  NAND2_X1 U6872 ( .A1(n5320), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5330) );
  INV_X1 U6873 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5328) );
  NAND2_X1 U6874 ( .A1(n5334), .A2(n5333), .ZN(n5335) );
  NAND2_X1 U6875 ( .A1(n5335), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5336) );
  INV_X1 U6876 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n10482) );
  XNOR2_X1 U6877 ( .A(n5336), .B(n10482), .ZN(n9251) );
  INV_X1 U6878 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6684) );
  OR2_X1 U6879 ( .A1(n5391), .A2(n6684), .ZN(n5343) );
  OR2_X1 U6880 ( .A1(n5338), .A2(n5337), .ZN(n5339) );
  NAND2_X1 U6881 ( .A1(n5340), .A2(n5339), .ZN(n6686) );
  OR2_X1 U6882 ( .A1(n5341), .A2(n6686), .ZN(n5342) );
  OAI211_X1 U6883 ( .C1(n6709), .C2(n9251), .A(n5343), .B(n5342), .ZN(n6991)
         );
  NAND2_X1 U6884 ( .A1(n7087), .A2(n6991), .ZN(n5717) );
  INV_X1 U6885 ( .A(n7087), .ZN(n9214) );
  NAND2_X1 U6886 ( .A1(n9764), .A2(n9763), .ZN(n5345) );
  NAND2_X1 U6887 ( .A1(n7087), .A2(n9796), .ZN(n5344) );
  NAND2_X1 U6888 ( .A1(n5345), .A2(n5344), .ZN(n7083) );
  INV_X2 U6889 ( .A(n5602), .ZN(n5798) );
  NAND2_X1 U6890 ( .A1(n5798), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5351) );
  NAND2_X1 U6891 ( .A1(n6334), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5350) );
  INV_X1 U6892 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U6893 ( .A1(n9758), .A2(n5346), .ZN(n5347) );
  AND2_X1 U6894 ( .A1(n5347), .A2(n5364), .ZN(n7167) );
  NAND2_X1 U6895 ( .A1(n4596), .A2(n7167), .ZN(n5349) );
  NAND2_X1 U6896 ( .A1(n5382), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U6897 ( .A1(n5352), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5353) );
  MUX2_X1 U6898 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5353), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5356) );
  NAND2_X1 U6899 ( .A1(n5356), .A2(n5355), .ZN(n9270) );
  INV_X1 U6900 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5357) );
  OR2_X1 U6901 ( .A1(n5391), .A2(n5357), .ZN(n5360) );
  XNOR2_X1 U6902 ( .A(n5358), .B(n5142), .ZN(n6689) );
  OR2_X1 U6903 ( .A1(n5341), .A2(n6689), .ZN(n5359) );
  OAI211_X1 U6904 ( .C1(n6709), .C2(n9270), .A(n5360), .B(n5359), .ZN(n9800)
         );
  NAND2_X1 U6905 ( .A1(n7263), .A2(n9800), .ZN(n6392) );
  INV_X1 U6906 ( .A(n7263), .ZN(n9213) );
  NAND2_X1 U6907 ( .A1(n9213), .A2(n4840), .ZN(n6496) );
  NAND2_X1 U6908 ( .A1(n6392), .A2(n6496), .ZN(n6354) );
  NAND2_X1 U6909 ( .A1(n7083), .A2(n6354), .ZN(n5362) );
  NAND2_X1 U6910 ( .A1(n7263), .A2(n4840), .ZN(n5361) );
  NAND2_X1 U6911 ( .A1(n5362), .A2(n5361), .ZN(n9747) );
  NAND2_X1 U6912 ( .A1(n5798), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5369) );
  NAND2_X1 U6913 ( .A1(n6334), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5368) );
  AND2_X1 U6914 ( .A1(n5364), .A2(n5363), .ZN(n5365) );
  NOR2_X1 U6915 ( .A1(n5380), .A2(n5365), .ZN(n9743) );
  NAND2_X1 U6916 ( .A1(n4596), .A2(n9743), .ZN(n5367) );
  NAND2_X1 U6917 ( .A1(n5382), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5366) );
  NAND2_X1 U6918 ( .A1(n5355), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5371) );
  INV_X1 U6919 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5370) );
  XNOR2_X1 U6920 ( .A(n5371), .B(n5370), .ZN(n6774) );
  OR2_X1 U6921 ( .A1(n5373), .A2(n5372), .ZN(n5374) );
  NAND2_X1 U6922 ( .A1(n5375), .A2(n5374), .ZN(n6693) );
  OR2_X1 U6923 ( .A1(n5341), .A2(n6693), .ZN(n5377) );
  INV_X1 U6924 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6694) );
  OR2_X1 U6925 ( .A1(n5391), .A2(n6694), .ZN(n5376) );
  OAI211_X1 U6926 ( .C1(n6709), .C2(n6774), .A(n5377), .B(n5376), .ZN(n7253)
         );
  NAND2_X1 U6927 ( .A1(n7260), .A2(n7253), .ZN(n6394) );
  INV_X1 U6928 ( .A(n7260), .ZN(n9212) );
  NAND2_X1 U6929 ( .A1(n9212), .A2(n9809), .ZN(n6500) );
  NAND2_X1 U6930 ( .A1(n6394), .A2(n6500), .ZN(n9746) );
  NAND2_X1 U6931 ( .A1(n9747), .A2(n9746), .ZN(n5379) );
  NAND2_X1 U6932 ( .A1(n7260), .A2(n9809), .ZN(n5378) );
  NAND2_X1 U6933 ( .A1(n5379), .A2(n5378), .ZN(n7245) );
  NAND2_X1 U6934 ( .A1(n6334), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5386) );
  NAND2_X1 U6935 ( .A1(n5798), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5385) );
  OR2_X1 U6936 ( .A1(n5380), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5381) );
  AND2_X1 U6937 ( .A1(n5409), .A2(n5381), .ZN(n7376) );
  NAND2_X1 U6938 ( .A1(n4596), .A2(n7376), .ZN(n5384) );
  NAND2_X1 U6939 ( .A1(n5382), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5383) );
  OR2_X1 U6940 ( .A1(n5388), .A2(n5387), .ZN(n5389) );
  NAND2_X1 U6941 ( .A1(n5390), .A2(n5389), .ZN(n6696) );
  OR2_X1 U6942 ( .A1(n6696), .A2(n5341), .ZN(n5398) );
  BUF_X1 U6943 ( .A(n5392), .Z(n5393) );
  NOR2_X1 U6944 ( .A1(n5393), .A2(n5282), .ZN(n5394) );
  NAND2_X1 U6945 ( .A1(n5394), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5396) );
  INV_X1 U6946 ( .A(n5394), .ZN(n5395) );
  INV_X1 U6947 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n10306) );
  NAND2_X1 U6948 ( .A1(n5395), .A2(n10306), .ZN(n5404) );
  AOI22_X1 U6949 ( .A1(n5594), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5593), .B2(
        n6792), .ZN(n5397) );
  NAND2_X1 U6950 ( .A1(n5398), .A2(n5397), .ZN(n7381) );
  NAND2_X1 U6951 ( .A1(n7345), .A2(n7381), .ZN(n6396) );
  INV_X1 U6952 ( .A(n7345), .ZN(n9211) );
  INV_X1 U6953 ( .A(n7381), .ZN(n9817) );
  NAND2_X1 U6954 ( .A1(n9211), .A2(n9817), .ZN(n7385) );
  NAND2_X1 U6955 ( .A1(n6396), .A2(n7385), .ZN(n7244) );
  NAND2_X1 U6956 ( .A1(n7245), .A2(n7244), .ZN(n5400) );
  NAND2_X1 U6957 ( .A1(n7345), .A2(n9817), .ZN(n5399) );
  NAND2_X1 U6958 ( .A1(n5400), .A2(n5399), .ZN(n7384) );
  OR2_X1 U6959 ( .A1(n6699), .A2(n5341), .ZN(n5407) );
  NAND2_X1 U6960 ( .A1(n5404), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5405) );
  XNOR2_X1 U6961 ( .A(n5405), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6793) );
  AOI22_X1 U6962 ( .A1(n5594), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5593), .B2(
        n6793), .ZN(n5406) );
  AND2_X2 U6963 ( .A1(n5407), .A2(n5406), .ZN(n9823) );
  NAND2_X1 U6964 ( .A1(n6334), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5414) );
  NAND2_X1 U6965 ( .A1(n5798), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5413) );
  NAND2_X1 U6966 ( .A1(n5409), .A2(n5408), .ZN(n5410) );
  AND2_X1 U6967 ( .A1(n5424), .A2(n5410), .ZN(n7396) );
  NAND2_X1 U6968 ( .A1(n4596), .A2(n7396), .ZN(n5412) );
  NAND2_X1 U6969 ( .A1(n5382), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5411) );
  NAND4_X1 U6970 ( .A1(n5414), .A2(n5413), .A3(n5412), .A4(n5411), .ZN(n9210)
         );
  NAND2_X1 U6971 ( .A1(n9823), .A2(n9210), .ZN(n6402) );
  INV_X1 U6972 ( .A(n9210), .ZN(n5415) );
  INV_X1 U6973 ( .A(n9823), .ZN(n7397) );
  NAND2_X1 U6974 ( .A1(n5415), .A2(n7397), .ZN(n7431) );
  NAND2_X1 U6975 ( .A1(n6402), .A2(n7431), .ZN(n7387) );
  NAND2_X1 U6976 ( .A1(n9823), .A2(n5415), .ZN(n5416) );
  XNOR2_X1 U6977 ( .A(n5418), .B(n5417), .ZN(n6705) );
  NAND2_X1 U6978 ( .A1(n6705), .A2(n6347), .ZN(n5422) );
  NOR2_X1 U6979 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5419) );
  NAND2_X1 U6980 ( .A1(n5393), .A2(n5419), .ZN(n5434) );
  NAND2_X1 U6981 ( .A1(n5434), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5420) );
  XNOR2_X1 U6982 ( .A(n5420), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6795) );
  AOI22_X1 U6983 ( .A1(n5594), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5593), .B2(
        n6795), .ZN(n5421) );
  NAND2_X1 U6984 ( .A1(n5422), .A2(n5421), .ZN(n7566) );
  NAND2_X1 U6985 ( .A1(n6334), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U6986 ( .A1(n5798), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5429) );
  NAND2_X1 U6987 ( .A1(n5382), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U6988 ( .A1(n5424), .A2(n5423), .ZN(n5425) );
  NAND2_X1 U6989 ( .A1(n5438), .A2(n5425), .ZN(n9728) );
  INV_X1 U6990 ( .A(n9728), .ZN(n5426) );
  NAND2_X1 U6991 ( .A1(n4596), .A2(n5426), .ZN(n5427) );
  NAND4_X1 U6992 ( .A1(n5430), .A2(n5429), .A3(n5428), .A4(n5427), .ZN(n9209)
         );
  NAND2_X1 U6993 ( .A1(n7566), .A2(n9209), .ZN(n7429) );
  XNOR2_X1 U6994 ( .A(n5433), .B(n5432), .ZN(n6720) );
  NAND2_X1 U6995 ( .A1(n6720), .A2(n6347), .ZN(n5437) );
  NAND2_X1 U6996 ( .A1(n5449), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5435) );
  XNOR2_X1 U6997 ( .A(n5435), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6892) );
  AOI22_X1 U6998 ( .A1(n5594), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5593), .B2(
        n6892), .ZN(n5436) );
  NAND2_X1 U6999 ( .A1(n5437), .A2(n5436), .ZN(n7576) );
  NAND2_X1 U7000 ( .A1(n6334), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5442) );
  NAND2_X1 U7001 ( .A1(n5798), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5441) );
  NOR2_X1 U7002 ( .A1(n5456), .A2(n5145), .ZN(n7585) );
  NAND2_X1 U7003 ( .A1(n4596), .A2(n7585), .ZN(n5440) );
  NAND2_X1 U7004 ( .A1(n5382), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5439) );
  OR2_X1 U7005 ( .A1(n7576), .A2(n7574), .ZN(n6409) );
  NAND2_X1 U7006 ( .A1(n7576), .A2(n7574), .ZN(n6421) );
  INV_X1 U7007 ( .A(n7574), .ZN(n9208) );
  OR2_X1 U7008 ( .A1(n7576), .A2(n9208), .ZN(n5443) );
  INV_X1 U7009 ( .A(n5444), .ZN(n5446) );
  NAND2_X1 U7010 ( .A1(n5446), .A2(n5445), .ZN(n5447) );
  NAND2_X1 U7011 ( .A1(n5448), .A2(n5447), .ZN(n6725) );
  OR2_X1 U7012 ( .A1(n6725), .A2(n5341), .ZN(n5455) );
  NAND2_X1 U7013 ( .A1(n5450), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5452) );
  INV_X1 U7014 ( .A(n5452), .ZN(n5451) );
  NAND2_X1 U7015 ( .A1(n5451), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5453) );
  INV_X1 U7016 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n10493) );
  NAND2_X1 U7017 ( .A1(n5452), .A2(n10493), .ZN(n5464) );
  AOI22_X1 U7018 ( .A1(n5594), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5593), .B2(
        n7019), .ZN(n5454) );
  NAND2_X1 U7019 ( .A1(n6334), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U7020 ( .A1(n5382), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U7021 ( .A1(n5798), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5459) );
  OR2_X1 U7022 ( .A1(n5456), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U7023 ( .A1(n5469), .A2(n5457), .ZN(n9706) );
  INV_X1 U7024 ( .A(n9706), .ZN(n7536) );
  NAND2_X1 U7025 ( .A1(n4596), .A2(n7536), .ZN(n5458) );
  OR2_X1 U7026 ( .A1(n9704), .A2(n7780), .ZN(n6508) );
  NAND2_X1 U7027 ( .A1(n9704), .A2(n7780), .ZN(n7689) );
  NAND2_X1 U7028 ( .A1(n6508), .A2(n7689), .ZN(n7530) );
  INV_X1 U7029 ( .A(n7780), .ZN(n9207) );
  XNOR2_X1 U7030 ( .A(n5463), .B(n5462), .ZN(n6736) );
  NAND2_X1 U7031 ( .A1(n6736), .A2(n6347), .ZN(n5467) );
  NAND2_X1 U7032 ( .A1(n5464), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5465) );
  XNOR2_X1 U7033 ( .A(n5465), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7109) );
  AOI22_X1 U7034 ( .A1(n5594), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5593), .B2(
        n7109), .ZN(n5466) );
  NAND2_X1 U7035 ( .A1(n5469), .A2(n5468), .ZN(n5470) );
  AND2_X1 U7036 ( .A1(n5495), .A2(n5470), .ZN(n9729) );
  NAND2_X1 U7037 ( .A1(n4596), .A2(n9729), .ZN(n5474) );
  NAND2_X1 U7038 ( .A1(n6334), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U7039 ( .A1(n5382), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U7040 ( .A1(n5798), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5471) );
  NAND2_X1 U7041 ( .A1(n9732), .A2(n7789), .ZN(n6423) );
  NAND2_X1 U7042 ( .A1(n7617), .A2(n6423), .ZN(n7694) );
  NAND2_X1 U7043 ( .A1(n7683), .A2(n7694), .ZN(n7682) );
  INV_X1 U7044 ( .A(n7789), .ZN(n9206) );
  OR2_X1 U7045 ( .A1(n9732), .A2(n9206), .ZN(n5475) );
  NAND2_X1 U7046 ( .A1(n7682), .A2(n5475), .ZN(n7615) );
  NAND2_X1 U7047 ( .A1(n5477), .A2(n5476), .ZN(n5479) );
  NAND2_X1 U7048 ( .A1(n5479), .A2(n5478), .ZN(n6741) );
  NOR2_X1 U7049 ( .A1(n5480), .A2(n5282), .ZN(n5481) );
  MUX2_X1 U7050 ( .A(n5282), .B(n5481), .S(P1_IR_REG_12__SCAN_IN), .Z(n5482)
         );
  INV_X1 U7051 ( .A(n7116), .ZN(n7361) );
  AOI22_X1 U7052 ( .A1(n5594), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5593), .B2(
        n7361), .ZN(n5483) );
  NAND2_X1 U7053 ( .A1(n6334), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U7054 ( .A1(n5382), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5487) );
  XNOR2_X1 U7055 ( .A(n5495), .B(P1_REG3_REG_12__SCAN_IN), .ZN(n9066) );
  NAND2_X1 U7056 ( .A1(n4596), .A2(n9066), .ZN(n5486) );
  NAND2_X1 U7057 ( .A1(n5798), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5485) );
  OR2_X1 U7058 ( .A1(n8011), .A2(n8009), .ZN(n6425) );
  NAND2_X1 U7059 ( .A1(n8011), .A2(n8009), .ZN(n6510) );
  NAND2_X1 U7060 ( .A1(n7615), .A2(n7618), .ZN(n7614) );
  INV_X1 U7061 ( .A(n8009), .ZN(n9205) );
  OR2_X1 U7062 ( .A1(n8011), .A2(n9205), .ZN(n5489) );
  NAND2_X1 U7063 ( .A1(n7614), .A2(n5489), .ZN(n7709) );
  XNOR2_X1 U7064 ( .A(n5491), .B(n5490), .ZN(n6834) );
  NAND2_X1 U7065 ( .A1(n6834), .A2(n6347), .ZN(n5494) );
  NAND2_X1 U7066 ( .A1(n5553), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5492) );
  XNOR2_X1 U7067 ( .A(n5492), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7547) );
  AOI22_X1 U7068 ( .A1(n5594), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5593), .B2(
        n7547), .ZN(n5493) );
  NAND2_X1 U7069 ( .A1(n6334), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5502) );
  NAND2_X1 U7070 ( .A1(n5382), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5501) );
  INV_X1 U7071 ( .A(n5495), .ZN(n5496) );
  AOI21_X1 U7072 ( .B1(n5496), .B2(P1_REG3_REG_12__SCAN_IN), .A(
        P1_REG3_REG_13__SCAN_IN), .ZN(n5497) );
  OR2_X1 U7073 ( .A1(n5497), .A2(n5510), .ZN(n9128) );
  INV_X1 U7074 ( .A(n9128), .ZN(n5498) );
  NAND2_X1 U7075 ( .A1(n4596), .A2(n5498), .ZN(n5500) );
  NAND2_X1 U7076 ( .A1(n5798), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5499) );
  NAND2_X1 U7077 ( .A1(n9137), .A2(n8018), .ZN(n6511) );
  NAND2_X1 U7078 ( .A1(n6514), .A2(n6511), .ZN(n7708) );
  INV_X1 U7079 ( .A(n8018), .ZN(n6729) );
  OR2_X1 U7080 ( .A1(n9137), .A2(n6729), .ZN(n5503) );
  XNOR2_X1 U7081 ( .A(n5504), .B(SI_14_), .ZN(n5505) );
  XNOR2_X1 U7082 ( .A(n5506), .B(n5505), .ZN(n6928) );
  NAND2_X1 U7083 ( .A1(n6928), .A2(n6347), .ZN(n5509) );
  OR2_X1 U7084 ( .A1(n5553), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U7085 ( .A1(n5507), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5520) );
  XNOR2_X1 U7086 ( .A(n5520), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7867) );
  AOI22_X1 U7087 ( .A1(n5594), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5593), .B2(
        n7867), .ZN(n5508) );
  NAND2_X1 U7088 ( .A1(n6334), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U7089 ( .A1(n5798), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5515) );
  OR2_X1 U7090 ( .A1(n5510), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5511) );
  AND2_X1 U7091 ( .A1(n5526), .A2(n5511), .ZN(n9028) );
  NAND2_X1 U7092 ( .A1(n4596), .A2(n9028), .ZN(n5514) );
  INV_X1 U7093 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n5512) );
  OR2_X1 U7094 ( .A1(n5171), .A2(n5512), .ZN(n5513) );
  XNOR2_X1 U7095 ( .A(n5517), .B(SI_15_), .ZN(n5518) );
  XNOR2_X1 U7096 ( .A(n5519), .B(n5518), .ZN(n6995) );
  NAND2_X1 U7097 ( .A1(n6995), .A2(n6347), .ZN(n5525) );
  NAND2_X1 U7098 ( .A1(n5520), .A2(n5555), .ZN(n5521) );
  NAND2_X1 U7099 ( .A1(n5521), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U7100 ( .A1(n5522), .A2(n10406), .ZN(n5538) );
  OR2_X1 U7101 ( .A1(n5522), .A2(n10406), .ZN(n5523) );
  AOI22_X1 U7102 ( .A1(n5594), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5593), .B2(
        n7860), .ZN(n5524) );
  NAND2_X2 U7103 ( .A1(n5525), .A2(n5524), .ZN(n9573) );
  NAND2_X1 U7104 ( .A1(n6334), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U7105 ( .A1(n5798), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U7106 ( .A1(n5526), .A2(n9184), .ZN(n5527) );
  AND2_X1 U7107 ( .A1(n5543), .A2(n5527), .ZN(n9564) );
  NAND2_X1 U7108 ( .A1(n4596), .A2(n9564), .ZN(n5529) );
  NAND2_X1 U7109 ( .A1(n5382), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5528) );
  NAND4_X1 U7110 ( .A1(n5531), .A2(n5530), .A3(n5529), .A4(n5528), .ZN(n9204)
         );
  NOR2_X1 U7111 ( .A1(n9573), .A2(n9204), .ZN(n5533) );
  NAND2_X1 U7112 ( .A1(n9573), .A2(n9204), .ZN(n5532) );
  INV_X1 U7113 ( .A(SI_16_), .ZN(n5534) );
  XNOR2_X1 U7114 ( .A(n5535), .B(n5534), .ZN(n5536) );
  NAND2_X1 U7115 ( .A1(n7075), .A2(n6347), .ZN(n5541) );
  NAND2_X1 U7116 ( .A1(n5538), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5539) );
  XNOR2_X1 U7117 ( .A(n5539), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9292) );
  AOI22_X1 U7118 ( .A1(n5594), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5593), .B2(
        n9292), .ZN(n5540) );
  NAND2_X1 U7119 ( .A1(n5798), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U7120 ( .A1(n6334), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5548) );
  AND2_X1 U7121 ( .A1(n5543), .A2(n5542), .ZN(n5544) );
  NOR2_X1 U7122 ( .A1(n9093), .A2(n5544), .ZN(n9551) );
  NAND2_X1 U7123 ( .A1(n4596), .A2(n9551), .ZN(n5547) );
  INV_X1 U7124 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n5545) );
  OR2_X1 U7125 ( .A1(n5171), .A2(n5545), .ZN(n5546) );
  OR2_X1 U7126 ( .A1(n9548), .A2(n9092), .ZN(n6521) );
  NAND2_X1 U7127 ( .A1(n9548), .A2(n9092), .ZN(n6522) );
  NAND2_X1 U7128 ( .A1(n6521), .A2(n6522), .ZN(n6364) );
  INV_X1 U7129 ( .A(n9092), .ZN(n9203) );
  NAND2_X1 U7130 ( .A1(n9548), .A2(n9203), .ZN(n5550) );
  XNOR2_X1 U7131 ( .A(n5552), .B(n5551), .ZN(n7235) );
  NAND2_X1 U7132 ( .A1(n7235), .A2(n6347), .ZN(n5564) );
  NAND2_X1 U7133 ( .A1(n10406), .A2(n10235), .ZN(n5557) );
  NAND2_X1 U7134 ( .A1(n5555), .A2(n5554), .ZN(n5556) );
  NAND2_X1 U7135 ( .A1(n5560), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5559) );
  MUX2_X1 U7136 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5559), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n5561) );
  NOR2_X2 U7137 ( .A1(n5560), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n5702) );
  INV_X1 U7138 ( .A(n5702), .ZN(n5573) );
  NAND2_X1 U7139 ( .A1(n5561), .A2(n5573), .ZN(n9313) );
  INV_X1 U7140 ( .A(n9313), .ZN(n5562) );
  AOI22_X1 U7141 ( .A1(n5594), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5593), .B2(
        n5562), .ZN(n5563) );
  NAND2_X1 U7142 ( .A1(n5798), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U7143 ( .A1(n6334), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5568) );
  NOR2_X1 U7144 ( .A1(n9093), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5565) );
  NAND2_X1 U7145 ( .A1(n4596), .A2(n5140), .ZN(n5567) );
  NAND2_X1 U7146 ( .A1(n5382), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5566) );
  NAND4_X1 U7147 ( .A1(n5569), .A2(n5568), .A3(n5567), .A4(n5566), .ZN(n9202)
         );
  OR2_X1 U7148 ( .A1(n9536), .A2(n9202), .ZN(n5570) );
  XNOR2_X1 U7149 ( .A(n5572), .B(n5571), .ZN(n7305) );
  NAND2_X1 U7150 ( .A1(n7305), .A2(n6347), .ZN(n5580) );
  INV_X1 U7151 ( .A(n5574), .ZN(n5575) );
  NAND2_X1 U7152 ( .A1(n5575), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n5578) );
  INV_X1 U7153 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U7154 ( .A1(n5577), .A2(n5576), .ZN(n5591) );
  AND2_X1 U7155 ( .A1(n5578), .A2(n5591), .ZN(n9329) );
  AOI22_X1 U7156 ( .A1(n5594), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5593), .B2(
        n9329), .ZN(n5579) );
  NAND2_X1 U7157 ( .A1(n5798), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5586) );
  NAND2_X1 U7158 ( .A1(n6334), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5585) );
  OR2_X1 U7159 ( .A1(n5581), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5582) );
  AND2_X1 U7160 ( .A1(n5599), .A2(n5582), .ZN(n9516) );
  NAND2_X1 U7161 ( .A1(n4596), .A2(n9516), .ZN(n5584) );
  NAND2_X1 U7162 ( .A1(n5382), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5583) );
  NAND4_X1 U7163 ( .A1(n5586), .A2(n5585), .A3(n5584), .A4(n5583), .ZN(n9201)
         );
  NAND2_X1 U7164 ( .A1(n9632), .A2(n9201), .ZN(n5587) );
  XNOR2_X1 U7165 ( .A(n5590), .B(n5589), .ZN(n7419) );
  NAND2_X1 U7166 ( .A1(n7419), .A2(n6347), .ZN(n5596) );
  AOI22_X1 U7167 ( .A1(n5594), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5593), .B2(
        n9344), .ZN(n5595) );
  INV_X1 U7168 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9332) );
  INV_X1 U7169 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9327) );
  OAI22_X1 U7170 ( .A1(n5597), .A2(n9332), .B1(n5171), .B2(n9327), .ZN(n5604)
         );
  NAND2_X1 U7171 ( .A1(n5599), .A2(n5598), .ZN(n5600) );
  NAND2_X1 U7172 ( .A1(n5612), .A2(n5600), .ZN(n9044) );
  INV_X1 U7173 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n5601) );
  OAI22_X1 U7174 ( .A1(n9044), .A2(n5650), .B1(n5602), .B2(n5601), .ZN(n5603)
         );
  AND2_X1 U7175 ( .A1(n9628), .A2(n9200), .ZN(n5605) );
  OR2_X1 U7176 ( .A1(n9628), .A2(n9200), .ZN(n5606) );
  XNOR2_X1 U7177 ( .A(n5607), .B(n10288), .ZN(n5608) );
  XNOR2_X1 U7178 ( .A(n5609), .B(n5608), .ZN(n7555) );
  NAND2_X1 U7179 ( .A1(n7555), .A2(n6347), .ZN(n5611) );
  INV_X1 U7180 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7559) );
  OR2_X1 U7181 ( .A1(n5391), .A2(n7559), .ZN(n5610) );
  NAND2_X1 U7182 ( .A1(n5612), .A2(n9120), .ZN(n5613) );
  NAND2_X1 U7183 ( .A1(n5621), .A2(n5613), .ZN(n9494) );
  AOI22_X1 U7184 ( .A1(n6334), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n5798), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n5615) );
  NAND2_X1 U7185 ( .A1(n5382), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5614) );
  OAI211_X1 U7186 ( .C1(n9494), .C2(n5650), .A(n5615), .B(n5614), .ZN(n9199)
         );
  XNOR2_X1 U7187 ( .A(n5616), .B(SI_21_), .ZN(n5617) );
  XNOR2_X1 U7188 ( .A(n5618), .B(n5617), .ZN(n7597) );
  NAND2_X1 U7189 ( .A1(n7597), .A2(n6347), .ZN(n5620) );
  OR2_X1 U7190 ( .A1(n5391), .A2(n7612), .ZN(n5619) );
  AND2_X1 U7191 ( .A1(n5621), .A2(n9053), .ZN(n5622) );
  OR2_X1 U7192 ( .A1(n5622), .A2(n5630), .ZN(n9479) );
  AOI22_X1 U7193 ( .A1(n6334), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n5798), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n5624) );
  NAND2_X1 U7194 ( .A1(n5382), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5623) );
  OAI211_X1 U7195 ( .C1(n9479), .C2(n5650), .A(n5624), .B(n5623), .ZN(n9198)
         );
  AND2_X1 U7196 ( .A1(n9478), .A2(n9198), .ZN(n5625) );
  XNOR2_X1 U7197 ( .A(n5627), .B(n5626), .ZN(n7716) );
  NAND2_X1 U7198 ( .A1(n7716), .A2(n6347), .ZN(n5629) );
  OR2_X1 U7199 ( .A1(n5391), .A2(n10446), .ZN(n5628) );
  NOR2_X1 U7200 ( .A1(n5630), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5631) );
  OR2_X1 U7201 ( .A1(n5643), .A2(n5631), .ZN(n9458) );
  INV_X1 U7202 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U7203 ( .A1(n5798), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5633) );
  NAND2_X1 U7204 ( .A1(n5382), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5632) );
  OAI211_X1 U7205 ( .C1(n5597), .C2(n5634), .A(n5633), .B(n5632), .ZN(n5635)
         );
  INV_X1 U7206 ( .A(n5635), .ZN(n5636) );
  OAI21_X1 U7207 ( .B1(n9458), .B2(n5650), .A(n5636), .ZN(n9197) );
  NOR2_X1 U7208 ( .A1(n9612), .A2(n9197), .ZN(n5637) );
  NAND2_X1 U7209 ( .A1(n9612), .A2(n9197), .ZN(n5638) );
  XNOR2_X1 U7210 ( .A(n5640), .B(n5639), .ZN(n7723) );
  NAND2_X1 U7211 ( .A1(n7723), .A2(n6347), .ZN(n5642) );
  OR2_X1 U7212 ( .A1(n5391), .A2(n10278), .ZN(n5641) );
  NOR2_X1 U7213 ( .A1(n5643), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5644) );
  OR2_X1 U7214 ( .A1(n5656), .A2(n5644), .ZN(n9033) );
  INV_X1 U7215 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5647) );
  NAND2_X1 U7216 ( .A1(n5382), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U7217 ( .A1(n5798), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5645) );
  OAI211_X1 U7218 ( .C1(n5597), .C2(n5647), .A(n5646), .B(n5645), .ZN(n5648)
         );
  INV_X1 U7219 ( .A(n5648), .ZN(n5649) );
  OAI21_X1 U7220 ( .B1(n9033), .B2(n5650), .A(n5649), .ZN(n9145) );
  AOI21_X1 U7221 ( .B1(n5651), .B2(n4523), .A(n4553), .ZN(n9430) );
  XNOR2_X1 U7222 ( .A(n5653), .B(n5652), .ZN(n7807) );
  NAND2_X1 U7223 ( .A1(n7807), .A2(n6347), .ZN(n5655) );
  OR2_X1 U7224 ( .A1(n5391), .A2(n7818), .ZN(n5654) );
  OR2_X1 U7225 ( .A1(n5656), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U7226 ( .A1(n5657), .A2(n5668), .ZN(n9110) );
  INV_X1 U7227 ( .A(n9110), .ZN(n9434) );
  INV_X1 U7228 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5660) );
  NAND2_X1 U7229 ( .A1(n5382), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5659) );
  NAND2_X1 U7230 ( .A1(n5798), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5658) );
  OAI211_X1 U7231 ( .C1(n5597), .C2(n5660), .A(n5659), .B(n5658), .ZN(n5661)
         );
  AOI21_X1 U7232 ( .B1(n9434), .B2(n4596), .A(n5661), .ZN(n9071) );
  NAND2_X1 U7233 ( .A1(n9601), .A2(n9071), .ZN(n6456) );
  NAND2_X1 U7234 ( .A1(n9430), .A2(n9429), .ZN(n9431) );
  INV_X1 U7235 ( .A(n9071), .ZN(n9196) );
  NAND2_X1 U7236 ( .A1(n9601), .A2(n9196), .ZN(n5662) );
  NAND2_X1 U7237 ( .A1(n9431), .A2(n5662), .ZN(n9414) );
  XNOR2_X1 U7238 ( .A(n5664), .B(n5663), .ZN(n7879) );
  NAND2_X1 U7239 ( .A1(n7879), .A2(n6347), .ZN(n5666) );
  OR2_X1 U7240 ( .A1(n5391), .A2(n10477), .ZN(n5665) );
  NAND2_X1 U7241 ( .A1(n6334), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U7242 ( .A1(n5798), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5672) );
  INV_X1 U7243 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5669) );
  INV_X1 U7244 ( .A(n5682), .ZN(n5667) );
  AOI21_X1 U7245 ( .B1(n5669), .B2(n5668), .A(n5667), .ZN(n9419) );
  NAND2_X1 U7246 ( .A1(n4596), .A2(n9419), .ZN(n5671) );
  NAND2_X1 U7247 ( .A1(n5382), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5670) );
  NAND4_X1 U7248 ( .A1(n5673), .A2(n5672), .A3(n5671), .A4(n5670), .ZN(n9195)
         );
  OR2_X1 U7249 ( .A1(n9418), .A2(n9195), .ZN(n5674) );
  NAND2_X1 U7250 ( .A1(n9414), .A2(n5674), .ZN(n5676) );
  NAND2_X1 U7251 ( .A1(n9418), .A2(n9195), .ZN(n5675) );
  NAND2_X1 U7252 ( .A1(n9014), .A2(n6347), .ZN(n5680) );
  OR2_X1 U7253 ( .A1(n5391), .A2(n10490), .ZN(n5679) );
  NAND2_X1 U7254 ( .A1(n6334), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U7255 ( .A1(n5319), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5685) );
  AOI21_X1 U7256 ( .B1(n9172), .B2(n5682), .A(n5681), .ZN(n9403) );
  NAND2_X1 U7257 ( .A1(n4596), .A2(n9403), .ZN(n5684) );
  NAND2_X1 U7258 ( .A1(n5382), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5683) );
  OR2_X1 U7259 ( .A1(n9402), .A2(n9072), .ZN(n6463) );
  NAND2_X1 U7260 ( .A1(n9402), .A2(n9072), .ZN(n6466) );
  NAND2_X1 U7261 ( .A1(n6463), .A2(n6466), .ZN(n6371) );
  INV_X1 U7262 ( .A(n9072), .ZN(n9194) );
  OR2_X1 U7263 ( .A1(n9390), .A2(n9169), .ZN(n6492) );
  NAND2_X1 U7264 ( .A1(n9390), .A2(n9169), .ZN(n6317) );
  MUX2_X1 U7265 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n4511), .Z(n5790) );
  XNOR2_X1 U7266 ( .A(n5790), .B(n5791), .ZN(n5788) );
  NAND2_X1 U7267 ( .A1(n6198), .A2(n6347), .ZN(n5691) );
  INV_X1 U7268 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7975) );
  OR2_X1 U7269 ( .A1(n5391), .A2(n7975), .ZN(n5690) );
  NAND2_X1 U7270 ( .A1(n6334), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5699) );
  NAND2_X1 U7271 ( .A1(n5319), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5698) );
  INV_X1 U7272 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5692) );
  NAND2_X1 U7273 ( .A1(n5692), .A2(n5693), .ZN(n5695) );
  INV_X1 U7274 ( .A(n5693), .ZN(n5694) );
  NAND2_X1 U7275 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(n5694), .ZN(n5740) );
  NAND2_X1 U7276 ( .A1(n4596), .A2(n9375), .ZN(n5697) );
  NAND2_X1 U7277 ( .A1(n5382), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5696) );
  NAND2_X1 U7278 ( .A1(n8368), .A2(n8357), .ZN(n6318) );
  INV_X1 U7279 ( .A(n6374), .ZN(n5700) );
  XNOR2_X1 U7280 ( .A(n5787), .B(n5700), .ZN(n9374) );
  NAND2_X1 U7281 ( .A1(n5702), .A2(n5701), .ZN(n5706) );
  NAND2_X1 U7282 ( .A1(n5705), .A2(n5704), .ZN(n5703) );
  INV_X1 U7283 ( .A(n6872), .ZN(n6349) );
  NAND2_X2 U7284 ( .A1(n5711), .A2(n7557), .ZN(n6555) );
  OR2_X1 U7285 ( .A1(n6349), .A2(n6555), .ZN(n5710) );
  INV_X1 U7286 ( .A(n6884), .ZN(n5709) );
  AND2_X1 U7287 ( .A1(n5710), .A2(n5709), .ZN(n7006) );
  NAND2_X1 U7288 ( .A1(n6551), .A2(n5711), .ZN(n6849) );
  NAND2_X1 U7289 ( .A1(n6849), .A2(n6555), .ZN(n5712) );
  NAND2_X1 U7290 ( .A1(n7006), .A2(n5712), .ZN(n7688) );
  NAND2_X1 U7291 ( .A1(n6842), .A2(n9344), .ZN(n6468) );
  OR2_X1 U7292 ( .A1(n6468), .A2(n6883), .ZN(n7681) );
  INV_X1 U7293 ( .A(n9783), .ZN(n7232) );
  NAND2_X1 U7294 ( .A1(n6494), .A2(n7232), .ZN(n5714) );
  INV_X1 U7295 ( .A(n5715), .ZN(n5716) );
  INV_X1 U7296 ( .A(n9763), .ZN(n9754) );
  NAND2_X1 U7297 ( .A1(n9753), .A2(n9754), .ZN(n9752) );
  NAND2_X1 U7298 ( .A1(n9752), .A2(n5717), .ZN(n7086) );
  NAND2_X1 U7299 ( .A1(n7086), .A2(n6496), .ZN(n6393) );
  AND2_X1 U7300 ( .A1(n6394), .A2(n6392), .ZN(n5718) );
  NAND2_X1 U7301 ( .A1(n6393), .A2(n5718), .ZN(n5719) );
  INV_X1 U7302 ( .A(n9209), .ZN(n5721) );
  NAND2_X1 U7303 ( .A1(n7566), .A2(n5721), .ZN(n6407) );
  NAND2_X1 U7304 ( .A1(n6421), .A2(n7406), .ZN(n5720) );
  OR2_X1 U7305 ( .A1(n7566), .A2(n5721), .ZN(n7404) );
  NAND3_X1 U7306 ( .A1(n6409), .A2(n7404), .A3(n6398), .ZN(n5722) );
  AND2_X1 U7307 ( .A1(n5722), .A2(n6421), .ZN(n6505) );
  INV_X1 U7308 ( .A(n7385), .ZN(n6397) );
  INV_X1 U7309 ( .A(n7530), .ZN(n6360) );
  INV_X1 U7310 ( .A(n7689), .ZN(n5723) );
  NOR2_X1 U7311 ( .A1(n7694), .A2(n5723), .ZN(n5724) );
  INV_X1 U7312 ( .A(n7617), .ZN(n5725) );
  NOR2_X1 U7313 ( .A1(n7618), .A2(n5725), .ZN(n5726) );
  OR2_X1 U7314 ( .A1(n7740), .A2(n8025), .ZN(n6515) );
  NAND2_X1 U7315 ( .A1(n7740), .A2(n8025), .ZN(n6416) );
  INV_X1 U7316 ( .A(n9204), .ZN(n5728) );
  OR2_X1 U7317 ( .A1(n9573), .A2(n5728), .ZN(n6520) );
  NAND2_X1 U7318 ( .A1(n9573), .A2(n5728), .ZN(n6417) );
  NAND2_X1 U7319 ( .A1(n9543), .A2(n6522), .ZN(n9529) );
  INV_X1 U7320 ( .A(n9202), .ZN(n5729) );
  OR2_X1 U7321 ( .A1(n9536), .A2(n5729), .ZN(n6351) );
  NAND2_X1 U7322 ( .A1(n9536), .A2(n5729), .ZN(n6352) );
  NAND2_X1 U7323 ( .A1(n6351), .A2(n6352), .ZN(n9528) );
  INV_X1 U7324 ( .A(n9201), .ZN(n5730) );
  OR2_X1 U7325 ( .A1(n9632), .A2(n5730), .ZN(n6432) );
  NAND2_X1 U7326 ( .A1(n9632), .A2(n5730), .ZN(n6441) );
  NAND2_X1 U7327 ( .A1(n6432), .A2(n6441), .ZN(n9519) );
  INV_X1 U7328 ( .A(n9200), .ZN(n5731) );
  NAND2_X1 U7329 ( .A1(n9628), .A2(n5731), .ZN(n6527) );
  NAND2_X1 U7330 ( .A1(n6433), .A2(n6527), .ZN(n9501) );
  INV_X1 U7331 ( .A(n9199), .ZN(n5732) );
  NAND2_X1 U7332 ( .A1(n9623), .A2(n5732), .ZN(n6387) );
  NAND2_X1 U7333 ( .A1(n9488), .A2(n9487), .ZN(n5733) );
  INV_X1 U7334 ( .A(n9198), .ZN(n6308) );
  XNOR2_X1 U7335 ( .A(n9478), .B(n6308), .ZN(n9474) );
  NAND2_X1 U7336 ( .A1(n9478), .A2(n6308), .ZN(n6443) );
  INV_X1 U7337 ( .A(n9197), .ZN(n5734) );
  OR2_X1 U7338 ( .A1(n9612), .A2(n5734), .ZN(n6305) );
  NAND2_X1 U7339 ( .A1(n9612), .A2(n5734), .ZN(n6311) );
  AND2_X2 U7340 ( .A1(n6305), .A2(n6311), .ZN(n9462) );
  NAND2_X1 U7341 ( .A1(n5735), .A2(n6311), .ZN(n9442) );
  INV_X1 U7342 ( .A(n9145), .ZN(n5736) );
  OR2_X1 U7343 ( .A1(n9608), .A2(n5736), .ZN(n6450) );
  NAND2_X1 U7344 ( .A1(n9608), .A2(n5736), .ZN(n6451) );
  NAND2_X1 U7345 ( .A1(n9442), .A2(n9443), .ZN(n5737) );
  NAND2_X1 U7346 ( .A1(n5737), .A2(n6451), .ZN(n9425) );
  AND2_X1 U7347 ( .A1(n9658), .A2(n9195), .ZN(n6461) );
  INV_X1 U7348 ( .A(n9195), .ZN(n8116) );
  NAND2_X1 U7349 ( .A1(n9418), .A2(n8116), .ZN(n6458) );
  XNOR2_X1 U7350 ( .A(n5797), .B(n6374), .ZN(n5739) );
  NAND2_X1 U7351 ( .A1(n6551), .A2(n9344), .ZN(n5738) );
  NAND2_X1 U7352 ( .A1(n6844), .A2(n6883), .ZN(n6552) );
  NAND2_X1 U7353 ( .A1(n6334), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U7354 ( .A1(n5319), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5743) );
  INV_X1 U7355 ( .A(n5740), .ZN(n9366) );
  NAND2_X1 U7356 ( .A1(n4596), .A2(n9366), .ZN(n5742) );
  NAND2_X1 U7357 ( .A1(n5382), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5741) );
  INV_X1 U7358 ( .A(n7973), .ZN(n9232) );
  OR2_X1 U7359 ( .A1(n7077), .A2(n9168), .ZN(n5746) );
  INV_X1 U7360 ( .A(n9181), .ZN(n9091) );
  OR2_X1 U7361 ( .A1(n9169), .A2(n9091), .ZN(n5745) );
  INV_X1 U7362 ( .A(n9601), .ZN(n9436) );
  INV_X1 U7363 ( .A(n9612), .ZN(n9461) );
  INV_X1 U7364 ( .A(n9632), .ZN(n9518) );
  NAND2_X1 U7365 ( .A1(n9783), .A2(n7228), .ZN(n7227) );
  NAND2_X1 U7366 ( .A1(n9767), .A2(n9796), .ZN(n9766) );
  INV_X1 U7367 ( .A(n9704), .ZN(n7593) );
  INV_X1 U7368 ( .A(n9732), .ZN(n7806) );
  NOR2_X1 U7369 ( .A1(n9478), .A2(n9492), .ZN(n9477) );
  NAND2_X1 U7370 ( .A1(n9461), .A2(n9477), .ZN(n9455) );
  INV_X1 U7371 ( .A(n5806), .ZN(n5749) );
  AOI211_X1 U7372 ( .C1(n8368), .C2(n9387), .A(n9850), .B(n5749), .ZN(n9378)
         );
  AOI21_X1 U7373 ( .B1(n9374), .B2(n9845), .A(n5751), .ZN(n9584) );
  NAND2_X1 U7374 ( .A1(n5752), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5753) );
  MUX2_X1 U7375 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5753), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5754) );
  NAND2_X1 U7376 ( .A1(n5759), .A2(n5758), .ZN(n5756) );
  INV_X1 U7377 ( .A(n5780), .ZN(n9690) );
  NAND3_X1 U7378 ( .A1(n7883), .A2(P1_B_REG_SCAN_IN), .A3(n7820), .ZN(n5760)
         );
  OAI211_X1 U7379 ( .C1(P1_B_REG_SCAN_IN), .C2(n7820), .A(n5780), .B(n5760), 
        .ZN(n5775) );
  INV_X1 U7380 ( .A(n7883), .ZN(n5761) );
  OAI22_X1 U7381 ( .A1(n5775), .A2(P1_D_REG_1__SCAN_IN), .B1(n5780), .B2(n5761), .ZN(n6866) );
  INV_X1 U7382 ( .A(n5775), .ZN(n9774) );
  NOR4_X1 U7383 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5770) );
  NOR4_X1 U7384 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5769) );
  INV_X1 U7385 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n9779) );
  INV_X1 U7386 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9778) );
  INV_X1 U7387 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10251) );
  INV_X1 U7388 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9777) );
  NAND4_X1 U7389 ( .A1(n9779), .A2(n9778), .A3(n10251), .A4(n9777), .ZN(n5767)
         );
  NOR4_X1 U7390 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5765) );
  NOR4_X1 U7391 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5764) );
  NOR4_X1 U7392 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5763) );
  NOR4_X1 U7393 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5762) );
  NAND4_X1 U7394 ( .A1(n5765), .A2(n5764), .A3(n5763), .A4(n5762), .ZN(n5766)
         );
  NOR4_X1 U7395 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n5767), .A4(n5766), .ZN(n5768) );
  NAND3_X1 U7396 ( .A1(n5770), .A2(n5769), .A3(n5768), .ZN(n5771) );
  NAND2_X1 U7397 ( .A1(n9774), .A2(n5771), .ZN(n6865) );
  AND2_X1 U7398 ( .A1(n6866), .A2(n6865), .ZN(n5772) );
  AND2_X1 U7399 ( .A1(n6886), .A2(n5772), .ZN(n5818) );
  INV_X1 U7400 ( .A(n7820), .ZN(n5773) );
  OAI22_X1 U7401 ( .A1(n5775), .A2(P1_D_REG_0__SCAN_IN), .B1(n5780), .B2(n5773), .ZN(n5816) );
  INV_X1 U7402 ( .A(n5816), .ZN(n6868) );
  OR2_X1 U7403 ( .A1(n6878), .A2(n6868), .ZN(n6999) );
  NAND2_X1 U7404 ( .A1(n5777), .A2(n5776), .ZN(n5778) );
  NAND2_X1 U7405 ( .A1(n5778), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5779) );
  NOR2_X1 U7406 ( .A1(n6999), .A2(n9775), .ZN(n5782) );
  NAND2_X1 U7407 ( .A1(n8368), .A2(n5784), .ZN(n5785) );
  NAND2_X1 U7408 ( .A1(n5786), .A2(n5785), .ZN(P1_U3518) );
  INV_X1 U7409 ( .A(n5790), .ZN(n5792) );
  MUX2_X1 U7410 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n4511), .Z(n6324) );
  INV_X1 U7411 ( .A(SI_29_), .ZN(n5793) );
  NAND2_X1 U7412 ( .A1(n8142), .A2(n6347), .ZN(n5795) );
  INV_X1 U7413 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10476) );
  OR2_X1 U7414 ( .A1(n5391), .A2(n10476), .ZN(n5794) );
  NAND2_X1 U7415 ( .A1(n5811), .A2(n7077), .ZN(n6477) );
  XNOR2_X1 U7416 ( .A(n5796), .B(n6474), .ZN(n9371) );
  INV_X1 U7417 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U7418 ( .A1(n5382), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U7419 ( .A1(n5798), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5799) );
  OAI211_X1 U7420 ( .C1(n5597), .C2(n5801), .A(n5800), .B(n5799), .ZN(n9191)
         );
  INV_X1 U7421 ( .A(P1_B_REG_SCAN_IN), .ZN(n5802) );
  NOR2_X1 U7422 ( .A1(n9684), .A2(n5802), .ZN(n5803) );
  NOR2_X1 U7423 ( .A1(n9168), .A2(n5803), .ZN(n6674) );
  AOI22_X1 U7424 ( .A1(n9192), .A2(n9181), .B1(n9191), .B2(n6674), .ZN(n5804)
         );
  OAI21_X1 U7425 ( .B1(n5805), .B2(n9504), .A(n5804), .ZN(n9364) );
  AOI21_X1 U7426 ( .B1(n5811), .B2(n5806), .A(n9850), .ZN(n5807) );
  AND2_X1 U7427 ( .A1(n5807), .A2(n9356), .ZN(n9365) );
  AOI21_X1 U7428 ( .B1(n9371), .B2(n9845), .A(n5808), .ZN(n5820) );
  OR2_X1 U7429 ( .A1(n5820), .A2(n5809), .ZN(n5815) );
  INV_X1 U7430 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5810) );
  NOR2_X1 U7431 ( .A1(n9858), .A2(n5810), .ZN(n5813) );
  NOR2_X1 U7432 ( .A1(n5813), .A2(n5812), .ZN(n5814) );
  NAND2_X1 U7433 ( .A1(n5815), .A2(n5814), .ZN(P1_U3519) );
  OR2_X1 U7434 ( .A1(n9775), .A2(n5816), .ZN(n6700) );
  NOR2_X1 U7435 ( .A1(n6700), .A2(n6878), .ZN(n5817) );
  OR2_X1 U7436 ( .A1(n5820), .A2(n5819), .ZN(n5825) );
  INV_X1 U7437 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5822) );
  NOR2_X1 U7438 ( .A1(n9875), .A2(n5822), .ZN(n5823) );
  NAND2_X1 U7439 ( .A1(n5825), .A2(n5824), .ZN(P1_U3551) );
  NOR2_X1 U7440 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5830) );
  NAND4_X1 U7441 ( .A1(n5830), .A2(n5829), .A3(n5828), .A4(n5827), .ZN(n5833)
         );
  NAND4_X1 U7442 ( .A1(n6003), .A2(n5921), .A3(n6007), .A4(n5831), .ZN(n5832)
         );
  INV_X1 U7443 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5840) );
  OR2_X2 U7444 ( .A1(n5845), .A2(n9002), .ZN(n5857) );
  NAND2_X1 U7445 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), 
        .ZN(n5841) );
  NAND2_X1 U7446 ( .A1(n5857), .A2(n5841), .ZN(n5843) );
  XNOR2_X2 U7447 ( .A(n5843), .B(n5842), .ZN(n5848) );
  NOR2_X1 U7448 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n5844) );
  NAND2_X1 U7449 ( .A1(n5845), .A2(n5844), .ZN(n9003) );
  INV_X1 U7450 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n5847) );
  OR2_X1 U7451 ( .A1(n5988), .A2(n5847), .ZN(n5855) );
  INV_X2 U7452 ( .A(n5848), .ZN(n8144) );
  INV_X1 U7453 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n5849) );
  OR2_X1 U7454 ( .A1(n5909), .A2(n5849), .ZN(n5854) );
  INV_X1 U7455 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5851) );
  OR2_X1 U7456 ( .A1(n5898), .A2(n5851), .ZN(n5853) );
  NAND2_X2 U7457 ( .A1(n9007), .A2(n5848), .ZN(n5883) );
  INV_X1 U7458 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9888) );
  XNOR2_X2 U7459 ( .A(n5857), .B(n5856), .ZN(n6226) );
  INV_X1 U7460 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6687) );
  MUX2_X1 U7461 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5860), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5862) );
  INV_X1 U7462 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7215) );
  INV_X1 U7463 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9878) );
  INV_X1 U7464 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7210) );
  NOR2_X1 U7465 ( .A1(n5865), .A2(n5864), .ZN(n5867) );
  NAND2_X1 U7466 ( .A1(n5952), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U7467 ( .A1(n5867), .A2(n5866), .ZN(n6830) );
  NAND2_X1 U7468 ( .A1(n4514), .A2(SI_0_), .ZN(n5868) );
  XNOR2_X1 U7469 ( .A(n5868), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9019) );
  NAND2_X1 U7470 ( .A1(n6830), .A2(n6575), .ZN(n7054) );
  NAND2_X1 U7471 ( .A1(n7055), .A2(n7054), .ZN(n5872) );
  OR2_X1 U7472 ( .A1(n6572), .A2(n5870), .ZN(n5871) );
  NAND2_X1 U7473 ( .A1(n5872), .A2(n5871), .ZN(n8821) );
  INV_X2 U7474 ( .A(n5909), .ZN(n6192) );
  NAND2_X1 U7475 ( .A1(n6192), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5877) );
  INV_X1 U7476 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7150) );
  OR2_X1 U7477 ( .A1(n4509), .A2(n7150), .ZN(n5876) );
  INV_X1 U7478 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5873) );
  OR2_X1 U7479 ( .A1(n5898), .A2(n5873), .ZN(n5875) );
  INV_X1 U7480 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6945) );
  OR2_X1 U7481 ( .A1(n5883), .A2(n6945), .ZN(n5874) );
  INV_X1 U7482 ( .A(n5878), .ZN(n5879) );
  INV_X1 U7483 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6691) );
  OR2_X1 U7484 ( .A1(n8207), .A2(n6578), .ZN(n5880) );
  NAND2_X1 U7485 ( .A1(n5952), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5887) );
  INV_X1 U7486 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5882) );
  OR2_X1 U7487 ( .A1(n7094), .A2(n5882), .ZN(n5886) );
  OR2_X1 U7488 ( .A1(n4509), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5885) );
  INV_X1 U7489 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9925) );
  OR2_X1 U7490 ( .A1(n5883), .A2(n9925), .ZN(n5884) );
  NOR2_X1 U7491 ( .A1(n5878), .A2(n9002), .ZN(n5888) );
  MUX2_X1 U7492 ( .A(n9002), .B(n5888), .S(P2_IR_REG_3__SCAN_IN), .Z(n5889) );
  INV_X1 U7493 ( .A(n5889), .ZN(n5892) );
  INV_X1 U7494 ( .A(n5890), .ZN(n5891) );
  NAND2_X1 U7495 ( .A1(n5892), .A2(n5891), .ZN(n6968) );
  OR2_X1 U7496 ( .A1(n6020), .A2(n6686), .ZN(n5894) );
  INV_X1 U7497 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6685) );
  OR2_X1 U7498 ( .A1(n5905), .A2(n6685), .ZN(n5893) );
  OAI211_X1 U7499 ( .C1(n6229), .C2(n6968), .A(n5894), .B(n5893), .ZN(n10033)
         );
  NOR2_X1 U7500 ( .A1(n4507), .A2(n10033), .ZN(n5896) );
  NAND2_X1 U7501 ( .A1(n4507), .A2(n10033), .ZN(n5895) );
  NAND2_X1 U7502 ( .A1(n6192), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5903) );
  INV_X1 U7503 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6944) );
  OR2_X1 U7504 ( .A1(n5883), .A2(n6944), .ZN(n5902) );
  NOR2_X1 U7505 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5913) );
  AND2_X1 U7506 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5897) );
  NOR2_X1 U7507 ( .A1(n5913), .A2(n5897), .ZN(n7309) );
  OR2_X1 U7508 ( .A1(n4509), .A2(n7309), .ZN(n5901) );
  INV_X1 U7509 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5899) );
  OR2_X1 U7510 ( .A1(n5898), .A2(n5899), .ZN(n5900) );
  NAND4_X1 U7511 ( .A1(n5903), .A2(n5902), .A3(n5901), .A4(n5900), .ZN(n8212)
         );
  OR2_X1 U7512 ( .A1(n5890), .A2(n9002), .ZN(n5904) );
  XNOR2_X1 U7513 ( .A(n5904), .B(n5920), .ZN(n7035) );
  OR2_X1 U7514 ( .A1(n6020), .A2(n6689), .ZN(n5907) );
  OR2_X1 U7515 ( .A1(n5905), .A2(n4611), .ZN(n5906) );
  OAI211_X1 U7516 ( .C1(n6229), .C2(n7035), .A(n5907), .B(n5906), .ZN(n10039)
         );
  OR2_X1 U7517 ( .A1(n8212), .A2(n10039), .ZN(n6239) );
  NAND2_X1 U7518 ( .A1(n7281), .A2(n6239), .ZN(n5908) );
  NAND2_X1 U7519 ( .A1(n8212), .A2(n10039), .ZN(n6238) );
  NAND2_X1 U7520 ( .A1(n5908), .A2(n6238), .ZN(n7423) );
  INV_X1 U7521 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5910) );
  OR2_X1 U7522 ( .A1(n7094), .A2(n5910), .ZN(n5918) );
  NAND2_X1 U7523 ( .A1(n5913), .A2(n5912), .ZN(n5929) );
  OR2_X1 U7524 ( .A1(n5913), .A2(n5912), .ZN(n5914) );
  AND2_X1 U7525 ( .A1(n5929), .A2(n5914), .ZN(n7448) );
  OR2_X1 U7526 ( .A1(n4509), .A2(n7448), .ZN(n5917) );
  INV_X1 U7527 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5915) );
  OR2_X1 U7528 ( .A1(n5898), .A2(n5915), .ZN(n5916) );
  NAND2_X1 U7529 ( .A1(n5890), .A2(n5920), .ZN(n5935) );
  NAND2_X1 U7530 ( .A1(n5935), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5922) );
  XNOR2_X1 U7531 ( .A(n5922), .B(n5921), .ZN(n7182) );
  OR2_X1 U7532 ( .A1(n6020), .A2(n6693), .ZN(n5924) );
  INV_X1 U7533 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6692) );
  OR2_X1 U7534 ( .A1(n5905), .A2(n6692), .ZN(n5923) );
  OAI211_X1 U7535 ( .C1(n6229), .C2(n7182), .A(n5924), .B(n5923), .ZN(n8217)
         );
  OR2_X1 U7536 ( .A1(n8527), .A2(n8217), .ZN(n5925) );
  NAND2_X1 U7537 ( .A1(n8527), .A2(n8217), .ZN(n5926) );
  NAND2_X1 U7538 ( .A1(n6192), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5934) );
  INV_X1 U7539 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5928) );
  OR2_X1 U7540 ( .A1(n5898), .A2(n5928), .ZN(n5933) );
  NAND2_X1 U7541 ( .A1(n5929), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5930) );
  AND2_X1 U7542 ( .A1(n5940), .A2(n5930), .ZN(n7599) );
  OR2_X1 U7543 ( .A1(n4509), .A2(n7599), .ZN(n5932) );
  INV_X1 U7544 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7180) );
  OR2_X1 U7545 ( .A1(n7096), .A2(n7180), .ZN(n5931) );
  NAND4_X1 U7546 ( .A1(n5934), .A2(n5933), .A3(n5932), .A4(n5931), .ZN(n8526)
         );
  NAND2_X1 U7547 ( .A1(n5947), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5937) );
  INV_X1 U7548 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5936) );
  XNOR2_X1 U7549 ( .A(n5937), .B(n5936), .ZN(n7464) );
  OR2_X1 U7550 ( .A1(n6020), .A2(n6696), .ZN(n5939) );
  INV_X1 U7551 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6695) );
  OR2_X1 U7552 ( .A1(n5905), .A2(n6695), .ZN(n5938) );
  OAI211_X1 U7553 ( .C1(n6229), .C2(n7464), .A(n5939), .B(n5938), .ZN(n10047)
         );
  NAND2_X1 U7554 ( .A1(n6231), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5946) );
  INV_X1 U7555 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7661) );
  OR2_X1 U7556 ( .A1(n7094), .A2(n7661), .ZN(n5945) );
  AND2_X1 U7557 ( .A1(n5940), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5941) );
  NOR2_X1 U7558 ( .A1(n5954), .A2(n5941), .ZN(n7660) );
  OR2_X1 U7559 ( .A1(n4509), .A2(n7660), .ZN(n5944) );
  INV_X1 U7560 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5942) );
  OR2_X1 U7561 ( .A1(n5898), .A2(n5942), .ZN(n5943) );
  NAND4_X1 U7562 ( .A1(n5946), .A2(n5945), .A3(n5944), .A4(n5943), .ZN(n8525)
         );
  NOR2_X1 U7563 ( .A1(n5947), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n6005) );
  OR2_X1 U7564 ( .A1(n6005), .A2(n9002), .ZN(n5968) );
  XNOR2_X1 U7565 ( .A(n5968), .B(n6003), .ZN(n7475) );
  OR2_X1 U7566 ( .A1(n6020), .A2(n6699), .ZN(n5949) );
  INV_X1 U7567 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6698) );
  OR2_X1 U7568 ( .A1(n5905), .A2(n6698), .ZN(n5948) );
  NOR2_X1 U7569 ( .A1(n8525), .A2(n7663), .ZN(n5951) );
  NAND2_X1 U7570 ( .A1(n8525), .A2(n7663), .ZN(n5950) );
  NAND2_X1 U7571 ( .A1(n5952), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5960) );
  INV_X1 U7572 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5953) );
  OR2_X1 U7573 ( .A1(n5883), .A2(n5953), .ZN(n5959) );
  INV_X1 U7574 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7513) );
  OR2_X1 U7575 ( .A1(n7094), .A2(n7513), .ZN(n5958) );
  NOR2_X1 U7576 ( .A1(n5954), .A2(n7518), .ZN(n5955) );
  OR2_X1 U7577 ( .A1(n5975), .A2(n5955), .ZN(n7678) );
  INV_X1 U7578 ( .A(n7678), .ZN(n5956) );
  OR2_X1 U7579 ( .A1(n4509), .A2(n5956), .ZN(n5957) );
  NAND4_X1 U7580 ( .A1(n5960), .A2(n5959), .A3(n5958), .A4(n5957), .ZN(n8524)
         );
  NAND2_X1 U7581 ( .A1(n6705), .A2(n8148), .ZN(n5964) );
  NAND2_X1 U7582 ( .A1(n5968), .A2(n6003), .ZN(n5961) );
  NAND2_X1 U7583 ( .A1(n5961), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5962) );
  XNOR2_X1 U7584 ( .A(n5962), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7519) );
  AOI22_X1 U7585 ( .A1(n8147), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6682), .B2(
        n7519), .ZN(n5963) );
  NAND2_X1 U7586 ( .A1(n5965), .A2(n10057), .ZN(n5966) );
  NAND2_X1 U7587 ( .A1(n6720), .A2(n8148), .ZN(n5973) );
  OAI21_X1 U7588 ( .B1(P2_IR_REG_7__SCAN_IN), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5967) );
  INV_X1 U7589 ( .A(n5970), .ZN(n5969) );
  NAND2_X1 U7590 ( .A1(n5969), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5971) );
  INV_X1 U7591 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7592 ( .A1(n5970), .A2(n6001), .ZN(n5981) );
  AOI22_X1 U7593 ( .A1(n8147), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6682), .B2(
        n7912), .ZN(n5972) );
  NAND2_X1 U7594 ( .A1(n5952), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5980) );
  OR2_X1 U7595 ( .A1(n5883), .A2(n10095), .ZN(n5979) );
  INV_X1 U7596 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7752) );
  OR2_X1 U7597 ( .A1(n7094), .A2(n7752), .ZN(n5978) );
  OR2_X1 U7598 ( .A1(n5975), .A2(n5974), .ZN(n5976) );
  AND2_X1 U7599 ( .A1(n5986), .A2(n5976), .ZN(n7847) );
  OR2_X1 U7600 ( .A1(n4509), .A2(n7847), .ZN(n5977) );
  NAND4_X1 U7601 ( .A1(n5980), .A2(n5979), .A3(n5978), .A4(n5977), .ZN(n8523)
         );
  NAND2_X1 U7602 ( .A1(n10065), .A2(n8523), .ZN(n7822) );
  OR2_X1 U7603 ( .A1(n6725), .A2(n6020), .ZN(n5984) );
  NAND2_X1 U7604 ( .A1(n5981), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5982) );
  XNOR2_X1 U7605 ( .A(n5982), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7949) );
  AOI22_X1 U7606 ( .A1(n8147), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6682), .B2(
        n7949), .ZN(n5983) );
  NAND2_X1 U7607 ( .A1(n5952), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5992) );
  INV_X1 U7608 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5985) );
  OR2_X1 U7609 ( .A1(n5883), .A2(n5985), .ZN(n5991) );
  INV_X1 U7610 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7914) );
  OR2_X1 U7611 ( .A1(n7094), .A2(n7914), .ZN(n5990) );
  NAND2_X1 U7612 ( .A1(n5986), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5987) );
  AND2_X1 U7613 ( .A1(n6013), .A2(n5987), .ZN(n7933) );
  OR2_X1 U7614 ( .A1(n4509), .A2(n7933), .ZN(n5989) );
  NAND4_X1 U7615 ( .A1(n5992), .A2(n5991), .A3(n5990), .A4(n5989), .ZN(n8522)
         );
  NAND2_X1 U7616 ( .A1(n10071), .A2(n8522), .ZN(n5994) );
  AND2_X1 U7617 ( .A1(n7822), .A2(n5994), .ZN(n5993) );
  NAND2_X1 U7618 ( .A1(n7810), .A2(n5993), .ZN(n5999) );
  INV_X1 U7619 ( .A(n5994), .ZN(n5997) );
  OR2_X1 U7620 ( .A1(n10065), .A2(n8523), .ZN(n7823) );
  OR2_X1 U7621 ( .A1(n10071), .A2(n8522), .ZN(n5995) );
  AND2_X1 U7622 ( .A1(n7823), .A2(n5995), .ZN(n5996) );
  OR2_X1 U7623 ( .A1(n5997), .A2(n5996), .ZN(n5998) );
  NAND2_X1 U7624 ( .A1(n6736), .A2(n8148), .ZN(n6012) );
  INV_X1 U7625 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6002) );
  INV_X1 U7626 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6000) );
  AND4_X1 U7627 ( .A1(n6003), .A2(n6002), .A3(n6001), .A4(n6000), .ZN(n6004)
         );
  AND2_X1 U7628 ( .A1(n6005), .A2(n6004), .ZN(n6008) );
  NOR2_X1 U7629 ( .A1(n6008), .A2(n9002), .ZN(n6006) );
  MUX2_X1 U7630 ( .A(n9002), .B(n6006), .S(P2_IR_REG_11__SCAN_IN), .Z(n6010)
         );
  NAND2_X1 U7631 ( .A1(n6008), .A2(n6007), .ZN(n6032) );
  INV_X1 U7632 ( .A(n6032), .ZN(n6009) );
  AOI22_X1 U7633 ( .A1(n8147), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6682), .B2(
        n7965), .ZN(n6011) );
  NAND2_X1 U7634 ( .A1(n6012), .A2(n6011), .ZN(n7839) );
  NAND2_X1 U7635 ( .A1(n5952), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6018) );
  OR2_X1 U7636 ( .A1(n7096), .A2(n10099), .ZN(n6017) );
  INV_X1 U7637 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7884) );
  OR2_X1 U7638 ( .A1(n7094), .A2(n7884), .ZN(n6016) );
  NAND2_X1 U7639 ( .A1(n6013), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6014) );
  AND2_X1 U7640 ( .A1(n6024), .A2(n6014), .ZN(n8477) );
  OR2_X1 U7641 ( .A1(n4509), .A2(n8477), .ZN(n6015) );
  OR2_X1 U7642 ( .A1(n7839), .A2(n8403), .ZN(n8254) );
  NAND2_X1 U7643 ( .A1(n7839), .A2(n8403), .ZN(n8255) );
  NAND2_X1 U7644 ( .A1(n7839), .A2(n8805), .ZN(n6019) );
  NAND2_X1 U7645 ( .A1(n6032), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6021) );
  XNOR2_X1 U7646 ( .A(n6021), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8570) );
  AOI22_X1 U7647 ( .A1(n8147), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6682), .B2(
        n8570), .ZN(n6022) );
  NAND2_X2 U7648 ( .A1(n6023), .A2(n6022), .ZN(n8996) );
  NAND2_X1 U7649 ( .A1(n5952), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6028) );
  INV_X1 U7650 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8899) );
  OR2_X1 U7651 ( .A1(n5883), .A2(n8899), .ZN(n6027) );
  INV_X1 U7652 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7898) );
  OR2_X1 U7653 ( .A1(n7094), .A2(n7898), .ZN(n6026) );
  NOR2_X1 U7654 ( .A1(n6036), .A2(n5137), .ZN(n8809) );
  OR2_X1 U7655 ( .A1(n4509), .A2(n8809), .ZN(n6025) );
  NAND4_X1 U7656 ( .A1(n6028), .A2(n6027), .A3(n6026), .A4(n6025), .ZN(n8786)
         );
  OR2_X1 U7657 ( .A1(n8996), .A2(n8786), .ZN(n6029) );
  NAND2_X1 U7658 ( .A1(n8804), .A2(n6029), .ZN(n6031) );
  NAND2_X1 U7659 ( .A1(n8996), .A2(n8786), .ZN(n6030) );
  NAND2_X1 U7660 ( .A1(n6834), .A2(n8148), .ZN(n6035) );
  OR2_X1 U7661 ( .A1(n6032), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6033) );
  NAND2_X1 U7662 ( .A1(n6033), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6044) );
  XNOR2_X1 U7663 ( .A(n6044), .B(P2_IR_REG_13__SCAN_IN), .ZN(n9942) );
  AOI22_X1 U7664 ( .A1(n8147), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6682), .B2(
        n9942), .ZN(n6034) );
  NAND2_X1 U7665 ( .A1(n5952), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6041) );
  INV_X1 U7666 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8797) );
  OR2_X1 U7667 ( .A1(n7094), .A2(n8797), .ZN(n6040) );
  OR2_X1 U7668 ( .A1(n6036), .A2(n10509), .ZN(n6037) );
  NAND2_X1 U7669 ( .A1(n6036), .A2(n10509), .ZN(n6051) );
  AND2_X1 U7670 ( .A1(n6037), .A2(n6051), .ZN(n8789) );
  OR2_X1 U7671 ( .A1(n4509), .A2(n8789), .ZN(n6039) );
  INV_X1 U7672 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8896) );
  OR2_X1 U7673 ( .A1(n5883), .A2(n8896), .ZN(n6038) );
  NAND4_X1 U7674 ( .A1(n6041), .A2(n6040), .A3(n6039), .A4(n6038), .ZN(n8806)
         );
  AND2_X1 U7675 ( .A1(n8990), .A2(n8806), .ZN(n6042) );
  NAND2_X1 U7676 ( .A1(n6928), .A2(n8148), .ZN(n6050) );
  INV_X1 U7677 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7678 ( .A1(n6044), .A2(n6043), .ZN(n6045) );
  NAND2_X1 U7679 ( .A1(n6045), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6047) );
  INV_X1 U7680 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6046) );
  NAND2_X1 U7681 ( .A1(n6047), .A2(n6046), .ZN(n6059) );
  OR2_X1 U7682 ( .A1(n6047), .A2(n6046), .ZN(n6048) );
  AOI22_X1 U7683 ( .A1(n8147), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6682), .B2(
        n9957), .ZN(n6049) );
  NAND2_X1 U7684 ( .A1(n5952), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6056) );
  INV_X1 U7685 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8893) );
  OR2_X1 U7686 ( .A1(n5883), .A2(n8893), .ZN(n6055) );
  INV_X1 U7687 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8784) );
  OR2_X1 U7688 ( .A1(n7094), .A2(n8784), .ZN(n6054) );
  NAND2_X1 U7689 ( .A1(n6051), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6052) );
  AND2_X1 U7690 ( .A1(n6075), .A2(n6052), .ZN(n8776) );
  OR2_X1 U7691 ( .A1(n4509), .A2(n8776), .ZN(n6053) );
  NAND4_X1 U7692 ( .A1(n6056), .A2(n6055), .A3(n6054), .A4(n6053), .ZN(n8787)
         );
  NOR2_X1 U7693 ( .A1(n8984), .A2(n8787), .ZN(n6057) );
  NAND2_X1 U7694 ( .A1(n8984), .A2(n8787), .ZN(n6058) );
  NAND2_X1 U7695 ( .A1(n6995), .A2(n8148), .ZN(n6062) );
  NAND2_X1 U7696 ( .A1(n6059), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6060) );
  XNOR2_X1 U7697 ( .A(n6060), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9974) );
  AOI22_X1 U7698 ( .A1(n8147), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6682), .B2(
        n9974), .ZN(n6061) );
  NAND2_X1 U7699 ( .A1(n5952), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6066) );
  INV_X1 U7700 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9983) );
  OR2_X1 U7701 ( .A1(n7094), .A2(n9983), .ZN(n6065) );
  XNOR2_X1 U7702 ( .A(n6075), .B(n10462), .ZN(n8768) );
  OR2_X1 U7703 ( .A1(n4509), .A2(n8768), .ZN(n6064) );
  INV_X1 U7704 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8890) );
  OR2_X1 U7705 ( .A1(n5883), .A2(n8890), .ZN(n6063) );
  NAND2_X1 U7706 ( .A1(n8978), .A2(n8754), .ZN(n8277) );
  NAND2_X1 U7707 ( .A1(n8272), .A2(n8277), .ZN(n8270) );
  NAND2_X1 U7708 ( .A1(n8765), .A2(n8270), .ZN(n6068) );
  NAND2_X1 U7709 ( .A1(n8978), .A2(n8774), .ZN(n6067) );
  NAND2_X1 U7710 ( .A1(n6068), .A2(n6067), .ZN(n8751) );
  NAND2_X1 U7711 ( .A1(n7075), .A2(n8148), .ZN(n6072) );
  NAND2_X1 U7712 ( .A1(n6069), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6070) );
  XNOR2_X1 U7713 ( .A(n6070), .B(P2_IR_REG_16__SCAN_IN), .ZN(n9990) );
  AOI22_X1 U7714 ( .A1(n8147), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6682), .B2(
        n9990), .ZN(n6071) );
  NAND2_X1 U7715 ( .A1(n5952), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6080) );
  INV_X1 U7716 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8759) );
  OR2_X1 U7717 ( .A1(n7094), .A2(n8759), .ZN(n6079) );
  OAI21_X1 U7718 ( .B1(n6075), .B2(P2_REG3_REG_15__SCAN_IN), .A(
        P2_REG3_REG_16__SCAN_IN), .ZN(n6073) );
  INV_X1 U7719 ( .A(n6073), .ZN(n6076) );
  INV_X1 U7720 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10520) );
  NAND2_X1 U7721 ( .A1(n10462), .A2(n10520), .ZN(n6074) );
  OR2_X1 U7722 ( .A1(n6076), .A2(n6086), .ZN(n8423) );
  INV_X1 U7723 ( .A(n8423), .ZN(n8758) );
  OR2_X1 U7724 ( .A1(n4509), .A2(n8758), .ZN(n6078) );
  INV_X1 U7725 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8888) );
  OR2_X1 U7726 ( .A1(n7096), .A2(n8888), .ZN(n6077) );
  OR2_X1 U7727 ( .A1(n8887), .A2(n8509), .ZN(n8278) );
  NAND2_X1 U7728 ( .A1(n8887), .A2(n8509), .ZN(n8273) );
  NAND2_X1 U7729 ( .A1(n8278), .A2(n8273), .ZN(n8752) );
  NAND2_X1 U7730 ( .A1(n8751), .A2(n8752), .ZN(n6082) );
  NAND2_X1 U7731 ( .A1(n8887), .A2(n8766), .ZN(n6081) );
  NAND2_X1 U7732 ( .A1(n6082), .A2(n6081), .ZN(n8743) );
  NAND2_X1 U7733 ( .A1(n7235), .A2(n8148), .ZN(n6085) );
  NAND2_X1 U7734 ( .A1(n4581), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6083) );
  XNOR2_X1 U7735 ( .A(n6083), .B(P2_IR_REG_17__SCAN_IN), .ZN(n10009) );
  AOI22_X1 U7736 ( .A1(n8147), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6682), .B2(
        n10009), .ZN(n6084) );
  NAND2_X1 U7737 ( .A1(n5952), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6091) );
  INV_X1 U7738 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8883) );
  OR2_X1 U7739 ( .A1(n5883), .A2(n8883), .ZN(n6090) );
  INV_X1 U7740 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n10020) );
  OR2_X1 U7741 ( .A1(n7094), .A2(n10020), .ZN(n6089) );
  NOR2_X1 U7742 ( .A1(n6086), .A2(n8429), .ZN(n6087) );
  OR2_X1 U7743 ( .A1(n6099), .A2(n6087), .ZN(n8746) );
  INV_X1 U7744 ( .A(n8746), .ZN(n8432) );
  OR2_X1 U7745 ( .A1(n4509), .A2(n8432), .ZN(n6088) );
  NAND2_X1 U7746 ( .A1(n8968), .A2(n8756), .ZN(n8274) );
  NAND2_X1 U7747 ( .A1(n8281), .A2(n8274), .ZN(n8741) );
  NAND2_X1 U7748 ( .A1(n8743), .A2(n8741), .ZN(n6093) );
  INV_X1 U7749 ( .A(n8756), .ZN(n8521) );
  NAND2_X1 U7750 ( .A1(n8968), .A2(n8521), .ZN(n6092) );
  NAND2_X1 U7751 ( .A1(n7305), .A2(n8148), .ZN(n6098) );
  NAND2_X1 U7752 ( .A1(n6094), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U7753 ( .A1(n6095), .A2(n5836), .ZN(n6107) );
  OR2_X1 U7754 ( .A1(n6095), .A2(n5836), .ZN(n6096) );
  AND2_X1 U7755 ( .A1(n6107), .A2(n6096), .ZN(n8587) );
  AOI22_X1 U7756 ( .A1(n8147), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6682), .B2(
        n8587), .ZN(n6097) );
  NAND2_X1 U7757 ( .A1(n6231), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6104) );
  INV_X1 U7758 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8735) );
  OR2_X1 U7759 ( .A1(n7094), .A2(n8735), .ZN(n6103) );
  OR2_X1 U7760 ( .A1(n6099), .A2(n10450), .ZN(n6100) );
  AND2_X1 U7761 ( .A1(n6111), .A2(n6100), .ZN(n8734) );
  OR2_X1 U7762 ( .A1(n4509), .A2(n8734), .ZN(n6102) );
  INV_X1 U7763 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8962) );
  OR2_X1 U7764 ( .A1(n5898), .A2(n8962), .ZN(n6101) );
  NAND4_X1 U7765 ( .A1(n6104), .A2(n6103), .A3(n6102), .A4(n6101), .ZN(n8744)
         );
  AND2_X1 U7766 ( .A1(n8483), .A2(n8744), .ZN(n6105) );
  OR2_X1 U7767 ( .A1(n8483), .A2(n8744), .ZN(n6106) );
  NAND2_X1 U7768 ( .A1(n7419), .A2(n8148), .ZN(n6110) );
  NAND2_X1 U7769 ( .A1(n6107), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6108) );
  AOI22_X1 U7770 ( .A1(n8147), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8344), .B2(
        n6682), .ZN(n6109) );
  NAND2_X1 U7771 ( .A1(n5952), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6116) );
  INV_X1 U7772 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8584) );
  OR2_X1 U7773 ( .A1(n7094), .A2(n8584), .ZN(n6115) );
  NAND2_X1 U7774 ( .A1(n6111), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6112) );
  AND2_X1 U7775 ( .A1(n6122), .A2(n6112), .ZN(n8389) );
  OR2_X1 U7776 ( .A1(n4509), .A2(n8389), .ZN(n6114) );
  INV_X1 U7777 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8589) );
  OR2_X1 U7778 ( .A1(n5883), .A2(n8589), .ZN(n6113) );
  NAND2_X1 U7779 ( .A1(n8391), .A2(n8729), .ZN(n8290) );
  INV_X1 U7780 ( .A(n8729), .ZN(n8719) );
  NAND2_X1 U7781 ( .A1(n8391), .A2(n8719), .ZN(n6119) );
  NAND2_X1 U7782 ( .A1(n7555), .A2(n8148), .ZN(n6121) );
  INV_X1 U7783 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7556) );
  OR2_X1 U7784 ( .A1(n5905), .A2(n7556), .ZN(n6120) );
  AND2_X1 U7785 ( .A1(n6122), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6123) );
  OR2_X1 U7786 ( .A1(n6123), .A2(n6133), .ZN(n8722) );
  NAND2_X1 U7787 ( .A1(n5911), .A2(n8722), .ZN(n6127) );
  INV_X1 U7788 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8724) );
  OR2_X1 U7789 ( .A1(n7094), .A2(n8724), .ZN(n6126) );
  INV_X1 U7790 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8875) );
  OR2_X1 U7791 ( .A1(n7096), .A2(n8875), .ZN(n6125) );
  INV_X1 U7792 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8958) );
  OR2_X1 U7793 ( .A1(n5898), .A2(n8958), .ZN(n6124) );
  OR2_X1 U7794 ( .A1(n8874), .A2(n8398), .ZN(n8192) );
  NAND2_X1 U7795 ( .A1(n8874), .A2(n8398), .ZN(n8296) );
  NAND2_X1 U7796 ( .A1(n8192), .A2(n8296), .ZN(n8716) );
  OR2_X1 U7797 ( .A1(n8874), .A2(n8705), .ZN(n6128) );
  NAND2_X1 U7798 ( .A1(n7597), .A2(n8148), .ZN(n6130) );
  OR2_X1 U7799 ( .A1(n5905), .A2(n7598), .ZN(n6129) );
  NAND2_X1 U7800 ( .A1(n6192), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U7801 ( .A1(n6231), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6131) );
  AND2_X1 U7802 ( .A1(n6132), .A2(n6131), .ZN(n6137) );
  NOR2_X1 U7803 ( .A1(n6133), .A2(n10491), .ZN(n6134) );
  OR2_X1 U7804 ( .A1(n6143), .A2(n6134), .ZN(n8708) );
  NAND2_X1 U7805 ( .A1(n8708), .A2(n5911), .ZN(n6136) );
  NAND2_X1 U7806 ( .A1(n5952), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7807 ( .A1(n8193), .A2(n8298), .ZN(n8703) );
  INV_X1 U7808 ( .A(n8691), .ZN(n8718) );
  OR2_X1 U7809 ( .A1(n8953), .A2(n8718), .ZN(n6138) );
  NAND2_X1 U7810 ( .A1(n6139), .A2(n6138), .ZN(n8688) );
  NAND2_X1 U7811 ( .A1(n7716), .A2(n8148), .ZN(n6141) );
  OR2_X1 U7812 ( .A1(n5905), .A2(n7718), .ZN(n6140) );
  INV_X1 U7813 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n6142) );
  OR2_X1 U7814 ( .A1(n6143), .A2(n6142), .ZN(n6144) );
  NAND2_X1 U7815 ( .A1(n6152), .A2(n6144), .ZN(n8696) );
  NAND2_X1 U7816 ( .A1(n8696), .A2(n5911), .ZN(n6147) );
  AOI22_X1 U7817 ( .A1(n6231), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n6192), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7818 ( .A1(n5952), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U7819 ( .A1(n8695), .A2(n6148), .ZN(n8301) );
  NAND2_X1 U7820 ( .A1(n8300), .A2(n8301), .ZN(n8693) );
  OR2_X1 U7821 ( .A1(n8695), .A2(n8704), .ZN(n6149) );
  NAND2_X1 U7822 ( .A1(n7723), .A2(n8148), .ZN(n6151) );
  OR2_X1 U7823 ( .A1(n5905), .A2(n7725), .ZN(n6150) );
  INV_X1 U7824 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8863) );
  NAND2_X1 U7825 ( .A1(n6152), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7826 ( .A1(n6160), .A2(n6153), .ZN(n8685) );
  NAND2_X1 U7827 ( .A1(n8685), .A2(n5911), .ZN(n6155) );
  AOI22_X1 U7828 ( .A1(n6192), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n5952), .B2(
        P2_REG0_REG_23__SCAN_IN), .ZN(n6154) );
  OAI211_X1 U7829 ( .C1(n7096), .C2(n8863), .A(n6155), .B(n6154), .ZN(n8672)
         );
  NAND2_X1 U7830 ( .A1(n8943), .A2(n8672), .ZN(n6156) );
  NAND2_X1 U7831 ( .A1(n6157), .A2(n6156), .ZN(n8669) );
  NAND2_X1 U7832 ( .A1(n7807), .A2(n8148), .ZN(n6159) );
  OR2_X1 U7833 ( .A1(n5905), .A2(n7808), .ZN(n6158) );
  NAND2_X1 U7834 ( .A1(n6160), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U7835 ( .A1(n6171), .A2(n6161), .ZN(n8676) );
  NAND2_X1 U7836 ( .A1(n8676), .A2(n5911), .ZN(n6166) );
  INV_X1 U7837 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8860) );
  NAND2_X1 U7838 ( .A1(n6192), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U7839 ( .A1(n5952), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6162) );
  OAI211_X1 U7840 ( .C1(n8860), .C2(n7096), .A(n6163), .B(n6162), .ZN(n6164)
         );
  INV_X1 U7841 ( .A(n6164), .ZN(n6165) );
  AND2_X1 U7842 ( .A1(n8937), .A2(n8682), .ZN(n6168) );
  NAND2_X1 U7843 ( .A1(n7879), .A2(n8148), .ZN(n6170) );
  OR2_X1 U7844 ( .A1(n5905), .A2(n7880), .ZN(n6169) );
  INV_X1 U7845 ( .A(n6182), .ZN(n6173) );
  NAND2_X1 U7846 ( .A1(n6171), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U7847 ( .A1(n6173), .A2(n6172), .ZN(n8662) );
  NAND2_X1 U7848 ( .A1(n8662), .A2(n5911), .ZN(n6178) );
  INV_X1 U7849 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8857) );
  NAND2_X1 U7850 ( .A1(n6192), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7851 ( .A1(n5952), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6174) );
  OAI211_X1 U7852 ( .C1(n5883), .C2(n8857), .A(n6175), .B(n6174), .ZN(n6176)
         );
  INV_X1 U7853 ( .A(n6176), .ZN(n6177) );
  NAND2_X1 U7854 ( .A1(n8931), .A2(n8647), .ZN(n8314) );
  NAND2_X1 U7855 ( .A1(n8315), .A2(n8314), .ZN(n8656) );
  NOR2_X1 U7856 ( .A1(n8931), .A2(n8671), .ZN(n6179) );
  NAND2_X1 U7857 ( .A1(n9014), .A2(n8148), .ZN(n6181) );
  OR2_X1 U7858 ( .A1(n5905), .A2(n9016), .ZN(n6180) );
  INV_X1 U7859 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10488) );
  NOR2_X1 U7860 ( .A1(n6182), .A2(n10488), .ZN(n6183) );
  INV_X1 U7861 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8854) );
  NAND2_X1 U7862 ( .A1(n5952), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6185) );
  NAND2_X1 U7863 ( .A1(n6192), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6184) );
  OAI211_X1 U7864 ( .C1(n5883), .C2(n8854), .A(n6185), .B(n6184), .ZN(n6186)
         );
  AOI21_X1 U7865 ( .B1(n8651), .B2(n5911), .A(n6186), .ZN(n6666) );
  NAND2_X1 U7866 ( .A1(n6641), .A2(n6666), .ZN(n6187) );
  NAND2_X1 U7867 ( .A1(n7991), .A2(n8148), .ZN(n6189) );
  OR2_X1 U7868 ( .A1(n5905), .A2(n7992), .ZN(n6188) );
  INV_X1 U7869 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6663) );
  OR2_X1 U7870 ( .A1(n6190), .A2(n6663), .ZN(n6191) );
  NAND2_X1 U7871 ( .A1(n6190), .A2(n6663), .ZN(n6203) );
  NAND2_X1 U7872 ( .A1(n6191), .A2(n6203), .ZN(n8639) );
  NAND2_X1 U7873 ( .A1(n8639), .A2(n5911), .ZN(n6197) );
  INV_X1 U7874 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8851) );
  NAND2_X1 U7875 ( .A1(n6192), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7876 ( .A1(n5952), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6193) );
  OAI211_X1 U7877 ( .C1(n8851), .C2(n7096), .A(n6194), .B(n6193), .ZN(n6195)
         );
  INV_X1 U7878 ( .A(n6195), .ZN(n6196) );
  NAND2_X1 U7879 ( .A1(n8919), .A2(n8645), .ZN(n6254) );
  NAND2_X1 U7880 ( .A1(n6198), .A2(n8148), .ZN(n6200) );
  INV_X1 U7881 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9013) );
  OR2_X1 U7882 ( .A1(n5905), .A2(n9013), .ZN(n6199) );
  NAND2_X1 U7883 ( .A1(n6231), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6208) );
  INV_X1 U7884 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8628) );
  OR2_X1 U7885 ( .A1(n7094), .A2(n8628), .ZN(n6207) );
  INV_X1 U7886 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6202) );
  INV_X1 U7887 ( .A(n6203), .ZN(n6201) );
  NAND2_X1 U7888 ( .A1(n6202), .A2(n6201), .ZN(n8606) );
  NAND2_X1 U7889 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(n6203), .ZN(n6204) );
  OR2_X1 U7890 ( .A1(n4509), .A2(n8629), .ZN(n6206) );
  INV_X1 U7891 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8912) );
  OR2_X1 U7892 ( .A1(n5898), .A2(n8912), .ZN(n6205) );
  NAND2_X1 U7893 ( .A1(n6210), .A2(n6209), .ZN(n6211) );
  NAND2_X1 U7894 ( .A1(n8142), .A2(n8148), .ZN(n6213) );
  INV_X1 U7895 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8143) );
  OR2_X1 U7896 ( .A1(n5905), .A2(n8143), .ZN(n6212) );
  INV_X1 U7897 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n6214) );
  OR2_X1 U7898 ( .A1(n7094), .A2(n6214), .ZN(n6217) );
  INV_X1 U7899 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8844) );
  OR2_X1 U7900 ( .A1(n7096), .A2(n8844), .ZN(n6216) );
  INV_X1 U7901 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6302) );
  OR2_X1 U7902 ( .A1(n5898), .A2(n6302), .ZN(n6215) );
  NAND2_X1 U7903 ( .A1(n8324), .A2(n8623), .ZN(n8152) );
  NAND2_X1 U7904 ( .A1(n8328), .A2(n8152), .ZN(n8188) );
  XNOR2_X1 U7905 ( .A(n6218), .B(n8188), .ZN(n6261) );
  NAND2_X1 U7906 ( .A1(n6219), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7907 ( .A1(n8348), .A2(n8344), .ZN(n6294) );
  NAND2_X1 U7908 ( .A1(n4661), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6222) );
  MUX2_X1 U7909 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6222), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n6223) );
  NAND2_X1 U7910 ( .A1(n4564), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U7911 ( .A1(n8195), .A2(n6293), .ZN(n6225) );
  NAND2_X1 U7912 ( .A1(n6939), .A2(n8346), .ZN(n6228) );
  NAND2_X1 U7913 ( .A1(n6229), .A2(n6228), .ZN(n6664) );
  NAND2_X2 U7914 ( .A1(n8348), .A2(n8195), .ZN(n8326) );
  AND2_X1 U7915 ( .A1(n6229), .A2(P2_B_REG_SCAN_IN), .ZN(n6230) );
  NOR2_X1 U7916 ( .A1(n8757), .A2(n6230), .ZN(n8604) );
  NAND2_X1 U7917 ( .A1(n6231), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6236) );
  INV_X1 U7918 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6232) );
  OR2_X1 U7919 ( .A1(n7094), .A2(n6232), .ZN(n6235) );
  INV_X1 U7920 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6233) );
  OR2_X1 U7921 ( .A1(n5898), .A2(n6233), .ZN(n6234) );
  NAND4_X1 U7922 ( .A1(n7101), .A2(n6236), .A3(n6235), .A4(n6234), .ZN(n8519)
         );
  INV_X1 U7923 ( .A(n6664), .ZN(n6662) );
  AOI22_X1 U7924 ( .A1(n8604), .A2(n8519), .B1(n8636), .B2(n8827), .ZN(n6260)
         );
  INV_X1 U7925 ( .A(n10047), .ZN(n7491) );
  NAND2_X1 U7926 ( .A1(n8526), .A2(n7491), .ZN(n8231) );
  INV_X1 U7927 ( .A(n6830), .ZN(n7135) );
  OR2_X1 U7928 ( .A1(n8207), .A2(n10028), .ZN(n8206) );
  NAND2_X1 U7929 ( .A1(n8817), .A2(n8206), .ZN(n7274) );
  INV_X1 U7930 ( .A(n10033), .ZN(n7277) );
  OR2_X1 U7931 ( .A1(n8825), .A2(n7277), .ZN(n8223) );
  NAND2_X1 U7932 ( .A1(n4507), .A2(n7277), .ZN(n8216) );
  NAND2_X1 U7933 ( .A1(n6239), .A2(n6238), .ZN(n8162) );
  INV_X1 U7934 ( .A(n10039), .ZN(n8211) );
  OR2_X1 U7935 ( .A1(n8212), .A2(n8211), .ZN(n8219) );
  NAND2_X1 U7936 ( .A1(n7425), .A2(n8218), .ZN(n6240) );
  INV_X1 U7937 ( .A(n8217), .ZN(n10044) );
  OR2_X1 U7938 ( .A1(n7425), .A2(n8218), .ZN(n7484) );
  OR2_X1 U7939 ( .A1(n8526), .A2(n7491), .ZN(n8229) );
  NAND2_X1 U7940 ( .A1(n6241), .A2(n8229), .ZN(n7655) );
  NAND2_X1 U7941 ( .A1(n8525), .A2(n10053), .ZN(n8237) );
  AND2_X1 U7942 ( .A1(n10057), .A2(n8524), .ZN(n8239) );
  NAND2_X1 U7943 ( .A1(n10065), .A2(n7676), .ZN(n8244) );
  NAND2_X1 U7944 ( .A1(n8240), .A2(n8244), .ZN(n8172) );
  INV_X1 U7945 ( .A(n8522), .ZN(n8475) );
  OR2_X1 U7946 ( .A1(n10071), .A2(n8475), .ZN(n8253) );
  NAND2_X1 U7947 ( .A1(n10071), .A2(n8475), .ZN(n8250) );
  NAND2_X1 U7948 ( .A1(n8253), .A2(n8250), .ZN(n8173) );
  OR2_X2 U7949 ( .A1(n8996), .A2(n8453), .ZN(n8261) );
  NAND2_X1 U7950 ( .A1(n8996), .A2(n8453), .ZN(n8260) );
  NAND2_X1 U7951 ( .A1(n8261), .A2(n8260), .ZN(n8798) );
  INV_X1 U7952 ( .A(n8255), .ZN(n8799) );
  NOR2_X1 U7953 ( .A1(n8990), .A2(n6609), .ZN(n8263) );
  NAND2_X1 U7954 ( .A1(n8990), .A2(n6609), .ZN(n8264) );
  INV_X1 U7955 ( .A(n8787), .ZN(n6612) );
  OR2_X1 U7956 ( .A1(n8984), .A2(n6612), .ZN(n8267) );
  AND2_X1 U7957 ( .A1(n8984), .A2(n6612), .ZN(n8269) );
  NAND2_X1 U7958 ( .A1(n8763), .A2(n8277), .ZN(n6243) );
  NAND2_X1 U7959 ( .A1(n8740), .A2(n8281), .ZN(n6244) );
  NAND2_X1 U7960 ( .A1(n6244), .A2(n8274), .ZN(n8732) );
  INV_X1 U7961 ( .A(n8732), .ZN(n6245) );
  NAND2_X1 U7962 ( .A1(n8483), .A2(n6620), .ZN(n8285) );
  NAND2_X1 U7963 ( .A1(n6246), .A2(n8286), .ZN(n7976) );
  NAND2_X1 U7964 ( .A1(n7976), .A2(n8290), .ZN(n8712) );
  AND2_X1 U7965 ( .A1(n8192), .A2(n8711), .ZN(n8289) );
  NAND2_X1 U7966 ( .A1(n6247), .A2(n8193), .ZN(n8694) );
  NAND2_X1 U7967 ( .A1(n8694), .A2(n8301), .ZN(n6248) );
  NAND2_X1 U7968 ( .A1(n8937), .A2(n8414), .ZN(n8308) );
  INV_X1 U7969 ( .A(n8672), .ZN(n8692) );
  NAND2_X1 U7970 ( .A1(n8943), .A2(n8692), .ZN(n8666) );
  NAND2_X1 U7971 ( .A1(n8679), .A2(n6249), .ZN(n6251) );
  INV_X1 U7972 ( .A(n6249), .ZN(n8306) );
  NAND2_X1 U7973 ( .A1(n6251), .A2(n8309), .ZN(n8655) );
  NOR2_X1 U7974 ( .A1(n8925), .A2(n6666), .ZN(n8318) );
  INV_X1 U7975 ( .A(n8318), .ZN(n6252) );
  NAND2_X1 U7976 ( .A1(n8925), .A2(n6666), .ZN(n8319) );
  NAND2_X1 U7977 ( .A1(n6253), .A2(n8319), .ZN(n8633) );
  INV_X1 U7978 ( .A(n8323), .ZN(n6255) );
  NAND2_X1 U7979 ( .A1(n8618), .A2(n8620), .ZN(n6257) );
  OR2_X1 U7980 ( .A1(n8913), .A2(n6209), .ZN(n6256) );
  NAND2_X1 U7981 ( .A1(n6257), .A2(n6256), .ZN(n8150) );
  NAND2_X1 U7982 ( .A1(n8348), .A2(n8596), .ZN(n7059) );
  INV_X1 U7983 ( .A(n7059), .ZN(n6258) );
  NOR2_X1 U7984 ( .A1(n8161), .A2(n6293), .ZN(n7275) );
  NAND2_X1 U7985 ( .A1(n6258), .A2(n7275), .ZN(n7208) );
  NAND2_X1 U7986 ( .A1(n8596), .A2(n8343), .ZN(n6650) );
  NAND2_X1 U7987 ( .A1(n7059), .A2(n6650), .ZN(n6259) );
  AND2_X1 U7988 ( .A1(n8344), .A2(n8343), .ZN(n6296) );
  NAND2_X1 U7989 ( .A1(n6291), .A2(n6292), .ZN(n6262) );
  XNOR2_X1 U7990 ( .A(n6276), .B(P2_B_REG_SCAN_IN), .ZN(n6273) );
  NAND2_X1 U7991 ( .A1(n4565), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6269) );
  MUX2_X1 U7992 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6269), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6272) );
  INV_X1 U7993 ( .A(n6270), .ZN(n6271) );
  INV_X1 U7994 ( .A(n9017), .ZN(n6274) );
  INV_X1 U7995 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6734) );
  NAND2_X1 U7996 ( .A1(n6275), .A2(n6734), .ZN(n6277) );
  NAND2_X1 U7997 ( .A1(n9017), .A2(n6276), .ZN(n6732) );
  AND2_X1 U7998 ( .A1(n7062), .A2(n6565), .ZN(n7204) );
  NOR2_X1 U7999 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6281) );
  NOR4_X1 U8000 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6280) );
  NOR4_X1 U8001 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6279) );
  NOR4_X1 U8002 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n6278) );
  NAND4_X1 U8003 ( .A1(n6281), .A2(n6280), .A3(n6279), .A4(n6278), .ZN(n6287)
         );
  NOR4_X1 U8004 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6285) );
  NOR4_X1 U8005 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6284) );
  NOR4_X1 U8006 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6283) );
  NOR4_X1 U8007 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6282) );
  NAND4_X1 U8008 ( .A1(n6285), .A2(n6284), .A3(n6283), .A4(n6282), .ZN(n6286)
         );
  NOR2_X1 U8009 ( .A1(n6287), .A2(n6286), .ZN(n6288) );
  NOR2_X1 U8010 ( .A1(n9017), .A2(n6276), .ZN(n6289) );
  AND2_X1 U8011 ( .A1(n8326), .A2(n10078), .ZN(n6295) );
  NAND2_X1 U8012 ( .A1(n8161), .A2(n6293), .ZN(n6566) );
  NAND2_X1 U8013 ( .A1(n6295), .A2(n6655), .ZN(n6644) );
  OR2_X1 U8014 ( .A1(n6661), .A2(n6651), .ZN(n6300) );
  INV_X1 U8015 ( .A(n6655), .ZN(n6298) );
  INV_X1 U8016 ( .A(n7208), .ZN(n6657) );
  NAND2_X1 U8017 ( .A1(n7068), .A2(n7067), .ZN(n6297) );
  OAI21_X1 U8018 ( .B1(n6298), .B2(n6657), .A(n6648), .ZN(n6299) );
  NOR2_X1 U8019 ( .A1(n10084), .A2(n6302), .ZN(n6303) );
  INV_X1 U8020 ( .A(n6455), .ZN(n6307) );
  NAND2_X1 U8021 ( .A1(n6450), .A2(n6305), .ZN(n6384) );
  AND3_X1 U8022 ( .A1(n6456), .A2(n6451), .A3(n6384), .ZN(n6306) );
  OR3_X1 U8023 ( .A1(n6461), .A2(n6307), .A3(n6306), .ZN(n6315) );
  INV_X1 U8024 ( .A(n6315), .ZN(n6310) );
  OR2_X1 U8025 ( .A1(n9478), .A2(n6308), .ZN(n6436) );
  NAND2_X1 U8026 ( .A1(n6436), .A2(n6386), .ZN(n6438) );
  INV_X1 U8027 ( .A(n6438), .ZN(n6309) );
  NAND3_X1 U8028 ( .A1(n6310), .A2(n6309), .A3(n6463), .ZN(n6532) );
  NOR2_X1 U8029 ( .A1(n6532), .A2(n9488), .ZN(n6322) );
  NAND2_X1 U8030 ( .A1(n6451), .A2(n6311), .ZN(n6385) );
  INV_X1 U8031 ( .A(n6385), .ZN(n6313) );
  NAND2_X1 U8032 ( .A1(n6443), .A2(n6387), .ZN(n6312) );
  NAND2_X1 U8033 ( .A1(n6312), .A2(n6436), .ZN(n6448) );
  AND3_X1 U8034 ( .A1(n6456), .A2(n6313), .A3(n6448), .ZN(n6314) );
  OAI21_X1 U8035 ( .B1(n6315), .B2(n6314), .A(n6458), .ZN(n6316) );
  AND3_X1 U8036 ( .A1(n6316), .A2(n6492), .A3(n6463), .ZN(n6321) );
  AND2_X1 U8037 ( .A1(n6318), .A2(n6317), .ZN(n6382) );
  INV_X1 U8038 ( .A(n6382), .ZN(n6472) );
  INV_X1 U8039 ( .A(n6466), .ZN(n6319) );
  AND2_X1 U8040 ( .A1(n6492), .A2(n6319), .ZN(n6320) );
  OR3_X1 U8041 ( .A1(n6321), .A2(n6472), .A3(n6320), .ZN(n6491) );
  AOI21_X1 U8042 ( .B1(n6322), .B2(n6492), .A(n6491), .ZN(n6338) );
  NAND2_X1 U8043 ( .A1(n6476), .A2(n4904), .ZN(n6490) );
  NAND2_X1 U8044 ( .A1(n6323), .A2(SI_29_), .ZN(n6328) );
  INV_X1 U8045 ( .A(n6324), .ZN(n6325) );
  INV_X1 U8046 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8141) );
  INV_X1 U8047 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9009) );
  MUX2_X1 U8048 ( .A(n8141), .B(n9009), .S(n4513), .Z(n6329) );
  INV_X1 U8049 ( .A(SI_30_), .ZN(n10327) );
  NAND2_X1 U8050 ( .A1(n6329), .A2(n10327), .ZN(n6340) );
  INV_X1 U8051 ( .A(n6329), .ZN(n6330) );
  NAND2_X1 U8052 ( .A1(n6330), .A2(SI_30_), .ZN(n6331) );
  NAND2_X1 U8053 ( .A1(n6340), .A2(n6331), .ZN(n6341) );
  NAND2_X1 U8054 ( .A1(n8146), .A2(n6347), .ZN(n6333) );
  OR2_X1 U8055 ( .A1(n5391), .A2(n8141), .ZN(n6332) );
  NAND2_X1 U8056 ( .A1(n6334), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6337) );
  NAND2_X1 U8057 ( .A1(n5382), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U8058 ( .A1(n5319), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6335) );
  NAND3_X1 U8059 ( .A1(n6337), .A2(n6336), .A3(n6335), .ZN(n9190) );
  OAI22_X1 U8060 ( .A1(n6338), .A2(n6490), .B1(n9649), .B2(n9190), .ZN(n6339)
         );
  INV_X1 U8061 ( .A(n9191), .ZN(n6480) );
  NAND2_X1 U8062 ( .A1(n9357), .A2(n6480), .ZN(n6375) );
  NAND2_X1 U8063 ( .A1(n6375), .A2(n6477), .ZN(n6536) );
  INV_X1 U8064 ( .A(n9190), .ZN(n6481) );
  OR2_X1 U8065 ( .A1(n9357), .A2(n6480), .ZN(n6377) );
  OAI22_X1 U8066 ( .A1(n6339), .A2(n6536), .B1(n6481), .B2(n6377), .ZN(n6350)
         );
  MUX2_X1 U8067 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n4514), .Z(n6343) );
  INV_X1 U8068 ( .A(SI_31_), .ZN(n10276) );
  XNOR2_X1 U8069 ( .A(n6343), .B(n10276), .ZN(n6344) );
  INV_X1 U8070 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6345) );
  NOR2_X1 U8071 ( .A1(n5391), .A2(n6345), .ZN(n6346) );
  AND2_X1 U8072 ( .A1(n9579), .A2(n9190), .ZN(n6483) );
  INV_X1 U8073 ( .A(n9579), .ZN(n6348) );
  AOI211_X1 U8074 ( .C1(n6350), .C2(n6554), .A(n6349), .B(n6549), .ZN(n6381)
         );
  AND2_X1 U8075 ( .A1(n6432), .A2(n6351), .ZN(n6439) );
  INV_X1 U8076 ( .A(n6439), .ZN(n6526) );
  AND2_X1 U8077 ( .A1(n6441), .A2(n6352), .ZN(n6524) );
  INV_X1 U8078 ( .A(n6524), .ZN(n6366) );
  INV_X1 U8079 ( .A(n6353), .ZN(n6503) );
  INV_X1 U8080 ( .A(n6354), .ZN(n7085) );
  INV_X1 U8081 ( .A(n7121), .ZN(n6355) );
  NAND4_X1 U8082 ( .A1(n7085), .A2(n9754), .A3(n6355), .A4(n7223), .ZN(n6357)
         );
  AND2_X1 U8083 ( .A1(n9218), .A2(n7228), .ZN(n6498) );
  NOR2_X1 U8084 ( .A1(n7222), .A2(n6498), .ZN(n7010) );
  INV_X1 U8085 ( .A(n9746), .ZN(n9739) );
  NAND4_X1 U8086 ( .A1(n7010), .A2(n9739), .A3(n6396), .A4(n6840), .ZN(n6356)
         );
  OR2_X1 U8087 ( .A1(n6357), .A2(n6356), .ZN(n6358) );
  NOR2_X1 U8088 ( .A1(n6398), .A2(n6358), .ZN(n6359) );
  NAND4_X1 U8089 ( .A1(n6360), .A2(n6503), .A3(n6359), .A4(n6421), .ZN(n6361)
         );
  NOR3_X1 U8090 ( .A1(n7618), .A2(n7694), .A3(n6361), .ZN(n6362) );
  NAND4_X1 U8091 ( .A1(n9562), .A2(n7730), .A3(n4923), .A4(n6362), .ZN(n6363)
         );
  OR2_X1 U8092 ( .A1(n6364), .A2(n6363), .ZN(n6365) );
  OR3_X1 U8093 ( .A1(n6526), .A2(n6366), .A3(n6365), .ZN(n6367) );
  NOR2_X1 U8094 ( .A1(n9501), .A2(n6367), .ZN(n6368) );
  INV_X1 U8095 ( .A(n9474), .ZN(n9469) );
  AND4_X1 U8096 ( .A1(n9462), .A2(n9487), .A3(n6368), .A4(n9469), .ZN(n6369)
         );
  NAND2_X1 U8097 ( .A1(n9443), .A2(n6369), .ZN(n6370) );
  OR2_X1 U8098 ( .A1(n6370), .A2(n9429), .ZN(n6372) );
  INV_X1 U8099 ( .A(n6458), .ZN(n6464) );
  OR4_X1 U8100 ( .A1(n6372), .A2(n9385), .A3(n9413), .A4(n6371), .ZN(n6373) );
  NOR2_X1 U8101 ( .A1(n6374), .A2(n6373), .ZN(n6376) );
  NAND4_X1 U8102 ( .A1(n6554), .A2(n4899), .A3(n6376), .A4(n6375), .ZN(n6379)
         );
  INV_X1 U8103 ( .A(n6549), .ZN(n6378) );
  NAND2_X1 U8104 ( .A1(n6378), .A2(n6377), .ZN(n6539) );
  OR2_X1 U8105 ( .A1(n6379), .A2(n6539), .ZN(n6486) );
  INV_X1 U8106 ( .A(n6486), .ZN(n6380) );
  NOR2_X1 U8107 ( .A1(n6381), .A2(n6380), .ZN(n6489) );
  INV_X1 U8108 ( .A(n6468), .ZN(n6550) );
  AOI211_X1 U8109 ( .C1(n9649), .C2(n6550), .A(n6480), .B(n9579), .ZN(n6485)
         );
  OR3_X1 U8110 ( .A1(n6382), .A2(n6470), .A3(n6550), .ZN(n6383) );
  NAND2_X1 U8111 ( .A1(n6383), .A2(n5135), .ZN(n6473) );
  MUX2_X1 U8112 ( .A(n6385), .B(n6384), .S(n6550), .Z(n6454) );
  INV_X1 U8113 ( .A(n9628), .ZN(n9510) );
  AOI22_X1 U8114 ( .A1(n9487), .A2(n9510), .B1(n6550), .B2(n6386), .ZN(n6390)
         );
  INV_X1 U8115 ( .A(n6433), .ZN(n6389) );
  NAND3_X1 U8116 ( .A1(n6387), .A2(n9200), .A3(n6468), .ZN(n6388) );
  OAI21_X1 U8117 ( .B1(n6390), .B2(n6389), .A(n6388), .ZN(n6437) );
  NAND2_X1 U8118 ( .A1(n6521), .A2(n4914), .ZN(n6391) );
  AND2_X1 U8119 ( .A1(n6391), .A2(n6522), .ZN(n6420) );
  NAND2_X1 U8120 ( .A1(n6393), .A2(n6392), .ZN(n9740) );
  NAND2_X1 U8121 ( .A1(n9740), .A2(n6500), .ZN(n6395) );
  INV_X1 U8122 ( .A(n7387), .ZN(n7389) );
  NAND4_X1 U8123 ( .A1(n6395), .A2(n7389), .A3(n6396), .A4(n6394), .ZN(n6401)
         );
  OAI21_X1 U8124 ( .B1(n7238), .B2(n6397), .A(n6396), .ZN(n6399) );
  AOI21_X1 U8125 ( .B1(n6399), .B2(n7389), .A(n6398), .ZN(n6400) );
  OAI211_X1 U8126 ( .C1(n7387), .C2(n7385), .A(n7404), .B(n6402), .ZN(n6403)
         );
  NAND2_X1 U8127 ( .A1(n6403), .A2(n6550), .ZN(n6404) );
  INV_X1 U8128 ( .A(n6405), .ZN(n6406) );
  MUX2_X1 U8129 ( .A(n6407), .B(n6406), .S(n6468), .Z(n6408) );
  INV_X1 U8130 ( .A(n6421), .ZN(n6410) );
  NAND2_X1 U8131 ( .A1(n6411), .A2(n7689), .ZN(n6412) );
  NAND3_X1 U8132 ( .A1(n6412), .A2(n7617), .A3(n6508), .ZN(n6413) );
  NAND3_X1 U8133 ( .A1(n6413), .A2(n6423), .A3(n6510), .ZN(n6414) );
  NAND3_X1 U8134 ( .A1(n6414), .A2(n6514), .A3(n6425), .ZN(n6415) );
  INV_X1 U8135 ( .A(n7730), .ZN(n7726) );
  AOI21_X1 U8136 ( .B1(n6415), .B2(n6511), .A(n7726), .ZN(n6418) );
  NAND2_X1 U8137 ( .A1(n6417), .A2(n6416), .ZN(n6493) );
  INV_X1 U8138 ( .A(n6521), .ZN(n6419) );
  NAND2_X1 U8139 ( .A1(n6422), .A2(n6421), .ZN(n6424) );
  NAND2_X1 U8140 ( .A1(n6423), .A2(n7689), .ZN(n6507) );
  AOI21_X1 U8141 ( .B1(n6424), .B2(n6508), .A(n6507), .ZN(n6426) );
  NAND2_X1 U8142 ( .A1(n6425), .A2(n7617), .ZN(n6512) );
  OAI21_X1 U8143 ( .B1(n6426), .B2(n6512), .A(n6510), .ZN(n6428) );
  NAND2_X1 U8144 ( .A1(n7730), .A2(n6511), .ZN(n6427) );
  AOI21_X1 U8145 ( .B1(n6428), .B2(n6514), .A(n6427), .ZN(n6430) );
  NAND4_X1 U8146 ( .A1(n6521), .A2(n6520), .A3(n6515), .A4(n6468), .ZN(n6429)
         );
  INV_X1 U8147 ( .A(n9528), .ZN(n9526) );
  NAND2_X1 U8148 ( .A1(n6431), .A2(n9526), .ZN(n6440) );
  NAND2_X1 U8149 ( .A1(n6440), .A2(n6524), .ZN(n6434) );
  AND2_X1 U8150 ( .A1(n6433), .A2(n6432), .ZN(n6530) );
  NAND3_X1 U8151 ( .A1(n6434), .A2(n6530), .A3(n6468), .ZN(n6435) );
  NAND3_X1 U8152 ( .A1(n6437), .A2(n6436), .A3(n6435), .ZN(n6447) );
  NAND2_X1 U8153 ( .A1(n6438), .A2(n6468), .ZN(n6446) );
  NAND2_X1 U8154 ( .A1(n6440), .A2(n6439), .ZN(n6442) );
  NAND4_X1 U8155 ( .A1(n6442), .A2(n6550), .A3(n6527), .A4(n6441), .ZN(n6444)
         );
  NAND2_X1 U8156 ( .A1(n6444), .A2(n6443), .ZN(n6445) );
  OAI21_X1 U8157 ( .B1(n6448), .B2(n6468), .A(n9462), .ZN(n6449) );
  INV_X1 U8158 ( .A(n9429), .ZN(n6453) );
  MUX2_X1 U8159 ( .A(n6451), .B(n6450), .S(n6468), .Z(n6452) );
  MUX2_X1 U8160 ( .A(n6456), .B(n6455), .S(n6550), .Z(n6457) );
  OAI211_X1 U8161 ( .C1(n6465), .C2(n6461), .A(n6466), .B(n6458), .ZN(n6459)
         );
  NAND2_X1 U8162 ( .A1(n6459), .A2(n6463), .ZN(n6460) );
  NAND2_X1 U8163 ( .A1(n6460), .A2(n6550), .ZN(n6471) );
  INV_X1 U8164 ( .A(n6461), .ZN(n6462) );
  OAI211_X1 U8165 ( .C1(n6465), .C2(n6464), .A(n6463), .B(n6462), .ZN(n6467)
         );
  AND2_X1 U8166 ( .A1(n6467), .A2(n6466), .ZN(n6469) );
  MUX2_X1 U8167 ( .A(n6477), .B(n6476), .S(n6550), .Z(n6478) );
  NAND2_X1 U8168 ( .A1(n6479), .A2(n6478), .ZN(n6484) );
  OAI22_X1 U8169 ( .A1(n9649), .A2(n6550), .B1(n6481), .B2(n6480), .ZN(n6482)
         );
  NAND2_X1 U8170 ( .A1(n6487), .A2(n6486), .ZN(n6488) );
  INV_X1 U8171 ( .A(n6490), .ZN(n6538) );
  INV_X1 U8172 ( .A(n6491), .ZN(n6535) );
  INV_X1 U8173 ( .A(n6492), .ZN(n6533) );
  INV_X1 U8174 ( .A(n6493), .ZN(n6518) );
  INV_X1 U8175 ( .A(n6494), .ZN(n9216) );
  NAND2_X1 U8176 ( .A1(n9216), .A2(n9783), .ZN(n6495) );
  NAND4_X1 U8177 ( .A1(n6497), .A2(n6496), .A3(n6844), .A4(n6495), .ZN(n6502)
         );
  INV_X1 U8178 ( .A(n6498), .ZN(n6499) );
  NOR2_X1 U8179 ( .A1(n6502), .A2(n6501), .ZN(n6504) );
  OAI21_X1 U8180 ( .B1(n7386), .B2(n6504), .A(n6503), .ZN(n6506) );
  NAND2_X1 U8181 ( .A1(n6506), .A2(n6505), .ZN(n6509) );
  AOI21_X1 U8182 ( .B1(n6509), .B2(n6508), .A(n6507), .ZN(n6513) );
  OAI211_X1 U8183 ( .C1(n6513), .C2(n6512), .A(n6511), .B(n6510), .ZN(n6516)
         );
  NAND3_X1 U8184 ( .A1(n6516), .A2(n6515), .A3(n6514), .ZN(n6517) );
  NAND2_X1 U8185 ( .A1(n6518), .A2(n6517), .ZN(n6519) );
  NAND3_X1 U8186 ( .A1(n6521), .A2(n6520), .A3(n6519), .ZN(n6523) );
  AND2_X1 U8187 ( .A1(n6523), .A2(n6522), .ZN(n6525) );
  OAI21_X1 U8188 ( .B1(n6526), .B2(n6525), .A(n6524), .ZN(n6529) );
  INV_X1 U8189 ( .A(n6527), .ZN(n6528) );
  AOI21_X1 U8190 ( .B1(n6530), .B2(n6529), .A(n6528), .ZN(n6531) );
  OR3_X1 U8191 ( .A1(n6533), .A2(n6532), .A3(n6531), .ZN(n6534) );
  NAND2_X1 U8192 ( .A1(n6535), .A2(n6534), .ZN(n6537) );
  AOI21_X1 U8193 ( .B1(n6538), .B2(n6537), .A(n6536), .ZN(n6540) );
  OR2_X1 U8194 ( .A1(n6540), .A2(n6539), .ZN(n6541) );
  NAND2_X1 U8195 ( .A1(n6541), .A2(n6554), .ZN(n6543) );
  OR2_X1 U8196 ( .A1(n6876), .A2(P1_U3086), .ZN(n7721) );
  AOI21_X1 U8197 ( .B1(n6543), .B2(n6845), .A(n7721), .ZN(n6544) );
  AOI21_X1 U8198 ( .B1(n6550), .B2(n6549), .A(n4577), .ZN(n6561) );
  NOR2_X1 U8199 ( .A1(n7721), .A2(n6551), .ZN(n6556) );
  INV_X1 U8200 ( .A(n6552), .ZN(n6553) );
  OAI211_X1 U8201 ( .C1(n6554), .C2(n5711), .A(n6556), .B(n6553), .ZN(n6560)
         );
  INV_X1 U8202 ( .A(n9684), .ZN(n6751) );
  INV_X1 U8203 ( .A(n6555), .ZN(n6843) );
  NAND3_X1 U8204 ( .A1(n9181), .A2(n6751), .A3(n6843), .ZN(n6558) );
  INV_X1 U8205 ( .A(n6556), .ZN(n6557) );
  OAI211_X1 U8206 ( .C1(n6558), .C2(n9775), .A(P1_B_REG_SCAN_IN), .B(n6557), 
        .ZN(n6559) );
  INV_X1 U8207 ( .A(n6565), .ZN(n6568) );
  INV_X1 U8208 ( .A(n6566), .ZN(n6567) );
  NAND2_X1 U8209 ( .A1(n6568), .A2(n6567), .ZN(n6571) );
  INV_X1 U8210 ( .A(n6650), .ZN(n6569) );
  NOR2_X1 U8211 ( .A1(n7275), .A2(n6569), .ZN(n6570) );
  OR2_X2 U8212 ( .A1(n6573), .A2(n6572), .ZN(n6577) );
  NAND2_X1 U8213 ( .A1(n6573), .A2(n6572), .ZN(n6574) );
  OR2_X1 U8214 ( .A1(n6582), .A2(n6575), .ZN(n6576) );
  NAND2_X1 U8215 ( .A1(n7048), .A2(n6576), .ZN(n7139) );
  NAND2_X1 U8216 ( .A1(n7137), .A2(n7139), .ZN(n7138) );
  NAND2_X1 U8217 ( .A1(n7138), .A2(n6577), .ZN(n7144) );
  INV_X1 U8218 ( .A(n8207), .ZN(n6579) );
  XNOR2_X1 U8219 ( .A(n6580), .B(n6579), .ZN(n7145) );
  NAND2_X1 U8220 ( .A1(n7144), .A2(n7145), .ZN(n7143) );
  OR2_X1 U8221 ( .A1(n6580), .A2(n8207), .ZN(n6581) );
  NAND2_X1 U8222 ( .A1(n7143), .A2(n6581), .ZN(n7300) );
  INV_X1 U8223 ( .A(n7300), .ZN(n6584) );
  XNOR2_X1 U8224 ( .A(n7997), .B(n10033), .ZN(n6586) );
  INV_X1 U8225 ( .A(n4507), .ZN(n6585) );
  XNOR2_X1 U8226 ( .A(n6586), .B(n6585), .ZN(n7301) );
  INV_X1 U8227 ( .A(n7301), .ZN(n6583) );
  OR2_X1 U8228 ( .A1(n6586), .A2(n6585), .ZN(n6587) );
  XNOR2_X1 U8229 ( .A(n7997), .B(n10039), .ZN(n6588) );
  INV_X1 U8230 ( .A(n8212), .ZN(n7297) );
  NAND2_X1 U8231 ( .A1(n6588), .A2(n7297), .ZN(n7454) );
  OR2_X1 U8232 ( .A1(n6588), .A2(n7297), .ZN(n6589) );
  AND2_X1 U8233 ( .A1(n6589), .A2(n7454), .ZN(n7307) );
  INV_X1 U8234 ( .A(n6590), .ZN(n6638) );
  XNOR2_X1 U8235 ( .A(n6638), .B(n8217), .ZN(n6592) );
  XNOR2_X1 U8236 ( .A(n6592), .B(n8527), .ZN(n7453) );
  NAND2_X1 U8237 ( .A1(n6592), .A2(n8218), .ZN(n6593) );
  XNOR2_X1 U8238 ( .A(n6638), .B(n10047), .ZN(n6595) );
  INV_X1 U8239 ( .A(n8526), .ZN(n7452) );
  XNOR2_X1 U8240 ( .A(n6595), .B(n7452), .ZN(n7607) );
  OR2_X1 U8241 ( .A1(n6595), .A2(n7452), .ZN(n6596) );
  XNOR2_X1 U8242 ( .A(n7997), .B(n7663), .ZN(n6597) );
  INV_X1 U8243 ( .A(n8525), .ZN(n7603) );
  NAND2_X1 U8244 ( .A1(n6597), .A2(n7603), .ZN(n7667) );
  OR2_X1 U8245 ( .A1(n6597), .A2(n7603), .ZN(n6598) );
  AND2_X1 U8246 ( .A1(n7667), .A2(n6598), .ZN(n7630) );
  NAND2_X1 U8247 ( .A1(n7629), .A2(n7667), .ZN(n6599) );
  XNOR2_X1 U8248 ( .A(n10057), .B(n6590), .ZN(n6600) );
  XNOR2_X1 U8249 ( .A(n6600), .B(n8524), .ZN(n7668) );
  NAND2_X1 U8250 ( .A1(n6600), .A2(n4862), .ZN(n6601) );
  XNOR2_X1 U8251 ( .A(n10065), .B(n6638), .ZN(n6603) );
  XNOR2_X1 U8252 ( .A(n6603), .B(n7676), .ZN(n7851) );
  INV_X1 U8253 ( .A(n7851), .ZN(n6602) );
  INV_X1 U8254 ( .A(n6603), .ZN(n6604) );
  NAND2_X1 U8255 ( .A1(n6604), .A2(n8523), .ZN(n6605) );
  XOR2_X1 U8256 ( .A(n6638), .B(n10071), .Z(n7929) );
  NOR2_X1 U8257 ( .A1(n6606), .A2(n8522), .ZN(n8469) );
  XNOR2_X1 U8258 ( .A(n8176), .B(n6590), .ZN(n8468) );
  AND2_X1 U8259 ( .A1(n8468), .A2(n8805), .ZN(n6607) );
  XNOR2_X1 U8260 ( .A(n8996), .B(n6638), .ZN(n6608) );
  XNOR2_X1 U8261 ( .A(n6608), .B(n8453), .ZN(n8402) );
  XNOR2_X1 U8262 ( .A(n8990), .B(n7997), .ZN(n6610) );
  NOR2_X1 U8263 ( .A1(n6610), .A2(n6609), .ZN(n8450) );
  XNOR2_X1 U8264 ( .A(n8984), .B(n6638), .ZN(n6611) );
  XNOR2_X1 U8265 ( .A(n6611), .B(n8787), .ZN(n8372) );
  XNOR2_X1 U8266 ( .A(n8978), .B(n7997), .ZN(n6613) );
  XNOR2_X1 U8267 ( .A(n6613), .B(n8774), .ZN(n8507) );
  NAND2_X1 U8268 ( .A1(n8508), .A2(n8507), .ZN(n8506) );
  NAND2_X1 U8269 ( .A1(n8506), .A2(n6614), .ZN(n8420) );
  XNOR2_X1 U8270 ( .A(n8887), .B(n6638), .ZN(n6615) );
  XNOR2_X1 U8271 ( .A(n6615), .B(n8766), .ZN(n8419) );
  XNOR2_X1 U8272 ( .A(n8968), .B(n7997), .ZN(n6617) );
  XNOR2_X1 U8273 ( .A(n6617), .B(n8756), .ZN(n8428) );
  INV_X1 U8274 ( .A(n6617), .ZN(n6618) );
  NOR2_X1 U8275 ( .A1(n6618), .A2(n8521), .ZN(n8486) );
  XNOR2_X1 U8276 ( .A(n8483), .B(n7997), .ZN(n6619) );
  XNOR2_X1 U8277 ( .A(n6619), .B(n8744), .ZN(n8485) );
  XNOR2_X1 U8278 ( .A(n8391), .B(n7997), .ZN(n6621) );
  XNOR2_X1 U8279 ( .A(n6621), .B(n8719), .ZN(n8386) );
  NAND2_X1 U8280 ( .A1(n8385), .A2(n8386), .ZN(n6623) );
  NAND2_X1 U8281 ( .A1(n6621), .A2(n8729), .ZN(n6622) );
  XOR2_X1 U8282 ( .A(n7997), .B(n8874), .Z(n6625) );
  INV_X1 U8283 ( .A(n6625), .ZN(n6624) );
  XNOR2_X1 U8284 ( .A(n6624), .B(n8705), .ZN(n8444) );
  XNOR2_X1 U8285 ( .A(n8953), .B(n7997), .ZN(n6626) );
  XNOR2_X1 U8286 ( .A(n6626), .B(n8691), .ZN(n8394) );
  NAND2_X1 U8287 ( .A1(n6626), .A2(n8691), .ZN(n6627) );
  XOR2_X1 U8288 ( .A(n7997), .B(n8695), .Z(n6629) );
  INV_X1 U8289 ( .A(n6629), .ZN(n6628) );
  XNOR2_X1 U8290 ( .A(n6628), .B(n8704), .ZN(n8461) );
  XNOR2_X1 U8291 ( .A(n8943), .B(n6638), .ZN(n6631) );
  NAND2_X1 U8292 ( .A1(n8379), .A2(n8692), .ZN(n6634) );
  INV_X1 U8293 ( .A(n6630), .ZN(n6632) );
  NAND2_X1 U8294 ( .A1(n6632), .A2(n6631), .ZN(n6633) );
  NAND2_X1 U8295 ( .A1(n6634), .A2(n6633), .ZN(n8436) );
  XNOR2_X1 U8296 ( .A(n8937), .B(n6638), .ZN(n6635) );
  NAND2_X1 U8297 ( .A1(n8436), .A2(n8437), .ZN(n6637) );
  NAND2_X1 U8298 ( .A1(n6635), .A2(n8414), .ZN(n6636) );
  XNOR2_X1 U8299 ( .A(n8931), .B(n6638), .ZN(n6639) );
  XNOR2_X1 U8300 ( .A(n6639), .B(n8671), .ZN(n8411) );
  NAND2_X1 U8301 ( .A1(n6639), .A2(n8647), .ZN(n6640) );
  XNOR2_X1 U8302 ( .A(n6641), .B(n7997), .ZN(n6642) );
  NAND2_X1 U8303 ( .A1(n6642), .A2(n8658), .ZN(n8494) );
  INV_X1 U8304 ( .A(n6642), .ZN(n6643) );
  NAND2_X1 U8305 ( .A1(n6643), .A2(n6666), .ZN(n8495) );
  XNOR2_X1 U8306 ( .A(n8919), .B(n7997), .ZN(n7993) );
  XNOR2_X1 U8307 ( .A(n7996), .B(n7995), .ZN(n6671) );
  INV_X1 U8308 ( .A(n6644), .ZN(n6645) );
  NAND2_X1 U8309 ( .A1(n6648), .A2(n6645), .ZN(n6646) );
  NAND2_X1 U8310 ( .A1(n6648), .A2(n10063), .ZN(n6649) );
  AND2_X1 U8311 ( .A1(n10076), .A2(n8161), .ZN(n7069) );
  NAND2_X1 U8312 ( .A1(n8919), .A2(n8501), .ZN(n6670) );
  INV_X1 U8313 ( .A(n6651), .ZN(n6653) );
  NAND2_X1 U8314 ( .A1(n8336), .A2(n6650), .ZN(n7066) );
  OAI211_X1 U8315 ( .C1(n7068), .C2(n6651), .A(n6679), .B(n7066), .ZN(n6652)
         );
  AOI21_X1 U8316 ( .B1(n7070), .B2(n6653), .A(n6652), .ZN(n6654) );
  OAI21_X1 U8317 ( .B1(n6658), .B2(n6655), .A(n6654), .ZN(n6656) );
  NAND2_X1 U8318 ( .A1(n6656), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6660) );
  NAND2_X1 U8319 ( .A1(n7067), .A2(n6657), .ZN(n8347) );
  OR2_X1 U8320 ( .A1(n6658), .A2(n8347), .ZN(n6659) );
  AND2_X1 U8321 ( .A1(n6660), .A2(n6659), .ZN(n7132) );
  OR2_X1 U8322 ( .A1(n6680), .A2(P2_U3151), .ZN(n8351) );
  OR2_X1 U8323 ( .A1(n6661), .A2(n7208), .ZN(n6665) );
  OAI22_X1 U8324 ( .A1(n8510), .A2(n6209), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6663), .ZN(n6668) );
  OR2_X1 U8325 ( .A1(n6665), .A2(n6664), .ZN(n8476) );
  NOR2_X1 U8326 ( .A1(n6666), .A2(n8476), .ZN(n6667) );
  AOI211_X1 U8327 ( .C1(n8639), .C2(n8497), .A(n6668), .B(n6667), .ZN(n6669)
         );
  OAI21_X1 U8328 ( .B1(n6671), .B2(n8503), .A(n5134), .ZN(P2_U3154) );
  INV_X1 U8329 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6672) );
  NOR2_X1 U8330 ( .A1(n9858), .A2(n6672), .ZN(n6673) );
  AOI21_X1 U8331 ( .B1(n6348), .B2(n5784), .A(n6673), .ZN(n6676) );
  AND2_X1 U8332 ( .A1(n9190), .A2(n6674), .ZN(n9353) );
  OR2_X1 U8333 ( .A1(n9576), .A2(n5809), .ZN(n6675) );
  NAND2_X1 U8334 ( .A1(n6676), .A2(n6675), .ZN(P1_U3521) );
  NOR2_X1 U8335 ( .A1(n6875), .A2(P1_U3086), .ZN(n6677) );
  INV_X1 U8336 ( .A(n6680), .ZN(n6678) );
  NAND2_X1 U8337 ( .A1(n8336), .A2(n6680), .ZN(n6681) );
  NAND2_X1 U8338 ( .A1(n6934), .A2(n6681), .ZN(n6956) );
  OR2_X1 U8339 ( .A1(n6956), .A2(n6682), .ZN(n6683) );
  NAND2_X1 U8340 ( .A1(n6683), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NAND2_X1 U8341 ( .A1(n4511), .A2(P1_U3086), .ZN(n9689) );
  AND2_X1 U8342 ( .A1(n4514), .A2(P1_U3086), .ZN(n9679) );
  INV_X2 U8343 ( .A(n9679), .ZN(n9687) );
  OAI222_X1 U8344 ( .A1(P1_U3086), .A2(n9270), .B1(n9689), .B2(n6689), .C1(
        n9687), .C2(n5357), .ZN(P1_U3351) );
  OAI222_X1 U8345 ( .A1(P1_U3086), .A2(n9251), .B1(n9689), .B2(n6686), .C1(
        n6684), .C2(n9687), .ZN(P1_U3352) );
  OAI222_X1 U8346 ( .A1(P1_U3086), .A2(n6753), .B1(n9689), .B2(n6690), .C1(
        n9687), .C2(n5316), .ZN(P1_U3353) );
  INV_X2 U8347 ( .A(n9010), .ZN(n9018) );
  NOR2_X1 U8348 ( .A1(n4513), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9005) );
  OAI222_X1 U8349 ( .A1(n9018), .A2(n6686), .B1(n6968), .B2(P2_U3151), .C1(
        n6685), .C2(n9015), .ZN(P2_U3292) );
  OAI222_X1 U8350 ( .A1(n9018), .A2(n6688), .B1(n9892), .B2(P2_U3151), .C1(
        n6687), .C2(n9015), .ZN(P2_U3294) );
  OAI222_X1 U8351 ( .A1(n9015), .A2(n4611), .B1(n9018), .B2(n6689), .C1(
        P2_U3151), .C2(n7035), .ZN(P2_U3291) );
  OAI222_X1 U8352 ( .A1(n9015), .A2(n6691), .B1(n9018), .B2(n6690), .C1(
        P2_U3151), .C2(n6966), .ZN(P2_U3293) );
  OAI222_X1 U8353 ( .A1(n9018), .A2(n6693), .B1(n7182), .B2(P2_U3151), .C1(
        n6692), .C2(n9015), .ZN(P2_U3290) );
  OAI222_X1 U8354 ( .A1(n9687), .A2(n6694), .B1(n9689), .B2(n6693), .C1(n6774), 
        .C2(P1_U3086), .ZN(P1_U3350) );
  OAI222_X1 U8355 ( .A1(n9018), .A2(n6696), .B1(n7464), .B2(P2_U3151), .C1(
        n6695), .C2(n9015), .ZN(P2_U3289) );
  INV_X1 U8356 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6697) );
  INV_X1 U8357 ( .A(n6792), .ZN(n6786) );
  OAI222_X1 U8358 ( .A1(n9687), .A2(n6697), .B1(n9689), .B2(n6696), .C1(n6786), 
        .C2(P1_U3086), .ZN(P1_U3349) );
  OAI222_X1 U8359 ( .A1(n9018), .A2(n6699), .B1(n7475), .B2(P2_U3151), .C1(
        n6698), .C2(n9015), .ZN(P2_U3288) );
  INV_X1 U8360 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10328) );
  INV_X1 U8361 ( .A(n9689), .ZN(n7720) );
  INV_X1 U8362 ( .A(n6793), .ZN(n6828) );
  OAI222_X1 U8363 ( .A1(n9687), .A2(n10328), .B1(n9686), .B2(n6699), .C1(n6828), .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U8364 ( .A(n9775), .ZN(n6870) );
  INV_X1 U8365 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6701) );
  OAI21_X1 U8366 ( .B1(n6870), .B2(n6701), .A(n6700), .ZN(P1_U3439) );
  INV_X1 U8367 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6704) );
  INV_X1 U8368 ( .A(n6866), .ZN(n6702) );
  NAND2_X1 U8369 ( .A1(n6870), .A2(n6702), .ZN(n6703) );
  OAI21_X1 U8370 ( .B1(n6870), .B2(n6704), .A(n6703), .ZN(P1_U3440) );
  INV_X1 U8371 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6706) );
  INV_X1 U8372 ( .A(n6705), .ZN(n6707) );
  OAI222_X1 U8373 ( .A1(n9015), .A2(n6706), .B1(n9018), .B2(n6707), .C1(
        P2_U3151), .C2(n7750), .ZN(P2_U3287) );
  INV_X1 U8374 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10440) );
  INV_X1 U8375 ( .A(n6795), .ZN(n6807) );
  OAI222_X1 U8376 ( .A1(n9687), .A2(n10440), .B1(n9689), .B2(n6707), .C1(
        P1_U3086), .C2(n6807), .ZN(P1_U3347) );
  INV_X1 U8377 ( .A(n6875), .ZN(n6852) );
  NAND2_X1 U8378 ( .A1(n6876), .A2(n6852), .ZN(n6708) );
  NAND2_X1 U8379 ( .A1(n6708), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6712) );
  INV_X1 U8380 ( .A(n6712), .ZN(n6711) );
  NAND2_X1 U8381 ( .A1(n6872), .A2(n6876), .ZN(n6710) );
  NAND2_X1 U8382 ( .A1(n6710), .A2(n6709), .ZN(n6713) );
  NAND2_X1 U8383 ( .A1(n6711), .A2(n6713), .ZN(n9263) );
  INV_X1 U8384 ( .A(n9263), .ZN(n9349) );
  NOR2_X1 U8385 ( .A1(n9349), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8386 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6719) );
  INV_X1 U8387 ( .A(n6752), .ZN(n6717) );
  INV_X1 U8388 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7014) );
  NAND2_X1 U8389 ( .A1(n6751), .A2(n7014), .ZN(n6714) );
  AND2_X1 U8390 ( .A1(n9232), .A2(n6714), .ZN(n9235) );
  OAI21_X1 U8391 ( .B1(n6751), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9235), .ZN(
        n6715) );
  XNOR2_X1 U8392 ( .A(n6715), .B(P1_IR_REG_0__SCAN_IN), .ZN(n6716) );
  AOI22_X1 U8393 ( .A1(n6717), .A2(n6716), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n6718) );
  OAI21_X1 U8394 ( .B1(n9263), .B2(n6719), .A(n6718), .ZN(P1_U3243) );
  INV_X1 U8395 ( .A(n6720), .ZN(n6723) );
  INV_X1 U8396 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6721) );
  OAI222_X1 U8397 ( .A1(n9018), .A2(n6723), .B1(n4983), .B2(P2_U3151), .C1(
        n6721), .C2(n9015), .ZN(P2_U3286) );
  INV_X1 U8398 ( .A(n7949), .ZN(n7915) );
  INV_X1 U8399 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6722) );
  OAI222_X1 U8400 ( .A1(n9018), .A2(n6725), .B1(n7915), .B2(P2_U3151), .C1(
        n6722), .C2(n9015), .ZN(P2_U3285) );
  INV_X1 U8401 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6724) );
  INV_X1 U8402 ( .A(n6892), .ZN(n6898) );
  OAI222_X1 U8403 ( .A1(n9687), .A2(n6724), .B1(n9689), .B2(n6723), .C1(n6898), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U8404 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10236) );
  INV_X1 U8405 ( .A(n7019), .ZN(n6904) );
  OAI222_X1 U8406 ( .A1(n9687), .A2(n10236), .B1(n9689), .B2(n6725), .C1(n6904), .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U8407 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6728) );
  INV_X1 U8408 ( .A(n7062), .ZN(n6726) );
  NAND2_X1 U8409 ( .A1(n6726), .A2(n7067), .ZN(n6727) );
  OAI21_X1 U8410 ( .B1(n7067), .B2(n6728), .A(n6727), .ZN(P2_U3377) );
  INV_X1 U8411 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6835) );
  NAND2_X1 U8412 ( .A1(n6729), .A2(P1_U3973), .ZN(n6730) );
  OAI21_X1 U8413 ( .B1(n6835), .B2(P1_U3973), .A(n6730), .ZN(P1_U3567) );
  AND2_X1 U8414 ( .A1(n6735), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8415 ( .A1(n6735), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8416 ( .A1(n6735), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8417 ( .A1(n6735), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8418 ( .A1(n6735), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8419 ( .A1(n6735), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8420 ( .A1(n6735), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8421 ( .A1(n6735), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8422 ( .A1(n6735), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8423 ( .A1(n6735), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8424 ( .A1(n6735), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8425 ( .A1(n6735), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8426 ( .A1(n6735), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8427 ( .A1(n6735), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8428 ( .A1(n6735), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8429 ( .A1(n6735), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8430 ( .A1(n6735), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8431 ( .A1(n6735), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8432 ( .A1(n6735), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8433 ( .A1(n6735), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8434 ( .A1(n6735), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8435 ( .A1(n6735), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8436 ( .A1(n6735), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8437 ( .A1(n6735), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8438 ( .A1(n6735), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8439 ( .A1(n6735), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8440 ( .A1(n6735), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8441 ( .A1(n6735), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8442 ( .A1(n6735), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8443 ( .A1(n6735), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  INV_X1 U8444 ( .A(n6732), .ZN(n6733) );
  AOI22_X1 U8445 ( .A1(n6735), .A2(n6734), .B1(n6733), .B2(n7131), .ZN(
        P2_U3376) );
  INV_X1 U8446 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6737) );
  INV_X1 U8447 ( .A(n6736), .ZN(n6738) );
  OAI222_X1 U8448 ( .A1(n9015), .A2(n6737), .B1(n9018), .B2(n6738), .C1(
        P2_U3151), .C2(n7917), .ZN(P2_U3284) );
  INV_X1 U8449 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10331) );
  INV_X1 U8450 ( .A(n7109), .ZN(n7028) );
  OAI222_X1 U8451 ( .A1(n9687), .A2(n10331), .B1(n9689), .B2(n6738), .C1(
        P1_U3086), .C2(n7028), .ZN(P1_U3344) );
  INV_X1 U8452 ( .A(n8570), .ZN(n8531) );
  INV_X1 U8453 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6739) );
  OAI222_X1 U8454 ( .A1(n9018), .A2(n6741), .B1(n8531), .B2(P2_U3151), .C1(
        n6739), .C2(n9015), .ZN(P2_U3283) );
  INV_X1 U8455 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6740) );
  OAI222_X1 U8456 ( .A1(P1_U3086), .A2(n7116), .B1(n9689), .B2(n6741), .C1(
        n6740), .C2(n9687), .ZN(P1_U3343) );
  OR2_X1 U8457 ( .A1(n6752), .A2(n9232), .ZN(n9337) );
  NAND2_X1 U8458 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7264) );
  NAND2_X1 U8459 ( .A1(n9349), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n6742) );
  OAI211_X1 U8460 ( .C1(n9337), .C2(n6774), .A(n7264), .B(n6742), .ZN(n6769)
         );
  INV_X1 U8461 ( .A(n9270), .ZN(n9266) );
  INV_X1 U8462 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7124) );
  MUX2_X1 U8463 ( .A(n7124), .B(P1_REG2_REG_2__SCAN_IN), .S(n6753), .Z(n9244)
         );
  INV_X1 U8464 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7229) );
  MUX2_X1 U8465 ( .A(n7229), .B(P1_REG2_REG_1__SCAN_IN), .S(n6756), .Z(n9223)
         );
  AND2_X1 U8466 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9231) );
  NAND2_X1 U8467 ( .A1(n9223), .A2(n9231), .ZN(n9222) );
  INV_X1 U8468 ( .A(n6756), .ZN(n9221) );
  NAND2_X1 U8469 ( .A1(n9221), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6743) );
  NAND2_X1 U8470 ( .A1(n9222), .A2(n6743), .ZN(n9243) );
  NAND2_X1 U8471 ( .A1(n9244), .A2(n9243), .ZN(n9242) );
  INV_X1 U8472 ( .A(n6753), .ZN(n9239) );
  NAND2_X1 U8473 ( .A1(n9239), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6744) );
  NAND2_X1 U8474 ( .A1(n9242), .A2(n6744), .ZN(n9249) );
  XNOR2_X1 U8475 ( .A(n9251), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9250) );
  NAND2_X1 U8476 ( .A1(n9249), .A2(n9250), .ZN(n9248) );
  INV_X1 U8477 ( .A(n9251), .ZN(n9256) );
  NAND2_X1 U8478 ( .A1(n9256), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6745) );
  NAND2_X1 U8479 ( .A1(n9248), .A2(n6745), .ZN(n9268) );
  INV_X1 U8480 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6746) );
  MUX2_X1 U8481 ( .A(n6746), .B(P1_REG2_REG_4__SCAN_IN), .S(n9270), .Z(n9269)
         );
  NAND2_X1 U8482 ( .A1(n9268), .A2(n9269), .ZN(n9267) );
  INV_X1 U8483 ( .A(n9267), .ZN(n6747) );
  XOR2_X1 U8484 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n6774), .Z(n6749) );
  NOR2_X1 U8485 ( .A1(n6750), .A2(n6749), .ZN(n6770) );
  OR2_X1 U8486 ( .A1(n7973), .A2(n9684), .ZN(n6748) );
  AOI211_X1 U8487 ( .C1(n6750), .C2(n6749), .A(n6770), .B(n9341), .ZN(n6768)
         );
  INV_X1 U8488 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6754) );
  MUX2_X1 U8489 ( .A(n6754), .B(P1_REG1_REG_2__SCAN_IN), .S(n6753), .Z(n9241)
         );
  INV_X1 U8490 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6755) );
  MUX2_X1 U8491 ( .A(n6755), .B(P1_REG1_REG_1__SCAN_IN), .S(n6756), .Z(n9225)
         );
  AND2_X1 U8492 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9226) );
  NAND2_X1 U8493 ( .A1(n9225), .A2(n9226), .ZN(n9224) );
  OR2_X1 U8494 ( .A1(n6756), .A2(n6755), .ZN(n6757) );
  NAND2_X1 U8495 ( .A1(n9224), .A2(n6757), .ZN(n9240) );
  NAND2_X1 U8496 ( .A1(n9241), .A2(n9240), .ZN(n9253) );
  NAND2_X1 U8497 ( .A1(n9239), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9252) );
  NAND2_X1 U8498 ( .A1(n9253), .A2(n9252), .ZN(n6760) );
  INV_X1 U8499 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6758) );
  MUX2_X1 U8500 ( .A(n6758), .B(P1_REG1_REG_3__SCAN_IN), .S(n9251), .Z(n6759)
         );
  NAND2_X1 U8501 ( .A1(n6760), .A2(n6759), .ZN(n9273) );
  NAND2_X1 U8502 ( .A1(n9256), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9272) );
  NAND2_X1 U8503 ( .A1(n9273), .A2(n9272), .ZN(n6763) );
  INV_X1 U8504 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6761) );
  MUX2_X1 U8505 ( .A(n6761), .B(P1_REG1_REG_4__SCAN_IN), .S(n9270), .Z(n6762)
         );
  NAND2_X1 U8506 ( .A1(n6763), .A2(n6762), .ZN(n9274) );
  NAND2_X1 U8507 ( .A1(n9266), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6765) );
  INV_X1 U8508 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9863) );
  MUX2_X1 U8509 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9863), .S(n6774), .Z(n6764)
         );
  AOI21_X1 U8510 ( .B1(n9274), .B2(n6765), .A(n6764), .ZN(n6778) );
  AND3_X1 U8511 ( .A1(n9274), .A2(n6765), .A3(n6764), .ZN(n6766) );
  NOR3_X1 U8512 ( .A1(n9339), .A2(n6778), .A3(n6766), .ZN(n6767) );
  OR3_X1 U8513 ( .A1(n6769), .A2(n6768), .A3(n6767), .ZN(P1_U3248) );
  INV_X1 U8514 ( .A(n6774), .ZN(n6771) );
  AOI21_X1 U8515 ( .B1(n6771), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6770), .ZN(
        n6773) );
  XNOR2_X1 U8516 ( .A(n6792), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n6772) );
  NOR2_X1 U8517 ( .A1(n6773), .A2(n6772), .ZN(n6791) );
  AOI211_X1 U8518 ( .C1(n6773), .C2(n6772), .A(n6791), .B(n9341), .ZN(n6782)
         );
  NOR2_X1 U8519 ( .A1(n6774), .A2(n9863), .ZN(n6777) );
  INV_X1 U8520 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6775) );
  MUX2_X1 U8521 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6775), .S(n6792), .Z(n6776)
         );
  OAI21_X1 U8522 ( .B1(n6778), .B2(n6777), .A(n6776), .ZN(n6820) );
  INV_X1 U8523 ( .A(n6820), .ZN(n6780) );
  NOR3_X1 U8524 ( .A1(n6778), .A2(n6777), .A3(n6776), .ZN(n6779) );
  NOR3_X1 U8525 ( .A1(n9339), .A2(n6780), .A3(n6779), .ZN(n6781) );
  NOR2_X1 U8526 ( .A1(n6782), .A2(n6781), .ZN(n6785) );
  AND2_X1 U8527 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6783) );
  AOI21_X1 U8528 ( .B1(n9349), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n6783), .ZN(
        n6784) );
  OAI211_X1 U8529 ( .C1(n6786), .C2(n9337), .A(n6785), .B(n6784), .ZN(P1_U3249) );
  NAND2_X1 U8530 ( .A1(n6795), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6788) );
  NAND2_X1 U8531 ( .A1(n6792), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6819) );
  INV_X1 U8532 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9866) );
  MUX2_X1 U8533 ( .A(n9866), .B(P1_REG1_REG_7__SCAN_IN), .S(n6793), .Z(n6818)
         );
  AOI21_X1 U8534 ( .B1(n6820), .B2(n6819), .A(n6818), .ZN(n6822) );
  AOI21_X1 U8535 ( .B1(n6793), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6822), .ZN(
        n6804) );
  INV_X1 U8536 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9868) );
  MUX2_X1 U8537 ( .A(n9868), .B(P1_REG1_REG_8__SCAN_IN), .S(n6795), .Z(n6805)
         );
  OR2_X1 U8538 ( .A1(n6804), .A2(n6805), .ZN(n6787) );
  NAND2_X1 U8539 ( .A1(n6788), .A2(n6787), .ZN(n6790) );
  INV_X1 U8540 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6897) );
  MUX2_X1 U8541 ( .A(n6897), .B(P1_REG1_REG_9__SCAN_IN), .S(n6892), .Z(n6789)
         );
  NOR2_X1 U8542 ( .A1(n6790), .A2(n6789), .ZN(n6896) );
  AOI21_X1 U8543 ( .B1(n6790), .B2(n6789), .A(n6896), .ZN(n6803) );
  XOR2_X1 U8544 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n6892), .Z(n6797) );
  XNOR2_X1 U8545 ( .A(n6793), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n6816) );
  NOR2_X1 U8546 ( .A1(n6817), .A2(n6816), .ZN(n6815) );
  AOI21_X1 U8547 ( .B1(n6793), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6815), .ZN(
        n6810) );
  NAND2_X1 U8548 ( .A1(n6795), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6794) );
  OAI21_X1 U8549 ( .B1(n6795), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6794), .ZN(
        n6809) );
  NOR2_X1 U8550 ( .A1(n6810), .A2(n6809), .ZN(n6808) );
  NAND2_X1 U8551 ( .A1(n6796), .A2(n6797), .ZN(n6891) );
  OAI21_X1 U8552 ( .B1(n6797), .B2(n6796), .A(n6891), .ZN(n6798) );
  NAND2_X1 U8553 ( .A1(n6798), .A2(n9319), .ZN(n6802) );
  NOR2_X1 U8554 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6799), .ZN(n7584) );
  NOR2_X1 U8555 ( .A1(n9337), .A2(n6898), .ZN(n6800) );
  AOI211_X1 U8556 ( .C1(n9349), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n7584), .B(
        n6800), .ZN(n6801) );
  OAI211_X1 U8557 ( .C1(n6803), .C2(n9339), .A(n6802), .B(n6801), .ZN(P1_U3252) );
  INV_X1 U8558 ( .A(n9339), .ZN(n9309) );
  XOR2_X1 U8559 ( .A(n6805), .B(n6804), .Z(n6813) );
  AND2_X1 U8560 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9718) );
  AOI21_X1 U8561 ( .B1(n9349), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n9718), .ZN(
        n6806) );
  OAI21_X1 U8562 ( .B1(n6807), .B2(n9337), .A(n6806), .ZN(n6812) );
  AOI211_X1 U8563 ( .C1(n6810), .C2(n6809), .A(n9341), .B(n6808), .ZN(n6811)
         );
  AOI211_X1 U8564 ( .C1(n9309), .C2(n6813), .A(n6812), .B(n6811), .ZN(n6814)
         );
  INV_X1 U8565 ( .A(n6814), .ZN(P1_U3251) );
  AOI211_X1 U8566 ( .C1(n6817), .C2(n6816), .A(n9341), .B(n6815), .ZN(n6824)
         );
  AND3_X1 U8567 ( .A1(n6820), .A2(n6819), .A3(n6818), .ZN(n6821) );
  NOR3_X1 U8568 ( .A1(n9339), .A2(n6822), .A3(n6821), .ZN(n6823) );
  NOR2_X1 U8569 ( .A1(n6824), .A2(n6823), .ZN(n6827) );
  NAND2_X1 U8570 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n7348) );
  INV_X1 U8571 ( .A(n7348), .ZN(n6825) );
  AOI21_X1 U8572 ( .B1(n9349), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n6825), .ZN(
        n6826) );
  OAI211_X1 U8573 ( .C1(n6828), .C2(n9337), .A(n6827), .B(n6826), .ZN(P1_U3250) );
  NAND2_X1 U8574 ( .A1(n8826), .A2(P2_U3893), .ZN(n6829) );
  OAI21_X1 U8575 ( .B1(P2_U3893), .B2(n5295), .A(n6829), .ZN(P2_U3492) );
  NAND2_X1 U8576 ( .A1(n6830), .A2(P2_U3893), .ZN(n6831) );
  OAI21_X1 U8577 ( .B1(P2_U3893), .B2(n5309), .A(n6831), .ZN(P2_U3491) );
  NAND2_X1 U8578 ( .A1(n8212), .A2(P2_U3893), .ZN(n6832) );
  OAI21_X1 U8579 ( .B1(P2_U3893), .B2(n5357), .A(n6832), .ZN(P2_U3495) );
  NAND2_X1 U8580 ( .A1(n8207), .A2(P2_U3893), .ZN(n6833) );
  OAI21_X1 U8581 ( .B1(P2_U3893), .B2(n5316), .A(n6833), .ZN(P2_U3493) );
  INV_X1 U8582 ( .A(n9942), .ZN(n8571) );
  INV_X1 U8583 ( .A(n6834), .ZN(n6836) );
  OAI222_X1 U8584 ( .A1(n8571), .A2(P2_U3151), .B1(n9018), .B2(n6836), .C1(
        n9015), .C2(n6835), .ZN(P2_U3282) );
  INV_X1 U8585 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10275) );
  INV_X1 U8586 ( .A(n7547), .ZN(n7543) );
  OAI222_X1 U8587 ( .A1(n9687), .A2(n10275), .B1(n9689), .B2(n6836), .C1(
        P1_U3086), .C2(n7543), .ZN(P1_U3342) );
  NAND2_X1 U8588 ( .A1(n9216), .A2(n9180), .ZN(n7007) );
  INV_X1 U8589 ( .A(n7007), .ZN(n6909) );
  AOI21_X1 U8590 ( .B1(n9805), .B2(n9504), .A(n7010), .ZN(n6837) );
  AOI211_X1 U8591 ( .C1(n6884), .C2(n7005), .A(n6909), .B(n6837), .ZN(n6931)
         );
  NAND2_X1 U8592 ( .A1(n5819), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6838) );
  OAI21_X1 U8593 ( .B1(n6931), .B2(n5819), .A(n6838), .ZN(P1_U3522) );
  NAND2_X1 U8594 ( .A1(n9145), .A2(P1_U3973), .ZN(n6839) );
  OAI21_X1 U8595 ( .B1(P1_U3973), .B2(n7725), .A(n6839), .ZN(P1_U3577) );
  INV_X1 U8596 ( .A(n6847), .ZN(n6841) );
  AND2_X1 U8597 ( .A1(n6847), .A2(n6875), .ZN(n6848) );
  NAND2_X1 U8598 ( .A1(n6849), .A2(n6848), .ZN(n7152) );
  NOR2_X1 U8599 ( .A1(n7228), .A2(n6981), .ZN(n6850) );
  NAND2_X1 U8600 ( .A1(n6852), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6851) );
  NAND2_X1 U8601 ( .A1(n6855), .A2(n6851), .ZN(n6907) );
  NAND2_X1 U8602 ( .A1(n9218), .A2(n8129), .ZN(n6854) );
  AOI22_X1 U8603 ( .A1(n7005), .A2(n6915), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n6852), .ZN(n6853) );
  NAND2_X1 U8604 ( .A1(n6854), .A2(n6853), .ZN(n6908) );
  NAND2_X1 U8605 ( .A1(n6907), .A2(n6908), .ZN(n6857) );
  INV_X2 U8606 ( .A(n7152), .ZN(n8354) );
  NAND2_X1 U8607 ( .A1(n6855), .A2(n8354), .ZN(n6856) );
  NAND2_X1 U8608 ( .A1(n6857), .A2(n6856), .ZN(n6919) );
  NAND2_X1 U8609 ( .A1(n6859), .A2(n6915), .ZN(n6858) );
  AOI22_X1 U8610 ( .A1(n9216), .A2(n8129), .B1(n6915), .B2(n7232), .ZN(n6861)
         );
  NAND2_X1 U8611 ( .A1(n6860), .A2(n6861), .ZN(n6918) );
  INV_X1 U8612 ( .A(n6860), .ZN(n6863) );
  INV_X1 U8613 ( .A(n6861), .ZN(n6862) );
  NAND2_X1 U8614 ( .A1(n6863), .A2(n6862), .ZN(n6920) );
  NAND2_X1 U8615 ( .A1(n6918), .A2(n6920), .ZN(n6864) );
  XOR2_X1 U8616 ( .A(n6919), .B(n6864), .Z(n6890) );
  INV_X1 U8617 ( .A(n6865), .ZN(n6867) );
  OR2_X1 U8618 ( .A1(n6867), .A2(n6866), .ZN(n7000) );
  INV_X1 U8619 ( .A(n7000), .ZN(n6869) );
  NAND2_X1 U8620 ( .A1(n6869), .A2(n6868), .ZN(n6874) );
  INV_X1 U8621 ( .A(n6874), .ZN(n6871) );
  AND2_X1 U8622 ( .A1(n6871), .A2(n6870), .ZN(n6882) );
  NOR2_X1 U8623 ( .A1(n9801), .A2(n6872), .ZN(n6873) );
  NAND2_X1 U8624 ( .A1(n6874), .A2(n6886), .ZN(n6880) );
  NAND2_X1 U8625 ( .A1(n6876), .A2(n6875), .ZN(n6877) );
  NOR2_X1 U8626 ( .A1(n6878), .A2(n6877), .ZN(n6879) );
  NAND2_X1 U8627 ( .A1(n6880), .A2(n6879), .ZN(n9094) );
  INV_X1 U8628 ( .A(n9094), .ZN(n6881) );
  NAND2_X1 U8629 ( .A1(n6881), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6925) );
  AOI22_X1 U8630 ( .A1(n9215), .A2(n9180), .B1(n9181), .B2(n9218), .ZN(n7226)
         );
  INV_X1 U8631 ( .A(n6882), .ZN(n6885) );
  NAND2_X1 U8632 ( .A1(n6884), .A2(n6883), .ZN(n7004) );
  OAI22_X1 U8633 ( .A1(n7226), .A2(n9694), .B1(n9783), .B2(n9722), .ZN(n6888)
         );
  AOI21_X1 U8634 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n6925), .A(n6888), .ZN(
        n6889) );
  OAI21_X1 U8635 ( .B1(n6890), .B2(n9699), .A(n6889), .ZN(P1_U3222) );
  OAI21_X1 U8636 ( .B1(n6892), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6891), .ZN(
        n6895) );
  NAND2_X1 U8637 ( .A1(n7019), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6893) );
  OAI21_X1 U8638 ( .B1(n7019), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6893), .ZN(
        n6894) );
  NOR2_X1 U8639 ( .A1(n6895), .A2(n6894), .ZN(n7015) );
  AOI211_X1 U8640 ( .C1(n6895), .C2(n6894), .A(n9341), .B(n7015), .ZN(n6906)
         );
  AOI21_X1 U8641 ( .B1(n6898), .B2(n6897), .A(n6896), .ZN(n6901) );
  INV_X1 U8642 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6899) );
  MUX2_X1 U8643 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6899), .S(n7019), .Z(n6900)
         );
  NAND2_X1 U8644 ( .A1(n6900), .A2(n6901), .ZN(n7020) );
  OAI211_X1 U8645 ( .C1(n6901), .C2(n6900), .A(n9309), .B(n7020), .ZN(n6903)
         );
  AND2_X1 U8646 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9692) );
  AOI21_X1 U8647 ( .B1(n9349), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n9692), .ZN(
        n6902) );
  OAI211_X1 U8648 ( .C1(n9337), .C2(n6904), .A(n6903), .B(n6902), .ZN(n6905)
         );
  OR2_X1 U8649 ( .A1(n6906), .A2(n6905), .ZN(P1_U3253) );
  XNOR2_X1 U8650 ( .A(n6907), .B(n6908), .ZN(n9230) );
  AOI22_X1 U8651 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n6925), .B1(n9719), .B2(
        n6909), .ZN(n6911) );
  NAND2_X1 U8652 ( .A1(n9703), .A2(n7005), .ZN(n6910) );
  OAI211_X1 U8653 ( .C1(n9230), .C2(n9699), .A(n6911), .B(n6910), .ZN(P1_U3232) );
  OR2_X1 U8654 ( .A1(n7087), .A2(n9168), .ZN(n6913) );
  NAND2_X1 U8655 ( .A1(n9216), .A2(n9181), .ZN(n6912) );
  AND2_X1 U8656 ( .A1(n6913), .A2(n6912), .ZN(n7118) );
  OAI22_X1 U8657 ( .A1(n9789), .A2(n6981), .B1(n6990), .B2(n8356), .ZN(n6914)
         );
  XNOR2_X1 U8658 ( .A(n6914), .B(n8354), .ZN(n6987) );
  OR2_X1 U8659 ( .A1(n6990), .A2(n8353), .ZN(n6917) );
  NAND2_X1 U8660 ( .A1(n7126), .A2(n8130), .ZN(n6916) );
  NAND2_X1 U8661 ( .A1(n6917), .A2(n6916), .ZN(n6985) );
  XNOR2_X1 U8662 ( .A(n6987), .B(n6985), .ZN(n6923) );
  NAND2_X1 U8663 ( .A1(n6919), .A2(n6918), .ZN(n6921) );
  AND2_X1 U8664 ( .A1(n6921), .A2(n6920), .ZN(n6922) );
  OAI21_X1 U8665 ( .B1(n6923), .B2(n6922), .A(n6989), .ZN(n6924) );
  NAND2_X1 U8666 ( .A1(n6924), .A2(n9724), .ZN(n6927) );
  AOI22_X1 U8667 ( .A1(n9703), .A2(n7126), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n6925), .ZN(n6926) );
  OAI211_X1 U8668 ( .C1(n7118), .C2(n9694), .A(n6927), .B(n6926), .ZN(P1_U3237) );
  INV_X1 U8669 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10508) );
  INV_X1 U8670 ( .A(n6928), .ZN(n6929) );
  INV_X1 U8671 ( .A(n7867), .ZN(n7859) );
  OAI222_X1 U8672 ( .A1(n9687), .A2(n10508), .B1(n9686), .B2(n6929), .C1(
        P1_U3086), .C2(n7859), .ZN(P1_U3341) );
  INV_X1 U8673 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6930) );
  OAI222_X1 U8674 ( .A1(n9015), .A2(n6930), .B1(n9018), .B2(n6929), .C1(
        P2_U3151), .C2(n8568), .ZN(P2_U3281) );
  INV_X1 U8675 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6933) );
  OR2_X1 U8676 ( .A1(n6931), .A2(n5809), .ZN(n6932) );
  OAI21_X1 U8677 ( .B1(n9858), .B2(n6933), .A(n6932), .ZN(P1_U3453) );
  INV_X1 U8678 ( .A(n6934), .ZN(n6958) );
  INV_X1 U8679 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6980) );
  MUX2_X1 U8680 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n4508), .Z(n6935) );
  XOR2_X1 U8681 ( .A(n9892), .B(n6935), .Z(n9899) );
  AOI22_X1 U8682 ( .A1(n9899), .A2(n9900), .B1(n6935), .B2(n9892), .ZN(n9918)
         );
  MUX2_X1 U8683 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n9876), .Z(n6936) );
  XNOR2_X1 U8684 ( .A(n6936), .B(n6966), .ZN(n9919) );
  INV_X1 U8685 ( .A(n6966), .ZN(n9913) );
  INV_X1 U8686 ( .A(n6936), .ZN(n6937) );
  OAI22_X1 U8687 ( .A1(n9918), .A2(n9919), .B1(n9913), .B2(n6937), .ZN(n9935)
         );
  MUX2_X1 U8688 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n9876), .Z(n6938) );
  XNOR2_X1 U8689 ( .A(n6938), .B(n6968), .ZN(n9936) );
  NOR2_X1 U8690 ( .A1(n6938), .A2(n6968), .ZN(n6941) );
  MUX2_X1 U8691 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n9876), .Z(n7032) );
  XNOR2_X1 U8692 ( .A(n7032), .B(n7035), .ZN(n6940) );
  INV_X1 U8693 ( .A(n7031), .ZN(n6943) );
  NOR2_X2 U8694 ( .A1(n8528), .A2(n6939), .ZN(n10016) );
  OAI21_X1 U8695 ( .B1(n9934), .B2(n6941), .A(n6940), .ZN(n6942) );
  NAND3_X1 U8696 ( .A1(n6943), .A2(n10016), .A3(n6942), .ZN(n6979) );
  OR2_X1 U8697 ( .A1(n6226), .A2(P2_U3151), .ZN(n9011) );
  NOR2_X1 U8698 ( .A1(n6956), .A2(n9011), .ZN(n9881) );
  NAND2_X1 U8699 ( .A1(n9881), .A2(n9876), .ZN(n9928) );
  MUX2_X1 U8700 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6944), .S(n7035), .Z(n6953)
         );
  MUX2_X1 U8701 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6945), .S(n6966), .Z(n9910)
         );
  AND2_X1 U8702 ( .A1(n9884), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6946) );
  NAND2_X1 U8703 ( .A1(n5861), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6947) );
  NAND2_X1 U8704 ( .A1(n9910), .A2(n9909), .ZN(n9908) );
  NAND2_X1 U8705 ( .A1(n6966), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6948) );
  NAND2_X1 U8706 ( .A1(n9908), .A2(n6948), .ZN(n6949) );
  XNOR2_X1 U8707 ( .A(n6949), .B(n4962), .ZN(n9926) );
  NAND2_X1 U8708 ( .A1(n9926), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6951) );
  NAND2_X1 U8709 ( .A1(n6949), .A2(n6968), .ZN(n6950) );
  NAND2_X1 U8710 ( .A1(n6951), .A2(n6950), .ZN(n6952) );
  NAND2_X1 U8711 ( .A1(n6952), .A2(n6953), .ZN(n7034) );
  OAI21_X1 U8712 ( .B1(n6953), .B2(n6952), .A(n7034), .ZN(n6977) );
  NOR2_X1 U8713 ( .A1(n9876), .A2(P2_U3151), .ZN(n6954) );
  NAND2_X1 U8714 ( .A1(n6954), .A2(n6226), .ZN(n6955) );
  OR2_X1 U8715 ( .A1(n6956), .A2(n6955), .ZN(n6960) );
  INV_X1 U8716 ( .A(n9011), .ZN(n6957) );
  NAND2_X1 U8717 ( .A1(n6958), .A2(n6957), .ZN(n6959) );
  INV_X1 U8718 ( .A(n10008), .ZN(n9885) );
  INV_X1 U8719 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6961) );
  NOR2_X1 U8720 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6961), .ZN(n7310) );
  INV_X1 U8721 ( .A(n7310), .ZN(n6962) );
  OAI21_X1 U8722 ( .B1(n9885), .B2(n7035), .A(n6962), .ZN(n6976) );
  INV_X1 U8723 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6963) );
  MUX2_X1 U8724 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6963), .S(n6966), .Z(n9906)
         );
  NAND2_X1 U8725 ( .A1(n5861), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6965) );
  NAND2_X1 U8726 ( .A1(n9887), .A2(n6965), .ZN(n9905) );
  NAND2_X1 U8727 ( .A1(n9906), .A2(n9905), .ZN(n9904) );
  NAND2_X1 U8728 ( .A1(n6966), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6967) );
  INV_X1 U8729 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7286) );
  MUX2_X1 U8730 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7286), .S(n7035), .Z(n6971)
         );
  INV_X1 U8731 ( .A(n6971), .ZN(n6973) );
  NAND3_X1 U8732 ( .A1(n9923), .A2(n6973), .A3(n6972), .ZN(n6974) );
  AOI21_X1 U8733 ( .B1(n7037), .B2(n6974), .A(n10023), .ZN(n6975) );
  AOI211_X1 U8734 ( .C1(n10017), .C2(n6977), .A(n6976), .B(n6975), .ZN(n6978)
         );
  OAI211_X1 U8735 ( .C1(n9941), .C2(n6980), .A(n6979), .B(n6978), .ZN(P2_U3186) );
  NAND2_X1 U8736 ( .A1(n6991), .A2(n8130), .ZN(n6983) );
  NAND2_X1 U8737 ( .A1(n6984), .A2(n6983), .ZN(n7158) );
  XNOR2_X1 U8738 ( .A(n7160), .B(n7158), .ZN(n7156) );
  INV_X1 U8739 ( .A(n6985), .ZN(n6986) );
  NAND2_X1 U8740 ( .A1(n6987), .A2(n6986), .ZN(n6988) );
  XOR2_X1 U8741 ( .A(n7156), .B(n7157), .Z(n6994) );
  OAI22_X1 U8742 ( .A1(n6990), .A2(n9091), .B1(n7263), .B2(n9168), .ZN(n9755)
         );
  AOI22_X1 U8743 ( .A1(n9755), .A2(n9719), .B1(n9703), .B2(n6991), .ZN(n6993)
         );
  MUX2_X1 U8744 ( .A(n9727), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n6992) );
  OAI211_X1 U8745 ( .C1(n6994), .C2(n9699), .A(n6993), .B(n6992), .ZN(P1_U3218) );
  INV_X1 U8746 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6996) );
  INV_X1 U8747 ( .A(n6995), .ZN(n6997) );
  INV_X1 U8748 ( .A(n9974), .ZN(n8574) );
  OAI222_X1 U8749 ( .A1(n9015), .A2(n6996), .B1(n9018), .B2(n6997), .C1(
        P2_U3151), .C2(n8574), .ZN(P2_U3280) );
  INV_X1 U8750 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6998) );
  INV_X1 U8751 ( .A(n7860), .ZN(n9280) );
  OAI222_X1 U8752 ( .A1(n9687), .A2(n6998), .B1(n9686), .B2(n6997), .C1(
        P1_U3086), .C2(n9280), .ZN(P1_U3340) );
  INV_X1 U8753 ( .A(n6999), .ZN(n7002) );
  NOR2_X1 U8754 ( .A1(n7000), .A2(n9775), .ZN(n7001) );
  NAND2_X1 U8755 ( .A1(n7002), .A2(n7001), .ZN(n7003) );
  INV_X1 U8756 ( .A(n9773), .ZN(n9452) );
  NOR2_X1 U8757 ( .A1(n9570), .A2(n9850), .ZN(n9438) );
  OAI21_X1 U8758 ( .B1(n9438), .B2(n9731), .A(n7005), .ZN(n7013) );
  INV_X1 U8759 ( .A(n7006), .ZN(n7009) );
  NAND2_X1 U8760 ( .A1(n9759), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7008) );
  OAI211_X1 U8761 ( .C1(n7010), .C2(n7009), .A(n7008), .B(n7007), .ZN(n7011)
         );
  NAND2_X1 U8762 ( .A1(n7011), .A2(n9452), .ZN(n7012) );
  OAI211_X1 U8763 ( .C1(n7014), .C2(n9452), .A(n7013), .B(n7012), .ZN(P1_U3293) );
  NAND2_X1 U8764 ( .A1(n7109), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7016) );
  OAI21_X1 U8765 ( .B1(n7109), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7016), .ZN(
        n7017) );
  NOR2_X1 U8766 ( .A1(n7018), .A2(n7017), .ZN(n7103) );
  AOI211_X1 U8767 ( .C1(n7018), .C2(n7017), .A(n7103), .B(n9341), .ZN(n7030)
         );
  NAND2_X1 U8768 ( .A1(n7019), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7021) );
  NAND2_X1 U8769 ( .A1(n7021), .A2(n7020), .ZN(n7024) );
  INV_X1 U8770 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7022) );
  MUX2_X1 U8771 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n7022), .S(n7109), .Z(n7023)
         );
  NAND2_X1 U8772 ( .A1(n7023), .A2(n7024), .ZN(n7107) );
  OAI211_X1 U8773 ( .C1(n7024), .C2(n7023), .A(n9309), .B(n7107), .ZN(n7027)
         );
  NAND2_X1 U8774 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n7801) );
  INV_X1 U8775 ( .A(n7801), .ZN(n7025) );
  AOI21_X1 U8776 ( .B1(n9349), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n7025), .ZN(
        n7026) );
  OAI211_X1 U8777 ( .C1(n9337), .C2(n7028), .A(n7027), .B(n7026), .ZN(n7029)
         );
  OR2_X1 U8778 ( .A1(n7030), .A2(n7029), .ZN(P1_U3254) );
  AOI21_X1 U8779 ( .B1(n7032), .B2(n7035), .A(n7031), .ZN(n7175) );
  MUX2_X1 U8780 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n9876), .Z(n7172) );
  XNOR2_X1 U8781 ( .A(n7172), .B(n7182), .ZN(n7174) );
  XNOR2_X1 U8782 ( .A(n7175), .B(n7174), .ZN(n7047) );
  NAND2_X1 U8783 ( .A1(n7035), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7033) );
  NAND2_X1 U8784 ( .A1(n7034), .A2(n7033), .ZN(n7183) );
  XNOR2_X1 U8785 ( .A(n7183), .B(n4960), .ZN(n7181) );
  XNOR2_X1 U8786 ( .A(n7181), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n7045) );
  NAND2_X1 U8787 ( .A1(n7035), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7036) );
  OAI21_X1 U8788 ( .B1(n7039), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7194), .ZN(
        n7040) );
  INV_X1 U8789 ( .A(n7040), .ZN(n7043) );
  NAND2_X1 U8790 ( .A1(n10007), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n7042) );
  NOR2_X1 U8791 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5912), .ZN(n7449) );
  AOI21_X1 U8792 ( .B1(n10008), .B2(n4960), .A(n7449), .ZN(n7041) );
  OAI211_X1 U8793 ( .C1(n7043), .C2(n10023), .A(n7042), .B(n7041), .ZN(n7044)
         );
  AOI21_X1 U8794 ( .B1(n10017), .B2(n7045), .A(n7044), .ZN(n7046) );
  OAI21_X1 U8795 ( .B1(n7047), .B2(n9937), .A(n7046), .ZN(P2_U3187) );
  INV_X1 U8796 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7051) );
  NAND2_X1 U8797 ( .A1(n6830), .A2(n7218), .ZN(n8200) );
  AND2_X1 U8798 ( .A1(n7048), .A2(n8200), .ZN(n8163) );
  INV_X1 U8799 ( .A(n8163), .ZN(n7213) );
  OAI21_X1 U8800 ( .B1(n8808), .B2(n10083), .A(n7213), .ZN(n7049) );
  NAND2_X1 U8801 ( .A1(n8826), .A2(n8824), .ZN(n7209) );
  OAI211_X1 U8802 ( .C1(n7218), .C2(n10078), .A(n7049), .B(n7209), .ZN(n8904)
         );
  NAND2_X1 U8803 ( .A1(n8904), .A2(n10084), .ZN(n7050) );
  OAI21_X1 U8804 ( .B1(n7051), .B2(n10084), .A(n7050), .ZN(P2_U3390) );
  OAI21_X1 U8805 ( .B1(n7052), .B2(n8196), .A(n7053), .ZN(n7293) );
  XNOR2_X1 U8806 ( .A(n7055), .B(n7054), .ZN(n7056) );
  NAND2_X1 U8807 ( .A1(n7056), .A2(n8808), .ZN(n7058) );
  AOI22_X1 U8808 ( .A1(n8827), .A2(n6830), .B1(n8207), .B2(n8824), .ZN(n7057)
         );
  NAND2_X1 U8809 ( .A1(n7058), .A2(n7057), .ZN(n7290) );
  AOI21_X1 U8810 ( .B1(n10083), .B2(n7293), .A(n7290), .ZN(n7082) );
  OR2_X1 U8811 ( .A1(n7059), .A2(n8343), .ZN(n7060) );
  NAND2_X1 U8812 ( .A1(n7060), .A2(n8326), .ZN(n7063) );
  INV_X1 U8813 ( .A(n7063), .ZN(n7061) );
  OR2_X1 U8814 ( .A1(n7062), .A2(n7061), .ZN(n7065) );
  NAND2_X1 U8815 ( .A1(n7065), .A2(n7064), .ZN(n7205) );
  NAND3_X1 U8816 ( .A1(n7068), .A2(n7067), .A3(n7066), .ZN(n7203) );
  NOR2_X1 U8817 ( .A1(n7203), .A2(n7069), .ZN(n7071) );
  NAND2_X1 U8818 ( .A1(n10101), .A2(n10063), .ZN(n8882) );
  OAI22_X1 U8819 ( .A1(n8882), .A2(n7072), .B1(n10101), .B2(n9888), .ZN(n7073)
         );
  INV_X1 U8820 ( .A(n7073), .ZN(n7074) );
  OAI21_X1 U8821 ( .B1(n7082), .B2(n10098), .A(n7074), .ZN(P2_U3460) );
  INV_X1 U8822 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10292) );
  INV_X1 U8823 ( .A(n7075), .ZN(n7078) );
  INV_X1 U8824 ( .A(n9292), .ZN(n9295) );
  OAI222_X1 U8825 ( .A1(n9687), .A2(n10292), .B1(n9686), .B2(n7078), .C1(n9295), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U8826 ( .A(P1_U3973), .ZN(n9217) );
  NAND2_X1 U8827 ( .A1(n9217), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7076) );
  OAI21_X1 U8828 ( .B1(n7077), .B2(n9217), .A(n7076), .ZN(P1_U3583) );
  INV_X1 U8829 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7079) );
  INV_X1 U8830 ( .A(n9990), .ZN(n8567) );
  OAI222_X1 U8831 ( .A1(n9015), .A2(n7079), .B1(n8567), .B2(P2_U3151), .C1(
        n9018), .C2(n7078), .ZN(P2_U3279) );
  OAI22_X1 U8832 ( .A1(n7072), .A2(n8964), .B1(n10084), .B2(n5851), .ZN(n7080)
         );
  INV_X1 U8833 ( .A(n7080), .ZN(n7081) );
  OAI21_X1 U8834 ( .B1(n7082), .B2(n10086), .A(n7081), .ZN(P2_U3393) );
  XNOR2_X1 U8835 ( .A(n7083), .B(n7085), .ZN(n9804) );
  AND2_X1 U8836 ( .A1(n7688), .A2(n7220), .ZN(n7084) );
  XNOR2_X1 U8837 ( .A(n7086), .B(n7085), .ZN(n7088) );
  OAI22_X1 U8838 ( .A1(n7087), .A2(n9091), .B1(n7260), .B2(n9168), .ZN(n7168)
         );
  AOI21_X1 U8839 ( .B1(n7088), .B2(n9756), .A(n7168), .ZN(n9803) );
  MUX2_X1 U8840 ( .A(n9803), .B(n6746), .S(n9773), .Z(n7092) );
  AOI211_X1 U8841 ( .C1(n9800), .C2(n9766), .A(n9850), .B(n4589), .ZN(n9799)
         );
  INV_X1 U8842 ( .A(n7167), .ZN(n7089) );
  OAI22_X1 U8843 ( .A1(n9761), .A2(n4840), .B1(n9565), .B2(n7089), .ZN(n7090)
         );
  AOI21_X1 U8844 ( .B1(n9799), .B2(n9769), .A(n7090), .ZN(n7091) );
  OAI211_X1 U8845 ( .C1(n9804), .C2(n9556), .A(n7092), .B(n7091), .ZN(P1_U3289) );
  INV_X1 U8846 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n7093) );
  OR2_X1 U8847 ( .A1(n7094), .A2(n7093), .ZN(n7100) );
  INV_X1 U8848 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7095) );
  OR2_X1 U8849 ( .A1(n7096), .A2(n7095), .ZN(n7099) );
  INV_X1 U8850 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n7097) );
  OR2_X1 U8851 ( .A1(n5898), .A2(n7097), .ZN(n7098) );
  NAND4_X1 U8852 ( .A1(n7101), .A2(n7100), .A3(n7099), .A4(n7098), .ZN(n8605)
         );
  NAND2_X1 U8853 ( .A1(n8605), .A2(P2_U3893), .ZN(n7102) );
  OAI21_X1 U8854 ( .B1(P2_U3893), .B2(n6345), .A(n7102), .ZN(P2_U3522) );
  XNOR2_X1 U8855 ( .A(n7116), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n7105) );
  AOI21_X1 U8856 ( .B1(n7109), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7103), .ZN(
        n7104) );
  NAND2_X1 U8857 ( .A1(n7105), .A2(n7104), .ZN(n7357) );
  OAI21_X1 U8858 ( .B1(n7105), .B2(n7104), .A(n7357), .ZN(n7113) );
  INV_X1 U8859 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7106) );
  MUX2_X1 U8860 ( .A(n7106), .B(P1_REG1_REG_12__SCAN_IN), .S(n7116), .Z(n7111)
         );
  INV_X1 U8861 ( .A(n7107), .ZN(n7108) );
  AOI21_X1 U8862 ( .B1(n7109), .B2(P1_REG1_REG_11__SCAN_IN), .A(n7108), .ZN(
        n7110) );
  NAND2_X1 U8863 ( .A1(n7110), .A2(n7111), .ZN(n7360) );
  OAI21_X1 U8864 ( .B1(n7111), .B2(n7110), .A(n7360), .ZN(n7112) );
  AOI22_X1 U8865 ( .A1(n9319), .A2(n7113), .B1(n9309), .B2(n7112), .ZN(n7115)
         );
  AND2_X1 U8866 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9065) );
  AOI21_X1 U8867 ( .B1(n9349), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n9065), .ZN(
        n7114) );
  OAI211_X1 U8868 ( .C1(n7116), .C2(n9337), .A(n7115), .B(n7114), .ZN(P1_U3255) );
  XNOR2_X1 U8869 ( .A(n7121), .B(n7117), .ZN(n7119) );
  OAI21_X1 U8870 ( .B1(n7119), .B2(n9504), .A(n7118), .ZN(n9790) );
  INV_X1 U8871 ( .A(n9790), .ZN(n7130) );
  XNOR2_X1 U8872 ( .A(n7121), .B(n7120), .ZN(n9792) );
  INV_X1 U8873 ( .A(n7227), .ZN(n7123) );
  INV_X1 U8874 ( .A(n9767), .ZN(n7122) );
  OAI211_X1 U8875 ( .C1(n9789), .C2(n7123), .A(n7122), .B(n9765), .ZN(n9788)
         );
  INV_X1 U8876 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9236) );
  OAI22_X1 U8877 ( .A1(n9452), .A2(n7124), .B1(n9236), .B2(n9565), .ZN(n7125)
         );
  AOI21_X1 U8878 ( .B1(n9731), .B2(n7126), .A(n7125), .ZN(n7127) );
  OAI21_X1 U8879 ( .B1(n9570), .B2(n9788), .A(n7127), .ZN(n7128) );
  AOI21_X1 U8880 ( .B1(n9770), .B2(n9792), .A(n7128), .ZN(n7129) );
  OAI21_X1 U8881 ( .B1(n7130), .B2(n9773), .A(n7129), .ZN(P1_U3291) );
  AND2_X1 U8882 ( .A1(n7132), .A2(n7131), .ZN(n7151) );
  OAI22_X1 U8883 ( .A1(n8503), .A2(n8163), .B1(n8517), .B2(n7218), .ZN(n7133)
         );
  AOI21_X1 U8884 ( .B1(n8480), .B2(n8826), .A(n7133), .ZN(n7134) );
  OAI21_X1 U8885 ( .B1(n7151), .B2(n7210), .A(n7134), .ZN(P2_U3172) );
  OAI22_X1 U8886 ( .A1(n8476), .A2(n7135), .B1(n8517), .B2(n7072), .ZN(n7136)
         );
  AOI21_X1 U8887 ( .B1(n8480), .B2(n8207), .A(n7136), .ZN(n7142) );
  OAI21_X1 U8888 ( .B1(n7137), .B2(n7139), .A(n7138), .ZN(n7140) );
  NAND2_X1 U8889 ( .A1(n7140), .A2(n8505), .ZN(n7141) );
  OAI211_X1 U8890 ( .C1(n7151), .C2(n5847), .A(n7142), .B(n7141), .ZN(P2_U3162) );
  OAI21_X1 U8891 ( .B1(n7145), .B2(n7144), .A(n7143), .ZN(n7146) );
  NAND2_X1 U8892 ( .A1(n7146), .A2(n8505), .ZN(n7149) );
  OAI22_X1 U8893 ( .A1(n8476), .A2(n5863), .B1(n8517), .B2(n10028), .ZN(n7147)
         );
  AOI21_X1 U8894 ( .B1(n8480), .B2(n4507), .A(n7147), .ZN(n7148) );
  OAI211_X1 U8895 ( .C1(n7151), .C2(n7150), .A(n7149), .B(n7148), .ZN(P2_U3177) );
  OAI22_X1 U8896 ( .A1(n7263), .A2(n8356), .B1(n4840), .B2(n8358), .ZN(n7153)
         );
  XNOR2_X1 U8897 ( .A(n7153), .B(n8128), .ZN(n7257) );
  OR2_X1 U8898 ( .A1(n7263), .A2(n8353), .ZN(n7155) );
  NAND2_X1 U8899 ( .A1(n9800), .A2(n8130), .ZN(n7154) );
  NAND2_X1 U8900 ( .A1(n7155), .A2(n7154), .ZN(n7256) );
  XNOR2_X1 U8901 ( .A(n7257), .B(n7256), .ZN(n7166) );
  INV_X1 U8902 ( .A(n7158), .ZN(n7159) );
  NAND2_X1 U8903 ( .A1(n7160), .A2(n7159), .ZN(n7161) );
  INV_X1 U8904 ( .A(n7259), .ZN(n7165) );
  AOI211_X1 U8905 ( .C1(n7166), .C2(n7162), .A(n9699), .B(n7165), .ZN(n7171)
         );
  AOI22_X1 U8906 ( .A1(n7168), .A2(n9719), .B1(n7167), .B2(n9187), .ZN(n7169)
         );
  NAND2_X1 U8907 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9261) );
  OAI211_X1 U8908 ( .C1(n4840), .C2(n9722), .A(n7169), .B(n9261), .ZN(n7170)
         );
  OR2_X1 U8909 ( .A1(n7171), .A2(n7170), .ZN(P1_U3230) );
  INV_X1 U8910 ( .A(n7172), .ZN(n7173) );
  INV_X1 U8911 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7189) );
  NOR2_X1 U8912 ( .A1(n9876), .A2(n7189), .ZN(n7176) );
  AOI21_X1 U8913 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n9876), .A(n7176), .ZN(
        n7177) );
  INV_X1 U8914 ( .A(n7464), .ZN(n7197) );
  NAND2_X1 U8915 ( .A1(n7177), .A2(n7197), .ZN(n7472) );
  OAI21_X1 U8916 ( .B1(n7177), .B2(n7197), .A(n7472), .ZN(n7178) );
  AOI21_X1 U8917 ( .B1(n7179), .B2(n7178), .A(n7474), .ZN(n7202) );
  MUX2_X1 U8918 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n7180), .S(n7464), .Z(n7187)
         );
  NAND2_X1 U8919 ( .A1(n7181), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7185) );
  NAND2_X1 U8920 ( .A1(n7183), .A2(n7182), .ZN(n7184) );
  NAND2_X1 U8921 ( .A1(n7185), .A2(n7184), .ZN(n7186) );
  NAND2_X1 U8922 ( .A1(n7186), .A2(n7187), .ZN(n7463) );
  OAI21_X1 U8923 ( .B1(n7187), .B2(n7186), .A(n7463), .ZN(n7200) );
  INV_X1 U8924 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7188) );
  NOR2_X1 U8925 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7188), .ZN(n7600) );
  XNOR2_X1 U8926 ( .A(n7464), .B(n7189), .ZN(n7191) );
  INV_X1 U8927 ( .A(n7191), .ZN(n7193) );
  NAND3_X1 U8928 ( .A1(n7194), .A2(n7193), .A3(n7192), .ZN(n7195) );
  AOI21_X1 U8929 ( .B1(n7466), .B2(n7195), .A(n10023), .ZN(n7196) );
  AOI211_X1 U8930 ( .C1(n7197), .C2(n10008), .A(n7600), .B(n7196), .ZN(n7198)
         );
  OAI21_X1 U8931 ( .B1(n10118), .B2(n9941), .A(n7198), .ZN(n7199) );
  AOI21_X1 U8932 ( .B1(n10017), .B2(n7200), .A(n7199), .ZN(n7201) );
  OAI21_X1 U8933 ( .B1(n7202), .B2(n9937), .A(n7201), .ZN(P2_U3188) );
  NOR2_X1 U8934 ( .A1(n7204), .A2(n7203), .ZN(n7207) );
  INV_X1 U8935 ( .A(n7205), .ZN(n7206) );
  NAND2_X1 U8936 ( .A1(n7207), .A2(n7206), .ZN(n7214) );
  AND2_X1 U8937 ( .A1(n7208), .A2(n10078), .ZN(n7212) );
  OAI21_X1 U8938 ( .B1(n8819), .B2(n7210), .A(n7209), .ZN(n7211) );
  AOI21_X1 U8939 ( .B1(n7213), .B2(n7212), .A(n7211), .ZN(n7216) );
  MUX2_X1 U8940 ( .A(n7216), .B(n7215), .S(n8812), .Z(n7217) );
  OAI21_X1 U8941 ( .B1(n8733), .B2(n7218), .A(n7217), .ZN(P2_U3233) );
  XNOR2_X1 U8942 ( .A(n7223), .B(n7219), .ZN(n9781) );
  NOR2_X1 U8943 ( .A1(n9730), .A2(n7220), .ZN(n9734) );
  INV_X1 U8944 ( .A(n9734), .ZN(n7447) );
  OAI21_X1 U8945 ( .B1(n7223), .B2(n7222), .A(n7221), .ZN(n7224) );
  NAND2_X1 U8946 ( .A1(n7224), .A2(n9756), .ZN(n7225) );
  OAI211_X1 U8947 ( .C1(n9781), .C2(n7688), .A(n7226), .B(n7225), .ZN(n9784)
         );
  NAND2_X1 U8948 ( .A1(n9784), .A2(n9452), .ZN(n7234) );
  OAI211_X1 U8949 ( .C1(n7228), .C2(n9783), .A(n9765), .B(n7227), .ZN(n9782)
         );
  NOR2_X1 U8950 ( .A1(n9570), .A2(n9782), .ZN(n7231) );
  INV_X1 U8951 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9219) );
  OAI22_X1 U8952 ( .A1(n9452), .A2(n7229), .B1(n9219), .B2(n9565), .ZN(n7230)
         );
  AOI211_X1 U8953 ( .C1(n9731), .C2(n7232), .A(n7231), .B(n7230), .ZN(n7233)
         );
  OAI211_X1 U8954 ( .C1(n9781), .C2(n7447), .A(n7234), .B(n7233), .ZN(P1_U3292) );
  INV_X1 U8955 ( .A(n7235), .ZN(n7237) );
  INV_X1 U8956 ( .A(n10009), .ZN(n8577) );
  OAI222_X1 U8957 ( .A1(n9015), .A2(n7236), .B1(n9018), .B2(n7237), .C1(
        P2_U3151), .C2(n8577), .ZN(P2_U3278) );
  OAI222_X1 U8958 ( .A1(n9687), .A2(n10447), .B1(n9686), .B2(n7237), .C1(
        P1_U3086), .C2(n9313), .ZN(P1_U3338) );
  XNOR2_X1 U8959 ( .A(n7238), .B(n7244), .ZN(n7239) );
  NAND2_X1 U8960 ( .A1(n7239), .A2(n9756), .ZN(n7243) );
  OR2_X1 U8961 ( .A1(n7260), .A2(n9091), .ZN(n7241) );
  NAND2_X1 U8962 ( .A1(n9210), .A2(n9180), .ZN(n7240) );
  NAND2_X1 U8963 ( .A1(n7241), .A2(n7240), .ZN(n7377) );
  INV_X1 U8964 ( .A(n7377), .ZN(n7242) );
  NAND2_X1 U8965 ( .A1(n7243), .A2(n7242), .ZN(n9820) );
  INV_X1 U8966 ( .A(n9820), .ZN(n7252) );
  XNOR2_X1 U8967 ( .A(n7245), .B(n7244), .ZN(n9815) );
  NAND2_X1 U8968 ( .A1(n9748), .A2(n7381), .ZN(n7246) );
  NAND2_X1 U8969 ( .A1(n7246), .A2(n9765), .ZN(n7247) );
  OR2_X1 U8970 ( .A1(n7247), .A2(n7395), .ZN(n9816) );
  AOI22_X1 U8971 ( .A1(n9730), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7376), .B2(
        n9759), .ZN(n7249) );
  NAND2_X1 U8972 ( .A1(n9731), .A2(n7381), .ZN(n7248) );
  OAI211_X1 U8973 ( .C1(n9816), .C2(n9570), .A(n7249), .B(n7248), .ZN(n7250)
         );
  AOI21_X1 U8974 ( .B1(n9815), .B2(n9770), .A(n7250), .ZN(n7251) );
  OAI21_X1 U8975 ( .B1(n7252), .B2(n9773), .A(n7251), .ZN(P1_U3287) );
  OR2_X1 U8976 ( .A1(n7260), .A2(n8353), .ZN(n7255) );
  NAND2_X1 U8977 ( .A1(n7253), .A2(n8130), .ZN(n7254) );
  NAND2_X1 U8978 ( .A1(n7255), .A2(n7254), .ZN(n7329) );
  INV_X1 U8979 ( .A(n7329), .ZN(n7333) );
  NAND2_X1 U8980 ( .A1(n7257), .A2(n7256), .ZN(n7258) );
  OAI22_X1 U8981 ( .A1(n7260), .A2(n8356), .B1(n9809), .B2(n8358), .ZN(n7261)
         );
  XNOR2_X1 U8982 ( .A(n7261), .B(n8128), .ZN(n7371) );
  INV_X1 U8983 ( .A(n7371), .ZN(n7332) );
  XNOR2_X1 U8984 ( .A(n7340), .B(n7332), .ZN(n7262) );
  NAND2_X1 U8985 ( .A1(n7262), .A2(n7333), .ZN(n7370) );
  OAI21_X1 U8986 ( .B1(n7333), .B2(n7262), .A(n7370), .ZN(n7267) );
  OAI22_X1 U8987 ( .A1(n7263), .A2(n9091), .B1(n7345), .B2(n9168), .ZN(n9741)
         );
  AOI22_X1 U8988 ( .A1(n9741), .A2(n9719), .B1(n9743), .B2(n9187), .ZN(n7265)
         );
  OAI211_X1 U8989 ( .C1(n9809), .C2(n9722), .A(n7265), .B(n7264), .ZN(n7266)
         );
  AOI21_X1 U8990 ( .B1(n7267), .B2(n9724), .A(n7266), .ZN(n7268) );
  INV_X1 U8991 ( .A(n7268), .ZN(P1_U3227) );
  INV_X1 U8992 ( .A(n8165), .ZN(n7269) );
  XNOR2_X1 U8993 ( .A(n7270), .B(n7269), .ZN(n7271) );
  NAND2_X1 U8994 ( .A1(n7271), .A2(n8808), .ZN(n7273) );
  AOI22_X1 U8995 ( .A1(n8827), .A2(n8207), .B1(n8212), .B2(n8824), .ZN(n7272)
         );
  AND2_X1 U8996 ( .A1(n7273), .A2(n7272), .ZN(n10035) );
  XNOR2_X1 U8997 ( .A(n7274), .B(n8165), .ZN(n10032) );
  AND2_X1 U8998 ( .A1(n7275), .A2(n8344), .ZN(n8833) );
  INV_X1 U8999 ( .A(n8816), .ZN(n8738) );
  NOR2_X1 U9000 ( .A1(n8835), .A2(n5882), .ZN(n7279) );
  OAI22_X1 U9001 ( .A1(n8733), .A2(n7277), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8819), .ZN(n7278) );
  AOI211_X1 U9002 ( .C1(n10032), .C2(n8738), .A(n7279), .B(n7278), .ZN(n7280)
         );
  OAI21_X1 U9003 ( .B1(n8812), .B2(n10035), .A(n7280), .ZN(P2_U3230) );
  XNOR2_X1 U9004 ( .A(n7281), .B(n8162), .ZN(n7282) );
  NAND2_X1 U9005 ( .A1(n7282), .A2(n8808), .ZN(n7284) );
  AOI22_X1 U9006 ( .A1(n8827), .A2(n4507), .B1(n8527), .B2(n8824), .ZN(n7283)
         );
  AND2_X1 U9007 ( .A1(n7284), .A2(n7283), .ZN(n10042) );
  XNOR2_X1 U9008 ( .A(n7285), .B(n8162), .ZN(n10038) );
  NOR2_X1 U9009 ( .A1(n8835), .A2(n7286), .ZN(n7288) );
  OAI22_X1 U9010 ( .A1(n8733), .A2(n8211), .B1(n7309), .B2(n8819), .ZN(n7287)
         );
  AOI211_X1 U9011 ( .C1(n10038), .C2(n8738), .A(n7288), .B(n7287), .ZN(n7289)
         );
  OAI21_X1 U9012 ( .B1(n8812), .B2(n10042), .A(n7289), .ZN(P2_U3229) );
  OAI22_X1 U9013 ( .A1(n8733), .A2(n7072), .B1(n5847), .B2(n8819), .ZN(n7292)
         );
  MUX2_X1 U9014 ( .A(n7290), .B(P2_REG2_REG_1__SCAN_IN), .S(n8812), .Z(n7291)
         );
  AOI211_X1 U9015 ( .C1(n8738), .C2(n7293), .A(n7292), .B(n7291), .ZN(n7294)
         );
  INV_X1 U9016 ( .A(n7294), .ZN(P2_U3232) );
  INV_X1 U9017 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10256) );
  NAND2_X1 U9018 ( .A1(n8514), .A2(n8207), .ZN(n7296) );
  NOR2_X1 U9019 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10256), .ZN(n9929) );
  AOI21_X1 U9020 ( .B1(n8501), .B2(n10033), .A(n9929), .ZN(n7295) );
  OAI211_X1 U9021 ( .C1(n7297), .C2(n8510), .A(n7296), .B(n7295), .ZN(n7303)
         );
  INV_X1 U9022 ( .A(n7298), .ZN(n7299) );
  AOI211_X1 U9023 ( .C1(n7301), .C2(n7300), .A(n8503), .B(n7299), .ZN(n7302)
         );
  AOI211_X1 U9024 ( .C1(n10256), .C2(n8497), .A(n7303), .B(n7302), .ZN(n7304)
         );
  INV_X1 U9025 ( .A(n7304), .ZN(P2_U3158) );
  INV_X1 U9026 ( .A(n9329), .ZN(n9303) );
  INV_X1 U9027 ( .A(n7305), .ZN(n7355) );
  INV_X1 U9028 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10505) );
  OAI222_X1 U9029 ( .A1(P1_U3086), .A2(n9303), .B1(n9686), .B2(n7355), .C1(
        n10505), .C2(n9687), .ZN(P1_U3337) );
  OAI21_X1 U9030 ( .B1(n7308), .B2(n7307), .A(n7306), .ZN(n7315) );
  NOR2_X1 U9031 ( .A1(n8511), .A2(n7309), .ZN(n7314) );
  NAND2_X1 U9032 ( .A1(n8514), .A2(n4507), .ZN(n7312) );
  AOI21_X1 U9033 ( .B1(n8501), .B2(n10039), .A(n7310), .ZN(n7311) );
  OAI211_X1 U9034 ( .C1(n8218), .C2(n8510), .A(n7312), .B(n7311), .ZN(n7313)
         );
  AOI211_X1 U9035 ( .C1(n7315), .C2(n8505), .A(n7314), .B(n7313), .ZN(n7316)
         );
  INV_X1 U9036 ( .A(n7316), .ZN(P2_U3170) );
  NAND2_X1 U9037 ( .A1(n9210), .A2(n8130), .ZN(n7317) );
  OAI21_X1 U9038 ( .B1(n9823), .B2(n8358), .A(n7317), .ZN(n7318) );
  XNOR2_X1 U9039 ( .A(n7318), .B(n8354), .ZN(n7321) );
  OR2_X1 U9040 ( .A1(n9823), .A2(n8356), .ZN(n7320) );
  NAND2_X1 U9041 ( .A1(n9210), .A2(n8129), .ZN(n7319) );
  AND2_X1 U9042 ( .A1(n7320), .A2(n7319), .ZN(n7322) );
  NAND2_X1 U9043 ( .A1(n7321), .A2(n7322), .ZN(n7560) );
  INV_X1 U9044 ( .A(n7321), .ZN(n7324) );
  INV_X1 U9045 ( .A(n7322), .ZN(n7323) );
  NAND2_X1 U9046 ( .A1(n7324), .A2(n7323), .ZN(n7325) );
  AND2_X1 U9047 ( .A1(n7560), .A2(n7325), .ZN(n7344) );
  OAI22_X1 U9048 ( .A1(n7345), .A2(n8356), .B1(n9817), .B2(n8358), .ZN(n7326)
         );
  XNOR2_X1 U9049 ( .A(n7326), .B(n8128), .ZN(n7334) );
  OR2_X1 U9050 ( .A1(n7345), .A2(n8353), .ZN(n7328) );
  NAND2_X1 U9051 ( .A1(n7381), .A2(n8130), .ZN(n7327) );
  NAND2_X1 U9052 ( .A1(n7328), .A2(n7327), .ZN(n7335) );
  AND2_X1 U9053 ( .A1(n7334), .A2(n7335), .ZN(n7331) );
  AND2_X1 U9054 ( .A1(n7371), .A2(n7329), .ZN(n7330) );
  INV_X1 U9055 ( .A(n7331), .ZN(n7373) );
  NAND3_X1 U9056 ( .A1(n7373), .A2(n7333), .A3(n7332), .ZN(n7338) );
  INV_X1 U9057 ( .A(n7334), .ZN(n7337) );
  INV_X1 U9058 ( .A(n7335), .ZN(n7336) );
  NAND2_X1 U9059 ( .A1(n7337), .A2(n7336), .ZN(n7372) );
  AND2_X1 U9060 ( .A1(n7338), .A2(n7372), .ZN(n7339) );
  OAI21_X1 U9061 ( .B1(n7344), .B2(n7341), .A(n7343), .ZN(n7353) );
  NOR2_X1 U9062 ( .A1(n9722), .A2(n9823), .ZN(n7352) );
  INV_X1 U9063 ( .A(n7396), .ZN(n7350) );
  OR2_X1 U9064 ( .A1(n7345), .A2(n9091), .ZN(n7347) );
  NAND2_X1 U9065 ( .A1(n9209), .A2(n9180), .ZN(n7346) );
  NAND2_X1 U9066 ( .A1(n7347), .A2(n7346), .ZN(n7391) );
  NAND2_X1 U9067 ( .A1(n7391), .A2(n9719), .ZN(n7349) );
  OAI211_X1 U9068 ( .C1(n9727), .C2(n7350), .A(n7349), .B(n7348), .ZN(n7351)
         );
  AOI211_X1 U9069 ( .C1(n7353), .C2(n9724), .A(n7352), .B(n7351), .ZN(n7354)
         );
  INV_X1 U9070 ( .A(n7354), .ZN(P1_U3213) );
  INV_X1 U9071 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7356) );
  INV_X1 U9072 ( .A(n8587), .ZN(n8597) );
  OAI222_X1 U9073 ( .A1(n9015), .A2(n7356), .B1(n8597), .B2(P2_U3151), .C1(
        n9018), .C2(n7355), .ZN(P2_U3277) );
  XNOR2_X1 U9074 ( .A(n7547), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n7359) );
  OAI21_X1 U9075 ( .B1(n7361), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7357), .ZN(
        n7358) );
  NOR2_X1 U9076 ( .A1(n7358), .A2(n7359), .ZN(n7546) );
  AOI211_X1 U9077 ( .C1(n7359), .C2(n7358), .A(n7546), .B(n9341), .ZN(n7366)
         );
  OAI21_X1 U9078 ( .B1(n7361), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7360), .ZN(
        n7364) );
  INV_X1 U9079 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9871) );
  MUX2_X1 U9080 ( .A(n9871), .B(P1_REG1_REG_13__SCAN_IN), .S(n7547), .Z(n7363)
         );
  OR2_X1 U9081 ( .A1(n7364), .A2(n7363), .ZN(n7542) );
  INV_X1 U9082 ( .A(n7542), .ZN(n7362) );
  AOI211_X1 U9083 ( .C1(n7364), .C2(n7363), .A(n7362), .B(n9339), .ZN(n7365)
         );
  NOR2_X1 U9084 ( .A1(n7366), .A2(n7365), .ZN(n7369) );
  NAND2_X1 U9085 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9126) );
  INV_X1 U9086 ( .A(n9126), .ZN(n7367) );
  AOI21_X1 U9087 ( .B1(n9349), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n7367), .ZN(
        n7368) );
  OAI211_X1 U9088 ( .C1(n7543), .C2(n9337), .A(n7369), .B(n7368), .ZN(P1_U3256) );
  OAI21_X1 U9089 ( .B1(n7371), .B2(n7340), .A(n7370), .ZN(n7375) );
  NAND2_X1 U9090 ( .A1(n7373), .A2(n7372), .ZN(n7374) );
  XNOR2_X1 U9091 ( .A(n7375), .B(n7374), .ZN(n7383) );
  INV_X1 U9092 ( .A(n7376), .ZN(n7379) );
  AOI22_X1 U9093 ( .A1(n7377), .A2(n9719), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n7378) );
  OAI21_X1 U9094 ( .B1(n7379), .B2(n9727), .A(n7378), .ZN(n7380) );
  AOI21_X1 U9095 ( .B1(n7381), .B2(n9703), .A(n7380), .ZN(n7382) );
  OAI21_X1 U9096 ( .B1(n7383), .B2(n9699), .A(n7382), .ZN(P1_U3239) );
  XNOR2_X1 U9097 ( .A(n7384), .B(n7389), .ZN(n7394) );
  NAND2_X1 U9098 ( .A1(n7386), .A2(n7385), .ZN(n7388) );
  INV_X1 U9099 ( .A(n7388), .ZN(n7390) );
  OR2_X1 U9100 ( .A1(n7388), .A2(n7387), .ZN(n7432) );
  OAI21_X1 U9101 ( .B1(n7390), .B2(n7389), .A(n7432), .ZN(n7392) );
  AOI21_X1 U9102 ( .B1(n7392), .B2(n9756), .A(n7391), .ZN(n7393) );
  OAI21_X1 U9103 ( .B1(n7394), .B2(n7688), .A(n7393), .ZN(n9824) );
  INV_X1 U9104 ( .A(n9824), .ZN(n7402) );
  INV_X1 U9105 ( .A(n7394), .ZN(n9826) );
  OAI211_X1 U9106 ( .C1(n7395), .C2(n9823), .A(n7440), .B(n9765), .ZN(n9822)
         );
  AOI22_X1 U9107 ( .A1(n9730), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7396), .B2(
        n9759), .ZN(n7399) );
  NAND2_X1 U9108 ( .A1(n9731), .A2(n7397), .ZN(n7398) );
  OAI211_X1 U9109 ( .C1(n9822), .C2(n9570), .A(n7399), .B(n7398), .ZN(n7400)
         );
  AOI21_X1 U9110 ( .B1(n9826), .B2(n9734), .A(n7400), .ZN(n7401) );
  OAI21_X1 U9111 ( .B1(n7402), .B2(n9773), .A(n7401), .ZN(P1_U3286) );
  XNOR2_X1 U9112 ( .A(n7403), .B(n7407), .ZN(n9835) );
  INV_X1 U9113 ( .A(n9835), .ZN(n7418) );
  INV_X1 U9114 ( .A(n7404), .ZN(n7405) );
  AOI21_X1 U9115 ( .B1(n7432), .B2(n7406), .A(n7405), .ZN(n7408) );
  XNOR2_X1 U9116 ( .A(n7408), .B(n7407), .ZN(n7409) );
  NAND2_X1 U9117 ( .A1(n7409), .A2(n9756), .ZN(n7410) );
  NAND2_X1 U9118 ( .A1(n9209), .A2(n9181), .ZN(n7581) );
  NAND2_X1 U9119 ( .A1(n7410), .A2(n7581), .ZN(n9839) );
  NAND2_X1 U9120 ( .A1(n7441), .A2(n7576), .ZN(n7411) );
  NAND2_X1 U9121 ( .A1(n7411), .A2(n9765), .ZN(n7412) );
  OR2_X1 U9122 ( .A1(n7412), .A2(n7534), .ZN(n7413) );
  OR2_X1 U9123 ( .A1(n7780), .A2(n9168), .ZN(n7582) );
  AND2_X1 U9124 ( .A1(n7413), .A2(n7582), .ZN(n9836) );
  AOI22_X1 U9125 ( .A1(n9730), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7585), .B2(
        n9759), .ZN(n7415) );
  NAND2_X1 U9126 ( .A1(n7576), .A2(n9731), .ZN(n7414) );
  OAI211_X1 U9127 ( .C1(n9836), .C2(n9570), .A(n7415), .B(n7414), .ZN(n7416)
         );
  AOI21_X1 U9128 ( .B1(n9839), .B2(n9452), .A(n7416), .ZN(n7417) );
  OAI21_X1 U9129 ( .B1(n9556), .B2(n7418), .A(n7417), .ZN(P1_U3284) );
  INV_X1 U9130 ( .A(n7419), .ZN(n7421) );
  OAI222_X1 U9131 ( .A1(n9015), .A2(n7420), .B1(n9018), .B2(n7421), .C1(n8596), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  OAI222_X1 U9132 ( .A1(n9687), .A2(n7422), .B1(n9686), .B2(n7421), .C1(
        P1_U3086), .C2(n5711), .ZN(P1_U3336) );
  XNOR2_X1 U9133 ( .A(n8527), .B(n10044), .ZN(n8168) );
  XOR2_X1 U9134 ( .A(n7423), .B(n8168), .Z(n7424) );
  AOI222_X1 U9135 ( .A1(n8808), .A2(n7424), .B1(n8526), .B2(n8824), .C1(n8212), 
        .C2(n8827), .ZN(n10043) );
  XOR2_X1 U9136 ( .A(n8168), .B(n7425), .Z(n10046) );
  NOR2_X1 U9137 ( .A1(n8835), .A2(n5910), .ZN(n7427) );
  OAI22_X1 U9138 ( .A1(n8733), .A2(n10044), .B1(n7448), .B2(n8819), .ZN(n7426)
         );
  AOI211_X1 U9139 ( .C1(n10046), .C2(n8738), .A(n7427), .B(n7426), .ZN(n7428)
         );
  OAI21_X1 U9140 ( .B1(n10043), .B2(n8812), .A(n7428), .ZN(P2_U3228) );
  NAND2_X1 U9141 ( .A1(n5136), .A2(n7429), .ZN(n7433) );
  XNOR2_X1 U9142 ( .A(n7430), .B(n7433), .ZN(n9828) );
  NAND2_X1 U9143 ( .A1(n7432), .A2(n7431), .ZN(n7434) );
  XNOR2_X1 U9144 ( .A(n7434), .B(n7433), .ZN(n7437) );
  OR2_X1 U9145 ( .A1(n7574), .A2(n9168), .ZN(n7436) );
  NAND2_X1 U9146 ( .A1(n9210), .A2(n9181), .ZN(n7435) );
  NAND2_X1 U9147 ( .A1(n7436), .A2(n7435), .ZN(n9720) );
  AOI21_X1 U9148 ( .B1(n7437), .B2(n9756), .A(n9720), .ZN(n7438) );
  OAI21_X1 U9149 ( .B1(n7688), .B2(n9828), .A(n7438), .ZN(n9831) );
  NAND2_X1 U9150 ( .A1(n9831), .A2(n9452), .ZN(n7446) );
  INV_X1 U9151 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7439) );
  OAI22_X1 U9152 ( .A1(n9452), .A2(n7439), .B1(n9728), .B2(n9565), .ZN(n7444)
         );
  INV_X1 U9153 ( .A(n7440), .ZN(n7442) );
  INV_X1 U9154 ( .A(n7566), .ZN(n9830) );
  OAI211_X1 U9155 ( .C1(n7442), .C2(n9830), .A(n9765), .B(n7441), .ZN(n9829)
         );
  NOR2_X1 U9156 ( .A1(n9829), .A2(n9570), .ZN(n7443) );
  AOI211_X1 U9157 ( .C1(n9731), .C2(n7566), .A(n7444), .B(n7443), .ZN(n7445)
         );
  OAI211_X1 U9158 ( .C1(n9828), .C2(n7447), .A(n7446), .B(n7445), .ZN(P1_U3285) );
  INV_X1 U9159 ( .A(n7448), .ZN(n7460) );
  NAND2_X1 U9160 ( .A1(n8514), .A2(n8212), .ZN(n7451) );
  AOI21_X1 U9161 ( .B1(n8501), .B2(n8217), .A(n7449), .ZN(n7450) );
  OAI211_X1 U9162 ( .C1(n7452), .C2(n8510), .A(n7451), .B(n7450), .ZN(n7459)
         );
  INV_X1 U9163 ( .A(n7453), .ZN(n7455) );
  NAND3_X1 U9164 ( .A1(n7306), .A2(n7455), .A3(n7454), .ZN(n7456) );
  AOI21_X1 U9165 ( .B1(n7457), .B2(n7456), .A(n8503), .ZN(n7458) );
  AOI211_X1 U9166 ( .C1(n7460), .C2(n8497), .A(n7459), .B(n7458), .ZN(n7461)
         );
  INV_X1 U9167 ( .A(n7461), .ZN(P2_U3167) );
  NAND2_X1 U9168 ( .A1(n7464), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7462) );
  NAND2_X1 U9169 ( .A1(n7463), .A2(n7462), .ZN(n7505) );
  XNOR2_X1 U9170 ( .A(n7505), .B(n7475), .ZN(n7508) );
  INV_X1 U9171 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7507) );
  XNOR2_X1 U9172 ( .A(n7508), .B(n7507), .ZN(n7481) );
  NAND2_X1 U9173 ( .A1(n7464), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7465) );
  OAI21_X1 U9174 ( .B1(n7467), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7512), .ZN(
        n7468) );
  INV_X1 U9175 ( .A(n10023), .ZN(n7516) );
  NAND2_X1 U9176 ( .A1(n7468), .A2(n7516), .ZN(n7471) );
  INV_X1 U9177 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10279) );
  NOR2_X1 U9178 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10279), .ZN(n7632) );
  AOI21_X1 U9179 ( .B1(n10008), .B2(n4959), .A(n7632), .ZN(n7470) );
  NAND2_X1 U9180 ( .A1(n10007), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7469) );
  NAND3_X1 U9181 ( .A1(n7471), .A2(n7470), .A3(n7469), .ZN(n7480) );
  INV_X1 U9182 ( .A(n7472), .ZN(n7473) );
  MUX2_X1 U9183 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n9876), .Z(n7496) );
  XNOR2_X1 U9184 ( .A(n7496), .B(n7475), .ZN(n7476) );
  AOI21_X1 U9185 ( .B1(n7477), .B2(n7476), .A(n7497), .ZN(n7478) );
  NOR2_X1 U9186 ( .A1(n7478), .A2(n9937), .ZN(n7479) );
  AOI211_X1 U9187 ( .C1(n10017), .C2(n7481), .A(n7480), .B(n7479), .ZN(n7482)
         );
  INV_X1 U9188 ( .A(n7482), .ZN(P2_U3189) );
  NAND2_X1 U9189 ( .A1(n7483), .A2(n7484), .ZN(n7485) );
  XNOR2_X1 U9190 ( .A(n8526), .B(n7491), .ZN(n8166) );
  XNOR2_X1 U9191 ( .A(n7485), .B(n8166), .ZN(n10050) );
  INV_X1 U9192 ( .A(n10050), .ZN(n7495) );
  INV_X1 U9193 ( .A(n8166), .ZN(n7486) );
  XNOR2_X1 U9194 ( .A(n7487), .B(n7486), .ZN(n7488) );
  NAND2_X1 U9195 ( .A1(n7488), .A2(n8808), .ZN(n7490) );
  AOI22_X1 U9196 ( .A1(n8827), .A2(n8527), .B1(n8525), .B2(n8824), .ZN(n7489)
         );
  NAND2_X1 U9197 ( .A1(n7490), .A2(n7489), .ZN(n10049) );
  NOR2_X1 U9198 ( .A1(n8835), .A2(n7189), .ZN(n7493) );
  OAI22_X1 U9199 ( .A1(n8733), .A2(n7491), .B1(n7599), .B2(n8819), .ZN(n7492)
         );
  AOI211_X1 U9200 ( .C1(n10049), .C2(n8835), .A(n7493), .B(n7492), .ZN(n7494)
         );
  OAI21_X1 U9201 ( .B1(n8816), .B2(n7495), .A(n7494), .ZN(P2_U3227) );
  INV_X1 U9202 ( .A(n7496), .ZN(n7498) );
  OR2_X1 U9203 ( .A1(n9876), .A2(n7513), .ZN(n7500) );
  NAND2_X1 U9204 ( .A1(n9876), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7499) );
  NAND2_X1 U9205 ( .A1(n7500), .A2(n7499), .ZN(n7501) );
  NOR2_X1 U9206 ( .A1(n7501), .A2(n7750), .ZN(n7759) );
  AOI21_X1 U9207 ( .B1(n7750), .B2(n7501), .A(n7759), .ZN(n7502) );
  INV_X1 U9208 ( .A(n7502), .ZN(n7503) );
  NOR2_X1 U9209 ( .A1(n7504), .A2(n7503), .ZN(n7758) );
  AOI21_X1 U9210 ( .B1(n7504), .B2(n7503), .A(n7758), .ZN(n7525) );
  INV_X1 U9211 ( .A(n7505), .ZN(n7506) );
  OAI22_X1 U9212 ( .A1(n7508), .A2(n7507), .B1(n4959), .B2(n7506), .ZN(n7510)
         );
  AOI22_X1 U9213 ( .A1(n7519), .A2(n5953), .B1(P2_REG1_REG_8__SCAN_IN), .B2(
        n7750), .ZN(n7509) );
  NAND2_X1 U9214 ( .A1(n7509), .A2(n7510), .ZN(n7746) );
  OAI21_X1 U9215 ( .B1(n7510), .B2(n7509), .A(n7746), .ZN(n7523) );
  INV_X1 U9216 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10124) );
  NAND2_X1 U9217 ( .A1(n7512), .A2(n7511), .ZN(n7515) );
  AOI21_X1 U9218 ( .B1(n7519), .B2(n7513), .A(n4558), .ZN(n7514) );
  NOR2_X1 U9219 ( .A1(n7515), .A2(n7514), .ZN(n7517) );
  OAI21_X1 U9220 ( .B1(n7749), .B2(n7517), .A(n7516), .ZN(n7521) );
  NOR2_X1 U9221 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7518), .ZN(n7674) );
  AOI21_X1 U9222 ( .B1(n10008), .B2(n7519), .A(n7674), .ZN(n7520) );
  OAI211_X1 U9223 ( .C1(n10124), .C2(n9941), .A(n7521), .B(n7520), .ZN(n7522)
         );
  AOI21_X1 U9224 ( .B1(n10017), .B2(n7523), .A(n7522), .ZN(n7524) );
  OAI21_X1 U9225 ( .B1(n7525), .B2(n9937), .A(n7524), .ZN(P2_U3190) );
  OAI21_X1 U9226 ( .B1(n7527), .B2(n7530), .A(n7526), .ZN(n7590) );
  INV_X1 U9227 ( .A(n7590), .ZN(n7541) );
  AOI21_X1 U9228 ( .B1(n7530), .B2(n4929), .A(n7529), .ZN(n7533) );
  OR2_X1 U9229 ( .A1(n7574), .A2(n9091), .ZN(n7532) );
  OR2_X1 U9230 ( .A1(n7789), .A2(n9168), .ZN(n7531) );
  AND2_X1 U9231 ( .A1(n7532), .A2(n7531), .ZN(n9695) );
  OAI21_X1 U9232 ( .B1(n7533), .B2(n9504), .A(n9695), .ZN(n7588) );
  INV_X1 U9233 ( .A(n7534), .ZN(n7535) );
  AOI211_X1 U9234 ( .C1(n9704), .C2(n7535), .A(n9850), .B(n7684), .ZN(n7589)
         );
  NAND2_X1 U9235 ( .A1(n7589), .A2(n9769), .ZN(n7538) );
  AOI22_X1 U9236 ( .A1(n9730), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7536), .B2(
        n9759), .ZN(n7537) );
  OAI211_X1 U9237 ( .C1(n7593), .C2(n9761), .A(n7538), .B(n7537), .ZN(n7539)
         );
  AOI21_X1 U9238 ( .B1(n7588), .B2(n9452), .A(n7539), .ZN(n7540) );
  OAI21_X1 U9239 ( .B1(n7541), .B2(n9556), .A(n7540), .ZN(P1_U3283) );
  OAI21_X1 U9240 ( .B1(n9871), .B2(n7543), .A(n7542), .ZN(n7857) );
  INV_X1 U9241 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9873) );
  MUX2_X1 U9242 ( .A(n9873), .B(P1_REG1_REG_14__SCAN_IN), .S(n7867), .Z(n7855)
         );
  XNOR2_X1 U9243 ( .A(n7857), .B(n7855), .ZN(n7553) );
  INV_X1 U9244 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9024) );
  NOR2_X1 U9245 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9024), .ZN(n7544) );
  AOI21_X1 U9246 ( .B1(n9349), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n7544), .ZN(
        n7545) );
  OAI21_X1 U9247 ( .B1(n7859), .B2(n9337), .A(n7545), .ZN(n7552) );
  NAND2_X1 U9248 ( .A1(n7867), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7548) );
  OAI21_X1 U9249 ( .B1(n7867), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7548), .ZN(
        n7549) );
  NOR2_X1 U9250 ( .A1(n7550), .A2(n7549), .ZN(n7866) );
  AOI211_X1 U9251 ( .C1(n7550), .C2(n7549), .A(n9341), .B(n7866), .ZN(n7551)
         );
  AOI211_X1 U9252 ( .C1(n7553), .C2(n9309), .A(n7552), .B(n7551), .ZN(n7554)
         );
  INV_X1 U9253 ( .A(n7554), .ZN(P1_U3257) );
  INV_X1 U9254 ( .A(n7555), .ZN(n7558) );
  OAI222_X1 U9255 ( .A1(n9018), .A2(n7558), .B1(P2_U3151), .B2(n8343), .C1(
        n7556), .C2(n9015), .ZN(P2_U3275) );
  OAI222_X1 U9256 ( .A1(n9687), .A2(n7559), .B1(n9686), .B2(n7558), .C1(n7557), 
        .C2(P1_U3086), .ZN(P1_U3335) );
  NAND2_X1 U9257 ( .A1(n7561), .A2(n7560), .ZN(n7570) );
  NAND2_X1 U9258 ( .A1(n7566), .A2(n8120), .ZN(n7563) );
  NAND2_X1 U9259 ( .A1(n9209), .A2(n8130), .ZN(n7562) );
  NAND2_X1 U9260 ( .A1(n7563), .A2(n7562), .ZN(n7564) );
  XNOR2_X1 U9261 ( .A(n7564), .B(n8128), .ZN(n7568) );
  XNOR2_X1 U9262 ( .A(n7570), .B(n7568), .ZN(n9715) );
  AND2_X1 U9263 ( .A1(n9209), .A2(n8129), .ZN(n7565) );
  AOI21_X1 U9264 ( .B1(n7566), .B2(n8130), .A(n7565), .ZN(n9717) );
  INV_X1 U9265 ( .A(n7568), .ZN(n7569) );
  NAND2_X1 U9266 ( .A1(n7570), .A2(n7569), .ZN(n7577) );
  AND2_X1 U9267 ( .A1(n7567), .A2(n7577), .ZN(n7580) );
  NAND2_X1 U9268 ( .A1(n7576), .A2(n8120), .ZN(n7572) );
  OR2_X1 U9269 ( .A1(n7574), .A2(n8356), .ZN(n7571) );
  NAND2_X1 U9270 ( .A1(n7572), .A2(n7571), .ZN(n7573) );
  XNOR2_X1 U9271 ( .A(n7573), .B(n8128), .ZN(n7772) );
  NOR2_X1 U9272 ( .A1(n7574), .A2(n8353), .ZN(n7575) );
  AOI21_X1 U9273 ( .B1(n7576), .B2(n8130), .A(n7575), .ZN(n7773) );
  XNOR2_X1 U9274 ( .A(n7772), .B(n7773), .ZN(n7579) );
  AND2_X1 U9275 ( .A1(n7577), .A2(n7579), .ZN(n7578) );
  OAI211_X1 U9276 ( .C1(n7580), .C2(n7579), .A(n9724), .B(n7776), .ZN(n7587)
         );
  AOI21_X1 U9277 ( .B1(n7582), .B2(n7581), .A(n9694), .ZN(n7583) );
  AOI211_X1 U9278 ( .C1(n9187), .C2(n7585), .A(n7584), .B(n7583), .ZN(n7586)
         );
  OAI211_X1 U9279 ( .C1(n4851), .C2(n9722), .A(n7587), .B(n7586), .ZN(P1_U3231) );
  AOI211_X1 U9280 ( .C1(n9845), .C2(n7590), .A(n7589), .B(n7588), .ZN(n7596)
         );
  INV_X1 U9281 ( .A(n9645), .ZN(n7701) );
  AOI22_X1 U9282 ( .A1(n9704), .A2(n7701), .B1(n5819), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7591) );
  OAI21_X1 U9283 ( .B1(n7596), .B2(n5819), .A(n7591), .ZN(P1_U3532) );
  INV_X1 U9284 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7592) );
  OAI22_X1 U9285 ( .A1(n7593), .A2(n9675), .B1(n9858), .B2(n7592), .ZN(n7594)
         );
  INV_X1 U9286 ( .A(n7594), .ZN(n7595) );
  OAI21_X1 U9287 ( .B1(n7596), .B2(n5809), .A(n7595), .ZN(P1_U3483) );
  INV_X1 U9288 ( .A(n7597), .ZN(n7613) );
  OAI222_X1 U9289 ( .A1(n9018), .A2(n7613), .B1(P2_U3151), .B2(n8161), .C1(
        n7598), .C2(n9015), .ZN(P2_U3274) );
  INV_X1 U9290 ( .A(n7599), .ZN(n7610) );
  NAND2_X1 U9291 ( .A1(n8514), .A2(n8527), .ZN(n7602) );
  AOI21_X1 U9292 ( .B1(n8501), .B2(n10047), .A(n7600), .ZN(n7601) );
  OAI211_X1 U9293 ( .C1(n7603), .C2(n8510), .A(n7602), .B(n7601), .ZN(n7609)
         );
  INV_X1 U9294 ( .A(n7604), .ZN(n7605) );
  AOI211_X1 U9295 ( .C1(n7607), .C2(n7606), .A(n8503), .B(n7605), .ZN(n7608)
         );
  AOI211_X1 U9296 ( .C1(n7610), .C2(n8497), .A(n7609), .B(n7608), .ZN(n7611)
         );
  INV_X1 U9297 ( .A(n7611), .ZN(P2_U3179) );
  OAI222_X1 U9298 ( .A1(P1_U3086), .A2(n6840), .B1(n9686), .B2(n7613), .C1(
        n7612), .C2(n9687), .ZN(P1_U3334) );
  OAI21_X1 U9299 ( .B1(n7615), .B2(n7618), .A(n7614), .ZN(n7647) );
  INV_X1 U9300 ( .A(n7616), .ZN(n7711) );
  AOI211_X1 U9301 ( .C1(n8011), .C2(n7685), .A(n9850), .B(n7711), .ZN(n7648)
         );
  NAND2_X1 U9302 ( .A1(n7691), .A2(n7617), .ZN(n7619) );
  XNOR2_X1 U9303 ( .A(n7619), .B(n7618), .ZN(n7620) );
  NAND2_X1 U9304 ( .A1(n7620), .A2(n9756), .ZN(n7623) );
  OR2_X1 U9305 ( .A1(n8018), .A2(n9168), .ZN(n7622) );
  OR2_X1 U9306 ( .A1(n7789), .A2(n9091), .ZN(n7621) );
  AND2_X1 U9307 ( .A1(n7622), .A2(n7621), .ZN(n9063) );
  NAND2_X1 U9308 ( .A1(n7623), .A2(n9063), .ZN(n7652) );
  AOI211_X1 U9309 ( .C1(n7647), .C2(n9845), .A(n7648), .B(n7652), .ZN(n7628)
         );
  INV_X1 U9310 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7624) );
  OAI22_X1 U9311 ( .A1(n4852), .A2(n9675), .B1(n9858), .B2(n7624), .ZN(n7625)
         );
  INV_X1 U9312 ( .A(n7625), .ZN(n7626) );
  OAI21_X1 U9313 ( .B1(n7628), .B2(n5809), .A(n7626), .ZN(P1_U3489) );
  AOI22_X1 U9314 ( .A1(n8011), .A2(n7701), .B1(n5819), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n7627) );
  OAI21_X1 U9315 ( .B1(n7628), .B2(n5819), .A(n7627), .ZN(P1_U3534) );
  OAI21_X1 U9316 ( .B1(n7631), .B2(n7630), .A(n7629), .ZN(n7637) );
  NOR2_X1 U9317 ( .A1(n8511), .A2(n7660), .ZN(n7636) );
  NAND2_X1 U9318 ( .A1(n8514), .A2(n8526), .ZN(n7634) );
  AOI21_X1 U9319 ( .B1(n8501), .B2(n7663), .A(n7632), .ZN(n7633) );
  OAI211_X1 U9320 ( .C1(n4862), .C2(n8510), .A(n7634), .B(n7633), .ZN(n7635)
         );
  AOI211_X1 U9321 ( .C1(n7637), .C2(n8505), .A(n7636), .B(n7635), .ZN(n7638)
         );
  INV_X1 U9322 ( .A(n7638), .ZN(P2_U3153) );
  INV_X1 U9323 ( .A(n8239), .ZN(n8233) );
  XNOR2_X1 U9324 ( .A(n7639), .B(n8170), .ZN(n10059) );
  XNOR2_X1 U9325 ( .A(n7640), .B(n8170), .ZN(n7641) );
  NAND2_X1 U9326 ( .A1(n7641), .A2(n8808), .ZN(n7643) );
  AOI22_X1 U9327 ( .A1(n8827), .A2(n8525), .B1(n8523), .B2(n8824), .ZN(n7642)
         );
  NAND2_X1 U9328 ( .A1(n7643), .A2(n7642), .ZN(n10061) );
  AOI22_X1 U9329 ( .A1(n8812), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n8769), .B2(
        n7678), .ZN(n7644) );
  OAI21_X1 U9330 ( .B1(n10057), .B2(n8733), .A(n7644), .ZN(n7645) );
  AOI21_X1 U9331 ( .B1(n10061), .B2(n8835), .A(n7645), .ZN(n7646) );
  OAI21_X1 U9332 ( .B1(n10059), .B2(n8816), .A(n7646), .ZN(P2_U3225) );
  INV_X1 U9333 ( .A(n7647), .ZN(n7654) );
  NAND2_X1 U9334 ( .A1(n7648), .A2(n9769), .ZN(n7650) );
  AOI22_X1 U9335 ( .A1(n9730), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9066), .B2(
        n9759), .ZN(n7649) );
  OAI211_X1 U9336 ( .C1(n4852), .C2(n9761), .A(n7650), .B(n7649), .ZN(n7651)
         );
  AOI21_X1 U9337 ( .B1(n9452), .B2(n7652), .A(n7651), .ZN(n7653) );
  OAI21_X1 U9338 ( .B1(n7654), .B2(n9556), .A(n7653), .ZN(P1_U3281) );
  XNOR2_X1 U9339 ( .A(n7655), .B(n4665), .ZN(n10056) );
  INV_X1 U9340 ( .A(n10056), .ZN(n7666) );
  NAND2_X1 U9341 ( .A1(n8835), .A2(n8833), .ZN(n8616) );
  XNOR2_X1 U9342 ( .A(n7656), .B(n4665), .ZN(n7659) );
  NAND2_X1 U9343 ( .A1(n10056), .A2(n8823), .ZN(n7658) );
  AOI22_X1 U9344 ( .A1(n8827), .A2(n8526), .B1(n8524), .B2(n8824), .ZN(n7657)
         );
  OAI211_X1 U9345 ( .C1(n8831), .C2(n7659), .A(n7658), .B(n7657), .ZN(n10054)
         );
  NAND2_X1 U9346 ( .A1(n10054), .A2(n8810), .ZN(n7665) );
  OAI22_X1 U9347 ( .A1(n8810), .A2(n7661), .B1(n7660), .B2(n8819), .ZN(n7662)
         );
  AOI21_X1 U9348 ( .B1(n8813), .B2(n7663), .A(n7662), .ZN(n7664) );
  OAI211_X1 U9349 ( .C1(n7666), .C2(n8616), .A(n7665), .B(n7664), .ZN(P2_U3226) );
  INV_X1 U9350 ( .A(n7629), .ZN(n7670) );
  INV_X1 U9351 ( .A(n7667), .ZN(n7669) );
  NOR3_X1 U9352 ( .A1(n7670), .A2(n7669), .A3(n7668), .ZN(n7673) );
  INV_X1 U9353 ( .A(n7671), .ZN(n7672) );
  OAI21_X1 U9354 ( .B1(n7673), .B2(n7672), .A(n8505), .ZN(n7680) );
  AOI21_X1 U9355 ( .B1(n8514), .B2(n8525), .A(n7674), .ZN(n7675) );
  OAI21_X1 U9356 ( .B1(n7676), .B2(n8510), .A(n7675), .ZN(n7677) );
  AOI21_X1 U9357 ( .B1(n7678), .B2(n8497), .A(n7677), .ZN(n7679) );
  OAI211_X1 U9358 ( .C1(n10057), .C2(n8517), .A(n7680), .B(n7679), .ZN(
        P2_U3161) );
  INV_X1 U9359 ( .A(n7681), .ZN(n9853) );
  OAI21_X1 U9360 ( .B1(n7683), .B2(n7694), .A(n7682), .ZN(n9735) );
  INV_X1 U9361 ( .A(n7684), .ZN(n7687) );
  INV_X1 U9362 ( .A(n7685), .ZN(n7686) );
  AOI211_X1 U9363 ( .C1(n9732), .C2(n7687), .A(n9850), .B(n7686), .ZN(n9733)
         );
  INV_X1 U9364 ( .A(n7688), .ZN(n7736) );
  AOI22_X1 U9365 ( .A1(n9181), .A2(n9207), .B1(n9205), .B2(n9180), .ZN(n7802)
         );
  INV_X1 U9366 ( .A(n7802), .ZN(n7696) );
  NAND2_X1 U9367 ( .A1(n7690), .A2(n7689), .ZN(n7693) );
  INV_X1 U9368 ( .A(n7691), .ZN(n7692) );
  AOI211_X1 U9369 ( .C1(n7694), .C2(n7693), .A(n9504), .B(n7692), .ZN(n7695)
         );
  AOI211_X1 U9370 ( .C1(n7736), .C2(n9735), .A(n7696), .B(n7695), .ZN(n9738)
         );
  INV_X1 U9371 ( .A(n9738), .ZN(n7697) );
  AOI211_X1 U9372 ( .C1(n9853), .C2(n9735), .A(n9733), .B(n7697), .ZN(n7703)
         );
  INV_X1 U9373 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7698) );
  OAI22_X1 U9374 ( .A1(n7806), .A2(n9675), .B1(n9858), .B2(n7698), .ZN(n7699)
         );
  INV_X1 U9375 ( .A(n7699), .ZN(n7700) );
  OAI21_X1 U9376 ( .B1(n7703), .B2(n5809), .A(n7700), .ZN(P1_U3486) );
  AOI22_X1 U9377 ( .A1(n9732), .A2(n7701), .B1(n5819), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7702) );
  OAI21_X1 U9378 ( .B1(n7703), .B2(n5819), .A(n7702), .ZN(P1_U3533) );
  XNOR2_X1 U9379 ( .A(n7704), .B(n4923), .ZN(n7706) );
  OR2_X1 U9380 ( .A1(n8009), .A2(n9091), .ZN(n7705) );
  OAI21_X1 U9381 ( .B1(n8025), .B2(n9168), .A(n7705), .ZN(n9125) );
  AOI21_X1 U9382 ( .B1(n7706), .B2(n9756), .A(n9125), .ZN(n9842) );
  OAI21_X1 U9383 ( .B1(n7709), .B2(n7708), .A(n7707), .ZN(n9846) );
  NAND2_X1 U9384 ( .A1(n9846), .A2(n9770), .ZN(n7715) );
  INV_X1 U9385 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7710) );
  OAI22_X1 U9386 ( .A1(n9452), .A2(n7710), .B1(n9128), .B2(n9565), .ZN(n7713)
         );
  INV_X1 U9387 ( .A(n9137), .ZN(n9843) );
  OAI211_X1 U9388 ( .C1(n7711), .C2(n9843), .A(n9765), .B(n7737), .ZN(n9841)
         );
  NOR2_X1 U9389 ( .A1(n9841), .A2(n9570), .ZN(n7712) );
  AOI211_X1 U9390 ( .C1(n9731), .C2(n9137), .A(n7713), .B(n7712), .ZN(n7714)
         );
  OAI211_X1 U9391 ( .C1(n9773), .C2(n9842), .A(n7715), .B(n7714), .ZN(P1_U3280) );
  INV_X1 U9392 ( .A(n7716), .ZN(n7719) );
  OAI222_X1 U9393 ( .A1(n9015), .A2(n7718), .B1(n9018), .B2(n7719), .C1(n7717), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U9394 ( .A1(n9687), .A2(n10446), .B1(n9686), .B2(n7719), .C1(
        P1_U3086), .C2(n6842), .ZN(P1_U3333) );
  NAND2_X1 U9395 ( .A1(n7723), .A2(n7720), .ZN(n7722) );
  OAI211_X1 U9396 ( .C1(n10278), .C2(n9687), .A(n7722), .B(n7721), .ZN(
        P1_U3332) );
  NAND2_X1 U9397 ( .A1(n7723), .A2(n9010), .ZN(n7724) );
  OAI211_X1 U9398 ( .C1(n7725), .C2(n9015), .A(n7724), .B(n8351), .ZN(P2_U3272) );
  XNOR2_X1 U9399 ( .A(n7727), .B(n7726), .ZN(n9854) );
  OAI21_X1 U9400 ( .B1(n7730), .B2(n7729), .A(n7728), .ZN(n7731) );
  NAND2_X1 U9401 ( .A1(n7731), .A2(n9756), .ZN(n7734) );
  OR2_X1 U9402 ( .A1(n8018), .A2(n9091), .ZN(n7733) );
  NAND2_X1 U9403 ( .A1(n9204), .A2(n9180), .ZN(n7732) );
  AND2_X1 U9404 ( .A1(n7733), .A2(n7732), .ZN(n9025) );
  NAND2_X1 U9405 ( .A1(n7734), .A2(n9025), .ZN(n7735) );
  AOI21_X1 U9406 ( .B1(n9854), .B2(n7736), .A(n7735), .ZN(n9856) );
  INV_X1 U9407 ( .A(n9569), .ZN(n7739) );
  NAND2_X1 U9408 ( .A1(n7740), .A2(n7737), .ZN(n7738) );
  NAND2_X1 U9409 ( .A1(n7739), .A2(n7738), .ZN(n9851) );
  INV_X1 U9410 ( .A(n9438), .ZN(n7743) );
  AOI22_X1 U9411 ( .A1(n9730), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9028), .B2(
        n9759), .ZN(n7742) );
  NAND2_X1 U9412 ( .A1(n7740), .A2(n9731), .ZN(n7741) );
  OAI211_X1 U9413 ( .C1(n9851), .C2(n7743), .A(n7742), .B(n7741), .ZN(n7744)
         );
  AOI21_X1 U9414 ( .B1(n9854), .B2(n9734), .A(n7744), .ZN(n7745) );
  OAI21_X1 U9415 ( .B1(n9856), .B2(n9773), .A(n7745), .ZN(P1_U3279) );
  NAND2_X1 U9416 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7750), .ZN(n7747) );
  NAND2_X1 U9417 ( .A1(n7747), .A2(n7746), .ZN(n7903) );
  XNOR2_X1 U9418 ( .A(n7912), .B(n7903), .ZN(n7748) );
  NAND2_X1 U9419 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(n7748), .ZN(n7904) );
  OAI21_X1 U9420 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n7748), .A(n7904), .ZN(
        n7770) );
  INV_X1 U9421 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10128) );
  NOR2_X1 U9422 ( .A1(n9941), .A2(n10128), .ZN(n7769) );
  AOI21_X1 U9423 ( .B1(n7751), .B2(n7752), .A(n7913), .ZN(n7767) );
  OR2_X1 U9424 ( .A1(n9876), .A2(n7752), .ZN(n7754) );
  NAND2_X1 U9425 ( .A1(n9876), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7753) );
  AND2_X1 U9426 ( .A1(n7754), .A2(n7753), .ZN(n7755) );
  AND2_X1 U9427 ( .A1(n7755), .A2(n7912), .ZN(n7890) );
  INV_X1 U9428 ( .A(n7755), .ZN(n7756) );
  AND2_X1 U9429 ( .A1(n7756), .A2(n4983), .ZN(n7757) );
  OR2_X1 U9430 ( .A1(n7890), .A2(n7757), .ZN(n7760) );
  NOR2_X1 U9431 ( .A1(n7759), .A2(n7758), .ZN(n7761) );
  NAND2_X1 U9432 ( .A1(n7760), .A2(n7761), .ZN(n7763) );
  INV_X1 U9433 ( .A(n7889), .ZN(n7762) );
  NAND2_X1 U9434 ( .A1(n7763), .A2(n7762), .ZN(n7764) );
  NOR2_X1 U9435 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5974), .ZN(n7844) );
  AOI21_X1 U9436 ( .B1(n7764), .B2(n10016), .A(n7844), .ZN(n7766) );
  NAND2_X1 U9437 ( .A1(n10008), .A2(n7912), .ZN(n7765) );
  OAI211_X1 U9438 ( .C1(n7767), .C2(n10023), .A(n7766), .B(n7765), .ZN(n7768)
         );
  AOI211_X1 U9439 ( .C1(n7770), .C2(n10017), .A(n7769), .B(n7768), .ZN(n7771)
         );
  INV_X1 U9440 ( .A(n7771), .ZN(P2_U3191) );
  INV_X1 U9441 ( .A(n7772), .ZN(n7774) );
  OR2_X1 U9442 ( .A1(n7774), .A2(n7773), .ZN(n7775) );
  NAND2_X1 U9443 ( .A1(n9704), .A2(n8120), .ZN(n7778) );
  OR2_X1 U9444 ( .A1(n7780), .A2(n8356), .ZN(n7777) );
  NAND2_X1 U9445 ( .A1(n7778), .A2(n7777), .ZN(n7779) );
  INV_X1 U9446 ( .A(n9697), .ZN(n7784) );
  NAND2_X1 U9447 ( .A1(n9704), .A2(n8130), .ZN(n7782) );
  OR2_X1 U9448 ( .A1(n7780), .A2(n8353), .ZN(n7781) );
  NAND2_X1 U9449 ( .A1(n7782), .A2(n7781), .ZN(n9698) );
  NAND2_X1 U9450 ( .A1(n7784), .A2(n7783), .ZN(n7796) );
  INV_X1 U9451 ( .A(n7785), .ZN(n9696) );
  INV_X1 U9452 ( .A(n7795), .ZN(n7794) );
  NAND2_X1 U9453 ( .A1(n9732), .A2(n8120), .ZN(n7787) );
  OR2_X1 U9454 ( .A1(n7789), .A2(n8356), .ZN(n7786) );
  NAND2_X1 U9455 ( .A1(n7787), .A2(n7786), .ZN(n7788) );
  XNOR2_X1 U9456 ( .A(n7788), .B(n8354), .ZN(n7792) );
  NOR2_X1 U9457 ( .A1(n7789), .A2(n8353), .ZN(n7790) );
  AOI21_X1 U9458 ( .B1(n9732), .B2(n6915), .A(n7790), .ZN(n7791) );
  NAND2_X1 U9459 ( .A1(n7792), .A2(n7791), .ZN(n9058) );
  OR2_X1 U9460 ( .A1(n7792), .A2(n7791), .ZN(n7793) );
  AND2_X1 U9461 ( .A1(n9058), .A2(n7793), .ZN(n7797) );
  NOR3_X1 U9462 ( .A1(n9696), .A2(n7794), .A3(n7797), .ZN(n7800) );
  NAND2_X1 U9463 ( .A1(n7796), .A2(n7795), .ZN(n7798) );
  NAND2_X1 U9464 ( .A1(n7798), .A2(n7797), .ZN(n8005) );
  INV_X1 U9465 ( .A(n7799), .ZN(n9060) );
  OAI21_X1 U9466 ( .B1(n7800), .B2(n9060), .A(n9724), .ZN(n7805) );
  OAI21_X1 U9467 ( .B1(n7802), .B2(n9694), .A(n7801), .ZN(n7803) );
  AOI21_X1 U9468 ( .B1(n9729), .B2(n9187), .A(n7803), .ZN(n7804) );
  OAI211_X1 U9469 ( .C1(n7806), .C2(n9722), .A(n7805), .B(n7804), .ZN(P1_U3236) );
  INV_X1 U9470 ( .A(n7807), .ZN(n7819) );
  XOR2_X1 U9471 ( .A(n8172), .B(n7809), .Z(n10069) );
  INV_X1 U9472 ( .A(n10069), .ZN(n7817) );
  XOR2_X1 U9473 ( .A(n7810), .B(n8172), .Z(n7813) );
  NAND2_X1 U9474 ( .A1(n10069), .A2(n8823), .ZN(n7812) );
  AOI22_X1 U9475 ( .A1(n8827), .A2(n8524), .B1(n8522), .B2(n8824), .ZN(n7811)
         );
  OAI211_X1 U9476 ( .C1(n8831), .C2(n7813), .A(n7812), .B(n7811), .ZN(n10067)
         );
  NAND2_X1 U9477 ( .A1(n10067), .A2(n8810), .ZN(n7816) );
  OAI22_X1 U9478 ( .A1(n8810), .A2(n7752), .B1(n7847), .B2(n8819), .ZN(n7814)
         );
  AOI21_X1 U9479 ( .B1(n8813), .B2(n10065), .A(n7814), .ZN(n7815) );
  OAI211_X1 U9480 ( .C1(n7817), .C2(n8616), .A(n7816), .B(n7815), .ZN(P2_U3224) );
  OAI222_X1 U9481 ( .A1(n7820), .A2(P1_U3086), .B1(n9686), .B2(n7819), .C1(
        n7818), .C2(n9687), .ZN(P1_U3331) );
  XNOR2_X1 U9482 ( .A(n7821), .B(n8173), .ZN(n10075) );
  INV_X1 U9483 ( .A(n10075), .ZN(n7832) );
  NAND2_X1 U9484 ( .A1(n7810), .A2(n7822), .ZN(n7824) );
  NAND2_X1 U9485 ( .A1(n7824), .A2(n7823), .ZN(n7825) );
  XOR2_X1 U9486 ( .A(n8173), .B(n7825), .Z(n7828) );
  NAND2_X1 U9487 ( .A1(n10075), .A2(n8823), .ZN(n7827) );
  AOI22_X1 U9488 ( .A1(n8805), .A2(n8824), .B1(n8827), .B2(n8523), .ZN(n7826)
         );
  OAI211_X1 U9489 ( .C1(n8831), .C2(n7828), .A(n7827), .B(n7826), .ZN(n10073)
         );
  NAND2_X1 U9490 ( .A1(n10073), .A2(n8810), .ZN(n7831) );
  OAI22_X1 U9491 ( .A1(n8810), .A2(n7914), .B1(n7933), .B2(n8819), .ZN(n7829)
         );
  AOI21_X1 U9492 ( .B1(n8813), .B2(n10071), .A(n7829), .ZN(n7830) );
  OAI211_X1 U9493 ( .C1(n7832), .C2(n8616), .A(n7831), .B(n7830), .ZN(P2_U3223) );
  OAI211_X1 U9494 ( .C1(n7834), .C2(n4817), .A(n8808), .B(n7833), .ZN(n7836)
         );
  AOI22_X1 U9495 ( .A1(n8824), .A2(n8786), .B1(n8522), .B2(n8827), .ZN(n7835)
         );
  NAND2_X1 U9496 ( .A1(n7836), .A2(n7835), .ZN(n10080) );
  INV_X1 U9497 ( .A(n10080), .ZN(n7843) );
  OAI21_X1 U9498 ( .B1(n7838), .B2(n8176), .A(n7837), .ZN(n10082) );
  INV_X1 U9499 ( .A(n7839), .ZN(n10079) );
  NOR2_X1 U9500 ( .A1(n10079), .A2(n8733), .ZN(n7841) );
  OAI22_X1 U9501 ( .A1(n8810), .A2(n7884), .B1(n8477), .B2(n8819), .ZN(n7840)
         );
  AOI211_X1 U9502 ( .C1(n10082), .C2(n8738), .A(n7841), .B(n7840), .ZN(n7842)
         );
  OAI21_X1 U9503 ( .B1(n8812), .B2(n7843), .A(n7842), .ZN(P2_U3222) );
  AOI21_X1 U9504 ( .B1(n8514), .B2(n8524), .A(n7844), .ZN(n7846) );
  NAND2_X1 U9505 ( .A1(n8480), .A2(n8522), .ZN(n7845) );
  OAI211_X1 U9506 ( .C1(n8511), .C2(n7847), .A(n7846), .B(n7845), .ZN(n7853)
         );
  INV_X1 U9507 ( .A(n7848), .ZN(n7849) );
  AOI211_X1 U9508 ( .C1(n7851), .C2(n7850), .A(n8503), .B(n7849), .ZN(n7852)
         );
  AOI211_X1 U9509 ( .C1(n10065), .C2(n8501), .A(n7853), .B(n7852), .ZN(n7854)
         );
  INV_X1 U9510 ( .A(n7854), .ZN(P2_U3171) );
  INV_X1 U9511 ( .A(n7855), .ZN(n7856) );
  NAND2_X1 U9512 ( .A1(n7857), .A2(n7856), .ZN(n7858) );
  OAI21_X1 U9513 ( .B1(n9873), .B2(n7859), .A(n7858), .ZN(n7861) );
  NAND2_X1 U9514 ( .A1(n7860), .A2(n7861), .ZN(n7862) );
  XNOR2_X1 U9515 ( .A(n9280), .B(n7861), .ZN(n9284) );
  NAND2_X1 U9516 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9284), .ZN(n9283) );
  NAND2_X1 U9517 ( .A1(n7862), .A2(n9283), .ZN(n7865) );
  INV_X1 U9518 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7863) );
  MUX2_X1 U9519 ( .A(n7863), .B(P1_REG1_REG_16__SCAN_IN), .S(n9292), .Z(n7864)
         );
  NOR2_X1 U9520 ( .A1(n7864), .A2(n7865), .ZN(n9294) );
  AOI21_X1 U9521 ( .B1(n7865), .B2(n7864), .A(n9294), .ZN(n7878) );
  NOR2_X1 U9522 ( .A1(n7868), .A2(n9280), .ZN(n7869) );
  INV_X1 U9523 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9567) );
  XNOR2_X1 U9524 ( .A(n9280), .B(n7868), .ZN(n9286) );
  NOR2_X1 U9525 ( .A1(n9567), .A2(n9286), .ZN(n9285) );
  NOR2_X1 U9526 ( .A1(n7869), .A2(n9285), .ZN(n7872) );
  NAND2_X1 U9527 ( .A1(n9292), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7870) );
  OAI21_X1 U9528 ( .B1(n9292), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7870), .ZN(
        n7871) );
  NOR2_X1 U9529 ( .A1(n7872), .A2(n7871), .ZN(n9291) );
  AOI211_X1 U9530 ( .C1(n7872), .C2(n7871), .A(n9291), .B(n9341), .ZN(n7873)
         );
  INV_X1 U9531 ( .A(n7873), .ZN(n7877) );
  INV_X1 U9532 ( .A(n9337), .ZN(n9265) );
  INV_X1 U9533 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7874) );
  NAND2_X1 U9534 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9082) );
  OAI21_X1 U9535 ( .B1(n9263), .B2(n7874), .A(n9082), .ZN(n7875) );
  AOI21_X1 U9536 ( .B1(n9292), .B2(n9265), .A(n7875), .ZN(n7876) );
  OAI211_X1 U9537 ( .C1(n7878), .C2(n9339), .A(n7877), .B(n7876), .ZN(P1_U3259) );
  INV_X1 U9538 ( .A(n7879), .ZN(n7882) );
  OAI222_X1 U9539 ( .A1(n9018), .A2(n7882), .B1(P2_U3151), .B2(n7881), .C1(
        n7880), .C2(n9015), .ZN(P2_U3270) );
  OAI222_X1 U9540 ( .A1(n7883), .A2(P1_U3086), .B1(n9686), .B2(n7882), .C1(
        n10477), .C2(n9687), .ZN(P1_U3330) );
  OR2_X1 U9541 ( .A1(n9876), .A2(n7884), .ZN(n7886) );
  NAND2_X1 U9542 ( .A1(n9876), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7885) );
  AND2_X1 U9543 ( .A1(n7886), .A2(n7885), .ZN(n7894) );
  AND2_X1 U9544 ( .A1(n7894), .A2(n7965), .ZN(n7897) );
  OR2_X1 U9545 ( .A1(n9876), .A2(n7914), .ZN(n7888) );
  NAND2_X1 U9546 ( .A1(n9876), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7887) );
  NAND2_X1 U9547 ( .A1(n7888), .A2(n7887), .ZN(n7891) );
  NOR2_X1 U9548 ( .A1(n7891), .A2(n7915), .ZN(n7893) );
  AOI21_X1 U9549 ( .B1(n7915), .B2(n7891), .A(n7893), .ZN(n7892) );
  INV_X1 U9550 ( .A(n7892), .ZN(n7945) );
  NOR2_X1 U9551 ( .A1(n7944), .A2(n7945), .ZN(n7943) );
  NOR2_X1 U9552 ( .A1(n7893), .A2(n7943), .ZN(n7959) );
  INV_X1 U9553 ( .A(n7894), .ZN(n7895) );
  AND2_X1 U9554 ( .A1(n7895), .A2(n7917), .ZN(n7896) );
  OR2_X1 U9555 ( .A1(n7897), .A2(n7896), .ZN(n7960) );
  OR2_X1 U9556 ( .A1(n9876), .A2(n7898), .ZN(n7900) );
  NAND2_X1 U9557 ( .A1(n9876), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7899) );
  AND2_X1 U9558 ( .A1(n7900), .A2(n7899), .ZN(n7901) );
  NOR2_X1 U9559 ( .A1(n7901), .A2(n8570), .ZN(n8548) );
  AND2_X1 U9560 ( .A1(n7901), .A2(n8570), .ZN(n8547) );
  NOR2_X1 U9561 ( .A1(n8548), .A2(n8547), .ZN(n7902) );
  XNOR2_X1 U9562 ( .A(n8550), .B(n7902), .ZN(n7927) );
  AOI22_X1 U9563 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8531), .B1(n8570), .B2(
        n8899), .ZN(n7909) );
  AOI22_X1 U9564 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7915), .B1(n7949), .B2(
        n5985), .ZN(n7942) );
  NAND2_X1 U9565 ( .A1(n4983), .A2(n7903), .ZN(n7905) );
  NAND2_X1 U9566 ( .A1(n7917), .A2(n7906), .ZN(n7907) );
  NAND2_X1 U9567 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n7956), .ZN(n7955) );
  OAI21_X1 U9568 ( .B1(n7909), .B2(n7908), .A(n8569), .ZN(n7925) );
  INV_X1 U9569 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n10140) );
  INV_X1 U9570 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10463) );
  NOR2_X1 U9571 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10463), .ZN(n8405) );
  AOI21_X1 U9572 ( .B1(n10008), .B2(n8570), .A(n8405), .ZN(n7910) );
  OAI21_X1 U9573 ( .B1(n9941), .B2(n10140), .A(n7910), .ZN(n7924) );
  MUX2_X1 U9574 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7914), .S(n7949), .Z(n7938)
         );
  NOR2_X1 U9575 ( .A1(n7965), .A2(n7916), .ZN(n7918) );
  MUX2_X1 U9576 ( .A(n7898), .B(P2_REG2_REG_12__SCAN_IN), .S(n8570), .Z(n7919)
         );
  INV_X1 U9577 ( .A(n7919), .ZN(n7920) );
  AOI21_X1 U9578 ( .B1(n7921), .B2(n7920), .A(n8530), .ZN(n7922) );
  NOR2_X1 U9579 ( .A1(n7922), .A2(n10023), .ZN(n7923) );
  AOI211_X1 U9580 ( .C1(n10017), .C2(n7925), .A(n7924), .B(n7923), .ZN(n7926)
         );
  OAI21_X1 U9581 ( .B1(n7927), .B2(n9937), .A(n7926), .ZN(P2_U3194) );
  AOI21_X1 U9582 ( .B1(n7929), .B2(n7928), .A(n8470), .ZN(n7936) );
  INV_X1 U9583 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7930) );
  NOR2_X1 U9584 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7930), .ZN(n7948) );
  AOI21_X1 U9585 ( .B1(n8514), .B2(n8523), .A(n7948), .ZN(n7932) );
  NAND2_X1 U9586 ( .A1(n8480), .A2(n8805), .ZN(n7931) );
  OAI211_X1 U9587 ( .C1(n8511), .C2(n7933), .A(n7932), .B(n7931), .ZN(n7934)
         );
  AOI21_X1 U9588 ( .B1(n10071), .B2(n8501), .A(n7934), .ZN(n7935) );
  OAI21_X1 U9589 ( .B1(n7936), .B2(n8503), .A(n7935), .ZN(P2_U3157) );
  AOI21_X1 U9590 ( .B1(n7939), .B2(n7938), .A(n7937), .ZN(n7954) );
  OAI21_X1 U9591 ( .B1(n7942), .B2(n7941), .A(n7940), .ZN(n7952) );
  INV_X1 U9592 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10132) );
  AOI21_X1 U9593 ( .B1(n7945), .B2(n7944), .A(n7943), .ZN(n7946) );
  NOR2_X1 U9594 ( .A1(n7946), .A2(n9937), .ZN(n7947) );
  AOI211_X1 U9595 ( .C1(n7949), .C2(n10008), .A(n7948), .B(n7947), .ZN(n7950)
         );
  OAI21_X1 U9596 ( .B1(n10132), .B2(n9941), .A(n7950), .ZN(n7951) );
  AOI21_X1 U9597 ( .B1(n7952), .B2(n10017), .A(n7951), .ZN(n7953) );
  OAI21_X1 U9598 ( .B1(n7954), .B2(n10023), .A(n7953), .ZN(P2_U3192) );
  OAI21_X1 U9599 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n7956), .A(n7955), .ZN(
        n7971) );
  INV_X1 U9600 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10136) );
  NOR2_X1 U9601 ( .A1(n9941), .A2(n10136), .ZN(n7970) );
  AOI21_X1 U9602 ( .B1(n7958), .B2(n7884), .A(n7957), .ZN(n7968) );
  NAND2_X1 U9603 ( .A1(n7960), .A2(n7959), .ZN(n7963) );
  INV_X1 U9604 ( .A(n7961), .ZN(n7962) );
  NAND2_X1 U9605 ( .A1(n7963), .A2(n7962), .ZN(n7964) );
  INV_X1 U9606 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10254) );
  NOR2_X1 U9607 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10254), .ZN(n8473) );
  AOI21_X1 U9608 ( .B1(n7964), .B2(n10016), .A(n8473), .ZN(n7967) );
  NAND2_X1 U9609 ( .A1(n10008), .A2(n7965), .ZN(n7966) );
  OAI211_X1 U9610 ( .C1(n7968), .C2(n10023), .A(n7967), .B(n7966), .ZN(n7969)
         );
  AOI211_X1 U9611 ( .C1(n7971), .C2(n10017), .A(n7970), .B(n7969), .ZN(n7972)
         );
  INV_X1 U9612 ( .A(n7972), .ZN(P2_U3193) );
  INV_X1 U9613 ( .A(n6198), .ZN(n7974) );
  OAI222_X1 U9614 ( .A1(n9687), .A2(n7975), .B1(n9686), .B2(n7974), .C1(n7973), 
        .C2(P1_U3086), .ZN(P1_U3327) );
  XNOR2_X1 U9615 ( .A(n7976), .B(n8180), .ZN(n7990) );
  INV_X1 U9616 ( .A(n10083), .ZN(n10058) );
  AOI21_X1 U9617 ( .B1(n7977), .B2(n8180), .A(n8831), .ZN(n7980) );
  OAI22_X1 U9618 ( .A1(n6620), .A2(n8755), .B1(n8398), .B2(n8757), .ZN(n7978)
         );
  AOI21_X1 U9619 ( .B1(n7980), .B2(n7979), .A(n7978), .ZN(n7986) );
  INV_X1 U9620 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n7981) );
  MUX2_X1 U9621 ( .A(n7986), .B(n7981), .S(n10086), .Z(n7983) );
  NAND2_X1 U9622 ( .A1(n8391), .A2(n6301), .ZN(n7982) );
  OAI211_X1 U9623 ( .C1(n7990), .C2(n8999), .A(n7983), .B(n7982), .ZN(P2_U3446) );
  MUX2_X1 U9624 ( .A(n7986), .B(n8589), .S(n10098), .Z(n7985) );
  NAND2_X1 U9625 ( .A1(n8391), .A2(n8900), .ZN(n7984) );
  OAI211_X1 U9626 ( .C1(n7990), .C2(n8903), .A(n7985), .B(n7984), .ZN(P2_U3478) );
  MUX2_X1 U9627 ( .A(n7986), .B(n8584), .S(n8812), .Z(n7989) );
  INV_X1 U9628 ( .A(n8389), .ZN(n7987) );
  AOI22_X1 U9629 ( .A1(n8391), .A2(n8813), .B1(n8769), .B2(n7987), .ZN(n7988)
         );
  OAI211_X1 U9630 ( .C1(n7990), .C2(n8816), .A(n7989), .B(n7988), .ZN(P2_U3214) );
  INV_X1 U9631 ( .A(n7991), .ZN(n9685) );
  OAI222_X1 U9632 ( .A1(n9018), .A2(n9685), .B1(n9876), .B2(P2_U3151), .C1(
        n7992), .C2(n9015), .ZN(P2_U3268) );
  OAI21_X1 U9633 ( .B1(n7996), .B2(n7995), .A(n7994), .ZN(n7999) );
  XNOR2_X1 U9634 ( .A(n8620), .B(n7997), .ZN(n7998) );
  XNOR2_X1 U9635 ( .A(n7999), .B(n7998), .ZN(n8004) );
  NOR2_X1 U9636 ( .A1(n8511), .A2(n8629), .ZN(n8002) );
  AOI22_X1 U9637 ( .A1(n8645), .A2(n8514), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8000) );
  OAI21_X1 U9638 ( .B1(n8623), .B2(n8510), .A(n8000), .ZN(n8001) );
  AOI211_X1 U9639 ( .C1(n8913), .C2(n8501), .A(n8002), .B(n8001), .ZN(n8003)
         );
  OAI21_X1 U9640 ( .B1(n8004), .B2(n8503), .A(n8003), .ZN(P2_U3160) );
  NAND2_X1 U9641 ( .A1(n8011), .A2(n8120), .ZN(n8007) );
  OR2_X1 U9642 ( .A1(n8009), .A2(n8356), .ZN(n8006) );
  NAND2_X1 U9643 ( .A1(n8007), .A2(n8006), .ZN(n8008) );
  XNOR2_X1 U9644 ( .A(n8008), .B(n8354), .ZN(n8013) );
  NOR2_X1 U9645 ( .A1(n8009), .A2(n8353), .ZN(n8010) );
  AOI21_X1 U9646 ( .B1(n8011), .B2(n8130), .A(n8010), .ZN(n8012) );
  NAND2_X1 U9647 ( .A1(n8013), .A2(n8012), .ZN(n9131) );
  OR2_X1 U9648 ( .A1(n8013), .A2(n8012), .ZN(n8014) );
  AND2_X1 U9649 ( .A1(n9131), .A2(n8014), .ZN(n9059) );
  NAND2_X1 U9650 ( .A1(n9137), .A2(n8120), .ZN(n8016) );
  OR2_X1 U9651 ( .A1(n8018), .A2(n8356), .ZN(n8015) );
  NAND2_X1 U9652 ( .A1(n8016), .A2(n8015), .ZN(n8017) );
  XNOR2_X1 U9653 ( .A(n8017), .B(n8354), .ZN(n8021) );
  NOR2_X1 U9654 ( .A1(n8018), .A2(n8353), .ZN(n8019) );
  AOI21_X1 U9655 ( .B1(n9137), .B2(n8130), .A(n8019), .ZN(n8020) );
  NAND2_X1 U9656 ( .A1(n8021), .A2(n8020), .ZN(n8023) );
  OR2_X1 U9657 ( .A1(n8021), .A2(n8020), .ZN(n8022) );
  AND2_X1 U9658 ( .A1(n8023), .A2(n8022), .ZN(n9129) );
  OAI22_X1 U9659 ( .A1(n9849), .A2(n8358), .B1(n8025), .B2(n8356), .ZN(n8024)
         );
  XNOR2_X1 U9660 ( .A(n8024), .B(n8354), .ZN(n8028) );
  NAND2_X1 U9661 ( .A1(n8029), .A2(n8028), .ZN(n9020) );
  OR2_X1 U9662 ( .A1(n9849), .A2(n8356), .ZN(n8027) );
  NAND2_X1 U9663 ( .A1(n4922), .A2(n8129), .ZN(n8026) );
  NAND2_X1 U9664 ( .A1(n8027), .A2(n8026), .ZN(n9023) );
  NAND2_X1 U9665 ( .A1(n9020), .A2(n9023), .ZN(n8030) );
  OR2_X2 U9666 ( .A1(n8029), .A2(n8028), .ZN(n9021) );
  NAND2_X1 U9667 ( .A1(n9573), .A2(n8120), .ZN(n8032) );
  NAND2_X1 U9668 ( .A1(n9204), .A2(n8130), .ZN(n8031) );
  NAND2_X1 U9669 ( .A1(n8032), .A2(n8031), .ZN(n8033) );
  XNOR2_X1 U9670 ( .A(n8033), .B(n8128), .ZN(n9176) );
  NAND2_X1 U9671 ( .A1(n9573), .A2(n8130), .ZN(n8035) );
  NAND2_X1 U9672 ( .A1(n9204), .A2(n8129), .ZN(n8034) );
  NAND2_X1 U9673 ( .A1(n8035), .A2(n8034), .ZN(n9177) );
  NAND2_X1 U9674 ( .A1(n9548), .A2(n8120), .ZN(n8037) );
  NAND2_X1 U9675 ( .A1(n9203), .A2(n8130), .ZN(n8036) );
  NAND2_X1 U9676 ( .A1(n8037), .A2(n8036), .ZN(n8038) );
  XNOR2_X1 U9677 ( .A(n8038), .B(n8354), .ZN(n8040) );
  NOR2_X1 U9678 ( .A1(n9092), .A2(n8353), .ZN(n8039) );
  AOI21_X1 U9679 ( .B1(n9548), .B2(n8130), .A(n8039), .ZN(n8041) );
  NAND2_X1 U9680 ( .A1(n8040), .A2(n8041), .ZN(n8046) );
  INV_X1 U9681 ( .A(n8040), .ZN(n8043) );
  INV_X1 U9682 ( .A(n8041), .ZN(n8042) );
  NAND2_X1 U9683 ( .A1(n8043), .A2(n8042), .ZN(n8044) );
  NAND2_X1 U9684 ( .A1(n8046), .A2(n8044), .ZN(n9080) );
  NAND2_X1 U9685 ( .A1(n9536), .A2(n8120), .ZN(n8048) );
  NAND2_X1 U9686 ( .A1(n9202), .A2(n8130), .ZN(n8047) );
  NAND2_X1 U9687 ( .A1(n8048), .A2(n8047), .ZN(n8049) );
  XNOR2_X1 U9688 ( .A(n8049), .B(n8128), .ZN(n8051) );
  AND2_X1 U9689 ( .A1(n9202), .A2(n8129), .ZN(n8050) );
  AOI21_X1 U9690 ( .B1(n9536), .B2(n8130), .A(n8050), .ZN(n8052) );
  XNOR2_X1 U9691 ( .A(n8051), .B(n8052), .ZN(n9088) );
  INV_X1 U9692 ( .A(n8051), .ZN(n8053) );
  NAND2_X1 U9693 ( .A1(n8053), .A2(n8052), .ZN(n8054) );
  NAND2_X1 U9694 ( .A1(n9632), .A2(n8120), .ZN(n8056) );
  NAND2_X1 U9695 ( .A1(n9201), .A2(n8130), .ZN(n8055) );
  NAND2_X1 U9696 ( .A1(n8056), .A2(n8055), .ZN(n8057) );
  XNOR2_X1 U9697 ( .A(n8057), .B(n8354), .ZN(n8059) );
  AND2_X1 U9698 ( .A1(n9201), .A2(n8129), .ZN(n8058) );
  AOI21_X1 U9699 ( .B1(n9632), .B2(n8130), .A(n8058), .ZN(n9153) );
  NAND2_X1 U9700 ( .A1(n9154), .A2(n9153), .ZN(n9152) );
  NAND2_X1 U9701 ( .A1(n9628), .A2(n8120), .ZN(n8062) );
  NAND2_X1 U9702 ( .A1(n9200), .A2(n8130), .ZN(n8061) );
  NAND2_X1 U9703 ( .A1(n8062), .A2(n8061), .ZN(n8063) );
  XNOR2_X1 U9704 ( .A(n8063), .B(n8128), .ZN(n8065) );
  AND2_X1 U9705 ( .A1(n9200), .A2(n8129), .ZN(n8064) );
  AOI21_X1 U9706 ( .B1(n9628), .B2(n6915), .A(n8064), .ZN(n8066) );
  XNOR2_X1 U9707 ( .A(n8065), .B(n8066), .ZN(n9042) );
  INV_X1 U9708 ( .A(n8065), .ZN(n8067) );
  NAND2_X1 U9709 ( .A1(n8067), .A2(n8066), .ZN(n8068) );
  NAND2_X1 U9710 ( .A1(n9623), .A2(n8120), .ZN(n8070) );
  NAND2_X1 U9711 ( .A1(n9199), .A2(n8130), .ZN(n8069) );
  NAND2_X1 U9712 ( .A1(n8070), .A2(n8069), .ZN(n8071) );
  XNOR2_X1 U9713 ( .A(n8071), .B(n8354), .ZN(n8073) );
  AND2_X1 U9714 ( .A1(n9199), .A2(n8129), .ZN(n8072) );
  AOI21_X1 U9715 ( .B1(n9623), .B2(n6915), .A(n8072), .ZN(n8074) );
  AND2_X1 U9716 ( .A1(n8073), .A2(n8074), .ZN(n9115) );
  INV_X1 U9717 ( .A(n8073), .ZN(n8076) );
  INV_X1 U9718 ( .A(n8074), .ZN(n8075) );
  NAND2_X1 U9719 ( .A1(n8076), .A2(n8075), .ZN(n9116) );
  NAND2_X1 U9720 ( .A1(n9478), .A2(n8120), .ZN(n8078) );
  NAND2_X1 U9721 ( .A1(n9198), .A2(n8130), .ZN(n8077) );
  NAND2_X1 U9722 ( .A1(n8078), .A2(n8077), .ZN(n8079) );
  XNOR2_X1 U9723 ( .A(n8079), .B(n8128), .ZN(n9049) );
  INV_X1 U9724 ( .A(n9049), .ZN(n8082) );
  NAND2_X1 U9725 ( .A1(n9478), .A2(n8130), .ZN(n8081) );
  NAND2_X1 U9726 ( .A1(n9198), .A2(n8129), .ZN(n8080) );
  NAND2_X1 U9727 ( .A1(n8081), .A2(n8080), .ZN(n8086) );
  INV_X1 U9728 ( .A(n8086), .ZN(n9048) );
  NAND2_X1 U9729 ( .A1(n8082), .A2(n9048), .ZN(n8090) );
  NAND2_X1 U9730 ( .A1(n9612), .A2(n8120), .ZN(n8084) );
  NAND2_X1 U9731 ( .A1(n9197), .A2(n8130), .ZN(n8083) );
  NAND2_X1 U9732 ( .A1(n8084), .A2(n8083), .ZN(n8085) );
  XNOR2_X1 U9733 ( .A(n8085), .B(n8128), .ZN(n8091) );
  AND2_X1 U9734 ( .A1(n9049), .A2(n8086), .ZN(n8089) );
  AND2_X1 U9735 ( .A1(n9197), .A2(n8129), .ZN(n8088) );
  AOI21_X1 U9736 ( .B1(n9612), .B2(n6915), .A(n8088), .ZN(n9140) );
  NOR2_X2 U9737 ( .A1(n9141), .A2(n9140), .ZN(n9139) );
  INV_X1 U9738 ( .A(n9051), .ZN(n8094) );
  INV_X1 U9739 ( .A(n8089), .ZN(n8093) );
  NAND2_X1 U9740 ( .A1(n8091), .A2(n8090), .ZN(n8092) );
  NAND2_X1 U9741 ( .A1(n9608), .A2(n8120), .ZN(n8096) );
  NAND2_X1 U9742 ( .A1(n9145), .A2(n8130), .ZN(n8095) );
  NAND2_X1 U9743 ( .A1(n8096), .A2(n8095), .ZN(n8097) );
  XNOR2_X1 U9744 ( .A(n8097), .B(n8354), .ZN(n8099) );
  AND2_X1 U9745 ( .A1(n9145), .A2(n8129), .ZN(n8098) );
  AOI21_X1 U9746 ( .B1(n9608), .B2(n6915), .A(n8098), .ZN(n8100) );
  NAND2_X1 U9747 ( .A1(n8099), .A2(n8100), .ZN(n9103) );
  INV_X1 U9748 ( .A(n8099), .ZN(n8102) );
  INV_X1 U9749 ( .A(n8100), .ZN(n8101) );
  NAND2_X1 U9750 ( .A1(n8102), .A2(n8101), .ZN(n8103) );
  NAND2_X1 U9751 ( .A1(n9103), .A2(n8103), .ZN(n9035) );
  NAND2_X1 U9752 ( .A1(n9601), .A2(n8120), .ZN(n8105) );
  OR2_X1 U9753 ( .A1(n9071), .A2(n8356), .ZN(n8104) );
  NAND2_X1 U9754 ( .A1(n8105), .A2(n8104), .ZN(n8106) );
  XNOR2_X1 U9755 ( .A(n8106), .B(n8354), .ZN(n8109) );
  NOR2_X1 U9756 ( .A1(n9071), .A2(n8353), .ZN(n8107) );
  AOI21_X1 U9757 ( .B1(n9601), .B2(n6915), .A(n8107), .ZN(n8108) );
  NAND2_X1 U9758 ( .A1(n8109), .A2(n8108), .ZN(n8111) );
  OR2_X1 U9759 ( .A1(n8109), .A2(n8108), .ZN(n8110) );
  NAND2_X1 U9760 ( .A1(n8111), .A2(n8110), .ZN(n9102) );
  INV_X1 U9761 ( .A(n8111), .ZN(n8112) );
  NAND2_X1 U9762 ( .A1(n9418), .A2(n8120), .ZN(n8114) );
  NAND2_X1 U9763 ( .A1(n9195), .A2(n8130), .ZN(n8113) );
  NAND2_X1 U9764 ( .A1(n8114), .A2(n8113), .ZN(n8115) );
  XNOR2_X1 U9765 ( .A(n8115), .B(n8128), .ZN(n8118) );
  OAI22_X1 U9766 ( .A1(n9658), .A2(n8356), .B1(n8116), .B2(n8353), .ZN(n8117)
         );
  XNOR2_X1 U9767 ( .A(n8118), .B(n8117), .ZN(n9069) );
  NOR2_X1 U9768 ( .A1(n8118), .A2(n8117), .ZN(n9166) );
  NOR2_X1 U9769 ( .A1(n9072), .A2(n8353), .ZN(n8119) );
  AOI21_X1 U9770 ( .B1(n9402), .B2(n8130), .A(n8119), .ZN(n8124) );
  NAND2_X1 U9771 ( .A1(n9402), .A2(n8120), .ZN(n8122) );
  OR2_X1 U9772 ( .A1(n9072), .A2(n8356), .ZN(n8121) );
  NAND2_X1 U9773 ( .A1(n8122), .A2(n8121), .ZN(n8123) );
  XNOR2_X1 U9774 ( .A(n8123), .B(n8128), .ZN(n8126) );
  XOR2_X1 U9775 ( .A(n8124), .B(n8126), .Z(n9165) );
  INV_X1 U9776 ( .A(n8124), .ZN(n8125) );
  OAI22_X1 U9777 ( .A1(n5748), .A2(n8358), .B1(n9169), .B2(n8356), .ZN(n8127)
         );
  XOR2_X1 U9778 ( .A(n8128), .B(n8127), .Z(n8132) );
  INV_X1 U9779 ( .A(n9169), .ZN(n9193) );
  AOI22_X1 U9780 ( .A1(n9390), .A2(n8130), .B1(n8129), .B2(n9193), .ZN(n8131)
         );
  NAND2_X1 U9781 ( .A1(n8132), .A2(n8131), .ZN(n8364) );
  OAI21_X1 U9782 ( .B1(n8132), .B2(n8131), .A(n8364), .ZN(n8133) );
  OR2_X1 U9783 ( .A1(n8357), .A2(n9168), .ZN(n8135) );
  OR2_X1 U9784 ( .A1(n9072), .A2(n9091), .ZN(n8134) );
  AND2_X1 U9785 ( .A1(n8135), .A2(n8134), .ZN(n9382) );
  INV_X1 U9786 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8136) );
  OAI22_X1 U9787 ( .A1(n9382), .A2(n9694), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8136), .ZN(n8137) );
  AOI21_X1 U9788 ( .B1(n9389), .B2(n9187), .A(n8137), .ZN(n8138) );
  OAI211_X1 U9789 ( .C1(n5748), .C2(n9722), .A(n8139), .B(n8138), .ZN(P1_U3214) );
  INV_X1 U9790 ( .A(n8146), .ZN(n9008) );
  OAI222_X1 U9791 ( .A1(n9687), .A2(n8141), .B1(n9689), .B2(n9008), .C1(n8140), 
        .C2(P1_U3086), .ZN(P1_U3325) );
  INV_X1 U9792 ( .A(n8142), .ZN(n9683) );
  OAI222_X1 U9793 ( .A1(n9018), .A2(n9683), .B1(P2_U3151), .B2(n8144), .C1(
        n8143), .C2(n9015), .ZN(P2_U3266) );
  NOR2_X1 U9794 ( .A1(n5905), .A2(n9009), .ZN(n8145) );
  AND2_X1 U9795 ( .A1(n8910), .A2(n8519), .ZN(n8334) );
  INV_X1 U9796 ( .A(n8907), .ZN(n8837) );
  INV_X1 U9797 ( .A(n8605), .ZN(n8149) );
  NAND2_X1 U9798 ( .A1(n8837), .A2(n8149), .ZN(n8340) );
  INV_X1 U9799 ( .A(n8150), .ZN(n8151) );
  NAND2_X1 U9800 ( .A1(n8151), .A2(n8328), .ZN(n8157) );
  OR2_X1 U9801 ( .A1(n8910), .A2(n8519), .ZN(n8335) );
  NAND2_X1 U9802 ( .A1(n8907), .A2(n8605), .ZN(n8338) );
  INV_X1 U9803 ( .A(n8335), .ZN(n8189) );
  INV_X1 U9804 ( .A(n8319), .ZN(n8158) );
  NAND2_X1 U9805 ( .A1(n8305), .A2(n8308), .ZN(n8670) );
  INV_X1 U9806 ( .A(n8693), .ZN(n8689) );
  INV_X1 U9807 ( .A(n8703), .ZN(n8183) );
  INV_X1 U9808 ( .A(n8741), .ZN(n8742) );
  INV_X1 U9809 ( .A(n8269), .ZN(n8159) );
  INV_X1 U9810 ( .A(n8264), .ZN(n8160) );
  OR2_X1 U9811 ( .A1(n8263), .A2(n8160), .ZN(n8259) );
  INV_X1 U9812 ( .A(n8798), .ZN(n8803) );
  AND2_X1 U9813 ( .A1(n8162), .A2(n8161), .ZN(n8164) );
  NAND4_X1 U9814 ( .A1(n7052), .A2(n8165), .A3(n8164), .A4(n8163), .ZN(n8167)
         );
  NOR2_X1 U9815 ( .A1(n8167), .A2(n8166), .ZN(n8171) );
  NOR2_X1 U9816 ( .A1(n8168), .A2(n8204), .ZN(n8169) );
  NAND4_X1 U9817 ( .A1(n8171), .A2(n8170), .A3(n8169), .A4(n4665), .ZN(n8174)
         );
  NOR3_X1 U9818 ( .A1(n8174), .A2(n8173), .A3(n8172), .ZN(n8175) );
  NAND3_X1 U9819 ( .A1(n8803), .A2(n8176), .A3(n8175), .ZN(n8177) );
  OR4_X1 U9820 ( .A1(n8781), .A2(n8270), .A3(n8259), .A4(n8177), .ZN(n8178) );
  NOR2_X1 U9821 ( .A1(n8752), .A2(n8178), .ZN(n8179) );
  NAND4_X1 U9822 ( .A1(n8180), .A2(n8742), .A3(n4515), .A4(n8179), .ZN(n8181)
         );
  NOR2_X1 U9823 ( .A1(n8716), .A2(n8181), .ZN(n8182) );
  NAND3_X1 U9824 ( .A1(n8689), .A2(n8183), .A3(n8182), .ZN(n8184) );
  NAND2_X1 U9825 ( .A1(n8665), .A2(n8666), .ZN(n8680) );
  OR4_X1 U9826 ( .A1(n8656), .A2(n8670), .A3(n8184), .A4(n8680), .ZN(n8185) );
  NOR2_X1 U9827 ( .A1(n8313), .A2(n8185), .ZN(n8186) );
  INV_X1 U9828 ( .A(n8634), .ZN(n8321) );
  NAND3_X1 U9829 ( .A1(n8620), .A2(n8186), .A3(n8321), .ZN(n8187) );
  NOR4_X1 U9830 ( .A1(n8189), .A2(n8334), .A3(n8188), .A4(n8187), .ZN(n8190)
         );
  MUX2_X1 U9831 ( .A(n8645), .B(n8919), .S(n8326), .Z(n8322) );
  INV_X1 U9832 ( .A(n8193), .ZN(n8299) );
  AND2_X1 U9833 ( .A1(n8193), .A2(n8192), .ZN(n8295) );
  INV_X1 U9834 ( .A(n8273), .ZN(n8194) );
  NOR2_X1 U9835 ( .A1(n8741), .A2(n8194), .ZN(n8275) );
  INV_X1 U9836 ( .A(n6237), .ZN(n8205) );
  OAI21_X1 U9837 ( .B1(n8196), .B2(n8195), .A(n8200), .ZN(n8198) );
  INV_X1 U9838 ( .A(n8199), .ZN(n8197) );
  AOI211_X1 U9839 ( .C1(n8198), .C2(n6237), .A(n8336), .B(n8197), .ZN(n8202)
         );
  AOI21_X1 U9840 ( .B1(n8200), .B2(n8199), .A(n8326), .ZN(n8201) );
  NOR2_X1 U9841 ( .A1(n8202), .A2(n8201), .ZN(n8203) );
  AOI211_X1 U9842 ( .C1(n8205), .C2(n8336), .A(n8204), .B(n8203), .ZN(n8215)
         );
  NAND2_X1 U9843 ( .A1(n8223), .A2(n8206), .ZN(n8210) );
  NAND2_X1 U9844 ( .A1(n8207), .A2(n10028), .ZN(n8208) );
  NAND2_X1 U9845 ( .A1(n8216), .A2(n8208), .ZN(n8209) );
  MUX2_X1 U9846 ( .A(n8210), .B(n8209), .S(n8336), .Z(n8214) );
  NAND2_X1 U9847 ( .A1(n8212), .A2(n8211), .ZN(n8224) );
  MUX2_X1 U9848 ( .A(n8219), .B(n8224), .S(n8326), .Z(n8213) );
  OAI21_X1 U9849 ( .B1(n8215), .B2(n8214), .A(n8213), .ZN(n8227) );
  INV_X1 U9850 ( .A(n8216), .ZN(n8220) );
  NAND2_X1 U9851 ( .A1(n8218), .A2(n8217), .ZN(n8228) );
  OAI211_X1 U9852 ( .C1(n8227), .C2(n8220), .A(n8228), .B(n8219), .ZN(n8221)
         );
  NAND2_X1 U9853 ( .A1(n8527), .A2(n10044), .ZN(n8225) );
  NAND3_X1 U9854 ( .A1(n8221), .A2(n8231), .A3(n8225), .ZN(n8222) );
  INV_X1 U9855 ( .A(n8223), .ZN(n8226) );
  OAI211_X1 U9856 ( .C1(n8227), .C2(n8226), .A(n8225), .B(n8224), .ZN(n8230)
         );
  NAND3_X1 U9857 ( .A1(n8230), .A2(n8229), .A3(n8228), .ZN(n8232) );
  NAND2_X1 U9858 ( .A1(n8233), .A2(n8240), .ZN(n8235) );
  NAND2_X1 U9859 ( .A1(n8244), .A2(n8243), .ZN(n8234) );
  MUX2_X1 U9860 ( .A(n8235), .B(n8234), .S(n8326), .Z(n8246) );
  INV_X1 U9861 ( .A(n8237), .ZN(n8238) );
  NOR2_X1 U9862 ( .A1(n8239), .A2(n8238), .ZN(n8241) );
  OAI211_X1 U9863 ( .C1(n8246), .C2(n8241), .A(n8240), .B(n8253), .ZN(n8248)
         );
  OR2_X1 U9864 ( .A1(n8525), .A2(n10053), .ZN(n8242) );
  AND2_X1 U9865 ( .A1(n8243), .A2(n8242), .ZN(n8245) );
  OAI211_X1 U9866 ( .C1(n8246), .C2(n8245), .A(n8250), .B(n8244), .ZN(n8247)
         );
  MUX2_X1 U9867 ( .A(n8248), .B(n8247), .S(n8336), .Z(n8249) );
  INV_X1 U9868 ( .A(n8257), .ZN(n8251) );
  NAND2_X1 U9869 ( .A1(n8251), .A2(n8250), .ZN(n8252) );
  NAND2_X1 U9870 ( .A1(n8254), .A2(n8253), .ZN(n8256) );
  OAI21_X1 U9871 ( .B1(n8257), .B2(n8256), .A(n8255), .ZN(n8258) );
  MUX2_X1 U9872 ( .A(n8261), .B(n8260), .S(n8326), .Z(n8262) );
  MUX2_X1 U9873 ( .A(n8264), .B(n4813), .S(n8326), .Z(n8265) );
  INV_X1 U9874 ( .A(n8267), .ZN(n8268) );
  MUX2_X1 U9875 ( .A(n8269), .B(n8268), .S(n8336), .Z(n8271) );
  INV_X1 U9876 ( .A(n8276), .ZN(n8280) );
  INV_X1 U9877 ( .A(n8277), .ZN(n8279) );
  OAI211_X1 U9878 ( .C1(n8280), .C2(n8279), .A(n8326), .B(n8278), .ZN(n8284)
         );
  INV_X1 U9879 ( .A(n8281), .ZN(n8283) );
  INV_X1 U9880 ( .A(n8286), .ZN(n8282) );
  AOI211_X1 U9881 ( .C1(n8287), .C2(n8284), .A(n8283), .B(n8282), .ZN(n8293)
         );
  NAND2_X1 U9882 ( .A1(n8290), .A2(n8285), .ZN(n8288) );
  MUX2_X1 U9883 ( .A(n8290), .B(n8289), .S(n8326), .Z(n8291) );
  OAI211_X1 U9884 ( .C1(n8293), .C2(n8292), .A(n8296), .B(n8291), .ZN(n8294)
         );
  AOI21_X1 U9885 ( .B1(n8298), .B2(n8296), .A(n8336), .ZN(n8297) );
  INV_X1 U9886 ( .A(n8300), .ZN(n8303) );
  NAND2_X1 U9887 ( .A1(n8666), .A2(n8301), .ZN(n8302) );
  MUX2_X1 U9888 ( .A(n8303), .B(n8302), .S(n8326), .Z(n8304) );
  NAND2_X1 U9889 ( .A1(n8305), .A2(n8665), .ZN(n8307) );
  MUX2_X1 U9890 ( .A(n8307), .B(n8306), .S(n8336), .Z(n8311) );
  INV_X1 U9891 ( .A(n8656), .ZN(n8654) );
  MUX2_X1 U9892 ( .A(n8309), .B(n8308), .S(n8326), .Z(n8310) );
  OAI211_X1 U9893 ( .C1(n8312), .C2(n8311), .A(n8654), .B(n8310), .ZN(n8317)
         );
  MUX2_X1 U9894 ( .A(n8315), .B(n8314), .S(n8336), .Z(n8316) );
  MUX2_X1 U9895 ( .A(n8319), .B(n6252), .S(n8336), .Z(n8320) );
  NAND2_X1 U9896 ( .A1(n8324), .A2(n8336), .ZN(n8325) );
  INV_X1 U9897 ( .A(n8623), .ZN(n8520) );
  AOI22_X1 U9898 ( .A1(n8328), .A2(n8325), .B1(n8336), .B2(n8520), .ZN(n8332)
         );
  MUX2_X1 U9899 ( .A(n6209), .B(n6210), .S(n8326), .Z(n8331) );
  INV_X1 U9900 ( .A(n8337), .ZN(n8329) );
  INV_X1 U9901 ( .A(n8334), .ZN(n8327) );
  NAND4_X1 U9902 ( .A1(n8329), .A2(n8336), .A3(n8328), .A4(n8327), .ZN(n8342)
         );
  OAI21_X1 U9903 ( .B1(n8333), .B2(n4766), .A(n4767), .ZN(n8339) );
  AOI21_X1 U9904 ( .B1(n8336), .B2(n8335), .A(n8334), .ZN(n8341) );
  XNOR2_X1 U9905 ( .A(n8345), .B(n8344), .ZN(n8352) );
  NOR3_X1 U9906 ( .A1(n8347), .A2(n8346), .A3(n6226), .ZN(n8350) );
  OAI21_X1 U9907 ( .B1(n8351), .B2(n8348), .A(P2_B_REG_SCAN_IN), .ZN(n8349) );
  OAI22_X1 U9908 ( .A1(n8352), .A2(n8351), .B1(n8350), .B2(n8349), .ZN(
        P2_U3296) );
  OAI22_X1 U9909 ( .A1(n4510), .A2(n8356), .B1(n8357), .B2(n8353), .ZN(n8355)
         );
  XNOR2_X1 U9910 ( .A(n8355), .B(n8354), .ZN(n8360) );
  OAI22_X1 U9911 ( .A1(n4510), .A2(n8358), .B1(n8357), .B2(n8356), .ZN(n8359)
         );
  XNOR2_X1 U9912 ( .A(n8360), .B(n8359), .ZN(n8361) );
  INV_X1 U9913 ( .A(n8361), .ZN(n8365) );
  NAND3_X1 U9914 ( .A1(n8365), .A2(n9724), .A3(n8364), .ZN(n8371) );
  NAND3_X1 U9915 ( .A1(n4551), .A2(n9724), .A3(n8361), .ZN(n8370) );
  INV_X1 U9916 ( .A(n9375), .ZN(n8363) );
  AOI22_X1 U9917 ( .A1(n4585), .A2(n9719), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n8362) );
  OAI21_X1 U9918 ( .B1(n8363), .B2(n9727), .A(n8362), .ZN(n8367) );
  NOR3_X1 U9919 ( .A1(n8365), .A2(n8364), .A3(n9699), .ZN(n8366) );
  AOI211_X1 U9920 ( .C1(n8368), .C2(n9703), .A(n8367), .B(n8366), .ZN(n8369)
         );
  OAI211_X1 U9921 ( .C1(n4551), .C2(n8371), .A(n8370), .B(n8369), .ZN(P1_U3220) );
  XOR2_X1 U9922 ( .A(n8373), .B(n8372), .Z(n8378) );
  AOI22_X1 U9923 ( .A1(n8480), .A2(n8774), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n8375) );
  NAND2_X1 U9924 ( .A1(n8514), .A2(n8806), .ZN(n8374) );
  OAI211_X1 U9925 ( .C1(n8511), .C2(n8776), .A(n8375), .B(n8374), .ZN(n8376)
         );
  AOI21_X1 U9926 ( .B1(n8984), .B2(n8501), .A(n8376), .ZN(n8377) );
  OAI21_X1 U9927 ( .B1(n8378), .B2(n8503), .A(n8377), .ZN(P2_U3155) );
  XNOR2_X1 U9928 ( .A(n8379), .B(n8672), .ZN(n8384) );
  NAND2_X1 U9929 ( .A1(n8497), .A2(n8685), .ZN(n8381) );
  AOI22_X1 U9930 ( .A1(n8514), .A2(n8704), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8380) );
  OAI211_X1 U9931 ( .C1(n8414), .C2(n8510), .A(n8381), .B(n8380), .ZN(n8382)
         );
  AOI21_X1 U9932 ( .B1(n8943), .B2(n8501), .A(n8382), .ZN(n8383) );
  OAI21_X1 U9933 ( .B1(n8384), .B2(n8503), .A(n8383), .ZN(P2_U3156) );
  XOR2_X1 U9934 ( .A(n8385), .B(n8386), .Z(n8393) );
  AOI22_X1 U9935 ( .A1(n8480), .A2(n8705), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3151), .ZN(n8388) );
  NAND2_X1 U9936 ( .A1(n8514), .A2(n8744), .ZN(n8387) );
  OAI211_X1 U9937 ( .C1(n8511), .C2(n8389), .A(n8388), .B(n8387), .ZN(n8390)
         );
  AOI21_X1 U9938 ( .B1(n8391), .B2(n8501), .A(n8390), .ZN(n8392) );
  OAI21_X1 U9939 ( .B1(n8393), .B2(n8503), .A(n8392), .ZN(P2_U3159) );
  XOR2_X1 U9940 ( .A(n8395), .B(n8394), .Z(n8401) );
  NAND2_X1 U9941 ( .A1(n8497), .A2(n8708), .ZN(n8397) );
  AOI22_X1 U9942 ( .A1(n8480), .A2(n8704), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8396) );
  OAI211_X1 U9943 ( .C1(n8398), .C2(n8476), .A(n8397), .B(n8396), .ZN(n8399)
         );
  AOI21_X1 U9944 ( .B1(n8953), .B2(n8501), .A(n8399), .ZN(n8400) );
  OAI21_X1 U9945 ( .B1(n8401), .B2(n8503), .A(n8400), .ZN(P2_U3163) );
  XNOR2_X1 U9946 ( .A(n4586), .B(n8402), .ZN(n8409) );
  NOR2_X1 U9947 ( .A1(n8476), .A2(n8403), .ZN(n8404) );
  AOI211_X1 U9948 ( .C1(n8480), .C2(n8806), .A(n8405), .B(n8404), .ZN(n8406)
         );
  OAI21_X1 U9949 ( .B1(n8809), .B2(n8511), .A(n8406), .ZN(n8407) );
  AOI21_X1 U9950 ( .B1(n8996), .B2(n8501), .A(n8407), .ZN(n8408) );
  OAI21_X1 U9951 ( .B1(n8409), .B2(n8503), .A(n8408), .ZN(P2_U3164) );
  XOR2_X1 U9952 ( .A(n8411), .B(n8410), .Z(n8417) );
  AOI22_X1 U9953 ( .A1(n8658), .A2(n8480), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8413) );
  NAND2_X1 U9954 ( .A1(n8497), .A2(n8662), .ZN(n8412) );
  OAI211_X1 U9955 ( .C1(n8414), .C2(n8476), .A(n8413), .B(n8412), .ZN(n8415)
         );
  AOI21_X1 U9956 ( .B1(n8931), .B2(n8501), .A(n8415), .ZN(n8416) );
  OAI21_X1 U9957 ( .B1(n8417), .B2(n8503), .A(n8416), .ZN(P2_U3165) );
  INV_X1 U9958 ( .A(n8887), .ZN(n8426) );
  OAI211_X1 U9959 ( .C1(n8420), .C2(n8419), .A(n8418), .B(n8505), .ZN(n8425)
         );
  NAND2_X1 U9960 ( .A1(n8514), .A2(n8774), .ZN(n8421) );
  NAND2_X1 U9961 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n10004) );
  OAI211_X1 U9962 ( .C1(n8756), .C2(n8510), .A(n8421), .B(n10004), .ZN(n8422)
         );
  AOI21_X1 U9963 ( .B1(n8423), .B2(n8497), .A(n8422), .ZN(n8424) );
  OAI211_X1 U9964 ( .C1(n8426), .C2(n8517), .A(n8425), .B(n8424), .ZN(P2_U3166) );
  AOI21_X1 U9965 ( .B1(n8428), .B2(n8427), .A(n4582), .ZN(n8435) );
  OAI22_X1 U9966 ( .A1(n8510), .A2(n6620), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8429), .ZN(n8430) );
  AOI21_X1 U9967 ( .B1(n8514), .B2(n8766), .A(n8430), .ZN(n8431) );
  OAI21_X1 U9968 ( .B1(n8432), .B2(n8511), .A(n8431), .ZN(n8433) );
  AOI21_X1 U9969 ( .B1(n8968), .B2(n8501), .A(n8433), .ZN(n8434) );
  OAI21_X1 U9970 ( .B1(n8435), .B2(n8503), .A(n8434), .ZN(P2_U3168) );
  XOR2_X1 U9971 ( .A(n8437), .B(n8436), .Z(n8442) );
  AOI22_X1 U9972 ( .A1(n8671), .A2(n8480), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8439) );
  NAND2_X1 U9973 ( .A1(n8497), .A2(n8676), .ZN(n8438) );
  OAI211_X1 U9974 ( .C1(n8692), .C2(n8476), .A(n8439), .B(n8438), .ZN(n8440)
         );
  AOI21_X1 U9975 ( .B1(n8937), .B2(n8501), .A(n8440), .ZN(n8441) );
  OAI21_X1 U9976 ( .B1(n8442), .B2(n8503), .A(n8441), .ZN(P2_U3169) );
  XOR2_X1 U9977 ( .A(n8443), .B(n8444), .Z(n8449) );
  NAND2_X1 U9978 ( .A1(n8497), .A2(n8722), .ZN(n8446) );
  AOI22_X1 U9979 ( .A1(n8480), .A2(n8718), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8445) );
  OAI211_X1 U9980 ( .C1(n8729), .C2(n8476), .A(n8446), .B(n8445), .ZN(n8447)
         );
  AOI21_X1 U9981 ( .B1(n8874), .B2(n8501), .A(n8447), .ZN(n8448) );
  OAI21_X1 U9982 ( .B1(n8449), .B2(n8503), .A(n8448), .ZN(P2_U3173) );
  NOR2_X1 U9983 ( .A1(n8450), .A2(n4587), .ZN(n8451) );
  XNOR2_X1 U9984 ( .A(n8452), .B(n8451), .ZN(n8459) );
  NAND2_X1 U9985 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9954) );
  INV_X1 U9986 ( .A(n9954), .ZN(n8455) );
  NOR2_X1 U9987 ( .A1(n8476), .A2(n8453), .ZN(n8454) );
  AOI211_X1 U9988 ( .C1(n8480), .C2(n8787), .A(n8455), .B(n8454), .ZN(n8456)
         );
  OAI21_X1 U9989 ( .B1(n8789), .B2(n8511), .A(n8456), .ZN(n8457) );
  AOI21_X1 U9990 ( .B1(n8990), .B2(n8501), .A(n8457), .ZN(n8458) );
  OAI21_X1 U9991 ( .B1(n8459), .B2(n8503), .A(n8458), .ZN(P2_U3174) );
  XOR2_X1 U9992 ( .A(n8461), .B(n8460), .Z(n8466) );
  NAND2_X1 U9993 ( .A1(n8497), .A2(n8696), .ZN(n8463) );
  AOI22_X1 U9994 ( .A1(n8514), .A2(n8718), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8462) );
  OAI211_X1 U9995 ( .C1(n8692), .C2(n8510), .A(n8463), .B(n8462), .ZN(n8464)
         );
  AOI21_X1 U9996 ( .B1(n8695), .B2(n8501), .A(n8464), .ZN(n8465) );
  OAI21_X1 U9997 ( .B1(n8466), .B2(n8503), .A(n8465), .ZN(P2_U3175) );
  INV_X1 U9998 ( .A(n8467), .ZN(n8472) );
  OAI21_X1 U9999 ( .B1(n8470), .B2(n8469), .A(n8468), .ZN(n8471) );
  NAND3_X1 U10000 ( .A1(n8472), .A2(n8505), .A3(n8471), .ZN(n8482) );
  INV_X1 U10001 ( .A(n8473), .ZN(n8474) );
  OAI21_X1 U10002 ( .B1(n8476), .B2(n8475), .A(n8474), .ZN(n8479) );
  NOR2_X1 U10003 ( .A1(n8511), .A2(n8477), .ZN(n8478) );
  AOI211_X1 U10004 ( .C1(n8480), .C2(n8786), .A(n8479), .B(n8478), .ZN(n8481)
         );
  OAI211_X1 U10005 ( .C1(n10079), .C2(n8517), .A(n8482), .B(n8481), .ZN(
        P2_U3176) );
  INV_X1 U10006 ( .A(n8484), .ZN(n8488) );
  NOR3_X1 U10007 ( .A1(n4582), .A2(n8486), .A3(n8485), .ZN(n8487) );
  OAI21_X1 U10008 ( .B1(n8488), .B2(n8487), .A(n8505), .ZN(n8492) );
  NAND2_X1 U10009 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8565) );
  OAI21_X1 U10010 ( .B1(n8510), .B2(n8729), .A(n8565), .ZN(n8490) );
  NOR2_X1 U10011 ( .A1(n8511), .A2(n8734), .ZN(n8489) );
  AOI211_X1 U10012 ( .C1(n8514), .C2(n8521), .A(n8490), .B(n8489), .ZN(n8491)
         );
  OAI211_X1 U10013 ( .C1(n8965), .C2(n8517), .A(n8492), .B(n8491), .ZN(
        P2_U3178) );
  NAND2_X1 U10014 ( .A1(n8495), .A2(n8494), .ZN(n8496) );
  XNOR2_X1 U10015 ( .A(n8493), .B(n8496), .ZN(n8504) );
  AOI22_X1 U10016 ( .A1(n8671), .A2(n8514), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8499) );
  NAND2_X1 U10017 ( .A1(n8497), .A2(n8651), .ZN(n8498) );
  OAI211_X1 U10018 ( .C1(n8622), .C2(n8510), .A(n8499), .B(n8498), .ZN(n8500)
         );
  AOI21_X1 U10019 ( .B1(n8925), .B2(n8501), .A(n8500), .ZN(n8502) );
  OAI21_X1 U10020 ( .B1(n8504), .B2(n8503), .A(n8502), .ZN(P2_U3180) );
  INV_X1 U10021 ( .A(n8978), .ZN(n8518) );
  OAI211_X1 U10022 ( .C1(n8508), .C2(n8507), .A(n8506), .B(n8505), .ZN(n8516)
         );
  NAND2_X1 U10023 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9987) );
  OAI21_X1 U10024 ( .B1(n8510), .B2(n8509), .A(n9987), .ZN(n8513) );
  NOR2_X1 U10025 ( .A1(n8511), .A2(n8768), .ZN(n8512) );
  AOI211_X1 U10026 ( .C1(n8514), .C2(n8787), .A(n8513), .B(n8512), .ZN(n8515)
         );
  OAI211_X1 U10027 ( .C1(n8518), .C2(n8517), .A(n8516), .B(n8515), .ZN(
        P2_U3181) );
  MUX2_X1 U10028 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8519), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10029 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8520), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10030 ( .A(n8636), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8528), .Z(
        P2_U3519) );
  MUX2_X1 U10031 ( .A(n8645), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8528), .Z(
        P2_U3518) );
  MUX2_X1 U10032 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8658), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10033 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8671), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10034 ( .A(n8682), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8528), .Z(
        P2_U3515) );
  MUX2_X1 U10035 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8672), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U10036 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8704), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10037 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8718), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10038 ( .A(n8705), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8528), .Z(
        P2_U3511) );
  MUX2_X1 U10039 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8719), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10040 ( .A(n8744), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8528), .Z(
        P2_U3509) );
  MUX2_X1 U10041 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8521), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10042 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8766), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10043 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8774), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10044 ( .A(n8787), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8528), .Z(
        P2_U3505) );
  MUX2_X1 U10045 ( .A(n8806), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8528), .Z(
        P2_U3504) );
  MUX2_X1 U10046 ( .A(n8786), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8528), .Z(
        P2_U3503) );
  MUX2_X1 U10047 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8805), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10048 ( .A(n8522), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8528), .Z(
        P2_U3501) );
  MUX2_X1 U10049 ( .A(n8523), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8528), .Z(
        P2_U3500) );
  MUX2_X1 U10050 ( .A(n8524), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8528), .Z(
        P2_U3499) );
  MUX2_X1 U10051 ( .A(n8525), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8528), .Z(
        P2_U3498) );
  MUX2_X1 U10052 ( .A(n8526), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8528), .Z(
        P2_U3497) );
  MUX2_X1 U10053 ( .A(n8527), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8528), .Z(
        P2_U3496) );
  MUX2_X1 U10054 ( .A(n4507), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8528), .Z(
        P2_U3494) );
  NOR2_X1 U10055 ( .A1(n8597), .A2(n8735), .ZN(n8529) );
  AOI21_X1 U10056 ( .B1(n8735), .B2(n8597), .A(n8529), .ZN(n8540) );
  NOR2_X1 U10057 ( .A1(n9942), .A2(n8532), .ZN(n8533) );
  NOR2_X1 U10058 ( .A1(n8797), .A2(n9951), .ZN(n9950) );
  NOR2_X1 U10059 ( .A1(n8533), .A2(n9950), .ZN(n9968) );
  MUX2_X1 U10060 ( .A(n8784), .B(P2_REG2_REG_14__SCAN_IN), .S(n9957), .Z(n8534) );
  INV_X1 U10061 ( .A(n8534), .ZN(n9967) );
  NAND2_X1 U10062 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8567), .ZN(n8536) );
  OAI21_X1 U10063 ( .B1(n8567), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8536), .ZN(
        n10000) );
  AOI21_X1 U10064 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8567), .A(n9999), .ZN(
        n8537) );
  NOR2_X1 U10065 ( .A1(n10009), .A2(n8537), .ZN(n8538) );
  XNOR2_X1 U10066 ( .A(n10009), .B(n8537), .ZN(n10021) );
  NOR2_X1 U10067 ( .A1(n10020), .A2(n10021), .ZN(n10019) );
  OR2_X1 U10068 ( .A1(n9876), .A2(n10020), .ZN(n8542) );
  NAND2_X1 U10069 ( .A1(n9876), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8541) );
  NAND2_X1 U10070 ( .A1(n8542), .A2(n8541), .ZN(n8543) );
  OR2_X1 U10071 ( .A1(n8543), .A2(n8577), .ZN(n8556) );
  XNOR2_X1 U10072 ( .A(n8543), .B(n10009), .ZN(n10014) );
  MUX2_X1 U10073 ( .A(n8759), .B(n8888), .S(n9876), .Z(n8544) );
  NAND2_X1 U10074 ( .A1(n9990), .A2(n8544), .ZN(n8555) );
  XNOR2_X1 U10075 ( .A(n8544), .B(n8567), .ZN(n9996) );
  MUX2_X1 U10076 ( .A(n9983), .B(n8890), .S(n9876), .Z(n8545) );
  NAND2_X1 U10077 ( .A1(n9974), .A2(n8545), .ZN(n8554) );
  XNOR2_X1 U10078 ( .A(n8545), .B(n8574), .ZN(n9979) );
  MUX2_X1 U10079 ( .A(n8784), .B(n8893), .S(n9876), .Z(n8546) );
  NAND2_X1 U10080 ( .A1(n9957), .A2(n8546), .ZN(n8553) );
  XNOR2_X1 U10081 ( .A(n8546), .B(n8568), .ZN(n9963) );
  MUX2_X1 U10082 ( .A(n8797), .B(n8896), .S(n9876), .Z(n8551) );
  NAND2_X1 U10083 ( .A1(n9942), .A2(n8551), .ZN(n8552) );
  INV_X1 U10084 ( .A(n8547), .ZN(n8549) );
  XNOR2_X1 U10085 ( .A(n8551), .B(n8571), .ZN(n9944) );
  NAND2_X1 U10086 ( .A1(n9945), .A2(n9944), .ZN(n9943) );
  NAND2_X1 U10087 ( .A1(n8552), .A2(n9943), .ZN(n9962) );
  NAND2_X1 U10088 ( .A1(n9979), .A2(n9978), .ZN(n9977) );
  NAND2_X1 U10089 ( .A1(n8554), .A2(n9977), .ZN(n9995) );
  NAND2_X1 U10090 ( .A1(n9996), .A2(n9995), .ZN(n9994) );
  OR2_X1 U10091 ( .A1(n9876), .A2(n8735), .ZN(n8558) );
  NAND2_X1 U10092 ( .A1(n9876), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8557) );
  NAND2_X1 U10093 ( .A1(n8558), .A2(n8557), .ZN(n8559) );
  NOR2_X1 U10094 ( .A1(n8560), .A2(n8559), .ZN(n8585) );
  NAND2_X1 U10095 ( .A1(n8560), .A2(n8559), .ZN(n8586) );
  INV_X1 U10096 ( .A(n8586), .ZN(n8561) );
  NOR2_X1 U10097 ( .A1(n8585), .A2(n8561), .ZN(n8562) );
  AOI21_X1 U10098 ( .B1(n8562), .B2(P2_U3893), .A(n10008), .ZN(n8566) );
  INV_X1 U10099 ( .A(n8562), .ZN(n8563) );
  NAND3_X1 U10100 ( .A1(n8563), .A2(n10016), .A3(n8597), .ZN(n8564) );
  OAI211_X1 U10101 ( .C1(n8566), .C2(n8597), .A(n8565), .B(n8564), .ZN(n8582)
         );
  XNOR2_X1 U10102 ( .A(n8587), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8598) );
  AOI22_X1 U10103 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8567), .B1(n9990), .B2(
        n8888), .ZN(n9993) );
  AOI22_X1 U10104 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8568), .B1(n9957), .B2(
        n8893), .ZN(n9960) );
  NAND2_X1 U10105 ( .A1(n8571), .A2(n8572), .ZN(n8573) );
  NAND2_X1 U10106 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n9947), .ZN(n9946) );
  NAND2_X1 U10107 ( .A1(n8574), .A2(n8575), .ZN(n8576) );
  NAND2_X1 U10108 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n9976), .ZN(n9975) );
  NAND2_X1 U10109 ( .A1(n8576), .A2(n9975), .ZN(n9992) );
  NAND2_X1 U10110 ( .A1(n8577), .A2(n8578), .ZN(n8579) );
  NAND2_X1 U10111 ( .A1(n8579), .A2(n10010), .ZN(n8599) );
  XOR2_X1 U10112 ( .A(n8598), .B(n8599), .Z(n8580) );
  NOR2_X1 U10113 ( .A1(n8580), .A2(n9928), .ZN(n8581) );
  AOI211_X1 U10114 ( .C1(n10007), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n8582), .B(
        n8581), .ZN(n8583) );
  XNOR2_X1 U10115 ( .A(n8596), .B(n8584), .ZN(n8588) );
  INV_X1 U10116 ( .A(n8588), .ZN(n8591) );
  XNOR2_X1 U10117 ( .A(n8596), .B(n8589), .ZN(n8600) );
  INV_X1 U10118 ( .A(n8600), .ZN(n8590) );
  MUX2_X1 U10119 ( .A(n8591), .B(n8590), .S(n9876), .Z(n8592) );
  XNOR2_X1 U10120 ( .A(n8593), .B(n8592), .ZN(n8602) );
  NAND2_X1 U10121 ( .A1(n10007), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8595) );
  NAND2_X1 U10122 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3151), .ZN(n8594) );
  OAI211_X1 U10123 ( .C1(n9885), .C2(n8596), .A(n8595), .B(n8594), .ZN(n8601)
         );
  NOR2_X1 U10124 ( .A1(n8819), .A2(n8606), .ZN(n8613) );
  AOI21_X1 U10125 ( .B1(n8810), .B2(n8905), .A(n8613), .ZN(n8609) );
  NAND2_X1 U10126 ( .A1(n8812), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8607) );
  OAI211_X1 U10127 ( .C1(n8907), .C2(n8733), .A(n8609), .B(n8607), .ZN(
        P2_U3202) );
  NAND2_X1 U10128 ( .A1(n8812), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8608) );
  OAI211_X1 U10129 ( .C1(n8910), .C2(n8733), .A(n8609), .B(n8608), .ZN(
        P2_U3203) );
  INV_X1 U10130 ( .A(n8610), .ZN(n8617) );
  NAND2_X1 U10131 ( .A1(n8611), .A2(n8835), .ZN(n8615) );
  NOR2_X1 U10132 ( .A1(n8847), .A2(n8733), .ZN(n8612) );
  AOI211_X1 U10133 ( .C1(n8812), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8613), .B(
        n8612), .ZN(n8614) );
  OAI211_X1 U10134 ( .C1(n8617), .C2(n8616), .A(n8615), .B(n8614), .ZN(
        P2_U3204) );
  XNOR2_X1 U10135 ( .A(n8618), .B(n8620), .ZN(n8916) );
  NOR2_X1 U10136 ( .A1(n8623), .A2(n8757), .ZN(n8624) );
  INV_X1 U10137 ( .A(n8848), .ZN(n8911) );
  MUX2_X1 U10138 ( .A(n8628), .B(n8911), .S(n8835), .Z(n8632) );
  INV_X1 U10139 ( .A(n8629), .ZN(n8630) );
  AOI22_X1 U10140 ( .A1(n8913), .A2(n8813), .B1(n8769), .B2(n8630), .ZN(n8631)
         );
  OAI211_X1 U10141 ( .C1(n8916), .C2(n8816), .A(n8632), .B(n8631), .ZN(
        P2_U3205) );
  XNOR2_X1 U10142 ( .A(n8633), .B(n8634), .ZN(n8922) );
  INV_X1 U10143 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8638) );
  XNOR2_X1 U10144 ( .A(n8635), .B(n8634), .ZN(n8637) );
  AOI222_X1 U10145 ( .A1(n8808), .A2(n8637), .B1(n8658), .B2(n8827), .C1(n8636), .C2(n8824), .ZN(n8917) );
  MUX2_X1 U10146 ( .A(n8638), .B(n8917), .S(n8835), .Z(n8641) );
  AOI22_X1 U10147 ( .A1(n8919), .A2(n8813), .B1(n8769), .B2(n8639), .ZN(n8640)
         );
  OAI211_X1 U10148 ( .C1(n8922), .C2(n8816), .A(n8641), .B(n8640), .ZN(
        P2_U3206) );
  XNOR2_X1 U10149 ( .A(n8642), .B(n8643), .ZN(n8928) );
  INV_X1 U10150 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8650) );
  XNOR2_X1 U10151 ( .A(n8644), .B(n8643), .ZN(n8649) );
  NAND2_X1 U10152 ( .A1(n8645), .A2(n8824), .ZN(n8646) );
  OAI21_X1 U10153 ( .B1(n8647), .B2(n8755), .A(n8646), .ZN(n8648) );
  AOI21_X1 U10154 ( .B1(n8649), .B2(n8808), .A(n8648), .ZN(n8923) );
  MUX2_X1 U10155 ( .A(n8650), .B(n8923), .S(n8835), .Z(n8653) );
  AOI22_X1 U10156 ( .A1(n8925), .A2(n8813), .B1(n8769), .B2(n8651), .ZN(n8652)
         );
  OAI211_X1 U10157 ( .C1(n8928), .C2(n8816), .A(n8653), .B(n8652), .ZN(
        P2_U3207) );
  XNOR2_X1 U10158 ( .A(n8655), .B(n8654), .ZN(n8934) );
  INV_X1 U10159 ( .A(n8931), .ZN(n8660) );
  XNOR2_X1 U10160 ( .A(n8657), .B(n8656), .ZN(n8659) );
  AOI222_X1 U10161 ( .A1(n8808), .A2(n8659), .B1(n8658), .B2(n8824), .C1(n8682), .C2(n8827), .ZN(n8929) );
  OAI21_X1 U10162 ( .B1(n8660), .B2(n8820), .A(n8929), .ZN(n8661) );
  NAND2_X1 U10163 ( .A1(n8661), .A2(n8835), .ZN(n8664) );
  AOI22_X1 U10164 ( .A1(n8662), .A2(n8769), .B1(n8812), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8663) );
  OAI211_X1 U10165 ( .C1(n8934), .C2(n8816), .A(n8664), .B(n8663), .ZN(
        P2_U3208) );
  INV_X1 U10166 ( .A(n8665), .ZN(n8667) );
  OAI21_X1 U10167 ( .B1(n8679), .B2(n8667), .A(n8666), .ZN(n8668) );
  XNOR2_X1 U10168 ( .A(n8668), .B(n8670), .ZN(n8940) );
  INV_X1 U10169 ( .A(n8937), .ZN(n8674) );
  XOR2_X1 U10170 ( .A(n8670), .B(n8669), .Z(n8673) );
  AOI222_X1 U10171 ( .A1(n8808), .A2(n8673), .B1(n8672), .B2(n8827), .C1(n8671), .C2(n8824), .ZN(n8935) );
  OAI21_X1 U10172 ( .B1(n8674), .B2(n8820), .A(n8935), .ZN(n8675) );
  NAND2_X1 U10173 ( .A1(n8675), .A2(n8810), .ZN(n8678) );
  AOI22_X1 U10174 ( .A1(n8812), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8769), .B2(
        n8676), .ZN(n8677) );
  OAI211_X1 U10175 ( .C1(n8940), .C2(n8816), .A(n8678), .B(n8677), .ZN(
        P2_U3209) );
  XOR2_X1 U10176 ( .A(n8680), .B(n8679), .Z(n8946) );
  INV_X1 U10177 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8684) );
  XNOR2_X1 U10178 ( .A(n8681), .B(n8680), .ZN(n8683) );
  AOI222_X1 U10179 ( .A1(n8808), .A2(n8683), .B1(n8704), .B2(n8827), .C1(n8682), .C2(n8824), .ZN(n8941) );
  MUX2_X1 U10180 ( .A(n8684), .B(n8941), .S(n8835), .Z(n8687) );
  AOI22_X1 U10181 ( .A1(n8943), .A2(n8813), .B1(n8769), .B2(n8685), .ZN(n8686)
         );
  OAI211_X1 U10182 ( .C1(n8946), .C2(n8816), .A(n8687), .B(n8686), .ZN(
        P2_U3210) );
  XNOR2_X1 U10183 ( .A(n8688), .B(n8689), .ZN(n8690) );
  OAI222_X1 U10184 ( .A1(n8757), .A2(n8692), .B1(n8755), .B2(n8691), .C1(n8831), .C2(n8690), .ZN(n8866) );
  INV_X1 U10185 ( .A(n8866), .ZN(n8700) );
  XNOR2_X1 U10186 ( .A(n8694), .B(n8693), .ZN(n8867) );
  INV_X1 U10187 ( .A(n8695), .ZN(n8950) );
  AOI22_X1 U10188 ( .A1(n8812), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8769), .B2(
        n8696), .ZN(n8697) );
  OAI21_X1 U10189 ( .B1(n8950), .B2(n8733), .A(n8697), .ZN(n8698) );
  AOI21_X1 U10190 ( .B1(n8867), .B2(n8738), .A(n8698), .ZN(n8699) );
  OAI21_X1 U10191 ( .B1(n8700), .B2(n8812), .A(n8699), .ZN(P2_U3211) );
  XNOR2_X1 U10192 ( .A(n8701), .B(n8703), .ZN(n8956) );
  INV_X1 U10193 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8707) );
  XNOR2_X1 U10194 ( .A(n8702), .B(n8703), .ZN(n8706) );
  AOI222_X1 U10195 ( .A1(n8808), .A2(n8706), .B1(n8705), .B2(n8827), .C1(n8704), .C2(n8824), .ZN(n8951) );
  MUX2_X1 U10196 ( .A(n8707), .B(n8951), .S(n8835), .Z(n8710) );
  AOI22_X1 U10197 ( .A1(n8953), .A2(n8813), .B1(n8769), .B2(n8708), .ZN(n8709)
         );
  OAI211_X1 U10198 ( .C1(n8956), .C2(n8816), .A(n8710), .B(n8709), .ZN(
        P2_U3212) );
  NAND2_X1 U10199 ( .A1(n8712), .A2(n8711), .ZN(n8714) );
  INV_X1 U10200 ( .A(n8716), .ZN(n8713) );
  XNOR2_X1 U10201 ( .A(n8714), .B(n8713), .ZN(n8960) );
  OAI21_X1 U10202 ( .B1(n8717), .B2(n8716), .A(n8715), .ZN(n8720) );
  AOI222_X1 U10203 ( .A1(n8808), .A2(n8720), .B1(n8719), .B2(n8827), .C1(n8718), .C2(n8824), .ZN(n8721) );
  INV_X1 U10204 ( .A(n8721), .ZN(n8873) );
  NAND2_X1 U10205 ( .A1(n8873), .A2(n8810), .ZN(n8727) );
  INV_X1 U10206 ( .A(n8722), .ZN(n8723) );
  OAI22_X1 U10207 ( .A1(n8810), .A2(n8724), .B1(n8723), .B2(n8819), .ZN(n8725)
         );
  AOI21_X1 U10208 ( .B1(n8874), .B2(n8813), .A(n8725), .ZN(n8726) );
  OAI211_X1 U10209 ( .C1(n8960), .C2(n8816), .A(n8727), .B(n8726), .ZN(
        P2_U3213) );
  XNOR2_X1 U10210 ( .A(n8728), .B(n4515), .ZN(n8731) );
  OAI22_X1 U10211 ( .A1(n8729), .A2(n8757), .B1(n8756), .B2(n8755), .ZN(n8730)
         );
  AOI21_X1 U10212 ( .B1(n8731), .B2(n8808), .A(n8730), .ZN(n8878) );
  XNOR2_X1 U10213 ( .A(n8732), .B(n4515), .ZN(n8877) );
  NOR2_X1 U10214 ( .A1(n8965), .A2(n8733), .ZN(n8737) );
  OAI22_X1 U10215 ( .A1(n8810), .A2(n8735), .B1(n8734), .B2(n8819), .ZN(n8736)
         );
  AOI211_X1 U10216 ( .C1(n8877), .C2(n8738), .A(n8737), .B(n8736), .ZN(n8739)
         );
  OAI21_X1 U10217 ( .B1(n8812), .B2(n8878), .A(n8739), .ZN(P2_U3215) );
  XNOR2_X1 U10218 ( .A(n8740), .B(n8741), .ZN(n8971) );
  XNOR2_X1 U10219 ( .A(n8743), .B(n8742), .ZN(n8745) );
  AOI222_X1 U10220 ( .A1(n8808), .A2(n8745), .B1(n8744), .B2(n8824), .C1(n8766), .C2(n8827), .ZN(n8966) );
  MUX2_X1 U10221 ( .A(n10020), .B(n8966), .S(n8835), .Z(n8748) );
  AOI22_X1 U10222 ( .A1(n8968), .A2(n8813), .B1(n8769), .B2(n8746), .ZN(n8747)
         );
  OAI211_X1 U10223 ( .C1(n8971), .C2(n8816), .A(n8748), .B(n8747), .ZN(
        P2_U3216) );
  INV_X1 U10224 ( .A(n8752), .ZN(n8749) );
  XNOR2_X1 U10225 ( .A(n8750), .B(n8749), .ZN(n8975) );
  XNOR2_X1 U10226 ( .A(n8751), .B(n8752), .ZN(n8753) );
  OAI222_X1 U10227 ( .A1(n8757), .A2(n8756), .B1(n8755), .B2(n8754), .C1(n8753), .C2(n8831), .ZN(n8886) );
  NAND2_X1 U10228 ( .A1(n8886), .A2(n8810), .ZN(n8762) );
  OAI22_X1 U10229 ( .A1(n8810), .A2(n8759), .B1(n8758), .B2(n8819), .ZN(n8760)
         );
  AOI21_X1 U10230 ( .B1(n8887), .B2(n8813), .A(n8760), .ZN(n8761) );
  OAI211_X1 U10231 ( .C1(n8975), .C2(n8816), .A(n8762), .B(n8761), .ZN(
        P2_U3217) );
  XNOR2_X1 U10232 ( .A(n8763), .B(n8764), .ZN(n8981) );
  XNOR2_X1 U10233 ( .A(n8765), .B(n8764), .ZN(n8767) );
  AOI222_X1 U10234 ( .A1(n8808), .A2(n8767), .B1(n8766), .B2(n8824), .C1(n8787), .C2(n8827), .ZN(n8976) );
  MUX2_X1 U10235 ( .A(n9983), .B(n8976), .S(n8810), .Z(n8772) );
  INV_X1 U10236 ( .A(n8768), .ZN(n8770) );
  AOI22_X1 U10237 ( .A1(n8978), .A2(n8813), .B1(n8770), .B2(n8769), .ZN(n8771)
         );
  OAI211_X1 U10238 ( .C1(n8981), .C2(n8816), .A(n8772), .B(n8771), .ZN(
        P2_U3218) );
  XNOR2_X1 U10239 ( .A(n8773), .B(n8781), .ZN(n8775) );
  AOI222_X1 U10240 ( .A1(n8808), .A2(n8775), .B1(n8774), .B2(n8824), .C1(n8806), .C2(n8827), .ZN(n8982) );
  INV_X1 U10241 ( .A(n8982), .ZN(n8779) );
  INV_X1 U10242 ( .A(n8984), .ZN(n8777) );
  OAI22_X1 U10243 ( .A1(n8777), .A2(n8820), .B1(n8776), .B2(n8819), .ZN(n8778)
         );
  OAI21_X1 U10244 ( .B1(n8779), .B2(n8778), .A(n8835), .ZN(n8783) );
  XNOR2_X1 U10245 ( .A(n8780), .B(n8781), .ZN(n8987) );
  OR2_X1 U10246 ( .A1(n8987), .A2(n8816), .ZN(n8782) );
  OAI211_X1 U10247 ( .C1(n8810), .C2(n8784), .A(n8783), .B(n8782), .ZN(
        P2_U3219) );
  XNOR2_X1 U10248 ( .A(n8785), .B(n8793), .ZN(n8788) );
  AOI222_X1 U10249 ( .A1(n8808), .A2(n8788), .B1(n8787), .B2(n8824), .C1(n8786), .C2(n8827), .ZN(n8988) );
  INV_X1 U10250 ( .A(n8988), .ZN(n8792) );
  INV_X1 U10251 ( .A(n8990), .ZN(n8790) );
  OAI22_X1 U10252 ( .A1(n8790), .A2(n8820), .B1(n8789), .B2(n8819), .ZN(n8791)
         );
  OAI21_X1 U10253 ( .B1(n8792), .B2(n8791), .A(n8835), .ZN(n8796) );
  XNOR2_X1 U10254 ( .A(n8794), .B(n8793), .ZN(n8993) );
  OR2_X1 U10255 ( .A1(n8993), .A2(n8816), .ZN(n8795) );
  OAI211_X1 U10256 ( .C1(n8810), .C2(n8797), .A(n8796), .B(n8795), .ZN(
        P2_U3220) );
  INV_X1 U10257 ( .A(n7837), .ZN(n8800) );
  OAI21_X1 U10258 ( .B1(n8800), .B2(n8799), .A(n8798), .ZN(n8802) );
  NAND2_X1 U10259 ( .A1(n8802), .A2(n8801), .ZN(n9000) );
  XNOR2_X1 U10260 ( .A(n8804), .B(n8803), .ZN(n8807) );
  AOI222_X1 U10261 ( .A1(n8808), .A2(n8807), .B1(n8806), .B2(n8824), .C1(n8805), .C2(n8827), .ZN(n8994) );
  OAI21_X1 U10262 ( .B1(n8809), .B2(n8819), .A(n8994), .ZN(n8811) );
  NAND2_X1 U10263 ( .A1(n8811), .A2(n8810), .ZN(n8815) );
  AOI22_X1 U10264 ( .A1(n8996), .A2(n8813), .B1(P2_REG2_REG_12__SCAN_IN), .B2(
        n8812), .ZN(n8814) );
  OAI211_X1 U10265 ( .C1(n9000), .C2(n8816), .A(n8815), .B(n8814), .ZN(
        P2_U3221) );
  OAI21_X1 U10266 ( .B1(n8818), .B2(n8822), .A(n8817), .ZN(n10031) );
  OAI22_X1 U10267 ( .A1(n10028), .A2(n8820), .B1(n7150), .B2(n8819), .ZN(n8832) );
  XNOR2_X1 U10268 ( .A(n8821), .B(n8822), .ZN(n8830) );
  NAND2_X1 U10269 ( .A1(n10031), .A2(n8823), .ZN(n8829) );
  AOI22_X1 U10270 ( .A1(n8827), .A2(n8826), .B1(n4507), .B2(n8824), .ZN(n8828)
         );
  OAI211_X1 U10271 ( .C1(n8831), .C2(n8830), .A(n8829), .B(n8828), .ZN(n10029)
         );
  AOI211_X1 U10272 ( .C1(n8833), .C2(n10031), .A(n8832), .B(n10029), .ZN(n8834) );
  INV_X1 U10273 ( .A(n8834), .ZN(n8836) );
  MUX2_X1 U10274 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n8836), .S(n8835), .Z(
        P2_U3231) );
  NAND2_X1 U10275 ( .A1(n8837), .A2(n8900), .ZN(n8838) );
  NAND2_X1 U10276 ( .A1(n10101), .A2(n8905), .ZN(n8840) );
  OAI211_X1 U10277 ( .C1(n10101), .C2(n7095), .A(n8838), .B(n8840), .ZN(
        P2_U3490) );
  INV_X1 U10278 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8842) );
  INV_X1 U10279 ( .A(n8910), .ZN(n8839) );
  NAND2_X1 U10280 ( .A1(n8839), .A2(n8900), .ZN(n8841) );
  OAI211_X1 U10281 ( .C1(n10101), .C2(n8842), .A(n8841), .B(n8840), .ZN(
        P2_U3489) );
  OAI21_X1 U10282 ( .B1(n8847), .B2(n8882), .A(n8846), .ZN(P2_U3488) );
  MUX2_X1 U10283 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8848), .S(n10101), .Z(
        n8850) );
  OAI22_X1 U10284 ( .A1(n8916), .A2(n8903), .B1(n6210), .B2(n8882), .ZN(n8849)
         );
  OR2_X1 U10285 ( .A1(n8850), .A2(n8849), .ZN(P2_U3487) );
  MUX2_X1 U10286 ( .A(n8851), .B(n8917), .S(n10101), .Z(n8853) );
  NAND2_X1 U10287 ( .A1(n8919), .A2(n8900), .ZN(n8852) );
  OAI211_X1 U10288 ( .C1(n8922), .C2(n8903), .A(n8853), .B(n8852), .ZN(
        P2_U3486) );
  MUX2_X1 U10289 ( .A(n8854), .B(n8923), .S(n10101), .Z(n8856) );
  NAND2_X1 U10290 ( .A1(n8925), .A2(n8900), .ZN(n8855) );
  OAI211_X1 U10291 ( .C1(n8928), .C2(n8903), .A(n8856), .B(n8855), .ZN(
        P2_U3485) );
  MUX2_X1 U10292 ( .A(n8857), .B(n8929), .S(n10101), .Z(n8859) );
  NAND2_X1 U10293 ( .A1(n8931), .A2(n8900), .ZN(n8858) );
  OAI211_X1 U10294 ( .C1(n8934), .C2(n8903), .A(n8859), .B(n8858), .ZN(
        P2_U3484) );
  MUX2_X1 U10295 ( .A(n8860), .B(n8935), .S(n10101), .Z(n8862) );
  NAND2_X1 U10296 ( .A1(n8937), .A2(n8900), .ZN(n8861) );
  OAI211_X1 U10297 ( .C1(n8903), .C2(n8940), .A(n8862), .B(n8861), .ZN(
        P2_U3483) );
  MUX2_X1 U10298 ( .A(n8863), .B(n8941), .S(n10101), .Z(n8865) );
  NAND2_X1 U10299 ( .A1(n8943), .A2(n8900), .ZN(n8864) );
  OAI211_X1 U10300 ( .C1(n8946), .C2(n8903), .A(n8865), .B(n8864), .ZN(
        P2_U3482) );
  INV_X1 U10301 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8868) );
  AOI21_X1 U10302 ( .B1(n10083), .B2(n8867), .A(n8866), .ZN(n8947) );
  MUX2_X1 U10303 ( .A(n8868), .B(n8947), .S(n10101), .Z(n8869) );
  OAI21_X1 U10304 ( .B1(n8950), .B2(n8882), .A(n8869), .ZN(P2_U3481) );
  INV_X1 U10305 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8870) );
  MUX2_X1 U10306 ( .A(n8870), .B(n8951), .S(n10101), .Z(n8872) );
  NAND2_X1 U10307 ( .A1(n8953), .A2(n8900), .ZN(n8871) );
  OAI211_X1 U10308 ( .C1(n8903), .C2(n8956), .A(n8872), .B(n8871), .ZN(
        P2_U3480) );
  AOI21_X1 U10309 ( .B1(n10063), .B2(n8874), .A(n8873), .ZN(n8957) );
  MUX2_X1 U10310 ( .A(n8875), .B(n8957), .S(n10101), .Z(n8876) );
  OAI21_X1 U10311 ( .B1(n8960), .B2(n8903), .A(n8876), .ZN(P2_U3479) );
  INV_X1 U10312 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8880) );
  NAND2_X1 U10313 ( .A1(n8877), .A2(n10083), .ZN(n8879) );
  AND2_X1 U10314 ( .A1(n8879), .A2(n8878), .ZN(n8961) );
  MUX2_X1 U10315 ( .A(n8880), .B(n8961), .S(n10101), .Z(n8881) );
  OAI21_X1 U10316 ( .B1(n8965), .B2(n8882), .A(n8881), .ZN(P2_U3477) );
  MUX2_X1 U10317 ( .A(n8883), .B(n8966), .S(n10101), .Z(n8885) );
  NAND2_X1 U10318 ( .A1(n8968), .A2(n8900), .ZN(n8884) );
  OAI211_X1 U10319 ( .C1(n8903), .C2(n8971), .A(n8885), .B(n8884), .ZN(
        P2_U3476) );
  AOI21_X1 U10320 ( .B1(n10063), .B2(n8887), .A(n8886), .ZN(n8972) );
  MUX2_X1 U10321 ( .A(n8888), .B(n8972), .S(n10101), .Z(n8889) );
  OAI21_X1 U10322 ( .B1(n8975), .B2(n8903), .A(n8889), .ZN(P2_U3475) );
  MUX2_X1 U10323 ( .A(n8890), .B(n8976), .S(n10101), .Z(n8892) );
  NAND2_X1 U10324 ( .A1(n8978), .A2(n8900), .ZN(n8891) );
  OAI211_X1 U10325 ( .C1(n8903), .C2(n8981), .A(n8892), .B(n8891), .ZN(
        P2_U3474) );
  MUX2_X1 U10326 ( .A(n8893), .B(n8982), .S(n10101), .Z(n8895) );
  NAND2_X1 U10327 ( .A1(n8984), .A2(n8900), .ZN(n8894) );
  OAI211_X1 U10328 ( .C1(n8903), .C2(n8987), .A(n8895), .B(n8894), .ZN(
        P2_U3473) );
  MUX2_X1 U10329 ( .A(n8896), .B(n8988), .S(n10101), .Z(n8898) );
  NAND2_X1 U10330 ( .A1(n8990), .A2(n8900), .ZN(n8897) );
  OAI211_X1 U10331 ( .C1(n8993), .C2(n8903), .A(n8898), .B(n8897), .ZN(
        P2_U3472) );
  MUX2_X1 U10332 ( .A(n8899), .B(n8994), .S(n10101), .Z(n8902) );
  NAND2_X1 U10333 ( .A1(n8996), .A2(n8900), .ZN(n8901) );
  OAI211_X1 U10334 ( .C1(n8903), .C2(n9000), .A(n8902), .B(n8901), .ZN(
        P2_U3471) );
  MUX2_X1 U10335 ( .A(n8904), .B(P2_REG1_REG_0__SCAN_IN), .S(n10098), .Z(
        P2_U3459) );
  NAND2_X1 U10336 ( .A1(n10084), .A2(n8905), .ZN(n8908) );
  NAND2_X1 U10337 ( .A1(n10086), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8906) );
  OAI211_X1 U10338 ( .C1(n8907), .C2(n8964), .A(n8908), .B(n8906), .ZN(
        P2_U3458) );
  NAND2_X1 U10339 ( .A1(n10086), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8909) );
  OAI211_X1 U10340 ( .C1(n8910), .C2(n8964), .A(n8909), .B(n8908), .ZN(
        P2_U3457) );
  MUX2_X1 U10341 ( .A(n8912), .B(n8911), .S(n10084), .Z(n8915) );
  NAND2_X1 U10342 ( .A1(n8913), .A2(n6301), .ZN(n8914) );
  OAI211_X1 U10343 ( .C1(n8916), .C2(n8999), .A(n8915), .B(n8914), .ZN(
        P2_U3455) );
  INV_X1 U10344 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8918) );
  MUX2_X1 U10345 ( .A(n8918), .B(n8917), .S(n10084), .Z(n8921) );
  NAND2_X1 U10346 ( .A1(n8919), .A2(n6301), .ZN(n8920) );
  OAI211_X1 U10347 ( .C1(n8922), .C2(n8999), .A(n8921), .B(n8920), .ZN(
        P2_U3454) );
  INV_X1 U10348 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8924) );
  MUX2_X1 U10349 ( .A(n8924), .B(n8923), .S(n10084), .Z(n8927) );
  NAND2_X1 U10350 ( .A1(n8925), .A2(n6301), .ZN(n8926) );
  OAI211_X1 U10351 ( .C1(n8928), .C2(n8999), .A(n8927), .B(n8926), .ZN(
        P2_U3453) );
  INV_X1 U10352 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8930) );
  MUX2_X1 U10353 ( .A(n8930), .B(n8929), .S(n10084), .Z(n8933) );
  NAND2_X1 U10354 ( .A1(n8931), .A2(n6301), .ZN(n8932) );
  OAI211_X1 U10355 ( .C1(n8934), .C2(n8999), .A(n8933), .B(n8932), .ZN(
        P2_U3452) );
  INV_X1 U10356 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8936) );
  MUX2_X1 U10357 ( .A(n8936), .B(n8935), .S(n10084), .Z(n8939) );
  NAND2_X1 U10358 ( .A1(n8937), .A2(n6301), .ZN(n8938) );
  OAI211_X1 U10359 ( .C1(n8940), .C2(n8999), .A(n8939), .B(n8938), .ZN(
        P2_U3451) );
  INV_X1 U10360 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8942) );
  MUX2_X1 U10361 ( .A(n8942), .B(n8941), .S(n10084), .Z(n8945) );
  NAND2_X1 U10362 ( .A1(n8943), .A2(n6301), .ZN(n8944) );
  OAI211_X1 U10363 ( .C1(n8946), .C2(n8999), .A(n8945), .B(n8944), .ZN(
        P2_U3450) );
  INV_X1 U10364 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8948) );
  MUX2_X1 U10365 ( .A(n8948), .B(n8947), .S(n10084), .Z(n8949) );
  OAI21_X1 U10366 ( .B1(n8950), .B2(n8964), .A(n8949), .ZN(P2_U3449) );
  INV_X1 U10367 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8952) );
  MUX2_X1 U10368 ( .A(n8952), .B(n8951), .S(n10084), .Z(n8955) );
  NAND2_X1 U10369 ( .A1(n8953), .A2(n6301), .ZN(n8954) );
  OAI211_X1 U10370 ( .C1(n8956), .C2(n8999), .A(n8955), .B(n8954), .ZN(
        P2_U3448) );
  MUX2_X1 U10371 ( .A(n8958), .B(n8957), .S(n10084), .Z(n8959) );
  OAI21_X1 U10372 ( .B1(n8960), .B2(n8999), .A(n8959), .ZN(P2_U3447) );
  MUX2_X1 U10373 ( .A(n8962), .B(n8961), .S(n10084), .Z(n8963) );
  OAI21_X1 U10374 ( .B1(n8965), .B2(n8964), .A(n8963), .ZN(P2_U3444) );
  INV_X1 U10375 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8967) );
  MUX2_X1 U10376 ( .A(n8967), .B(n8966), .S(n10084), .Z(n8970) );
  NAND2_X1 U10377 ( .A1(n8968), .A2(n6301), .ZN(n8969) );
  OAI211_X1 U10378 ( .C1(n8971), .C2(n8999), .A(n8970), .B(n8969), .ZN(
        P2_U3441) );
  INV_X1 U10379 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8973) );
  MUX2_X1 U10380 ( .A(n8973), .B(n8972), .S(n10084), .Z(n8974) );
  OAI21_X1 U10381 ( .B1(n8975), .B2(n8999), .A(n8974), .ZN(P2_U3438) );
  INV_X1 U10382 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8977) );
  MUX2_X1 U10383 ( .A(n8977), .B(n8976), .S(n10084), .Z(n8980) );
  NAND2_X1 U10384 ( .A1(n8978), .A2(n6301), .ZN(n8979) );
  OAI211_X1 U10385 ( .C1(n8981), .C2(n8999), .A(n8980), .B(n8979), .ZN(
        P2_U3435) );
  INV_X1 U10386 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8983) );
  MUX2_X1 U10387 ( .A(n8983), .B(n8982), .S(n10084), .Z(n8986) );
  NAND2_X1 U10388 ( .A1(n8984), .A2(n6301), .ZN(n8985) );
  OAI211_X1 U10389 ( .C1(n8987), .C2(n8999), .A(n8986), .B(n8985), .ZN(
        P2_U3432) );
  INV_X1 U10390 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8989) );
  MUX2_X1 U10391 ( .A(n8989), .B(n8988), .S(n10084), .Z(n8992) );
  NAND2_X1 U10392 ( .A1(n8990), .A2(n6301), .ZN(n8991) );
  OAI211_X1 U10393 ( .C1(n8993), .C2(n8999), .A(n8992), .B(n8991), .ZN(
        P2_U3429) );
  INV_X1 U10394 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n8995) );
  MUX2_X1 U10395 ( .A(n8995), .B(n8994), .S(n10084), .Z(n8998) );
  NAND2_X1 U10396 ( .A1(n8996), .A2(n6301), .ZN(n8997) );
  OAI211_X1 U10397 ( .C1(n9000), .C2(n8999), .A(n8998), .B(n8997), .ZN(
        P2_U3426) );
  INV_X1 U10398 ( .A(n9001), .ZN(n9681) );
  NOR4_X1 U10399 ( .A1(n9003), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n9002), .ZN(n9004) );
  AOI21_X1 U10400 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n9005), .A(n9004), .ZN(
        n9006) );
  OAI21_X1 U10401 ( .B1(n9681), .B2(n9018), .A(n9006), .ZN(P2_U3264) );
  OAI222_X1 U10402 ( .A1(n9015), .A2(n9009), .B1(n9018), .B2(n9008), .C1(
        P2_U3151), .C2(n9007), .ZN(P2_U3265) );
  NAND2_X1 U10403 ( .A1(n6198), .A2(n9010), .ZN(n9012) );
  OAI211_X1 U10404 ( .C1(n9015), .C2(n9013), .A(n9012), .B(n9011), .ZN(
        P2_U3267) );
  INV_X1 U10405 ( .A(n9014), .ZN(n9688) );
  OAI222_X1 U10406 ( .A1(n9018), .A2(n9688), .B1(P2_U3151), .B2(n9017), .C1(
        n9016), .C2(n9015), .ZN(P2_U3269) );
  NAND2_X1 U10407 ( .A1(n9021), .A2(n9020), .ZN(n9022) );
  XOR2_X1 U10408 ( .A(n9023), .B(n9022), .Z(n9030) );
  OAI22_X1 U10409 ( .A1(n9025), .A2(n9694), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9024), .ZN(n9027) );
  NOR2_X1 U10410 ( .A1(n9849), .A2(n9722), .ZN(n9026) );
  AOI211_X1 U10411 ( .C1(n9187), .C2(n9028), .A(n9027), .B(n9026), .ZN(n9029)
         );
  OAI21_X1 U10412 ( .B1(n9030), .B2(n9699), .A(n9029), .ZN(P1_U3215) );
  OR2_X1 U10413 ( .A1(n9071), .A2(n9168), .ZN(n9032) );
  NAND2_X1 U10414 ( .A1(n9197), .A2(n9181), .ZN(n9031) );
  AND2_X1 U10415 ( .A1(n9032), .A2(n9031), .ZN(n9444) );
  INV_X1 U10416 ( .A(n9033), .ZN(n9447) );
  AOI22_X1 U10417 ( .A1(n9447), .A2(n9187), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9034) );
  OAI21_X1 U10418 ( .B1(n9444), .B2(n9694), .A(n9034), .ZN(n9038) );
  OAI21_X1 U10419 ( .B1(n9139), .B2(n9143), .A(n9035), .ZN(n9036) );
  AOI21_X1 U10420 ( .B1(n9036), .B2(n9104), .A(n9699), .ZN(n9037) );
  AOI211_X1 U10421 ( .C1(n9608), .C2(n9703), .A(n9038), .B(n9037), .ZN(n9039)
         );
  INV_X1 U10422 ( .A(n9039), .ZN(P1_U3216) );
  OAI21_X1 U10423 ( .B1(n9042), .B2(n9041), .A(n9040), .ZN(n9043) );
  NAND2_X1 U10424 ( .A1(n9043), .A2(n9724), .ZN(n9047) );
  INV_X1 U10425 ( .A(n9044), .ZN(n9507) );
  AOI22_X1 U10426 ( .A1(n9199), .A2(n9180), .B1(n9181), .B2(n9201), .ZN(n9503)
         );
  NAND2_X1 U10427 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9347) );
  OAI21_X1 U10428 ( .B1(n9503), .B2(n9694), .A(n9347), .ZN(n9045) );
  AOI21_X1 U10429 ( .B1(n9507), .B2(n9187), .A(n9045), .ZN(n9046) );
  OAI211_X1 U10430 ( .C1(n9510), .C2(n9722), .A(n9047), .B(n9046), .ZN(
        P1_U3219) );
  XNOR2_X1 U10431 ( .A(n9049), .B(n9048), .ZN(n9050) );
  XNOR2_X1 U10432 ( .A(n9051), .B(n9050), .ZN(n9057) );
  AND2_X1 U10433 ( .A1(n9199), .A2(n9181), .ZN(n9052) );
  AOI21_X1 U10434 ( .B1(n9197), .B2(n9180), .A(n9052), .ZN(n9475) );
  NOR2_X1 U10435 ( .A1(n9475), .A2(n9694), .ZN(n9055) );
  OAI22_X1 U10436 ( .A1(n9727), .A2(n9479), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9053), .ZN(n9054) );
  AOI211_X1 U10437 ( .C1(n9478), .C2(n9703), .A(n9055), .B(n9054), .ZN(n9056)
         );
  OAI21_X1 U10438 ( .B1(n9057), .B2(n9699), .A(n9056), .ZN(P1_U3223) );
  NOR3_X1 U10439 ( .A1(n9060), .A2(n5053), .A3(n9059), .ZN(n9062) );
  INV_X1 U10440 ( .A(n9132), .ZN(n9061) );
  OAI21_X1 U10441 ( .B1(n9062), .B2(n9061), .A(n9724), .ZN(n9068) );
  NOR2_X1 U10442 ( .A1(n9063), .A2(n9694), .ZN(n9064) );
  AOI211_X1 U10443 ( .C1(n9187), .C2(n9066), .A(n9065), .B(n9064), .ZN(n9067)
         );
  OAI211_X1 U10444 ( .C1(n4852), .C2(n9722), .A(n9068), .B(n9067), .ZN(
        P1_U3224) );
  AOI21_X1 U10445 ( .B1(n9070), .B2(n9069), .A(n4530), .ZN(n9078) );
  OR2_X1 U10446 ( .A1(n9071), .A2(n9091), .ZN(n9074) );
  OR2_X1 U10447 ( .A1(n9072), .A2(n9168), .ZN(n9073) );
  AND2_X1 U10448 ( .A1(n9074), .A2(n9073), .ZN(n9411) );
  AOI22_X1 U10449 ( .A1(n9187), .A2(n9419), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9075) );
  OAI21_X1 U10450 ( .B1(n9411), .B2(n9694), .A(n9075), .ZN(n9076) );
  AOI21_X1 U10451 ( .B1(n9418), .B2(n9703), .A(n9076), .ZN(n9077) );
  OAI21_X1 U10452 ( .B1(n9078), .B2(n9699), .A(n9077), .ZN(P1_U3225) );
  AOI21_X1 U10453 ( .B1(n9080), .B2(n9079), .A(n8045), .ZN(n9085) );
  AOI22_X1 U10454 ( .A1(n9181), .A2(n9204), .B1(n9202), .B2(n9180), .ZN(n9546)
         );
  NAND2_X1 U10455 ( .A1(n9187), .A2(n9551), .ZN(n9081) );
  OAI211_X1 U10456 ( .C1(n9546), .C2(n9694), .A(n9082), .B(n9081), .ZN(n9083)
         );
  AOI21_X1 U10457 ( .B1(n9548), .B2(n9703), .A(n9083), .ZN(n9084) );
  OAI21_X1 U10458 ( .B1(n9085), .B2(n9699), .A(n9084), .ZN(P1_U3226) );
  OAI21_X1 U10459 ( .B1(n9088), .B2(n9087), .A(n9086), .ZN(n9089) );
  NAND2_X1 U10460 ( .A1(n9089), .A2(n9724), .ZN(n9101) );
  NAND2_X1 U10461 ( .A1(n9201), .A2(n9180), .ZN(n9090) );
  OAI21_X1 U10462 ( .B1(n9092), .B2(n9091), .A(n9090), .ZN(n9532) );
  INV_X1 U10463 ( .A(n9093), .ZN(n9097) );
  AOI21_X1 U10464 ( .B1(n9094), .B2(n9097), .A(P1_U3086), .ZN(n9096) );
  INV_X1 U10465 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9095) );
  NOR2_X1 U10466 ( .A1(n9096), .A2(n9095), .ZN(n9099) );
  NOR3_X1 U10467 ( .A1(n9727), .A2(P1_REG3_REG_17__SCAN_IN), .A3(n9097), .ZN(
        n9098) );
  AOI211_X1 U10468 ( .C1(n9719), .C2(n9532), .A(n9099), .B(n9098), .ZN(n9100)
         );
  OAI211_X1 U10469 ( .C1(n4855), .C2(n9722), .A(n9101), .B(n9100), .ZN(
        P1_U3228) );
  AND3_X1 U10470 ( .A1(n9104), .A2(n9103), .A3(n9102), .ZN(n9105) );
  OAI21_X1 U10471 ( .B1(n9106), .B2(n9105), .A(n9724), .ZN(n9113) );
  NAND2_X1 U10472 ( .A1(n9145), .A2(n9181), .ZN(n9108) );
  NAND2_X1 U10473 ( .A1(n9195), .A2(n9180), .ZN(n9107) );
  NAND2_X1 U10474 ( .A1(n9108), .A2(n9107), .ZN(n9426) );
  INV_X1 U10475 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9109) );
  OAI22_X1 U10476 ( .A1(n9110), .A2(n9727), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9109), .ZN(n9111) );
  AOI21_X1 U10477 ( .B1(n9426), .B2(n9719), .A(n9111), .ZN(n9112) );
  OAI211_X1 U10478 ( .C1(n9436), .C2(n9722), .A(n9113), .B(n9112), .ZN(
        P1_U3229) );
  INV_X1 U10479 ( .A(n9115), .ZN(n9117) );
  NAND2_X1 U10480 ( .A1(n9117), .A2(n9116), .ZN(n9118) );
  XNOR2_X1 U10481 ( .A(n9114), .B(n9118), .ZN(n9124) );
  AND2_X1 U10482 ( .A1(n9200), .A2(n9181), .ZN(n9119) );
  AOI21_X1 U10483 ( .B1(n9198), .B2(n9180), .A(n9119), .ZN(n9489) );
  NOR2_X1 U10484 ( .A1(n9489), .A2(n9694), .ZN(n9122) );
  OAI22_X1 U10485 ( .A1(n9727), .A2(n9494), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9120), .ZN(n9121) );
  AOI211_X1 U10486 ( .C1(n9623), .C2(n9703), .A(n9122), .B(n9121), .ZN(n9123)
         );
  OAI21_X1 U10487 ( .B1(n9124), .B2(n9699), .A(n9123), .ZN(P1_U3233) );
  NAND2_X1 U10488 ( .A1(n9125), .A2(n9719), .ZN(n9127) );
  OAI211_X1 U10489 ( .C1(n9727), .C2(n9128), .A(n9127), .B(n9126), .ZN(n9136)
         );
  INV_X1 U10490 ( .A(n9129), .ZN(n9130) );
  NAND3_X1 U10491 ( .A1(n9132), .A2(n9131), .A3(n9130), .ZN(n9133) );
  AOI21_X1 U10492 ( .B1(n9134), .B2(n9133), .A(n9699), .ZN(n9135) );
  AOI211_X1 U10493 ( .C1(n9137), .C2(n9703), .A(n9136), .B(n9135), .ZN(n9138)
         );
  INV_X1 U10494 ( .A(n9138), .ZN(P1_U3234) );
  INV_X1 U10495 ( .A(n9139), .ZN(n9144) );
  OAI21_X1 U10496 ( .B1(n9141), .B2(n9143), .A(n9140), .ZN(n9142) );
  OAI211_X1 U10497 ( .C1(n9144), .C2(n9143), .A(n9724), .B(n9142), .ZN(n9151)
         );
  NAND2_X1 U10498 ( .A1(n9145), .A2(n9180), .ZN(n9147) );
  NAND2_X1 U10499 ( .A1(n9198), .A2(n9181), .ZN(n9146) );
  NAND2_X1 U10500 ( .A1(n9147), .A2(n9146), .ZN(n9464) );
  INV_X1 U10501 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9148) );
  OAI22_X1 U10502 ( .A1(n9458), .A2(n9727), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9148), .ZN(n9149) );
  AOI21_X1 U10503 ( .B1(n9464), .B2(n9719), .A(n9149), .ZN(n9150) );
  OAI211_X1 U10504 ( .C1(n9461), .C2(n9722), .A(n9151), .B(n9150), .ZN(
        P1_U3235) );
  INV_X1 U10505 ( .A(n9152), .ZN(n9157) );
  AOI21_X1 U10506 ( .B1(n9154), .B2(n9156), .A(n9153), .ZN(n9155) );
  AOI21_X1 U10507 ( .B1(n9157), .B2(n9156), .A(n9155), .ZN(n9164) );
  INV_X1 U10508 ( .A(n9516), .ZN(n9161) );
  NAND2_X1 U10509 ( .A1(n9200), .A2(n9180), .ZN(n9159) );
  NAND2_X1 U10510 ( .A1(n9202), .A2(n9181), .ZN(n9158) );
  NAND2_X1 U10511 ( .A1(n9159), .A2(n9158), .ZN(n9521) );
  AOI22_X1 U10512 ( .A1(n9719), .A2(n9521), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n9160) );
  OAI21_X1 U10513 ( .B1(n9161), .B2(n9727), .A(n9160), .ZN(n9162) );
  AOI21_X1 U10514 ( .B1(n9632), .B2(n9703), .A(n9162), .ZN(n9163) );
  OAI21_X1 U10515 ( .B1(n9164), .B2(n9699), .A(n9163), .ZN(P1_U3238) );
  OAI21_X1 U10516 ( .B1(n4530), .B2(n9166), .A(n9165), .ZN(n9167) );
  NAND3_X1 U10517 ( .A1(n4563), .A2(n9724), .A3(n9167), .ZN(n9175) );
  OR2_X1 U10518 ( .A1(n9169), .A2(n9168), .ZN(n9171) );
  NAND2_X1 U10519 ( .A1(n9195), .A2(n9181), .ZN(n9170) );
  AND2_X1 U10520 ( .A1(n9171), .A2(n9170), .ZN(n9398) );
  OAI22_X1 U10521 ( .A1(n9398), .A2(n9694), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9172), .ZN(n9173) );
  AOI21_X1 U10522 ( .B1(n9403), .B2(n9187), .A(n9173), .ZN(n9174) );
  OAI211_X1 U10523 ( .C1(n9654), .C2(n9722), .A(n9175), .B(n9174), .ZN(
        P1_U3240) );
  XOR2_X1 U10524 ( .A(n9177), .B(n9176), .Z(n9178) );
  XNOR2_X1 U10525 ( .A(n9179), .B(n9178), .ZN(n9189) );
  NAND2_X1 U10526 ( .A1(n9203), .A2(n9180), .ZN(n9183) );
  NAND2_X1 U10527 ( .A1(n4922), .A2(n9181), .ZN(n9182) );
  AND2_X1 U10528 ( .A1(n9183), .A2(n9182), .ZN(n9559) );
  OAI22_X1 U10529 ( .A1(n9559), .A2(n9694), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9184), .ZN(n9186) );
  NOR2_X1 U10530 ( .A1(n9709), .A2(n9722), .ZN(n9185) );
  AOI211_X1 U10531 ( .C1(n9187), .C2(n9564), .A(n9186), .B(n9185), .ZN(n9188)
         );
  OAI21_X1 U10532 ( .B1(n9189), .B2(n9699), .A(n9188), .ZN(P1_U3241) );
  MUX2_X1 U10533 ( .A(n9190), .B(P1_DATAO_REG_31__SCAN_IN), .S(n9217), .Z(
        P1_U3585) );
  MUX2_X1 U10534 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9191), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10535 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9192), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10536 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9193), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10537 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9194), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10538 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9195), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10539 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9196), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10540 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9197), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10541 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9198), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10542 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9199), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10543 ( .A(n9200), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9217), .Z(
        P1_U3573) );
  MUX2_X1 U10544 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9201), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10545 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9202), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10546 ( .A(n9203), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9217), .Z(
        P1_U3570) );
  MUX2_X1 U10547 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9204), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10548 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n4922), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10549 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9205), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10550 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9206), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10551 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9207), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10552 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9208), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10553 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9209), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10554 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9210), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10555 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9211), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10556 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9212), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10557 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9213), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10558 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9214), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10559 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9215), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10560 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9216), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10561 ( .A(n9218), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9217), .Z(
        P1_U3554) );
  INV_X1 U10562 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10103) );
  OAI22_X1 U10563 ( .A1(n9263), .A2(n10103), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9219), .ZN(n9220) );
  AOI21_X1 U10564 ( .B1(n9221), .B2(n9265), .A(n9220), .ZN(n9229) );
  OAI211_X1 U10565 ( .C1(n9231), .C2(n9223), .A(n9319), .B(n9222), .ZN(n9228)
         );
  OAI211_X1 U10566 ( .C1(n9226), .C2(n9225), .A(n9309), .B(n9224), .ZN(n9227)
         );
  NAND3_X1 U10567 ( .A1(n9229), .A2(n9228), .A3(n9227), .ZN(P1_U3244) );
  MUX2_X1 U10568 ( .A(n9231), .B(n9230), .S(n9684), .Z(n9233) );
  NAND2_X1 U10569 ( .A1(n9233), .A2(n9232), .ZN(n9234) );
  OAI211_X1 U10570 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9235), .A(n9234), .B(
        P1_U3973), .ZN(n9279) );
  INV_X1 U10571 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9237) );
  OAI22_X1 U10572 ( .A1(n9263), .A2(n9237), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9236), .ZN(n9238) );
  AOI21_X1 U10573 ( .B1(n9239), .B2(n9265), .A(n9238), .ZN(n9247) );
  OAI211_X1 U10574 ( .C1(n9241), .C2(n9240), .A(n9309), .B(n9253), .ZN(n9246)
         );
  OAI211_X1 U10575 ( .C1(n9244), .C2(n9243), .A(n9319), .B(n9242), .ZN(n9245)
         );
  NAND4_X1 U10576 ( .A1(n9279), .A2(n9247), .A3(n9246), .A4(n9245), .ZN(
        P1_U3245) );
  OAI211_X1 U10577 ( .C1(n9250), .C2(n9249), .A(n9319), .B(n9248), .ZN(n9260)
         );
  MUX2_X1 U10578 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6758), .S(n9251), .Z(n9254)
         );
  NAND3_X1 U10579 ( .A1(n9254), .A2(n9253), .A3(n9252), .ZN(n9255) );
  NAND3_X1 U10580 ( .A1(n9309), .A2(n9273), .A3(n9255), .ZN(n9259) );
  AOI22_X1 U10581 ( .A1(n9349), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(P1_U3086), .ZN(n9258) );
  NAND2_X1 U10582 ( .A1(n9265), .A2(n9256), .ZN(n9257) );
  NAND4_X1 U10583 ( .A1(n9260), .A2(n9259), .A3(n9258), .A4(n9257), .ZN(
        P1_U3246) );
  INV_X1 U10584 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9262) );
  OAI21_X1 U10585 ( .B1(n9263), .B2(n9262), .A(n9261), .ZN(n9264) );
  AOI21_X1 U10586 ( .B1(n9266), .B2(n9265), .A(n9264), .ZN(n9278) );
  OAI211_X1 U10587 ( .C1(n9269), .C2(n9268), .A(n9319), .B(n9267), .ZN(n9277)
         );
  MUX2_X1 U10588 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6761), .S(n9270), .Z(n9271)
         );
  NAND3_X1 U10589 ( .A1(n9273), .A2(n9272), .A3(n9271), .ZN(n9275) );
  NAND3_X1 U10590 ( .A1(n9309), .A2(n9275), .A3(n9274), .ZN(n9276) );
  NAND4_X1 U10591 ( .A1(n9279), .A2(n9278), .A3(n9277), .A4(n9276), .ZN(
        P1_U3247) );
  AND2_X1 U10592 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9282) );
  NOR2_X1 U10593 ( .A1(n9337), .A2(n9280), .ZN(n9281) );
  AOI211_X1 U10594 ( .C1(n9349), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n9282), .B(
        n9281), .ZN(n9290) );
  OAI211_X1 U10595 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n9284), .A(n9309), .B(
        n9283), .ZN(n9289) );
  AOI211_X1 U10596 ( .C1(n9567), .C2(n9286), .A(n9285), .B(n9341), .ZN(n9287)
         );
  INV_X1 U10597 ( .A(n9287), .ZN(n9288) );
  NAND3_X1 U10598 ( .A1(n9290), .A2(n9289), .A3(n9288), .ZN(P1_U3258) );
  XNOR2_X1 U10599 ( .A(n9313), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n9316) );
  XNOR2_X1 U10600 ( .A(n9316), .B(n9315), .ZN(n9300) );
  NAND2_X1 U10601 ( .A1(n9313), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9293) );
  OAI21_X1 U10602 ( .B1(n9313), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9293), .ZN(
        n9298) );
  AOI21_X1 U10603 ( .B1(n9295), .B2(n7863), .A(n9294), .ZN(n9296) );
  INV_X1 U10604 ( .A(n9296), .ZN(n9297) );
  NAND2_X1 U10605 ( .A1(n9298), .A2(n9297), .ZN(n9308) );
  OAI21_X1 U10606 ( .B1(n9298), .B2(n9297), .A(n9308), .ZN(n9299) );
  AOI22_X1 U10607 ( .A1(n9319), .A2(n9300), .B1(n9309), .B2(n9299), .ZN(n9302)
         );
  AOI22_X1 U10608 ( .A1(n9349), .A2(P1_ADDR_REG_17__SCAN_IN), .B1(
        P1_REG3_REG_17__SCAN_IN), .B2(P1_U3086), .ZN(n9301) );
  OAI211_X1 U10609 ( .C1(n9313), .C2(n9337), .A(n9302), .B(n9301), .ZN(
        P1_U3260) );
  AND2_X1 U10610 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9305) );
  NOR2_X1 U10611 ( .A1(n9337), .A2(n9303), .ZN(n9304) );
  AOI211_X1 U10612 ( .C1(n9349), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9305), .B(
        n9304), .ZN(n9324) );
  INV_X1 U10613 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9306) );
  XNOR2_X1 U10614 ( .A(n9329), .B(n9306), .ZN(n9311) );
  INV_X1 U10615 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9639) );
  NAND2_X1 U10616 ( .A1(n9313), .A2(n9639), .ZN(n9307) );
  AND2_X1 U10617 ( .A1(n9308), .A2(n9307), .ZN(n9310) );
  NAND2_X1 U10618 ( .A1(n9310), .A2(n9311), .ZN(n9331) );
  OAI211_X1 U10619 ( .C1(n9311), .C2(n9310), .A(n9309), .B(n9331), .ZN(n9323)
         );
  INV_X1 U10620 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9312) );
  AND2_X1 U10621 ( .A1(n9313), .A2(n9312), .ZN(n9314) );
  AOI21_X1 U10622 ( .B1(n9316), .B2(n9315), .A(n9314), .ZN(n9321) );
  INV_X1 U10623 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9318) );
  NAND2_X1 U10624 ( .A1(n9329), .A2(n9318), .ZN(n9317) );
  OAI21_X1 U10625 ( .B1(n9329), .B2(n9318), .A(n9317), .ZN(n9320) );
  NAND2_X1 U10626 ( .A1(n9321), .A2(n9320), .ZN(n9326) );
  OAI211_X1 U10627 ( .C1(n9321), .C2(n9320), .A(n9319), .B(n9326), .ZN(n9322)
         );
  NAND3_X1 U10628 ( .A1(n9324), .A2(n9323), .A3(n9322), .ZN(P1_U3261) );
  NAND2_X1 U10629 ( .A1(n9329), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9325) );
  NAND2_X1 U10630 ( .A1(n9326), .A2(n9325), .ZN(n9328) );
  INV_X1 U10631 ( .A(n9340), .ZN(n9335) );
  NAND2_X1 U10632 ( .A1(n9329), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9330) );
  NAND2_X1 U10633 ( .A1(n9331), .A2(n9330), .ZN(n9333) );
  XNOR2_X1 U10634 ( .A(n9333), .B(n9332), .ZN(n9338) );
  INV_X1 U10635 ( .A(n9338), .ZN(n9334) );
  OAI22_X1 U10636 ( .A1(n9335), .A2(n9341), .B1(n9339), .B2(n9334), .ZN(n9336)
         );
  INV_X1 U10637 ( .A(n9336), .ZN(n9346) );
  OAI21_X1 U10638 ( .B1(n9339), .B2(n9338), .A(n9337), .ZN(n9343) );
  NOR2_X1 U10639 ( .A1(n9341), .A2(n9340), .ZN(n9342) );
  NOR2_X1 U10640 ( .A1(n9343), .A2(n9342), .ZN(n9345) );
  MUX2_X1 U10641 ( .A(n9346), .B(n9345), .S(n9344), .Z(n9351) );
  INV_X1 U10642 ( .A(n9347), .ZN(n9348) );
  AOI21_X1 U10643 ( .B1(n9349), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9348), .ZN(
        n9350) );
  NAND2_X1 U10644 ( .A1(n9351), .A2(n9350), .ZN(P1_U3262) );
  NAND2_X1 U10645 ( .A1(n9352), .A2(n9769), .ZN(n9355) );
  INV_X1 U10646 ( .A(n9353), .ZN(n9580) );
  NOR2_X1 U10647 ( .A1(n9580), .A2(n9773), .ZN(n9362) );
  AOI21_X1 U10648 ( .B1(n9773), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9362), .ZN(
        n9354) );
  OAI211_X1 U10649 ( .C1(n9579), .C2(n9761), .A(n9355), .B(n9354), .ZN(
        P1_U3263) );
  NAND2_X1 U10650 ( .A1(n9357), .A2(n9356), .ZN(n9358) );
  NAND2_X1 U10651 ( .A1(n9358), .A2(n9765), .ZN(n9359) );
  NOR2_X1 U10652 ( .A1(n9649), .A2(n9761), .ZN(n9361) );
  AOI211_X1 U10653 ( .C1(n9773), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9362), .B(
        n9361), .ZN(n9363) );
  OAI21_X1 U10654 ( .B1(n9581), .B2(n9570), .A(n9363), .ZN(P1_U3264) );
  INV_X1 U10655 ( .A(n9364), .ZN(n9373) );
  NAND2_X1 U10656 ( .A1(n9365), .A2(n9769), .ZN(n9368) );
  AOI22_X1 U10657 ( .A1(n9773), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9366), .B2(
        n9759), .ZN(n9367) );
  OAI211_X1 U10658 ( .C1(n9369), .C2(n9761), .A(n9368), .B(n9367), .ZN(n9370)
         );
  AOI21_X1 U10659 ( .B1(n9371), .B2(n9770), .A(n9370), .ZN(n9372) );
  OAI21_X1 U10660 ( .B1(n9373), .B2(n9773), .A(n9372), .ZN(P1_U3356) );
  NAND2_X1 U10661 ( .A1(n9374), .A2(n9770), .ZN(n9380) );
  AOI22_X1 U10662 ( .A1(n9730), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9375), .B2(
        n9759), .ZN(n9376) );
  OAI21_X1 U10663 ( .B1(n4510), .B2(n9761), .A(n9376), .ZN(n9377) );
  AOI21_X1 U10664 ( .B1(n9378), .B2(n9769), .A(n9377), .ZN(n9379) );
  OAI211_X1 U10665 ( .C1(n5139), .C2(n9773), .A(n9380), .B(n9379), .ZN(
        P1_U3265) );
  XNOR2_X1 U10666 ( .A(n9381), .B(n4937), .ZN(n9384) );
  INV_X1 U10667 ( .A(n9382), .ZN(n9383) );
  AOI21_X1 U10668 ( .B1(n9384), .B2(n9756), .A(n9383), .ZN(n9588) );
  AOI21_X1 U10669 ( .B1(n9390), .B2(n4846), .A(n9850), .ZN(n9388) );
  NAND2_X1 U10670 ( .A1(n9388), .A2(n9387), .ZN(n9587) );
  AOI22_X1 U10671 ( .A1(n9773), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9389), .B2(
        n9759), .ZN(n9392) );
  NAND2_X1 U10672 ( .A1(n9390), .A2(n9731), .ZN(n9391) );
  OAI211_X1 U10673 ( .C1(n9587), .C2(n9570), .A(n9392), .B(n9391), .ZN(n9393)
         );
  AOI21_X1 U10674 ( .B1(n9586), .B2(n9770), .A(n9393), .ZN(n9394) );
  OAI21_X1 U10675 ( .B1(n9773), .B2(n9588), .A(n9394), .ZN(P1_U3266) );
  OAI21_X1 U10676 ( .B1(n9400), .B2(n9396), .A(n9395), .ZN(n9397) );
  NAND2_X1 U10677 ( .A1(n9397), .A2(n9756), .ZN(n9399) );
  NAND2_X1 U10678 ( .A1(n9399), .A2(n9398), .ZN(n9590) );
  INV_X1 U10679 ( .A(n9590), .ZN(n9408) );
  XNOR2_X1 U10680 ( .A(n9401), .B(n9400), .ZN(n9592) );
  NAND2_X1 U10681 ( .A1(n9592), .A2(n9770), .ZN(n9407) );
  AOI211_X1 U10682 ( .C1(n9402), .C2(n9415), .A(n9850), .B(n9386), .ZN(n9591)
         );
  AOI22_X1 U10683 ( .A1(n9730), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9403), .B2(
        n9759), .ZN(n9404) );
  OAI21_X1 U10684 ( .B1(n9654), .B2(n9761), .A(n9404), .ZN(n9405) );
  AOI21_X1 U10685 ( .B1(n9591), .B2(n9769), .A(n9405), .ZN(n9406) );
  OAI211_X1 U10686 ( .C1(n9773), .C2(n9408), .A(n9407), .B(n9406), .ZN(
        P1_U3267) );
  XNOR2_X1 U10687 ( .A(n9409), .B(n9413), .ZN(n9410) );
  NAND2_X1 U10688 ( .A1(n9410), .A2(n9756), .ZN(n9412) );
  NAND2_X1 U10689 ( .A1(n9412), .A2(n9411), .ZN(n9595) );
  INV_X1 U10690 ( .A(n9595), .ZN(n9424) );
  XOR2_X1 U10691 ( .A(n9414), .B(n9413), .Z(n9597) );
  NAND2_X1 U10692 ( .A1(n9597), .A2(n9770), .ZN(n9423) );
  INV_X1 U10693 ( .A(n9432), .ZN(n9417) );
  INV_X1 U10694 ( .A(n9415), .ZN(n9416) );
  AOI211_X1 U10695 ( .C1(n9418), .C2(n9417), .A(n9850), .B(n9416), .ZN(n9596)
         );
  AOI22_X1 U10696 ( .A1(n9730), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9419), .B2(
        n9759), .ZN(n9420) );
  OAI21_X1 U10697 ( .B1(n9658), .B2(n9761), .A(n9420), .ZN(n9421) );
  AOI21_X1 U10698 ( .B1(n9596), .B2(n9769), .A(n9421), .ZN(n9422) );
  OAI211_X1 U10699 ( .C1(n9773), .C2(n9424), .A(n9423), .B(n9422), .ZN(
        P1_U3268) );
  AOI21_X1 U10700 ( .B1(n9425), .B2(n9429), .A(n9504), .ZN(n9428) );
  AOI21_X1 U10701 ( .B1(n9428), .B2(n9427), .A(n9426), .ZN(n9604) );
  OR2_X1 U10702 ( .A1(n9430), .A2(n9429), .ZN(n9600) );
  NAND3_X1 U10703 ( .A1(n9600), .A2(n9770), .A3(n9431), .ZN(n9440) );
  INV_X1 U10704 ( .A(n9446), .ZN(n9433) );
  AOI21_X1 U10705 ( .B1(n9601), .B2(n9433), .A(n9432), .ZN(n9602) );
  AOI22_X1 U10706 ( .A1(n9434), .A2(n9759), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9773), .ZN(n9435) );
  OAI21_X1 U10707 ( .B1(n9436), .B2(n9761), .A(n9435), .ZN(n9437) );
  AOI21_X1 U10708 ( .B1(n9602), .B2(n9438), .A(n9437), .ZN(n9439) );
  OAI211_X1 U10709 ( .C1(n9773), .C2(n9604), .A(n9440), .B(n9439), .ZN(
        P1_U3269) );
  XOR2_X1 U10710 ( .A(n9441), .B(n9443), .Z(n9610) );
  XOR2_X1 U10711 ( .A(n9442), .B(n9443), .Z(n9445) );
  OAI21_X1 U10712 ( .B1(n9445), .B2(n9504), .A(n9444), .ZN(n9606) );
  INV_X1 U10713 ( .A(n9608), .ZN(n9450) );
  AOI211_X1 U10714 ( .C1(n9608), .C2(n9455), .A(n9850), .B(n9446), .ZN(n9607)
         );
  NAND2_X1 U10715 ( .A1(n9607), .A2(n9769), .ZN(n9449) );
  AOI22_X1 U10716 ( .A1(n9447), .A2(n9759), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9773), .ZN(n9448) );
  OAI211_X1 U10717 ( .C1(n9450), .C2(n9761), .A(n9449), .B(n9448), .ZN(n9451)
         );
  AOI21_X1 U10718 ( .B1(n9452), .B2(n9606), .A(n9451), .ZN(n9453) );
  OAI21_X1 U10719 ( .B1(n9610), .B2(n9556), .A(n9453), .ZN(P1_U3270) );
  XNOR2_X1 U10720 ( .A(n9454), .B(n9462), .ZN(n9615) );
  INV_X1 U10721 ( .A(n9477), .ZN(n9457) );
  INV_X1 U10722 ( .A(n9455), .ZN(n9456) );
  AOI211_X1 U10723 ( .C1(n9612), .C2(n9457), .A(n9850), .B(n9456), .ZN(n9611)
         );
  INV_X1 U10724 ( .A(n9458), .ZN(n9459) );
  AOI22_X1 U10725 ( .A1(n9459), .A2(n9759), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9773), .ZN(n9460) );
  OAI21_X1 U10726 ( .B1(n9461), .B2(n9761), .A(n9460), .ZN(n9467) );
  XNOR2_X1 U10727 ( .A(n9463), .B(n9462), .ZN(n9465) );
  AOI21_X1 U10728 ( .B1(n9465), .B2(n9756), .A(n9464), .ZN(n9614) );
  NOR2_X1 U10729 ( .A1(n9614), .A2(n9730), .ZN(n9466) );
  AOI211_X1 U10730 ( .C1(n9611), .C2(n9769), .A(n9467), .B(n9466), .ZN(n9468)
         );
  OAI21_X1 U10731 ( .B1(n9615), .B2(n9556), .A(n9468), .ZN(P1_U3271) );
  XNOR2_X1 U10732 ( .A(n9470), .B(n9469), .ZN(n9618) );
  INV_X1 U10733 ( .A(n9618), .ZN(n9485) );
  INV_X1 U10734 ( .A(n9471), .ZN(n9472) );
  AOI21_X1 U10735 ( .B1(n9474), .B2(n9473), .A(n9472), .ZN(n9476) );
  OAI21_X1 U10736 ( .B1(n9476), .B2(n9504), .A(n9475), .ZN(n9616) );
  INV_X1 U10737 ( .A(n9478), .ZN(n9665) );
  AOI211_X1 U10738 ( .C1(n9478), .C2(n9492), .A(n9850), .B(n9477), .ZN(n9617)
         );
  NAND2_X1 U10739 ( .A1(n9617), .A2(n9769), .ZN(n9482) );
  INV_X1 U10740 ( .A(n9479), .ZN(n9480) );
  AOI22_X1 U10741 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(n9730), .B1(n9480), .B2(
        n9759), .ZN(n9481) );
  OAI211_X1 U10742 ( .C1(n9665), .C2(n9761), .A(n9482), .B(n9481), .ZN(n9483)
         );
  AOI21_X1 U10743 ( .B1(n9616), .B2(n9452), .A(n9483), .ZN(n9484) );
  OAI21_X1 U10744 ( .B1(n9485), .B2(n9556), .A(n9484), .ZN(P1_U3272) );
  XNOR2_X1 U10745 ( .A(n9486), .B(n9487), .ZN(n9625) );
  XNOR2_X1 U10746 ( .A(n9488), .B(n9487), .ZN(n9490) );
  OAI21_X1 U10747 ( .B1(n9490), .B2(n9504), .A(n9489), .ZN(n9621) );
  INV_X1 U10748 ( .A(n9492), .ZN(n9493) );
  AOI211_X1 U10749 ( .C1(n9623), .C2(n9506), .A(n9850), .B(n9493), .ZN(n9622)
         );
  NAND2_X1 U10750 ( .A1(n9622), .A2(n9769), .ZN(n9497) );
  INV_X1 U10751 ( .A(n9494), .ZN(n9495) );
  AOI22_X1 U10752 ( .A1(n9730), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9495), .B2(
        n9759), .ZN(n9496) );
  OAI211_X1 U10753 ( .C1(n5747), .C2(n9761), .A(n9497), .B(n9496), .ZN(n9498)
         );
  AOI21_X1 U10754 ( .B1(n9621), .B2(n9452), .A(n9498), .ZN(n9499) );
  OAI21_X1 U10755 ( .B1(n9625), .B2(n9556), .A(n9499), .ZN(P1_U3273) );
  XNOR2_X1 U10756 ( .A(n9500), .B(n9501), .ZN(n9630) );
  XNOR2_X1 U10757 ( .A(n9502), .B(n9501), .ZN(n9505) );
  OAI21_X1 U10758 ( .B1(n9505), .B2(n9504), .A(n9503), .ZN(n9626) );
  AOI211_X1 U10759 ( .C1(n9628), .C2(n9514), .A(n9850), .B(n9491), .ZN(n9627)
         );
  NAND2_X1 U10760 ( .A1(n9627), .A2(n9769), .ZN(n9509) );
  AOI22_X1 U10761 ( .A1(n9730), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9507), .B2(
        n9759), .ZN(n9508) );
  OAI211_X1 U10762 ( .C1(n9510), .C2(n9761), .A(n9509), .B(n9508), .ZN(n9511)
         );
  AOI21_X1 U10763 ( .B1(n9626), .B2(n9452), .A(n9511), .ZN(n9512) );
  OAI21_X1 U10764 ( .B1(n9630), .B2(n9556), .A(n9512), .ZN(P1_U3274) );
  XOR2_X1 U10765 ( .A(n9519), .B(n9513), .Z(n9635) );
  INV_X1 U10766 ( .A(n9514), .ZN(n9515) );
  AOI211_X1 U10767 ( .C1(n9632), .C2(n4857), .A(n9850), .B(n9515), .ZN(n9631)
         );
  AOI22_X1 U10768 ( .A1(n9730), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9516), .B2(
        n9759), .ZN(n9517) );
  OAI21_X1 U10769 ( .B1(n9518), .B2(n9761), .A(n9517), .ZN(n9524) );
  XNOR2_X1 U10770 ( .A(n9520), .B(n9519), .ZN(n9522) );
  AOI21_X1 U10771 ( .B1(n9522), .B2(n9756), .A(n9521), .ZN(n9634) );
  NOR2_X1 U10772 ( .A1(n9634), .A2(n9773), .ZN(n9523) );
  AOI211_X1 U10773 ( .C1(n9631), .C2(n9769), .A(n9524), .B(n9523), .ZN(n9525)
         );
  OAI21_X1 U10774 ( .B1(n9635), .B2(n9556), .A(n9525), .ZN(P1_U3275) );
  XNOR2_X1 U10775 ( .A(n9527), .B(n9526), .ZN(n9638) );
  INV_X1 U10776 ( .A(n9638), .ZN(n9541) );
  NAND2_X1 U10777 ( .A1(n9529), .A2(n9528), .ZN(n9530) );
  NAND3_X1 U10778 ( .A1(n9531), .A2(n9756), .A3(n9530), .ZN(n9534) );
  INV_X1 U10779 ( .A(n9532), .ZN(n9533) );
  NAND2_X1 U10780 ( .A1(n9534), .A2(n9533), .ZN(n9636) );
  AOI211_X1 U10781 ( .C1(n9536), .C2(n9549), .A(n9850), .B(n9535), .ZN(n9637)
         );
  NAND2_X1 U10782 ( .A1(n9637), .A2(n9769), .ZN(n9538) );
  AOI22_X1 U10783 ( .A1(n9730), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n5140), .B2(
        n9759), .ZN(n9537) );
  OAI211_X1 U10784 ( .C1(n4855), .C2(n9761), .A(n9538), .B(n9537), .ZN(n9539)
         );
  AOI21_X1 U10785 ( .B1(n9452), .B2(n9636), .A(n9539), .ZN(n9540) );
  OAI21_X1 U10786 ( .B1(n9541), .B2(n9556), .A(n9540), .ZN(P1_U3276) );
  XNOR2_X1 U10787 ( .A(n9542), .B(n4647), .ZN(n9643) );
  INV_X1 U10788 ( .A(n9643), .ZN(n9557) );
  OAI21_X1 U10789 ( .B1(n4647), .B2(n9544), .A(n9543), .ZN(n9545) );
  NAND2_X1 U10790 ( .A1(n9545), .A2(n9756), .ZN(n9547) );
  NAND2_X1 U10791 ( .A1(n9547), .A2(n9546), .ZN(n9641) );
  INV_X1 U10792 ( .A(n9548), .ZN(n9676) );
  AOI21_X1 U10793 ( .B1(n9548), .B2(n9568), .A(n9850), .ZN(n9550) );
  AND2_X1 U10794 ( .A1(n9550), .A2(n9549), .ZN(n9642) );
  NAND2_X1 U10795 ( .A1(n9642), .A2(n9769), .ZN(n9553) );
  AOI22_X1 U10796 ( .A1(n9730), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9551), .B2(
        n9759), .ZN(n9552) );
  OAI211_X1 U10797 ( .C1(n9676), .C2(n9761), .A(n9553), .B(n9552), .ZN(n9554)
         );
  AOI21_X1 U10798 ( .B1(n9641), .B2(n9452), .A(n9554), .ZN(n9555) );
  OAI21_X1 U10799 ( .B1(n9557), .B2(n9556), .A(n9555), .ZN(P1_U3277) );
  XNOR2_X1 U10800 ( .A(n9558), .B(n9562), .ZN(n9561) );
  INV_X1 U10801 ( .A(n9559), .ZN(n9560) );
  AOI21_X1 U10802 ( .B1(n9561), .B2(n9756), .A(n9560), .ZN(n9708) );
  XOR2_X1 U10803 ( .A(n9563), .B(n9562), .Z(n9711) );
  NAND2_X1 U10804 ( .A1(n9711), .A2(n9770), .ZN(n9575) );
  INV_X1 U10805 ( .A(n9564), .ZN(n9566) );
  OAI22_X1 U10806 ( .A1(n9452), .A2(n9567), .B1(n9566), .B2(n9565), .ZN(n9572)
         );
  OAI211_X1 U10807 ( .C1(n9709), .C2(n9569), .A(n9765), .B(n9568), .ZN(n9707)
         );
  NOR2_X1 U10808 ( .A1(n9707), .A2(n9570), .ZN(n9571) );
  AOI211_X1 U10809 ( .C1(n9731), .C2(n9573), .A(n9572), .B(n9571), .ZN(n9574)
         );
  OAI211_X1 U10810 ( .C1(n9773), .C2(n9708), .A(n9575), .B(n9574), .ZN(
        P1_U3278) );
  INV_X1 U10811 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9577) );
  MUX2_X1 U10812 ( .A(n9577), .B(n9576), .S(n9875), .Z(n9578) );
  OAI21_X1 U10813 ( .B1(n9579), .B2(n9645), .A(n9578), .ZN(P1_U3553) );
  NAND2_X1 U10814 ( .A1(n9581), .A2(n9580), .ZN(n9646) );
  MUX2_X1 U10815 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9646), .S(n9875), .Z(n9582) );
  INV_X1 U10816 ( .A(n9582), .ZN(n9583) );
  OAI21_X1 U10817 ( .B1(n9649), .B2(n9645), .A(n9583), .ZN(P1_U3552) );
  INV_X1 U10818 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9585) );
  NAND2_X1 U10819 ( .A1(n9586), .A2(n9845), .ZN(n9589) );
  INV_X1 U10820 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9593) );
  AOI211_X1 U10821 ( .C1(n9592), .C2(n9845), .A(n9591), .B(n9590), .ZN(n9651)
         );
  MUX2_X1 U10822 ( .A(n9593), .B(n9651), .S(n9875), .Z(n9594) );
  OAI21_X1 U10823 ( .B1(n9654), .B2(n9645), .A(n9594), .ZN(P1_U3548) );
  INV_X1 U10824 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9598) );
  AOI211_X1 U10825 ( .C1(n9597), .C2(n9845), .A(n9596), .B(n9595), .ZN(n9655)
         );
  MUX2_X1 U10826 ( .A(n9598), .B(n9655), .S(n9875), .Z(n9599) );
  OAI21_X1 U10827 ( .B1(n9658), .B2(n9645), .A(n9599), .ZN(P1_U3547) );
  NAND3_X1 U10828 ( .A1(n9600), .A2(n9845), .A3(n9431), .ZN(n9605) );
  AOI22_X1 U10829 ( .A1(n9602), .A2(n9765), .B1(n9801), .B2(n9601), .ZN(n9603)
         );
  NAND3_X1 U10830 ( .A1(n9605), .A2(n9604), .A3(n9603), .ZN(n9659) );
  MUX2_X1 U10831 ( .A(n9659), .B(P1_REG1_REG_24__SCAN_IN), .S(n5819), .Z(
        P1_U3546) );
  AOI211_X1 U10832 ( .C1(n9801), .C2(n9608), .A(n9607), .B(n9606), .ZN(n9609)
         );
  OAI21_X1 U10833 ( .B1(n9610), .B2(n9805), .A(n9609), .ZN(n9660) );
  MUX2_X1 U10834 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9660), .S(n9875), .Z(
        P1_U3545) );
  AOI21_X1 U10835 ( .B1(n9801), .B2(n9612), .A(n9611), .ZN(n9613) );
  OAI211_X1 U10836 ( .C1(n9615), .C2(n9805), .A(n9614), .B(n9613), .ZN(n9661)
         );
  MUX2_X1 U10837 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9661), .S(n9875), .Z(
        P1_U3544) );
  INV_X1 U10838 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9619) );
  AOI211_X1 U10839 ( .C1(n9845), .C2(n9618), .A(n9617), .B(n9616), .ZN(n9662)
         );
  MUX2_X1 U10840 ( .A(n9619), .B(n9662), .S(n9875), .Z(n9620) );
  OAI21_X1 U10841 ( .B1(n9665), .B2(n9645), .A(n9620), .ZN(P1_U3543) );
  AOI211_X1 U10842 ( .C1(n9801), .C2(n9623), .A(n9622), .B(n9621), .ZN(n9624)
         );
  OAI21_X1 U10843 ( .B1(n9625), .B2(n9805), .A(n9624), .ZN(n9666) );
  MUX2_X1 U10844 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9666), .S(n9875), .Z(
        P1_U3542) );
  AOI211_X1 U10845 ( .C1(n9801), .C2(n9628), .A(n9627), .B(n9626), .ZN(n9629)
         );
  OAI21_X1 U10846 ( .B1(n9805), .B2(n9630), .A(n9629), .ZN(n9667) );
  MUX2_X1 U10847 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9667), .S(n9875), .Z(
        P1_U3541) );
  AOI21_X1 U10848 ( .B1(n9801), .B2(n9632), .A(n9631), .ZN(n9633) );
  OAI211_X1 U10849 ( .C1(n9635), .C2(n9805), .A(n9634), .B(n9633), .ZN(n9668)
         );
  MUX2_X1 U10850 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9668), .S(n9875), .Z(
        P1_U3540) );
  AOI211_X1 U10851 ( .C1(n9638), .C2(n9845), .A(n9637), .B(n9636), .ZN(n9669)
         );
  MUX2_X1 U10852 ( .A(n9639), .B(n9669), .S(n9875), .Z(n9640) );
  OAI21_X1 U10853 ( .B1(n4855), .B2(n9645), .A(n9640), .ZN(P1_U3539) );
  AOI211_X1 U10854 ( .C1(n9643), .C2(n9845), .A(n9642), .B(n9641), .ZN(n9672)
         );
  MUX2_X1 U10855 ( .A(n7863), .B(n9672), .S(n9875), .Z(n9644) );
  OAI21_X1 U10856 ( .B1(n9676), .B2(n9645), .A(n9644), .ZN(P1_U3538) );
  MUX2_X1 U10857 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9646), .S(n9858), .Z(n9647) );
  INV_X1 U10858 ( .A(n9647), .ZN(n9648) );
  OAI21_X1 U10859 ( .B1(n9649), .B2(n9675), .A(n9648), .ZN(P1_U3520) );
  INV_X1 U10860 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9652) );
  MUX2_X1 U10861 ( .A(n9652), .B(n9651), .S(n9858), .Z(n9653) );
  OAI21_X1 U10862 ( .B1(n9654), .B2(n9675), .A(n9653), .ZN(P1_U3516) );
  INV_X1 U10863 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9656) );
  MUX2_X1 U10864 ( .A(n9656), .B(n9655), .S(n9858), .Z(n9657) );
  OAI21_X1 U10865 ( .B1(n9658), .B2(n9675), .A(n9657), .ZN(P1_U3515) );
  MUX2_X1 U10866 ( .A(n9659), .B(P1_REG0_REG_24__SCAN_IN), .S(n5809), .Z(
        P1_U3514) );
  MUX2_X1 U10867 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9660), .S(n9858), .Z(
        P1_U3513) );
  MUX2_X1 U10868 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9661), .S(n9858), .Z(
        P1_U3512) );
  INV_X1 U10869 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9663) );
  MUX2_X1 U10870 ( .A(n9663), .B(n9662), .S(n9858), .Z(n9664) );
  OAI21_X1 U10871 ( .B1(n9665), .B2(n9675), .A(n9664), .ZN(P1_U3511) );
  MUX2_X1 U10872 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9666), .S(n9858), .Z(
        P1_U3510) );
  MUX2_X1 U10873 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9667), .S(n9858), .Z(
        P1_U3509) );
  MUX2_X1 U10874 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9668), .S(n9858), .Z(
        P1_U3507) );
  INV_X1 U10875 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9670) );
  MUX2_X1 U10876 ( .A(n9670), .B(n9669), .S(n9858), .Z(n9671) );
  OAI21_X1 U10877 ( .B1(n4855), .B2(n9675), .A(n9671), .ZN(P1_U3504) );
  INV_X1 U10878 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9673) );
  MUX2_X1 U10879 ( .A(n9673), .B(n9672), .S(n9858), .Z(n9674) );
  OAI21_X1 U10880 ( .B1(n9676), .B2(n9675), .A(n9674), .ZN(P1_U3501) );
  NOR4_X1 U10881 ( .A1(n9677), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5282), .A4(
        P1_U3086), .ZN(n9678) );
  AOI21_X1 U10882 ( .B1(n9679), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9678), .ZN(
        n9680) );
  OAI21_X1 U10883 ( .B1(n9681), .B2(n9686), .A(n9680), .ZN(P1_U3324) );
  OAI222_X1 U10884 ( .A1(n9687), .A2(n10476), .B1(P1_U3086), .B2(n9682), .C1(
        n9689), .C2(n9683), .ZN(P1_U3326) );
  OAI222_X1 U10885 ( .A1(n9687), .A2(n10317), .B1(n9686), .B2(n9685), .C1(
        n9684), .C2(P1_U3086), .ZN(P1_U3328) );
  OAI222_X1 U10886 ( .A1(n9690), .A2(P1_U3086), .B1(n9689), .B2(n9688), .C1(
        n10490), .C2(n9687), .ZN(P1_U3329) );
  MUX2_X1 U10887 ( .A(n9691), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U10888 ( .A(n9692), .ZN(n9693) );
  OAI21_X1 U10889 ( .B1(n9695), .B2(n9694), .A(n9693), .ZN(n9702) );
  AOI21_X1 U10890 ( .B1(n9698), .B2(n9697), .A(n9696), .ZN(n9700) );
  NOR2_X1 U10891 ( .A1(n9700), .A2(n9699), .ZN(n9701) );
  AOI211_X1 U10892 ( .C1(n9704), .C2(n9703), .A(n9702), .B(n9701), .ZN(n9705)
         );
  OAI21_X1 U10893 ( .B1(n9706), .B2(n9727), .A(n9705), .ZN(P1_U3217) );
  INV_X1 U10894 ( .A(n9801), .ZN(n9848) );
  OAI211_X1 U10895 ( .C1(n9709), .C2(n9848), .A(n9708), .B(n9707), .ZN(n9710)
         );
  AOI21_X1 U10896 ( .B1(n9711), .B2(n9845), .A(n9710), .ZN(n9714) );
  INV_X1 U10897 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9712) );
  AOI22_X1 U10898 ( .A1(n9875), .A2(n9714), .B1(n9712), .B2(n5819), .ZN(
        P1_U3537) );
  INV_X1 U10899 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9713) );
  AOI22_X1 U10900 ( .A1(n9858), .A2(n9714), .B1(n9713), .B2(n5809), .ZN(
        P1_U3498) );
  XNOR2_X1 U10901 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XOR2_X1 U10902 ( .A(n4759), .B(P1_RD_REG_SCAN_IN), .Z(U126) );
  BUF_X1 U10903 ( .A(n9715), .Z(n9716) );
  OAI21_X1 U10904 ( .B1(n9717), .B2(n9716), .A(n7567), .ZN(n9725) );
  AOI21_X1 U10905 ( .B1(n9720), .B2(n9719), .A(n9718), .ZN(n9721) );
  OAI21_X1 U10906 ( .B1(n9830), .B2(n9722), .A(n9721), .ZN(n9723) );
  AOI21_X1 U10907 ( .B1(n9725), .B2(n9724), .A(n9723), .ZN(n9726) );
  OAI21_X1 U10908 ( .B1(n9728), .B2(n9727), .A(n9726), .ZN(P1_U3221) );
  AOI222_X1 U10909 ( .A1(n9732), .A2(n9731), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n9730), .C1(n9759), .C2(n9729), .ZN(n9737) );
  AOI22_X1 U10910 ( .A1(n9735), .A2(n9734), .B1(n9769), .B2(n9733), .ZN(n9736)
         );
  OAI211_X1 U10911 ( .C1(n9773), .C2(n9738), .A(n9737), .B(n9736), .ZN(
        P1_U3282) );
  XNOR2_X1 U10912 ( .A(n9740), .B(n9739), .ZN(n9742) );
  AOI21_X1 U10913 ( .B1(n9742), .B2(n9756), .A(n9741), .ZN(n9810) );
  AOI22_X1 U10914 ( .A1(n9773), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n9743), .B2(
        n9759), .ZN(n9744) );
  OAI21_X1 U10915 ( .B1(n9761), .B2(n9809), .A(n9744), .ZN(n9745) );
  INV_X1 U10916 ( .A(n9745), .ZN(n9751) );
  XNOR2_X1 U10917 ( .A(n9747), .B(n9746), .ZN(n9813) );
  OAI211_X1 U10918 ( .C1(n4589), .C2(n9809), .A(n9765), .B(n9748), .ZN(n9808)
         );
  INV_X1 U10919 ( .A(n9808), .ZN(n9749) );
  AOI22_X1 U10920 ( .A1(n9813), .A2(n9770), .B1(n9769), .B2(n9749), .ZN(n9750)
         );
  OAI211_X1 U10921 ( .C1(n9773), .C2(n9810), .A(n9751), .B(n9750), .ZN(
        P1_U3288) );
  OAI21_X1 U10922 ( .B1(n9754), .B2(n9753), .A(n9752), .ZN(n9757) );
  AOI21_X1 U10923 ( .B1(n9757), .B2(n9756), .A(n9755), .ZN(n9795) );
  AOI22_X1 U10924 ( .A1(n9773), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9759), .B2(
        n9758), .ZN(n9760) );
  OAI21_X1 U10925 ( .B1(n9761), .B2(n9796), .A(n9760), .ZN(n9762) );
  INV_X1 U10926 ( .A(n9762), .ZN(n9772) );
  XNOR2_X1 U10927 ( .A(n9764), .B(n9763), .ZN(n9798) );
  OAI211_X1 U10928 ( .C1(n9767), .C2(n9796), .A(n9766), .B(n9765), .ZN(n9794)
         );
  INV_X1 U10929 ( .A(n9794), .ZN(n9768) );
  AOI22_X1 U10930 ( .A1(n9798), .A2(n9770), .B1(n9769), .B2(n9768), .ZN(n9771)
         );
  OAI211_X1 U10931 ( .C1(n9773), .C2(n9795), .A(n9772), .B(n9771), .ZN(
        P1_U3290) );
  AND2_X1 U10932 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9776), .ZN(P1_U3294) );
  AND2_X1 U10933 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9776), .ZN(P1_U3295) );
  AND2_X1 U10934 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9776), .ZN(P1_U3296) );
  AND2_X1 U10935 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9776), .ZN(P1_U3297) );
  AND2_X1 U10936 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9776), .ZN(P1_U3298) );
  AND2_X1 U10937 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9776), .ZN(P1_U3299) );
  AND2_X1 U10938 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9776), .ZN(P1_U3300) );
  AND2_X1 U10939 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9776), .ZN(P1_U3301) );
  AND2_X1 U10940 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9776), .ZN(P1_U3302) );
  AND2_X1 U10941 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9776), .ZN(P1_U3303) );
  AND2_X1 U10942 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9776), .ZN(P1_U3304) );
  AND2_X1 U10943 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9776), .ZN(P1_U3305) );
  AND2_X1 U10944 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9776), .ZN(P1_U3306) );
  AND2_X1 U10945 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9776), .ZN(P1_U3307) );
  AND2_X1 U10946 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9776), .ZN(P1_U3308) );
  AND2_X1 U10947 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9776), .ZN(P1_U3309) );
  AND2_X1 U10948 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9776), .ZN(P1_U3310) );
  AND2_X1 U10949 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9776), .ZN(P1_U3311) );
  AND2_X1 U10950 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9776), .ZN(P1_U3312) );
  AND2_X1 U10951 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9776), .ZN(P1_U3313) );
  AND2_X1 U10952 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9776), .ZN(P1_U3314) );
  AND2_X1 U10953 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9776), .ZN(P1_U3315) );
  AND2_X1 U10954 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9776), .ZN(P1_U3316) );
  AND2_X1 U10955 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9776), .ZN(P1_U3317) );
  AND2_X1 U10956 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9776), .ZN(P1_U3318) );
  AND2_X1 U10957 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9776), .ZN(P1_U3319) );
  INV_X1 U10958 ( .A(n9776), .ZN(n9780) );
  NOR2_X1 U10959 ( .A1(n9780), .A2(n10251), .ZN(P1_U3320) );
  NOR2_X1 U10960 ( .A1(n9780), .A2(n9777), .ZN(P1_U3321) );
  NOR2_X1 U10961 ( .A1(n9780), .A2(n9778), .ZN(P1_U3322) );
  NOR2_X1 U10962 ( .A1(n9780), .A2(n9779), .ZN(P1_U3323) );
  INV_X1 U10963 ( .A(n9781), .ZN(n9786) );
  OAI21_X1 U10964 ( .B1(n9783), .B2(n9848), .A(n9782), .ZN(n9785) );
  AOI211_X1 U10965 ( .C1(n9853), .C2(n9786), .A(n9785), .B(n9784), .ZN(n9859)
         );
  INV_X1 U10966 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9787) );
  AOI22_X1 U10967 ( .A1(n9858), .A2(n9859), .B1(n9787), .B2(n5809), .ZN(
        P1_U3456) );
  OAI21_X1 U10968 ( .B1(n9789), .B2(n9848), .A(n9788), .ZN(n9791) );
  AOI211_X1 U10969 ( .C1(n9845), .C2(n9792), .A(n9791), .B(n9790), .ZN(n9860)
         );
  INV_X1 U10970 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9793) );
  AOI22_X1 U10971 ( .A1(n9858), .A2(n9860), .B1(n9793), .B2(n5809), .ZN(
        P1_U3459) );
  OAI211_X1 U10972 ( .C1(n9796), .C2(n9848), .A(n9795), .B(n9794), .ZN(n9797)
         );
  AOI21_X1 U10973 ( .B1(n9845), .B2(n9798), .A(n9797), .ZN(n9861) );
  AOI22_X1 U10974 ( .A1(n9858), .A2(n9861), .B1(n5328), .B2(n5809), .ZN(
        P1_U3462) );
  AOI21_X1 U10975 ( .B1(n9801), .B2(n9800), .A(n9799), .ZN(n9802) );
  OAI211_X1 U10976 ( .C1(n9805), .C2(n9804), .A(n9803), .B(n9802), .ZN(n9806)
         );
  INV_X1 U10977 ( .A(n9806), .ZN(n9862) );
  INV_X1 U10978 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9807) );
  AOI22_X1 U10979 ( .A1(n9858), .A2(n9862), .B1(n9807), .B2(n5809), .ZN(
        P1_U3465) );
  OAI21_X1 U10980 ( .B1(n9809), .B2(n9848), .A(n9808), .ZN(n9812) );
  INV_X1 U10981 ( .A(n9810), .ZN(n9811) );
  AOI211_X1 U10982 ( .C1(n9845), .C2(n9813), .A(n9812), .B(n9811), .ZN(n9864)
         );
  INV_X1 U10983 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9814) );
  AOI22_X1 U10984 ( .A1(n9858), .A2(n9864), .B1(n9814), .B2(n5809), .ZN(
        P1_U3468) );
  AND2_X1 U10985 ( .A1(n9815), .A2(n9845), .ZN(n9819) );
  OAI21_X1 U10986 ( .B1(n9817), .B2(n9848), .A(n9816), .ZN(n9818) );
  NOR3_X1 U10987 ( .A1(n9820), .A2(n9819), .A3(n9818), .ZN(n9865) );
  INV_X1 U10988 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9821) );
  AOI22_X1 U10989 ( .A1(n9858), .A2(n9865), .B1(n9821), .B2(n5809), .ZN(
        P1_U3471) );
  OAI21_X1 U10990 ( .B1(n9823), .B2(n9848), .A(n9822), .ZN(n9825) );
  AOI211_X1 U10991 ( .C1(n9853), .C2(n9826), .A(n9825), .B(n9824), .ZN(n9867)
         );
  INV_X1 U10992 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9827) );
  AOI22_X1 U10993 ( .A1(n9858), .A2(n9867), .B1(n9827), .B2(n5809), .ZN(
        P1_U3474) );
  INV_X1 U10994 ( .A(n9828), .ZN(n9833) );
  OAI21_X1 U10995 ( .B1(n9830), .B2(n9848), .A(n9829), .ZN(n9832) );
  AOI211_X1 U10996 ( .C1(n9853), .C2(n9833), .A(n9832), .B(n9831), .ZN(n9869)
         );
  INV_X1 U10997 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9834) );
  AOI22_X1 U10998 ( .A1(n9858), .A2(n9869), .B1(n9834), .B2(n5809), .ZN(
        P1_U3477) );
  AND2_X1 U10999 ( .A1(n9835), .A2(n9845), .ZN(n9838) );
  OAI21_X1 U11000 ( .B1(n4851), .B2(n9848), .A(n9836), .ZN(n9837) );
  NOR3_X1 U11001 ( .A1(n9839), .A2(n9838), .A3(n9837), .ZN(n9870) );
  INV_X1 U11002 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9840) );
  AOI22_X1 U11003 ( .A1(n9858), .A2(n9870), .B1(n9840), .B2(n5809), .ZN(
        P1_U3480) );
  OAI211_X1 U11004 ( .C1(n9843), .C2(n9848), .A(n9842), .B(n9841), .ZN(n9844)
         );
  AOI21_X1 U11005 ( .B1(n9846), .B2(n9845), .A(n9844), .ZN(n9872) );
  INV_X1 U11006 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9847) );
  AOI22_X1 U11007 ( .A1(n9858), .A2(n9872), .B1(n9847), .B2(n5809), .ZN(
        P1_U3492) );
  OAI22_X1 U11008 ( .A1(n9851), .A2(n9850), .B1(n9849), .B2(n9848), .ZN(n9852)
         );
  AOI21_X1 U11009 ( .B1(n9854), .B2(n9853), .A(n9852), .ZN(n9855) );
  AND2_X1 U11010 ( .A1(n9856), .A2(n9855), .ZN(n9874) );
  INV_X1 U11011 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9857) );
  AOI22_X1 U11012 ( .A1(n9858), .A2(n9874), .B1(n9857), .B2(n5809), .ZN(
        P1_U3495) );
  AOI22_X1 U11013 ( .A1(n9875), .A2(n9859), .B1(n6755), .B2(n5819), .ZN(
        P1_U3523) );
  AOI22_X1 U11014 ( .A1(n9875), .A2(n9860), .B1(n6754), .B2(n5819), .ZN(
        P1_U3524) );
  AOI22_X1 U11015 ( .A1(n9875), .A2(n9861), .B1(n6758), .B2(n5819), .ZN(
        P1_U3525) );
  AOI22_X1 U11016 ( .A1(n9875), .A2(n9862), .B1(n6761), .B2(n5819), .ZN(
        P1_U3526) );
  AOI22_X1 U11017 ( .A1(n9875), .A2(n9864), .B1(n9863), .B2(n5819), .ZN(
        P1_U3527) );
  AOI22_X1 U11018 ( .A1(n9875), .A2(n9865), .B1(n6775), .B2(n5819), .ZN(
        P1_U3528) );
  AOI22_X1 U11019 ( .A1(n9875), .A2(n9867), .B1(n9866), .B2(n5819), .ZN(
        P1_U3529) );
  AOI22_X1 U11020 ( .A1(n9875), .A2(n9869), .B1(n9868), .B2(n5819), .ZN(
        P1_U3530) );
  AOI22_X1 U11021 ( .A1(n9875), .A2(n9870), .B1(n6897), .B2(n5819), .ZN(
        P1_U3531) );
  AOI22_X1 U11022 ( .A1(n9875), .A2(n9872), .B1(n9871), .B2(n5819), .ZN(
        P1_U3535) );
  AOI22_X1 U11023 ( .A1(n9875), .A2(n9874), .B1(n9873), .B2(n5819), .ZN(
        P1_U3536) );
  AOI22_X1 U11024 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n10007), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n9883) );
  NOR2_X1 U11025 ( .A1(n9876), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9877) );
  INV_X1 U11026 ( .A(n9900), .ZN(n9879) );
  OAI22_X1 U11027 ( .A1(n10016), .A2(n9881), .B1(n9880), .B2(n9879), .ZN(n9882) );
  OAI211_X1 U11028 ( .C1(n9885), .C2(n9884), .A(n9883), .B(n9882), .ZN(
        P2_U3182) );
  AND2_X1 U11029 ( .A1(n9887), .A2(n9886), .ZN(n9897) );
  NAND2_X1 U11030 ( .A1(n9889), .A2(n9888), .ZN(n9890) );
  NAND2_X1 U11031 ( .A1(n9891), .A2(n9890), .ZN(n9894) );
  INV_X1 U11032 ( .A(n9892), .ZN(n9893) );
  AOI22_X1 U11033 ( .A1(n10017), .A2(n9894), .B1(n9893), .B2(n10008), .ZN(
        n9896) );
  NAND2_X1 U11034 ( .A1(n10007), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n9895) );
  OAI211_X1 U11035 ( .C1(n9897), .C2(n10023), .A(n9896), .B(n9895), .ZN(n9898)
         );
  INV_X1 U11036 ( .A(n9898), .ZN(n9903) );
  XOR2_X1 U11037 ( .A(n9900), .B(n9899), .Z(n9901) );
  NAND2_X1 U11038 ( .A1(n9901), .A2(n10016), .ZN(n9902) );
  OAI211_X1 U11039 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n5847), .A(n9903), .B(
        n9902), .ZN(P2_U3183) );
  INV_X1 U11040 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10109) );
  OAI21_X1 U11041 ( .B1(n9906), .B2(n9905), .A(n9904), .ZN(n9907) );
  INV_X1 U11042 ( .A(n9907), .ZN(n9916) );
  OAI21_X1 U11043 ( .B1(n9910), .B2(n9909), .A(n9908), .ZN(n9911) );
  NAND2_X1 U11044 ( .A1(n10017), .A2(n9911), .ZN(n9915) );
  NOR2_X1 U11045 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7150), .ZN(n9912) );
  AOI21_X1 U11046 ( .B1(n10008), .B2(n9913), .A(n9912), .ZN(n9914) );
  OAI211_X1 U11047 ( .C1(n9916), .C2(n10023), .A(n9915), .B(n9914), .ZN(n9917)
         );
  INV_X1 U11048 ( .A(n9917), .ZN(n9922) );
  XOR2_X1 U11049 ( .A(n9919), .B(n9918), .Z(n9920) );
  NAND2_X1 U11050 ( .A1(n9920), .A2(n10016), .ZN(n9921) );
  OAI211_X1 U11051 ( .C1(n10109), .C2(n9941), .A(n9922), .B(n9921), .ZN(
        P2_U3184) );
  INV_X1 U11052 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10105) );
  OAI21_X1 U11053 ( .B1(n4592), .B2(P2_REG2_REG_3__SCAN_IN), .A(n9923), .ZN(
        n9924) );
  INV_X1 U11054 ( .A(n9924), .ZN(n9932) );
  XNOR2_X1 U11055 ( .A(n9926), .B(n9925), .ZN(n9927) );
  OR2_X1 U11056 ( .A1(n9928), .A2(n9927), .ZN(n9931) );
  AOI21_X1 U11057 ( .B1(n10008), .B2(n4962), .A(n9929), .ZN(n9930) );
  OAI211_X1 U11058 ( .C1(n10023), .C2(n9932), .A(n9931), .B(n9930), .ZN(n9933)
         );
  INV_X1 U11059 ( .A(n9933), .ZN(n9940) );
  AOI21_X1 U11060 ( .B1(n9936), .B2(n9935), .A(n9934), .ZN(n9938) );
  OR2_X1 U11061 ( .A1(n9938), .A2(n9937), .ZN(n9939) );
  OAI211_X1 U11062 ( .C1(n10105), .C2(n9941), .A(n9940), .B(n9939), .ZN(
        P2_U3185) );
  AOI22_X1 U11063 ( .A1(n9942), .A2(n10008), .B1(n10007), .B2(
        P2_ADDR_REG_13__SCAN_IN), .ZN(n9956) );
  OAI21_X1 U11064 ( .B1(n9945), .B2(n9944), .A(n9943), .ZN(n9949) );
  OAI21_X1 U11065 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n9947), .A(n9946), .ZN(
        n9948) );
  AOI22_X1 U11066 ( .A1(n9949), .A2(n10016), .B1(n10017), .B2(n9948), .ZN(
        n9955) );
  AOI21_X1 U11067 ( .B1(n9951), .B2(n8797), .A(n9950), .ZN(n9952) );
  OR2_X1 U11068 ( .A1(n10023), .A2(n9952), .ZN(n9953) );
  NAND4_X1 U11069 ( .A1(n9956), .A2(n9955), .A3(n9954), .A4(n9953), .ZN(
        P2_U3195) );
  AOI22_X1 U11070 ( .A1(n9957), .A2(n10008), .B1(n10007), .B2(
        P2_ADDR_REG_14__SCAN_IN), .ZN(n9973) );
  OAI21_X1 U11071 ( .B1(n9960), .B2(n9959), .A(n9958), .ZN(n9965) );
  OAI21_X1 U11072 ( .B1(n9963), .B2(n9962), .A(n9961), .ZN(n9964) );
  AOI22_X1 U11073 ( .A1(n9965), .A2(n10017), .B1(n10016), .B2(n9964), .ZN(
        n9972) );
  NAND2_X1 U11074 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3151), .ZN(n9971) );
  AOI21_X1 U11075 ( .B1(n9968), .B2(n9967), .A(n9966), .ZN(n9969) );
  OR2_X1 U11076 ( .A1(n9969), .A2(n10023), .ZN(n9970) );
  NAND4_X1 U11077 ( .A1(n9973), .A2(n9972), .A3(n9971), .A4(n9970), .ZN(
        P2_U3196) );
  AOI22_X1 U11078 ( .A1(n9974), .A2(n10008), .B1(n10007), .B2(
        P2_ADDR_REG_15__SCAN_IN), .ZN(n9989) );
  OAI21_X1 U11079 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n9976), .A(n9975), .ZN(
        n9981) );
  OAI21_X1 U11080 ( .B1(n9979), .B2(n9978), .A(n9977), .ZN(n9980) );
  AOI22_X1 U11081 ( .A1(n9981), .A2(n10017), .B1(n10016), .B2(n9980), .ZN(
        n9988) );
  AOI21_X1 U11082 ( .B1(n9984), .B2(n9983), .A(n9982), .ZN(n9985) );
  OR2_X1 U11083 ( .A1(n10023), .A2(n9985), .ZN(n9986) );
  NAND4_X1 U11084 ( .A1(n9989), .A2(n9988), .A3(n9987), .A4(n9986), .ZN(
        P2_U3197) );
  AOI22_X1 U11085 ( .A1(n9990), .A2(n10008), .B1(n10007), .B2(
        P2_ADDR_REG_16__SCAN_IN), .ZN(n10006) );
  OAI21_X1 U11086 ( .B1(n9993), .B2(n9992), .A(n9991), .ZN(n9998) );
  OAI21_X1 U11087 ( .B1(n9996), .B2(n9995), .A(n9994), .ZN(n9997) );
  AOI22_X1 U11088 ( .A1(n9998), .A2(n10017), .B1(n10016), .B2(n9997), .ZN(
        n10005) );
  AOI21_X1 U11089 ( .B1(n10001), .B2(n10000), .A(n9999), .ZN(n10002) );
  OR2_X1 U11090 ( .A1(n10002), .A2(n10023), .ZN(n10003) );
  NAND4_X1 U11091 ( .A1(n10006), .A2(n10005), .A3(n10004), .A4(n10003), .ZN(
        P2_U3198) );
  AOI22_X1 U11092 ( .A1(n10009), .A2(n10008), .B1(n10007), .B2(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n10027) );
  OAI21_X1 U11093 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n10011), .A(n10010), 
        .ZN(n10018) );
  OAI21_X1 U11094 ( .B1(n10014), .B2(n10013), .A(n10012), .ZN(n10015) );
  AOI22_X1 U11095 ( .A1(n10018), .A2(n10017), .B1(n10016), .B2(n10015), .ZN(
        n10026) );
  NAND2_X1 U11096 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3151), .ZN(n10025)
         );
  AOI21_X1 U11097 ( .B1(n10021), .B2(n10020), .A(n10019), .ZN(n10022) );
  OR2_X1 U11098 ( .A1(n10023), .A2(n10022), .ZN(n10024) );
  NAND4_X1 U11099 ( .A1(n10027), .A2(n10026), .A3(n10025), .A4(n10024), .ZN(
        P2_U3199) );
  NOR2_X1 U11100 ( .A1(n10028), .A2(n10078), .ZN(n10030) );
  AOI211_X1 U11101 ( .C1(n10076), .C2(n10031), .A(n10030), .B(n10029), .ZN(
        n10087) );
  AOI22_X1 U11102 ( .A1(n10086), .A2(n5873), .B1(n10087), .B2(n10084), .ZN(
        P2_U3396) );
  INV_X1 U11103 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10037) );
  NAND2_X1 U11104 ( .A1(n10032), .A2(n10083), .ZN(n10036) );
  NAND2_X1 U11105 ( .A1(n10033), .A2(n10063), .ZN(n10034) );
  AND3_X1 U11106 ( .A1(n10036), .A2(n10035), .A3(n10034), .ZN(n10088) );
  AOI22_X1 U11107 ( .A1(n10086), .A2(n10037), .B1(n10088), .B2(n10084), .ZN(
        P2_U3399) );
  NAND2_X1 U11108 ( .A1(n10038), .A2(n10083), .ZN(n10041) );
  NAND2_X1 U11109 ( .A1(n10039), .A2(n10063), .ZN(n10040) );
  AND3_X1 U11110 ( .A1(n10042), .A2(n10041), .A3(n10040), .ZN(n10089) );
  AOI22_X1 U11111 ( .A1(n10086), .A2(n5899), .B1(n10089), .B2(n10084), .ZN(
        P2_U3402) );
  OAI21_X1 U11112 ( .B1(n10044), .B2(n10078), .A(n10043), .ZN(n10045) );
  AOI21_X1 U11113 ( .B1(n10083), .B2(n10046), .A(n10045), .ZN(n10091) );
  AOI22_X1 U11114 ( .A1(n10086), .A2(n5915), .B1(n10091), .B2(n10084), .ZN(
        P2_U3405) );
  AND2_X1 U11115 ( .A1(n10047), .A2(n10063), .ZN(n10048) );
  NOR2_X1 U11116 ( .A1(n10049), .A2(n10048), .ZN(n10052) );
  NAND2_X1 U11117 ( .A1(n10050), .A2(n10083), .ZN(n10051) );
  AOI22_X1 U11118 ( .A1(n10086), .A2(n5928), .B1(n10092), .B2(n10084), .ZN(
        P2_U3408) );
  NOR2_X1 U11119 ( .A1(n10053), .A2(n10078), .ZN(n10055) );
  AOI211_X1 U11120 ( .C1(n10076), .C2(n10056), .A(n10055), .B(n10054), .ZN(
        n10093) );
  AOI22_X1 U11121 ( .A1(n10086), .A2(n5942), .B1(n10093), .B2(n10084), .ZN(
        P2_U3411) );
  INV_X1 U11122 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10064) );
  INV_X1 U11123 ( .A(n10057), .ZN(n10062) );
  NOR2_X1 U11124 ( .A1(n10059), .A2(n10058), .ZN(n10060) );
  AOI211_X1 U11125 ( .C1(n10063), .C2(n10062), .A(n10061), .B(n10060), .ZN(
        n10094) );
  AOI22_X1 U11126 ( .A1(n10086), .A2(n10064), .B1(n10094), .B2(n10084), .ZN(
        P2_U3414) );
  INV_X1 U11127 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10070) );
  INV_X1 U11128 ( .A(n10065), .ZN(n10066) );
  NOR2_X1 U11129 ( .A1(n10066), .A2(n10078), .ZN(n10068) );
  AOI211_X1 U11130 ( .C1(n10069), .C2(n10076), .A(n10068), .B(n10067), .ZN(
        n10096) );
  AOI22_X1 U11131 ( .A1(n10086), .A2(n10070), .B1(n10096), .B2(n10084), .ZN(
        P2_U3417) );
  INV_X1 U11132 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10077) );
  INV_X1 U11133 ( .A(n10071), .ZN(n10072) );
  NOR2_X1 U11134 ( .A1(n10072), .A2(n10078), .ZN(n10074) );
  AOI211_X1 U11135 ( .C1(n10076), .C2(n10075), .A(n10074), .B(n10073), .ZN(
        n10097) );
  AOI22_X1 U11136 ( .A1(n10086), .A2(n10077), .B1(n10097), .B2(n10084), .ZN(
        P2_U3420) );
  INV_X1 U11137 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10085) );
  NOR2_X1 U11138 ( .A1(n10079), .A2(n10078), .ZN(n10081) );
  AOI211_X1 U11139 ( .C1(n10083), .C2(n10082), .A(n10081), .B(n10080), .ZN(
        n10100) );
  AOI22_X1 U11140 ( .A1(n10086), .A2(n10085), .B1(n10100), .B2(n10084), .ZN(
        P2_U3423) );
  AOI22_X1 U11141 ( .A1(n10101), .A2(n10087), .B1(n6945), .B2(n10098), .ZN(
        P2_U3461) );
  AOI22_X1 U11142 ( .A1(n10101), .A2(n10088), .B1(n9925), .B2(n10098), .ZN(
        P2_U3462) );
  AOI22_X1 U11143 ( .A1(n10101), .A2(n10089), .B1(n6944), .B2(n10098), .ZN(
        P2_U3463) );
  INV_X1 U11144 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10090) );
  AOI22_X1 U11145 ( .A1(n10101), .A2(n10091), .B1(n10090), .B2(n10098), .ZN(
        P2_U3464) );
  AOI22_X1 U11146 ( .A1(n10101), .A2(n10092), .B1(n7180), .B2(n10098), .ZN(
        P2_U3465) );
  AOI22_X1 U11147 ( .A1(n10101), .A2(n10093), .B1(n7507), .B2(n10098), .ZN(
        P2_U3466) );
  AOI22_X1 U11148 ( .A1(n10101), .A2(n10094), .B1(n5953), .B2(n10098), .ZN(
        P2_U3467) );
  INV_X1 U11149 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10095) );
  AOI22_X1 U11150 ( .A1(n10101), .A2(n10096), .B1(n10095), .B2(n10098), .ZN(
        P2_U3468) );
  AOI22_X1 U11151 ( .A1(n10101), .A2(n10097), .B1(n5985), .B2(n10098), .ZN(
        P2_U3469) );
  INV_X1 U11152 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10099) );
  AOI22_X1 U11153 ( .A1(n10101), .A2(n10100), .B1(n10099), .B2(n10098), .ZN(
        P2_U3470) );
  AOI21_X1 U11154 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10108) );
  NAND2_X1 U11155 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n10102) );
  NOR2_X1 U11156 ( .A1(n10103), .A2(n10102), .ZN(n10106) );
  NOR2_X1 U11157 ( .A1(n10108), .A2(n10106), .ZN(n10104) );
  XOR2_X1 U11158 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10104), .Z(ADD_1068_U5) );
  XOR2_X1 U11159 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11160 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10153) );
  NOR2_X1 U11161 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10151) );
  NOR2_X1 U11162 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10149) );
  NOR2_X1 U11163 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10147) );
  NOR2_X1 U11164 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10145) );
  NOR2_X1 U11165 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10143) );
  NOR2_X1 U11166 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10139) );
  NOR2_X1 U11167 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10135) );
  NOR2_X1 U11168 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10131) );
  NOR2_X1 U11169 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10127) );
  NOR2_X1 U11170 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10123) );
  NOR2_X1 U11171 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n10120) );
  NOR2_X1 U11172 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10117) );
  NOR2_X1 U11173 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10115) );
  NAND2_X1 U11174 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10113) );
  XNOR2_X1 U11175 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n10105), .ZN(n10560) );
  NAND2_X1 U11176 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10111) );
  NOR2_X1 U11177 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10106), .ZN(n10107) );
  NOR2_X1 U11178 ( .A1(n10108), .A2(n10107), .ZN(n10550) );
  XNOR2_X1 U11179 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n10109), .ZN(n10549) );
  NAND2_X1 U11180 ( .A1(n10550), .A2(n10549), .ZN(n10110) );
  NAND2_X1 U11181 ( .A1(n10111), .A2(n10110), .ZN(n10559) );
  NAND2_X1 U11182 ( .A1(n10560), .A2(n10559), .ZN(n10112) );
  NAND2_X1 U11183 ( .A1(n10113), .A2(n10112), .ZN(n10562) );
  XNOR2_X1 U11184 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10561) );
  NOR2_X1 U11185 ( .A1(n10562), .A2(n10561), .ZN(n10114) );
  NOR2_X1 U11186 ( .A1(n10115), .A2(n10114), .ZN(n10552) );
  XNOR2_X1 U11187 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10551) );
  NOR2_X1 U11188 ( .A1(n10552), .A2(n10551), .ZN(n10116) );
  NOR2_X1 U11189 ( .A1(n10117), .A2(n10116), .ZN(n10558) );
  XOR2_X1 U11190 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n10118), .Z(n10557) );
  NOR2_X1 U11191 ( .A1(n10558), .A2(n10557), .ZN(n10119) );
  NOR2_X1 U11192 ( .A1(n10120), .A2(n10119), .ZN(n10554) );
  INV_X1 U11193 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10121) );
  XOR2_X1 U11194 ( .A(n10121), .B(P1_ADDR_REG_7__SCAN_IN), .Z(n10553) );
  NOR2_X1 U11195 ( .A1(n10554), .A2(n10553), .ZN(n10122) );
  NOR2_X1 U11196 ( .A1(n10123), .A2(n10122), .ZN(n10556) );
  INV_X1 U11197 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10125) );
  AOI22_X1 U11198 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10125), .B1(
        P1_ADDR_REG_8__SCAN_IN), .B2(n10124), .ZN(n10555) );
  NOR2_X1 U11199 ( .A1(n10556), .A2(n10555), .ZN(n10126) );
  NOR2_X1 U11200 ( .A1(n10127), .A2(n10126), .ZN(n10548) );
  INV_X1 U11201 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10129) );
  AOI22_X1 U11202 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10129), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n10128), .ZN(n10547) );
  NOR2_X1 U11203 ( .A1(n10548), .A2(n10547), .ZN(n10130) );
  NOR2_X1 U11204 ( .A1(n10131), .A2(n10130), .ZN(n10171) );
  INV_X1 U11205 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10133) );
  AOI22_X1 U11206 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n10133), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n10132), .ZN(n10170) );
  NOR2_X1 U11207 ( .A1(n10171), .A2(n10170), .ZN(n10134) );
  NOR2_X1 U11208 ( .A1(n10135), .A2(n10134), .ZN(n10169) );
  INV_X1 U11209 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10137) );
  AOI22_X1 U11210 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n10137), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n10136), .ZN(n10168) );
  NOR2_X1 U11211 ( .A1(n10169), .A2(n10168), .ZN(n10138) );
  NOR2_X1 U11212 ( .A1(n10139), .A2(n10138), .ZN(n10167) );
  INV_X1 U11213 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10141) );
  AOI22_X1 U11214 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n10141), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n10140), .ZN(n10166) );
  NOR2_X1 U11215 ( .A1(n10167), .A2(n10166), .ZN(n10142) );
  NOR2_X1 U11216 ( .A1(n10143), .A2(n10142), .ZN(n10165) );
  XNOR2_X1 U11217 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10164) );
  NOR2_X1 U11218 ( .A1(n10165), .A2(n10164), .ZN(n10144) );
  NOR2_X1 U11219 ( .A1(n10145), .A2(n10144), .ZN(n10163) );
  XNOR2_X1 U11220 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10162) );
  NOR2_X1 U11221 ( .A1(n10163), .A2(n10162), .ZN(n10146) );
  NOR2_X1 U11222 ( .A1(n10147), .A2(n10146), .ZN(n10161) );
  XNOR2_X1 U11223 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10160) );
  NOR2_X1 U11224 ( .A1(n10161), .A2(n10160), .ZN(n10148) );
  NOR2_X1 U11225 ( .A1(n10149), .A2(n10148), .ZN(n10159) );
  XNOR2_X1 U11226 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10158) );
  NOR2_X1 U11227 ( .A1(n10159), .A2(n10158), .ZN(n10150) );
  NOR2_X1 U11228 ( .A1(n10151), .A2(n10150), .ZN(n10157) );
  XNOR2_X1 U11229 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10156) );
  NOR2_X1 U11230 ( .A1(n10157), .A2(n10156), .ZN(n10152) );
  NOR2_X1 U11231 ( .A1(n10153), .A2(n10152), .ZN(n10154) );
  NOR2_X1 U11232 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10154), .ZN(n10174) );
  AND2_X1 U11233 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10154), .ZN(n10172) );
  NOR2_X1 U11234 ( .A1(n10174), .A2(n10172), .ZN(n10155) );
  XOR2_X1 U11235 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n10155), .Z(ADD_1068_U55)
         );
  XNOR2_X1 U11236 ( .A(n10157), .B(n10156), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11237 ( .A(n10159), .B(n10158), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11238 ( .A(n10161), .B(n10160), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11239 ( .A(n10163), .B(n10162), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11240 ( .A(n10165), .B(n10164), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11241 ( .A(n10167), .B(n10166), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11242 ( .A(n10169), .B(n10168), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11243 ( .A(n10171), .B(n10170), .ZN(ADD_1068_U63) );
  NOR2_X1 U11244 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10172), .ZN(n10173) );
  NOR2_X1 U11245 ( .A1(n10174), .A2(n10173), .ZN(n10546) );
  XOR2_X1 U11246 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_g37), .Z(n10181)
         );
  AOI22_X1 U11247 ( .A1(SI_1_), .A2(keyinput_g31), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_g79), .ZN(n10175) );
  OAI221_X1 U11248 ( .B1(SI_1_), .B2(keyinput_g31), .C1(
        P2_DATAO_REG_17__SCAN_IN), .C2(keyinput_g79), .A(n10175), .ZN(n10180)
         );
  AOI22_X1 U11249 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_g61), .B1(
        P1_IR_REG_27__SCAN_IN), .B2(keyinput_g117), .ZN(n10176) );
  OAI221_X1 U11250 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .C1(
        P1_IR_REG_27__SCAN_IN), .C2(keyinput_g117), .A(n10176), .ZN(n10179) );
  AOI22_X1 U11251 ( .A1(SI_28_), .A2(keyinput_g4), .B1(P1_D_REG_4__SCAN_IN), 
        .B2(keyinput_g126), .ZN(n10177) );
  OAI221_X1 U11252 ( .B1(SI_28_), .B2(keyinput_g4), .C1(P1_D_REG_4__SCAN_IN), 
        .C2(keyinput_g126), .A(n10177), .ZN(n10178) );
  NOR4_X1 U11253 ( .A1(n10181), .A2(n10180), .A3(n10179), .A4(n10178), .ZN(
        n10209) );
  AOI22_X1 U11254 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_g0), .B1(
        P1_D_REG_2__SCAN_IN), .B2(keyinput_g124), .ZN(n10182) );
  OAI221_X1 U11255 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_g0), .C1(
        P1_D_REG_2__SCAN_IN), .C2(keyinput_g124), .A(n10182), .ZN(n10189) );
  AOI22_X1 U11256 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(keyinput_g113), .B1(
        P1_IR_REG_3__SCAN_IN), .B2(keyinput_g93), .ZN(n10183) );
  OAI221_X1 U11257 ( .B1(P1_IR_REG_23__SCAN_IN), .B2(keyinput_g113), .C1(
        P1_IR_REG_3__SCAN_IN), .C2(keyinput_g93), .A(n10183), .ZN(n10188) );
  AOI22_X1 U11258 ( .A1(SI_29_), .A2(keyinput_g3), .B1(SI_3_), .B2(
        keyinput_g29), .ZN(n10184) );
  OAI221_X1 U11259 ( .B1(SI_29_), .B2(keyinput_g3), .C1(SI_3_), .C2(
        keyinput_g29), .A(n10184), .ZN(n10187) );
  AOI22_X1 U11260 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_g63), .B1(SI_6_), .B2(keyinput_g26), .ZN(n10185) );
  OAI221_X1 U11261 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .C1(
        SI_6_), .C2(keyinput_g26), .A(n10185), .ZN(n10186) );
  NOR4_X1 U11262 ( .A1(n10189), .A2(n10188), .A3(n10187), .A4(n10186), .ZN(
        n10208) );
  AOI22_X1 U11263 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput_g87), .B1(
        SI_14_), .B2(keyinput_g18), .ZN(n10190) );
  OAI221_X1 U11264 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_g87), .C1(
        SI_14_), .C2(keyinput_g18), .A(n10190), .ZN(n10197) );
  AOI22_X1 U11265 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(
        P2_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .ZN(n10191) );
  OAI221_X1 U11266 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_g42), .A(n10191), .ZN(n10196)
         );
  AOI22_X1 U11267 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(keyinput_g84), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(keyinput_g77), .ZN(n10192) );
  OAI221_X1 U11268 ( .B1(P2_DATAO_REG_12__SCAN_IN), .B2(keyinput_g84), .C1(
        P2_DATAO_REG_19__SCAN_IN), .C2(keyinput_g77), .A(n10192), .ZN(n10195)
         );
  AOI22_X1 U11269 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(keyinput_g76), .B1(
        P1_IR_REG_7__SCAN_IN), .B2(keyinput_g97), .ZN(n10193) );
  OAI221_X1 U11270 ( .B1(P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_g76), .C1(
        P1_IR_REG_7__SCAN_IN), .C2(keyinput_g97), .A(n10193), .ZN(n10194) );
  NOR4_X1 U11271 ( .A1(n10197), .A2(n10196), .A3(n10195), .A4(n10194), .ZN(
        n10207) );
  AOI22_X1 U11272 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_g39), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(keyinput_g82), .ZN(n10198) );
  OAI221_X1 U11273 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .C1(
        P2_DATAO_REG_14__SCAN_IN), .C2(keyinput_g82), .A(n10198), .ZN(n10205)
         );
  AOI22_X1 U11274 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(keyinput_g68), .B1(
        P1_IR_REG_20__SCAN_IN), .B2(keyinput_g110), .ZN(n10199) );
  OAI221_X1 U11275 ( .B1(P2_DATAO_REG_28__SCAN_IN), .B2(keyinput_g68), .C1(
        P1_IR_REG_20__SCAN_IN), .C2(keyinput_g110), .A(n10199), .ZN(n10204) );
  AOI22_X1 U11276 ( .A1(SI_13_), .A2(keyinput_g19), .B1(SI_16_), .B2(
        keyinput_g16), .ZN(n10200) );
  OAI221_X1 U11277 ( .B1(SI_13_), .B2(keyinput_g19), .C1(SI_16_), .C2(
        keyinput_g16), .A(n10200), .ZN(n10203) );
  AOI22_X1 U11278 ( .A1(SI_12_), .A2(keyinput_g20), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(keyinput_g71), .ZN(n10201) );
  OAI221_X1 U11279 ( .B1(SI_12_), .B2(keyinput_g20), .C1(
        P2_DATAO_REG_25__SCAN_IN), .C2(keyinput_g71), .A(n10201), .ZN(n10202)
         );
  NOR4_X1 U11280 ( .A1(n10205), .A2(n10204), .A3(n10203), .A4(n10202), .ZN(
        n10206) );
  NAND4_X1 U11281 ( .A1(n10209), .A2(n10208), .A3(n10207), .A4(n10206), .ZN(
        n10355) );
  AOI22_X1 U11282 ( .A1(P1_D_REG_0__SCAN_IN), .A2(keyinput_g122), .B1(
        P1_IR_REG_22__SCAN_IN), .B2(keyinput_g112), .ZN(n10210) );
  OAI221_X1 U11283 ( .B1(P1_D_REG_0__SCAN_IN), .B2(keyinput_g122), .C1(
        P1_IR_REG_22__SCAN_IN), .C2(keyinput_g112), .A(n10210), .ZN(n10217) );
  AOI22_X1 U11284 ( .A1(SI_9_), .A2(keyinput_g23), .B1(SI_15_), .B2(
        keyinput_g17), .ZN(n10211) );
  OAI221_X1 U11285 ( .B1(SI_9_), .B2(keyinput_g23), .C1(SI_15_), .C2(
        keyinput_g17), .A(n10211), .ZN(n10216) );
  AOI22_X1 U11286 ( .A1(SI_17_), .A2(keyinput_g15), .B1(SI_27_), .B2(
        keyinput_g5), .ZN(n10212) );
  OAI221_X1 U11287 ( .B1(SI_17_), .B2(keyinput_g15), .C1(SI_27_), .C2(
        keyinput_g5), .A(n10212), .ZN(n10215) );
  AOI22_X1 U11288 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_g50), .B1(
        P1_IR_REG_11__SCAN_IN), .B2(keyinput_g101), .ZN(n10213) );
  OAI221_X1 U11289 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .C1(
        P1_IR_REG_11__SCAN_IN), .C2(keyinput_g101), .A(n10213), .ZN(n10214) );
  NOR4_X1 U11290 ( .A1(n10217), .A2(n10216), .A3(n10215), .A4(n10214), .ZN(
        n10249) );
  AOI22_X1 U11291 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_g36), .B1(SI_4_), .B2(keyinput_g28), .ZN(n10218) );
  OAI221_X1 U11292 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .C1(
        SI_4_), .C2(keyinput_g28), .A(n10218), .ZN(n10225) );
  AOI22_X1 U11293 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(keyinput_g78), .B1(
        P1_D_REG_1__SCAN_IN), .B2(keyinput_g123), .ZN(n10219) );
  OAI221_X1 U11294 ( .B1(P2_DATAO_REG_18__SCAN_IN), .B2(keyinput_g78), .C1(
        P1_D_REG_1__SCAN_IN), .C2(keyinput_g123), .A(n10219), .ZN(n10224) );
  AOI22_X1 U11295 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_g43), .B1(SI_18_), .B2(keyinput_g14), .ZN(n10220) );
  OAI221_X1 U11296 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_g43), .C1(
        SI_18_), .C2(keyinput_g14), .A(n10220), .ZN(n10223) );
  AOI22_X1 U11297 ( .A1(SI_8_), .A2(keyinput_g24), .B1(P1_D_REG_3__SCAN_IN), 
        .B2(keyinput_g125), .ZN(n10221) );
  OAI221_X1 U11298 ( .B1(SI_8_), .B2(keyinput_g24), .C1(P1_D_REG_3__SCAN_IN), 
        .C2(keyinput_g125), .A(n10221), .ZN(n10222) );
  NOR4_X1 U11299 ( .A1(n10225), .A2(n10224), .A3(n10223), .A4(n10222), .ZN(
        n10248) );
  AOI22_X1 U11300 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_g44), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(keyinput_g81), .ZN(n10226) );
  OAI221_X1 U11301 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .C1(
        P2_DATAO_REG_15__SCAN_IN), .C2(keyinput_g81), .A(n10226), .ZN(n10233)
         );
  AOI22_X1 U11302 ( .A1(SI_10_), .A2(keyinput_g22), .B1(P1_IR_REG_14__SCAN_IN), 
        .B2(keyinput_g104), .ZN(n10227) );
  OAI221_X1 U11303 ( .B1(SI_10_), .B2(keyinput_g22), .C1(P1_IR_REG_14__SCAN_IN), .C2(keyinput_g104), .A(n10227), .ZN(n10232) );
  AOI22_X1 U11304 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_g57), .B1(
        P2_B_REG_SCAN_IN), .B2(keyinput_g64), .ZN(n10228) );
  OAI221_X1 U11305 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .C1(
        P2_B_REG_SCAN_IN), .C2(keyinput_g64), .A(n10228), .ZN(n10231) );
  AOI22_X1 U11306 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(keyinput_g72), .B1(
        P1_IR_REG_8__SCAN_IN), .B2(keyinput_g98), .ZN(n10229) );
  OAI221_X1 U11307 ( .B1(P2_DATAO_REG_24__SCAN_IN), .B2(keyinput_g72), .C1(
        P1_IR_REG_8__SCAN_IN), .C2(keyinput_g98), .A(n10229), .ZN(n10230) );
  NOR4_X1 U11308 ( .A1(n10233), .A2(n10232), .A3(n10231), .A4(n10230), .ZN(
        n10247) );
  AOI22_X1 U11309 ( .A1(n10236), .A2(keyinput_g86), .B1(n10235), .B2(
        keyinput_g106), .ZN(n10234) );
  OAI221_X1 U11310 ( .B1(n10236), .B2(keyinput_g86), .C1(n10235), .C2(
        keyinput_g106), .A(n10234), .ZN(n10245) );
  AOI22_X1 U11311 ( .A1(n10493), .A2(keyinput_g100), .B1(keyinput_g56), .B2(
        n10509), .ZN(n10237) );
  OAI221_X1 U11312 ( .B1(n10493), .B2(keyinput_g100), .C1(n10509), .C2(
        keyinput_g56), .A(n10237), .ZN(n10244) );
  AOI22_X1 U11313 ( .A1(n10450), .A2(keyinput_g60), .B1(n10239), .B2(
        keyinput_g6), .ZN(n10238) );
  OAI221_X1 U11314 ( .B1(n10450), .B2(keyinput_g60), .C1(n10239), .C2(
        keyinput_g6), .A(n10238), .ZN(n10243) );
  XOR2_X1 U11315 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_g52), .Z(n10241) );
  XNOR2_X1 U11316 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_g103), .ZN(n10240)
         );
  NAND2_X1 U11317 ( .A1(n10241), .A2(n10240), .ZN(n10242) );
  NOR4_X1 U11318 ( .A1(n10245), .A2(n10244), .A3(n10243), .A4(n10242), .ZN(
        n10246) );
  NAND4_X1 U11319 ( .A1(n10249), .A2(n10248), .A3(n10247), .A4(n10246), .ZN(
        n10354) );
  INV_X1 U11320 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10439) );
  AOI22_X1 U11321 ( .A1(n10439), .A2(keyinput_g55), .B1(n10251), .B2(
        keyinput_g127), .ZN(n10250) );
  OAI221_X1 U11322 ( .B1(n10439), .B2(keyinput_g55), .C1(n10251), .C2(
        keyinput_g127), .A(n10250), .ZN(n10262) );
  AOI22_X1 U11323 ( .A1(n10254), .A2(keyinput_g58), .B1(n10253), .B2(
        keyinput_g13), .ZN(n10252) );
  OAI221_X1 U11324 ( .B1(n10254), .B2(keyinput_g58), .C1(n10253), .C2(
        keyinput_g13), .A(n10252), .ZN(n10261) );
  AOI22_X1 U11325 ( .A1(n10256), .A2(keyinput_g40), .B1(n10440), .B2(
        keyinput_g88), .ZN(n10255) );
  OAI221_X1 U11326 ( .B1(n10256), .B2(keyinput_g40), .C1(n10440), .C2(
        keyinput_g88), .A(n10255), .ZN(n10260) );
  INV_X1 U11327 ( .A(SI_21_), .ZN(n10459) );
  XOR2_X1 U11328 ( .A(n10459), .B(keyinput_g11), .Z(n10258) );
  XNOR2_X1 U11329 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_g91), .ZN(n10257) );
  NAND2_X1 U11330 ( .A1(n10258), .A2(n10257), .ZN(n10259) );
  NOR4_X1 U11331 ( .A1(n10262), .A2(n10261), .A3(n10260), .A4(n10259), .ZN(
        n10304) );
  AOI22_X1 U11332 ( .A1(P2_U3151), .A2(keyinput_g34), .B1(keyinput_g67), .B2(
        n10476), .ZN(n10263) );
  OAI221_X1 U11333 ( .B1(P2_U3151), .B2(keyinput_g34), .C1(n10476), .C2(
        keyinput_g67), .A(n10263), .ZN(n10273) );
  INV_X1 U11334 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10266) );
  AOI22_X1 U11335 ( .A1(n10266), .A2(keyinput_g51), .B1(n10517), .B2(
        keyinput_g10), .ZN(n10265) );
  OAI221_X1 U11336 ( .B1(n10266), .B2(keyinput_g51), .C1(n10517), .C2(
        keyinput_g10), .A(n10265), .ZN(n10272) );
  XOR2_X1 U11337 ( .A(n5912), .B(keyinput_g49), .Z(n10270) );
  XNOR2_X1 U11338 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_g111), .ZN(n10269)
         );
  XNOR2_X1 U11339 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_g121), .ZN(n10268)
         );
  XNOR2_X1 U11340 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_g115), .ZN(n10267)
         );
  NAND4_X1 U11341 ( .A1(n10270), .A2(n10269), .A3(n10268), .A4(n10267), .ZN(
        n10271) );
  NOR3_X1 U11342 ( .A1(n10273), .A2(n10272), .A3(n10271), .ZN(n10303) );
  AOI22_X1 U11343 ( .A1(n10276), .A2(keyinput_g1), .B1(n10275), .B2(
        keyinput_g83), .ZN(n10274) );
  OAI221_X1 U11344 ( .B1(n10276), .B2(keyinput_g1), .C1(n10275), .C2(
        keyinput_g83), .A(n10274), .ZN(n10286) );
  AOI22_X1 U11345 ( .A1(n10488), .A2(keyinput_g62), .B1(n10278), .B2(
        keyinput_g73), .ZN(n10277) );
  OAI221_X1 U11346 ( .B1(n10488), .B2(keyinput_g62), .C1(n10278), .C2(
        keyinput_g73), .A(n10277), .ZN(n10285) );
  XOR2_X1 U11347 ( .A(n10279), .B(keyinput_g35), .Z(n10283) );
  XNOR2_X1 U11348 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_g75), .ZN(n10282) );
  XNOR2_X1 U11349 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_g94), .ZN(n10281) );
  XNOR2_X1 U11350 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_g114), .ZN(n10280)
         );
  NAND4_X1 U11351 ( .A1(n10283), .A2(n10282), .A3(n10281), .A4(n10280), .ZN(
        n10284) );
  NOR3_X1 U11352 ( .A1(n10286), .A2(n10285), .A3(n10284), .ZN(n10302) );
  INV_X1 U11353 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U11354 ( .A1(n10289), .A2(keyinput_g38), .B1(n10288), .B2(
        keyinput_g12), .ZN(n10287) );
  OAI221_X1 U11355 ( .B1(n10289), .B2(keyinput_g38), .C1(n10288), .C2(
        keyinput_g12), .A(n10287), .ZN(n10300) );
  AOI22_X1 U11356 ( .A1(n10292), .A2(keyinput_g80), .B1(n10291), .B2(
        keyinput_g7), .ZN(n10290) );
  OAI221_X1 U11357 ( .B1(n10292), .B2(keyinput_g80), .C1(n10291), .C2(
        keyinput_g7), .A(n10290), .ZN(n10299) );
  INV_X1 U11358 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10293) );
  XOR2_X1 U11359 ( .A(n10293), .B(keyinput_g47), .Z(n10297) );
  XNOR2_X1 U11360 ( .A(SI_2_), .B(keyinput_g30), .ZN(n10296) );
  XNOR2_X1 U11361 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_g54), .ZN(n10295)
         );
  XNOR2_X1 U11362 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_g108), .ZN(n10294)
         );
  NAND4_X1 U11363 ( .A1(n10297), .A2(n10296), .A3(n10295), .A4(n10294), .ZN(
        n10298) );
  NOR3_X1 U11364 ( .A1(n10300), .A2(n10299), .A3(n10298), .ZN(n10301) );
  NAND4_X1 U11365 ( .A1(n10304), .A2(n10303), .A3(n10302), .A4(n10301), .ZN(
        n10353) );
  AOI22_X1 U11366 ( .A1(n10306), .A2(keyinput_g96), .B1(keyinput_g45), .B2(
        n10491), .ZN(n10305) );
  OAI221_X1 U11367 ( .B1(n10306), .B2(keyinput_g96), .C1(n10491), .C2(
        keyinput_g45), .A(n10305), .ZN(n10315) );
  XOR2_X1 U11368 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_g107), .Z(n10314) );
  XNOR2_X1 U11369 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_g109), .ZN(n10310)
         );
  XNOR2_X1 U11370 ( .A(SI_24_), .B(keyinput_g8), .ZN(n10309) );
  XNOR2_X1 U11371 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_g48), .ZN(n10308)
         );
  XNOR2_X1 U11372 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_g99), .ZN(n10307) );
  NAND4_X1 U11373 ( .A1(n10310), .A2(n10309), .A3(n10308), .A4(n10307), .ZN(
        n10313) );
  INV_X1 U11374 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10311) );
  XNOR2_X1 U11375 ( .A(keyinput_g41), .B(n10311), .ZN(n10312) );
  NOR4_X1 U11376 ( .A1(n10315), .A2(n10314), .A3(n10313), .A4(n10312), .ZN(
        n10351) );
  AOI22_X1 U11377 ( .A1(n10317), .A2(keyinput_g69), .B1(keyinput_g25), .B2(
        n10449), .ZN(n10316) );
  OAI221_X1 U11378 ( .B1(n10317), .B2(keyinput_g69), .C1(n10449), .C2(
        keyinput_g25), .A(n10316), .ZN(n10325) );
  AOI22_X1 U11379 ( .A1(n10446), .A2(keyinput_g74), .B1(n10406), .B2(
        keyinput_g105), .ZN(n10318) );
  OAI221_X1 U11380 ( .B1(n10446), .B2(keyinput_g74), .C1(n10406), .C2(
        keyinput_g105), .A(n10318), .ZN(n10324) );
  XNOR2_X1 U11381 ( .A(SI_11_), .B(keyinput_g21), .ZN(n10322) );
  XNOR2_X1 U11382 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_g120), .ZN(n10321)
         );
  XNOR2_X1 U11383 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_g102), .ZN(n10320)
         );
  XNOR2_X1 U11384 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_g66), .ZN(n10319) );
  NAND4_X1 U11385 ( .A1(n10322), .A2(n10321), .A3(n10320), .A4(n10319), .ZN(
        n10323) );
  NOR3_X1 U11386 ( .A1(n10325), .A2(n10324), .A3(n10323), .ZN(n10350) );
  AOI22_X1 U11387 ( .A1(n10328), .A2(keyinput_g89), .B1(keyinput_g2), .B2(
        n10327), .ZN(n10326) );
  OAI221_X1 U11388 ( .B1(n10328), .B2(keyinput_g89), .C1(n10327), .C2(
        keyinput_g2), .A(n10326), .ZN(n10338) );
  AOI22_X1 U11389 ( .A1(n10331), .A2(keyinput_g85), .B1(keyinput_g27), .B2(
        n10330), .ZN(n10329) );
  OAI221_X1 U11390 ( .B1(n10331), .B2(keyinput_g85), .C1(n10330), .C2(
        keyinput_g27), .A(n10329), .ZN(n10337) );
  XOR2_X1 U11391 ( .A(n4759), .B(keyinput_g33), .Z(n10335) );
  XNOR2_X1 U11392 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_g92), .ZN(n10334) );
  XNOR2_X1 U11393 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_g119), .ZN(n10333)
         );
  XNOR2_X1 U11394 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_g90), .ZN(n10332) );
  NAND4_X1 U11395 ( .A1(n10335), .A2(n10334), .A3(n10333), .A4(n10332), .ZN(
        n10336) );
  NOR3_X1 U11396 ( .A1(n10338), .A2(n10337), .A3(n10336), .ZN(n10349) );
  AOI22_X1 U11397 ( .A1(n6345), .A2(keyinput_g65), .B1(n10490), .B2(
        keyinput_g70), .ZN(n10339) );
  OAI221_X1 U11398 ( .B1(n6345), .B2(keyinput_g65), .C1(n10490), .C2(
        keyinput_g70), .A(n10339), .ZN(n10347) );
  XNOR2_X1 U11399 ( .A(keyinput_g53), .B(n5974), .ZN(n10346) );
  XNOR2_X1 U11400 ( .A(keyinput_g46), .B(n10463), .ZN(n10345) );
  XNOR2_X1 U11401 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_g95), .ZN(n10343) );
  XNOR2_X1 U11402 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_g118), .ZN(n10342)
         );
  XNOR2_X1 U11403 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_g116), .ZN(n10341)
         );
  XNOR2_X1 U11404 ( .A(SI_23_), .B(keyinput_g9), .ZN(n10340) );
  NAND4_X1 U11405 ( .A1(n10343), .A2(n10342), .A3(n10341), .A4(n10340), .ZN(
        n10344) );
  NOR4_X1 U11406 ( .A1(n10347), .A2(n10346), .A3(n10345), .A4(n10344), .ZN(
        n10348) );
  NAND4_X1 U11407 ( .A1(n10351), .A2(n10350), .A3(n10349), .A4(n10348), .ZN(
        n10352) );
  NOR4_X1 U11408 ( .A1(n10355), .A2(n10354), .A3(n10353), .A4(n10352), .ZN(
        n10541) );
  OAI22_X1 U11409 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput_f99), .B1(SI_26_), 
        .B2(keyinput_f6), .ZN(n10356) );
  AOI221_X1 U11410 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput_f99), .C1(
        keyinput_f6), .C2(SI_26_), .A(n10356), .ZN(n10363) );
  OAI22_X1 U11411 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(keyinput_f68), .B1(
        P2_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .ZN(n10357) );
  AOI221_X1 U11412 ( .B1(P2_DATAO_REG_28__SCAN_IN), .B2(keyinput_f68), .C1(
        keyinput_f51), .C2(P2_REG3_REG_24__SCAN_IN), .A(n10357), .ZN(n10362)
         );
  OAI22_X1 U11413 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(keyinput_f86), .B1(
        keyinput_f59), .B2(P2_REG3_REG_2__SCAN_IN), .ZN(n10358) );
  AOI221_X1 U11414 ( .B1(P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_f86), .C1(
        P2_REG3_REG_2__SCAN_IN), .C2(keyinput_f59), .A(n10358), .ZN(n10361) );
  OAI22_X1 U11415 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput_f123), .B1(SI_8_), 
        .B2(keyinput_f24), .ZN(n10359) );
  AOI221_X1 U11416 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput_f123), .C1(
        keyinput_f24), .C2(SI_8_), .A(n10359), .ZN(n10360) );
  NAND4_X1 U11417 ( .A1(n10363), .A2(n10362), .A3(n10361), .A4(n10360), .ZN(
        n10391) );
  OAI22_X1 U11418 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(keyinput_f117), .B1(
        keyinput_f43), .B2(P2_REG3_REG_8__SCAN_IN), .ZN(n10364) );
  AOI221_X1 U11419 ( .B1(P1_IR_REG_27__SCAN_IN), .B2(keyinput_f117), .C1(
        P2_REG3_REG_8__SCAN_IN), .C2(keyinput_f43), .A(n10364), .ZN(n10371) );
  OAI22_X1 U11420 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(keyinput_f119), .B1(
        keyinput_f3), .B2(SI_29_), .ZN(n10365) );
  AOI221_X1 U11421 ( .B1(P1_IR_REG_29__SCAN_IN), .B2(keyinput_f119), .C1(
        SI_29_), .C2(keyinput_f3), .A(n10365), .ZN(n10370) );
  OAI22_X1 U11422 ( .A1(SI_17_), .A2(keyinput_f15), .B1(keyinput_f35), .B2(
        P2_REG3_REG_7__SCAN_IN), .ZN(n10366) );
  AOI221_X1 U11423 ( .B1(SI_17_), .B2(keyinput_f15), .C1(
        P2_REG3_REG_7__SCAN_IN), .C2(keyinput_f35), .A(n10366), .ZN(n10369) );
  OAI22_X1 U11424 ( .A1(SI_13_), .A2(keyinput_f19), .B1(keyinput_f40), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n10367) );
  AOI221_X1 U11425 ( .B1(SI_13_), .B2(keyinput_f19), .C1(
        P2_REG3_REG_3__SCAN_IN), .C2(keyinput_f40), .A(n10367), .ZN(n10368) );
  NAND4_X1 U11426 ( .A1(n10371), .A2(n10370), .A3(n10369), .A4(n10368), .ZN(
        n10390) );
  OAI22_X1 U11427 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(keyinput_f121), .B1(
        keyinput_f125), .B2(P1_D_REG_3__SCAN_IN), .ZN(n10372) );
  AOI221_X1 U11428 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(keyinput_f121), .C1(
        P1_D_REG_3__SCAN_IN), .C2(keyinput_f125), .A(n10372), .ZN(n10379) );
  OAI22_X1 U11429 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput_f112), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_f69), .ZN(n10373) );
  AOI221_X1 U11430 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(keyinput_f112), .C1(
        keyinput_f69), .C2(P2_DATAO_REG_27__SCAN_IN), .A(n10373), .ZN(n10378)
         );
  OAI22_X1 U11431 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(keyinput_f116), .B1(
        keyinput_f57), .B2(P2_REG3_REG_22__SCAN_IN), .ZN(n10374) );
  AOI221_X1 U11432 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(keyinput_f116), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_f57), .A(n10374), .ZN(n10377)
         );
  OAI22_X1 U11433 ( .A1(P1_D_REG_5__SCAN_IN), .A2(keyinput_f127), .B1(
        keyinput_f84), .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n10375) );
  AOI221_X1 U11434 ( .B1(P1_D_REG_5__SCAN_IN), .B2(keyinput_f127), .C1(
        P2_DATAO_REG_12__SCAN_IN), .C2(keyinput_f84), .A(n10375), .ZN(n10376)
         );
  NAND4_X1 U11435 ( .A1(n10379), .A2(n10378), .A3(n10377), .A4(n10376), .ZN(
        n10389) );
  OAI22_X1 U11436 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(keyinput_f72), .B1(
        keyinput_f28), .B2(SI_4_), .ZN(n10380) );
  AOI221_X1 U11437 ( .B1(P2_DATAO_REG_24__SCAN_IN), .B2(keyinput_f72), .C1(
        SI_4_), .C2(keyinput_f28), .A(n10380), .ZN(n10387) );
  OAI22_X1 U11438 ( .A1(SI_3_), .A2(keyinput_f29), .B1(P2_WR_REG_SCAN_IN), 
        .B2(keyinput_f0), .ZN(n10381) );
  AOI221_X1 U11439 ( .B1(SI_3_), .B2(keyinput_f29), .C1(keyinput_f0), .C2(
        P2_WR_REG_SCAN_IN), .A(n10381), .ZN(n10386) );
  OAI22_X1 U11440 ( .A1(SI_14_), .A2(keyinput_f18), .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .ZN(n10382) );
  AOI221_X1 U11441 ( .B1(SI_14_), .B2(keyinput_f18), .C1(keyinput_f53), .C2(
        P2_REG3_REG_9__SCAN_IN), .A(n10382), .ZN(n10385) );
  OAI22_X1 U11442 ( .A1(SI_30_), .A2(keyinput_f2), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(keyinput_f66), .ZN(n10383) );
  AOI221_X1 U11443 ( .B1(SI_30_), .B2(keyinput_f2), .C1(keyinput_f66), .C2(
        P2_DATAO_REG_30__SCAN_IN), .A(n10383), .ZN(n10384) );
  NAND4_X1 U11444 ( .A1(n10387), .A2(n10386), .A3(n10385), .A4(n10384), .ZN(
        n10388) );
  NOR4_X1 U11445 ( .A1(n10391), .A2(n10390), .A3(n10389), .A4(n10388), .ZN(
        n10537) );
  OAI22_X1 U11446 ( .A1(SI_19_), .A2(keyinput_f13), .B1(SI_5_), .B2(
        keyinput_f27), .ZN(n10392) );
  AOI221_X1 U11447 ( .B1(SI_19_), .B2(keyinput_f13), .C1(keyinput_f27), .C2(
        SI_5_), .A(n10392), .ZN(n10399) );
  OAI22_X1 U11448 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(keyinput_f118), .B1(
        keyinput_f38), .B2(P2_REG3_REG_23__SCAN_IN), .ZN(n10393) );
  AOI221_X1 U11449 ( .B1(P1_IR_REG_28__SCAN_IN), .B2(keyinput_f118), .C1(
        P2_REG3_REG_23__SCAN_IN), .C2(keyinput_f38), .A(n10393), .ZN(n10398)
         );
  OAI22_X1 U11450 ( .A1(SI_27_), .A2(keyinput_f5), .B1(keyinput_f23), .B2(
        SI_9_), .ZN(n10394) );
  AOI221_X1 U11451 ( .B1(SI_27_), .B2(keyinput_f5), .C1(SI_9_), .C2(
        keyinput_f23), .A(n10394), .ZN(n10397) );
  OAI22_X1 U11452 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput_f110), .B1(
        keyinput_f58), .B2(P2_REG3_REG_11__SCAN_IN), .ZN(n10395) );
  AOI221_X1 U11453 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput_f110), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_f58), .A(n10395), .ZN(n10396)
         );
  NAND4_X1 U11454 ( .A1(n10399), .A2(n10398), .A3(n10397), .A4(n10396), .ZN(
        n10535) );
  OAI22_X1 U11455 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(keyinput_f98), .B1(
        P1_D_REG_0__SCAN_IN), .B2(keyinput_f122), .ZN(n10400) );
  AOI221_X1 U11456 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(keyinput_f98), .C1(
        keyinput_f122), .C2(P1_D_REG_0__SCAN_IN), .A(n10400), .ZN(n10426) );
  OAI22_X1 U11457 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(keyinput_f108), .B1(
        keyinput_f20), .B2(SI_12_), .ZN(n10401) );
  AOI221_X1 U11458 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(keyinput_f108), .C1(
        SI_12_), .C2(keyinput_f20), .A(n10401), .ZN(n10404) );
  OAI22_X1 U11459 ( .A1(P1_D_REG_2__SCAN_IN), .A2(keyinput_f124), .B1(
        P2_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .ZN(n10402) );
  AOI221_X1 U11460 ( .B1(P1_D_REG_2__SCAN_IN), .B2(keyinput_f124), .C1(
        keyinput_f61), .C2(P2_REG3_REG_6__SCAN_IN), .A(n10402), .ZN(n10403) );
  OAI211_X1 U11461 ( .C1(n10406), .C2(keyinput_f105), .A(n10404), .B(n10403), 
        .ZN(n10405) );
  AOI21_X1 U11462 ( .B1(n10406), .B2(keyinput_f105), .A(n10405), .ZN(n10425)
         );
  AOI22_X1 U11463 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput_f52), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_f85), .ZN(n10407) );
  OAI221_X1 U11464 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_f52), .C1(
        P2_DATAO_REG_11__SCAN_IN), .C2(keyinput_f85), .A(n10407), .ZN(n10414)
         );
  AOI22_X1 U11465 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput_f65), .B1(
        P1_IR_REG_11__SCAN_IN), .B2(keyinput_f101), .ZN(n10408) );
  OAI221_X1 U11466 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(keyinput_f65), .C1(
        P1_IR_REG_11__SCAN_IN), .C2(keyinput_f101), .A(n10408), .ZN(n10413) );
  AOI22_X1 U11467 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_f47), .B1(
        SI_20_), .B2(keyinput_f12), .ZN(n10409) );
  OAI221_X1 U11468 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .C1(
        SI_20_), .C2(keyinput_f12), .A(n10409), .ZN(n10412) );
  AOI22_X1 U11469 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(keyinput_f89), .B1(
        SI_10_), .B2(keyinput_f22), .ZN(n10410) );
  OAI221_X1 U11470 ( .B1(P2_DATAO_REG_7__SCAN_IN), .B2(keyinput_f89), .C1(
        SI_10_), .C2(keyinput_f22), .A(n10410), .ZN(n10411) );
  NOR4_X1 U11471 ( .A1(n10414), .A2(n10413), .A3(n10412), .A4(n10411), .ZN(
        n10424) );
  AOI22_X1 U11472 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(keyinput_f83), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_f76), .ZN(n10415) );
  OAI221_X1 U11473 ( .B1(P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_f83), .C1(
        P2_DATAO_REG_20__SCAN_IN), .C2(keyinput_f76), .A(n10415), .ZN(n10422)
         );
  AOI22_X1 U11474 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_f37), .B1(
        P1_IR_REG_25__SCAN_IN), .B2(keyinput_f115), .ZN(n10416) );
  OAI221_X1 U11475 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_f37), .C1(
        P1_IR_REG_25__SCAN_IN), .C2(keyinput_f115), .A(n10416), .ZN(n10421) );
  AOI22_X1 U11476 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_f42), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(keyinput_f81), .ZN(n10417) );
  OAI221_X1 U11477 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .C1(
        P2_DATAO_REG_15__SCAN_IN), .C2(keyinput_f81), .A(n10417), .ZN(n10420)
         );
  AOI22_X1 U11478 ( .A1(SI_23_), .A2(keyinput_f9), .B1(P1_IR_REG_14__SCAN_IN), 
        .B2(keyinput_f104), .ZN(n10418) );
  OAI221_X1 U11479 ( .B1(SI_23_), .B2(keyinput_f9), .C1(P1_IR_REG_14__SCAN_IN), 
        .C2(keyinput_f104), .A(n10418), .ZN(n10419) );
  NOR4_X1 U11480 ( .A1(n10422), .A2(n10421), .A3(n10420), .A4(n10419), .ZN(
        n10423) );
  NAND4_X1 U11481 ( .A1(n10426), .A2(n10425), .A3(n10424), .A4(n10423), .ZN(
        n10534) );
  AOI22_X1 U11482 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput_f80), .B1(
        SI_25_), .B2(keyinput_f7), .ZN(n10427) );
  OAI221_X1 U11483 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput_f80), .C1(
        SI_25_), .C2(keyinput_f7), .A(n10427), .ZN(n10434) );
  AOI22_X1 U11484 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_f34), .B1(
        P1_D_REG_4__SCAN_IN), .B2(keyinput_f126), .ZN(n10428) );
  OAI221_X1 U11485 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_f34), .C1(
        P1_D_REG_4__SCAN_IN), .C2(keyinput_f126), .A(n10428), .ZN(n10433) );
  AOI22_X1 U11486 ( .A1(SI_1_), .A2(keyinput_f31), .B1(P1_IR_REG_0__SCAN_IN), 
        .B2(keyinput_f90), .ZN(n10429) );
  OAI221_X1 U11487 ( .B1(SI_1_), .B2(keyinput_f31), .C1(P1_IR_REG_0__SCAN_IN), 
        .C2(keyinput_f90), .A(n10429), .ZN(n10432) );
  AOI22_X1 U11488 ( .A1(SI_2_), .A2(keyinput_f30), .B1(P1_IR_REG_21__SCAN_IN), 
        .B2(keyinput_f111), .ZN(n10430) );
  OAI221_X1 U11489 ( .B1(SI_2_), .B2(keyinput_f30), .C1(P1_IR_REG_21__SCAN_IN), 
        .C2(keyinput_f111), .A(n10430), .ZN(n10431) );
  NOR4_X1 U11490 ( .A1(n10434), .A2(n10433), .A3(n10432), .A4(n10431), .ZN(
        n10474) );
  AOI22_X1 U11491 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_f41), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_f87), .ZN(n10435) );
  OAI221_X1 U11492 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .C1(
        P2_DATAO_REG_9__SCAN_IN), .C2(keyinput_f87), .A(n10435), .ZN(n10444)
         );
  AOI22_X1 U11493 ( .A1(SI_6_), .A2(keyinput_f26), .B1(P1_IR_REG_6__SCAN_IN), 
        .B2(keyinput_f96), .ZN(n10436) );
  OAI221_X1 U11494 ( .B1(SI_6_), .B2(keyinput_f26), .C1(P1_IR_REG_6__SCAN_IN), 
        .C2(keyinput_f96), .A(n10436), .ZN(n10443) );
  AOI22_X1 U11495 ( .A1(SI_31_), .A2(keyinput_f1), .B1(SI_15_), .B2(
        keyinput_f17), .ZN(n10437) );
  OAI221_X1 U11496 ( .B1(SI_31_), .B2(keyinput_f1), .C1(SI_15_), .C2(
        keyinput_f17), .A(n10437), .ZN(n10442) );
  AOI22_X1 U11497 ( .A1(n10440), .A2(keyinput_f88), .B1(keyinput_f55), .B2(
        n10439), .ZN(n10438) );
  OAI221_X1 U11498 ( .B1(n10440), .B2(keyinput_f88), .C1(n10439), .C2(
        keyinput_f55), .A(n10438), .ZN(n10441) );
  NOR4_X1 U11499 ( .A1(n10444), .A2(n10443), .A3(n10442), .A4(n10441), .ZN(
        n10473) );
  AOI22_X1 U11500 ( .A1(n10447), .A2(keyinput_f79), .B1(n10446), .B2(
        keyinput_f74), .ZN(n10445) );
  OAI221_X1 U11501 ( .B1(n10447), .B2(keyinput_f79), .C1(n10446), .C2(
        keyinput_f74), .A(n10445), .ZN(n10457) );
  AOI22_X1 U11502 ( .A1(n10450), .A2(keyinput_f60), .B1(n10449), .B2(
        keyinput_f25), .ZN(n10448) );
  OAI221_X1 U11503 ( .B1(n10450), .B2(keyinput_f60), .C1(n10449), .C2(
        keyinput_f25), .A(n10448), .ZN(n10456) );
  XOR2_X1 U11504 ( .A(n8429), .B(keyinput_f50), .Z(n10454) );
  XNOR2_X1 U11505 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_f39), .ZN(n10453)
         );
  XNOR2_X1 U11506 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_f114), .ZN(n10452)
         );
  XNOR2_X1 U11507 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_f94), .ZN(n10451) );
  NAND4_X1 U11508 ( .A1(n10454), .A2(n10453), .A3(n10452), .A4(n10451), .ZN(
        n10455) );
  NOR3_X1 U11509 ( .A1(n10457), .A2(n10456), .A3(n10455), .ZN(n10472) );
  AOI22_X1 U11510 ( .A1(n10460), .A2(keyinput_f14), .B1(n10459), .B2(
        keyinput_f11), .ZN(n10458) );
  OAI221_X1 U11511 ( .B1(n10460), .B2(keyinput_f14), .C1(n10459), .C2(
        keyinput_f11), .A(n10458), .ZN(n10470) );
  AOI22_X1 U11512 ( .A1(n10463), .A2(keyinput_f46), .B1(n10462), .B2(
        keyinput_f63), .ZN(n10461) );
  OAI221_X1 U11513 ( .B1(n10463), .B2(keyinput_f46), .C1(n10462), .C2(
        keyinput_f63), .A(n10461), .ZN(n10469) );
  XOR2_X1 U11514 ( .A(n5791), .B(keyinput_f4), .Z(n10467) );
  XNOR2_X1 U11515 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_f102), .ZN(n10466)
         );
  XNOR2_X1 U11516 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_f77), .ZN(n10465) );
  XNOR2_X1 U11517 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_f103), .ZN(n10464)
         );
  NAND4_X1 U11518 ( .A1(n10467), .A2(n10466), .A3(n10465), .A4(n10464), .ZN(
        n10468) );
  NOR3_X1 U11519 ( .A1(n10470), .A2(n10469), .A3(n10468), .ZN(n10471) );
  NAND4_X1 U11520 ( .A1(n10474), .A2(n10473), .A3(n10472), .A4(n10471), .ZN(
        n10533) );
  AOI22_X1 U11521 ( .A1(n10477), .A2(keyinput_f71), .B1(keyinput_f67), .B2(
        n10476), .ZN(n10475) );
  OAI221_X1 U11522 ( .B1(n10477), .B2(keyinput_f71), .C1(n10476), .C2(
        keyinput_f67), .A(n10475), .ZN(n10486) );
  XOR2_X1 U11523 ( .A(SI_11_), .B(keyinput_f21), .Z(n10485) );
  XNOR2_X1 U11524 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_f75), .ZN(n10481) );
  XNOR2_X1 U11525 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_f54), .ZN(n10480)
         );
  XNOR2_X1 U11526 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_f107), .ZN(n10479)
         );
  XNOR2_X1 U11527 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_f95), .ZN(n10478) );
  NAND4_X1 U11528 ( .A1(n10481), .A2(n10480), .A3(n10479), .A4(n10478), .ZN(
        n10484) );
  XNOR2_X1 U11529 ( .A(n10482), .B(keyinput_f93), .ZN(n10483) );
  NOR4_X1 U11530 ( .A1(n10486), .A2(n10485), .A3(n10484), .A4(n10483), .ZN(
        n10531) );
  AOI22_X1 U11531 ( .A1(n10488), .A2(keyinput_f62), .B1(n4759), .B2(
        keyinput_f33), .ZN(n10487) );
  OAI221_X1 U11532 ( .B1(n10488), .B2(keyinput_f62), .C1(n4759), .C2(
        keyinput_f33), .A(n10487), .ZN(n10501) );
  AOI22_X1 U11533 ( .A1(n10491), .A2(keyinput_f45), .B1(n10490), .B2(
        keyinput_f70), .ZN(n10489) );
  OAI221_X1 U11534 ( .B1(n10491), .B2(keyinput_f45), .C1(n10490), .C2(
        keyinput_f70), .A(n10489), .ZN(n10500) );
  AOI22_X1 U11535 ( .A1(n10494), .A2(keyinput_f97), .B1(n10493), .B2(
        keyinput_f100), .ZN(n10492) );
  OAI221_X1 U11536 ( .B1(n10494), .B2(keyinput_f97), .C1(n10493), .C2(
        keyinput_f100), .A(n10492), .ZN(n10499) );
  XNOR2_X1 U11537 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_f106), .ZN(n10497)
         );
  XNOR2_X1 U11538 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_f91), .ZN(n10496) );
  NAND2_X1 U11539 ( .A1(n10497), .A2(n10496), .ZN(n10498) );
  NOR4_X1 U11540 ( .A1(n10501), .A2(n10500), .A3(n10499), .A4(n10498), .ZN(
        n10530) );
  INV_X1 U11541 ( .A(P2_B_REG_SCAN_IN), .ZN(n10503) );
  AOI22_X1 U11542 ( .A1(n10503), .A2(keyinput_f64), .B1(keyinput_f49), .B2(
        n5912), .ZN(n10502) );
  OAI221_X1 U11543 ( .B1(n10503), .B2(keyinput_f64), .C1(n5912), .C2(
        keyinput_f49), .A(n10502), .ZN(n10515) );
  AOI22_X1 U11544 ( .A1(n10506), .A2(keyinput_f8), .B1(keyinput_f78), .B2(
        n10505), .ZN(n10504) );
  OAI221_X1 U11545 ( .B1(n10506), .B2(keyinput_f8), .C1(n10505), .C2(
        keyinput_f78), .A(n10504), .ZN(n10514) );
  AOI22_X1 U11546 ( .A1(n10509), .A2(keyinput_f56), .B1(n10508), .B2(
        keyinput_f82), .ZN(n10507) );
  OAI221_X1 U11547 ( .B1(n10509), .B2(keyinput_f56), .C1(n10508), .C2(
        keyinput_f82), .A(n10507), .ZN(n10513) );
  XNOR2_X1 U11548 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_f120), .ZN(n10511)
         );
  XNOR2_X1 U11549 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_f36), .ZN(n10510)
         );
  NAND2_X1 U11550 ( .A1(n10511), .A2(n10510), .ZN(n10512) );
  NOR4_X1 U11551 ( .A1(n10515), .A2(n10514), .A3(n10513), .A4(n10512), .ZN(
        n10529) );
  AOI22_X1 U11552 ( .A1(n10517), .A2(keyinput_f10), .B1(keyinput_f16), .B2(
        n5534), .ZN(n10516) );
  OAI221_X1 U11553 ( .B1(n10517), .B2(keyinput_f10), .C1(n5534), .C2(
        keyinput_f16), .A(n10516), .ZN(n10527) );
  AOI22_X1 U11554 ( .A1(n10520), .A2(keyinput_f48), .B1(n10519), .B2(
        keyinput_f113), .ZN(n10518) );
  OAI221_X1 U11555 ( .B1(n10520), .B2(keyinput_f48), .C1(n10519), .C2(
        keyinput_f113), .A(n10518), .ZN(n10526) );
  XOR2_X1 U11556 ( .A(n5847), .B(keyinput_f44), .Z(n10524) );
  XNOR2_X1 U11557 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_f109), .ZN(n10523)
         );
  XNOR2_X1 U11558 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_f73), .ZN(n10522) );
  XNOR2_X1 U11559 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_f92), .ZN(n10521) );
  NAND4_X1 U11560 ( .A1(n10524), .A2(n10523), .A3(n10522), .A4(n10521), .ZN(
        n10525) );
  NOR3_X1 U11561 ( .A1(n10527), .A2(n10526), .A3(n10525), .ZN(n10528) );
  NAND4_X1 U11562 ( .A1(n10531), .A2(n10530), .A3(n10529), .A4(n10528), .ZN(
        n10532) );
  NOR4_X1 U11563 ( .A1(n10535), .A2(n10534), .A3(n10533), .A4(n10532), .ZN(
        n10536) );
  AOI22_X1 U11564 ( .A1(n10537), .A2(n10536), .B1(keyinput_f32), .B2(SI_0_), 
        .ZN(n10538) );
  OAI21_X1 U11565 ( .B1(keyinput_f32), .B2(SI_0_), .A(n10538), .ZN(n10539) );
  OAI21_X1 U11566 ( .B1(n5308), .B2(keyinput_g32), .A(n10539), .ZN(n10540) );
  AOI211_X1 U11567 ( .C1(n5308), .C2(keyinput_g32), .A(n10541), .B(n10540), 
        .ZN(n10544) );
  XNOR2_X1 U11568 ( .A(n10542), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n10543) );
  XNOR2_X1 U11569 ( .A(n10544), .B(n10543), .ZN(n10545) );
  XNOR2_X1 U11570 ( .A(n10546), .B(n10545), .ZN(ADD_1068_U4) );
  XNOR2_X1 U11571 ( .A(n10548), .B(n10547), .ZN(ADD_1068_U47) );
  XOR2_X1 U11572 ( .A(n10550), .B(n10549), .Z(ADD_1068_U54) );
  XNOR2_X1 U11573 ( .A(n10552), .B(n10551), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11574 ( .A(n10554), .B(n10553), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11575 ( .A(n10556), .B(n10555), .ZN(ADD_1068_U48) );
  XNOR2_X1 U11576 ( .A(n10558), .B(n10557), .ZN(ADD_1068_U50) );
  XOR2_X1 U11577 ( .A(n10560), .B(n10559), .Z(ADD_1068_U53) );
  XNOR2_X1 U11578 ( .A(n10562), .B(n10561), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U5031 ( .A(n7152), .Z(n8128) );
  CLKBUF_X1 U5230 ( .A(n5883), .Z(n7096) );
endmodule

