

module b15_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, 
        DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, 
        DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, 
        DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, 
        DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, 
        DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, 
        HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712;

  XNOR2_X1 U3692 ( .A(n4881), .B(n4880), .ZN(n6579) );
  OR2_X1 U3693 ( .A1(n4936), .A2(n4879), .ZN(n4881) );
  NAND2_X1 U3694 ( .A1(n4613), .A2(n4612), .ZN(n6651) );
  NAND2_X1 U3695 ( .A1(n6936), .A2(n4178), .ZN(n4181) );
  AND2_X2 U3696 ( .A1(n3941), .A2(n3924), .ZN(n5085) );
  CLKBUF_X2 U3697 ( .A(n3850), .Z(n3660) );
  CLKBUF_X2 U3698 ( .A(n3974), .Z(n4730) );
  CLKBUF_X2 U3699 ( .A(n3968), .Z(n4718) );
  AND2_X1 U3700 ( .A1(n3940), .A2(n5172), .ZN(n4885) );
  BUF_X2 U3701 ( .A(n3909), .Z(n5172) );
  AND2_X1 U3702 ( .A1(n5027), .A2(n5307), .ZN(n3855) );
  AND2_X1 U3703 ( .A1(n6513), .A2(n5033), .ZN(n3968) );
  AND2_X1 U3704 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5308) );
  CLKBUF_X1 U3705 ( .A(n7611), .Z(n3658) );
  NOR2_X1 U3706 ( .A1(n7309), .A2(n7135), .ZN(n7611) );
  NOR2_X1 U3707 ( .A1(n3924), .A2(n7616), .ZN(n3918) );
  OAI21_X1 U3708 ( .B1(n4956), .B2(n3918), .A(n4784), .ZN(n3903) );
  AND2_X1 U3709 ( .A1(n5030), .A2(n3926), .ZN(n3953) );
  AND2_X1 U3710 ( .A1(n3941), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4208) );
  NOR2_X1 U3711 ( .A1(n3923), .A2(n3945), .ZN(n4887) );
  AND2_X2 U3712 ( .A1(n5039), .A2(n6513), .ZN(n3850) );
  NAND2_X2 U3713 ( .A1(n4932), .A2(n5085), .ZN(n4795) );
  NOR2_X1 U3714 ( .A1(n3941), .A2(n3924), .ZN(n5088) );
  INV_X1 U3716 ( .A(n4187), .ZN(n7066) );
  INV_X1 U3717 ( .A(n3924), .ZN(n5228) );
  INV_X1 U3718 ( .A(n7541), .ZN(n7504) );
  NAND2_X1 U3719 ( .A1(n7384), .A2(n4904), .ZN(n7383) );
  NOR2_X2 U3720 ( .A1(n3785), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5039)
         );
  INV_X1 U3721 ( .A(n7521), .ZN(n7535) );
  AND2_X4 U3722 ( .A1(n5039), .A2(n5308), .ZN(n3866) );
  OAI222_X1 U3723 ( .A1(n5809), .A2(n5125), .B1(n5805), .B2(n5719), .C1(n5718), 
        .C2(n7129), .ZN(U3463) );
  BUF_X8 U3724 ( .A(n3871), .Z(n3665) );
  OAI21_X2 U3725 ( .B1(n6861), .B2(n3683), .A(n3747), .ZN(n6852) );
  NAND2_X2 U3726 ( .A1(n6882), .A2(n4184), .ZN(n6861) );
  OR2_X1 U3727 ( .A1(n4086), .A2(n7349), .ZN(n7268) );
  AOI21_X2 U3728 ( .B1(n6432), .B2(n6433), .A(n6435), .ZN(n7288) );
  AND2_X4 U3729 ( .A1(n3799), .A2(n5310), .ZN(n4000) );
  OAI21_X2 U3730 ( .B1(n6637), .B2(n6635), .A(n6636), .ZN(n6846) );
  NOR2_X4 U3731 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3708) );
  NOR2_X1 U3732 ( .A1(n3919), .A2(n5177), .ZN(n3925) );
  OAI21_X2 U3733 ( .B1(n6024), .B2(n6023), .A(n4134), .ZN(n6432) );
  OR2_X1 U3734 ( .A1(n6638), .A2(n6639), .ZN(n6641) );
  NOR3_X1 U3735 ( .A1(n6709), .A2(n3724), .A3(n3723), .ZN(n3722) );
  BUF_X1 U3736 ( .A(n5124), .Z(n3661) );
  OR2_X1 U3737 ( .A1(n3675), .A2(n6707), .ZN(n6709) );
  OR2_X1 U3738 ( .A1(n6745), .A2(n6744), .ZN(n6747) );
  NOR2_X1 U3739 ( .A1(n6484), .A2(n6483), .ZN(n6503) );
  NAND2_X1 U3740 ( .A1(n5083), .A2(n5085), .ZN(n3710) );
  NAND2_X1 U3741 ( .A1(n4256), .A2(n6575), .ZN(n3905) );
  INV_X4 U3742 ( .A(n4874), .ZN(n4932) );
  INV_X1 U3743 ( .A(n3901), .ZN(n3904) );
  BUF_X2 U3744 ( .A(n4367), .Z(n4727) );
  BUF_X2 U3745 ( .A(n3865), .Z(n4732) );
  BUF_X2 U3746 ( .A(n3855), .Z(n4731) );
  AND2_X2 U3747 ( .A1(n5027), .A2(n6513), .ZN(n4367) );
  OR2_X1 U3748 ( .A1(n6581), .A2(n6976), .ZN(n3748) );
  OAI21_X1 U3749 ( .B1(n7040), .B2(n7066), .A(n7032), .ZN(n6888) );
  XNOR2_X1 U3750 ( .A(n3730), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4949)
         );
  OR2_X1 U3751 ( .A1(n6880), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6868)
         );
  OR2_X1 U3752 ( .A1(n6521), .A2(n6520), .ZN(n3707) );
  AND2_X1 U3753 ( .A1(n3674), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3706)
         );
  OAI21_X1 U3754 ( .B1(n6522), .B2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n4187), 
        .ZN(n6539) );
  AND2_X2 U3755 ( .A1(n6501), .A2(n3755), .ZN(n6730) );
  AND2_X1 U3756 ( .A1(n4929), .A2(n4928), .ZN(n4930) );
  INV_X1 U3757 ( .A(n3697), .ZN(n3695) );
  NAND2_X1 U3758 ( .A1(n3743), .A2(n3676), .ZN(n3740) );
  NAND2_X1 U3759 ( .A1(n3743), .A2(n3742), .ZN(n3741) );
  OR2_X1 U3760 ( .A1(n4295), .A2(n4432), .ZN(n4300) );
  OAI21_X1 U3761 ( .B1(n4295), .B2(n4222), .A(n4132), .ZN(n4133) );
  AND2_X1 U3762 ( .A1(n4154), .A2(n4153), .ZN(n4307) );
  OAI21_X1 U3763 ( .B1(n4301), .B2(n4432), .A(n4306), .ZN(n5597) );
  NAND2_X2 U3764 ( .A1(n4167), .A2(n4166), .ZN(n4171) );
  NAND2_X1 U3765 ( .A1(n3727), .A2(n3750), .ZN(n4167) );
  OR2_X1 U3766 ( .A1(n7062), .A2(n4900), .ZN(n7353) );
  NAND2_X1 U3767 ( .A1(n4254), .A2(n4607), .ZN(n5098) );
  AND2_X1 U3768 ( .A1(n5080), .A2(n5079), .ZN(n5099) );
  NAND2_X1 U3769 ( .A1(n4051), .A2(n4050), .ZN(n5158) );
  NAND2_X1 U3770 ( .A1(n4782), .A2(n7581), .ZN(n4909) );
  NAND2_X1 U3771 ( .A1(n4993), .A2(n4269), .ZN(n5079) );
  INV_X2 U3772 ( .A(n6780), .ZN(n3659) );
  OR2_X1 U3773 ( .A1(n4995), .A2(n4996), .ZN(n4993) );
  NAND2_X2 U3775 ( .A1(n4073), .A2(n4072), .ZN(n5487) );
  OR3_X1 U3776 ( .A1(n5837), .A2(n6451), .A3(n6450), .ZN(n6484) );
  NAND2_X1 U3777 ( .A1(n4069), .A2(n4068), .ZN(n4073) );
  AND2_X1 U3778 ( .A1(n5813), .A2(n5812), .ZN(n5839) );
  AND2_X1 U3779 ( .A1(n5654), .A2(n3680), .ZN(n5813) );
  AND2_X1 U3780 ( .A1(n3998), .A2(n3997), .ZN(n3983) );
  AND2_X1 U3781 ( .A1(n5652), .A2(n5651), .ZN(n5654) );
  AND2_X1 U3782 ( .A1(n3956), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4033) );
  NOR2_X1 U3783 ( .A1(n5722), .A2(n5110), .ZN(n5652) );
  AND4_X1 U3784 ( .A1(n3953), .A2(n3952), .A3(n3951), .A4(n3950), .ZN(n3954)
         );
  AND2_X1 U3785 ( .A1(n3689), .A2(n3688), .ZN(n3927) );
  NAND2_X1 U3786 ( .A1(n4861), .A2(n6653), .ZN(n3723) );
  OR2_X1 U3787 ( .A1(n4068), .A2(n4071), .ZN(n4072) );
  NAND2_X1 U3788 ( .A1(n4791), .A2(n4790), .ZN(n4794) );
  AND2_X2 U3789 ( .A1(n3924), .A2(n5172), .ZN(n4232) );
  INV_X2 U3790 ( .A(n4713), .ZN(n4749) );
  NAND2_X2 U3791 ( .A1(n4029), .A2(n4027), .ZN(n4231) );
  AND2_X1 U3792 ( .A1(n4261), .A2(n3945), .ZN(n3908) );
  OAI21_X1 U3793 ( .B1(n3909), .B2(n3904), .A(n4237), .ZN(n3919) );
  NAND2_X1 U3794 ( .A1(n3904), .A2(n4237), .ZN(n4261) );
  AND2_X1 U3795 ( .A1(n3798), .A2(n3797), .ZN(n3811) );
  INV_X4 U3796 ( .A(n3941), .ZN(n5140) );
  OR2_X2 U3797 ( .A1(n3839), .A2(n3838), .ZN(n5177) );
  AND4_X1 U3798 ( .A1(n3815), .A2(n3814), .A3(n3813), .A4(n3812), .ZN(n3821)
         );
  AND4_X1 U3799 ( .A1(n3887), .A2(n3886), .A3(n3885), .A4(n3884), .ZN(n3899)
         );
  AND4_X1 U3800 ( .A1(n3891), .A2(n3890), .A3(n3889), .A4(n3888), .ZN(n3898)
         );
  AND4_X1 U3801 ( .A1(n3883), .A2(n3882), .A3(n3881), .A4(n3880), .ZN(n3900)
         );
  AND4_X1 U3802 ( .A1(n3803), .A2(n3802), .A3(n3801), .A4(n3800), .ZN(n3810)
         );
  AND4_X1 U3803 ( .A1(n3808), .A2(n3807), .A3(n3806), .A4(n3805), .ZN(n3809)
         );
  AND4_X1 U3804 ( .A1(n3819), .A2(n3818), .A3(n3817), .A4(n3816), .ZN(n3820)
         );
  INV_X2 U3805 ( .A(n6976), .ZN(n7297) );
  BUF_X2 U3806 ( .A(n4655), .Z(n4721) );
  BUF_X2 U3807 ( .A(n4118), .Z(n4719) );
  BUF_X4 U3808 ( .A(n3871), .Z(n3666) );
  BUF_X2 U3809 ( .A(n3975), .Z(n4539) );
  CLKBUF_X1 U3810 ( .A(n3892), .Z(n4722) );
  AND2_X2 U3811 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5033) );
  AOI21_X1 U3812 ( .B1(n4263), .B2(n7318), .A(n4024), .ZN(n4069) );
  NAND2_X2 U3813 ( .A1(n4770), .A2(n3910), .ZN(n4783) );
  INV_X2 U3814 ( .A(n3927), .ZN(n4770) );
  NAND2_X1 U3815 ( .A1(n3706), .A2(n3707), .ZN(n6834) );
  OR2_X2 U3816 ( .A1(n3681), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6978)
         );
  XNOR2_X1 U3817 ( .A(n5329), .B(n5330), .ZN(n5124) );
  NAND2_X1 U3818 ( .A1(n6942), .A2(n4177), .ZN(n6936) );
  XNOR2_X1 U3819 ( .A(n6556), .B(n4950), .ZN(n6581) );
  AND2_X2 U3820 ( .A1(n6852), .A2(n6853), .ZN(n6519) );
  NAND2_X2 U3821 ( .A1(n3821), .A2(n3820), .ZN(n3901) );
  AOI21_X2 U3822 ( .B1(n5066), .B2(n5065), .A(n4113), .ZN(n6024) );
  AND2_X4 U3823 ( .A1(n5068), .A2(n5107), .ZN(n5106) );
  AND2_X2 U3824 ( .A1(n5007), .A2(n5067), .ZN(n5068) );
  NAND2_X2 U3825 ( .A1(n6730), .A2(n6782), .ZN(n6716) );
  XNOR2_X2 U3826 ( .A(n4059), .B(n4058), .ZN(n4255) );
  NAND2_X2 U3827 ( .A1(n3996), .A2(n3995), .ZN(n4059) );
  NAND2_X2 U3828 ( .A1(n3962), .A2(n3964), .ZN(n5329) );
  AND2_X2 U3829 ( .A1(n6681), .A2(n6684), .ZN(n6682) );
  NOR2_X2 U3830 ( .A1(n6716), .A2(n3759), .ZN(n6681) );
  NOR2_X1 U3831 ( .A1(n6651), .A2(n3769), .ZN(n6625) );
  AND2_X1 U3832 ( .A1(n6513), .A2(n5033), .ZN(n3662) );
  AND2_X1 U3833 ( .A1(n6513), .A2(n5033), .ZN(n3663) );
  NAND2_X4 U3834 ( .A1(n3776), .A2(n3700), .ZN(n4237) );
  NOR2_X2 U3835 ( .A1(n3702), .A2(n3701), .ZN(n3700) );
  NOR2_X2 U3836 ( .A1(n5147), .A2(n3751), .ZN(n5831) );
  NAND2_X2 U3837 ( .A1(n5106), .A2(n4317), .ZN(n5147) );
  XNOR2_X2 U3838 ( .A(n4414), .B(n4415), .ZN(n6481) );
  NAND2_X2 U3839 ( .A1(n5329), .A2(n3966), .ZN(n5125) );
  AND2_X4 U3840 ( .A1(n5027), .A2(n5308), .ZN(n4702) );
  AND2_X4 U3841 ( .A1(n5033), .A2(n3804), .ZN(n3664) );
  INV_X1 U3842 ( .A(n6425), .ZN(n3743) );
  AND2_X1 U3843 ( .A1(n4232), .A2(n4165), .ZN(n4166) );
  BUF_X1 U3844 ( .A(n4702), .Z(n4729) );
  INV_X1 U3845 ( .A(n4232), .ZN(n4222) );
  INV_X1 U3846 ( .A(n6705), .ZN(n3760) );
  XNOR2_X1 U3847 ( .A(n4167), .B(n4159), .ZN(n4301) );
  NAND2_X1 U3848 ( .A1(n5082), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4713) );
  NAND2_X1 U3849 ( .A1(n4103), .A2(n4147), .ZN(n4294) );
  INV_X1 U3850 ( .A(n7289), .ZN(n3742) );
  INV_X1 U3851 ( .A(n5051), .ZN(n4931) );
  NAND2_X1 U3852 ( .A1(n3746), .A2(n3672), .ZN(n6522) );
  NAND2_X1 U3853 ( .A1(n4187), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4178) );
  NAND2_X1 U3854 ( .A1(n4175), .A2(n3733), .ZN(n3732) );
  AND2_X1 U3855 ( .A1(n6951), .A2(n4187), .ZN(n3733) );
  NAND2_X1 U3856 ( .A1(n4176), .A2(n3734), .ZN(n3731) );
  AND2_X1 U3857 ( .A1(n6951), .A2(n3778), .ZN(n3734) );
  NAND2_X1 U3858 ( .A1(n3740), .A2(n3679), .ZN(n3697) );
  AOI22_X1 U3859 ( .A1(n4201), .A2(n4200), .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n5481), .ZN(n4197) );
  XNOR2_X1 U3860 ( .A(n6573), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4196)
         );
  INV_X1 U3861 ( .A(n4231), .ZN(n4203) );
  NOR2_X1 U3862 ( .A1(n7130), .A2(n4192), .ZN(n4193) );
  OR2_X1 U3863 ( .A1(n4146), .A2(n4145), .ZN(n4161) );
  OR2_X1 U3864 ( .A1(n4124), .A2(n4123), .ZN(n4135) );
  NAND2_X1 U3865 ( .A1(n3967), .A2(n5094), .ZN(n3929) );
  NAND2_X1 U3866 ( .A1(n3927), .A2(n5140), .ZN(n3930) );
  NOR2_X1 U3867 ( .A1(n3922), .A2(n4236), .ZN(n3931) );
  AND2_X1 U3868 ( .A1(n3866), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3796) );
  INV_X1 U3869 ( .A(n7311), .ZN(n7131) );
  AND2_X1 U3870 ( .A1(n3768), .A2(n6626), .ZN(n3767) );
  INV_X1 U3871 ( .A(n3769), .ZN(n3768) );
  INV_X1 U3872 ( .A(n6716), .ZN(n3761) );
  AND2_X1 U3873 ( .A1(n4428), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4433)
         );
  NOR2_X1 U3874 ( .A1(n6742), .A2(n3758), .ZN(n3757) );
  INV_X1 U3875 ( .A(n6500), .ZN(n3758) );
  NAND2_X1 U3876 ( .A1(n3754), .A2(n4333), .ZN(n3753) );
  INV_X1 U3877 ( .A(n5810), .ZN(n3754) );
  NAND2_X1 U3878 ( .A1(n3683), .A2(n3747), .ZN(n3745) );
  OR2_X1 U3879 ( .A1(n3725), .A2(n6698), .ZN(n3724) );
  NAND2_X1 U3880 ( .A1(n5215), .A2(n3941), .ZN(n4871) );
  AND2_X1 U3881 ( .A1(n4151), .A2(n4101), .ZN(n3750) );
  INV_X1 U3882 ( .A(n5701), .ZN(n3714) );
  OAI22_X1 U3883 ( .A1(n4294), .A2(n4222), .B1(n4136), .B2(n4110), .ZN(n4112)
         );
  OR2_X1 U3884 ( .A1(n3994), .A2(n3993), .ZN(n4060) );
  NOR2_X1 U3885 ( .A1(n4236), .A2(n4239), .ZN(n4786) );
  INV_X1 U3886 ( .A(n4060), .ZN(n4028) );
  NAND2_X1 U3887 ( .A1(n3940), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U3888 ( .A1(n3855), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3819) );
  INV_X1 U3889 ( .A(n4054), .ZN(n6594) );
  CLKBUF_X1 U3890 ( .A(n4956), .Z(n4957) );
  NAND2_X1 U3891 ( .A1(n7320), .A2(n4961), .ZN(n7436) );
  AND3_X1 U3892 ( .A1(n7088), .A2(n7603), .A3(n7589), .ZN(n4961) );
  CLKBUF_X1 U3893 ( .A(n4768), .Z(n4769) );
  AND2_X1 U3894 ( .A1(n6593), .A2(n7581), .ZN(n7631) );
  XNOR2_X1 U3895 ( .A(n4247), .B(n4246), .ZN(n4966) );
  AND2_X1 U3896 ( .A1(n7584), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4748) );
  OR2_X1 U3897 ( .A1(n4696), .A2(n4695), .ZN(n4716) );
  OR2_X1 U3898 ( .A1(n6620), .A2(n4284), .ZN(n4694) );
  OR2_X1 U3899 ( .A1(n4636), .A2(n6845), .ZN(n4653) );
  OR2_X1 U3900 ( .A1(n4653), .A2(n6835), .ZN(n4674) );
  NAND2_X1 U3901 ( .A1(n6694), .A2(n3671), .ZN(n3759) );
  AND2_X1 U3902 ( .A1(n5597), .A2(n5598), .ZN(n4317) );
  INV_X1 U3903 ( .A(n5085), .ZN(n5075) );
  AND2_X1 U3904 ( .A1(n4937), .A2(n6532), .ZN(n3715) );
  NOR2_X1 U3905 ( .A1(n7056), .A2(n6878), .ZN(n7017) );
  OR2_X1 U3906 ( .A1(n6723), .A2(n6774), .ZN(n3719) );
  NOR2_X1 U3907 ( .A1(n3773), .A2(n4179), .ZN(n3739) );
  NAND2_X1 U3908 ( .A1(n7066), .A2(n7092), .ZN(n4177) );
  NAND2_X1 U3909 ( .A1(n3694), .A2(n3693), .ZN(n3699) );
  AOI21_X1 U3910 ( .B1(n3695), .B2(n3741), .A(n6465), .ZN(n3694) );
  NAND2_X1 U3911 ( .A1(n7288), .A2(n3695), .ZN(n3693) );
  NOR2_X1 U3912 ( .A1(n7288), .A2(n3741), .ZN(n3698) );
  OR2_X1 U3913 ( .A1(n4769), .A2(n6594), .ZN(n7554) );
  NAND2_X1 U3914 ( .A1(n4899), .A2(n6589), .ZN(n7079) );
  AND2_X1 U3915 ( .A1(n4786), .A2(n4885), .ZN(n6583) );
  INV_X1 U3916 ( .A(n4909), .ZN(n4899) );
  INV_X1 U3917 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5338) );
  INV_X1 U3918 ( .A(n5317), .ZN(n7132) );
  AND2_X1 U3919 ( .A1(n6593), .A2(n6583), .ZN(n7575) );
  INV_X1 U3920 ( .A(READY_N), .ZN(n7634) );
  INV_X1 U3921 ( .A(n7529), .ZN(n7519) );
  AND2_X1 U3922 ( .A1(n6829), .A2(n4256), .ZN(n7706) );
  OAI21_X1 U3923 ( .B1(n5091), .B2(n5090), .A(n7581), .ZN(n5092) );
  INV_X1 U3924 ( .A(n7302), .ZN(n7278) );
  NAND2_X1 U3925 ( .A1(n7283), .A2(n4997), .ZN(n7302) );
  INV_X1 U3926 ( .A(n4189), .ZN(n3730) );
  XNOR2_X1 U3927 ( .A(n4756), .B(n4940), .ZN(n4955) );
  AND2_X1 U3928 ( .A1(n4231), .A2(n4198), .ZN(n4218) );
  OAI22_X1 U3929 ( .A1(n4197), .A2(n4196), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6573), .ZN(n4195) );
  OAI22_X1 U3930 ( .A1(n4195), .A2(n4190), .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n7566), .ZN(n4191) );
  NOR2_X1 U3931 ( .A1(n6518), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4190)
         );
  INV_X1 U3932 ( .A(n4088), .ZN(n3728) );
  NAND2_X1 U3933 ( .A1(n3727), .A2(n4101), .ZN(n4147) );
  OR2_X1 U3934 ( .A1(n4098), .A2(n4097), .ZN(n4108) );
  NAND2_X1 U3935 ( .A1(n5140), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4029) );
  AND2_X1 U3936 ( .A1(n3915), .A2(n3914), .ZN(n3932) );
  NAND2_X1 U3937 ( .A1(n3909), .A2(n3904), .ZN(n3928) );
  NAND2_X1 U3938 ( .A1(n3943), .A2(n3942), .ZN(n4894) );
  NAND2_X1 U3939 ( .A1(n3923), .A2(n3928), .ZN(n3949) );
  NAND2_X1 U3940 ( .A1(n3789), .A2(n3788), .ZN(n3790) );
  AOI22_X1 U3941 ( .A1(n4367), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U3942 ( .A1(n3855), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3846) );
  OAI21_X1 U3943 ( .B1(n3967), .B2(n4226), .A(n4225), .ZN(n4227) );
  OR2_X1 U3944 ( .A1(n6857), .A2(n4284), .ZN(n4635) );
  NAND2_X1 U3945 ( .A1(n3770), .A2(n6637), .ZN(n3769) );
  AND2_X1 U3946 ( .A1(n4514), .A2(n3763), .ZN(n3762) );
  INV_X1 U3947 ( .A(n6718), .ZN(n3763) );
  INV_X1 U3948 ( .A(n4691), .ZN(n4744) );
  AND2_X1 U3949 ( .A1(n4442), .A2(n4409), .ZN(n4415) );
  INV_X1 U3950 ( .A(n4307), .ZN(n4308) );
  INV_X1 U3951 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4241) );
  NAND2_X1 U3952 ( .A1(n7066), .A2(n3686), .ZN(n3747) );
  OR2_X1 U3953 ( .A1(n4010), .A2(n4009), .ZN(n4165) );
  OR2_X1 U3954 ( .A1(n7066), .A2(n4183), .ZN(n4184) );
  OR2_X1 U3955 ( .A1(n6732), .A2(n3721), .ZN(n3720) );
  INV_X1 U3956 ( .A(n6784), .ZN(n3721) );
  INV_X1 U3957 ( .A(n4167), .ZN(n4155) );
  OR2_X1 U3958 ( .A1(n4049), .A2(n4048), .ZN(n4104) );
  OR2_X1 U3959 ( .A1(n3981), .A2(n3980), .ZN(n4082) );
  OR2_X1 U3960 ( .A1(n4020), .A2(n4019), .ZN(n4074) );
  AND2_X1 U3961 ( .A1(STATE2_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3936) );
  INV_X1 U3962 ( .A(n5121), .ZN(n5132) );
  AOI21_X1 U3963 ( .B1(n7586), .B2(n7596), .A(n7598), .ZN(n5121) );
  NAND2_X1 U3964 ( .A1(n4515), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4532)
         );
  OR2_X1 U3965 ( .A1(n5487), .A2(n4261), .ZN(n4262) );
  AND2_X1 U3966 ( .A1(n4832), .A2(n4831), .ZN(n6502) );
  AND2_X1 U3967 ( .A1(n4824), .A2(n4823), .ZN(n6451) );
  NAND2_X1 U3968 ( .A1(n5015), .A2(n5014), .ZN(n5091) );
  AND2_X1 U3969 ( .A1(n7631), .A2(n7133), .ZN(n7153) );
  AND2_X1 U3970 ( .A1(n3765), .A2(n3767), .ZN(n3764) );
  INV_X1 U3971 ( .A(n6527), .ZN(n3765) );
  NAND2_X1 U3972 ( .A1(n3766), .A2(n3767), .ZN(n6525) );
  NOR2_X1 U3973 ( .A1(n4596), .A2(n6671), .ZN(n4614) );
  AND2_X1 U3974 ( .A1(n4595), .A2(n4594), .ZN(n6876) );
  NAND2_X1 U3975 ( .A1(n4550), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4566)
         );
  NOR2_X1 U3976 ( .A1(n4532), .A2(n6897), .ZN(n4550) );
  NOR2_X1 U3977 ( .A1(n4493), .A2(n6720), .ZN(n4496) );
  AND2_X1 U3978 ( .A1(n4496), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4515)
         );
  NOR2_X1 U3979 ( .A1(n4449), .A2(n4243), .ZN(n4463) );
  NAND2_X1 U3980 ( .A1(n4463), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4493)
         );
  NAND2_X1 U3981 ( .A1(n4433), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4449)
         );
  NOR2_X1 U3982 ( .A1(n3756), .A2(n6731), .ZN(n3755) );
  INV_X1 U3983 ( .A(n3757), .ZN(n3756) );
  INV_X1 U3984 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4242) );
  NAND2_X1 U3985 ( .A1(n6501), .A2(n6500), .ZN(n6741) );
  NOR2_X1 U3986 ( .A1(n4366), .A2(n5858), .ZN(n4382) );
  INV_X1 U3987 ( .A(n4414), .ZN(n6447) );
  NAND2_X1 U3988 ( .A1(n4350), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4366)
         );
  CLKBUF_X1 U3989 ( .A(n5850), .Z(n5851) );
  OR2_X1 U3990 ( .A1(n3753), .A2(n3752), .ZN(n3751) );
  INV_X1 U3991 ( .A(n5832), .ZN(n3752) );
  OR2_X1 U3992 ( .A1(n4328), .A2(n5798), .ZN(n4334) );
  NOR2_X1 U3993 ( .A1(n5147), .A2(n3753), .ZN(n5833) );
  AND4_X1 U3994 ( .A1(n4332), .A2(n4331), .A3(n4330), .A4(n4329), .ZN(n5148)
         );
  INV_X1 U3995 ( .A(n4305), .ZN(n4306) );
  NAND2_X1 U3996 ( .A1(n4296), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4309)
         );
  NOR2_X1 U3997 ( .A1(n4309), .A2(n7479), .ZN(n4310) );
  CLKBUF_X1 U3998 ( .A(n5007), .Z(n5008) );
  OR2_X1 U3999 ( .A1(n5098), .A2(n5099), .ZN(n4276) );
  NAND2_X1 U4000 ( .A1(n6851), .A2(n6855), .ZN(n6843) );
  INV_X1 U4001 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6842) );
  NOR3_X1 U4002 ( .A1(n6709), .A2(n3724), .A3(n3726), .ZN(n6677) );
  AND2_X1 U4003 ( .A1(n4171), .A2(n3687), .ZN(n6866) );
  AND2_X1 U4004 ( .A1(n4853), .A2(n4852), .ZN(n6686) );
  NOR2_X1 U4005 ( .A1(n6709), .A2(n3724), .ZN(n7014) );
  AND2_X1 U4006 ( .A1(n7066), .A2(n7023), .ZN(n6863) );
  NOR2_X1 U4007 ( .A1(n6747), .A2(n6732), .ZN(n6785) );
  AND2_X1 U4008 ( .A1(n4836), .A2(n4835), .ZN(n6744) );
  INV_X1 U4009 ( .A(n5150), .ZN(n3713) );
  NAND2_X1 U4010 ( .A1(n5654), .A2(n3677), .ZN(n5704) );
  NAND2_X1 U4011 ( .A1(n5654), .A2(n5154), .ZN(n5702) );
  NOR2_X1 U4012 ( .A1(n3711), .A2(n5720), .ZN(n3709) );
  OR2_X1 U4013 ( .A1(n4027), .A2(n4028), .ZN(n3995) );
  INV_X1 U4014 ( .A(n5043), .ZN(n5034) );
  AND2_X1 U4015 ( .A1(n4770), .A2(n4886), .ZN(n5317) );
  NAND2_X1 U4016 ( .A1(n4039), .A2(n4038), .ZN(n5330) );
  AND2_X1 U4017 ( .A1(n5480), .A2(n5617), .ZN(n5489) );
  NOR2_X1 U4018 ( .A1(n5259), .A2(n5258), .ZN(n5339) );
  NAND2_X1 U4019 ( .A1(n7318), .A2(n5132), .ZN(n5399) );
  NOR2_X1 U4020 ( .A1(n5193), .A2(n4255), .ZN(n5340) );
  INV_X1 U4021 ( .A(n5747), .ZN(n5668) );
  NOR2_X1 U4022 ( .A1(n5193), .A2(n5258), .ZN(n5404) );
  NAND2_X1 U4023 ( .A1(n7584), .A2(n5044), .ZN(n5870) );
  AOI21_X1 U4024 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n3937), .A(n5399), .ZN(
        n5873) );
  INV_X1 U4025 ( .A(n6593), .ZN(n5026) );
  AND2_X1 U4026 ( .A1(n5338), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4240) );
  INV_X1 U4027 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6361) );
  AND2_X1 U4028 ( .A1(n7632), .A2(n4990), .ZN(n7320) );
  INV_X1 U4029 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n7318) );
  INV_X1 U4030 ( .A(n7514), .ZN(n7487) );
  AND2_X1 U4031 ( .A1(n7436), .A2(STATE2_REG_3__SCAN_IN), .ZN(n7501) );
  OR2_X1 U4032 ( .A1(n6597), .A2(n4980), .ZN(n7529) );
  OR2_X1 U4033 ( .A1(n6597), .A2(n4970), .ZN(n7457) );
  INV_X1 U4034 ( .A(n7501), .ZN(n7531) );
  INV_X1 U4035 ( .A(n7256), .ZN(n6793) );
  NAND2_X2 U4036 ( .A1(n7259), .A2(n4237), .ZN(n7256) );
  INV_X1 U4037 ( .A(n6831), .ZN(n7707) );
  AND2_X1 U4038 ( .A1(n6829), .A2(n6576), .ZN(n7710) );
  NAND2_X2 U4039 ( .A1(n6829), .A2(n5095), .ZN(n6831) );
  NAND2_X1 U4040 ( .A1(n6829), .A2(n5096), .ZN(n6833) );
  NOR2_X1 U4041 ( .A1(n7580), .A2(n7153), .ZN(n7164) );
  INV_X1 U4042 ( .A(n7632), .ZN(n7633) );
  AND2_X2 U4043 ( .A1(n7631), .A2(n5087), .ZN(n7692) );
  CLKBUF_X1 U4044 ( .A(n7666), .Z(n7691) );
  AND2_X1 U4045 ( .A1(n4674), .A2(n4654), .ZN(n6837) );
  INV_X1 U4046 ( .A(n6700), .ZN(n6899) );
  INV_X1 U4047 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6897) );
  XNOR2_X1 U4048 ( .A(n3716), .B(n4938), .ZN(n6755) );
  OR2_X1 U4049 ( .A1(n4936), .A2(n3717), .ZN(n3716) );
  AND2_X1 U4050 ( .A1(n6533), .A2(n3715), .ZN(n3717) );
  INV_X1 U4051 ( .A(n6542), .ZN(n6545) );
  AND2_X1 U4052 ( .A1(n6996), .A2(n4925), .ZN(n6549) );
  OAI21_X1 U4053 ( .B1(n6834), .B2(n6842), .A(n6523), .ZN(n6524) );
  AND2_X1 U4054 ( .A1(n7017), .A2(n4924), .ZN(n6996) );
  NAND2_X1 U4055 ( .A1(n4181), .A2(n3739), .ZN(n3736) );
  AND2_X1 U4056 ( .A1(n3732), .A2(n3731), .ZN(n6944) );
  OR2_X1 U4057 ( .A1(n7079), .A2(n7077), .ZN(n4904) );
  OR2_X1 U4058 ( .A1(n7081), .A2(n7080), .ZN(n7396) );
  NOR2_X1 U4059 ( .A1(n3698), .A2(n3697), .ZN(n6466) );
  NAND2_X1 U4060 ( .A1(n3696), .A2(n3740), .ZN(n6423) );
  NOR2_X1 U4061 ( .A1(n3744), .A2(n3676), .ZN(n6424) );
  NAND2_X1 U4062 ( .A1(n4899), .A2(n4882), .ZN(n7090) );
  AOI221_X1 U4063 ( .B1(n7353), .B2(n7079), .C1(n5820), .C2(n7079), .A(n5818), 
        .ZN(n6472) );
  AND2_X1 U4064 ( .A1(n3710), .A2(n3712), .ZN(n5116) );
  OR2_X1 U4065 ( .A1(n3692), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n7261)
         );
  NAND2_X1 U4066 ( .A1(n4899), .A2(n4789), .ZN(n7350) );
  INV_X1 U4067 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5481) );
  INV_X1 U4068 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5049) );
  INV_X1 U4069 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n5044) );
  INV_X1 U4070 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3785) );
  INV_X1 U4071 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n6573) );
  INV_X1 U4072 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n6518) );
  NOR2_X1 U4073 ( .A1(n7593), .A2(n7549), .ZN(n6572) );
  INV_X1 U4074 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n7551) );
  NOR2_X1 U4075 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n7548) );
  INV_X1 U4076 ( .A(n6572), .ZN(n7552) );
  OR2_X1 U4077 ( .A1(n5499), .A2(n5804), .ZN(n5899) );
  INV_X1 U4078 ( .A(n6420), .ZN(n6019) );
  OAI21_X1 U4079 ( .B1(n5567), .B2(n5566), .A(n5565), .ZN(n5589) );
  INV_X1 U4080 ( .A(n5964), .ZN(n5748) );
  INV_X1 U4081 ( .A(n5971), .ZN(n5772) );
  INV_X1 U4082 ( .A(n5979), .ZN(n5753) );
  INV_X1 U4083 ( .A(n5957), .ZN(n5764) );
  NAND2_X1 U4084 ( .A1(n5618), .A2(n5128), .ZN(n5590) );
  NOR2_X1 U4085 ( .A1(n5399), .A2(n5602), .ZN(n6416) );
  NOR2_X1 U4086 ( .A1(n5399), .A2(n5230), .ZN(n5971) );
  INV_X1 U4087 ( .A(n5776), .ZN(n5973) );
  NOR2_X1 U4088 ( .A1(n5399), .A2(n6250), .ZN(n5979) );
  INV_X1 U4089 ( .A(n5755), .ZN(n5983) );
  NOR2_X1 U4090 ( .A1(n5399), .A2(n5217), .ZN(n5957) );
  INV_X1 U4091 ( .A(n5766), .ZN(n5959) );
  NAND2_X1 U4092 ( .A1(n5340), .A2(n5804), .ZN(n5918) );
  NOR2_X1 U4093 ( .A1(n5229), .A2(n5228), .ZN(n5776) );
  INV_X1 U4094 ( .A(n5759), .ZN(n6005) );
  NAND2_X1 U4095 ( .A1(n5260), .A2(DATAI_5_), .ZN(n5997) );
  INV_X1 U4096 ( .A(n5789), .ZN(n5991) );
  NAND2_X1 U4097 ( .A1(n5260), .A2(DATAI_6_), .ZN(n6004) );
  INV_X1 U4098 ( .A(n5780), .ZN(n5998) );
  NAND2_X1 U4099 ( .A1(n5404), .A2(n5804), .ZN(n5603) );
  INV_X1 U4100 ( .A(n6413), .ZN(n6014) );
  NOR2_X1 U4101 ( .A1(n5026), .A2(n5044), .ZN(n7598) );
  NAND2_X1 U4102 ( .A1(n4240), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7605) );
  INV_X1 U4103 ( .A(STATE_REG_0__SCAN_IN), .ZN(n7619) );
  NOR2_X1 U4104 ( .A1(n7709), .A2(n4237), .ZN(n6796) );
  OAI21_X1 U4105 ( .B1(n4949), .B2(n7543), .A(n3670), .ZN(U2955) );
  INV_X1 U4106 ( .A(n4253), .ZN(n3729) );
  OAI211_X1 U4107 ( .C1(n4955), .C2(n7543), .A(n3748), .B(n4954), .ZN(U2956)
         );
  AND2_X2 U4108 ( .A1(n5039), .A2(n5307), .ZN(n4655) );
  INV_X1 U4109 ( .A(n4171), .ZN(n4187) );
  AND2_X1 U4110 ( .A1(n3761), .A2(n3671), .ZN(n3667) );
  NAND2_X1 U4111 ( .A1(n6501), .A2(n3757), .ZN(n6729) );
  OR2_X1 U4112 ( .A1(n6747), .A2(n3720), .ZN(n3668) );
  NAND2_X1 U4113 ( .A1(n3761), .A2(n3762), .ZN(n6704) );
  AND2_X1 U4114 ( .A1(n3736), .A2(n3682), .ZN(n3669) );
  INV_X1 U4115 ( .A(n3682), .ZN(n3738) );
  AND2_X1 U4116 ( .A1(n4753), .A2(n3729), .ZN(n3670) );
  NAND2_X1 U4117 ( .A1(n3728), .A2(n5158), .ZN(n4102) );
  INV_X1 U4118 ( .A(n4102), .ZN(n3727) );
  OR2_X2 U4119 ( .A1(n3861), .A2(n3860), .ZN(n3945) );
  INV_X1 U4120 ( .A(n3945), .ZN(n3906) );
  AND2_X1 U4121 ( .A1(n3762), .A2(n3760), .ZN(n3671) );
  NAND2_X1 U4122 ( .A1(n5600), .A2(n4333), .ZN(n5146) );
  AND2_X1 U4123 ( .A1(n3685), .A2(n3745), .ZN(n3672) );
  AND2_X1 U4124 ( .A1(n6532), .A2(n4877), .ZN(n3673) );
  AND2_X2 U4125 ( .A1(n5228), .A2(n3941), .ZN(n4054) );
  OR2_X1 U4126 ( .A1(n7066), .A2(n6519), .ZN(n3674) );
  OR3_X1 U4127 ( .A1(n6747), .A2(n3720), .A3(n3719), .ZN(n3675) );
  OR2_X1 U4128 ( .A1(n3849), .A2(n3848), .ZN(n3923) );
  NOR2_X1 U4129 ( .A1(n6716), .A2(n6718), .ZN(n6717) );
  AND2_X1 U4130 ( .A1(n4164), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3676)
         );
  AND2_X1 U4131 ( .A1(n5154), .A2(n3714), .ZN(n3677) );
  NAND2_X1 U4132 ( .A1(n6862), .A2(n7052), .ZN(n7051) );
  NAND4_X1 U4133 ( .A1(n3931), .A2(n3953), .A3(n3930), .A4(n3929), .ZN(n3956)
         );
  OAI21_X1 U4134 ( .B1(n3984), .B2(n3983), .A(n3955), .ZN(n3963) );
  NAND2_X1 U4135 ( .A1(n4187), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3678)
         );
  INV_X1 U4136 ( .A(n6519), .ZN(n6851) );
  NAND2_X1 U4137 ( .A1(n4170), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3679)
         );
  INV_X1 U4138 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5042) );
  AND2_X1 U4139 ( .A1(n3677), .A2(n3713), .ZN(n3680) );
  AND2_X1 U4140 ( .A1(n3707), .A2(n3674), .ZN(n3681) );
  INV_X1 U4141 ( .A(n4237), .ZN(n5082) );
  NAND2_X1 U4142 ( .A1(n3921), .A2(n3906), .ZN(n4236) );
  NAND2_X1 U4143 ( .A1(n4187), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3682) );
  AND2_X1 U4144 ( .A1(n4187), .A2(n3777), .ZN(n3683) );
  NAND2_X1 U4145 ( .A1(n4181), .A2(n4180), .ZN(n6927) );
  NAND2_X1 U4146 ( .A1(n5140), .A2(n3924), .ZN(n4884) );
  OAI21_X1 U4147 ( .B1(n4025), .B2(n4100), .A(n4099), .ZN(n4101) );
  INV_X1 U4148 ( .A(n4101), .ZN(n3749) );
  INV_X1 U4149 ( .A(n3718), .ZN(n6775) );
  NOR3_X1 U4150 ( .A1(n6747), .A2(n3720), .A3(n6723), .ZN(n3718) );
  NOR2_X1 U4151 ( .A1(n7288), .A2(n7289), .ZN(n3744) );
  INV_X1 U4152 ( .A(n4179), .ZN(n4180) );
  NOR2_X1 U4153 ( .A1(n4187), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4179)
         );
  NAND2_X1 U4154 ( .A1(n7066), .A2(n7408), .ZN(n3684) );
  AOI21_X1 U4155 ( .B1(n7278), .B2(n4967), .A(n4953), .ZN(n4954) );
  OAI21_X1 U4156 ( .B1(n3739), .B2(n3738), .A(n3684), .ZN(n3737) );
  NAND2_X1 U4157 ( .A1(n5839), .A2(n5838), .ZN(n5837) );
  NOR2_X2 U4158 ( .A1(n3901), .A2(n7584), .ZN(n4442) );
  INV_X1 U4159 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5798) );
  INV_X1 U4160 ( .A(n6650), .ZN(n3770) );
  NAND2_X1 U4161 ( .A1(n3692), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n7260)
         );
  NAND2_X1 U4162 ( .A1(n7575), .A2(n7581), .ZN(n7543) );
  INV_X1 U4163 ( .A(n7543), .ZN(n7298) );
  AND2_X1 U4164 ( .A1(n6853), .A2(n4186), .ZN(n3685) );
  INV_X1 U4165 ( .A(n3708), .ZN(n5327) );
  INV_X1 U4166 ( .A(n3712), .ZN(n3711) );
  OR2_X1 U4167 ( .A1(n6878), .A2(n4920), .ZN(n3686) );
  AND2_X1 U4168 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3687) );
  NAND3_X1 U4169 ( .A1(n3925), .A2(n3908), .A3(n3949), .ZN(n3688) );
  NAND3_X1 U4170 ( .A1(n3907), .A2(n3949), .A3(n3906), .ZN(n3689) );
  OAI21_X1 U4171 ( .B1(n3692), .B2(n3691), .A(n3690), .ZN(n4086) );
  NAND2_X1 U4172 ( .A1(n7263), .A2(n4078), .ZN(n3690) );
  NOR2_X1 U4173 ( .A1(n7263), .A2(n4078), .ZN(n3691) );
  NAND2_X1 U4174 ( .A1(n4064), .A2(n4063), .ZN(n3692) );
  INV_X1 U4175 ( .A(n3698), .ZN(n3696) );
  INV_X1 U4176 ( .A(n3699), .ZN(n6464) );
  AND2_X2 U4177 ( .A1(n3699), .A2(n3678), .ZN(n6970) );
  NAND3_X1 U4178 ( .A1(n3732), .A2(n3731), .A3(n6943), .ZN(n6942) );
  AND2_X2 U4179 ( .A1(n3901), .A2(n4237), .ZN(n4256) );
  NAND2_X1 U4180 ( .A1(n3827), .A2(n3826), .ZN(n3701) );
  NAND2_X1 U4181 ( .A1(n3829), .A2(n3828), .ZN(n3702) );
  AND2_X2 U4182 ( .A1(n3704), .A2(n3703), .ZN(n5066) );
  NAND2_X1 U4183 ( .A1(n5003), .A2(n5004), .ZN(n3703) );
  NAND2_X1 U4184 ( .A1(n3705), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n5003)
         );
  OR2_X1 U4185 ( .A1(n3705), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3704)
         );
  AOI21_X1 U4186 ( .B1(n7268), .B2(n7269), .A(n4087), .ZN(n3705) );
  AND2_X4 U4187 ( .A1(n3708), .A2(n5307), .ZN(n3864) );
  AND2_X2 U4188 ( .A1(n5308), .A2(n3708), .ZN(n3974) );
  AND2_X2 U4189 ( .A1(n3708), .A2(n3804), .ZN(n4118) );
  AND2_X2 U4190 ( .A1(n3708), .A2(n6513), .ZN(n3865) );
  XNOR2_X1 U4191 ( .A(n4794), .B(n5050), .ZN(n5083) );
  NAND3_X1 U4192 ( .A1(n3710), .A2(n5115), .A3(n3712), .ZN(n5114) );
  NAND3_X1 U4193 ( .A1(n3710), .A2(n3709), .A3(n5115), .ZN(n5722) );
  INV_X1 U4194 ( .A(n4794), .ZN(n3712) );
  AND2_X1 U4195 ( .A1(n6533), .A2(n6532), .ZN(n6546) );
  AOI21_X1 U4196 ( .B1(n6533), .B2(n3673), .A(n4932), .ZN(n4936) );
  INV_X1 U4197 ( .A(n3722), .ZN(n6638) );
  NOR2_X1 U4198 ( .A1(n6709), .A2(n6698), .ZN(n6697) );
  INV_X1 U4199 ( .A(n6686), .ZN(n3725) );
  INV_X1 U4200 ( .A(n4861), .ZN(n3726) );
  INV_X1 U4201 ( .A(n4181), .ZN(n3735) );
  AOI21_X2 U4202 ( .B1(n3735), .B2(n3682), .A(n3737), .ZN(n6911) );
  NAND2_X1 U4203 ( .A1(n6861), .A2(n3747), .ZN(n3746) );
  NOR2_X4 U4204 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5307) );
  NOR2_X1 U4205 ( .A1(n6651), .A2(n6650), .ZN(n6635) );
  NAND2_X2 U4206 ( .A1(n3766), .A2(n3764), .ZN(n6558) );
  INV_X2 U4207 ( .A(n6651), .ZN(n3766) );
  AOI21_X2 U4208 ( .B1(n6865), .B2(n6864), .A(n6863), .ZN(n6896) );
  INV_X1 U4209 ( .A(n7051), .ZN(n6865) );
  NAND2_X1 U4210 ( .A1(n6797), .A2(n6796), .ZN(n6799) );
  NAND2_X1 U4211 ( .A1(n6797), .A2(n7297), .ZN(n4753) );
  INV_X1 U4212 ( .A(n6521), .ZN(n6541) );
  NAND2_X1 U4213 ( .A1(n6682), .A2(n6876), .ZN(n6665) );
  INV_X1 U4214 ( .A(n6665), .ZN(n4613) );
  NAND2_X1 U4215 ( .A1(n3935), .A2(n3955), .ZN(n3984) );
  NAND2_X1 U4216 ( .A1(n5124), .A2(n7318), .ZN(n4051) );
  NOR2_X2 U4217 ( .A1(n6519), .A2(n6988), .ZN(n6521) );
  NAND2_X1 U4218 ( .A1(n5404), .A2(n5487), .ZN(n5786) );
  NAND2_X1 U4219 ( .A1(n5340), .A2(n5487), .ZN(n5894) );
  OR2_X1 U4220 ( .A1(n5499), .A2(n5487), .ZN(n5926) );
  INV_X1 U4221 ( .A(n5487), .ZN(n5804) );
  NAND2_X1 U4222 ( .A1(n3956), .A2(n3936), .ZN(n3939) );
  OR2_X1 U4223 ( .A1(n6579), .A2(n7535), .ZN(n3771) );
  AND3_X1 U4224 ( .A1(n4174), .A2(n4173), .A3(n4172), .ZN(n3772) );
  AND2_X1 U4225 ( .A1(n7066), .A2(n7401), .ZN(n3773) );
  AND2_X1 U4226 ( .A1(n3775), .A2(n4031), .ZN(n3774) );
  OR2_X1 U4227 ( .A1(n4025), .A2(n4026), .ZN(n3775) );
  AND4_X1 U4228 ( .A1(n3825), .A2(n3824), .A3(n3823), .A4(n3822), .ZN(n3776)
         );
  INV_X2 U4229 ( .A(n7627), .ZN(n7309) );
  NAND2_X1 U4230 ( .A1(n5093), .A2(n5092), .ZN(n6829) );
  INV_X1 U4231 ( .A(n6829), .ZN(n7709) );
  NAND2_X1 U4232 ( .A1(n4185), .A2(n6867), .ZN(n3777) );
  AND2_X1 U4233 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3778) );
  OR2_X1 U4234 ( .A1(n7541), .A2(n4968), .ZN(n3779) );
  INV_X1 U4235 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4565) );
  INV_X1 U4236 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4243) );
  AND2_X2 U4237 ( .A1(n5078), .A2(n7581), .ZN(n7259) );
  INV_X1 U4238 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n7130) );
  INV_X1 U4239 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4111) );
  AND2_X1 U4240 ( .A1(n3857), .A2(n3856), .ZN(n3780) );
  OR2_X1 U4241 ( .A1(n6581), .A2(n7537), .ZN(n3781) );
  OR2_X1 U4242 ( .A1(n3916), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3782)
         );
  INV_X1 U4243 ( .A(n3879), .ZN(n3969) );
  INV_X1 U4244 ( .A(n3925), .ZN(n4773) );
  INV_X1 U4245 ( .A(n4205), .ZN(n4200) );
  NOR2_X1 U4246 ( .A1(n5088), .A2(n4199), .ZN(n4223) );
  INV_X1 U4247 ( .A(n3948), .ZN(n3921) );
  NAND3_X1 U4248 ( .A1(n4887), .A2(n3902), .A3(n5088), .ZN(n4784) );
  INV_X1 U4249 ( .A(n4759), .ZN(n4226) );
  OAI21_X1 U4250 ( .B1(n4713), .B2(n4304), .A(n4303), .ZN(n4305) );
  AND3_X1 U4251 ( .A1(n4892), .A2(n4891), .A3(n4890), .ZN(n4893) );
  AOI21_X1 U4252 ( .B1(n4232), .B2(n4203), .A(n4760), .ZN(n4228) );
  INV_X1 U4253 ( .A(n4674), .ZN(n4244) );
  INV_X1 U4254 ( .A(n6771), .ZN(n4514) );
  NAND2_X1 U4255 ( .A1(n5034), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4691) );
  NAND2_X1 U4256 ( .A1(n4382), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4410)
         );
  NAND2_X1 U4257 ( .A1(n4127), .A2(n4150), .ZN(n4154) );
  INV_X1 U4258 ( .A(n3997), .ZN(n3999) );
  OR2_X1 U4259 ( .A1(n5094), .A2(n4238), .ZN(n5043) );
  INV_X1 U4260 ( .A(n4071), .ZN(n4024) );
  INV_X1 U4261 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3937) );
  AND2_X1 U4262 ( .A1(n4894), .A2(n4893), .ZN(n5032) );
  NOR2_X1 U4263 ( .A1(n4278), .A2(n4241), .ZN(n4279) );
  AND2_X1 U4264 ( .A1(n4830), .A2(n4829), .ZN(n6483) );
  INV_X1 U4265 ( .A(n6667), .ZN(n4612) );
  OR2_X1 U4266 ( .A1(n4783), .A2(n5013), .ZN(n5014) );
  NAND2_X1 U4267 ( .A1(n4244), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4696)
         );
  OR2_X1 U4268 ( .A1(n7542), .A2(n4284), .ZN(n4595) );
  INV_X1 U4269 ( .A(n6717), .ZN(n6772) );
  NOR2_X1 U4270 ( .A1(n4410), .A2(n4242), .ZN(n4428) );
  NOR2_X1 U4271 ( .A1(n4334), .A2(n5826), .ZN(n4350) );
  INV_X1 U4272 ( .A(n5148), .ZN(n4333) );
  INV_X1 U4273 ( .A(n6548), .ZN(n6540) );
  OR2_X1 U4274 ( .A1(n4915), .A2(n4914), .ZN(n7053) );
  NAND2_X1 U4275 ( .A1(n4133), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4134)
         );
  INV_X1 U4276 ( .A(n4255), .ZN(n5258) );
  AND2_X1 U4277 ( .A1(n5395), .A2(n3958), .ZN(n5134) );
  INV_X1 U4278 ( .A(n5614), .ZN(n5501) );
  INV_X1 U4279 ( .A(n5229), .ZN(n5182) );
  AND2_X1 U4280 ( .A1(n5032), .A2(n4898), .ZN(n6589) );
  INV_X1 U4281 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6671) );
  INV_X1 U4282 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6720) );
  INV_X1 U4283 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5858) );
  INV_X1 U4284 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5826) );
  AND2_X1 U4285 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n4279), .ZN(n4296)
         );
  NAND2_X1 U4286 ( .A1(n7436), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6597) );
  NAND2_X1 U4287 ( .A1(n4614), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4636)
         );
  INV_X1 U4288 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n7479) );
  OR2_X1 U4289 ( .A1(n6522), .A2(n4171), .ZN(n6523) );
  INV_X1 U4290 ( .A(n7370), .ZN(n7088) );
  INV_X1 U4291 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3786) );
  AND2_X1 U4292 ( .A1(n5168), .A2(n5167), .ZN(n5351) );
  NAND2_X1 U4293 ( .A1(n5339), .A2(n5804), .ZN(n5950) );
  NAND2_X1 U4294 ( .A1(n5339), .A2(n5487), .ZN(n6411) );
  NOR2_X1 U4295 ( .A1(n5126), .A2(n4255), .ZN(n5480) );
  AND2_X1 U4296 ( .A1(n3913), .A2(n3957), .ZN(n5281) );
  NAND2_X1 U4297 ( .A1(n5132), .A2(n7593), .ZN(n5229) );
  INV_X1 U4298 ( .A(n4267), .ZN(n4284) );
  INV_X1 U4299 ( .A(n4957), .ZN(n6582) );
  OR2_X1 U4300 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n7586), .ZN(n7322) );
  OR2_X1 U4301 ( .A1(n4566), .A2(n4565), .ZN(n4596) );
  NOR2_X1 U4302 ( .A1(n5870), .A2(STATE2_REG_1__SCAN_IN), .ZN(n7305) );
  INV_X1 U4303 ( .A(n7537), .ZN(n7522) );
  INV_X1 U4304 ( .A(n7457), .ZN(n7468) );
  AND2_X1 U4305 ( .A1(n4963), .A2(n4962), .ZN(n7521) );
  AND2_X1 U4306 ( .A1(n7259), .A2(n5082), .ZN(n6780) );
  INV_X1 U4307 ( .A(n7692), .ZN(n5093) );
  OAI21_X1 U4308 ( .B1(n4054), .B2(n7634), .A(n7633), .ZN(n7666) );
  NAND2_X1 U4309 ( .A1(n4310), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4328)
         );
  INV_X1 U4310 ( .A(n7605), .ZN(n7581) );
  INV_X1 U4311 ( .A(n7283), .ZN(n7296) );
  INV_X1 U4312 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n7401) );
  XNOR2_X1 U4313 ( .A(n4112), .B(n4111), .ZN(n5065) );
  INV_X1 U4314 ( .A(n7350), .ZN(n7419) );
  INV_X1 U4315 ( .A(n7090), .ZN(n7418) );
  OAI21_X1 U4316 ( .B1(n5742), .B2(n5741), .A(n5740), .ZN(n5785) );
  OAI211_X1 U4317 ( .C1(n5663), .C2(n5664), .A(n5662), .B(n5661), .ZN(n5693)
         );
  AND2_X1 U4318 ( .A1(n5489), .A2(n5487), .ZN(n5657) );
  AND2_X1 U4319 ( .A1(n5618), .A2(n5617), .ZN(n5697) );
  INV_X1 U4320 ( .A(n5128), .ZN(n5617) );
  OAI21_X1 U4321 ( .B1(n5166), .B2(n5165), .A(n5164), .ZN(n5350) );
  INV_X1 U4322 ( .A(n5950), .ZN(n5376) );
  OAI21_X1 U4323 ( .B1(n5289), .B2(n5288), .A(n5287), .ZN(n5373) );
  OAI21_X1 U4324 ( .B1(n5264), .B2(n5263), .A(n5262), .ZN(n6409) );
  INV_X1 U4325 ( .A(n6016), .ZN(n5593) );
  NOR2_X1 U4326 ( .A1(n5399), .A2(n5141), .ZN(n5964) );
  OAI211_X1 U4327 ( .C1(n5875), .C2(n5442), .A(n5441), .B(n5873), .ZN(n5466)
         );
  AND2_X1 U4328 ( .A1(n5157), .A2(n5128), .ZN(n5465) );
  INV_X1 U4329 ( .A(n5894), .ZN(n5920) );
  NOR2_X1 U4330 ( .A1(n5229), .A2(n5140), .ZN(n5750) );
  OAI21_X1 U4331 ( .B1(n5196), .B2(n5195), .A(n5194), .ZN(n5214) );
  NOR2_X1 U4332 ( .A1(n5229), .A2(n5215), .ZN(n5766) );
  INV_X1 U4333 ( .A(n5399), .ZN(n5260) );
  INV_X2 U4334 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n7584) );
  AOI21_X1 U4335 ( .B1(n7583), .B2(n7630), .A(n7582), .ZN(n7597) );
  AND2_X1 U4336 ( .A1(n7616), .A2(n7619), .ZN(n7311) );
  NAND2_X1 U4337 ( .A1(n7631), .A2(n6582), .ZN(n7632) );
  INV_X1 U4338 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n7608) );
  OR2_X1 U4339 ( .A1(n4966), .A2(n4964), .ZN(n7537) );
  NAND2_X1 U4340 ( .A1(n4966), .A2(n4965), .ZN(n7541) );
  NAND2_X1 U4341 ( .A1(n7153), .A2(n3941), .ZN(n7171) );
  INV_X1 U4342 ( .A(n7153), .ZN(n7152) );
  NAND2_X2 U4343 ( .A1(n7631), .A2(n7630), .ZN(n7694) );
  NAND2_X1 U4344 ( .A1(n7543), .A2(n4249), .ZN(n7283) );
  OR2_X1 U4345 ( .A1(n7314), .A2(n5870), .ZN(n6976) );
  INV_X1 U4346 ( .A(n7383), .ZN(n7414) );
  INV_X1 U4347 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n7566) );
  NAND2_X1 U4348 ( .A1(n5489), .A2(n5804), .ZN(n5956) );
  INV_X1 U4349 ( .A(n5657), .ZN(n5989) );
  AOI22_X1 U4350 ( .A1(n5616), .A2(n5621), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5615), .ZN(n5649) );
  NAND2_X1 U4351 ( .A1(n5157), .A2(n5617), .ZN(n5643) );
  INV_X1 U4352 ( .A(n5923), .ZN(n5557) );
  OR2_X1 U4353 ( .A1(n5868), .A2(n5487), .ZN(n6420) );
  OR2_X1 U4354 ( .A1(n5868), .A2(n5804), .ZN(n6016) );
  AOI22_X1 U4355 ( .A1(n5562), .A2(n5567), .B1(n5743), .B2(n5561), .ZN(n5596)
         );
  INV_X1 U4356 ( .A(n5434), .ZN(n5469) );
  AND2_X1 U4357 ( .A1(n5131), .A2(n5130), .ZN(n5394) );
  INV_X1 U4358 ( .A(n5750), .ZN(n5966) );
  AND2_X1 U4359 ( .A1(n5192), .A2(n5191), .ZN(n5216) );
  NAND2_X1 U4360 ( .A1(n5260), .A2(DATAI_4_), .ZN(n6011) );
  INV_X1 U4361 ( .A(n6416), .ZN(n6021) );
  CLKBUF_X1 U4362 ( .A(n7230), .Z(n7219) );
  AND2_X4 U4363 ( .A1(n5042), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5027)
         );
  NAND2_X1 U4364 ( .A1(n3855), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3784) );
  NAND2_X1 U4365 ( .A1(n3974), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3783)
         );
  NAND2_X1 U4366 ( .A1(n3784), .A2(n3783), .ZN(n3791) );
  AND2_X2 U4367 ( .A1(n3786), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n6513)
         );
  NAND2_X1 U4368 ( .A1(n3850), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3789)
         );
  INV_X1 U4369 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3787) );
  AND2_X2 U4370 ( .A1(n3787), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3804)
         );
  AND2_X4 U4371 ( .A1(n5027), .A2(n3804), .ZN(n3871) );
  NAND2_X1 U4372 ( .A1(n3665), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3788) );
  NOR2_X1 U4373 ( .A1(n3791), .A2(n3790), .ZN(n3798) );
  NAND2_X1 U4374 ( .A1(n3968), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3794)
         );
  NAND2_X1 U4375 ( .A1(n4367), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3793) );
  AND2_X4 U4376 ( .A1(n5033), .A2(n3804), .ZN(n3879) );
  NAND2_X1 U4377 ( .A1(n3879), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3792) );
  NAND3_X1 U4378 ( .A1(n3794), .A2(n3793), .A3(n3792), .ZN(n3795) );
  NOR2_X1 U4379 ( .A1(n3796), .A2(n3795), .ZN(n3797) );
  NAND2_X1 U4380 ( .A1(n4655), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3803) );
  AND2_X4 U4381 ( .A1(n5307), .A2(n5033), .ZN(n3892) );
  NAND2_X1 U4382 ( .A1(n3892), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3802) );
  NAND2_X1 U4383 ( .A1(n3864), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3801) );
  NOR2_X2 U4384 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3799) );
  AND2_X2 U4385 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5310) );
  BUF_X4 U4386 ( .A(n4000), .Z(n4534) );
  NAND2_X1 U4387 ( .A1(n4534), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3800) );
  NAND2_X1 U4388 ( .A1(n3865), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3808) );
  NAND2_X1 U4389 ( .A1(n4702), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3807)
         );
  NAND2_X1 U4390 ( .A1(n4118), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3806) );
  AND2_X2 U4391 ( .A1(n5033), .A2(n5308), .ZN(n3975) );
  NAND2_X1 U4392 ( .A1(n3975), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3805)
         );
  NAND3_X2 U4393 ( .A1(n3811), .A2(n3810), .A3(n3809), .ZN(n3909) );
  AOI22_X1 U4394 ( .A1(n4655), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3815) );
  AOI22_X1 U4395 ( .A1(n4702), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3892), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3814) );
  AOI22_X1 U4396 ( .A1(n3865), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3813) );
  AOI22_X1 U4397 ( .A1(n3850), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3871), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4398 ( .A1(n4367), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4399 ( .A1(n4118), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4400 ( .A1(n3662), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3816) );
  AOI22_X1 U4401 ( .A1(n3866), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3663), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4402 ( .A1(n4367), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4403 ( .A1(n4655), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4404 ( .A1(n3892), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4405 ( .A1(n3665), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4406 ( .A1(n4702), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4407 ( .A1(n4118), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3865), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4408 ( .A1(n3850), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4409 ( .A1(n4655), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4410 ( .A1(n4367), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4411 ( .A1(n3866), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3968), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4412 ( .A1(n3892), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3830) );
  NAND4_X1 U4413 ( .A1(n3833), .A2(n3832), .A3(n3831), .A4(n3830), .ZN(n3839)
         );
  AOI22_X1 U4414 ( .A1(n3666), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4415 ( .A1(n3865), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4416 ( .A1(n3850), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4417 ( .A1(n4702), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3834) );
  NAND4_X1 U4418 ( .A1(n3837), .A2(n3836), .A3(n3835), .A4(n3834), .ZN(n3838)
         );
  AOI22_X1 U4419 ( .A1(n3892), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4420 ( .A1(n3850), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4421 ( .A1(n4655), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3840) );
  NAND4_X1 U4422 ( .A1(n3843), .A2(n3842), .A3(n3841), .A4(n3840), .ZN(n3849)
         );
  AOI22_X1 U4423 ( .A1(n3866), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3968), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4424 ( .A1(n3865), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4425 ( .A1(n4702), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3844) );
  NAND4_X1 U4426 ( .A1(n3847), .A2(n3846), .A3(n3845), .A4(n3844), .ZN(n3848)
         );
  INV_X1 U4427 ( .A(n3949), .ZN(n3863) );
  AOI22_X1 U4428 ( .A1(n3968), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3892), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4429 ( .A1(n4655), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3850), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3853) );
  AOI22_X1 U4430 ( .A1(n3865), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3852) );
  AOI22_X1 U4431 ( .A1(n3864), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3851) );
  NAND4_X1 U4432 ( .A1(n3854), .A2(n3853), .A3(n3852), .A4(n3851), .ZN(n3861)
         );
  AOI22_X1 U4433 ( .A1(n4728), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3855), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4434 ( .A1(n3665), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4702), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4435 ( .A1(n4118), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4436 ( .A1(n4367), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3856) );
  NAND3_X1 U4437 ( .A1(n3859), .A2(n3858), .A3(n3780), .ZN(n3860) );
  NOR2_X1 U4438 ( .A1(n3945), .A2(n3901), .ZN(n3862) );
  NAND3_X1 U4439 ( .A1(n3925), .A2(n3863), .A3(n3862), .ZN(n4768) );
  INV_X1 U4440 ( .A(n4768), .ZN(n3878) );
  BUF_X8 U4441 ( .A(n3864), .Z(n4720) );
  AOI22_X1 U4442 ( .A1(n4655), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4720), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4443 ( .A1(n3865), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3892), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3869) );
  AOI22_X1 U4444 ( .A1(n3866), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3968), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4445 ( .A1(n4367), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3867) );
  NAND4_X1 U4446 ( .A1(n3870), .A2(n3869), .A3(n3868), .A4(n3867), .ZN(n3877)
         );
  AOI22_X1 U4447 ( .A1(n4702), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4118), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4448 ( .A1(n3666), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3974), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4449 ( .A1(n3850), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4450 ( .A1(n3855), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3872) );
  NAND4_X1 U4451 ( .A1(n3875), .A2(n3874), .A3(n3873), .A4(n3872), .ZN(n3876)
         );
  OR2_X4 U4452 ( .A1(n3877), .A2(n3876), .ZN(n3941) );
  NAND2_X1 U4453 ( .A1(n3878), .A2(n3941), .ZN(n4956) );
  NAND2_X1 U4454 ( .A1(n3866), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3883)
         );
  NAND2_X1 U4455 ( .A1(n3663), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3882)
         );
  NAND2_X1 U4456 ( .A1(n4367), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3881) );
  NAND2_X1 U4457 ( .A1(n3879), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3880) );
  NAND2_X1 U4458 ( .A1(n3850), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3887)
         );
  NAND2_X1 U4459 ( .A1(n3666), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3886) );
  NAND2_X1 U4460 ( .A1(n3855), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3885) );
  NAND2_X1 U4461 ( .A1(n3974), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3884)
         );
  NAND2_X1 U4462 ( .A1(n4702), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3891)
         );
  NAND2_X1 U4463 ( .A1(n3865), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3890) );
  NAND2_X1 U4464 ( .A1(n4118), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3889) );
  NAND2_X1 U4465 ( .A1(n3975), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3888)
         );
  NAND2_X1 U4466 ( .A1(n4655), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3896) );
  NAND2_X1 U4467 ( .A1(n3892), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3895) );
  NAND2_X1 U4468 ( .A1(n3864), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3894) );
  NAND2_X1 U4469 ( .A1(n4534), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3893) );
  AND4_X2 U4470 ( .A1(n3896), .A2(n3895), .A3(n3894), .A4(n3893), .ZN(n3897)
         );
  NAND4_X4 U4471 ( .A1(n3900), .A2(n3899), .A3(n3898), .A4(n3897), .ZN(n3924)
         );
  XNOR2_X1 U4472 ( .A(n6361), .B(STATE_REG_2__SCAN_IN), .ZN(n7616) );
  INV_X1 U4473 ( .A(n3909), .ZN(n6575) );
  INV_X1 U4474 ( .A(n3905), .ZN(n3902) );
  INV_X1 U4475 ( .A(n3903), .ZN(n3911) );
  INV_X2 U4476 ( .A(n5177), .ZN(n3940) );
  OAI21_X1 U4477 ( .B1(n3940), .B2(n4261), .A(n3905), .ZN(n3907) );
  AND2_X1 U4478 ( .A1(n4885), .A2(n5140), .ZN(n4771) );
  AND2_X1 U4479 ( .A1(n5228), .A2(n4771), .ZN(n3910) );
  NAND2_X1 U4480 ( .A1(n3911), .A2(n4783), .ZN(n3912) );
  NAND2_X1 U4481 ( .A1(n3912), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3933) );
  INV_X1 U4482 ( .A(n3933), .ZN(n3917) );
  NAND2_X1 U4483 ( .A1(n7548), .A2(n7318), .ZN(n4248) );
  INV_X1 U4484 ( .A(n4248), .ZN(n4037) );
  NAND2_X1 U4485 ( .A1(n3937), .A2(n5481), .ZN(n3913) );
  NAND2_X1 U4486 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3957) );
  NAND2_X1 U4487 ( .A1(n4037), .A2(n5281), .ZN(n3915) );
  INV_X1 U4488 ( .A(n4240), .ZN(n3959) );
  NAND2_X1 U4489 ( .A1(n3959), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3914) );
  INV_X1 U4490 ( .A(n3932), .ZN(n3916) );
  NAND2_X1 U4491 ( .A1(n3917), .A2(n3782), .ZN(n3935) );
  OAI21_X1 U4492 ( .B1(n3918), .B2(n5172), .A(n4884), .ZN(n3922) );
  INV_X1 U4493 ( .A(n3919), .ZN(n3920) );
  OAI211_X1 U4494 ( .C1(n3928), .C2(n5177), .A(n3920), .B(n3923), .ZN(n3948)
         );
  AND2_X4 U4495 ( .A1(n3924), .A2(n3923), .ZN(n4874) );
  NAND2_X1 U4496 ( .A1(n4885), .A2(n4874), .ZN(n5030) );
  NAND2_X1 U4497 ( .A1(n4773), .A2(n4054), .ZN(n3926) );
  NAND2_X2 U4498 ( .A1(n4208), .A2(n5177), .ZN(n4025) );
  INV_X2 U4499 ( .A(n4025), .ZN(n3967) );
  NAND3_X1 U4500 ( .A1(n3956), .A2(STATE2_REG_0__SCAN_IN), .A3(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3934) );
  NAND3_X1 U4501 ( .A1(n3934), .A2(n3933), .A3(n3932), .ZN(n3955) );
  MUX2_X1 U4502 ( .A(n4240), .B(n4248), .S(n3937), .Z(n3938) );
  NAND2_X1 U4503 ( .A1(n3939), .A2(n3938), .ZN(n3998) );
  NAND2_X1 U4504 ( .A1(n4770), .A2(n5228), .ZN(n3943) );
  AOI21_X1 U4505 ( .B1(n4232), .B2(n3940), .A(n3941), .ZN(n3942) );
  INV_X1 U4506 ( .A(n4261), .ZN(n3944) );
  NAND2_X1 U4507 ( .A1(n4887), .A2(n3944), .ZN(n4895) );
  NAND2_X1 U4508 ( .A1(n7548), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7585) );
  AOI21_X1 U4509 ( .B1(n3941), .B2(n3945), .A(n7585), .ZN(n3946) );
  AND2_X1 U4510 ( .A1(n4895), .A2(n3946), .ZN(n3952) );
  AND2_X1 U4511 ( .A1(n5094), .A2(n5177), .ZN(n3947) );
  OAI21_X1 U4512 ( .B1(n3948), .B2(n3947), .A(n3924), .ZN(n3951) );
  NAND2_X1 U4513 ( .A1(n3949), .A2(n4054), .ZN(n3950) );
  NAND2_X1 U4514 ( .A1(n4894), .A2(n3954), .ZN(n3997) );
  INV_X1 U4515 ( .A(n3963), .ZN(n3962) );
  NAND2_X1 U4516 ( .A1(n4033), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3961) );
  INV_X1 U4517 ( .A(n3957), .ZN(n5612) );
  NAND2_X1 U4518 ( .A1(n5612), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5395) );
  INV_X1 U4519 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5718) );
  NAND2_X1 U4520 ( .A1(n3957), .A2(n5718), .ZN(n3958) );
  AOI22_X1 U4521 ( .A1(n5134), .A2(n4037), .B1(n3959), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3960) );
  NAND2_X1 U4522 ( .A1(n3961), .A2(n3960), .ZN(n3964) );
  INV_X1 U4523 ( .A(n3964), .ZN(n3965) );
  NAND2_X1 U4524 ( .A1(n3963), .A2(n3965), .ZN(n3966) );
  BUF_X4 U4525 ( .A(n3866), .Z(n4728) );
  AOI22_X1 U4526 ( .A1(n4728), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4527 ( .A1(n4727), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4528 ( .A1(n4721), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4720), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3971) );
  AOI22_X1 U4529 ( .A1(n3892), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3970) );
  NAND4_X1 U4530 ( .A1(n3973), .A2(n3972), .A3(n3971), .A4(n3970), .ZN(n3981)
         );
  AOI22_X1 U4531 ( .A1(n3665), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4532 ( .A1(n4732), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4533 ( .A1(n3660), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4534 ( .A1(n4702), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3976) );
  NAND4_X1 U4535 ( .A1(n3979), .A2(n3978), .A3(n3977), .A4(n3976), .ZN(n3980)
         );
  AOI22_X1 U4536 ( .A1(n3967), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4231), 
        .B2(n4082), .ZN(n3982) );
  OAI21_X2 U4537 ( .B1(n5125), .B2(STATE2_REG_0__SCAN_IN), .A(n3982), .ZN(
        n4079) );
  XNOR2_X1 U4538 ( .A(n3984), .B(n3983), .ZN(n5028) );
  NAND2_X1 U4539 ( .A1(n5028), .A2(n7318), .ZN(n3996) );
  AOI22_X1 U4540 ( .A1(n4728), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3988) );
  AOI22_X1 U4541 ( .A1(n4727), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3987) );
  AOI22_X1 U4542 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n3666), .B1(n3865), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3986) );
  AOI22_X1 U4543 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n4721), .B1(n4720), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3985) );
  NAND4_X1 U4544 ( .A1(n3988), .A2(n3987), .A3(n3986), .A4(n3985), .ZN(n3994)
         );
  AOI22_X1 U4545 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n3660), .B1(n4702), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U4546 ( .A1(n3879), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U4547 ( .A1(n3892), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3990) );
  AOI22_X1 U4548 ( .A1(n4118), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3989) );
  NAND4_X1 U4549 ( .A1(n3992), .A2(n3991), .A3(n3990), .A4(n3989), .ZN(n3993)
         );
  XNOR2_X2 U4550 ( .A(n3999), .B(n3998), .ZN(n4263) );
  INV_X1 U4551 ( .A(n4027), .ZN(n4023) );
  AOI22_X1 U4552 ( .A1(n4728), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4553 ( .A1(n4727), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U4554 ( .A1(n4721), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4720), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4555 ( .A1(n3892), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4001) );
  NAND4_X1 U4556 ( .A1(n4004), .A2(n4003), .A3(n4002), .A4(n4001), .ZN(n4010)
         );
  AOI22_X1 U4557 ( .A1(n3665), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4558 ( .A1(n4732), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U4559 ( .A1(n3850), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U4560 ( .A1(n4702), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4005) );
  NAND4_X1 U4561 ( .A1(n4008), .A2(n4007), .A3(n4006), .A4(n4005), .ZN(n4009)
         );
  INV_X1 U4562 ( .A(n4165), .ZN(n4021) );
  AOI22_X1 U4563 ( .A1(n4721), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U4564 ( .A1(n4727), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4702), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4565 ( .A1(n4720), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4566 ( .A1(n4719), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4011) );
  NAND4_X1 U4567 ( .A1(n4014), .A2(n4013), .A3(n4012), .A4(n4011), .ZN(n4020)
         );
  AOI22_X1 U4568 ( .A1(n3660), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U4569 ( .A1(n3666), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4732), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4570 ( .A1(n4728), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3892), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U4571 ( .A1(n3664), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4015) );
  NAND4_X1 U4572 ( .A1(n4018), .A2(n4017), .A3(n4016), .A4(n4015), .ZN(n4019)
         );
  XNOR2_X1 U4573 ( .A(n4021), .B(n4074), .ZN(n4022) );
  NAND2_X1 U4574 ( .A1(n4023), .A2(n4022), .ZN(n4071) );
  INV_X1 U4575 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4026) );
  OAI21_X1 U4576 ( .B1(n4029), .B2(n4028), .A(n4027), .ZN(n4030) );
  INV_X1 U4577 ( .A(n4030), .ZN(n4031) );
  NAND2_X1 U4578 ( .A1(n4069), .A2(n3774), .ZN(n4057) );
  NAND2_X1 U4579 ( .A1(n4059), .A2(n4057), .ZN(n4080) );
  INV_X1 U4580 ( .A(n4080), .ZN(n4032) );
  NAND2_X1 U4581 ( .A1(n4079), .A2(n4032), .ZN(n4088) );
  NAND2_X1 U4582 ( .A1(n4033), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4039) );
  INV_X1 U4583 ( .A(n5395), .ZN(n4034) );
  NAND2_X1 U4584 ( .A1(n4034), .A2(n7566), .ZN(n5955) );
  NAND2_X1 U4585 ( .A1(n5395), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4035) );
  NAND2_X1 U4586 ( .A1(n5955), .A2(n4035), .ZN(n5162) );
  NOR2_X1 U4587 ( .A1(n4240), .A2(n7566), .ZN(n4036) );
  AOI21_X1 U4588 ( .B1(n5162), .B2(n4037), .A(n4036), .ZN(n4038) );
  AOI22_X1 U4589 ( .A1(n4721), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U4590 ( .A1(n4728), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U4591 ( .A1(n3660), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4729), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U4592 ( .A1(n4732), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4040) );
  NAND4_X1 U4593 ( .A1(n4043), .A2(n4042), .A3(n4041), .A4(n4040), .ZN(n4049)
         );
  AOI22_X1 U4594 ( .A1(n4727), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U4595 ( .A1(n3664), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4722), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4046) );
  AOI22_X1 U4596 ( .A1(n4118), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U4597 ( .A1(n4720), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4044) );
  NAND4_X1 U4598 ( .A1(n4047), .A2(n4046), .A3(n4045), .A4(n4044), .ZN(n4048)
         );
  AOI22_X1 U4599 ( .A1(n3967), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4231), 
        .B2(n4104), .ZN(n4050) );
  XNOR2_X2 U4600 ( .A(n4088), .B(n5158), .ZN(n5128) );
  NAND2_X1 U4601 ( .A1(n4060), .A2(n4074), .ZN(n4083) );
  INV_X1 U4602 ( .A(n4082), .ZN(n4052) );
  NAND2_X1 U4603 ( .A1(n4083), .A2(n4052), .ZN(n4105) );
  INV_X1 U4604 ( .A(n4104), .ZN(n4053) );
  XNOR2_X1 U4605 ( .A(n4105), .B(n4053), .ZN(n4055) );
  AND2_X1 U4606 ( .A1(n4055), .A2(n4054), .ZN(n4056) );
  AOI21_X1 U4607 ( .B1(n5128), .B2(n4232), .A(n4056), .ZN(n5004) );
  INV_X1 U4608 ( .A(n4057), .ZN(n4058) );
  NAND2_X1 U4609 ( .A1(n4255), .A2(n3924), .ZN(n4064) );
  INV_X1 U4610 ( .A(n4074), .ZN(n4066) );
  XNOR2_X1 U4611 ( .A(n4066), .B(n4060), .ZN(n4062) );
  NAND2_X1 U4612 ( .A1(n3923), .A2(n5172), .ZN(n4061) );
  AOI21_X1 U4613 ( .B1(n4062), .B2(n4054), .A(n4061), .ZN(n4063) );
  NAND2_X1 U4614 ( .A1(n3940), .A2(n4165), .ZN(n4065) );
  OAI211_X1 U4615 ( .C1(n4066), .C2(n3941), .A(n4065), .B(
        STATE2_REG_0__SCAN_IN), .ZN(n4067) );
  AOI21_X1 U4616 ( .B1(n3967), .B2(INSTQUEUE_REG_0__0__SCAN_IN), .A(n4067), 
        .ZN(n4070) );
  INV_X1 U4617 ( .A(n4070), .ZN(n4068) );
  NAND2_X1 U4618 ( .A1(n5487), .A2(n4232), .ZN(n4077) );
  NAND2_X1 U4619 ( .A1(n5140), .A2(n3923), .ZN(n4896) );
  OAI21_X1 U4620 ( .B1(n6594), .B2(n4074), .A(n4896), .ZN(n4075) );
  INV_X1 U4621 ( .A(n4075), .ZN(n4076) );
  NAND2_X1 U4622 ( .A1(n4077), .A2(n4076), .ZN(n4998) );
  NAND2_X1 U4623 ( .A1(n4998), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n7263)
         );
  INV_X1 U4624 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4078) );
  INV_X1 U4625 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n7349) );
  INV_X1 U4626 ( .A(n4079), .ZN(n4081) );
  NAND2_X1 U4627 ( .A1(n4081), .A2(n4080), .ZN(n5127) );
  AND2_X2 U4628 ( .A1(n4088), .A2(n5127), .ZN(n5126) );
  XNOR2_X1 U4629 ( .A(n4083), .B(n4082), .ZN(n4084) );
  OAI21_X1 U4630 ( .B1(n4084), .B2(n6594), .A(n4896), .ZN(n4085) );
  AOI21_X1 U4631 ( .B1(n5126), .B2(n4232), .A(n4085), .ZN(n7269) );
  NAND2_X1 U4632 ( .A1(n4086), .A2(n7349), .ZN(n7267) );
  INV_X1 U4633 ( .A(n7267), .ZN(n4087) );
  INV_X1 U4634 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4100) );
  AOI22_X1 U4635 ( .A1(n4728), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4092) );
  AOI22_X1 U4636 ( .A1(n4727), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U4637 ( .A1(n4721), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4720), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4090) );
  AOI22_X1 U4638 ( .A1(n3892), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4089) );
  NAND4_X1 U4639 ( .A1(n4092), .A2(n4091), .A3(n4090), .A4(n4089), .ZN(n4098)
         );
  AOI22_X1 U4640 ( .A1(n3665), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4096) );
  AOI22_X1 U4641 ( .A1(n4732), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4095) );
  AOI22_X1 U4642 ( .A1(n3660), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4094) );
  AOI22_X1 U4643 ( .A1(n4702), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4093) );
  NAND4_X1 U4644 ( .A1(n4096), .A2(n4095), .A3(n4094), .A4(n4093), .ZN(n4097)
         );
  NAND2_X1 U4645 ( .A1(n4231), .A2(n4108), .ZN(n4099) );
  NAND2_X1 U4646 ( .A1(n4102), .A2(n3749), .ZN(n4103) );
  AND2_X1 U4647 ( .A1(n4105), .A2(n4104), .ZN(n4109) );
  INV_X1 U4648 ( .A(n4109), .ZN(n4107) );
  INV_X1 U4649 ( .A(n4108), .ZN(n4106) );
  NOR2_X1 U4650 ( .A1(n4107), .A2(n4106), .ZN(n4136) );
  OAI21_X1 U4651 ( .B1(n4109), .B2(n4108), .A(n4054), .ZN(n4110) );
  AND2_X1 U4652 ( .A1(n4112), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4113)
         );
  INV_X1 U4653 ( .A(n4147), .ZN(n4127) );
  INV_X1 U4654 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4126) );
  AOI22_X1 U4655 ( .A1(n3666), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4117) );
  AOI22_X1 U4656 ( .A1(n4729), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4732), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4116) );
  AOI22_X1 U4657 ( .A1(n4720), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4115) );
  AOI22_X1 U4658 ( .A1(n4721), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4114) );
  NAND4_X1 U4659 ( .A1(n4117), .A2(n4116), .A3(n4115), .A4(n4114), .ZN(n4124)
         );
  AOI22_X1 U4660 ( .A1(n4728), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4122) );
  AOI22_X1 U4661 ( .A1(n3660), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4121) );
  AOI22_X1 U4662 ( .A1(n4718), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4722), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4120) );
  AOI22_X1 U4663 ( .A1(n4118), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4119) );
  NAND4_X1 U4664 ( .A1(n4122), .A2(n4121), .A3(n4120), .A4(n4119), .ZN(n4123)
         );
  NAND2_X1 U4665 ( .A1(n4231), .A2(n4135), .ZN(n4125) );
  OAI21_X1 U4666 ( .B1(n4126), .B2(n4025), .A(n4125), .ZN(n4150) );
  INV_X1 U4667 ( .A(n4150), .ZN(n4128) );
  NAND2_X1 U4668 ( .A1(n4147), .A2(n4128), .ZN(n4129) );
  NAND2_X1 U4669 ( .A1(n4154), .A2(n4129), .ZN(n4295) );
  INV_X1 U4670 ( .A(n4136), .ZN(n4130) );
  XNOR2_X1 U4671 ( .A(n4130), .B(n4135), .ZN(n4131) );
  NAND2_X1 U4672 ( .A1(n4131), .A2(n4054), .ZN(n4132) );
  XNOR2_X1 U4673 ( .A(n4133), .B(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6023)
         );
  INV_X1 U4674 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6438) );
  NAND2_X1 U4675 ( .A1(n4136), .A2(n4135), .ZN(n4160) );
  AOI22_X1 U4676 ( .A1(n4728), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4140) );
  AOI22_X1 U4677 ( .A1(n4727), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4139) );
  AOI22_X1 U4678 ( .A1(n4721), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4720), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4138) );
  AOI22_X1 U4679 ( .A1(n3892), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4137) );
  NAND4_X1 U4680 ( .A1(n4140), .A2(n4139), .A3(n4138), .A4(n4137), .ZN(n4146)
         );
  AOI22_X1 U4681 ( .A1(n3665), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4144) );
  AOI22_X1 U4682 ( .A1(n4732), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4143) );
  AOI22_X1 U4683 ( .A1(n3660), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4142) );
  AOI22_X1 U4684 ( .A1(n4729), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4141) );
  NAND4_X1 U4685 ( .A1(n4144), .A2(n4143), .A3(n4142), .A4(n4141), .ZN(n4145)
         );
  XNOR2_X1 U4686 ( .A(n4160), .B(n4161), .ZN(n4157) );
  INV_X1 U4687 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4149) );
  NAND2_X1 U4688 ( .A1(n4231), .A2(n4161), .ZN(n4148) );
  OAI21_X1 U4689 ( .B1(n4149), .B2(n4025), .A(n4148), .ZN(n4152) );
  AND2_X1 U4690 ( .A1(n4152), .A2(n4150), .ZN(n4151) );
  INV_X1 U4691 ( .A(n4152), .ZN(n4153) );
  NOR3_X1 U4692 ( .A1(n4155), .A2(n4307), .A3(n4222), .ZN(n4156) );
  AOI21_X1 U4693 ( .B1(n4054), .B2(n4157), .A(n4156), .ZN(n4158) );
  INV_X1 U4694 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6440) );
  NAND2_X1 U4695 ( .A1(n4158), .A2(n6440), .ZN(n6433) );
  NOR2_X1 U4696 ( .A1(n4158), .A2(n6440), .ZN(n6435) );
  AOI22_X1 U4697 ( .A1(n3967), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4231), 
        .B2(n4165), .ZN(n4159) );
  INV_X1 U4698 ( .A(n4160), .ZN(n4162) );
  NAND2_X1 U4699 ( .A1(n4162), .A2(n4161), .ZN(n4169) );
  XOR2_X1 U4700 ( .A(n4165), .B(n4169), .Z(n4163) );
  OAI22_X1 U4701 ( .A1(n4301), .A2(n4222), .B1(n4163), .B2(n6594), .ZN(n4164)
         );
  XNOR2_X1 U4702 ( .A(n4164), .B(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n7289)
         );
  NAND2_X1 U4703 ( .A1(n4054), .A2(n4165), .ZN(n4168) );
  OAI21_X1 U4704 ( .B1(n4169), .B2(n4168), .A(n4171), .ZN(n4170) );
  XNOR2_X1 U4705 ( .A(n4170), .B(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6425)
         );
  XOR2_X1 U4706 ( .A(n4171), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .Z(n6465) );
  INV_X1 U4707 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4174) );
  INV_X1 U4708 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4173) );
  INV_X1 U4709 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4172) );
  NAND2_X1 U4710 ( .A1(n6970), .A2(n3772), .ZN(n4175) );
  INV_X1 U4711 ( .A(n6970), .ZN(n4176) );
  NAND2_X1 U4712 ( .A1(n7066), .A2(n4172), .ZN(n6951) );
  XNOR2_X1 U4713 ( .A(n7066), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6943)
         );
  INV_X1 U4714 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n7330) );
  INV_X1 U4715 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n7408) );
  INV_X1 U4716 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n7423) );
  INV_X1 U4717 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n7073) );
  OAI21_X1 U4718 ( .B1(n7423), .B2(n7073), .A(n7066), .ZN(n4182) );
  NAND2_X1 U4719 ( .A1(n6911), .A2(n4182), .ZN(n6882) );
  NOR3_X1 U4720 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A3(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n4183) );
  NOR4_X1 U4721 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4185) );
  NOR2_X1 U4722 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6867) );
  AND2_X1 U4723 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4905) );
  AND2_X1 U4724 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4917) );
  NAND2_X1 U4725 ( .A1(n4905), .A2(n4917), .ZN(n6878) );
  NAND2_X1 U4726 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4920) );
  NAND2_X1 U4727 ( .A1(n4187), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6853) );
  NAND2_X1 U4728 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6988) );
  INV_X1 U4729 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4940) );
  INV_X1 U4730 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6986) );
  AND2_X1 U4731 ( .A1(n6986), .A2(n6842), .ZN(n4186) );
  AND2_X1 U4732 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6548) );
  NAND2_X1 U4733 ( .A1(n6548), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4941) );
  INV_X1 U4734 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6552) );
  NAND2_X1 U4735 ( .A1(n4187), .A2(n6552), .ZN(n4754) );
  OAI21_X1 U4736 ( .B1(n4941), .B2(n4940), .A(n4754), .ZN(n4188) );
  OAI211_X1 U4737 ( .C1(n6521), .C2(n4940), .A(n6539), .B(n4188), .ZN(n4189)
         );
  XNOR2_X1 U4738 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4201) );
  NAND2_X1 U4739 ( .A1(n3937), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4205) );
  AOI222_X1 U4740 ( .A1(n4191), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B1(
        n4191), .B2(n7551), .C1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n7551), 
        .ZN(n4761) );
  NAND2_X1 U4741 ( .A1(n4191), .A2(n7551), .ZN(n4192) );
  AOI22_X1 U4742 ( .A1(n4193), .A2(n3967), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n7318), .ZN(n4229) );
  INV_X1 U4743 ( .A(n4193), .ZN(n4760) );
  XNOR2_X1 U4744 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4194) );
  XNOR2_X1 U4745 ( .A(n4195), .B(n4194), .ZN(n4759) );
  XNOR2_X1 U4746 ( .A(n4197), .B(n4196), .ZN(n4758) );
  INV_X1 U4747 ( .A(n4758), .ZN(n4198) );
  INV_X1 U4748 ( .A(n4218), .ZN(n4224) );
  AND2_X1 U4749 ( .A1(n5228), .A2(n5172), .ZN(n4199) );
  XNOR2_X1 U4750 ( .A(n4201), .B(n4200), .ZN(n4757) );
  INV_X1 U4751 ( .A(n4757), .ZN(n4202) );
  NOR2_X1 U4752 ( .A1(n4025), .A2(n4222), .ZN(n4207) );
  AOI21_X1 U4753 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n4202), .A(n4207), .ZN(
        n4211) );
  INV_X1 U4754 ( .A(n4211), .ZN(n4217) );
  OAI21_X1 U4755 ( .B1(n4203), .B2(n5228), .A(n5172), .ZN(n4204) );
  AOI21_X1 U4756 ( .B1(n3967), .B2(n4757), .A(n4204), .ZN(n4212) );
  INV_X1 U4757 ( .A(n4212), .ZN(n4216) );
  OAI21_X1 U4758 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n3937), .A(n4205), 
        .ZN(n4209) );
  INV_X1 U4759 ( .A(n4209), .ZN(n4206) );
  NAND2_X1 U4760 ( .A1(n4231), .A2(n4206), .ZN(n4214) );
  INV_X1 U4761 ( .A(n4207), .ZN(n4213) );
  OAI21_X1 U4762 ( .B1(n4885), .B2(n4209), .A(n4208), .ZN(n4210) );
  AOI222_X1 U4763 ( .A1(n4214), .A2(n4213), .B1(n4212), .B2(n4211), .C1(n4210), 
        .C2(n4223), .ZN(n4215) );
  AOI21_X1 U4764 ( .B1(n4217), .B2(n4216), .A(n4215), .ZN(n4221) );
  INV_X1 U4765 ( .A(n4223), .ZN(n4219) );
  AOI211_X1 U4766 ( .C1(n3967), .C2(n4758), .A(n4219), .B(n4218), .ZN(n4220)
         );
  OAI222_X1 U4767 ( .A1(n4224), .A2(n4223), .B1(n4222), .B2(n4226), .C1(n4221), 
        .C2(n4220), .ZN(n4225) );
  AOI222_X1 U4768 ( .A1(n4229), .A2(n4228), .B1(n4229), .B2(n4227), .C1(n4228), 
        .C2(n4227), .ZN(n4230) );
  AOI21_X1 U4769 ( .B1(n4231), .B2(n4761), .A(n4230), .ZN(n4235) );
  NAND2_X1 U4770 ( .A1(n4232), .A2(n4761), .ZN(n4233) );
  NOR2_X1 U4771 ( .A1(n4025), .A2(n4233), .ZN(n4234) );
  OR2_X2 U4772 ( .A1(n4235), .A2(n4234), .ZN(n6593) );
  NAND2_X1 U4773 ( .A1(n5177), .A2(n4237), .ZN(n4238) );
  AND2_X1 U4774 ( .A1(n5043), .A2(n5140), .ZN(n4239) );
  NAND2_X1 U4775 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4278) );
  INV_X1 U4776 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6845) );
  INV_X1 U4777 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6835) );
  INV_X1 U4778 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4695) );
  INV_X1 U4779 ( .A(n4716), .ZN(n4245) );
  NAND2_X1 U4780 ( .A1(n4245), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4247)
         );
  INV_X1 U4781 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4246) );
  AND2_X1 U4782 ( .A1(n4248), .A2(n5870), .ZN(n7321) );
  OR2_X1 U4783 ( .A1(n7321), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4249) );
  NAND2_X1 U4784 ( .A1(n7318), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4251) );
  NAND2_X1 U4785 ( .A1(n7608), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4250) );
  NAND2_X1 U4786 ( .A1(n4251), .A2(n4250), .ZN(n4997) );
  AND2_X2 U4787 ( .A1(n7305), .A2(n7318), .ZN(n7370) );
  NAND2_X1 U4788 ( .A1(n7370), .A2(REIP_REG_31__SCAN_IN), .ZN(n4944) );
  NAND2_X1 U4789 ( .A1(n7296), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4252)
         );
  OAI211_X1 U4790 ( .C1(n4966), .C2(n7302), .A(n4944), .B(n4252), .ZN(n4253)
         );
  NAND2_X1 U4791 ( .A1(n5126), .A2(n4442), .ZN(n4254) );
  INV_X1 U4792 ( .A(n4748), .ZN(n4607) );
  NAND2_X1 U4793 ( .A1(n4255), .A2(n4442), .ZN(n4260) );
  AOI22_X1 U4794 ( .A1(n4749), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n7584), .ZN(n4258) );
  AND2_X1 U4795 ( .A1(n4256), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4270) );
  NAND2_X1 U4796 ( .A1(n4270), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4257) );
  AND2_X1 U4797 ( .A1(n4258), .A2(n4257), .ZN(n4259) );
  NAND2_X1 U4798 ( .A1(n4260), .A2(n4259), .ZN(n5080) );
  NAND2_X1 U4799 ( .A1(n4262), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4995) );
  INV_X1 U4800 ( .A(n4270), .ZN(n4291) );
  NAND2_X1 U4801 ( .A1(n4749), .A2(EAX_REG_0__SCAN_IN), .ZN(n4265) );
  NAND2_X1 U4802 ( .A1(n7584), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4264)
         );
  OAI211_X1 U4803 ( .C1(n4291), .C2(n5049), .A(n4265), .B(n4264), .ZN(n4266)
         );
  AOI21_X1 U4804 ( .B1(n4263), .B2(n4442), .A(n4266), .ZN(n4996) );
  INV_X1 U4805 ( .A(n4996), .ZN(n4268) );
  NOR2_X2 U4806 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4267) );
  OR2_X1 U4807 ( .A1(n4268), .A2(n4284), .ZN(n4269) );
  NAND2_X1 U4808 ( .A1(n5098), .A2(n5099), .ZN(n4275) );
  NAND2_X1 U4809 ( .A1(n4270), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4274) );
  INV_X1 U4810 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5728) );
  INV_X1 U4811 ( .A(n4284), .ZN(n4960) );
  OAI21_X1 U4812 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n4278), .ZN(n7275) );
  NAND2_X1 U4813 ( .A1(n4960), .A2(n7275), .ZN(n4271) );
  OAI21_X1 U4814 ( .B1(n4607), .B2(n5728), .A(n4271), .ZN(n4272) );
  AOI21_X1 U4815 ( .B1(n4749), .B2(EAX_REG_2__SCAN_IN), .A(n4272), .ZN(n4273)
         );
  AND2_X1 U4816 ( .A1(n4274), .A2(n4273), .ZN(n5101) );
  NAND2_X1 U4817 ( .A1(n4275), .A2(n5101), .ZN(n4277) );
  NAND2_X1 U4818 ( .A1(n4277), .A2(n4276), .ZN(n5006) );
  INV_X1 U4819 ( .A(n4278), .ZN(n4280) );
  INV_X1 U4820 ( .A(n4279), .ZN(n4285) );
  OAI21_X1 U4821 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n4280), .A(n4285), 
        .ZN(n7447) );
  AOI22_X1 U4822 ( .A1(n4960), .A2(n7447), .B1(n4748), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4282) );
  NAND2_X1 U4823 ( .A1(n4749), .A2(EAX_REG_3__SCAN_IN), .ZN(n4281) );
  OAI211_X1 U4824 ( .C1(n4291), .C2(n6518), .A(n4282), .B(n4281), .ZN(n4283)
         );
  AOI21_X1 U4825 ( .B1(n5128), .B2(n4442), .A(n4283), .ZN(n5009) );
  NOR2_X2 U4826 ( .A1(n5006), .A2(n5009), .ZN(n5007) );
  INV_X1 U4827 ( .A(n4442), .ZN(n4432) );
  INV_X1 U4828 ( .A(n4296), .ZN(n4288) );
  INV_X1 U4829 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4286) );
  NAND2_X1 U4830 ( .A1(n4286), .A2(n4285), .ZN(n4287) );
  NAND2_X1 U4831 ( .A1(n4288), .A2(n4287), .ZN(n7465) );
  OAI21_X1 U4832 ( .B1(n7608), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n7584), 
        .ZN(n4290) );
  NAND2_X1 U4833 ( .A1(n4749), .A2(EAX_REG_4__SCAN_IN), .ZN(n4289) );
  OAI211_X1 U4834 ( .C1(n4291), .C2(n7551), .A(n4290), .B(n4289), .ZN(n4292)
         );
  OAI21_X1 U4835 ( .B1(n4284), .B2(n7465), .A(n4292), .ZN(n4293) );
  OAI21_X1 U4836 ( .B1(n4294), .B2(n4432), .A(n4293), .ZN(n5067) );
  INV_X1 U4837 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n7282) );
  OAI21_X1 U4838 ( .B1(n4296), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n4309), 
        .ZN(n7277) );
  NAND2_X1 U4839 ( .A1(n7277), .A2(n4960), .ZN(n4297) );
  OAI21_X1 U4840 ( .B1(n7282), .B2(n4607), .A(n4297), .ZN(n4298) );
  AOI21_X1 U4841 ( .B1(n4749), .B2(EAX_REG_5__SCAN_IN), .A(n4298), .ZN(n4299)
         );
  NAND2_X1 U4842 ( .A1(n4300), .A2(n4299), .ZN(n5107) );
  INV_X1 U4843 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4304) );
  OR2_X1 U4844 ( .A1(n4310), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4302) );
  NAND2_X1 U4845 ( .A1(n4328), .A2(n4302), .ZN(n7500) );
  AOI22_X1 U4846 ( .A1(n7500), .A2(n4267), .B1(n4748), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4303) );
  NAND2_X1 U4847 ( .A1(n4308), .A2(n4442), .ZN(n4316) );
  AND2_X1 U4848 ( .A1(n4309), .A2(n7479), .ZN(n4311) );
  OR2_X1 U4849 ( .A1(n4311), .A2(n4310), .ZN(n7486) );
  INV_X1 U4850 ( .A(n7486), .ZN(n4314) );
  NOR2_X1 U4851 ( .A1(n7479), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4312) );
  AOI21_X1 U4852 ( .B1(n4749), .B2(EAX_REG_6__SCAN_IN), .A(n4312), .ZN(n4313)
         );
  MUX2_X1 U4853 ( .A(n4314), .B(n4313), .S(n4284), .Z(n4315) );
  NAND2_X1 U4854 ( .A1(n4316), .A2(n4315), .ZN(n5598) );
  AOI22_X1 U4855 ( .A1(n4728), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4729), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4321) );
  AOI22_X1 U4856 ( .A1(n3665), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4320) );
  AOI22_X1 U4857 ( .A1(n4720), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4319) );
  AOI22_X1 U4858 ( .A1(n4721), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4318) );
  NAND4_X1 U4859 ( .A1(n4321), .A2(n4320), .A3(n4319), .A4(n4318), .ZN(n4327)
         );
  AOI22_X1 U4860 ( .A1(n4727), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4325) );
  AOI22_X1 U4861 ( .A1(n4731), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4732), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4324) );
  AOI22_X1 U4862 ( .A1(n3660), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4323) );
  AOI22_X1 U4863 ( .A1(n3892), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4322) );
  NAND4_X1 U4864 ( .A1(n4325), .A2(n4324), .A3(n4323), .A4(n4322), .ZN(n4326)
         );
  OAI21_X1 U4865 ( .B1(n4327), .B2(n4326), .A(n4442), .ZN(n4332) );
  NAND2_X1 U4866 ( .A1(n4749), .A2(EAX_REG_8__SCAN_IN), .ZN(n4331) );
  XNOR2_X1 U4867 ( .A(n4328), .B(n5798), .ZN(n6426) );
  NAND2_X1 U4868 ( .A1(n6426), .A2(n4267), .ZN(n4330) );
  NAND2_X1 U4869 ( .A1(n4748), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4329)
         );
  XNOR2_X1 U4870 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n4334), .ZN(n6468) );
  INV_X1 U4871 ( .A(n6468), .ZN(n4349) );
  AOI22_X1 U4872 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n3666), .B1(n4731), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4338) );
  AOI22_X1 U4873 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n4729), .B1(n4719), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4337) );
  AOI22_X1 U4874 ( .A1(n3660), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4336) );
  AOI22_X1 U4875 ( .A1(n4727), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4335) );
  NAND4_X1 U4876 ( .A1(n4338), .A2(n4337), .A3(n4336), .A4(n4335), .ZN(n4344)
         );
  AOI22_X1 U4877 ( .A1(n4721), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4342) );
  AOI22_X1 U4878 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(n3866), .B1(n3664), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4341) );
  AOI22_X1 U4879 ( .A1(INSTQUEUE_REG_2__1__SCAN_IN), .A2(n4720), .B1(n4722), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4340) );
  AOI22_X1 U4880 ( .A1(n4732), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4339) );
  NAND4_X1 U4881 ( .A1(n4342), .A2(n4341), .A3(n4340), .A4(n4339), .ZN(n4343)
         );
  OAI21_X1 U4882 ( .B1(n4344), .B2(n4343), .A(n4442), .ZN(n4347) );
  NAND2_X1 U4883 ( .A1(n4749), .A2(EAX_REG_9__SCAN_IN), .ZN(n4346) );
  NAND2_X1 U4884 ( .A1(n4748), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4345)
         );
  NAND3_X1 U4885 ( .A1(n4347), .A2(n4346), .A3(n4345), .ZN(n4348) );
  AOI21_X1 U4886 ( .B1(n4349), .B2(n4267), .A(n4348), .ZN(n5810) );
  XNOR2_X1 U4887 ( .A(n4350), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6971)
         );
  NAND2_X1 U4888 ( .A1(n6971), .A2(n4267), .ZN(n4365) );
  AOI22_X1 U4889 ( .A1(n4727), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4354) );
  AOI22_X1 U4890 ( .A1(n3660), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4729), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4353) );
  AOI22_X1 U4891 ( .A1(n4721), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4352) );
  AOI22_X1 U4892 ( .A1(n4718), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4351) );
  NAND4_X1 U4893 ( .A1(n4354), .A2(n4353), .A3(n4352), .A4(n4351), .ZN(n4360)
         );
  AOI22_X1 U4894 ( .A1(n4732), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4358) );
  AOI22_X1 U4895 ( .A1(n4728), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4720), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4357) );
  AOI22_X1 U4896 ( .A1(n3666), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4722), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4356) );
  AOI22_X1 U4897 ( .A1(n4730), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4355) );
  NAND4_X1 U4898 ( .A1(n4358), .A2(n4357), .A3(n4356), .A4(n4355), .ZN(n4359)
         );
  OAI21_X1 U4899 ( .B1(n4360), .B2(n4359), .A(n4442), .ZN(n4363) );
  NAND2_X1 U4900 ( .A1(n4749), .A2(EAX_REG_10__SCAN_IN), .ZN(n4362) );
  NAND2_X1 U4901 ( .A1(n4748), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4361)
         );
  AND3_X1 U4902 ( .A1(n4363), .A2(n4362), .A3(n4361), .ZN(n4364) );
  NAND2_X1 U4903 ( .A1(n4365), .A2(n4364), .ZN(n5832) );
  XNOR2_X1 U4904 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n4366), .ZN(n6964)
         );
  AOI22_X1 U4905 ( .A1(n4721), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4367), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4371) );
  AOI22_X1 U4906 ( .A1(n3660), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4370) );
  AOI22_X1 U4907 ( .A1(n3892), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4369) );
  AOI22_X1 U4908 ( .A1(n4729), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4368) );
  NAND4_X1 U4909 ( .A1(n4371), .A2(n4370), .A3(n4369), .A4(n4368), .ZN(n4377)
         );
  AOI22_X1 U4910 ( .A1(n4728), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4375) );
  AOI22_X1 U4911 ( .A1(n4732), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4374) );
  AOI22_X1 U4912 ( .A1(n4718), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4720), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4373) );
  AOI22_X1 U4913 ( .A1(n3666), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4372) );
  NAND4_X1 U4914 ( .A1(n4375), .A2(n4374), .A3(n4373), .A4(n4372), .ZN(n4376)
         );
  OAI21_X1 U4915 ( .B1(n4377), .B2(n4376), .A(n4442), .ZN(n4380) );
  NAND2_X1 U4916 ( .A1(n4749), .A2(EAX_REG_11__SCAN_IN), .ZN(n4379) );
  NAND2_X1 U4917 ( .A1(n4748), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4378)
         );
  AND3_X1 U4918 ( .A1(n4380), .A2(n4379), .A3(n4378), .ZN(n4381) );
  OAI21_X1 U4919 ( .B1(n6964), .B2(n4284), .A(n4381), .ZN(n5852) );
  NAND2_X1 U4920 ( .A1(n5831), .A2(n5852), .ZN(n5850) );
  INV_X1 U4921 ( .A(n5850), .ZN(n4398) );
  XNOR2_X1 U4922 ( .A(n4382), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6955)
         );
  AOI22_X1 U4923 ( .A1(n4721), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4386) );
  AOI22_X1 U4924 ( .A1(n4732), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4385) );
  AOI22_X1 U4925 ( .A1(n3892), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4384) );
  AOI22_X1 U4926 ( .A1(n4729), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4383) );
  NAND4_X1 U4927 ( .A1(n4386), .A2(n4385), .A3(n4384), .A4(n4383), .ZN(n4392)
         );
  AOI22_X1 U4928 ( .A1(n4728), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4390) );
  AOI22_X1 U4929 ( .A1(n3665), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4389) );
  AOI22_X1 U4930 ( .A1(n4718), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4720), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4388) );
  AOI22_X1 U4931 ( .A1(n3660), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4387) );
  NAND4_X1 U4932 ( .A1(n4390), .A2(n4389), .A3(n4388), .A4(n4387), .ZN(n4391)
         );
  OAI21_X1 U4933 ( .B1(n4392), .B2(n4391), .A(n4442), .ZN(n4395) );
  NAND2_X1 U4934 ( .A1(n4749), .A2(EAX_REG_12__SCAN_IN), .ZN(n4394) );
  NAND2_X1 U4935 ( .A1(n4748), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4393)
         );
  NAND3_X1 U4936 ( .A1(n4395), .A2(n4394), .A3(n4393), .ZN(n4396) );
  AOI21_X1 U4937 ( .B1(n6955), .B2(n4267), .A(n4396), .ZN(n6448) );
  INV_X1 U4938 ( .A(n6448), .ZN(n4397) );
  NAND2_X1 U4939 ( .A1(n4398), .A2(n4397), .ZN(n4414) );
  AOI22_X1 U4940 ( .A1(n4727), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4402) );
  AOI22_X1 U4941 ( .A1(n3660), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4401) );
  AOI22_X1 U4942 ( .A1(n4732), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4400) );
  AOI22_X1 U4943 ( .A1(n4729), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4722), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4399) );
  NAND4_X1 U4944 ( .A1(n4402), .A2(n4401), .A3(n4400), .A4(n4399), .ZN(n4408)
         );
  AOI22_X1 U4945 ( .A1(n3666), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4406) );
  AOI22_X1 U4946 ( .A1(n3866), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4720), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4405) );
  AOI22_X1 U4947 ( .A1(n4721), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4404) );
  AOI22_X1 U4948 ( .A1(n4730), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4403) );
  NAND4_X1 U4949 ( .A1(n4406), .A2(n4405), .A3(n4404), .A4(n4403), .ZN(n4407)
         );
  OR2_X1 U4950 ( .A1(n4408), .A2(n4407), .ZN(n4409) );
  NAND2_X1 U4951 ( .A1(n4749), .A2(EAX_REG_13__SCAN_IN), .ZN(n4413) );
  INV_X1 U4952 ( .A(n4410), .ZN(n4411) );
  XNOR2_X1 U4953 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(n4411), .ZN(n6947)
         );
  AOI22_X1 U4954 ( .A1(n4960), .A2(n6947), .B1(n4748), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4412) );
  NAND2_X1 U4955 ( .A1(n4413), .A2(n4412), .ZN(n6482) );
  NAND2_X1 U4956 ( .A1(n6481), .A2(n6482), .ZN(n4417) );
  NAND2_X1 U4957 ( .A1(n6447), .A2(n4415), .ZN(n4416) );
  NAND2_X2 U4958 ( .A1(n4417), .A2(n4416), .ZN(n6501) );
  AOI22_X1 U4959 ( .A1(n4721), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4421) );
  AOI22_X1 U4960 ( .A1(n3665), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4420) );
  AOI22_X1 U4961 ( .A1(n4720), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4419) );
  AOI22_X1 U4962 ( .A1(n4729), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4418) );
  NAND4_X1 U4963 ( .A1(n4421), .A2(n4420), .A3(n4419), .A4(n4418), .ZN(n4427)
         );
  AOI22_X1 U4964 ( .A1(n4727), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4425) );
  AOI22_X1 U4965 ( .A1(n4732), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4424) );
  AOI22_X1 U4966 ( .A1(n4718), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4722), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4423) );
  AOI22_X1 U4967 ( .A1(n3850), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4422) );
  NAND4_X1 U4968 ( .A1(n4425), .A2(n4424), .A3(n4423), .A4(n4422), .ZN(n4426)
         );
  NOR2_X1 U4969 ( .A1(n4427), .A2(n4426), .ZN(n4431) );
  XNOR2_X1 U4970 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4428), .ZN(n6937)
         );
  AOI22_X1 U4971 ( .A1(n4267), .A2(n6937), .B1(n4748), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4430) );
  NAND2_X1 U4972 ( .A1(n4749), .A2(EAX_REG_14__SCAN_IN), .ZN(n4429) );
  OAI211_X1 U4973 ( .C1(n4432), .C2(n4431), .A(n4430), .B(n4429), .ZN(n6500)
         );
  XOR2_X1 U4974 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n4433), .Z(n6929) );
  INV_X1 U4975 ( .A(n6929), .ZN(n6751) );
  AOI22_X1 U4976 ( .A1(n3660), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4729), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4437) );
  AOI22_X1 U4977 ( .A1(n3665), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4436) );
  AOI22_X1 U4978 ( .A1(n4731), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4722), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4435) );
  AOI22_X1 U4979 ( .A1(n4721), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4434) );
  NAND4_X1 U4980 ( .A1(n4437), .A2(n4436), .A3(n4435), .A4(n4434), .ZN(n4444)
         );
  AOI22_X1 U4981 ( .A1(n3866), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4441) );
  AOI22_X1 U4982 ( .A1(n4727), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4440) );
  AOI22_X1 U4983 ( .A1(n4732), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4439) );
  AOI22_X1 U4984 ( .A1(n4720), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4438) );
  NAND4_X1 U4985 ( .A1(n4441), .A2(n4440), .A3(n4439), .A4(n4438), .ZN(n4443)
         );
  OAI21_X1 U4986 ( .B1(n4444), .B2(n4443), .A(n4442), .ZN(n4447) );
  NAND2_X1 U4987 ( .A1(n4749), .A2(EAX_REG_15__SCAN_IN), .ZN(n4446) );
  NAND2_X1 U4988 ( .A1(n4748), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4445)
         );
  NAND3_X1 U4989 ( .A1(n4447), .A2(n4446), .A3(n4445), .ZN(n4448) );
  AOI21_X1 U4990 ( .B1(n6751), .B2(n4267), .A(n4448), .ZN(n6742) );
  XNOR2_X1 U4991 ( .A(n4449), .B(n4243), .ZN(n6922) );
  AOI22_X1 U4992 ( .A1(n3665), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4453) );
  AOI22_X1 U4993 ( .A1(n4729), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4452) );
  AOI22_X1 U4994 ( .A1(n4727), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4722), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4451) );
  AOI22_X1 U4995 ( .A1(n3660), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4450) );
  NAND4_X1 U4996 ( .A1(n4453), .A2(n4452), .A3(n4451), .A4(n4450), .ZN(n4459)
         );
  AOI22_X1 U4997 ( .A1(n4721), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4457) );
  AOI22_X1 U4998 ( .A1(n3866), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4456) );
  AOI22_X1 U4999 ( .A1(n4720), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4455) );
  AOI22_X1 U5000 ( .A1(n4732), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4454) );
  NAND4_X1 U5001 ( .A1(n4457), .A2(n4456), .A3(n4455), .A4(n4454), .ZN(n4458)
         );
  NOR2_X1 U5002 ( .A1(n4459), .A2(n4458), .ZN(n4461) );
  AOI22_X1 U5003 ( .A1(n4749), .A2(EAX_REG_16__SCAN_IN), .B1(n4748), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4460) );
  OAI21_X1 U5004 ( .B1(n4691), .B2(n4461), .A(n4460), .ZN(n4462) );
  AOI21_X1 U5005 ( .B1(n6922), .B2(n4267), .A(n4462), .ZN(n6731) );
  OR2_X1 U5006 ( .A1(n4463), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4464)
         );
  NAND2_X1 U5007 ( .A1(n4464), .A2(n4493), .ZN(n7295) );
  INV_X1 U5008 ( .A(n7295), .ZN(n7505) );
  AOI22_X1 U5009 ( .A1(n3850), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4468) );
  AOI22_X1 U5010 ( .A1(n3665), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4729), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4467) );
  AOI22_X1 U5011 ( .A1(n4721), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4466) );
  AOI22_X1 U5012 ( .A1(n4732), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4465) );
  NAND4_X1 U5013 ( .A1(n4468), .A2(n4467), .A3(n4466), .A4(n4465), .ZN(n4474)
         );
  AOI22_X1 U5014 ( .A1(n3866), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4472) );
  AOI22_X1 U5015 ( .A1(n4727), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4471) );
  AOI22_X1 U5016 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n4720), .B1(n4722), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4470) );
  AOI22_X1 U5017 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n4719), .B1(n4730), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4469) );
  NAND4_X1 U5018 ( .A1(n4472), .A2(n4471), .A3(n4470), .A4(n4469), .ZN(n4473)
         );
  OR2_X1 U5019 ( .A1(n4474), .A2(n4473), .ZN(n4478) );
  INV_X1 U5020 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4476) );
  NAND2_X1 U5021 ( .A1(n7584), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4475)
         );
  OAI211_X1 U5022 ( .C1(n4713), .C2(n4476), .A(n4284), .B(n4475), .ZN(n4477)
         );
  AOI21_X1 U5023 ( .B1(n4744), .B2(n4478), .A(n4477), .ZN(n4479) );
  AOI21_X1 U5024 ( .B1(n7505), .B2(n4267), .A(n4479), .ZN(n6782) );
  AOI22_X1 U5025 ( .A1(n4721), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4483) );
  AOI22_X1 U5026 ( .A1(n3866), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4482) );
  AOI22_X1 U5027 ( .A1(n4731), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4729), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4481) );
  AOI22_X1 U5028 ( .A1(n3850), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4480) );
  NAND4_X1 U5029 ( .A1(n4483), .A2(n4482), .A3(n4481), .A4(n4480), .ZN(n4489)
         );
  AOI22_X1 U5030 ( .A1(n4732), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4487) );
  AOI22_X1 U5031 ( .A1(n3664), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4720), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4486) );
  AOI22_X1 U5032 ( .A1(n4722), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4485) );
  AOI22_X1 U5033 ( .A1(n3666), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4484) );
  NAND4_X1 U5034 ( .A1(n4487), .A2(n4486), .A3(n4485), .A4(n4484), .ZN(n4488)
         );
  NOR2_X1 U5035 ( .A1(n4489), .A2(n4488), .ZN(n4492) );
  AOI21_X1 U5036 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n6720), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4490) );
  AOI21_X1 U5037 ( .B1(n4749), .B2(EAX_REG_18__SCAN_IN), .A(n4490), .ZN(n4491)
         );
  OAI21_X1 U5038 ( .B1(n4691), .B2(n4492), .A(n4491), .ZN(n4495) );
  XNOR2_X1 U5039 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n4493), .ZN(n6724)
         );
  NAND2_X1 U5040 ( .A1(n4960), .A2(n6724), .ZN(n4494) );
  NAND2_X1 U5041 ( .A1(n4495), .A2(n4494), .ZN(n6718) );
  INV_X1 U5042 ( .A(n4515), .ZN(n4498) );
  OR2_X1 U5043 ( .A1(n4496), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4497)
         );
  NAND2_X1 U5044 ( .A1(n4498), .A2(n4497), .ZN(n7525) );
  AOI22_X1 U5045 ( .A1(n3866), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4502) );
  AOI22_X1 U5046 ( .A1(n4729), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4732), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4501) );
  AOI22_X1 U5047 ( .A1(n3666), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4500) );
  AOI22_X1 U5048 ( .A1(n3864), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3892), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4499) );
  NAND4_X1 U5049 ( .A1(n4502), .A2(n4501), .A3(n4500), .A4(n4499), .ZN(n4508)
         );
  AOI22_X1 U5050 ( .A1(n3660), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4506) );
  AOI22_X1 U5051 ( .A1(n4718), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4505) );
  AOI22_X1 U5052 ( .A1(n4721), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4504) );
  AOI22_X1 U5053 ( .A1(n4719), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4503) );
  NAND4_X1 U5054 ( .A1(n4506), .A2(n4505), .A3(n4504), .A4(n4503), .ZN(n4507)
         );
  NOR2_X1 U5055 ( .A1(n4508), .A2(n4507), .ZN(n4509) );
  NOR2_X1 U5056 ( .A1(n4691), .A2(n4509), .ZN(n4513) );
  INV_X1 U5057 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4511) );
  NAND2_X1 U5058 ( .A1(n7584), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4510)
         );
  OAI211_X1 U5059 ( .C1(n4713), .C2(n4511), .A(n4284), .B(n4510), .ZN(n4512)
         );
  OAI22_X1 U5060 ( .A1(n7525), .A2(n4284), .B1(n4513), .B2(n4512), .ZN(n6771)
         );
  INV_X1 U5061 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6905) );
  XNOR2_X1 U5062 ( .A(n4515), .B(n6905), .ZN(n6909) );
  NAND2_X1 U5063 ( .A1(n6909), .A2(n4267), .ZN(n4531) );
  AOI22_X1 U5064 ( .A1(n4731), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4729), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4519) );
  AOI22_X1 U5065 ( .A1(n4727), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4518) );
  AOI22_X1 U5066 ( .A1(n3866), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4720), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4517) );
  AOI22_X1 U5067 ( .A1(n4732), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3892), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4516) );
  NAND4_X1 U5068 ( .A1(n4519), .A2(n4518), .A3(n4517), .A4(n4516), .ZN(n4525)
         );
  AOI22_X1 U5069 ( .A1(n4721), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4523) );
  AOI22_X1 U5070 ( .A1(n3666), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4522) );
  AOI22_X1 U5071 ( .A1(n4718), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4521) );
  AOI22_X1 U5072 ( .A1(n4730), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4520) );
  NAND4_X1 U5073 ( .A1(n4523), .A2(n4522), .A3(n4521), .A4(n4520), .ZN(n4524)
         );
  NOR2_X1 U5074 ( .A1(n4525), .A2(n4524), .ZN(n4529) );
  NAND2_X1 U5075 ( .A1(n7584), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4526)
         );
  NAND2_X1 U5076 ( .A1(n4284), .A2(n4526), .ZN(n4527) );
  AOI21_X1 U5077 ( .B1(n4749), .B2(EAX_REG_20__SCAN_IN), .A(n4527), .ZN(n4528)
         );
  OAI21_X1 U5078 ( .B1(n4691), .B2(n4529), .A(n4528), .ZN(n4530) );
  NAND2_X1 U5079 ( .A1(n4531), .A2(n4530), .ZN(n6705) );
  AND2_X1 U5080 ( .A1(n4532), .A2(n6897), .ZN(n4533) );
  OR2_X1 U5081 ( .A1(n4533), .A2(n4550), .ZN(n6700) );
  AOI22_X1 U5082 ( .A1(n3666), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4538) );
  AOI22_X1 U5083 ( .A1(n3660), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4537) );
  AOI22_X1 U5084 ( .A1(n3879), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4720), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4536) );
  AOI22_X1 U5085 ( .A1(n4721), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4535) );
  NAND4_X1 U5086 ( .A1(n4538), .A2(n4537), .A3(n4536), .A4(n4535), .ZN(n4545)
         );
  AOI22_X1 U5087 ( .A1(n3866), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4543) );
  AOI22_X1 U5088 ( .A1(n4732), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4722), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4542) );
  AOI22_X1 U5089 ( .A1(n4731), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4541) );
  AOI22_X1 U5090 ( .A1(n4729), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4540) );
  NAND4_X1 U5091 ( .A1(n4543), .A2(n4542), .A3(n4541), .A4(n4540), .ZN(n4544)
         );
  OR2_X1 U5092 ( .A1(n4545), .A2(n4544), .ZN(n4548) );
  NAND2_X1 U5093 ( .A1(n4749), .A2(EAX_REG_21__SCAN_IN), .ZN(n4546) );
  OAI211_X1 U5094 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6897), .A(n4546), .B(
        n4284), .ZN(n4547) );
  AOI21_X1 U5095 ( .B1(n4744), .B2(n4548), .A(n4547), .ZN(n4549) );
  AOI21_X1 U5096 ( .B1(n6899), .B2(n4267), .A(n4549), .ZN(n6694) );
  INV_X1 U5097 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6889) );
  XNOR2_X1 U5098 ( .A(n4550), .B(n6889), .ZN(n6893) );
  AOI22_X1 U5099 ( .A1(n4728), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4554) );
  AOI22_X1 U5100 ( .A1(n3665), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4729), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4553) );
  AOI22_X1 U5101 ( .A1(n4732), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4720), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4552) );
  AOI22_X1 U5102 ( .A1(n3664), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4551) );
  NAND4_X1 U5103 ( .A1(n4554), .A2(n4553), .A3(n4552), .A4(n4551), .ZN(n4560)
         );
  AOI22_X1 U5104 ( .A1(n4731), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4558) );
  AOI22_X1 U5105 ( .A1(n3660), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3892), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4557) );
  AOI22_X1 U5106 ( .A1(n4721), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4556) );
  AOI22_X1 U5107 ( .A1(n4727), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4555) );
  NAND4_X1 U5108 ( .A1(n4558), .A2(n4557), .A3(n4556), .A4(n4555), .ZN(n4559)
         );
  OR2_X1 U5109 ( .A1(n4560), .A2(n4559), .ZN(n4563) );
  NAND2_X1 U5110 ( .A1(n4749), .A2(EAX_REG_22__SCAN_IN), .ZN(n4561) );
  OAI211_X1 U5111 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6889), .A(n4561), .B(
        n4284), .ZN(n4562) );
  AOI21_X1 U5112 ( .B1(n4744), .B2(n4563), .A(n4562), .ZN(n4564) );
  AOI21_X1 U5113 ( .B1(n6893), .B2(n4267), .A(n4564), .ZN(n6684) );
  NAND2_X1 U5114 ( .A1(n4566), .A2(n4565), .ZN(n4567) );
  NAND2_X1 U5115 ( .A1(n4596), .A2(n4567), .ZN(n7542) );
  AOI22_X1 U5116 ( .A1(n4728), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4571) );
  AOI22_X1 U5117 ( .A1(n4727), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4570) );
  AOI22_X1 U5118 ( .A1(n4655), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4569) );
  AOI22_X1 U5119 ( .A1(n3892), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4568) );
  NAND4_X1 U5120 ( .A1(n4571), .A2(n4570), .A3(n4569), .A4(n4568), .ZN(n4577)
         );
  AOI22_X1 U5121 ( .A1(n3666), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4575) );
  AOI22_X1 U5122 ( .A1(n4732), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4574) );
  AOI22_X1 U5123 ( .A1(n3660), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4573) );
  AOI22_X1 U5124 ( .A1(n4729), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4572) );
  NAND4_X1 U5125 ( .A1(n4575), .A2(n4574), .A3(n4573), .A4(n4572), .ZN(n4576)
         );
  OR2_X1 U5126 ( .A1(n4577), .A2(n4576), .ZN(n4589) );
  AOI22_X1 U5127 ( .A1(n4728), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4581) );
  AOI22_X1 U5128 ( .A1(n4727), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4580) );
  AOI22_X1 U5129 ( .A1(n4655), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4579) );
  AOI22_X1 U5130 ( .A1(n3892), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4578) );
  NAND4_X1 U5131 ( .A1(n4581), .A2(n4580), .A3(n4579), .A4(n4578), .ZN(n4587)
         );
  AOI22_X1 U5132 ( .A1(n3666), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4585) );
  AOI22_X1 U5133 ( .A1(n4732), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4584) );
  AOI22_X1 U5134 ( .A1(n3660), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4583) );
  AOI22_X1 U5135 ( .A1(n4729), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4582) );
  NAND4_X1 U5136 ( .A1(n4585), .A2(n4584), .A3(n4583), .A4(n4582), .ZN(n4586)
         );
  OR2_X1 U5137 ( .A1(n4587), .A2(n4586), .ZN(n4588) );
  NAND2_X1 U5138 ( .A1(n4588), .A2(n4589), .ZN(n4628) );
  OAI21_X1 U5139 ( .B1(n4589), .B2(n4588), .A(n4628), .ZN(n4593) );
  NAND2_X1 U5140 ( .A1(n7584), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4590)
         );
  NAND2_X1 U5141 ( .A1(n4284), .A2(n4590), .ZN(n4591) );
  AOI21_X1 U5142 ( .B1(n4749), .B2(EAX_REG_23__SCAN_IN), .A(n4591), .ZN(n4592)
         );
  OAI21_X1 U5143 ( .B1(n4691), .B2(n4593), .A(n4592), .ZN(n4594) );
  XNOR2_X1 U5144 ( .A(n4596), .B(n6671), .ZN(n6872) );
  AOI22_X1 U5145 ( .A1(n4727), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4729), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4600) );
  AOI22_X1 U5146 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n3665), .B1(n4732), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4599) );
  AOI22_X1 U5147 ( .A1(n4728), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4598) );
  AOI22_X1 U5148 ( .A1(n4718), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4597) );
  NAND4_X1 U5149 ( .A1(n4600), .A2(n4599), .A3(n4598), .A4(n4597), .ZN(n4606)
         );
  AOI22_X1 U5150 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n3660), .B1(n3879), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4604) );
  AOI22_X1 U5151 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n4731), .B1(n4719), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4603) );
  AOI22_X1 U5152 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n4721), .B1(n4720), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4602) );
  AOI22_X1 U5153 ( .A1(n4722), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4601) );
  NAND4_X1 U5154 ( .A1(n4604), .A2(n4603), .A3(n4602), .A4(n4601), .ZN(n4605)
         );
  NOR2_X1 U5155 ( .A1(n4606), .A2(n4605), .ZN(n4629) );
  XNOR2_X1 U5156 ( .A(n4628), .B(n4629), .ZN(n4610) );
  NOR2_X1 U5157 ( .A1(n4607), .A2(n6671), .ZN(n4608) );
  AOI21_X1 U5158 ( .B1(n4749), .B2(EAX_REG_24__SCAN_IN), .A(n4608), .ZN(n4609)
         );
  OAI21_X1 U5159 ( .B1(n4691), .B2(n4610), .A(n4609), .ZN(n4611) );
  AOI21_X1 U5160 ( .B1(n6872), .B2(n4267), .A(n4611), .ZN(n6667) );
  INV_X1 U5161 ( .A(n4614), .ZN(n4616) );
  INV_X1 U5162 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4615) );
  NAND2_X1 U5163 ( .A1(n4616), .A2(n4615), .ZN(n4617) );
  NAND2_X1 U5164 ( .A1(n4636), .A2(n4617), .ZN(n6857) );
  AOI22_X1 U5165 ( .A1(n4728), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4621) );
  AOI22_X1 U5166 ( .A1(n4727), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4620) );
  AOI22_X1 U5167 ( .A1(n4721), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4720), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4619) );
  AOI22_X1 U5168 ( .A1(n3892), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4618) );
  NAND4_X1 U5169 ( .A1(n4621), .A2(n4620), .A3(n4619), .A4(n4618), .ZN(n4627)
         );
  AOI22_X1 U5170 ( .A1(n3665), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4625) );
  AOI22_X1 U5171 ( .A1(n4732), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4624) );
  AOI22_X1 U5172 ( .A1(n3850), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4623) );
  AOI22_X1 U5173 ( .A1(n4702), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4622) );
  NAND4_X1 U5174 ( .A1(n4625), .A2(n4624), .A3(n4623), .A4(n4622), .ZN(n4626)
         );
  OR2_X1 U5175 ( .A1(n4627), .A2(n4626), .ZN(n4647) );
  NOR2_X1 U5176 ( .A1(n4629), .A2(n4628), .ZN(n4648) );
  XNOR2_X1 U5177 ( .A(n4647), .B(n4648), .ZN(n4633) );
  NAND2_X1 U5178 ( .A1(n7584), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4630)
         );
  NAND2_X1 U5179 ( .A1(n4284), .A2(n4630), .ZN(n4631) );
  AOI21_X1 U5180 ( .B1(n4749), .B2(EAX_REG_25__SCAN_IN), .A(n4631), .ZN(n4632)
         );
  OAI21_X1 U5181 ( .B1(n4691), .B2(n4633), .A(n4632), .ZN(n4634) );
  NAND2_X1 U5182 ( .A1(n4635), .A2(n4634), .ZN(n6650) );
  XNOR2_X1 U5183 ( .A(n4636), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6849)
         );
  AOI22_X1 U5184 ( .A1(n4721), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4640) );
  AOI22_X1 U5185 ( .A1(n4732), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4639) );
  AOI22_X1 U5186 ( .A1(n3660), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4638) );
  AOI22_X1 U5187 ( .A1(n3864), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4637) );
  NAND4_X1 U5188 ( .A1(n4640), .A2(n4639), .A3(n4638), .A4(n4637), .ZN(n4646)
         );
  AOI22_X1 U5189 ( .A1(n3665), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4644) );
  AOI22_X1 U5190 ( .A1(n4727), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4643) );
  AOI22_X1 U5191 ( .A1(n4718), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4722), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4642) );
  AOI22_X1 U5192 ( .A1(n4702), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4641) );
  NAND4_X1 U5193 ( .A1(n4644), .A2(n4643), .A3(n4642), .A4(n4641), .ZN(n4645)
         );
  NOR2_X1 U5194 ( .A1(n4646), .A2(n4645), .ZN(n4667) );
  NAND2_X1 U5195 ( .A1(n4648), .A2(n4647), .ZN(n4666) );
  XOR2_X1 U5196 ( .A(n4667), .B(n4666), .Z(n4651) );
  NAND2_X1 U5197 ( .A1(n4749), .A2(EAX_REG_26__SCAN_IN), .ZN(n4649) );
  OAI211_X1 U5198 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6845), .A(n4649), .B(
        n4284), .ZN(n4650) );
  AOI21_X1 U5199 ( .B1(n4651), .B2(n4744), .A(n4650), .ZN(n4652) );
  AOI21_X1 U5200 ( .B1(n6849), .B2(n4267), .A(n4652), .ZN(n6637) );
  NAND2_X1 U5201 ( .A1(n4653), .A2(n6835), .ZN(n4654) );
  AOI22_X1 U5202 ( .A1(n4655), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4659) );
  AOI22_X1 U5203 ( .A1(n4728), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4658) );
  AOI22_X1 U5204 ( .A1(n3666), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4657) );
  AOI22_X1 U5205 ( .A1(n4720), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4656) );
  NAND4_X1 U5206 ( .A1(n4659), .A2(n4658), .A3(n4657), .A4(n4656), .ZN(n4665)
         );
  AOI22_X1 U5207 ( .A1(n3660), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4731), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4663) );
  AOI22_X1 U5208 ( .A1(n3865), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4662) );
  AOI22_X1 U5209 ( .A1(n4727), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3892), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4661) );
  AOI22_X1 U5210 ( .A1(n4702), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4660) );
  NAND4_X1 U5211 ( .A1(n4663), .A2(n4662), .A3(n4661), .A4(n4660), .ZN(n4664)
         );
  OR2_X1 U5212 ( .A1(n4665), .A2(n4664), .ZN(n4677) );
  NOR2_X1 U5213 ( .A1(n4667), .A2(n4666), .ZN(n4676) );
  XOR2_X1 U5214 ( .A(n4677), .B(n4676), .Z(n4671) );
  INV_X1 U5215 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4669) );
  NAND2_X1 U5216 ( .A1(n7584), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4668)
         );
  OAI211_X1 U5217 ( .C1(n4713), .C2(n4669), .A(n4284), .B(n4668), .ZN(n4670)
         );
  AOI21_X1 U5218 ( .B1(n4671), .B2(n4744), .A(n4670), .ZN(n4672) );
  AOI21_X1 U5219 ( .B1(n6837), .B2(n4267), .A(n4672), .ZN(n6626) );
  INV_X1 U5220 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4673) );
  NAND2_X1 U5221 ( .A1(n4674), .A2(n4673), .ZN(n4675) );
  NAND2_X1 U5222 ( .A1(n4696), .A2(n4675), .ZN(n6620) );
  NAND2_X1 U5223 ( .A1(n4677), .A2(n4676), .ZN(n4740) );
  AOI22_X1 U5224 ( .A1(n4728), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4718), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4681) );
  AOI22_X1 U5225 ( .A1(n4731), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4680) );
  AOI22_X1 U5226 ( .A1(n3892), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4679) );
  AOI22_X1 U5227 ( .A1(n4702), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4678) );
  NAND4_X1 U5228 ( .A1(n4681), .A2(n4680), .A3(n4679), .A4(n4678), .ZN(n4687)
         );
  AOI22_X1 U5229 ( .A1(n4727), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4685) );
  AOI22_X1 U5230 ( .A1(n3660), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3665), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4684) );
  AOI22_X1 U5231 ( .A1(n4732), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4683) );
  AOI22_X1 U5232 ( .A1(n4721), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4682) );
  NAND4_X1 U5233 ( .A1(n4685), .A2(n4684), .A3(n4683), .A4(n4682), .ZN(n4686)
         );
  NOR2_X1 U5234 ( .A1(n4687), .A2(n4686), .ZN(n4739) );
  XNOR2_X1 U5235 ( .A(n4740), .B(n4739), .ZN(n4692) );
  NAND2_X1 U5236 ( .A1(n7584), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4688)
         );
  NAND2_X1 U5237 ( .A1(n4284), .A2(n4688), .ZN(n4689) );
  AOI21_X1 U5238 ( .B1(n4749), .B2(EAX_REG_28__SCAN_IN), .A(n4689), .ZN(n4690)
         );
  OAI21_X1 U5239 ( .B1(n4692), .B2(n4691), .A(n4690), .ZN(n4693) );
  NAND2_X1 U5240 ( .A1(n4694), .A2(n4693), .ZN(n6527) );
  NAND2_X1 U5241 ( .A1(n4696), .A2(n4695), .ZN(n4697) );
  NAND2_X1 U5242 ( .A1(n4716), .A2(n4697), .ZN(n6610) );
  NOR2_X1 U5243 ( .A1(n4740), .A2(n4739), .ZN(n4709) );
  AOI22_X1 U5244 ( .A1(n4721), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4701) );
  AOI22_X1 U5245 ( .A1(n4732), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4700) );
  AOI22_X1 U5246 ( .A1(n3660), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4699) );
  AOI22_X1 U5247 ( .A1(n4731), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4698) );
  NAND4_X1 U5248 ( .A1(n4701), .A2(n4700), .A3(n4699), .A4(n4698), .ZN(n4708)
         );
  AOI22_X1 U5249 ( .A1(n3666), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4702), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4706) );
  AOI22_X1 U5250 ( .A1(n4727), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3879), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4705) );
  AOI22_X1 U5251 ( .A1(n4718), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4704) );
  AOI22_X1 U5252 ( .A1(n4722), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4703) );
  NAND4_X1 U5253 ( .A1(n4706), .A2(n4705), .A3(n4704), .A4(n4703), .ZN(n4707)
         );
  NOR2_X1 U5254 ( .A1(n4708), .A2(n4707), .ZN(n4741) );
  XNOR2_X1 U5255 ( .A(n4709), .B(n4741), .ZN(n4710) );
  AND2_X1 U5256 ( .A1(n4710), .A2(n4744), .ZN(n4715) );
  INV_X1 U5257 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4712) );
  NAND2_X1 U5258 ( .A1(n7584), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4711)
         );
  OAI211_X1 U5259 ( .C1(n4713), .C2(n4712), .A(n4284), .B(n4711), .ZN(n4714)
         );
  OAI22_X1 U5260 ( .A1(n6610), .A2(n4284), .B1(n4715), .B2(n4714), .ZN(n6557)
         );
  NOR2_X4 U5261 ( .A1(n6558), .A2(n6557), .ZN(n6556) );
  XNOR2_X1 U5262 ( .A(n4716), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4967)
         );
  INV_X1 U5263 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4952) );
  NOR2_X1 U5264 ( .A1(n4952), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4717) );
  AOI211_X1 U5265 ( .C1(n4749), .C2(EAX_REG_30__SCAN_IN), .A(n4267), .B(n4717), 
        .ZN(n4747) );
  AOI22_X1 U5266 ( .A1(n4718), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4726) );
  AOI22_X1 U5267 ( .A1(n3660), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4719), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4725) );
  AOI22_X1 U5268 ( .A1(n4721), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4720), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4724) );
  AOI22_X1 U5269 ( .A1(n4722), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4723) );
  NAND4_X1 U5270 ( .A1(n4726), .A2(n4725), .A3(n4724), .A4(n4723), .ZN(n4738)
         );
  AOI22_X1 U5271 ( .A1(n4728), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4727), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4736) );
  AOI22_X1 U5272 ( .A1(n3665), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4729), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4735) );
  AOI22_X1 U5273 ( .A1(n4731), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4730), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4734) );
  AOI22_X1 U5274 ( .A1(n4732), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4539), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4733) );
  NAND4_X1 U5275 ( .A1(n4736), .A2(n4735), .A3(n4734), .A4(n4733), .ZN(n4737)
         );
  NOR2_X1 U5276 ( .A1(n4738), .A2(n4737), .ZN(n4743) );
  NOR3_X1 U5277 ( .A1(n4741), .A2(n4740), .A3(n4739), .ZN(n4742) );
  XNOR2_X1 U5278 ( .A(n4743), .B(n4742), .ZN(n4745) );
  NAND2_X1 U5279 ( .A1(n4745), .A2(n4744), .ZN(n4746) );
  AOI22_X1 U5280 ( .A1(n4967), .A2(n4267), .B1(n4747), .B2(n4746), .ZN(n4950)
         );
  NAND2_X1 U5281 ( .A1(n6556), .A2(n4950), .ZN(n4752) );
  AOI22_X1 U5282 ( .A1(n4749), .A2(EAX_REG_31__SCAN_IN), .B1(n4748), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4750) );
  INV_X1 U5283 ( .A(n4750), .ZN(n4751) );
  XNOR2_X2 U5284 ( .A(n4752), .B(n4751), .ZN(n6797) );
  NAND3_X1 U5285 ( .A1(n7318), .A2(STATE2_REG_1__SCAN_IN), .A3(
        STATEBS16_REG_SCAN_IN), .ZN(n7314) );
  INV_X1 U5286 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6995) );
  NAND2_X1 U5287 ( .A1(n4171), .A2(n6995), .ZN(n6855) );
  NOR3_X1 U5288 ( .A1(n6843), .A2(n6842), .A3(n4941), .ZN(n4755) );
  INV_X1 U5289 ( .A(n4754), .ZN(n6543) );
  OAI21_X1 U5290 ( .B1(n4755), .B2(n6543), .A(n6539), .ZN(n4756) );
  NAND2_X1 U5291 ( .A1(n3924), .A2(n7131), .ZN(n4764) );
  NOR3_X1 U5292 ( .A1(n4759), .A2(n4758), .A3(n4757), .ZN(n4762) );
  OAI21_X1 U5293 ( .B1(n4762), .B2(n4761), .A(n4760), .ZN(n6586) );
  NAND2_X1 U5294 ( .A1(n7634), .A2(n6586), .ZN(n5013) );
  INV_X1 U5295 ( .A(n5013), .ZN(n4763) );
  NAND2_X1 U5296 ( .A1(n4764), .A2(n4763), .ZN(n4766) );
  OAI21_X1 U5297 ( .B1(n5140), .B2(n4256), .A(n6593), .ZN(n4765) );
  MUX2_X1 U5298 ( .A(n4766), .B(n4765), .S(n3906), .Z(n4781) );
  AOI21_X1 U5299 ( .B1(n5228), .B2(n7131), .A(READY_N), .ZN(n4767) );
  NAND2_X1 U5300 ( .A1(n6593), .A2(n4767), .ZN(n5016) );
  NOR2_X1 U5301 ( .A1(n5043), .A2(n5228), .ZN(n4898) );
  NAND2_X1 U5302 ( .A1(n5026), .A2(n4898), .ZN(n4778) );
  NAND2_X1 U5303 ( .A1(n4770), .A2(n4771), .ZN(n4958) );
  INV_X1 U5304 ( .A(n5094), .ZN(n4772) );
  OR2_X1 U5305 ( .A1(n4773), .A2(n4772), .ZN(n4776) );
  NAND2_X1 U5306 ( .A1(n5094), .A2(n3941), .ZN(n4774) );
  NAND2_X1 U5307 ( .A1(n6594), .A2(n4774), .ZN(n4775) );
  NAND2_X1 U5308 ( .A1(n4776), .A2(n4775), .ZN(n4890) );
  NAND2_X1 U5309 ( .A1(n4786), .A2(n4890), .ZN(n4777) );
  NAND2_X1 U5310 ( .A1(n4958), .A2(n4777), .ZN(n5021) );
  OAI211_X1 U5311 ( .C1(n5016), .C2(n4769), .A(n4778), .B(n5021), .ZN(n4779)
         );
  INV_X1 U5312 ( .A(n4779), .ZN(n4780) );
  NAND2_X1 U5313 ( .A1(n4781), .A2(n4780), .ZN(n4782) );
  OAI22_X1 U5314 ( .A1(n4769), .A2(n5075), .B1(n3940), .B2(n4784), .ZN(n4785)
         );
  NOR2_X1 U5315 ( .A1(n6583), .A2(n4785), .ZN(n4788) );
  AND2_X1 U5316 ( .A1(n4786), .A2(n5088), .ZN(n6584) );
  INV_X1 U5317 ( .A(n6584), .ZN(n4787) );
  NAND3_X1 U5318 ( .A1(n4783), .A2(n4788), .A3(n4787), .ZN(n4789) );
  MUX2_X1 U5319 ( .A(n4795), .B(n4932), .S(EBX_REG_1__SCAN_IN), .Z(n4791) );
  INV_X1 U5320 ( .A(n3923), .ZN(n5215) );
  AND2_X2 U5321 ( .A1(n4932), .A2(n4871), .ZN(n5051) );
  NAND2_X1 U5322 ( .A1(n5051), .A2(n4078), .ZN(n4790) );
  INV_X1 U5323 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4793) );
  NAND2_X1 U5324 ( .A1(n4874), .A2(n4793), .ZN(n4792) );
  OAI21_X1 U5325 ( .B1(n4871), .B2(n4793), .A(n4792), .ZN(n5050) );
  MUX2_X1 U5326 ( .A(n4795), .B(n4932), .S(EBX_REG_2__SCAN_IN), .Z(n4797) );
  NAND2_X1 U5327 ( .A1(n5051), .A2(n7349), .ZN(n4796) );
  AND2_X1 U5328 ( .A1(n4797), .A2(n4796), .ZN(n5115) );
  NAND2_X1 U5329 ( .A1(n4871), .A2(n7102), .ZN(n4799) );
  INV_X1 U5330 ( .A(EBX_REG_3__SCAN_IN), .ZN(n7439) );
  NAND2_X1 U5331 ( .A1(n5085), .A2(n7439), .ZN(n4798) );
  NAND3_X1 U5332 ( .A1(n4799), .A2(n4932), .A3(n4798), .ZN(n4801) );
  NAND2_X1 U5333 ( .A1(n4874), .A2(n7439), .ZN(n4800) );
  AND2_X1 U5334 ( .A1(n4801), .A2(n4800), .ZN(n5720) );
  MUX2_X1 U5335 ( .A(n4795), .B(n4932), .S(EBX_REG_4__SCAN_IN), .Z(n4802) );
  OAI21_X1 U5336 ( .B1(INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n4931), .A(n4802), 
        .ZN(n5110) );
  NAND2_X1 U5337 ( .A1(n4871), .A2(n6438), .ZN(n4804) );
  INV_X1 U5338 ( .A(EBX_REG_5__SCAN_IN), .ZN(n7470) );
  NAND2_X1 U5339 ( .A1(n5085), .A2(n7470), .ZN(n4803) );
  NAND3_X1 U5340 ( .A1(n4804), .A2(n4932), .A3(n4803), .ZN(n4806) );
  NAND2_X1 U5341 ( .A1(n4874), .A2(n7470), .ZN(n4805) );
  NAND2_X1 U5342 ( .A1(n4806), .A2(n4805), .ZN(n5651) );
  MUX2_X1 U5343 ( .A(n4795), .B(n4932), .S(EBX_REG_6__SCAN_IN), .Z(n4808) );
  NAND2_X1 U5344 ( .A1(n5051), .A2(n6440), .ZN(n4807) );
  AND2_X1 U5345 ( .A1(n4808), .A2(n4807), .ZN(n5154) );
  INV_X1 U5346 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4809) );
  NAND2_X1 U5347 ( .A1(n4871), .A2(n4809), .ZN(n4811) );
  INV_X1 U5348 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5705) );
  NAND2_X1 U5349 ( .A1(n5085), .A2(n5705), .ZN(n4810) );
  NAND3_X1 U5350 ( .A1(n4811), .A2(n4932), .A3(n4810), .ZN(n4813) );
  NAND2_X1 U5351 ( .A1(n4874), .A2(n5705), .ZN(n4812) );
  AND2_X1 U5352 ( .A1(n4813), .A2(n4812), .ZN(n5701) );
  MUX2_X1 U5353 ( .A(n4795), .B(n4932), .S(EBX_REG_8__SCAN_IN), .Z(n4814) );
  OAI21_X1 U5354 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n4931), .A(n4814), 
        .ZN(n5150) );
  INV_X1 U5355 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4901) );
  NAND2_X1 U5356 ( .A1(n4871), .A2(n4901), .ZN(n4816) );
  INV_X1 U5357 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5815) );
  NAND2_X1 U5358 ( .A1(n5085), .A2(n5815), .ZN(n4815) );
  NAND3_X1 U5359 ( .A1(n4816), .A2(n4932), .A3(n4815), .ZN(n4818) );
  NAND2_X1 U5360 ( .A1(n4874), .A2(n5815), .ZN(n4817) );
  NAND2_X1 U5361 ( .A1(n4818), .A2(n4817), .ZN(n5812) );
  MUX2_X1 U5362 ( .A(n4795), .B(n4932), .S(EBX_REG_10__SCAN_IN), .Z(n4820) );
  NAND2_X1 U5363 ( .A1(n5051), .A2(n4173), .ZN(n4819) );
  AND2_X1 U5364 ( .A1(n4820), .A2(n4819), .ZN(n5838) );
  NAND2_X1 U5365 ( .A1(n4871), .A2(n4174), .ZN(n4822) );
  INV_X1 U5366 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5853) );
  NAND2_X1 U5367 ( .A1(n5085), .A2(n5853), .ZN(n4821) );
  NAND3_X1 U5368 ( .A1(n4822), .A2(n4932), .A3(n4821), .ZN(n4824) );
  NAND2_X1 U5369 ( .A1(n4874), .A2(n5853), .ZN(n4823) );
  INV_X1 U5370 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U5371 ( .A1(n5085), .A2(n6458), .ZN(n4825) );
  OAI211_X1 U5372 ( .C1(n4874), .C2(n4172), .A(n4825), .B(n4871), .ZN(n4826)
         );
  OAI21_X1 U5373 ( .B1(n4795), .B2(EBX_REG_12__SCAN_IN), .A(n4826), .ZN(n6450)
         );
  INV_X1 U5374 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n7092) );
  NAND2_X1 U5375 ( .A1(n4871), .A2(n7092), .ZN(n4828) );
  INV_X1 U5376 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U5377 ( .A1(n5085), .A2(n6487), .ZN(n4827) );
  NAND3_X1 U5378 ( .A1(n4828), .A2(n4932), .A3(n4827), .ZN(n4830) );
  NAND2_X1 U5379 ( .A1(n4874), .A2(n6487), .ZN(n4829) );
  MUX2_X1 U5380 ( .A(n4795), .B(n4932), .S(EBX_REG_14__SCAN_IN), .Z(n4832) );
  NAND2_X1 U5381 ( .A1(n5051), .A2(n7330), .ZN(n4831) );
  NAND2_X1 U5382 ( .A1(n6503), .A2(n6502), .ZN(n6745) );
  NAND2_X1 U5383 ( .A1(n4871), .A2(n7401), .ZN(n4834) );
  INV_X1 U5384 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6791) );
  NAND2_X1 U5385 ( .A1(n5085), .A2(n6791), .ZN(n4833) );
  NAND3_X1 U5386 ( .A1(n4834), .A2(n4932), .A3(n4833), .ZN(n4836) );
  NAND2_X1 U5387 ( .A1(n4874), .A2(n6791), .ZN(n4835) );
  MUX2_X1 U5388 ( .A(n4795), .B(n4932), .S(EBX_REG_16__SCAN_IN), .Z(n4838) );
  NAND2_X1 U5389 ( .A1(n5051), .A2(n7408), .ZN(n4837) );
  NAND2_X1 U5390 ( .A1(n4838), .A2(n4837), .ZN(n6732) );
  OAI21_X1 U5391 ( .B1(n4874), .B2(n7073), .A(n4871), .ZN(n4840) );
  INV_X1 U5392 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6786) );
  NAND2_X1 U5393 ( .A1(n5085), .A2(n6786), .ZN(n4839) );
  NAND2_X1 U5394 ( .A1(n4840), .A2(n4839), .ZN(n4842) );
  NAND2_X1 U5395 ( .A1(n4874), .A2(n6786), .ZN(n4841) );
  NAND2_X1 U5396 ( .A1(n4842), .A2(n4841), .ZN(n6784) );
  MUX2_X1 U5397 ( .A(n4795), .B(n4932), .S(EBX_REG_18__SCAN_IN), .Z(n4844) );
  NAND2_X1 U5398 ( .A1(n5051), .A2(n7423), .ZN(n4843) );
  NAND2_X1 U5399 ( .A1(n4844), .A2(n4843), .ZN(n6723) );
  INV_X1 U5400 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n7044) );
  OAI21_X1 U5401 ( .B1(n4874), .B2(n7044), .A(n4871), .ZN(n4846) );
  INV_X1 U5402 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6778) );
  NAND2_X1 U5403 ( .A1(n5085), .A2(n6778), .ZN(n4845) );
  AOI22_X1 U5404 ( .A1(n4846), .A2(n4845), .B1(n4874), .B2(n6778), .ZN(n6774)
         );
  INV_X1 U5405 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4848) );
  INV_X1 U5406 ( .A(EBX_REG_20__SCAN_IN), .ZN(n6768) );
  NAND2_X1 U5407 ( .A1(n5085), .A2(n6768), .ZN(n4847) );
  OAI211_X1 U5408 ( .C1(n4874), .C2(n4848), .A(n4847), .B(n4871), .ZN(n4849)
         );
  OAI21_X1 U5409 ( .B1(n4795), .B2(EBX_REG_20__SCAN_IN), .A(n4849), .ZN(n6707)
         );
  INV_X1 U5410 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n7040) );
  OAI21_X1 U5411 ( .B1(n4874), .B2(n7040), .A(n4871), .ZN(n4851) );
  INV_X1 U5412 ( .A(EBX_REG_21__SCAN_IN), .ZN(n6767) );
  NAND2_X1 U5413 ( .A1(n5085), .A2(n6767), .ZN(n4850) );
  AOI22_X1 U5414 ( .A1(n4851), .A2(n4850), .B1(n4874), .B2(n6767), .ZN(n6698)
         );
  MUX2_X1 U5415 ( .A(n4795), .B(n4932), .S(EBX_REG_22__SCAN_IN), .Z(n4853) );
  INV_X1 U5416 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n7024) );
  NAND2_X1 U5417 ( .A1(n5051), .A2(n7024), .ZN(n4852) );
  MUX2_X1 U5418 ( .A(n4795), .B(n4932), .S(EBX_REG_24__SCAN_IN), .Z(n4856) );
  INV_X1 U5419 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4854) );
  NAND2_X1 U5420 ( .A1(n5051), .A2(n4854), .ZN(n4855) );
  NAND2_X1 U5421 ( .A1(n4856), .A2(n4855), .ZN(n6674) );
  INV_X1 U5422 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n7016) );
  NAND2_X1 U5423 ( .A1(n4871), .A2(n7016), .ZN(n4858) );
  INV_X1 U5424 ( .A(EBX_REG_23__SCAN_IN), .ZN(n7530) );
  NAND2_X1 U5425 ( .A1(n5085), .A2(n7530), .ZN(n4857) );
  NAND3_X1 U5426 ( .A1(n4858), .A2(n4932), .A3(n4857), .ZN(n4860) );
  NAND2_X1 U5427 ( .A1(n4874), .A2(n7530), .ZN(n4859) );
  AND2_X1 U5428 ( .A1(n4860), .A2(n4859), .ZN(n6673) );
  NOR2_X1 U5429 ( .A1(n6674), .A2(n6673), .ZN(n4861) );
  NAND2_X1 U5430 ( .A1(n4871), .A2(n6995), .ZN(n4863) );
  INV_X1 U5431 ( .A(EBX_REG_25__SCAN_IN), .ZN(n6764) );
  NAND2_X1 U5432 ( .A1(n5085), .A2(n6764), .ZN(n4862) );
  NAND3_X1 U5433 ( .A1(n4863), .A2(n4932), .A3(n4862), .ZN(n4865) );
  NAND2_X1 U5434 ( .A1(n4874), .A2(n6764), .ZN(n4864) );
  NAND2_X1 U5435 ( .A1(n4865), .A2(n4864), .ZN(n6653) );
  MUX2_X1 U5436 ( .A(n4795), .B(n4932), .S(EBX_REG_26__SCAN_IN), .Z(n4867) );
  NAND2_X1 U5437 ( .A1(n5051), .A2(n6842), .ZN(n4866) );
  NAND2_X1 U5438 ( .A1(n4867), .A2(n4866), .ZN(n6639) );
  OAI21_X1 U5439 ( .B1(n4874), .B2(n6986), .A(n4871), .ZN(n4869) );
  INV_X1 U5440 ( .A(EBX_REG_27__SCAN_IN), .ZN(n6762) );
  NAND2_X1 U5441 ( .A1(n5085), .A2(n6762), .ZN(n4868) );
  AOI22_X1 U5442 ( .A1(n4869), .A2(n4868), .B1(n4874), .B2(n6762), .ZN(n6624)
         );
  NOR2_X2 U5443 ( .A1(n6641), .A2(n6624), .ZN(n6533) );
  INV_X1 U5444 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4870) );
  NAND2_X1 U5445 ( .A1(n4871), .A2(n4870), .ZN(n4873) );
  INV_X1 U5446 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6761) );
  NAND2_X1 U5447 ( .A1(n5085), .A2(n6761), .ZN(n4872) );
  NAND3_X1 U5448 ( .A1(n4873), .A2(n4932), .A3(n4872), .ZN(n4876) );
  NAND2_X1 U5449 ( .A1(n4874), .A2(n6761), .ZN(n4875) );
  NAND2_X1 U5450 ( .A1(n4876), .A2(n4875), .ZN(n6532) );
  INV_X1 U5451 ( .A(EBX_REG_29__SCAN_IN), .ZN(n6759) );
  AND2_X1 U5452 ( .A1(n5085), .A2(n6759), .ZN(n4877) );
  INV_X1 U5453 ( .A(n4877), .ZN(n4934) );
  OAI21_X1 U5454 ( .B1(n4931), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n4934), 
        .ZN(n4933) );
  INV_X1 U5455 ( .A(n4933), .ZN(n4878) );
  AND2_X1 U5456 ( .A1(n6546), .A2(n4878), .ZN(n4879) );
  AOI22_X1 U5457 ( .A1(n4931), .A2(EBX_REG_30__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5075), .ZN(n4935) );
  INV_X1 U5458 ( .A(n4935), .ZN(n4880) );
  INV_X1 U5459 ( .A(n6579), .ZN(n4883) );
  OAI21_X1 U5460 ( .B1(n4784), .B2(n5177), .A(n7554), .ZN(n4882) );
  NAND2_X1 U5461 ( .A1(n4883), .A2(n7418), .ZN(n4929) );
  INV_X1 U5462 ( .A(n4884), .ZN(n4889) );
  AND2_X1 U5463 ( .A1(n4889), .A2(n4885), .ZN(n4886) );
  NAND2_X1 U5464 ( .A1(n4899), .A2(n5317), .ZN(n5060) );
  NAND2_X1 U5465 ( .A1(n4236), .A2(n4931), .ZN(n4892) );
  NAND2_X1 U5466 ( .A1(n4256), .A2(n5140), .ZN(n4888) );
  AOI22_X1 U5467 ( .A1(n4889), .A2(n4887), .B1(n4888), .B2(n3945), .ZN(n4891)
         );
  OAI211_X1 U5468 ( .C1(n5177), .C2(n4896), .A(n5032), .B(n4895), .ZN(n4897)
         );
  NAND2_X1 U5469 ( .A1(n4899), .A2(n4897), .ZN(n5054) );
  AND2_X2 U5470 ( .A1(n5060), .A2(n5054), .ZN(n7062) );
  NAND2_X1 U5471 ( .A1(n7062), .A2(n7079), .ZN(n7340) );
  INV_X1 U5472 ( .A(n7340), .ZN(n7095) );
  INV_X1 U5473 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5059) );
  NAND2_X1 U5474 ( .A1(n5060), .A2(n5059), .ZN(n7341) );
  INV_X1 U5475 ( .A(n7341), .ZN(n4900) );
  INV_X1 U5476 ( .A(n7353), .ZN(n4903) );
  NAND3_X1 U5477 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .ZN(n6437) );
  NOR2_X1 U5478 ( .A1(n6440), .A2(n6437), .ZN(n6474) );
  INV_X1 U5479 ( .A(n6474), .ZN(n4902) );
  NAND2_X1 U5480 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n7362) );
  NAND2_X1 U5481 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5820) );
  NOR2_X1 U5482 ( .A1(n4173), .A2(n4901), .ZN(n7061) );
  INV_X1 U5483 ( .A(n7061), .ZN(n7378) );
  NOR4_X1 U5484 ( .A1(n4902), .A2(n7362), .A3(n5820), .A4(n7378), .ZN(n4908)
         );
  NAND2_X1 U5485 ( .A1(n4903), .A2(n4908), .ZN(n7384) );
  OAI21_X1 U5486 ( .B1(n4078), .B2(n5059), .A(n7349), .ZN(n7345) );
  NAND2_X1 U5487 ( .A1(n6474), .A2(n7345), .ZN(n7359) );
  NOR2_X1 U5488 ( .A1(n7362), .A2(n7359), .ZN(n6475) );
  NAND2_X1 U5489 ( .A1(n7061), .A2(n6475), .ZN(n7077) );
  NAND2_X1 U5490 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n7385) );
  NOR2_X1 U5491 ( .A1(n7092), .A2(n7385), .ZN(n7331) );
  NAND2_X1 U5492 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n7331), .ZN(n7400) );
  NOR3_X1 U5493 ( .A1(n7408), .A2(n7401), .A3(n7400), .ZN(n7059) );
  NAND2_X1 U5494 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n7059), .ZN(n7413) );
  NOR2_X1 U5495 ( .A1(n7423), .A2(n7413), .ZN(n4907) );
  NAND2_X1 U5496 ( .A1(n7383), .A2(n4907), .ZN(n7056) );
  INV_X1 U5497 ( .A(n7056), .ZN(n4906) );
  INV_X1 U5498 ( .A(n4905), .ZN(n7023) );
  NAND2_X1 U5499 ( .A1(n4906), .A2(n7023), .ZN(n7045) );
  AOI21_X1 U5500 ( .B1(n4908), .B2(n4907), .A(n7062), .ZN(n4915) );
  OR2_X1 U5501 ( .A1(n5054), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4910)
         );
  NAND2_X1 U5502 ( .A1(n7088), .A2(n4909), .ZN(n7336) );
  NAND2_X1 U5503 ( .A1(n4910), .A2(n7336), .ZN(n5819) );
  INV_X1 U5504 ( .A(n5819), .ZN(n4913) );
  INV_X1 U5505 ( .A(n7079), .ZN(n7386) );
  NOR2_X1 U5506 ( .A1(n7077), .A2(n7413), .ZN(n7065) );
  NAND2_X1 U5507 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n7065), .ZN(n4911) );
  NAND2_X1 U5508 ( .A1(n7386), .A2(n4911), .ZN(n4912) );
  NAND2_X1 U5509 ( .A1(n4913), .A2(n4912), .ZN(n4914) );
  INV_X1 U5510 ( .A(n7053), .ZN(n4916) );
  NAND2_X1 U5511 ( .A1(n7045), .A2(n4916), .ZN(n7048) );
  INV_X1 U5512 ( .A(n4917), .ZN(n4918) );
  AND2_X1 U5513 ( .A1(n7340), .A2(n4918), .ZN(n4919) );
  OR2_X2 U5514 ( .A1(n7048), .A2(n4919), .ZN(n7020) );
  INV_X1 U5515 ( .A(n4920), .ZN(n4924) );
  AOI21_X1 U5516 ( .B1(n7353), .B2(n7079), .A(n4924), .ZN(n4921) );
  NOR2_X1 U5517 ( .A1(n7020), .A2(n4921), .ZN(n7006) );
  NAND2_X1 U5518 ( .A1(n7340), .A2(n6988), .ZN(n4922) );
  NAND2_X1 U5519 ( .A1(n7006), .A2(n4922), .ZN(n6977) );
  AND2_X1 U5520 ( .A1(n7340), .A2(n6540), .ZN(n4923) );
  NOR2_X1 U5521 ( .A1(n6977), .A2(n4923), .ZN(n6553) );
  OAI21_X1 U5522 ( .B1(n7095), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n6553), 
        .ZN(n4939) );
  NAND2_X1 U5523 ( .A1(n7370), .A2(REIP_REG_30__SCAN_IN), .ZN(n4951) );
  INV_X1 U5524 ( .A(n4951), .ZN(n4927) );
  INV_X1 U5525 ( .A(n6988), .ZN(n4925) );
  INV_X1 U5526 ( .A(n6549), .ZN(n6981) );
  NOR3_X1 U5527 ( .A1(n6981), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n4941), 
        .ZN(n4926) );
  AOI211_X1 U5528 ( .C1(n4939), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n4927), .B(n4926), .ZN(n4928) );
  OAI21_X1 U5529 ( .B1(n4955), .B2(n7350), .A(n4930), .ZN(U2988) );
  AOI22_X1 U5530 ( .A1(n4931), .A2(EBX_REG_31__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5075), .ZN(n4938) );
  MUX2_X1 U5531 ( .A(n4934), .B(n4933), .S(n4932), .Z(n6547) );
  NOR2_X1 U5532 ( .A1(n6547), .A2(n4935), .ZN(n4937) );
  AOI21_X1 U5533 ( .B1(n7340), .B2(n4940), .A(n4939), .ZN(n4946) );
  INV_X1 U5534 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4945) );
  INV_X1 U5535 ( .A(n4941), .ZN(n4942) );
  NAND4_X1 U5536 ( .A1(n6549), .A2(n4942), .A3(INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n4945), .ZN(n4943) );
  OAI211_X1 U5537 ( .C1(n4946), .C2(n4945), .A(n4944), .B(n4943), .ZN(n4947)
         );
  AOI21_X1 U5538 ( .B1(n6755), .B2(n7418), .A(n4947), .ZN(n4948) );
  OAI21_X1 U5539 ( .B1(n4949), .B2(n7350), .A(n4948), .ZN(U2987) );
  OAI21_X1 U5540 ( .B1(n7283), .B2(n4952), .A(n4951), .ZN(n4953) );
  INV_X1 U5541 ( .A(n4958), .ZN(n6588) );
  AND2_X1 U5542 ( .A1(n6588), .A2(n6586), .ZN(n4986) );
  NAND2_X1 U5543 ( .A1(n4986), .A2(n7581), .ZN(n4990) );
  NAND2_X1 U5544 ( .A1(n7584), .A2(n5338), .ZN(n7596) );
  NOR2_X1 U5545 ( .A1(n7318), .A2(n7596), .ZN(n4987) );
  NAND2_X1 U5546 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4987), .ZN(n7603) );
  AND2_X1 U5547 ( .A1(n7318), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4959) );
  NAND2_X1 U5548 ( .A1(n4960), .A2(n4959), .ZN(n7589) );
  NAND2_X1 U5549 ( .A1(n7436), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4964) );
  INV_X1 U5550 ( .A(n6597), .ZN(n4963) );
  NAND2_X1 U5551 ( .A1(n7608), .A2(n7634), .ZN(n4978) );
  AND3_X1 U5552 ( .A1(n5085), .A2(EBX_REG_31__SCAN_IN), .A3(n4978), .ZN(n4962)
         );
  INV_X1 U5553 ( .A(n4964), .ZN(n4965) );
  INV_X1 U5554 ( .A(n4967), .ZN(n4968) );
  AND2_X1 U5555 ( .A1(n3941), .A2(n7311), .ZN(n4969) );
  INV_X1 U5556 ( .A(n4978), .ZN(n4977) );
  OAI21_X1 U5557 ( .B1(n5085), .B2(n4969), .A(n4977), .ZN(n4970) );
  AND2_X1 U5558 ( .A1(n7457), .A2(n7436), .ZN(n7429) );
  INV_X1 U5559 ( .A(n7429), .ZN(n5860) );
  INV_X1 U5560 ( .A(REIP_REG_25__SCAN_IN), .ZN(n7214) );
  INV_X1 U5561 ( .A(REIP_REG_23__SCAN_IN), .ZN(n7526) );
  INV_X1 U5562 ( .A(REIP_REG_19__SCAN_IN), .ZN(n7203) );
  NAND3_X1 U5563 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .ZN(n7456) );
  INV_X1 U5564 ( .A(REIP_REG_4__SCAN_IN), .ZN(n7453) );
  NOR2_X1 U5565 ( .A1(n7456), .A2(n7453), .ZN(n7469) );
  NAND2_X1 U5566 ( .A1(n7469), .A2(REIP_REG_5__SCAN_IN), .ZN(n7467) );
  NAND2_X1 U5567 ( .A1(REIP_REG_6__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .ZN(
        n7491) );
  INV_X1 U5568 ( .A(REIP_REG_8__SCAN_IN), .ZN(n7181) );
  NOR3_X1 U5569 ( .A1(n7467), .A2(n7491), .A3(n7181), .ZN(n6506) );
  NAND2_X1 U5570 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n6492) );
  NAND3_X1 U5571 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_11__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .ZN(n5861) );
  NOR2_X1 U5572 ( .A1(n6492), .A2(n5861), .ZN(n6505) );
  NAND3_X1 U5573 ( .A1(n6506), .A2(n6505), .A3(REIP_REG_14__SCAN_IN), .ZN(
        n6721) );
  INV_X1 U5574 ( .A(REIP_REG_17__SCAN_IN), .ZN(n7199) );
  INV_X1 U5575 ( .A(REIP_REG_16__SCAN_IN), .ZN(n7198) );
  INV_X1 U5576 ( .A(REIP_REG_15__SCAN_IN), .ZN(n7196) );
  NOR3_X1 U5577 ( .A1(n7199), .A2(n7198), .A3(n7196), .ZN(n6722) );
  NAND2_X1 U5578 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6722), .ZN(n7511) );
  NOR3_X1 U5579 ( .A1(n7203), .A2(n6721), .A3(n7511), .ZN(n6710) );
  NAND2_X1 U5580 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6710), .ZN(n6689) );
  NAND2_X1 U5581 ( .A1(REIP_REG_21__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .ZN(
        n7528) );
  NOR3_X1 U5582 ( .A1(n7526), .A2(n6689), .A3(n7528), .ZN(n6669) );
  NAND2_X1 U5583 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6669), .ZN(n6655) );
  NOR2_X1 U5584 ( .A1(n7214), .A2(n6655), .ZN(n6642) );
  NAND2_X1 U5585 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6642), .ZN(n6628) );
  INV_X1 U5586 ( .A(n6628), .ZN(n4974) );
  NAND2_X1 U5587 ( .A1(n7436), .A2(n4974), .ZN(n4971) );
  NAND2_X1 U5588 ( .A1(n5860), .A2(n4971), .ZN(n6644) );
  INV_X1 U5589 ( .A(REIP_REG_28__SCAN_IN), .ZN(n7222) );
  INV_X1 U5590 ( .A(REIP_REG_27__SCAN_IN), .ZN(n7221) );
  OAI21_X1 U5591 ( .B1(n7222), .B2(n7221), .A(n7468), .ZN(n4972) );
  AND2_X1 U5592 ( .A1(n6644), .A2(n4972), .ZN(n6615) );
  INV_X1 U5593 ( .A(REIP_REG_30__SCAN_IN), .ZN(n7227) );
  INV_X1 U5594 ( .A(REIP_REG_29__SCAN_IN), .ZN(n7224) );
  OAI21_X1 U5595 ( .B1(n7227), .B2(n7224), .A(n7468), .ZN(n4973) );
  AND2_X1 U5596 ( .A1(n6615), .A2(n4973), .ZN(n6602) );
  NAND2_X1 U5597 ( .A1(n4974), .A2(REIP_REG_27__SCAN_IN), .ZN(n4975) );
  NOR2_X1 U5598 ( .A1(n7457), .A2(n4975), .ZN(n6617) );
  NAND2_X1 U5599 ( .A1(n6617), .A2(REIP_REG_28__SCAN_IN), .ZN(n6607) );
  INV_X1 U5600 ( .A(n6607), .ZN(n4976) );
  AOI21_X1 U5601 ( .B1(n4976), .B2(REIP_REG_29__SCAN_IN), .A(
        REIP_REG_30__SCAN_IN), .ZN(n4983) );
  NAND2_X1 U5602 ( .A1(n7311), .A2(n4977), .ZN(n7553) );
  NAND2_X1 U5603 ( .A1(n4054), .A2(n7553), .ZN(n6596) );
  INV_X1 U5604 ( .A(EBX_REG_31__SCAN_IN), .ZN(n6756) );
  NAND3_X1 U5605 ( .A1(n3941), .A2(n4978), .A3(n6756), .ZN(n4979) );
  AND2_X1 U5606 ( .A1(n6596), .A2(n4979), .ZN(n4980) );
  NAND2_X1 U5607 ( .A1(n7519), .A2(EBX_REG_30__SCAN_IN), .ZN(n4982) );
  NAND2_X1 U5608 ( .A1(n7501), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4981)
         );
  OAI211_X1 U5609 ( .C1(n6602), .C2(n4983), .A(n4982), .B(n4981), .ZN(n4984)
         );
  INV_X1 U5610 ( .A(n4984), .ZN(n4985) );
  NAND4_X1 U5611 ( .A1(n3781), .A2(n3771), .A3(n3779), .A4(n4985), .ZN(U2797)
         );
  OAI22_X1 U5612 ( .A1(n6593), .A2(n5088), .B1(n6582), .B2(n4986), .ZN(n6595)
         );
  OAI21_X1 U5613 ( .B1(n6595), .B2(n7605), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n4989) );
  NAND2_X1 U5614 ( .A1(n4987), .A2(n5044), .ZN(n4988) );
  NAND2_X1 U5615 ( .A1(n4989), .A2(n4988), .ZN(U2790) );
  INV_X1 U5616 ( .A(n4990), .ZN(n4992) );
  INV_X1 U5617 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n7629) );
  INV_X1 U5618 ( .A(n7305), .ZN(n4991) );
  OAI211_X1 U5619 ( .C1(n4992), .C2(n7629), .A(n7632), .B(n4991), .ZN(U2788)
         );
  INV_X1 U5620 ( .A(n4993), .ZN(n4994) );
  AOI21_X1 U5621 ( .B1(n4996), .B2(n4995), .A(n4994), .ZN(n7431) );
  INV_X1 U5622 ( .A(n7431), .ZN(n5113) );
  OAI21_X1 U5623 ( .B1(n7296), .B2(n4997), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5002) );
  OAI21_X1 U5624 ( .B1(n4998), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n7263), 
        .ZN(n5064) );
  INV_X1 U5625 ( .A(n5064), .ZN(n5000) );
  INV_X1 U5626 ( .A(REIP_REG_0__SCAN_IN), .ZN(n4999) );
  NOR2_X1 U5627 ( .A1(n7088), .A2(n4999), .ZN(n5056) );
  AOI21_X1 U5628 ( .B1(n7298), .B2(n5000), .A(n5056), .ZN(n5001) );
  OAI211_X1 U5629 ( .C1(n5113), .C2(n6976), .A(n5002), .B(n5001), .ZN(U2986)
         );
  NAND2_X1 U5630 ( .A1(n3704), .A2(n5003), .ZN(n5005) );
  XNOR2_X1 U5631 ( .A(n5005), .B(n5004), .ZN(n5824) );
  AOI21_X1 U5632 ( .B1(n5009), .B2(n5006), .A(n5008), .ZN(n7449) );
  AOI22_X1 U5633 ( .A1(n7296), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n7370), 
        .B2(REIP_REG_3__SCAN_IN), .ZN(n5010) );
  OAI21_X1 U5634 ( .B1(n7447), .B2(n7302), .A(n5010), .ZN(n5011) );
  AOI21_X1 U5635 ( .B1(n7449), .B2(n7297), .A(n5011), .ZN(n5012) );
  OAI21_X1 U5636 ( .B1(n5824), .B2(n7543), .A(n5012), .ZN(U2983) );
  NOR2_X1 U5637 ( .A1(n5044), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7593) );
  NAND2_X1 U5638 ( .A1(n6593), .A2(n6584), .ZN(n5015) );
  INV_X1 U5639 ( .A(n5091), .ZN(n5024) );
  INV_X1 U5640 ( .A(n5016), .ZN(n5019) );
  OAI22_X1 U5641 ( .A1(n5317), .A2(n3878), .B1(n7311), .B2(n6582), .ZN(n5017)
         );
  INV_X1 U5642 ( .A(n5017), .ZN(n5018) );
  NAND2_X1 U5643 ( .A1(n5019), .A2(n5018), .ZN(n5023) );
  OR2_X1 U5644 ( .A1(n4884), .A2(n3945), .ZN(n5020) );
  AND2_X1 U5645 ( .A1(n5021), .A2(n5020), .ZN(n5022) );
  NAND2_X1 U5646 ( .A1(n5026), .A2(n6589), .ZN(n5077) );
  NAND4_X1 U5647 ( .A1(n5024), .A2(n5023), .A3(n5022), .A4(n5077), .ZN(n5328)
         );
  INV_X1 U5648 ( .A(n5328), .ZN(n7560) );
  NAND2_X1 U5649 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .ZN(n7586) );
  NOR2_X1 U5650 ( .A1(n7318), .A2(n7586), .ZN(n7592) );
  INV_X1 U5651 ( .A(n7592), .ZN(n5025) );
  INV_X1 U5652 ( .A(FLUSH_REG_SCAN_IN), .ZN(n7571) );
  OAI22_X1 U5653 ( .A1(n7560), .A2(n7605), .B1(n5025), .B2(n7571), .ZN(n7549)
         );
  INV_X1 U5654 ( .A(n7598), .ZN(n6566) );
  INV_X1 U5655 ( .A(n5027), .ZN(n5038) );
  AOI22_X1 U5656 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n4945), .B2(n4078), .ZN(n6565)
         );
  NAND2_X1 U5657 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5045) );
  INV_X1 U5658 ( .A(n7548), .ZN(n5037) );
  INV_X1 U5659 ( .A(n4887), .ZN(n5029) );
  AND3_X1 U5660 ( .A1(n5030), .A2(n5029), .A3(n4769), .ZN(n5031) );
  AND3_X1 U5661 ( .A1(n5032), .A2(n5031), .A3(n4783), .ZN(n5315) );
  INV_X1 U5662 ( .A(n5315), .ZN(n5306) );
  INV_X1 U5663 ( .A(n5033), .ZN(n6567) );
  NAND3_X1 U5664 ( .A1(n5034), .A2(n6567), .A3(n5327), .ZN(n5035) );
  OAI21_X1 U5665 ( .B1(n7132), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n5035), 
        .ZN(n5036) );
  AOI21_X1 U5666 ( .B1(n5028), .B2(n5306), .A(n5036), .ZN(n7559) );
  OAI222_X1 U5667 ( .A1(n6566), .A2(n5038), .B1(n6565), .B2(n5045), .C1(n5037), 
        .C2(n7559), .ZN(n5040) );
  AOI22_X1 U5668 ( .A1(n7552), .A2(n5040), .B1(n5039), .B2(n7598), .ZN(n5041)
         );
  OAI21_X1 U5669 ( .B1(n5042), .B2(n7552), .A(n5041), .ZN(U3460) );
  INV_X1 U5670 ( .A(n4263), .ZN(n7425) );
  OAI22_X1 U5671 ( .A1(n7425), .A2(n5315), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5043), .ZN(n7557) );
  AOI21_X1 U5672 ( .B1(n7557), .B2(n5044), .A(STATE2_REG_1__SCAN_IN), .ZN(
        n5046) );
  INV_X1 U5673 ( .A(n5045), .ZN(n6564) );
  OAI22_X1 U5674 ( .A1(n5046), .A2(n6564), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6566), .ZN(n5047) );
  NOR2_X1 U5675 ( .A1(n7132), .A2(n5049), .ZN(n7556) );
  AOI22_X1 U5676 ( .A1(n7552), .A2(n5047), .B1(n7548), .B2(n7556), .ZN(n5048)
         );
  OAI21_X1 U5677 ( .B1(n5049), .B2(n7552), .A(n5048), .ZN(U3461) );
  INV_X1 U5678 ( .A(n5050), .ZN(n5053) );
  NAND2_X1 U5679 ( .A1(n5051), .A2(n5059), .ZN(n5052) );
  NAND2_X1 U5680 ( .A1(n5053), .A2(n5052), .ZN(n7426) );
  INV_X1 U5681 ( .A(n7426), .ZN(n5058) );
  INV_X1 U5682 ( .A(n5054), .ZN(n5055) );
  NOR2_X1 U5683 ( .A1(n7386), .A2(n5055), .ZN(n7337) );
  NOR2_X1 U5684 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n7337), .ZN(n5057)
         );
  AOI211_X1 U5685 ( .C1(n7418), .C2(n5058), .A(n5057), .B(n5056), .ZN(n5063)
         );
  AOI21_X1 U5686 ( .B1(n5060), .B2(n7336), .A(n5059), .ZN(n5061) );
  INV_X1 U5687 ( .A(n5061), .ZN(n5062) );
  OAI211_X1 U5688 ( .C1(n7350), .C2(n5064), .A(n5063), .B(n5062), .ZN(U3018)
         );
  XNOR2_X1 U5689 ( .A(n5066), .B(n5065), .ZN(n7107) );
  INV_X1 U5690 ( .A(n5067), .ZN(n5070) );
  INV_X1 U5691 ( .A(n5008), .ZN(n5069) );
  AOI21_X1 U5692 ( .B1(n5070), .B2(n5069), .A(n5068), .ZN(n7462) );
  NAND2_X1 U5693 ( .A1(n7370), .A2(REIP_REG_4__SCAN_IN), .ZN(n7099) );
  NAND2_X1 U5694 ( .A1(n7296), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5071)
         );
  OAI211_X1 U5695 ( .C1(n7302), .C2(n7465), .A(n7099), .B(n5071), .ZN(n5072)
         );
  AOI21_X1 U5696 ( .B1(n7462), .B2(n7297), .A(n5072), .ZN(n5073) );
  OAI21_X1 U5697 ( .B1(n7107), .B2(n7543), .A(n5073), .ZN(U2982) );
  AND4_X1 U5698 ( .A1(n6575), .A2(n5082), .A3(n3940), .A4(n3901), .ZN(n5074)
         );
  NAND2_X1 U5699 ( .A1(n5074), .A2(n4887), .ZN(n5089) );
  OR2_X1 U5700 ( .A1(n5089), .A2(n5075), .ZN(n5076) );
  NAND2_X1 U5701 ( .A1(n5077), .A2(n5076), .ZN(n5078) );
  NOR2_X1 U5702 ( .A1(n5080), .A2(n5079), .ZN(n5081) );
  NOR2_X1 U5703 ( .A1(n5099), .A2(n5081), .ZN(n7264) );
  INV_X1 U5704 ( .A(n7264), .ZN(n5104) );
  XNOR2_X1 U5705 ( .A(n5083), .B(n5085), .ZN(n7335) );
  INV_X1 U5706 ( .A(n7259), .ZN(n5152) );
  AOI22_X1 U5707 ( .A1(n6780), .A2(n7335), .B1(EBX_REG_1__SCAN_IN), .B2(n5152), 
        .ZN(n5084) );
  OAI21_X1 U5708 ( .B1(n7256), .B2(n5104), .A(n5084), .ZN(U2858) );
  NAND2_X1 U5709 ( .A1(n5085), .A2(n7634), .ZN(n5086) );
  NOR2_X1 U5710 ( .A1(n4769), .A2(n5086), .ZN(n5087) );
  INV_X1 U5711 ( .A(n5088), .ZN(n5708) );
  NOR2_X1 U5712 ( .A1(n5089), .A2(n5708), .ZN(n5090) );
  NAND2_X1 U5713 ( .A1(n5094), .A2(n4237), .ZN(n5095) );
  INV_X1 U5714 ( .A(n5095), .ZN(n5096) );
  INV_X1 U5715 ( .A(DATAI_0_), .ZN(n5141) );
  INV_X1 U5716 ( .A(EAX_REG_0__SCAN_IN), .ZN(n7638) );
  OAI222_X1 U5717 ( .A1(n5113), .A2(n6831), .B1(n6833), .B2(n5141), .C1(n6829), 
        .C2(n7638), .ZN(U2891) );
  INV_X1 U5718 ( .A(n7462), .ZN(n5112) );
  INV_X1 U5719 ( .A(EAX_REG_4__SCAN_IN), .ZN(n7652) );
  INV_X1 U5720 ( .A(DATAI_4_), .ZN(n5097) );
  OAI222_X1 U5721 ( .A1(n5112), .A2(n6831), .B1(n6829), .B2(n7652), .C1(n6833), 
        .C2(n5097), .ZN(U2887) );
  INV_X1 U5722 ( .A(DATAI_2_), .ZN(n6250) );
  INV_X1 U5723 ( .A(EAX_REG_2__SCAN_IN), .ZN(n7645) );
  INV_X1 U5724 ( .A(n5098), .ZN(n5102) );
  INV_X1 U5725 ( .A(n5099), .ZN(n5100) );
  NAND3_X1 U5726 ( .A1(n5102), .A2(n5101), .A3(n5100), .ZN(n5103) );
  AND2_X1 U5727 ( .A1(n5006), .A2(n5103), .ZN(n7271) );
  INV_X1 U5728 ( .A(n7271), .ZN(n5118) );
  OAI222_X1 U5729 ( .A1(n6833), .A2(n6250), .B1(n6829), .B2(n7645), .C1(n6831), 
        .C2(n5118), .ZN(U2889) );
  INV_X1 U5730 ( .A(DATAI_1_), .ZN(n5230) );
  INV_X1 U5731 ( .A(EAX_REG_1__SCAN_IN), .ZN(n7641) );
  OAI222_X1 U5732 ( .A1(n5230), .A2(n6833), .B1(n6829), .B2(n7641), .C1(n6831), 
        .C2(n5104), .ZN(U2890) );
  INV_X1 U5733 ( .A(DATAI_3_), .ZN(n5217) );
  INV_X1 U5734 ( .A(EAX_REG_3__SCAN_IN), .ZN(n7648) );
  INV_X1 U5735 ( .A(n7449), .ZN(n5105) );
  OAI222_X1 U5736 ( .A1(n5217), .A2(n6833), .B1(n6829), .B2(n7648), .C1(n6831), 
        .C2(n5105), .ZN(U2888) );
  INV_X1 U5737 ( .A(DATAI_5_), .ZN(n5109) );
  INV_X1 U5738 ( .A(EAX_REG_5__SCAN_IN), .ZN(n7656) );
  NOR2_X1 U5739 ( .A1(n5068), .A2(n5107), .ZN(n5108) );
  OR2_X1 U5740 ( .A1(n5106), .A2(n5108), .ZN(n5650) );
  OAI222_X1 U5741 ( .A1(n5109), .A2(n6833), .B1(n6829), .B2(n7656), .C1(n6831), 
        .C2(n5650), .ZN(U2886) );
  INV_X1 U5742 ( .A(EBX_REG_4__SCAN_IN), .ZN(n7458) );
  AND2_X1 U5743 ( .A1(n5722), .A2(n5110), .ZN(n5111) );
  OR2_X1 U5744 ( .A1(n5111), .A2(n5652), .ZN(n7459) );
  OAI222_X1 U5745 ( .A1(n5112), .A2(n7256), .B1(n7458), .B2(n7259), .C1(n7459), 
        .C2(n3659), .ZN(U2855) );
  OAI222_X1 U5746 ( .A1(n7426), .A2(n3659), .B1(n4793), .B2(n7259), .C1(n5113), 
        .C2(n7256), .ZN(U2859) );
  OR2_X1 U5747 ( .A1(n5116), .A2(n5115), .ZN(n5117) );
  AND2_X1 U5748 ( .A1(n5114), .A2(n5117), .ZN(n7347) );
  INV_X1 U5749 ( .A(n7347), .ZN(n5119) );
  INV_X1 U5750 ( .A(EBX_REG_2__SCAN_IN), .ZN(n5729) );
  OAI222_X1 U5751 ( .A1(n5119), .A2(n3659), .B1(n5729), .B2(n7259), .C1(n5118), 
        .C2(n7256), .ZN(U2857) );
  NAND3_X1 U5752 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n5481), .ZN(n5519) );
  NOR2_X1 U5753 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5519), .ZN(n5390)
         );
  INV_X1 U5754 ( .A(n5390), .ZN(n5123) );
  INV_X1 U5755 ( .A(n5281), .ZN(n5120) );
  NAND2_X1 U5756 ( .A1(n5162), .A2(n5120), .ZN(n5266) );
  AND2_X1 U5757 ( .A1(n5266), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5261) );
  INV_X1 U5758 ( .A(n5134), .ZN(n5122) );
  NAND2_X1 U5759 ( .A1(n5122), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5560) );
  NAND2_X1 U5760 ( .A1(n5260), .A2(n5560), .ZN(n5285) );
  AOI211_X1 U5761 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5123), .A(n5261), .B(
        n5285), .ZN(n5131) );
  OR2_X1 U5762 ( .A1(n3661), .A2(n5870), .ZN(n5747) );
  NOR2_X1 U5763 ( .A1(n5125), .A2(n5028), .ZN(n5516) );
  NOR2_X1 U5764 ( .A1(n5516), .A2(n5870), .ZN(n5161) );
  NAND2_X1 U5765 ( .A1(n5126), .A2(n5158), .ZN(n5193) );
  INV_X1 U5766 ( .A(n5918), .ZN(n5184) );
  NOR2_X1 U5767 ( .A1(n5127), .A2(n5258), .ZN(n5436) );
  AND2_X1 U5768 ( .A1(n5436), .A2(n5487), .ZN(n5157) );
  OAI21_X1 U5769 ( .B1(n5184), .B2(n5465), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5129) );
  OAI21_X1 U5770 ( .B1(n5668), .B2(n5161), .A(n5129), .ZN(n5130) );
  INV_X1 U5771 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5139) );
  NAND2_X1 U5772 ( .A1(n5182), .A2(n4237), .ZN(n6413) );
  NAND2_X1 U5773 ( .A1(n7297), .A2(DATAI_23_), .ZN(n6419) );
  INV_X1 U5774 ( .A(n6419), .ZN(n5698) );
  AOI22_X1 U5775 ( .A1(n6014), .A2(n5390), .B1(n5698), .B2(n5184), .ZN(n5138)
         );
  INV_X1 U5776 ( .A(DATAI_7_), .ZN(n5602) );
  INV_X1 U5777 ( .A(n5516), .ZN(n5133) );
  INV_X1 U5778 ( .A(n5870), .ZN(n5875) );
  NAND2_X1 U5779 ( .A1(n3661), .A2(n5875), .ZN(n5265) );
  OR2_X1 U5780 ( .A1(n5133), .A2(n5265), .ZN(n5136) );
  NAND2_X1 U5781 ( .A1(n5134), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5282) );
  OR2_X1 U5782 ( .A1(n5266), .A2(n5282), .ZN(n5135) );
  NAND2_X1 U5783 ( .A1(n5136), .A2(n5135), .ZN(n5185) );
  NAND2_X1 U5784 ( .A1(n7297), .A2(DATAI_31_), .ZN(n6410) );
  INV_X1 U5785 ( .A(n6410), .ZN(n6018) );
  AOI22_X1 U5786 ( .A1(n6416), .A2(n5185), .B1(n6018), .B2(n5465), .ZN(n5137)
         );
  OAI211_X1 U5787 ( .C1(n5394), .C2(n5139), .A(n5138), .B(n5137), .ZN(U3123)
         );
  INV_X1 U5788 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5145) );
  NAND2_X1 U5789 ( .A1(n7297), .A2(DATAI_16_), .ZN(n5970) );
  INV_X1 U5790 ( .A(n5185), .ZN(n5388) );
  OAI22_X1 U5791 ( .A1(n5918), .A2(n5970), .B1(n5388), .B2(n5748), .ZN(n5142)
         );
  AOI21_X1 U5792 ( .B1(n5750), .B2(n5390), .A(n5142), .ZN(n5144) );
  NAND2_X1 U5793 ( .A1(n7297), .A2(DATAI_24_), .ZN(n5942) );
  INV_X1 U5794 ( .A(n5942), .ZN(n5968) );
  NAND2_X1 U5795 ( .A1(n5465), .A2(n5968), .ZN(n5143) );
  OAI211_X1 U5796 ( .C1(n5394), .C2(n5145), .A(n5144), .B(n5143), .ZN(U3116)
         );
  NAND2_X1 U5797 ( .A1(n5147), .A2(n5148), .ZN(n5149) );
  NAND2_X1 U5798 ( .A1(n5146), .A2(n5149), .ZN(n6430) );
  AND2_X1 U5799 ( .A1(n5704), .A2(n5150), .ZN(n5151) );
  NOR2_X1 U5800 ( .A1(n5813), .A2(n5151), .ZN(n7361) );
  AOI22_X1 U5801 ( .A1(n6780), .A2(n7361), .B1(EBX_REG_8__SCAN_IN), .B2(n5152), 
        .ZN(n5153) );
  OAI21_X1 U5802 ( .B1(n6430), .B2(n7256), .A(n5153), .ZN(U2851) );
  OAI21_X1 U5803 ( .B1(n5654), .B2(n5154), .A(n5702), .ZN(n7480) );
  INV_X1 U5804 ( .A(n5598), .ZN(n5155) );
  XNOR2_X1 U5805 ( .A(n5106), .B(n5155), .ZN(n7484) );
  INV_X1 U5806 ( .A(n7484), .ZN(n5239) );
  INV_X1 U5807 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5156) );
  OAI222_X1 U5808 ( .A1(n7480), .A2(n3659), .B1(n7256), .B2(n5239), .C1(n5156), 
        .C2(n7259), .ZN(U2853) );
  INV_X1 U5809 ( .A(n5158), .ZN(n5159) );
  NAND2_X1 U5810 ( .A1(n5126), .A2(n5159), .ZN(n5259) );
  INV_X1 U5811 ( .A(n5259), .ZN(n5160) );
  NAND2_X1 U5812 ( .A1(n5160), .A2(n5258), .ZN(n5499) );
  AOI21_X1 U5813 ( .B1(n5926), .B2(n5643), .A(n7608), .ZN(n5166) );
  INV_X1 U5814 ( .A(n5265), .ZN(n5734) );
  NOR2_X1 U5815 ( .A1(n5161), .A2(n5734), .ZN(n5165) );
  NAND3_X1 U5816 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n7566), .A3(n5481), .ZN(n5506) );
  NOR2_X1 U5817 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5506), .ZN(n5353)
         );
  INV_X1 U5818 ( .A(n5353), .ZN(n5163) );
  NOR2_X1 U5819 ( .A1(n5162), .A2(n5281), .ZN(n5744) );
  NOR2_X1 U5820 ( .A1(n5744), .A2(n7584), .ZN(n5739) );
  AOI211_X1 U5821 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5163), .A(n5739), .B(
        n5285), .ZN(n5164) );
  NAND2_X1 U5822 ( .A1(n5350), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5171) );
  NAND2_X1 U5823 ( .A1(n5668), .A2(n5516), .ZN(n5168) );
  INV_X1 U5824 ( .A(n5282), .ZN(n5190) );
  NAND2_X1 U5825 ( .A1(n5744), .A2(n5190), .ZN(n5167) );
  OAI22_X1 U5826 ( .A1(n5926), .A2(n5970), .B1(n5351), .B2(n5748), .ZN(n5169)
         );
  AOI21_X1 U5827 ( .B1(n5750), .B2(n5353), .A(n5169), .ZN(n5170) );
  OAI211_X1 U5828 ( .C1(n5643), .C2(n5942), .A(n5171), .B(n5170), .ZN(U3052)
         );
  INV_X1 U5829 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5176) );
  NAND2_X1 U5830 ( .A1(n5182), .A2(n5172), .ZN(n5789) );
  INV_X1 U5831 ( .A(DATAI_21_), .ZN(n5173) );
  NOR2_X1 U5832 ( .A1(n6976), .A2(n5173), .ZN(n5673) );
  AOI22_X1 U5833 ( .A1(n5991), .A2(n5390), .B1(n5673), .B2(n5184), .ZN(n5175)
         );
  INV_X1 U5834 ( .A(n5997), .ZN(n5792) );
  NAND2_X1 U5835 ( .A1(n7297), .A2(DATAI_29_), .ZN(n5787) );
  INV_X1 U5836 ( .A(n5787), .ZN(n5995) );
  AOI22_X1 U5837 ( .A1(n5792), .A2(n5185), .B1(n5995), .B2(n5465), .ZN(n5174)
         );
  OAI211_X1 U5838 ( .C1(n5394), .C2(n5176), .A(n5175), .B(n5174), .ZN(U3121)
         );
  INV_X1 U5839 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5181) );
  NAND2_X1 U5840 ( .A1(n5182), .A2(n5177), .ZN(n5759) );
  INV_X1 U5841 ( .A(DATAI_20_), .ZN(n5178) );
  NOR2_X1 U5842 ( .A1(n6976), .A2(n5178), .ZN(n5681) );
  AOI22_X1 U5843 ( .A1(n6005), .A2(n5390), .B1(n5681), .B2(n5184), .ZN(n5180)
         );
  INV_X1 U5844 ( .A(n6011), .ZN(n5761) );
  NAND2_X1 U5845 ( .A1(n7297), .A2(DATAI_28_), .ZN(n5758) );
  INV_X1 U5846 ( .A(n5758), .ZN(n6009) );
  AOI22_X1 U5847 ( .A1(n5761), .A2(n5185), .B1(n6009), .B2(n5465), .ZN(n5179)
         );
  OAI211_X1 U5848 ( .C1(n5394), .C2(n5181), .A(n5180), .B(n5179), .ZN(U3120)
         );
  INV_X1 U5849 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5188) );
  NAND2_X1 U5850 ( .A1(n5182), .A2(n3901), .ZN(n5780) );
  INV_X1 U5851 ( .A(DATAI_22_), .ZN(n5183) );
  NOR2_X1 U5852 ( .A1(n6976), .A2(n5183), .ZN(n5677) );
  AOI22_X1 U5853 ( .A1(n5998), .A2(n5390), .B1(n5677), .B2(n5184), .ZN(n5187)
         );
  INV_X1 U5854 ( .A(n6004), .ZN(n5782) );
  NAND2_X1 U5855 ( .A1(n7297), .A2(DATAI_30_), .ZN(n5779) );
  INV_X1 U5856 ( .A(n5779), .ZN(n6002) );
  AOI22_X1 U5857 ( .A1(n5782), .A2(n5185), .B1(n6002), .B2(n5465), .ZN(n5186)
         );
  OAI211_X1 U5858 ( .C1(n5394), .C2(n5188), .A(n5187), .B(n5186), .ZN(U3122)
         );
  INV_X1 U5859 ( .A(n5028), .ZN(n5711) );
  NOR2_X1 U5860 ( .A1(n5125), .A2(n5711), .ZN(n5470) );
  INV_X1 U5861 ( .A(n5470), .ZN(n5189) );
  OR2_X1 U5862 ( .A1(n5189), .A2(n5265), .ZN(n5192) );
  AND2_X1 U5863 ( .A1(n5281), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5561)
         );
  NAND2_X1 U5864 ( .A1(n5190), .A2(n5561), .ZN(n5191) );
  AOI21_X1 U5865 ( .B1(n5894), .B2(n5603), .A(n7608), .ZN(n5196) );
  NOR2_X1 U5866 ( .A1(n5470), .A2(n5870), .ZN(n5284) );
  NOR2_X1 U5867 ( .A1(n5284), .A2(n5668), .ZN(n5195) );
  NAND3_X1 U5868 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5400) );
  NOR2_X1 U5869 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5400), .ZN(n5235)
         );
  INV_X1 U5870 ( .A(n5235), .ZN(n5204) );
  AOI21_X1 U5871 ( .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n5281), .A(n7584), 
        .ZN(n5564) );
  AOI211_X1 U5872 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5204), .A(n5564), .B(
        n5285), .ZN(n5194) );
  NAND2_X1 U5873 ( .A1(n5214), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5199)
         );
  OAI22_X1 U5874 ( .A1(n6419), .A2(n5603), .B1(n5894), .B2(n6410), .ZN(n5197)
         );
  AOI21_X1 U5875 ( .B1(n6014), .B2(n5235), .A(n5197), .ZN(n5198) );
  OAI211_X1 U5876 ( .C1(n5216), .C2(n6021), .A(n5199), .B(n5198), .ZN(U3139)
         );
  NAND2_X1 U5877 ( .A1(n5214), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5203)
         );
  INV_X1 U5878 ( .A(n5970), .ZN(n5944) );
  INV_X1 U5879 ( .A(n5603), .ZN(n5201) );
  OAI22_X1 U5880 ( .A1(n5894), .A2(n5942), .B1(n5216), .B2(n5748), .ZN(n5200)
         );
  AOI21_X1 U5881 ( .B1(n5944), .B2(n5201), .A(n5200), .ZN(n5202) );
  OAI211_X1 U5882 ( .C1(n5966), .C2(n5204), .A(n5203), .B(n5202), .ZN(U3132)
         );
  NAND2_X1 U5883 ( .A1(n5214), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5207)
         );
  INV_X1 U5884 ( .A(n5681), .ZN(n6007) );
  OAI22_X1 U5885 ( .A1(n6007), .A2(n5603), .B1(n5894), .B2(n5758), .ZN(n5205)
         );
  AOI21_X1 U5886 ( .B1(n6005), .B2(n5235), .A(n5205), .ZN(n5206) );
  OAI211_X1 U5887 ( .C1(n5216), .C2(n6011), .A(n5207), .B(n5206), .ZN(U3136)
         );
  NAND2_X1 U5888 ( .A1(n5214), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5210)
         );
  INV_X1 U5889 ( .A(n5677), .ZN(n6000) );
  OAI22_X1 U5890 ( .A1(n6000), .A2(n5603), .B1(n5894), .B2(n5779), .ZN(n5208)
         );
  AOI21_X1 U5891 ( .B1(n5998), .B2(n5235), .A(n5208), .ZN(n5209) );
  OAI211_X1 U5892 ( .C1(n5216), .C2(n6004), .A(n5210), .B(n5209), .ZN(U3138)
         );
  NAND2_X1 U5893 ( .A1(n5214), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5213)
         );
  INV_X1 U5894 ( .A(n5673), .ZN(n5993) );
  OAI22_X1 U5895 ( .A1(n5993), .A2(n5603), .B1(n5894), .B2(n5787), .ZN(n5211)
         );
  AOI21_X1 U5896 ( .B1(n5991), .B2(n5235), .A(n5211), .ZN(n5212) );
  OAI211_X1 U5897 ( .C1(n5216), .C2(n5997), .A(n5213), .B(n5212), .ZN(U3137)
         );
  INV_X1 U5898 ( .A(n5214), .ZN(n5238) );
  INV_X1 U5899 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5222) );
  NAND2_X1 U5900 ( .A1(n7297), .A2(DATAI_27_), .ZN(n5932) );
  NAND2_X1 U5901 ( .A1(n7297), .A2(DATAI_19_), .ZN(n5963) );
  OR2_X1 U5902 ( .A1(n5603), .A2(n5963), .ZN(n5219) );
  INV_X1 U5903 ( .A(n5216), .ZN(n5231) );
  NAND2_X1 U5904 ( .A1(n5231), .A2(n5957), .ZN(n5218) );
  OAI211_X1 U5905 ( .C1(n5894), .C2(n5932), .A(n5219), .B(n5218), .ZN(n5220)
         );
  AOI21_X1 U5906 ( .B1(n5766), .B2(n5235), .A(n5220), .ZN(n5221) );
  OAI21_X1 U5907 ( .B1(n5238), .B2(n5222), .A(n5221), .ZN(U3135) );
  INV_X1 U5908 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5227) );
  NOR2_X1 U5909 ( .A1(n5229), .A2(n3906), .ZN(n5755) );
  NAND2_X1 U5910 ( .A1(n7297), .A2(DATAI_26_), .ZN(n5937) );
  NAND2_X1 U5911 ( .A1(n7297), .A2(DATAI_18_), .ZN(n5988) );
  OR2_X1 U5912 ( .A1(n5603), .A2(n5988), .ZN(n5224) );
  NAND2_X1 U5913 ( .A1(n5231), .A2(n5979), .ZN(n5223) );
  OAI211_X1 U5914 ( .C1(n5894), .C2(n5937), .A(n5224), .B(n5223), .ZN(n5225)
         );
  AOI21_X1 U5915 ( .B1(n5755), .B2(n5235), .A(n5225), .ZN(n5226) );
  OAI21_X1 U5916 ( .B1(n5238), .B2(n5227), .A(n5226), .ZN(U3134) );
  INV_X1 U5917 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U5918 ( .A1(n7297), .A2(DATAI_25_), .ZN(n5949) );
  NAND2_X1 U5919 ( .A1(n7297), .A2(DATAI_17_), .ZN(n5977) );
  OR2_X1 U5920 ( .A1(n5603), .A2(n5977), .ZN(n5233) );
  NAND2_X1 U5921 ( .A1(n5231), .A2(n5971), .ZN(n5232) );
  OAI211_X1 U5922 ( .C1(n5894), .C2(n5949), .A(n5233), .B(n5232), .ZN(n5234)
         );
  AOI21_X1 U5923 ( .B1(n5776), .B2(n5235), .A(n5234), .ZN(n5236) );
  OAI21_X1 U5924 ( .B1(n5238), .B2(n5237), .A(n5236), .ZN(U3133) );
  INV_X1 U5925 ( .A(DATAI_6_), .ZN(n5240) );
  INV_X1 U5926 ( .A(EAX_REG_6__SCAN_IN), .ZN(n7660) );
  OAI222_X1 U5927 ( .A1(n6833), .A2(n5240), .B1(n6829), .B2(n7660), .C1(n6831), 
        .C2(n5239), .ZN(U2885) );
  INV_X1 U5928 ( .A(DATAI_8_), .ZN(n5241) );
  INV_X1 U5929 ( .A(EAX_REG_8__SCAN_IN), .ZN(n7668) );
  OAI222_X1 U5930 ( .A1(n6833), .A2(n5241), .B1(n6829), .B2(n7668), .C1(n6831), 
        .C2(n6430), .ZN(U2883) );
  INV_X1 U5931 ( .A(n5350), .ZN(n5257) );
  INV_X1 U5932 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5244) );
  INV_X1 U5933 ( .A(n5926), .ZN(n5251) );
  AOI22_X1 U5934 ( .A1(n5998), .A2(n5353), .B1(n5677), .B2(n5251), .ZN(n5243)
         );
  INV_X1 U5935 ( .A(n5351), .ZN(n5253) );
  INV_X1 U5936 ( .A(n5643), .ZN(n5252) );
  AOI22_X1 U5937 ( .A1(n5782), .A2(n5253), .B1(n6002), .B2(n5252), .ZN(n5242)
         );
  OAI211_X1 U5938 ( .C1(n5257), .C2(n5244), .A(n5243), .B(n5242), .ZN(U3058)
         );
  INV_X1 U5939 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5247) );
  AOI22_X1 U5940 ( .A1(n6014), .A2(n5353), .B1(n5698), .B2(n5251), .ZN(n5246)
         );
  AOI22_X1 U5941 ( .A1(n6416), .A2(n5253), .B1(n6018), .B2(n5252), .ZN(n5245)
         );
  OAI211_X1 U5942 ( .C1(n5257), .C2(n5247), .A(n5246), .B(n5245), .ZN(U3059)
         );
  INV_X1 U5943 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5250) );
  AOI22_X1 U5944 ( .A1(n6005), .A2(n5353), .B1(n5681), .B2(n5251), .ZN(n5249)
         );
  AOI22_X1 U5945 ( .A1(n5761), .A2(n5253), .B1(n6009), .B2(n5252), .ZN(n5248)
         );
  OAI211_X1 U5946 ( .C1(n5257), .C2(n5250), .A(n5249), .B(n5248), .ZN(U3056)
         );
  INV_X1 U5947 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5256) );
  AOI22_X1 U5948 ( .A1(n5991), .A2(n5353), .B1(n5673), .B2(n5251), .ZN(n5255)
         );
  AOI22_X1 U5949 ( .A1(n5792), .A2(n5253), .B1(n5995), .B2(n5252), .ZN(n5254)
         );
  OAI211_X1 U5950 ( .C1(n5257), .C2(n5256), .A(n5255), .B(n5254), .ZN(U3057)
         );
  NAND2_X1 U5951 ( .A1(n5480), .A2(n5128), .ZN(n5868) );
  AOI21_X1 U5952 ( .B1(n6420), .B2(n6411), .A(n7608), .ZN(n5264) );
  AND2_X1 U5953 ( .A1(n5125), .A2(n5711), .ZN(n5866) );
  NOR2_X1 U5954 ( .A1(n5866), .A2(n5870), .ZN(n5735) );
  NOR2_X1 U5955 ( .A1(n5735), .A2(n5668), .ZN(n5263) );
  NOR3_X1 U5956 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n7566), .ZN(n5874) );
  NAND2_X1 U5957 ( .A1(n5874), .A2(n3937), .ZN(n6412) );
  NAND2_X1 U5958 ( .A1(n5260), .A2(n5282), .ZN(n5738) );
  AOI211_X1 U5959 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6412), .A(n5261), .B(
        n5738), .ZN(n5262) );
  NAND2_X1 U5960 ( .A1(n6409), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5271) );
  INV_X1 U5961 ( .A(n5866), .ZN(n5746) );
  OR2_X1 U5962 ( .A1(n5265), .A2(n5746), .ZN(n5268) );
  OR2_X1 U5963 ( .A1(n5266), .A2(n5560), .ZN(n5267) );
  NAND2_X1 U5964 ( .A1(n5268), .A2(n5267), .ZN(n6415) );
  OAI22_X1 U5965 ( .A1(n5759), .A2(n6412), .B1(n6411), .B2(n5758), .ZN(n5269)
         );
  AOI21_X1 U5966 ( .B1(n5761), .B2(n6415), .A(n5269), .ZN(n5270) );
  OAI211_X1 U5967 ( .C1(n6007), .C2(n6420), .A(n5271), .B(n5270), .ZN(U3088)
         );
  NAND2_X1 U5968 ( .A1(n6409), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5274) );
  OAI22_X1 U5969 ( .A1(n5780), .A2(n6412), .B1(n6411), .B2(n5779), .ZN(n5272)
         );
  AOI21_X1 U5970 ( .B1(n5782), .B2(n6415), .A(n5272), .ZN(n5273) );
  OAI211_X1 U5971 ( .C1(n6000), .C2(n6420), .A(n5274), .B(n5273), .ZN(U3090)
         );
  NAND2_X1 U5972 ( .A1(n6409), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5277) );
  OAI22_X1 U5973 ( .A1(n5789), .A2(n6412), .B1(n6411), .B2(n5787), .ZN(n5275)
         );
  AOI21_X1 U5974 ( .B1(n5792), .B2(n6415), .A(n5275), .ZN(n5276) );
  OAI211_X1 U5975 ( .C1(n5993), .C2(n6420), .A(n5277), .B(n5276), .ZN(U3089)
         );
  NAND2_X1 U5976 ( .A1(n6409), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5280) );
  INV_X1 U5977 ( .A(n6412), .ZN(n5367) );
  INV_X1 U5978 ( .A(n6415), .ZN(n5365) );
  OAI22_X1 U5979 ( .A1(n6411), .A2(n5942), .B1(n5365), .B2(n5748), .ZN(n5278)
         );
  AOI21_X1 U5980 ( .B1(n5750), .B2(n5367), .A(n5278), .ZN(n5279) );
  OAI211_X1 U5981 ( .C1(n5970), .C2(n6420), .A(n5280), .B(n5279), .ZN(U3084)
         );
  NAND2_X1 U5982 ( .A1(n5281), .A2(n7566), .ZN(n5665) );
  NOR2_X1 U5983 ( .A1(n5282), .A2(n5665), .ZN(n5283) );
  AOI21_X1 U5984 ( .B1(n5668), .B2(n5470), .A(n5283), .ZN(n5374) );
  AOI21_X1 U5985 ( .B1(n5950), .B2(n5899), .A(n7608), .ZN(n5289) );
  NOR2_X1 U5986 ( .A1(n5284), .A2(n5734), .ZN(n5288) );
  NAND3_X1 U5987 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n7566), .ZN(n5473) );
  NOR2_X1 U5988 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5473), .ZN(n5303)
         );
  INV_X1 U5989 ( .A(n5303), .ZN(n5379) );
  NAND2_X1 U5990 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5665), .ZN(n5662) );
  INV_X1 U5991 ( .A(n5662), .ZN(n5286) );
  AOI211_X1 U5992 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5379), .A(n5286), .B(
        n5285), .ZN(n5287) );
  NAND2_X1 U5993 ( .A1(n5373), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5292) );
  OAI22_X1 U5994 ( .A1(n6007), .A2(n5950), .B1(n5899), .B2(n5758), .ZN(n5290)
         );
  AOI21_X1 U5995 ( .B1(n6005), .B2(n5303), .A(n5290), .ZN(n5291) );
  OAI211_X1 U5996 ( .C1(n5374), .C2(n6011), .A(n5292), .B(n5291), .ZN(U3072)
         );
  NAND2_X1 U5997 ( .A1(n5373), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5295) );
  OAI22_X1 U5998 ( .A1(n5993), .A2(n5950), .B1(n5899), .B2(n5787), .ZN(n5293)
         );
  AOI21_X1 U5999 ( .B1(n5991), .B2(n5303), .A(n5293), .ZN(n5294) );
  OAI211_X1 U6000 ( .C1(n5374), .C2(n5997), .A(n5295), .B(n5294), .ZN(U3073)
         );
  NAND2_X1 U6001 ( .A1(n5373), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n5298) );
  OAI22_X1 U6002 ( .A1(n5899), .A2(n5942), .B1(n5374), .B2(n5748), .ZN(n5296)
         );
  AOI21_X1 U6003 ( .B1(n5376), .B2(n5944), .A(n5296), .ZN(n5297) );
  OAI211_X1 U6004 ( .C1(n5966), .C2(n5379), .A(n5298), .B(n5297), .ZN(U3068)
         );
  NAND2_X1 U6005 ( .A1(n5373), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5301) );
  OAI22_X1 U6006 ( .A1(n6419), .A2(n5950), .B1(n5899), .B2(n6410), .ZN(n5299)
         );
  AOI21_X1 U6007 ( .B1(n6014), .B2(n5303), .A(n5299), .ZN(n5300) );
  OAI211_X1 U6008 ( .C1(n5374), .C2(n6021), .A(n5301), .B(n5300), .ZN(U3075)
         );
  NAND2_X1 U6009 ( .A1(n5373), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5305) );
  OAI22_X1 U6010 ( .A1(n6000), .A2(n5950), .B1(n5899), .B2(n5779), .ZN(n5302)
         );
  AOI21_X1 U6011 ( .B1(n5998), .B2(n5303), .A(n5302), .ZN(n5304) );
  OAI211_X1 U6012 ( .C1(n5374), .C2(n6004), .A(n5305), .B(n5304), .ZN(U3074)
         );
  NAND2_X1 U6013 ( .A1(n3661), .A2(n5306), .ZN(n5314) );
  OR2_X1 U6014 ( .A1(n6589), .A2(n6584), .ZN(n5319) );
  MUX2_X1 U6015 ( .A(n5307), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n5033), 
        .Z(n5309) );
  NOR2_X1 U6016 ( .A1(n5309), .A2(n5308), .ZN(n5312) );
  XNOR2_X1 U6017 ( .A(n5310), .B(n6518), .ZN(n5311) );
  AOI22_X1 U6018 ( .A1(n5319), .A2(n5312), .B1(n5317), .B2(n5311), .ZN(n5313)
         );
  NAND2_X1 U6019 ( .A1(n5314), .A2(n5313), .ZN(n6515) );
  MUX2_X1 U6020 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6515), .S(n5328), 
        .Z(n7565) );
  OR2_X1 U6021 ( .A1(n5328), .A2(n6573), .ZN(n5323) );
  OR2_X1 U6022 ( .A1(n5125), .A2(n5315), .ZN(n5321) );
  XNOR2_X1 U6023 ( .A(n5033), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5318)
         );
  XNOR2_X1 U6024 ( .A(n6573), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5316)
         );
  AOI22_X1 U6025 ( .A1(n5319), .A2(n5318), .B1(n5317), .B2(n5316), .ZN(n5320)
         );
  NAND2_X1 U6026 ( .A1(n5321), .A2(n5320), .ZN(n6570) );
  NAND2_X1 U6027 ( .A1(n5328), .A2(n6570), .ZN(n5322) );
  NAND2_X1 U6028 ( .A1(n5323), .A2(n5322), .ZN(n7555) );
  NAND3_X1 U6029 ( .A1(n7565), .A2(n5338), .A3(n7555), .ZN(n5326) );
  NOR2_X1 U6030 ( .A1(FLUSH_REG_SCAN_IN), .A2(n5338), .ZN(n5324) );
  NAND2_X1 U6031 ( .A1(n5308), .A2(n5324), .ZN(n5325) );
  NAND2_X1 U6032 ( .A1(n5326), .A2(n5325), .ZN(n7576) );
  NAND2_X1 U6033 ( .A1(n7576), .A2(n5327), .ZN(n5336) );
  MUX2_X1 U6034 ( .A(n5328), .B(FLUSH_REG_SCAN_IN), .S(STATE2_REG_1__SCAN_IN), 
        .Z(n5334) );
  INV_X1 U6035 ( .A(n5330), .ZN(n5331) );
  NOR2_X1 U6036 ( .A1(n5329), .A2(n5331), .ZN(n5332) );
  XNOR2_X1 U6037 ( .A(n5332), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n7545)
         );
  OR3_X1 U6038 ( .A1(n7545), .A2(STATE2_REG_1__SCAN_IN), .A3(n4783), .ZN(n5333) );
  OAI21_X1 U6039 ( .B1(n5334), .B2(n7551), .A(n5333), .ZN(n7578) );
  INV_X1 U6040 ( .A(n7578), .ZN(n5335) );
  NAND2_X1 U6041 ( .A1(n5336), .A2(n5335), .ZN(n5803) );
  OAI21_X1 U6042 ( .B1(n5803), .B2(FLUSH_REG_SCAN_IN), .A(n7592), .ZN(n5337)
         );
  NAND2_X1 U6043 ( .A1(n5337), .A2(n5399), .ZN(n7129) );
  OAI21_X1 U6044 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5338), .A(n7129), .ZN(
        n5809) );
  INV_X1 U6045 ( .A(n3661), .ZN(n7438) );
  NAND2_X1 U6046 ( .A1(n7129), .A2(n5875), .ZN(n5805) );
  AND2_X1 U6047 ( .A1(n5339), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5471) );
  AND2_X1 U6048 ( .A1(n5340), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5517) );
  AOI21_X1 U6049 ( .B1(n5126), .B2(STATEBS16_REG_SCAN_IN), .A(n5617), .ZN(
        n5341) );
  NOR3_X1 U6050 ( .A1(n5471), .A2(n5517), .A3(n5341), .ZN(n5342) );
  OAI222_X1 U6051 ( .A1(n7129), .A2(n7566), .B1(n5809), .B2(n7438), .C1(n5805), 
        .C2(n5342), .ZN(U3462) );
  XNOR2_X1 U6052 ( .A(n4255), .B(STATEBS16_REG_SCAN_IN), .ZN(n5343) );
  OAI222_X1 U6053 ( .A1(n5809), .A2(n5711), .B1(n7129), .B2(n5481), .C1(n5805), 
        .C2(n5343), .ZN(U3464) );
  NAND2_X1 U6054 ( .A1(n5350), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5346) );
  OAI22_X1 U6055 ( .A1(n5926), .A2(n5963), .B1(n5351), .B2(n5764), .ZN(n5344)
         );
  AOI21_X1 U6056 ( .B1(n5766), .B2(n5353), .A(n5344), .ZN(n5345) );
  OAI211_X1 U6057 ( .C1(n5643), .C2(n5932), .A(n5346), .B(n5345), .ZN(U3055)
         );
  NAND2_X1 U6058 ( .A1(n5350), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5349) );
  OAI22_X1 U6059 ( .A1(n5926), .A2(n5988), .B1(n5351), .B2(n5753), .ZN(n5347)
         );
  AOI21_X1 U6060 ( .B1(n5755), .B2(n5353), .A(n5347), .ZN(n5348) );
  OAI211_X1 U6061 ( .C1(n5643), .C2(n5937), .A(n5349), .B(n5348), .ZN(U3054)
         );
  NAND2_X1 U6062 ( .A1(n5350), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5355) );
  OAI22_X1 U6063 ( .A1(n5926), .A2(n5977), .B1(n5351), .B2(n5772), .ZN(n5352)
         );
  AOI21_X1 U6064 ( .B1(n5776), .B2(n5353), .A(n5352), .ZN(n5354) );
  OAI211_X1 U6065 ( .C1(n5643), .C2(n5949), .A(n5355), .B(n5354), .ZN(U3053)
         );
  NAND2_X1 U6066 ( .A1(n6409), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5358) );
  OAI22_X1 U6067 ( .A1(n6411), .A2(n5949), .B1(n5365), .B2(n5772), .ZN(n5356)
         );
  AOI21_X1 U6068 ( .B1(n5776), .B2(n5367), .A(n5356), .ZN(n5357) );
  OAI211_X1 U6069 ( .C1(n5977), .C2(n6420), .A(n5358), .B(n5357), .ZN(U3085)
         );
  NAND2_X1 U6070 ( .A1(n6409), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5361) );
  OAI22_X1 U6071 ( .A1(n6411), .A2(n5937), .B1(n5365), .B2(n5753), .ZN(n5359)
         );
  AOI21_X1 U6072 ( .B1(n5755), .B2(n5367), .A(n5359), .ZN(n5360) );
  OAI211_X1 U6073 ( .C1(n5988), .C2(n6420), .A(n5361), .B(n5360), .ZN(U3086)
         );
  NAND2_X1 U6074 ( .A1(n5373), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5364) );
  INV_X1 U6075 ( .A(n5977), .ZN(n5952) );
  OAI22_X1 U6076 ( .A1(n5899), .A2(n5949), .B1(n5374), .B2(n5772), .ZN(n5362)
         );
  AOI21_X1 U6077 ( .B1(n5376), .B2(n5952), .A(n5362), .ZN(n5363) );
  OAI211_X1 U6078 ( .C1(n5379), .C2(n5973), .A(n5364), .B(n5363), .ZN(U3069)
         );
  NAND2_X1 U6079 ( .A1(n6409), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5369) );
  OAI22_X1 U6080 ( .A1(n6411), .A2(n5932), .B1(n5365), .B2(n5764), .ZN(n5366)
         );
  AOI21_X1 U6081 ( .B1(n5766), .B2(n5367), .A(n5366), .ZN(n5368) );
  OAI211_X1 U6082 ( .C1(n5963), .C2(n6420), .A(n5369), .B(n5368), .ZN(U3087)
         );
  NAND2_X1 U6083 ( .A1(n5373), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5372) );
  INV_X1 U6084 ( .A(n5988), .ZN(n5939) );
  OAI22_X1 U6085 ( .A1(n5899), .A2(n5937), .B1(n5374), .B2(n5753), .ZN(n5370)
         );
  AOI21_X1 U6086 ( .B1(n5376), .B2(n5939), .A(n5370), .ZN(n5371) );
  OAI211_X1 U6087 ( .C1(n5379), .C2(n5983), .A(n5372), .B(n5371), .ZN(U3070)
         );
  NAND2_X1 U6088 ( .A1(n5373), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5378) );
  INV_X1 U6089 ( .A(n5963), .ZN(n5934) );
  OAI22_X1 U6090 ( .A1(n5899), .A2(n5932), .B1(n5374), .B2(n5764), .ZN(n5375)
         );
  AOI21_X1 U6091 ( .B1(n5376), .B2(n5934), .A(n5375), .ZN(n5377) );
  OAI211_X1 U6092 ( .C1(n5379), .C2(n5959), .A(n5378), .B(n5377), .ZN(U3071)
         );
  INV_X1 U6093 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5383) );
  OAI22_X1 U6094 ( .A1(n5918), .A2(n5963), .B1(n5388), .B2(n5764), .ZN(n5380)
         );
  AOI21_X1 U6095 ( .B1(n5766), .B2(n5390), .A(n5380), .ZN(n5382) );
  INV_X1 U6096 ( .A(n5932), .ZN(n5961) );
  NAND2_X1 U6097 ( .A1(n5465), .A2(n5961), .ZN(n5381) );
  OAI211_X1 U6098 ( .C1(n5394), .C2(n5383), .A(n5382), .B(n5381), .ZN(U3119)
         );
  INV_X1 U6099 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5387) );
  OAI22_X1 U6100 ( .A1(n5918), .A2(n5988), .B1(n5388), .B2(n5753), .ZN(n5384)
         );
  AOI21_X1 U6101 ( .B1(n5755), .B2(n5390), .A(n5384), .ZN(n5386) );
  INV_X1 U6102 ( .A(n5937), .ZN(n5985) );
  NAND2_X1 U6103 ( .A1(n5465), .A2(n5985), .ZN(n5385) );
  OAI211_X1 U6104 ( .C1(n5394), .C2(n5387), .A(n5386), .B(n5385), .ZN(U3118)
         );
  INV_X1 U6105 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5393) );
  OAI22_X1 U6106 ( .A1(n5918), .A2(n5977), .B1(n5388), .B2(n5772), .ZN(n5389)
         );
  AOI21_X1 U6107 ( .B1(n5776), .B2(n5390), .A(n5389), .ZN(n5392) );
  INV_X1 U6108 ( .A(n5949), .ZN(n5975) );
  NAND2_X1 U6109 ( .A1(n5465), .A2(n5975), .ZN(n5391) );
  OAI211_X1 U6110 ( .C1(n5394), .C2(n5393), .A(n5392), .B(n5391), .ZN(U3117)
         );
  AND2_X1 U6111 ( .A1(n3661), .A2(n4263), .ZN(n5867) );
  NOR2_X1 U6112 ( .A1(n5395), .A2(n7566), .ZN(n5605) );
  AOI21_X1 U6113 ( .B1(n5867), .B2(n5470), .A(n5605), .ZN(n5402) );
  OR2_X1 U6114 ( .A1(n5402), .A2(n5870), .ZN(n5398) );
  INV_X1 U6115 ( .A(n5400), .ZN(n5396) );
  NAND2_X1 U6116 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5396), .ZN(n5397) );
  NAND2_X1 U6117 ( .A1(n5398), .A2(n5397), .ZN(n5604) );
  INV_X1 U6118 ( .A(n5604), .ZN(n5417) );
  OR2_X1 U6119 ( .A1(n5870), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5869) );
  OAI21_X1 U6120 ( .B1(n5404), .B2(n6976), .A(n5869), .ZN(n5401) );
  AOI22_X1 U6121 ( .A1(n5402), .A2(n5401), .B1(n5870), .B2(n5400), .ZN(n5403)
         );
  NAND2_X1 U6122 ( .A1(n5873), .A2(n5403), .ZN(n5609) );
  NAND2_X1 U6123 ( .A1(n5609), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5407)
         );
  OAI22_X1 U6124 ( .A1(n5993), .A2(n5786), .B1(n5603), .B2(n5787), .ZN(n5405)
         );
  AOI21_X1 U6125 ( .B1(n5991), .B2(n5605), .A(n5405), .ZN(n5406) );
  OAI211_X1 U6126 ( .C1(n5417), .C2(n5997), .A(n5407), .B(n5406), .ZN(U3145)
         );
  NAND2_X1 U6127 ( .A1(n5609), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5410)
         );
  OAI22_X1 U6128 ( .A1(n6000), .A2(n5786), .B1(n5603), .B2(n5779), .ZN(n5408)
         );
  AOI21_X1 U6129 ( .B1(n5998), .B2(n5605), .A(n5408), .ZN(n5409) );
  OAI211_X1 U6130 ( .C1(n5417), .C2(n6004), .A(n5410), .B(n5409), .ZN(U3146)
         );
  NAND2_X1 U6131 ( .A1(n5609), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5413)
         );
  OAI22_X1 U6132 ( .A1(n6419), .A2(n5786), .B1(n5603), .B2(n6410), .ZN(n5411)
         );
  AOI21_X1 U6133 ( .B1(n6014), .B2(n5605), .A(n5411), .ZN(n5412) );
  OAI211_X1 U6134 ( .C1(n5417), .C2(n6021), .A(n5413), .B(n5412), .ZN(U3147)
         );
  NAND2_X1 U6135 ( .A1(n5609), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5416)
         );
  OAI22_X1 U6136 ( .A1(n6007), .A2(n5786), .B1(n5603), .B2(n5758), .ZN(n5414)
         );
  AOI21_X1 U6137 ( .B1(n6005), .B2(n5605), .A(n5414), .ZN(n5415) );
  OAI211_X1 U6138 ( .C1(n5417), .C2(n6011), .A(n5416), .B(n5415), .ZN(U3144)
         );
  INV_X1 U6139 ( .A(n5609), .ZN(n5433) );
  INV_X1 U6140 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n5422) );
  OR2_X1 U6141 ( .A1(n5603), .A2(n5932), .ZN(n5419) );
  NAND2_X1 U6142 ( .A1(n5604), .A2(n5957), .ZN(n5418) );
  OAI211_X1 U6143 ( .C1(n5786), .C2(n5963), .A(n5419), .B(n5418), .ZN(n5420)
         );
  AOI21_X1 U6144 ( .B1(n5766), .B2(n5605), .A(n5420), .ZN(n5421) );
  OAI21_X1 U6145 ( .B1(n5433), .B2(n5422), .A(n5421), .ZN(U3143) );
  INV_X1 U6146 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n5427) );
  OR2_X1 U6147 ( .A1(n5603), .A2(n5949), .ZN(n5424) );
  NAND2_X1 U6148 ( .A1(n5604), .A2(n5971), .ZN(n5423) );
  OAI211_X1 U6149 ( .C1(n5786), .C2(n5977), .A(n5424), .B(n5423), .ZN(n5425)
         );
  AOI21_X1 U6150 ( .B1(n5776), .B2(n5605), .A(n5425), .ZN(n5426) );
  OAI21_X1 U6151 ( .B1(n5433), .B2(n5427), .A(n5426), .ZN(U3141) );
  INV_X1 U6152 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n5432) );
  OR2_X1 U6153 ( .A1(n5603), .A2(n5937), .ZN(n5429) );
  NAND2_X1 U6154 ( .A1(n5604), .A2(n5979), .ZN(n5428) );
  OAI211_X1 U6155 ( .C1(n5786), .C2(n5988), .A(n5429), .B(n5428), .ZN(n5430)
         );
  AOI21_X1 U6156 ( .B1(n5755), .B2(n5605), .A(n5430), .ZN(n5431) );
  OAI21_X1 U6157 ( .B1(n5433), .B2(n5432), .A(n5431), .ZN(U3142) );
  NAND2_X1 U6158 ( .A1(n4255), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5717) );
  NOR2_X1 U6159 ( .A1(n5126), .A2(n5717), .ZN(n5716) );
  INV_X1 U6160 ( .A(n5716), .ZN(n5611) );
  OAI21_X1 U6161 ( .B1(n5611), .B2(n5617), .A(n5875), .ZN(n5438) );
  AND2_X1 U6162 ( .A1(n5028), .A2(n5125), .ZN(n5667) );
  AND2_X1 U6163 ( .A1(n5667), .A2(n3661), .ZN(n5567) );
  NAND3_X1 U6164 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n5718), .ZN(n5563) );
  NOR2_X1 U6165 ( .A1(n3937), .A2(n5563), .ZN(n5435) );
  AOI21_X1 U6166 ( .B1(n5567), .B2(n4263), .A(n5435), .ZN(n5439) );
  OAI22_X1 U6167 ( .A1(n5438), .A2(n5439), .B1(n5563), .B2(n7584), .ZN(n5434)
         );
  INV_X1 U6168 ( .A(n5435), .ZN(n5463) );
  AND2_X1 U6169 ( .A1(n5436), .A2(n5804), .ZN(n5618) );
  OAI22_X1 U6170 ( .A1(n5966), .A2(n5463), .B1(n5942), .B2(n5590), .ZN(n5437)
         );
  AOI21_X1 U6171 ( .B1(n5944), .B2(n5465), .A(n5437), .ZN(n5444) );
  INV_X1 U6172 ( .A(n5563), .ZN(n5442) );
  INV_X1 U6173 ( .A(n5438), .ZN(n5440) );
  NAND2_X1 U6174 ( .A1(n5440), .A2(n5439), .ZN(n5441) );
  NAND2_X1 U6175 ( .A1(n5466), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n5443)
         );
  OAI211_X1 U6176 ( .C1(n5469), .C2(n5748), .A(n5444), .B(n5443), .ZN(U3108)
         );
  OAI22_X1 U6177 ( .A1(n5789), .A2(n5463), .B1(n5787), .B2(n5590), .ZN(n5445)
         );
  AOI21_X1 U6178 ( .B1(n5673), .B2(n5465), .A(n5445), .ZN(n5447) );
  NAND2_X1 U6179 ( .A1(n5466), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n5446)
         );
  OAI211_X1 U6180 ( .C1(n5469), .C2(n5997), .A(n5447), .B(n5446), .ZN(U3113)
         );
  OAI22_X1 U6181 ( .A1(n6413), .A2(n5463), .B1(n6410), .B2(n5590), .ZN(n5448)
         );
  AOI21_X1 U6182 ( .B1(n5698), .B2(n5465), .A(n5448), .ZN(n5450) );
  NAND2_X1 U6183 ( .A1(n5466), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n5449)
         );
  OAI211_X1 U6184 ( .C1(n5469), .C2(n6021), .A(n5450), .B(n5449), .ZN(U3115)
         );
  OAI22_X1 U6185 ( .A1(n5959), .A2(n5463), .B1(n5932), .B2(n5590), .ZN(n5451)
         );
  AOI21_X1 U6186 ( .B1(n5934), .B2(n5465), .A(n5451), .ZN(n5453) );
  NAND2_X1 U6187 ( .A1(n5466), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n5452)
         );
  OAI211_X1 U6188 ( .C1(n5469), .C2(n5764), .A(n5453), .B(n5452), .ZN(U3111)
         );
  OAI22_X1 U6189 ( .A1(n5759), .A2(n5463), .B1(n5758), .B2(n5590), .ZN(n5454)
         );
  AOI21_X1 U6190 ( .B1(n5681), .B2(n5465), .A(n5454), .ZN(n5456) );
  NAND2_X1 U6191 ( .A1(n5466), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n5455)
         );
  OAI211_X1 U6192 ( .C1(n5469), .C2(n6011), .A(n5456), .B(n5455), .ZN(U3112)
         );
  OAI22_X1 U6193 ( .A1(n5973), .A2(n5463), .B1(n5949), .B2(n5590), .ZN(n5457)
         );
  AOI21_X1 U6194 ( .B1(n5952), .B2(n5465), .A(n5457), .ZN(n5459) );
  NAND2_X1 U6195 ( .A1(n5466), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n5458)
         );
  OAI211_X1 U6196 ( .C1(n5469), .C2(n5772), .A(n5459), .B(n5458), .ZN(U3109)
         );
  OAI22_X1 U6197 ( .A1(n5780), .A2(n5463), .B1(n5779), .B2(n5590), .ZN(n5460)
         );
  AOI21_X1 U6198 ( .B1(n5677), .B2(n5465), .A(n5460), .ZN(n5462) );
  NAND2_X1 U6199 ( .A1(n5466), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n5461)
         );
  OAI211_X1 U6200 ( .C1(n5469), .C2(n6004), .A(n5462), .B(n5461), .ZN(U3114)
         );
  OAI22_X1 U6201 ( .A1(n5983), .A2(n5463), .B1(n5937), .B2(n5590), .ZN(n5464)
         );
  AOI21_X1 U6202 ( .B1(n5939), .B2(n5465), .A(n5464), .ZN(n5468) );
  NAND2_X1 U6203 ( .A1(n5466), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n5467)
         );
  OAI211_X1 U6204 ( .C1(n5469), .C2(n5753), .A(n5468), .B(n5467), .ZN(U3110)
         );
  OR2_X1 U6205 ( .A1(n3661), .A2(n7425), .ZN(n5614) );
  INV_X1 U6206 ( .A(n5955), .ZN(n5536) );
  AOI21_X1 U6207 ( .B1(n5501), .B2(n5470), .A(n5536), .ZN(n5474) );
  NOR2_X1 U6208 ( .A1(n5471), .A2(n5870), .ZN(n5475) );
  INV_X1 U6209 ( .A(n5475), .ZN(n5472) );
  OAI22_X1 U6210 ( .A1(n5474), .A2(n5472), .B1(n5473), .B2(n7584), .ZN(n5946)
         );
  INV_X1 U6211 ( .A(n5946), .ZN(n5539) );
  AOI22_X1 U6212 ( .A1(n5475), .A2(n5474), .B1(n5870), .B2(n5473), .ZN(n5476)
         );
  NAND2_X1 U6213 ( .A1(n5873), .A2(n5476), .ZN(n5947) );
  NAND2_X1 U6214 ( .A1(n5947), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n5479) );
  OAI22_X1 U6215 ( .A1(n6411), .A2(n5993), .B1(n5950), .B2(n5787), .ZN(n5477)
         );
  AOI21_X1 U6216 ( .B1(n5991), .B2(n5536), .A(n5477), .ZN(n5478) );
  OAI211_X1 U6217 ( .C1(n5539), .C2(n5997), .A(n5479), .B(n5478), .ZN(U3081)
         );
  OAI21_X1 U6218 ( .B1(n5489), .B2(n5870), .A(n5869), .ZN(n5484) );
  INV_X1 U6219 ( .A(n5484), .ZN(n5482) );
  NOR2_X1 U6220 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5736) );
  NAND2_X1 U6221 ( .A1(n5736), .A2(n5481), .ZN(n5483) );
  NOR2_X1 U6222 ( .A1(n3937), .A2(n5483), .ZN(n5488) );
  AOI21_X1 U6223 ( .B1(n5501), .B2(n5866), .A(n5488), .ZN(n5485) );
  OAI22_X1 U6224 ( .A1(n5482), .A2(n5485), .B1(n5483), .B2(n7584), .ZN(n5978)
         );
  INV_X1 U6225 ( .A(n5978), .ZN(n5553) );
  AOI22_X1 U6226 ( .A1(n5485), .A2(n5484), .B1(n5870), .B2(n5483), .ZN(n5486)
         );
  NAND2_X1 U6227 ( .A1(n5873), .A2(n5486), .ZN(n5980) );
  NAND2_X1 U6228 ( .A1(n5980), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n5492) );
  INV_X1 U6229 ( .A(n5488), .ZN(n5982) );
  OAI22_X1 U6230 ( .A1(n5789), .A2(n5982), .B1(n5956), .B2(n5787), .ZN(n5490)
         );
  AOI21_X1 U6231 ( .B1(n5657), .B2(n5673), .A(n5490), .ZN(n5491) );
  OAI211_X1 U6232 ( .C1(n5553), .C2(n5997), .A(n5492), .B(n5491), .ZN(U3033)
         );
  NAND2_X1 U6233 ( .A1(n5947), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n5495) );
  OAI22_X1 U6234 ( .A1(n6411), .A2(n6419), .B1(n5950), .B2(n6410), .ZN(n5493)
         );
  AOI21_X1 U6235 ( .B1(n6014), .B2(n5536), .A(n5493), .ZN(n5494) );
  OAI211_X1 U6236 ( .C1(n5539), .C2(n6021), .A(n5495), .B(n5494), .ZN(U3083)
         );
  NAND2_X1 U6237 ( .A1(n5980), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n5498) );
  OAI22_X1 U6238 ( .A1(n5759), .A2(n5982), .B1(n5758), .B2(n5956), .ZN(n5496)
         );
  AOI21_X1 U6239 ( .B1(n5657), .B2(n5681), .A(n5496), .ZN(n5497) );
  OAI211_X1 U6240 ( .C1(n5553), .C2(n6011), .A(n5498), .B(n5497), .ZN(U3032)
         );
  NAND2_X1 U6241 ( .A1(n5499), .A2(n5875), .ZN(n5500) );
  NAND2_X1 U6242 ( .A1(n5500), .A2(n5869), .ZN(n5507) );
  NOR2_X1 U6243 ( .A1(n3937), .A2(n5506), .ZN(n5898) );
  AOI21_X1 U6244 ( .B1(n5501), .B2(n5516), .A(n5898), .ZN(n5508) );
  INV_X1 U6245 ( .A(n5508), .ZN(n5502) );
  NAND2_X1 U6246 ( .A1(n5507), .A2(n5502), .ZN(n5505) );
  INV_X1 U6247 ( .A(n5506), .ZN(n5503) );
  NAND2_X1 U6248 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5503), .ZN(n5504) );
  NAND2_X1 U6249 ( .A1(n5505), .A2(n5504), .ZN(n5923) );
  AOI22_X1 U6250 ( .A1(n5508), .A2(n5507), .B1(n5870), .B2(n5506), .ZN(n5509)
         );
  NAND2_X1 U6251 ( .A1(n5873), .A2(n5509), .ZN(n5924) );
  NAND2_X1 U6252 ( .A1(n5924), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n5512) );
  OAI22_X1 U6253 ( .A1(n6007), .A2(n5899), .B1(n5926), .B2(n5758), .ZN(n5510)
         );
  AOI21_X1 U6254 ( .B1(n6005), .B2(n5898), .A(n5510), .ZN(n5511) );
  OAI211_X1 U6255 ( .C1(n5557), .C2(n6011), .A(n5512), .B(n5511), .ZN(U3064)
         );
  NAND2_X1 U6256 ( .A1(n5947), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n5515) );
  OAI22_X1 U6257 ( .A1(n6411), .A2(n6007), .B1(n5950), .B2(n5758), .ZN(n5513)
         );
  AOI21_X1 U6258 ( .B1(n6005), .B2(n5536), .A(n5513), .ZN(n5514) );
  OAI211_X1 U6259 ( .C1(n5539), .C2(n6011), .A(n5515), .B(n5514), .ZN(U3080)
         );
  NOR2_X1 U6260 ( .A1(n3937), .A2(n5519), .ZN(n5893) );
  AOI21_X1 U6261 ( .B1(n5867), .B2(n5516), .A(n5893), .ZN(n5521) );
  NOR2_X1 U6262 ( .A1(n5517), .A2(n5870), .ZN(n5520) );
  INV_X1 U6263 ( .A(n5520), .ZN(n5518) );
  OAI22_X1 U6264 ( .A1(n5521), .A2(n5518), .B1(n5519), .B2(n7584), .ZN(n5915)
         );
  INV_X1 U6265 ( .A(n5915), .ZN(n5546) );
  AOI22_X1 U6266 ( .A1(n5521), .A2(n5520), .B1(n5870), .B2(n5519), .ZN(n5522)
         );
  NAND2_X1 U6267 ( .A1(n5873), .A2(n5522), .ZN(n5916) );
  NAND2_X1 U6268 ( .A1(n5916), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n5525)
         );
  OAI22_X1 U6269 ( .A1(n5993), .A2(n5894), .B1(n5918), .B2(n5787), .ZN(n5523)
         );
  AOI21_X1 U6270 ( .B1(n5991), .B2(n5893), .A(n5523), .ZN(n5524) );
  OAI211_X1 U6271 ( .C1(n5546), .C2(n5997), .A(n5525), .B(n5524), .ZN(U3129)
         );
  NAND2_X1 U6272 ( .A1(n5916), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n5528)
         );
  OAI22_X1 U6273 ( .A1(n6007), .A2(n5894), .B1(n5918), .B2(n5758), .ZN(n5526)
         );
  AOI21_X1 U6274 ( .B1(n6005), .B2(n5893), .A(n5526), .ZN(n5527) );
  OAI211_X1 U6275 ( .C1(n5546), .C2(n6011), .A(n5528), .B(n5527), .ZN(U3128)
         );
  NAND2_X1 U6276 ( .A1(n5924), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n5531) );
  OAI22_X1 U6277 ( .A1(n5993), .A2(n5899), .B1(n5926), .B2(n5787), .ZN(n5529)
         );
  AOI21_X1 U6278 ( .B1(n5991), .B2(n5898), .A(n5529), .ZN(n5530) );
  OAI211_X1 U6279 ( .C1(n5557), .C2(n5997), .A(n5531), .B(n5530), .ZN(U3065)
         );
  NAND2_X1 U6280 ( .A1(n5924), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5534) );
  OAI22_X1 U6281 ( .A1(n6419), .A2(n5899), .B1(n5926), .B2(n6410), .ZN(n5532)
         );
  AOI21_X1 U6282 ( .B1(n6014), .B2(n5898), .A(n5532), .ZN(n5533) );
  OAI211_X1 U6283 ( .C1(n5557), .C2(n6021), .A(n5534), .B(n5533), .ZN(U3067)
         );
  NAND2_X1 U6284 ( .A1(n5947), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n5538) );
  OAI22_X1 U6285 ( .A1(n6411), .A2(n6000), .B1(n5950), .B2(n5779), .ZN(n5535)
         );
  AOI21_X1 U6286 ( .B1(n5998), .B2(n5536), .A(n5535), .ZN(n5537) );
  OAI211_X1 U6287 ( .C1(n5539), .C2(n6004), .A(n5538), .B(n5537), .ZN(U3082)
         );
  NAND2_X1 U6288 ( .A1(n5916), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n5542)
         );
  OAI22_X1 U6289 ( .A1(n6419), .A2(n5894), .B1(n5918), .B2(n6410), .ZN(n5540)
         );
  AOI21_X1 U6290 ( .B1(n6014), .B2(n5893), .A(n5540), .ZN(n5541) );
  OAI211_X1 U6291 ( .C1(n5546), .C2(n6021), .A(n5542), .B(n5541), .ZN(U3131)
         );
  NAND2_X1 U6292 ( .A1(n5916), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n5545)
         );
  OAI22_X1 U6293 ( .A1(n6000), .A2(n5894), .B1(n5918), .B2(n5779), .ZN(n5543)
         );
  AOI21_X1 U6294 ( .B1(n5998), .B2(n5893), .A(n5543), .ZN(n5544) );
  OAI211_X1 U6295 ( .C1(n5546), .C2(n6004), .A(n5545), .B(n5544), .ZN(U3130)
         );
  NAND2_X1 U6296 ( .A1(n5980), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5549) );
  OAI22_X1 U6297 ( .A1(n5780), .A2(n5982), .B1(n5956), .B2(n5779), .ZN(n5547)
         );
  AOI21_X1 U6298 ( .B1(n5657), .B2(n5677), .A(n5547), .ZN(n5548) );
  OAI211_X1 U6299 ( .C1(n5553), .C2(n6004), .A(n5549), .B(n5548), .ZN(U3034)
         );
  NAND2_X1 U6300 ( .A1(n5980), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5552) );
  OAI22_X1 U6301 ( .A1(n6413), .A2(n5982), .B1(n6410), .B2(n5956), .ZN(n5550)
         );
  AOI21_X1 U6302 ( .B1(n5698), .B2(n5657), .A(n5550), .ZN(n5551) );
  OAI211_X1 U6303 ( .C1(n5553), .C2(n6021), .A(n5552), .B(n5551), .ZN(U3035)
         );
  NAND2_X1 U6304 ( .A1(n5924), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5556) );
  OAI22_X1 U6305 ( .A1(n6000), .A2(n5899), .B1(n5926), .B2(n5779), .ZN(n5554)
         );
  AOI21_X1 U6306 ( .B1(n5998), .B2(n5898), .A(n5554), .ZN(n5555) );
  OAI211_X1 U6307 ( .C1(n5557), .C2(n6004), .A(n5556), .B(n5555), .ZN(U3066)
         );
  NAND2_X1 U6308 ( .A1(n6016), .A2(n5590), .ZN(n5558) );
  NAND2_X1 U6309 ( .A1(n5558), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5559) );
  NAND2_X1 U6310 ( .A1(n5559), .A2(n5875), .ZN(n5566) );
  INV_X1 U6311 ( .A(n5566), .ZN(n5562) );
  INV_X1 U6312 ( .A(n5560), .ZN(n5743) );
  OR2_X1 U6313 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5563), .ZN(n5591)
         );
  AOI211_X1 U6314 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5591), .A(n5564), .B(
        n5738), .ZN(n5565) );
  NAND2_X1 U6315 ( .A1(n5589), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5570)
         );
  OAI22_X1 U6316 ( .A1(n5759), .A2(n5591), .B1(n6007), .B2(n5590), .ZN(n5568)
         );
  AOI21_X1 U6317 ( .B1(n6009), .B2(n5593), .A(n5568), .ZN(n5569) );
  OAI211_X1 U6318 ( .C1(n5596), .C2(n6011), .A(n5570), .B(n5569), .ZN(U3104)
         );
  NAND2_X1 U6319 ( .A1(n5589), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5573)
         );
  OAI22_X1 U6320 ( .A1(n5973), .A2(n5591), .B1(n5977), .B2(n5590), .ZN(n5571)
         );
  AOI21_X1 U6321 ( .B1(n5975), .B2(n5593), .A(n5571), .ZN(n5572) );
  OAI211_X1 U6322 ( .C1(n5596), .C2(n5772), .A(n5573), .B(n5572), .ZN(U3101)
         );
  NAND2_X1 U6323 ( .A1(n5589), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5576)
         );
  OAI22_X1 U6324 ( .A1(n5966), .A2(n5591), .B1(n5970), .B2(n5590), .ZN(n5574)
         );
  AOI21_X1 U6325 ( .B1(n5968), .B2(n5593), .A(n5574), .ZN(n5575) );
  OAI211_X1 U6326 ( .C1(n5596), .C2(n5748), .A(n5576), .B(n5575), .ZN(U3100)
         );
  NAND2_X1 U6327 ( .A1(n5589), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5579)
         );
  OAI22_X1 U6328 ( .A1(n5983), .A2(n5591), .B1(n5988), .B2(n5590), .ZN(n5577)
         );
  AOI21_X1 U6329 ( .B1(n5985), .B2(n5593), .A(n5577), .ZN(n5578) );
  OAI211_X1 U6330 ( .C1(n5596), .C2(n5753), .A(n5579), .B(n5578), .ZN(U3102)
         );
  NAND2_X1 U6331 ( .A1(n5589), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5582)
         );
  OAI22_X1 U6332 ( .A1(n5789), .A2(n5591), .B1(n5993), .B2(n5590), .ZN(n5580)
         );
  AOI21_X1 U6333 ( .B1(n5995), .B2(n5593), .A(n5580), .ZN(n5581) );
  OAI211_X1 U6334 ( .C1(n5596), .C2(n5997), .A(n5582), .B(n5581), .ZN(U3105)
         );
  NAND2_X1 U6335 ( .A1(n5589), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5585)
         );
  OAI22_X1 U6336 ( .A1(n5959), .A2(n5591), .B1(n5963), .B2(n5590), .ZN(n5583)
         );
  AOI21_X1 U6337 ( .B1(n5961), .B2(n5593), .A(n5583), .ZN(n5584) );
  OAI211_X1 U6338 ( .C1(n5596), .C2(n5764), .A(n5585), .B(n5584), .ZN(U3103)
         );
  NAND2_X1 U6339 ( .A1(n5589), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5588)
         );
  OAI22_X1 U6340 ( .A1(n5780), .A2(n5591), .B1(n6000), .B2(n5590), .ZN(n5586)
         );
  AOI21_X1 U6341 ( .B1(n6002), .B2(n5593), .A(n5586), .ZN(n5587) );
  OAI211_X1 U6342 ( .C1(n5596), .C2(n6004), .A(n5588), .B(n5587), .ZN(U3106)
         );
  NAND2_X1 U6343 ( .A1(n5589), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5595)
         );
  OAI22_X1 U6344 ( .A1(n6413), .A2(n5591), .B1(n6419), .B2(n5590), .ZN(n5592)
         );
  AOI21_X1 U6345 ( .B1(n6018), .B2(n5593), .A(n5592), .ZN(n5594) );
  OAI211_X1 U6346 ( .C1(n5596), .C2(n6021), .A(n5595), .B(n5594), .ZN(U3107)
         );
  INV_X1 U6347 ( .A(n5147), .ZN(n5600) );
  AOI21_X1 U6348 ( .B1(n5106), .B2(n5598), .A(n5597), .ZN(n5599) );
  NOR2_X1 U6349 ( .A1(n5600), .A2(n5599), .ZN(n7498) );
  INV_X1 U6350 ( .A(n7498), .ZN(n5601) );
  OAI222_X1 U6351 ( .A1(n6833), .A2(n5602), .B1(n6829), .B2(n4304), .C1(n6831), 
        .C2(n5601), .ZN(U2884) );
  NOR2_X1 U6352 ( .A1(n5603), .A2(n5942), .ZN(n5608) );
  AOI22_X1 U6353 ( .A1(n5750), .A2(n5605), .B1(n5964), .B2(n5604), .ZN(n5606)
         );
  OAI21_X1 U6354 ( .B1(n5786), .B2(n5970), .A(n5606), .ZN(n5607) );
  AOI211_X1 U6355 ( .C1(n5609), .C2(INSTQUEUE_REG_15__0__SCAN_IN), .A(n5608), 
        .B(n5607), .ZN(n5610) );
  INV_X1 U6356 ( .A(n5610), .ZN(U3140) );
  OAI21_X1 U6357 ( .B1(n5611), .B2(n5128), .A(n5875), .ZN(n5622) );
  INV_X1 U6358 ( .A(n5622), .ZN(n5616) );
  INV_X1 U6359 ( .A(n5667), .ZN(n5613) );
  NAND2_X1 U6360 ( .A1(n5736), .A2(n5612), .ZN(n5644) );
  OAI21_X1 U6361 ( .B1(n5614), .B2(n5613), .A(n5644), .ZN(n5621) );
  NAND2_X1 U6362 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n5736), .ZN(n5660) );
  INV_X1 U6363 ( .A(n5660), .ZN(n5615) );
  OAI22_X1 U6364 ( .A1(n6413), .A2(n5644), .B1(n6419), .B2(n5643), .ZN(n5619)
         );
  AOI21_X1 U6365 ( .B1(n6018), .B2(n5697), .A(n5619), .ZN(n5624) );
  NAND2_X1 U6366 ( .A1(n5660), .A2(n5870), .ZN(n5620) );
  OAI211_X1 U6367 ( .C1(n5622), .C2(n5621), .A(n5873), .B(n5620), .ZN(n5646)
         );
  NAND2_X1 U6368 ( .A1(n5646), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5623) );
  OAI211_X1 U6369 ( .C1(n5649), .C2(n6021), .A(n5624), .B(n5623), .ZN(U3051)
         );
  OAI22_X1 U6370 ( .A1(n5780), .A2(n5644), .B1(n6000), .B2(n5643), .ZN(n5625)
         );
  AOI21_X1 U6371 ( .B1(n6002), .B2(n5697), .A(n5625), .ZN(n5627) );
  NAND2_X1 U6372 ( .A1(n5646), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5626) );
  OAI211_X1 U6373 ( .C1(n5649), .C2(n6004), .A(n5627), .B(n5626), .ZN(U3050)
         );
  OAI22_X1 U6374 ( .A1(n5983), .A2(n5644), .B1(n5988), .B2(n5643), .ZN(n5628)
         );
  AOI21_X1 U6375 ( .B1(n5985), .B2(n5697), .A(n5628), .ZN(n5630) );
  NAND2_X1 U6376 ( .A1(n5646), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n5629) );
  OAI211_X1 U6377 ( .C1(n5649), .C2(n5753), .A(n5630), .B(n5629), .ZN(U3046)
         );
  OAI22_X1 U6378 ( .A1(n5759), .A2(n5644), .B1(n6007), .B2(n5643), .ZN(n5631)
         );
  AOI21_X1 U6379 ( .B1(n6009), .B2(n5697), .A(n5631), .ZN(n5633) );
  NAND2_X1 U6380 ( .A1(n5646), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5632) );
  OAI211_X1 U6381 ( .C1(n5649), .C2(n6011), .A(n5633), .B(n5632), .ZN(U3048)
         );
  OAI22_X1 U6382 ( .A1(n5789), .A2(n5644), .B1(n5993), .B2(n5643), .ZN(n5634)
         );
  AOI21_X1 U6383 ( .B1(n5995), .B2(n5697), .A(n5634), .ZN(n5636) );
  NAND2_X1 U6384 ( .A1(n5646), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5635) );
  OAI211_X1 U6385 ( .C1(n5649), .C2(n5997), .A(n5636), .B(n5635), .ZN(U3049)
         );
  OAI22_X1 U6386 ( .A1(n5973), .A2(n5644), .B1(n5977), .B2(n5643), .ZN(n5637)
         );
  AOI21_X1 U6387 ( .B1(n5975), .B2(n5697), .A(n5637), .ZN(n5639) );
  NAND2_X1 U6388 ( .A1(n5646), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n5638) );
  OAI211_X1 U6389 ( .C1(n5649), .C2(n5772), .A(n5639), .B(n5638), .ZN(U3045)
         );
  OAI22_X1 U6390 ( .A1(n5966), .A2(n5644), .B1(n5970), .B2(n5643), .ZN(n5640)
         );
  AOI21_X1 U6391 ( .B1(n5968), .B2(n5697), .A(n5640), .ZN(n5642) );
  NAND2_X1 U6392 ( .A1(n5646), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n5641) );
  OAI211_X1 U6393 ( .C1(n5649), .C2(n5748), .A(n5642), .B(n5641), .ZN(U3044)
         );
  OAI22_X1 U6394 ( .A1(n5959), .A2(n5644), .B1(n5963), .B2(n5643), .ZN(n5645)
         );
  AOI21_X1 U6395 ( .B1(n5961), .B2(n5697), .A(n5645), .ZN(n5648) );
  NAND2_X1 U6396 ( .A1(n5646), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5647) );
  OAI211_X1 U6397 ( .C1(n5649), .C2(n5764), .A(n5648), .B(n5647), .ZN(U3047)
         );
  INV_X1 U6398 ( .A(n5650), .ZN(n7475) );
  NOR2_X1 U6399 ( .A1(n5652), .A2(n5651), .ZN(n5653) );
  OR2_X1 U6400 ( .A1(n5654), .A2(n5653), .ZN(n7471) );
  OAI22_X1 U6401 ( .A1(n3659), .A2(n7471), .B1(n7470), .B2(n7259), .ZN(n5655)
         );
  AOI21_X1 U6402 ( .B1(n7475), .B2(n6793), .A(n5655), .ZN(n5656) );
  INV_X1 U6403 ( .A(n5656), .ZN(U2854) );
  OAI21_X1 U6404 ( .B1(n5657), .B2(n5697), .A(n5869), .ZN(n5659) );
  NAND2_X1 U6405 ( .A1(n7438), .A2(n5667), .ZN(n5658) );
  AOI21_X1 U6406 ( .B1(n5659), .B2(n5658), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n5663) );
  NOR2_X1 U6407 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5660), .ZN(n5664)
         );
  INV_X1 U6408 ( .A(n5738), .ZN(n5661) );
  NAND2_X1 U6409 ( .A1(n5693), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5671) );
  INV_X1 U6410 ( .A(n5664), .ZN(n5694) );
  INV_X1 U6411 ( .A(n5665), .ZN(n5666) );
  AOI22_X1 U6412 ( .A1(n5668), .A2(n5667), .B1(n5743), .B2(n5666), .ZN(n5695)
         );
  OAI22_X1 U6413 ( .A1(n5959), .A2(n5694), .B1(n5695), .B2(n5764), .ZN(n5669)
         );
  AOI21_X1 U6414 ( .B1(n5934), .B2(n5697), .A(n5669), .ZN(n5670) );
  OAI211_X1 U6415 ( .C1(n5932), .C2(n5989), .A(n5671), .B(n5670), .ZN(U3039)
         );
  NAND2_X1 U6416 ( .A1(n5693), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5675) );
  OAI22_X1 U6417 ( .A1(n5997), .A2(n5695), .B1(n5789), .B2(n5694), .ZN(n5672)
         );
  AOI21_X1 U6418 ( .B1(n5673), .B2(n5697), .A(n5672), .ZN(n5674) );
  OAI211_X1 U6419 ( .C1(n5787), .C2(n5989), .A(n5675), .B(n5674), .ZN(U3041)
         );
  NAND2_X1 U6420 ( .A1(n5693), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5679) );
  OAI22_X1 U6421 ( .A1(n6004), .A2(n5695), .B1(n5780), .B2(n5694), .ZN(n5676)
         );
  AOI21_X1 U6422 ( .B1(n5677), .B2(n5697), .A(n5676), .ZN(n5678) );
  OAI211_X1 U6423 ( .C1(n5779), .C2(n5989), .A(n5679), .B(n5678), .ZN(U3042)
         );
  NAND2_X1 U6424 ( .A1(n5693), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5683) );
  OAI22_X1 U6425 ( .A1(n6011), .A2(n5695), .B1(n5759), .B2(n5694), .ZN(n5680)
         );
  AOI21_X1 U6426 ( .B1(n5681), .B2(n5697), .A(n5680), .ZN(n5682) );
  OAI211_X1 U6427 ( .C1(n5758), .C2(n5989), .A(n5683), .B(n5682), .ZN(U3040)
         );
  NAND2_X1 U6428 ( .A1(n5693), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5686) );
  OAI22_X1 U6429 ( .A1(n5983), .A2(n5694), .B1(n5695), .B2(n5753), .ZN(n5684)
         );
  AOI21_X1 U6430 ( .B1(n5939), .B2(n5697), .A(n5684), .ZN(n5685) );
  OAI211_X1 U6431 ( .C1(n5937), .C2(n5989), .A(n5686), .B(n5685), .ZN(U3038)
         );
  NAND2_X1 U6432 ( .A1(n5693), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5689) );
  OAI22_X1 U6433 ( .A1(n5973), .A2(n5694), .B1(n5695), .B2(n5772), .ZN(n5687)
         );
  AOI21_X1 U6434 ( .B1(n5952), .B2(n5697), .A(n5687), .ZN(n5688) );
  OAI211_X1 U6435 ( .C1(n5949), .C2(n5989), .A(n5689), .B(n5688), .ZN(U3037)
         );
  NAND2_X1 U6436 ( .A1(n5693), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5692) );
  OAI22_X1 U6437 ( .A1(n5966), .A2(n5694), .B1(n5695), .B2(n5748), .ZN(n5690)
         );
  AOI21_X1 U6438 ( .B1(n5944), .B2(n5697), .A(n5690), .ZN(n5691) );
  OAI211_X1 U6439 ( .C1(n5942), .C2(n5989), .A(n5692), .B(n5691), .ZN(U3036)
         );
  NAND2_X1 U6440 ( .A1(n5693), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5700) );
  OAI22_X1 U6441 ( .A1(n6021), .A2(n5695), .B1(n6413), .B2(n5694), .ZN(n5696)
         );
  AOI21_X1 U6442 ( .B1(n5698), .B2(n5697), .A(n5696), .ZN(n5699) );
  OAI211_X1 U6443 ( .C1(n5989), .C2(n6410), .A(n5700), .B(n5699), .ZN(U3043)
         );
  NAND2_X1 U6444 ( .A1(n5702), .A2(n5701), .ZN(n5703) );
  AND2_X1 U6445 ( .A1(n5704), .A2(n5703), .ZN(n7369) );
  INV_X1 U6446 ( .A(n7369), .ZN(n7490) );
  OAI22_X1 U6447 ( .A1(n3659), .A2(n7490), .B1(n5705), .B2(n7259), .ZN(n5706)
         );
  AOI21_X1 U6448 ( .B1(n7498), .B2(n6793), .A(n5706), .ZN(n5707) );
  INV_X1 U6449 ( .A(n5707), .ZN(U2852) );
  OAI21_X1 U6450 ( .B1(n5708), .B2(n6597), .A(n7537), .ZN(n7474) );
  NAND2_X1 U6451 ( .A1(n7474), .A2(n7264), .ZN(n5715) );
  INV_X1 U6452 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5710) );
  INV_X1 U6453 ( .A(n7436), .ZN(n7466) );
  AOI22_X1 U6454 ( .A1(EBX_REG_1__SCAN_IN), .A2(n7519), .B1(n7466), .B2(
        REIP_REG_1__SCAN_IN), .ZN(n5709) );
  OAI21_X1 U6455 ( .B1(n7531), .B2(n5710), .A(n5709), .ZN(n5713) );
  OR2_X1 U6456 ( .A1(n6597), .A2(n4884), .ZN(n7452) );
  OAI22_X1 U6457 ( .A1(n5711), .A2(n7452), .B1(n7457), .B2(REIP_REG_1__SCAN_IN), .ZN(n5712) );
  AOI211_X1 U6458 ( .C1(n7521), .C2(n7335), .A(n5713), .B(n5712), .ZN(n5714)
         );
  OAI211_X1 U6459 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n7541), .A(n5715), 
        .B(n5714), .ZN(U2826) );
  AOI21_X1 U6460 ( .B1(n5126), .B2(n5717), .A(n5716), .ZN(n5719) );
  NAND2_X1 U6461 ( .A1(n5114), .A2(n5720), .ZN(n5721) );
  NAND2_X1 U6462 ( .A1(n5722), .A2(n5721), .ZN(n7441) );
  OAI22_X1 U6463 ( .A1(n3659), .A2(n7441), .B1(n7439), .B2(n7259), .ZN(n5723)
         );
  AOI21_X1 U6464 ( .B1(n7449), .B2(n6793), .A(n5723), .ZN(n5724) );
  INV_X1 U6465 ( .A(n5724), .ZN(U2856) );
  NAND2_X1 U6466 ( .A1(n7474), .A2(n7271), .ZN(n5733) );
  INV_X1 U6467 ( .A(REIP_REG_2__SCAN_IN), .ZN(n7434) );
  NAND3_X1 U6468 ( .A1(REIP_REG_1__SCAN_IN), .A2(n7468), .A3(n7434), .ZN(n5727) );
  OAI21_X1 U6469 ( .B1(REIP_REG_1__SCAN_IN), .B2(n7457), .A(n7436), .ZN(n5725)
         );
  NAND2_X1 U6470 ( .A1(REIP_REG_2__SCAN_IN), .A2(n5725), .ZN(n5726) );
  OAI211_X1 U6471 ( .C1(n7531), .C2(n5728), .A(n5727), .B(n5726), .ZN(n5731)
         );
  OAI22_X1 U6472 ( .A1(n5125), .A2(n7452), .B1(n7529), .B2(n5729), .ZN(n5730)
         );
  AOI211_X1 U6473 ( .C1(n7521), .C2(n7347), .A(n5731), .B(n5730), .ZN(n5732)
         );
  OAI211_X1 U6474 ( .C1(n7275), .C2(n7541), .A(n5733), .B(n5732), .ZN(U2825)
         );
  AOI21_X1 U6475 ( .B1(n5956), .B2(n5786), .A(n7608), .ZN(n5742) );
  NOR2_X1 U6476 ( .A1(n5735), .A2(n5734), .ZN(n5741) );
  INV_X1 U6477 ( .A(n5736), .ZN(n5737) );
  NOR3_X1 U6478 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n5737), .ZN(n5775) );
  INV_X1 U6479 ( .A(n5775), .ZN(n5788) );
  AOI211_X1 U6480 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5788), .A(n5739), .B(
        n5738), .ZN(n5740) );
  NAND2_X1 U6481 ( .A1(n5785), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5752) );
  NAND2_X1 U6482 ( .A1(n5744), .A2(n5743), .ZN(n5745) );
  OAI21_X1 U6483 ( .B1(n5747), .B2(n5746), .A(n5745), .ZN(n5791) );
  INV_X1 U6484 ( .A(n5791), .ZN(n5773) );
  OAI22_X1 U6485 ( .A1(n5786), .A2(n5942), .B1(n5773), .B2(n5748), .ZN(n5749)
         );
  AOI21_X1 U6486 ( .B1(n5750), .B2(n5775), .A(n5749), .ZN(n5751) );
  OAI211_X1 U6487 ( .C1(n5956), .C2(n5970), .A(n5752), .B(n5751), .ZN(U3020)
         );
  NAND2_X1 U6488 ( .A1(n5785), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5757) );
  OAI22_X1 U6489 ( .A1(n5786), .A2(n5937), .B1(n5773), .B2(n5753), .ZN(n5754)
         );
  AOI21_X1 U6490 ( .B1(n5775), .B2(n5755), .A(n5754), .ZN(n5756) );
  OAI211_X1 U6491 ( .C1(n5956), .C2(n5988), .A(n5757), .B(n5756), .ZN(U3022)
         );
  NAND2_X1 U6492 ( .A1(n5785), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5763) );
  OAI22_X1 U6493 ( .A1(n5759), .A2(n5788), .B1(n5758), .B2(n5786), .ZN(n5760)
         );
  AOI21_X1 U6494 ( .B1(n5761), .B2(n5791), .A(n5760), .ZN(n5762) );
  OAI211_X1 U6495 ( .C1(n5956), .C2(n6007), .A(n5763), .B(n5762), .ZN(U3024)
         );
  NAND2_X1 U6496 ( .A1(n5785), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5768) );
  OAI22_X1 U6497 ( .A1(n5786), .A2(n5932), .B1(n5773), .B2(n5764), .ZN(n5765)
         );
  AOI21_X1 U6498 ( .B1(n5775), .B2(n5766), .A(n5765), .ZN(n5767) );
  OAI211_X1 U6499 ( .C1(n5956), .C2(n5963), .A(n5768), .B(n5767), .ZN(U3023)
         );
  NAND2_X1 U6500 ( .A1(n5785), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5771) );
  OAI22_X1 U6501 ( .A1(n6413), .A2(n5788), .B1(n6410), .B2(n5786), .ZN(n5769)
         );
  AOI21_X1 U6502 ( .B1(n6416), .B2(n5791), .A(n5769), .ZN(n5770) );
  OAI211_X1 U6503 ( .C1(n5956), .C2(n6419), .A(n5771), .B(n5770), .ZN(U3027)
         );
  NAND2_X1 U6504 ( .A1(n5785), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5778) );
  OAI22_X1 U6505 ( .A1(n5786), .A2(n5949), .B1(n5773), .B2(n5772), .ZN(n5774)
         );
  AOI21_X1 U6506 ( .B1(n5776), .B2(n5775), .A(n5774), .ZN(n5777) );
  OAI211_X1 U6507 ( .C1(n5956), .C2(n5977), .A(n5778), .B(n5777), .ZN(U3021)
         );
  NAND2_X1 U6508 ( .A1(n5785), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5784) );
  OAI22_X1 U6509 ( .A1(n5780), .A2(n5788), .B1(n5779), .B2(n5786), .ZN(n5781)
         );
  AOI21_X1 U6510 ( .B1(n5782), .B2(n5791), .A(n5781), .ZN(n5783) );
  OAI211_X1 U6511 ( .C1(n6000), .C2(n5956), .A(n5784), .B(n5783), .ZN(U3026)
         );
  NAND2_X1 U6512 ( .A1(n5785), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5794) );
  OAI22_X1 U6513 ( .A1(n5789), .A2(n5788), .B1(n5787), .B2(n5786), .ZN(n5790)
         );
  AOI21_X1 U6514 ( .B1(n5792), .B2(n5791), .A(n5790), .ZN(n5793) );
  OAI211_X1 U6515 ( .C1(n5993), .C2(n5956), .A(n5794), .B(n5793), .ZN(U3025)
         );
  OAI21_X1 U6517 ( .B1(n6506), .B2(n7457), .A(n7436), .ZN(n5859) );
  INV_X1 U6518 ( .A(n5859), .ZN(n5835) );
  NAND3_X1 U6519 ( .A1(n7468), .A2(n7469), .A3(REIP_REG_5__SCAN_IN), .ZN(n7493) );
  OAI33_X1 U6520 ( .A1(1'b0), .A2(n5835), .A3(n7181), .B1(REIP_REG_8__SCAN_IN), 
        .B2(n7491), .B3(n7493), .ZN(n5796) );
  INV_X1 U6521 ( .A(n5796), .ZN(n5802) );
  INV_X1 U6522 ( .A(n6426), .ZN(n5800) );
  AOI22_X1 U6523 ( .A1(n7519), .A2(EBX_REG_8__SCAN_IN), .B1(n7521), .B2(n7361), 
        .ZN(n5797) );
  NAND2_X1 U6524 ( .A1(n7436), .A2(n7305), .ZN(n7514) );
  OAI211_X1 U6525 ( .C1(n7531), .C2(n5798), .A(n5797), .B(n7514), .ZN(n5799)
         );
  AOI21_X1 U6526 ( .B1(n7504), .B2(n5800), .A(n5799), .ZN(n5801) );
  OAI211_X1 U6527 ( .C1(n6430), .C2(n7537), .A(n5802), .B(n5801), .ZN(U2819)
         );
  NOR2_X1 U6528 ( .A1(n5803), .A2(n7586), .ZN(n7602) );
  NOR2_X1 U6529 ( .A1(n7129), .A2(n3937), .ZN(n5807) );
  NOR2_X1 U6530 ( .A1(n5805), .A2(n5804), .ZN(n5806) );
  AOI211_X1 U6531 ( .C1(n7602), .C2(n7129), .A(n5807), .B(n5806), .ZN(n5808)
         );
  OAI21_X1 U6532 ( .B1(n7425), .B2(n5809), .A(n5808), .ZN(U3465) );
  AND2_X1 U6533 ( .A1(n5146), .A2(n5810), .ZN(n5811) );
  OR2_X1 U6534 ( .A1(n5811), .A2(n5833), .ZN(n6471) );
  NOR2_X1 U6535 ( .A1(n5813), .A2(n5812), .ZN(n5814) );
  OR2_X1 U6536 ( .A1(n5839), .A2(n5814), .ZN(n6476) );
  OAI22_X1 U6537 ( .A1(n3659), .A2(n6476), .B1(n5815), .B2(n7259), .ZN(n5816)
         );
  INV_X1 U6538 ( .A(n5816), .ZN(n5817) );
  OAI21_X1 U6539 ( .B1(n6471), .B2(n7256), .A(n5817), .ZN(U2850) );
  INV_X1 U6540 ( .A(n7345), .ZN(n5818) );
  INV_X1 U6541 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n7102) );
  NAND2_X1 U6542 ( .A1(n6472), .A2(n7102), .ZN(n5823) );
  INV_X1 U6543 ( .A(n7062), .ZN(n7063) );
  AOI21_X1 U6544 ( .B1(n7063), .B2(n5820), .A(n5819), .ZN(n7357) );
  OAI21_X1 U6545 ( .B1(n7079), .B2(n7345), .A(n7357), .ZN(n6025) );
  INV_X1 U6546 ( .A(REIP_REG_3__SCAN_IN), .ZN(n7174) );
  OAI22_X1 U6547 ( .A1(n7090), .A2(n7441), .B1(n7174), .B2(n7088), .ZN(n5821)
         );
  AOI21_X1 U6548 ( .B1(n6025), .B2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n5821), 
        .ZN(n5822) );
  OAI211_X1 U6549 ( .C1(n5824), .C2(n7350), .A(n5823), .B(n5822), .ZN(U3015)
         );
  NAND2_X1 U6550 ( .A1(n7468), .A2(n6506), .ZN(n5836) );
  OAI22_X1 U6551 ( .A1(n5836), .A2(REIP_REG_9__SCAN_IN), .B1(n7535), .B2(n6476), .ZN(n5828) );
  AOI22_X1 U6552 ( .A1(EBX_REG_9__SCAN_IN), .A2(n7519), .B1(
        REIP_REG_9__SCAN_IN), .B2(n5859), .ZN(n5825) );
  OAI211_X1 U6553 ( .C1(n7531), .C2(n5826), .A(n5825), .B(n7514), .ZN(n5827)
         );
  AOI211_X1 U6554 ( .C1(n6468), .C2(n7504), .A(n5828), .B(n5827), .ZN(n5829)
         );
  OAI21_X1 U6555 ( .B1(n7537), .B2(n6471), .A(n5829), .ZN(U2818) );
  INV_X1 U6556 ( .A(DATAI_9_), .ZN(n5830) );
  INV_X1 U6557 ( .A(EAX_REG_9__SCAN_IN), .ZN(n7672) );
  OAI222_X1 U6558 ( .A1(n6833), .A2(n5830), .B1(n6829), .B2(n7672), .C1(n6831), 
        .C2(n6471), .ZN(U2882) );
  NOR2_X1 U6559 ( .A1(n5833), .A2(n5832), .ZN(n5834) );
  OR2_X1 U6560 ( .A1(n5831), .A2(n5834), .ZN(n6975) );
  INV_X1 U6561 ( .A(REIP_REG_9__SCAN_IN), .ZN(n7184) );
  NOR2_X1 U6562 ( .A1(n7184), .A2(n5836), .ZN(n6449) );
  OAI211_X1 U6563 ( .C1(REIP_REG_9__SCAN_IN), .C2(n5836), .A(
        REIP_REG_10__SCAN_IN), .B(n5835), .ZN(n5862) );
  OAI21_X1 U6564 ( .B1(REIP_REG_10__SCAN_IN), .B2(n6449), .A(n5862), .ZN(n5846) );
  INV_X1 U6565 ( .A(n6971), .ZN(n5844) );
  INV_X1 U6566 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5842) );
  OR2_X1 U6567 ( .A1(n5839), .A2(n5838), .ZN(n5840) );
  NAND2_X1 U6568 ( .A1(n5837), .A2(n5840), .ZN(n5849) );
  INV_X1 U6569 ( .A(n5849), .ZN(n7375) );
  AOI22_X1 U6570 ( .A1(n7521), .A2(n7375), .B1(n7519), .B2(EBX_REG_10__SCAN_IN), .ZN(n5841) );
  OAI211_X1 U6571 ( .C1(n7531), .C2(n5842), .A(n5841), .B(n7514), .ZN(n5843)
         );
  AOI21_X1 U6572 ( .B1(n7504), .B2(n5844), .A(n5843), .ZN(n5845) );
  OAI211_X1 U6573 ( .C1(n6975), .C2(n7537), .A(n5846), .B(n5845), .ZN(U2817)
         );
  INV_X1 U6574 ( .A(DATAI_10_), .ZN(n5847) );
  INV_X1 U6575 ( .A(EAX_REG_10__SCAN_IN), .ZN(n7676) );
  OAI222_X1 U6576 ( .A1(n6975), .A2(n6831), .B1(n6833), .B2(n5847), .C1(n6829), 
        .C2(n7676), .ZN(U2881) );
  INV_X1 U6577 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5848) );
  OAI222_X1 U6578 ( .A1(n5849), .A2(n3659), .B1(n5848), .B2(n7259), .C1(n6975), 
        .C2(n7256), .ZN(U2849) );
  OAI21_X1 U6579 ( .B1(n5831), .B2(n5852), .A(n5851), .ZN(n6967) );
  XNOR2_X1 U6580 ( .A(n5837), .B(n6451), .ZN(n5856) );
  OAI22_X1 U6581 ( .A1(n3659), .A2(n5856), .B1(n5853), .B2(n7259), .ZN(n5854)
         );
  INV_X1 U6582 ( .A(n5854), .ZN(n5855) );
  OAI21_X1 U6583 ( .B1(n6967), .B2(n7256), .A(n5855), .ZN(U2848) );
  INV_X1 U6584 ( .A(n5856), .ZN(n7395) );
  AOI22_X1 U6585 ( .A1(n7519), .A2(EBX_REG_11__SCAN_IN), .B1(n7521), .B2(n7395), .ZN(n5857) );
  OAI211_X1 U6586 ( .C1(n7531), .C2(n5858), .A(n5857), .B(n7514), .ZN(n5864)
         );
  INV_X1 U6587 ( .A(REIP_REG_11__SCAN_IN), .ZN(n7188) );
  AOI21_X1 U6588 ( .B1(n5861), .B2(n5860), .A(n5859), .ZN(n6495) );
  AOI21_X1 U6589 ( .B1(n7188), .B2(n5862), .A(n6495), .ZN(n5863) );
  AOI211_X1 U6590 ( .C1(n6964), .C2(n7504), .A(n5864), .B(n5863), .ZN(n5865)
         );
  OAI21_X1 U6591 ( .B1(n7537), .B2(n6967), .A(n5865), .ZN(U2816) );
  INV_X1 U6592 ( .A(n5874), .ZN(n5877) );
  NOR2_X1 U6593 ( .A1(n3937), .A2(n5877), .ZN(n6013) );
  INV_X1 U6594 ( .A(n6013), .ZN(n5890) );
  AOI21_X1 U6595 ( .B1(n5867), .B2(n5866), .A(n6013), .ZN(n5878) );
  INV_X1 U6596 ( .A(n5868), .ZN(n5871) );
  OAI21_X1 U6597 ( .B1(n5871), .B2(n5870), .A(n5869), .ZN(n5876) );
  NAND2_X1 U6598 ( .A1(n5878), .A2(n5876), .ZN(n5872) );
  OAI211_X1 U6599 ( .C1(n5875), .C2(n5874), .A(n5873), .B(n5872), .ZN(n6012)
         );
  INV_X1 U6600 ( .A(n5876), .ZN(n5879) );
  OAI22_X1 U6601 ( .A1(n5879), .A2(n5878), .B1(n5877), .B2(n7584), .ZN(n5990)
         );
  AOI22_X1 U6602 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n6012), .B1(n5971), 
        .B2(n5990), .ZN(n5880) );
  OAI21_X1 U6603 ( .B1(n5973), .B2(n5890), .A(n5880), .ZN(n5881) );
  AOI21_X1 U6604 ( .B1(n6019), .B2(n5975), .A(n5881), .ZN(n5882) );
  OAI21_X1 U6605 ( .B1(n5977), .B2(n6016), .A(n5882), .ZN(U3093) );
  AOI22_X1 U6606 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n6012), .B1(n5979), 
        .B2(n5990), .ZN(n5883) );
  OAI21_X1 U6607 ( .B1(n5983), .B2(n5890), .A(n5883), .ZN(n5884) );
  AOI21_X1 U6608 ( .B1(n6019), .B2(n5985), .A(n5884), .ZN(n5885) );
  OAI21_X1 U6609 ( .B1(n5988), .B2(n6016), .A(n5885), .ZN(U3094) );
  AOI22_X1 U6610 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n6012), .B1(n5957), 
        .B2(n5990), .ZN(n5886) );
  OAI21_X1 U6611 ( .B1(n5959), .B2(n5890), .A(n5886), .ZN(n5887) );
  AOI21_X1 U6612 ( .B1(n6019), .B2(n5961), .A(n5887), .ZN(n5888) );
  OAI21_X1 U6613 ( .B1(n5963), .B2(n6016), .A(n5888), .ZN(U3095) );
  AOI22_X1 U6614 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n6012), .B1(n5964), 
        .B2(n5990), .ZN(n5889) );
  OAI21_X1 U6615 ( .B1(n5966), .B2(n5890), .A(n5889), .ZN(n5891) );
  AOI21_X1 U6616 ( .B1(n6019), .B2(n5968), .A(n5891), .ZN(n5892) );
  OAI21_X1 U6617 ( .B1(n5970), .B2(n6016), .A(n5892), .ZN(U3092) );
  INV_X1 U6618 ( .A(n5893), .ZN(n5922) );
  AOI22_X1 U6619 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n5916), .B1(n5957), 
        .B2(n5915), .ZN(n5895) );
  OAI21_X1 U6620 ( .B1(n5918), .B2(n5932), .A(n5895), .ZN(n5896) );
  AOI21_X1 U6621 ( .B1(n5920), .B2(n5934), .A(n5896), .ZN(n5897) );
  OAI21_X1 U6622 ( .B1(n5922), .B2(n5959), .A(n5897), .ZN(U3127) );
  INV_X1 U6623 ( .A(n5898), .ZN(n5930) );
  INV_X1 U6624 ( .A(n5899), .ZN(n5928) );
  AOI22_X1 U6625 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n5924), .B1(n5957), 
        .B2(n5923), .ZN(n5900) );
  OAI21_X1 U6626 ( .B1(n5926), .B2(n5932), .A(n5900), .ZN(n5901) );
  AOI21_X1 U6627 ( .B1(n5928), .B2(n5934), .A(n5901), .ZN(n5902) );
  OAI21_X1 U6628 ( .B1(n5930), .B2(n5959), .A(n5902), .ZN(U3063) );
  AOI22_X1 U6629 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n5916), .B1(n5971), 
        .B2(n5915), .ZN(n5903) );
  OAI21_X1 U6630 ( .B1(n5918), .B2(n5949), .A(n5903), .ZN(n5904) );
  AOI21_X1 U6631 ( .B1(n5920), .B2(n5952), .A(n5904), .ZN(n5905) );
  OAI21_X1 U6632 ( .B1(n5922), .B2(n5973), .A(n5905), .ZN(U3125) );
  AOI22_X1 U6633 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n5924), .B1(n5979), 
        .B2(n5923), .ZN(n5906) );
  OAI21_X1 U6634 ( .B1(n5926), .B2(n5937), .A(n5906), .ZN(n5907) );
  AOI21_X1 U6635 ( .B1(n5928), .B2(n5939), .A(n5907), .ZN(n5908) );
  OAI21_X1 U6636 ( .B1(n5930), .B2(n5983), .A(n5908), .ZN(U3062) );
  AOI22_X1 U6637 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n5916), .B1(n5979), 
        .B2(n5915), .ZN(n5909) );
  OAI21_X1 U6638 ( .B1(n5918), .B2(n5937), .A(n5909), .ZN(n5910) );
  AOI21_X1 U6639 ( .B1(n5920), .B2(n5939), .A(n5910), .ZN(n5911) );
  OAI21_X1 U6640 ( .B1(n5922), .B2(n5983), .A(n5911), .ZN(U3126) );
  AOI22_X1 U6641 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n5924), .B1(n5971), 
        .B2(n5923), .ZN(n5912) );
  OAI21_X1 U6642 ( .B1(n5926), .B2(n5949), .A(n5912), .ZN(n5913) );
  AOI21_X1 U6643 ( .B1(n5928), .B2(n5952), .A(n5913), .ZN(n5914) );
  OAI21_X1 U6644 ( .B1(n5930), .B2(n5973), .A(n5914), .ZN(U3061) );
  AOI22_X1 U6645 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n5916), .B1(n5964), 
        .B2(n5915), .ZN(n5917) );
  OAI21_X1 U6646 ( .B1(n5918), .B2(n5942), .A(n5917), .ZN(n5919) );
  AOI21_X1 U6647 ( .B1(n5920), .B2(n5944), .A(n5919), .ZN(n5921) );
  OAI21_X1 U6648 ( .B1(n5966), .B2(n5922), .A(n5921), .ZN(U3124) );
  AOI22_X1 U6649 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n5924), .B1(n5964), 
        .B2(n5923), .ZN(n5925) );
  OAI21_X1 U6650 ( .B1(n5926), .B2(n5942), .A(n5925), .ZN(n5927) );
  AOI21_X1 U6651 ( .B1(n5928), .B2(n5944), .A(n5927), .ZN(n5929) );
  OAI21_X1 U6652 ( .B1(n5966), .B2(n5930), .A(n5929), .ZN(U3060) );
  INV_X1 U6653 ( .A(n6411), .ZN(n5953) );
  AOI22_X1 U6654 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n5947), .B1(n5957), 
        .B2(n5946), .ZN(n5931) );
  OAI21_X1 U6655 ( .B1(n5950), .B2(n5932), .A(n5931), .ZN(n5933) );
  AOI21_X1 U6656 ( .B1(n5953), .B2(n5934), .A(n5933), .ZN(n5935) );
  OAI21_X1 U6657 ( .B1(n5955), .B2(n5959), .A(n5935), .ZN(U3079) );
  AOI22_X1 U6658 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n5947), .B1(n5979), 
        .B2(n5946), .ZN(n5936) );
  OAI21_X1 U6659 ( .B1(n5950), .B2(n5937), .A(n5936), .ZN(n5938) );
  AOI21_X1 U6660 ( .B1(n5953), .B2(n5939), .A(n5938), .ZN(n5940) );
  OAI21_X1 U6661 ( .B1(n5955), .B2(n5983), .A(n5940), .ZN(U3078) );
  AOI22_X1 U6662 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n5947), .B1(n5964), 
        .B2(n5946), .ZN(n5941) );
  OAI21_X1 U6663 ( .B1(n5950), .B2(n5942), .A(n5941), .ZN(n5943) );
  AOI21_X1 U6664 ( .B1(n5953), .B2(n5944), .A(n5943), .ZN(n5945) );
  OAI21_X1 U6665 ( .B1(n5966), .B2(n5955), .A(n5945), .ZN(U3076) );
  AOI22_X1 U6666 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n5947), .B1(n5971), 
        .B2(n5946), .ZN(n5948) );
  OAI21_X1 U6667 ( .B1(n5950), .B2(n5949), .A(n5948), .ZN(n5951) );
  AOI21_X1 U6668 ( .B1(n5953), .B2(n5952), .A(n5951), .ZN(n5954) );
  OAI21_X1 U6669 ( .B1(n5955), .B2(n5973), .A(n5954), .ZN(U3077) );
  INV_X1 U6670 ( .A(n5956), .ZN(n5986) );
  AOI22_X1 U6671 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n5980), .B1(n5957), 
        .B2(n5978), .ZN(n5958) );
  OAI21_X1 U6672 ( .B1(n5959), .B2(n5982), .A(n5958), .ZN(n5960) );
  AOI21_X1 U6673 ( .B1(n5986), .B2(n5961), .A(n5960), .ZN(n5962) );
  OAI21_X1 U6674 ( .B1(n5989), .B2(n5963), .A(n5962), .ZN(U3031) );
  AOI22_X1 U6675 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n5980), .B1(n5964), 
        .B2(n5978), .ZN(n5965) );
  OAI21_X1 U6676 ( .B1(n5966), .B2(n5982), .A(n5965), .ZN(n5967) );
  AOI21_X1 U6677 ( .B1(n5986), .B2(n5968), .A(n5967), .ZN(n5969) );
  OAI21_X1 U6678 ( .B1(n5989), .B2(n5970), .A(n5969), .ZN(U3028) );
  AOI22_X1 U6679 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n5980), .B1(n5971), 
        .B2(n5978), .ZN(n5972) );
  OAI21_X1 U6680 ( .B1(n5973), .B2(n5982), .A(n5972), .ZN(n5974) );
  AOI21_X1 U6681 ( .B1(n5986), .B2(n5975), .A(n5974), .ZN(n5976) );
  OAI21_X1 U6682 ( .B1(n5989), .B2(n5977), .A(n5976), .ZN(U3029) );
  AOI22_X1 U6683 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n5980), .B1(n5979), 
        .B2(n5978), .ZN(n5981) );
  OAI21_X1 U6684 ( .B1(n5983), .B2(n5982), .A(n5981), .ZN(n5984) );
  AOI21_X1 U6685 ( .B1(n5986), .B2(n5985), .A(n5984), .ZN(n5987) );
  OAI21_X1 U6686 ( .B1(n5989), .B2(n5988), .A(n5987), .ZN(U3030) );
  INV_X1 U6687 ( .A(n5990), .ZN(n6022) );
  AOI22_X1 U6688 ( .A1(n5991), .A2(n6013), .B1(INSTQUEUE_REG_9__5__SCAN_IN), 
        .B2(n6012), .ZN(n5992) );
  OAI21_X1 U6689 ( .B1(n5993), .B2(n6016), .A(n5992), .ZN(n5994) );
  AOI21_X1 U6690 ( .B1(n6019), .B2(n5995), .A(n5994), .ZN(n5996) );
  OAI21_X1 U6691 ( .B1(n6022), .B2(n5997), .A(n5996), .ZN(U3097) );
  AOI22_X1 U6692 ( .A1(n5998), .A2(n6013), .B1(INSTQUEUE_REG_9__6__SCAN_IN), 
        .B2(n6012), .ZN(n5999) );
  OAI21_X1 U6693 ( .B1(n6000), .B2(n6016), .A(n5999), .ZN(n6001) );
  AOI21_X1 U6694 ( .B1(n6019), .B2(n6002), .A(n6001), .ZN(n6003) );
  OAI21_X1 U6695 ( .B1(n6022), .B2(n6004), .A(n6003), .ZN(U3098) );
  AOI22_X1 U6696 ( .A1(n6005), .A2(n6013), .B1(INSTQUEUE_REG_9__4__SCAN_IN), 
        .B2(n6012), .ZN(n6006) );
  OAI21_X1 U6697 ( .B1(n6007), .B2(n6016), .A(n6006), .ZN(n6008) );
  AOI21_X1 U6698 ( .B1(n6019), .B2(n6009), .A(n6008), .ZN(n6010) );
  OAI21_X1 U6699 ( .B1(n6022), .B2(n6011), .A(n6010), .ZN(U3096) );
  AOI22_X1 U6700 ( .A1(n6014), .A2(n6013), .B1(INSTQUEUE_REG_9__7__SCAN_IN), 
        .B2(n6012), .ZN(n6015) );
  OAI21_X1 U6701 ( .B1(n6419), .B2(n6016), .A(n6015), .ZN(n6017) );
  AOI21_X1 U6702 ( .B1(n6019), .B2(n6018), .A(n6017), .ZN(n6020) );
  OAI21_X1 U6703 ( .B1(n6022), .B2(n6021), .A(n6020), .ZN(U3099) );
  XNOR2_X1 U6704 ( .A(n6024), .B(n6023), .ZN(n7276) );
  NAND2_X1 U6705 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6026) );
  NOR2_X1 U6706 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6026), .ZN(n6439)
         );
  NAND2_X1 U6707 ( .A1(n7370), .A2(REIP_REG_5__SCAN_IN), .ZN(n7280) );
  OAI21_X1 U6708 ( .B1(n7090), .B2(n7471), .A(n7280), .ZN(n6028) );
  AOI21_X1 U6709 ( .B1(n6472), .B2(n6026), .A(n6025), .ZN(n7100) );
  NOR2_X1 U6710 ( .A1(n7100), .A2(n6438), .ZN(n6027) );
  AOI211_X1 U6711 ( .C1(n6472), .C2(n6439), .A(n6028), .B(n6027), .ZN(n6029)
         );
  OAI21_X1 U6712 ( .B1(n7350), .B2(n7276), .A(n6029), .ZN(U3013) );
  XOR2_X1 U6713 ( .A(DATAI_30_), .B(keyinput_1), .Z(n6032) );
  XOR2_X1 U6714 ( .A(DATAI_31_), .B(keyinput_0), .Z(n6031) );
  XNOR2_X1 U6715 ( .A(DATAI_28_), .B(keyinput_3), .ZN(n6030) );
  AOI21_X1 U6716 ( .B1(n6032), .B2(n6031), .A(n6030), .ZN(n6035) );
  XOR2_X1 U6717 ( .A(DATAI_27_), .B(keyinput_4), .Z(n6034) );
  XOR2_X1 U6718 ( .A(DATAI_29_), .B(keyinput_2), .Z(n6033) );
  NAND3_X1 U6719 ( .A1(n6035), .A2(n6034), .A3(n6033), .ZN(n6038) );
  XOR2_X1 U6720 ( .A(DATAI_26_), .B(keyinput_5), .Z(n6037) );
  XNOR2_X1 U6721 ( .A(DATAI_25_), .B(keyinput_6), .ZN(n6036) );
  AOI21_X1 U6722 ( .B1(n6038), .B2(n6037), .A(n6036), .ZN(n6041) );
  XOR2_X1 U6723 ( .A(DATAI_24_), .B(keyinput_7), .Z(n6040) );
  XNOR2_X1 U6724 ( .A(DATAI_23_), .B(keyinput_8), .ZN(n6039) );
  NOR3_X1 U6725 ( .A1(n6041), .A2(n6040), .A3(n6039), .ZN(n6044) );
  XOR2_X1 U6726 ( .A(DATAI_22_), .B(keyinput_9), .Z(n6043) );
  XOR2_X1 U6727 ( .A(DATAI_21_), .B(keyinput_10), .Z(n6042) );
  NOR3_X1 U6728 ( .A1(n6044), .A2(n6043), .A3(n6042), .ZN(n6047) );
  XNOR2_X1 U6729 ( .A(DATAI_20_), .B(keyinput_11), .ZN(n6046) );
  XNOR2_X1 U6730 ( .A(DATAI_19_), .B(keyinput_12), .ZN(n6045) );
  NOR3_X1 U6731 ( .A1(n6047), .A2(n6046), .A3(n6045), .ZN(n6050) );
  XNOR2_X1 U6732 ( .A(DATAI_18_), .B(keyinput_13), .ZN(n6049) );
  XOR2_X1 U6733 ( .A(DATAI_17_), .B(keyinput_14), .Z(n6048) );
  OAI21_X1 U6734 ( .B1(n6050), .B2(n6049), .A(n6048), .ZN(n6053) );
  XOR2_X1 U6735 ( .A(DATAI_16_), .B(keyinput_15), .Z(n6052) );
  XOR2_X1 U6736 ( .A(DATAI_15_), .B(keyinput_16), .Z(n6051) );
  AOI21_X1 U6737 ( .B1(n6053), .B2(n6052), .A(n6051), .ZN(n6056) );
  XOR2_X1 U6738 ( .A(DATAI_14_), .B(keyinput_17), .Z(n6055) );
  XOR2_X1 U6739 ( .A(DATAI_13_), .B(keyinput_18), .Z(n6054) );
  OAI21_X1 U6740 ( .B1(n6056), .B2(n6055), .A(n6054), .ZN(n6064) );
  XOR2_X1 U6741 ( .A(DATAI_12_), .B(keyinput_19), .Z(n6063) );
  INV_X1 U6742 ( .A(keyinput_21), .ZN(n6057) );
  XNOR2_X1 U6743 ( .A(n6057), .B(DATAI_10_), .ZN(n6061) );
  XNOR2_X1 U6744 ( .A(DATAI_9_), .B(keyinput_22), .ZN(n6060) );
  XNOR2_X1 U6745 ( .A(DATAI_8_), .B(keyinput_23), .ZN(n6059) );
  XNOR2_X1 U6746 ( .A(DATAI_11_), .B(keyinput_20), .ZN(n6058) );
  NAND4_X1 U6747 ( .A1(n6061), .A2(n6060), .A3(n6059), .A4(n6058), .ZN(n6062)
         );
  AOI21_X1 U6748 ( .B1(n6064), .B2(n6063), .A(n6062), .ZN(n6075) );
  XNOR2_X1 U6749 ( .A(DATAI_6_), .B(keyinput_25), .ZN(n6068) );
  XNOR2_X1 U6750 ( .A(DATAI_7_), .B(keyinput_24), .ZN(n6067) );
  XNOR2_X1 U6751 ( .A(DATAI_4_), .B(keyinput_27), .ZN(n6066) );
  XNOR2_X1 U6752 ( .A(DATAI_5_), .B(keyinput_26), .ZN(n6065) );
  NAND4_X1 U6753 ( .A1(n6068), .A2(n6067), .A3(n6066), .A4(n6065), .ZN(n6074)
         );
  XOR2_X1 U6754 ( .A(DATAI_1_), .B(keyinput_30), .Z(n6072) );
  XOR2_X1 U6755 ( .A(DATAI_3_), .B(keyinput_28), .Z(n6071) );
  XOR2_X1 U6756 ( .A(DATAI_2_), .B(keyinput_29), .Z(n6070) );
  XNOR2_X1 U6757 ( .A(n5141), .B(keyinput_31), .ZN(n6069) );
  NAND4_X1 U6758 ( .A1(n6072), .A2(n6071), .A3(n6070), .A4(n6069), .ZN(n6073)
         );
  NOR3_X1 U6759 ( .A1(n6075), .A2(n6074), .A3(n6073), .ZN(n6077) );
  XNOR2_X1 U6760 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(keyinput_32), .ZN(n6076) );
  NOR2_X1 U6761 ( .A1(n6077), .A2(n6076), .ZN(n6081) );
  INV_X1 U6762 ( .A(BS16_N), .ZN(n7108) );
  XNOR2_X1 U6763 ( .A(n7108), .B(keyinput_34), .ZN(n6080) );
  XNOR2_X1 U6764 ( .A(n7634), .B(keyinput_35), .ZN(n6079) );
  XNOR2_X1 U6765 ( .A(NA_N), .B(keyinput_33), .ZN(n6078) );
  NOR4_X1 U6766 ( .A1(n6081), .A2(n6080), .A3(n6079), .A4(n6078), .ZN(n6087)
         );
  INV_X1 U6767 ( .A(HOLD), .ZN(n7310) );
  XNOR2_X1 U6768 ( .A(n7310), .B(keyinput_36), .ZN(n6086) );
  XOR2_X1 U6769 ( .A(READREQUEST_REG_SCAN_IN), .B(keyinput_37), .Z(n6084) );
  XOR2_X1 U6770 ( .A(CODEFETCH_REG_SCAN_IN), .B(keyinput_39), .Z(n6083) );
  XNOR2_X1 U6771 ( .A(ADS_N_REG_SCAN_IN), .B(keyinput_38), .ZN(n6082) );
  NOR3_X1 U6772 ( .A1(n6084), .A2(n6083), .A3(n6082), .ZN(n6085) );
  OAI21_X1 U6773 ( .B1(n6087), .B2(n6086), .A(n6085), .ZN(n6090) );
  INV_X1 U6774 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n7628) );
  XNOR2_X1 U6775 ( .A(n7628), .B(keyinput_40), .ZN(n6089) );
  XNOR2_X1 U6776 ( .A(D_C_N_REG_SCAN_IN), .B(keyinput_41), .ZN(n6088) );
  AOI21_X1 U6777 ( .B1(n6090), .B2(n6089), .A(n6088), .ZN(n6093) );
  XNOR2_X1 U6778 ( .A(n7608), .B(keyinput_43), .ZN(n6092) );
  XNOR2_X1 U6779 ( .A(REQUESTPENDING_REG_SCAN_IN), .B(keyinput_42), .ZN(n6091)
         );
  NOR3_X1 U6780 ( .A1(n6093), .A2(n6092), .A3(n6091), .ZN(n6096) );
  XOR2_X1 U6781 ( .A(MORE_REG_SCAN_IN), .B(keyinput_44), .Z(n6095) );
  XOR2_X1 U6782 ( .A(FLUSH_REG_SCAN_IN), .B(keyinput_45), .Z(n6094) );
  NOR3_X1 U6783 ( .A1(n6096), .A2(n6095), .A3(n6094), .ZN(n6102) );
  INV_X1 U6784 ( .A(W_R_N_REG_SCAN_IN), .ZN(n7308) );
  XNOR2_X1 U6785 ( .A(n7308), .B(keyinput_46), .ZN(n6101) );
  XOR2_X1 U6786 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(keyinput_49), .Z(n6100) );
  OAI22_X1 U6787 ( .A1(BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_48), .B1(
        BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_47), .ZN(n6098) );
  AND2_X1 U6788 ( .A1(BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_48), .ZN(n6097)
         );
  AOI211_X1 U6789 ( .C1(BYTEENABLE_REG_0__SCAN_IN), .C2(keyinput_47), .A(n6098), .B(n6097), .ZN(n6099) );
  OAI211_X1 U6790 ( .C1(n6102), .C2(n6101), .A(n6100), .B(n6099), .ZN(n6106)
         );
  INV_X1 U6791 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n7232) );
  XNOR2_X1 U6792 ( .A(n7232), .B(keyinput_50), .ZN(n6105) );
  XOR2_X1 U6793 ( .A(REIP_REG_31__SCAN_IN), .B(keyinput_51), .Z(n6104) );
  XOR2_X1 U6794 ( .A(REIP_REG_30__SCAN_IN), .B(keyinput_52), .Z(n6103) );
  AOI211_X1 U6795 ( .C1(n6106), .C2(n6105), .A(n6104), .B(n6103), .ZN(n6114)
         );
  XNOR2_X1 U6796 ( .A(REIP_REG_28__SCAN_IN), .B(keyinput_54), .ZN(n6113) );
  XNOR2_X1 U6797 ( .A(REIP_REG_26__SCAN_IN), .B(keyinput_56), .ZN(n6112) );
  XOR2_X1 U6798 ( .A(REIP_REG_25__SCAN_IN), .B(keyinput_57), .Z(n6110) );
  XNOR2_X1 U6799 ( .A(REIP_REG_29__SCAN_IN), .B(keyinput_53), .ZN(n6109) );
  XNOR2_X1 U6800 ( .A(REIP_REG_24__SCAN_IN), .B(keyinput_58), .ZN(n6108) );
  XNOR2_X1 U6801 ( .A(REIP_REG_27__SCAN_IN), .B(keyinput_55), .ZN(n6107) );
  NAND4_X1 U6802 ( .A1(n6110), .A2(n6109), .A3(n6108), .A4(n6107), .ZN(n6111)
         );
  NOR4_X1 U6803 ( .A1(n6114), .A2(n6113), .A3(n6112), .A4(n6111), .ZN(n6118)
         );
  XNOR2_X1 U6804 ( .A(REIP_REG_23__SCAN_IN), .B(keyinput_59), .ZN(n6117) );
  XOR2_X1 U6805 ( .A(REIP_REG_22__SCAN_IN), .B(keyinput_60), .Z(n6116) );
  XNOR2_X1 U6806 ( .A(REIP_REG_21__SCAN_IN), .B(keyinput_61), .ZN(n6115) );
  OAI211_X1 U6807 ( .C1(n6118), .C2(n6117), .A(n6116), .B(n6115), .ZN(n6121)
         );
  XOR2_X1 U6808 ( .A(REIP_REG_19__SCAN_IN), .B(keyinput_63), .Z(n6120) );
  XNOR2_X1 U6809 ( .A(REIP_REG_20__SCAN_IN), .B(keyinput_62), .ZN(n6119) );
  NAND3_X1 U6810 ( .A1(n6121), .A2(n6120), .A3(n6119), .ZN(n6128) );
  XOR2_X1 U6811 ( .A(REIP_REG_16__SCAN_IN), .B(keyinput_66), .Z(n6124) );
  XNOR2_X1 U6812 ( .A(n7199), .B(keyinput_65), .ZN(n6123) );
  XNOR2_X1 U6813 ( .A(REIP_REG_18__SCAN_IN), .B(keyinput_64), .ZN(n6122) );
  NOR3_X1 U6814 ( .A1(n6124), .A2(n6123), .A3(n6122), .ZN(n6127) );
  INV_X1 U6815 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n7231) );
  XNOR2_X1 U6816 ( .A(n7231), .B(keyinput_67), .ZN(n6126) );
  XNOR2_X1 U6817 ( .A(BE_N_REG_2__SCAN_IN), .B(keyinput_68), .ZN(n6125) );
  AOI211_X1 U6818 ( .C1(n6128), .C2(n6127), .A(n6126), .B(n6125), .ZN(n6132)
         );
  INV_X1 U6819 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n7248) );
  XNOR2_X1 U6820 ( .A(n7248), .B(keyinput_69), .ZN(n6131) );
  XOR2_X1 U6821 ( .A(BE_N_REG_0__SCAN_IN), .B(keyinput_70), .Z(n6130) );
  INV_X1 U6822 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n7228) );
  XNOR2_X1 U6823 ( .A(n7228), .B(keyinput_71), .ZN(n6129) );
  OAI211_X1 U6824 ( .C1(n6132), .C2(n6131), .A(n6130), .B(n6129), .ZN(n6135)
         );
  INV_X1 U6825 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n7225) );
  XNOR2_X1 U6826 ( .A(n7225), .B(keyinput_72), .ZN(n6134) );
  XNOR2_X1 U6827 ( .A(ADDRESS_REG_27__SCAN_IN), .B(keyinput_73), .ZN(n6133) );
  AOI21_X1 U6828 ( .B1(n6135), .B2(n6134), .A(n6133), .ZN(n6138) );
  INV_X1 U6829 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n7220) );
  XNOR2_X1 U6830 ( .A(n7220), .B(keyinput_74), .ZN(n6137) );
  XNOR2_X1 U6831 ( .A(ADDRESS_REG_25__SCAN_IN), .B(keyinput_75), .ZN(n6136) );
  OAI21_X1 U6832 ( .B1(n6138), .B2(n6137), .A(n6136), .ZN(n6142) );
  XNOR2_X1 U6833 ( .A(ADDRESS_REG_24__SCAN_IN), .B(keyinput_76), .ZN(n6141) );
  XNOR2_X1 U6834 ( .A(ADDRESS_REG_23__SCAN_IN), .B(keyinput_77), .ZN(n6140) );
  XNOR2_X1 U6835 ( .A(ADDRESS_REG_22__SCAN_IN), .B(keyinput_78), .ZN(n6139) );
  AOI211_X1 U6836 ( .C1(n6142), .C2(n6141), .A(n6140), .B(n6139), .ZN(n6145)
         );
  XNOR2_X1 U6837 ( .A(ADDRESS_REG_21__SCAN_IN), .B(keyinput_79), .ZN(n6144) );
  XNOR2_X1 U6838 ( .A(ADDRESS_REG_20__SCAN_IN), .B(keyinput_80), .ZN(n6143) );
  NOR3_X1 U6839 ( .A1(n6145), .A2(n6144), .A3(n6143), .ZN(n6158) );
  XOR2_X1 U6840 ( .A(ADDRESS_REG_16__SCAN_IN), .B(keyinput_84), .Z(n6155) );
  INV_X1 U6841 ( .A(keyinput_87), .ZN(n6146) );
  NAND2_X1 U6842 ( .A1(n6146), .A2(ADDRESS_REG_13__SCAN_IN), .ZN(n6151) );
  INV_X1 U6843 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n7195) );
  INV_X1 U6844 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n7194) );
  AOI22_X1 U6845 ( .A1(n7195), .A2(keyinput_86), .B1(n7194), .B2(keyinput_87), 
        .ZN(n6149) );
  AOI22_X1 U6846 ( .A1(ADDRESS_REG_15__SCAN_IN), .A2(keyinput_85), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(keyinput_83), .ZN(n6148) );
  AOI22_X1 U6847 ( .A1(ADDRESS_REG_18__SCAN_IN), .A2(keyinput_82), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(keyinput_81), .ZN(n6147) );
  AND3_X1 U6848 ( .A1(n6149), .A2(n6148), .A3(n6147), .ZN(n6150) );
  OAI211_X1 U6849 ( .C1(ADDRESS_REG_19__SCAN_IN), .C2(keyinput_81), .A(n6151), 
        .B(n6150), .ZN(n6154) );
  OAI22_X1 U6850 ( .A1(ADDRESS_REG_18__SCAN_IN), .A2(keyinput_82), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(keyinput_85), .ZN(n6153) );
  OAI22_X1 U6851 ( .A1(n7195), .A2(keyinput_86), .B1(ADDRESS_REG_17__SCAN_IN), 
        .B2(keyinput_83), .ZN(n6152) );
  OR4_X1 U6852 ( .A1(n6155), .A2(n6154), .A3(n6153), .A4(n6152), .ZN(n6157) );
  XOR2_X1 U6853 ( .A(ADDRESS_REG_12__SCAN_IN), .B(keyinput_88), .Z(n6156) );
  OAI21_X1 U6854 ( .B1(n6158), .B2(n6157), .A(n6156), .ZN(n6161) );
  INV_X1 U6855 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n7189) );
  XNOR2_X1 U6856 ( .A(n7189), .B(keyinput_89), .ZN(n6160) );
  XOR2_X1 U6857 ( .A(ADDRESS_REG_10__SCAN_IN), .B(keyinput_90), .Z(n6159) );
  AOI21_X1 U6858 ( .B1(n6161), .B2(n6160), .A(n6159), .ZN(n6170) );
  INV_X1 U6859 ( .A(keyinput_93), .ZN(n6162) );
  XNOR2_X1 U6860 ( .A(n6162), .B(ADDRESS_REG_7__SCAN_IN), .ZN(n6166) );
  XNOR2_X1 U6861 ( .A(ADDRESS_REG_8__SCAN_IN), .B(keyinput_92), .ZN(n6165) );
  XNOR2_X1 U6862 ( .A(ADDRESS_REG_6__SCAN_IN), .B(keyinput_94), .ZN(n6164) );
  XNOR2_X1 U6863 ( .A(ADDRESS_REG_9__SCAN_IN), .B(keyinput_91), .ZN(n6163) );
  NAND4_X1 U6864 ( .A1(n6166), .A2(n6165), .A3(n6164), .A4(n6163), .ZN(n6169)
         );
  XNOR2_X1 U6865 ( .A(ADDRESS_REG_4__SCAN_IN), .B(keyinput_96), .ZN(n6168) );
  XNOR2_X1 U6866 ( .A(ADDRESS_REG_5__SCAN_IN), .B(keyinput_95), .ZN(n6167) );
  OAI211_X1 U6867 ( .C1(n6170), .C2(n6169), .A(n6168), .B(n6167), .ZN(n6179)
         );
  XOR2_X1 U6868 ( .A(ADDRESS_REG_3__SCAN_IN), .B(keyinput_97), .Z(n6178) );
  XOR2_X1 U6869 ( .A(STATE_REG_2__SCAN_IN), .B(keyinput_101), .Z(n6173) );
  XNOR2_X1 U6870 ( .A(n6361), .B(keyinput_102), .ZN(n6172) );
  XNOR2_X1 U6871 ( .A(ADDRESS_REG_0__SCAN_IN), .B(keyinput_100), .ZN(n6171) );
  NOR3_X1 U6872 ( .A1(n6173), .A2(n6172), .A3(n6171), .ZN(n6176) );
  XOR2_X1 U6873 ( .A(ADDRESS_REG_1__SCAN_IN), .B(keyinput_99), .Z(n6175) );
  XOR2_X1 U6874 ( .A(ADDRESS_REG_2__SCAN_IN), .B(keyinput_98), .Z(n6174) );
  NAND3_X1 U6875 ( .A1(n6176), .A2(n6175), .A3(n6174), .ZN(n6177) );
  AOI21_X1 U6876 ( .B1(n6179), .B2(n6178), .A(n6177), .ZN(n6186) );
  XNOR2_X1 U6877 ( .A(n7619), .B(keyinput_103), .ZN(n6185) );
  INV_X1 U6878 ( .A(DATAWIDTH_REG_2__SCAN_IN), .ZN(n7110) );
  OAI22_X1 U6879 ( .A1(n7110), .A2(keyinput_106), .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(keyinput_104), .ZN(n6182) );
  INV_X1 U6880 ( .A(keyinput_106), .ZN(n6180) );
  NOR2_X1 U6881 ( .A1(n6180), .A2(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6181) );
  AOI211_X1 U6882 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(keyinput_104), .A(n6182), .B(n6181), .ZN(n6184) );
  XNOR2_X1 U6883 ( .A(DATAWIDTH_REG_1__SCAN_IN), .B(keyinput_105), .ZN(n6183)
         );
  OAI211_X1 U6884 ( .C1(n6186), .C2(n6185), .A(n6184), .B(n6183), .ZN(n6193)
         );
  XNOR2_X1 U6885 ( .A(DATAWIDTH_REG_3__SCAN_IN), .B(keyinput_107), .ZN(n6192)
         );
  XOR2_X1 U6886 ( .A(DATAWIDTH_REG_7__SCAN_IN), .B(keyinput_111), .Z(n6190) );
  INV_X1 U6887 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n7113) );
  XNOR2_X1 U6888 ( .A(n7113), .B(keyinput_110), .ZN(n6189) );
  INV_X1 U6889 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n7111) );
  XNOR2_X1 U6890 ( .A(n7111), .B(keyinput_108), .ZN(n6188) );
  INV_X1 U6891 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n7112) );
  XNOR2_X1 U6892 ( .A(n7112), .B(keyinput_109), .ZN(n6187) );
  NAND4_X1 U6893 ( .A1(n6190), .A2(n6189), .A3(n6188), .A4(n6187), .ZN(n6191)
         );
  AOI21_X1 U6894 ( .B1(n6193), .B2(n6192), .A(n6191), .ZN(n6200) );
  XOR2_X1 U6895 ( .A(DATAWIDTH_REG_8__SCAN_IN), .B(keyinput_112), .Z(n6199) );
  XNOR2_X1 U6896 ( .A(DATAWIDTH_REG_10__SCAN_IN), .B(keyinput_114), .ZN(n6197)
         );
  XNOR2_X1 U6897 ( .A(DATAWIDTH_REG_9__SCAN_IN), .B(keyinput_113), .ZN(n6196)
         );
  XNOR2_X1 U6898 ( .A(DATAWIDTH_REG_11__SCAN_IN), .B(keyinput_115), .ZN(n6195)
         );
  XNOR2_X1 U6899 ( .A(DATAWIDTH_REG_12__SCAN_IN), .B(keyinput_116), .ZN(n6194)
         );
  NOR4_X1 U6900 ( .A1(n6197), .A2(n6196), .A3(n6195), .A4(n6194), .ZN(n6198)
         );
  OAI21_X1 U6901 ( .B1(n6200), .B2(n6199), .A(n6198), .ZN(n6203) );
  XNOR2_X1 U6902 ( .A(DATAWIDTH_REG_13__SCAN_IN), .B(keyinput_117), .ZN(n6202)
         );
  INV_X1 U6903 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n7119) );
  XNOR2_X1 U6904 ( .A(n7119), .B(keyinput_118), .ZN(n6201) );
  AOI21_X1 U6905 ( .B1(n6203), .B2(n6202), .A(n6201), .ZN(n6206) );
  XNOR2_X1 U6906 ( .A(DATAWIDTH_REG_15__SCAN_IN), .B(keyinput_119), .ZN(n6205)
         );
  INV_X1 U6907 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n7121) );
  XNOR2_X1 U6908 ( .A(n7121), .B(keyinput_120), .ZN(n6204) );
  OAI21_X1 U6909 ( .B1(n6206), .B2(n6205), .A(n6204), .ZN(n6209) );
  XNOR2_X1 U6910 ( .A(DATAWIDTH_REG_17__SCAN_IN), .B(keyinput_121), .ZN(n6208)
         );
  INV_X1 U6911 ( .A(DATAWIDTH_REG_18__SCAN_IN), .ZN(n7123) );
  XNOR2_X1 U6912 ( .A(n7123), .B(keyinput_122), .ZN(n6207) );
  AOI21_X1 U6913 ( .B1(n6209), .B2(n6208), .A(n6207), .ZN(n6212) );
  INV_X1 U6914 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n7124) );
  XNOR2_X1 U6915 ( .A(n7124), .B(keyinput_123), .ZN(n6211) );
  XNOR2_X1 U6916 ( .A(DATAWIDTH_REG_20__SCAN_IN), .B(keyinput_124), .ZN(n6210)
         );
  OAI21_X1 U6917 ( .B1(n6212), .B2(n6211), .A(n6210), .ZN(n6215) );
  INV_X1 U6918 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n7126) );
  XNOR2_X1 U6919 ( .A(n7126), .B(keyinput_125), .ZN(n6214) );
  XNOR2_X1 U6920 ( .A(DATAWIDTH_REG_22__SCAN_IN), .B(keyinput_126), .ZN(n6213)
         );
  NAND3_X1 U6921 ( .A1(n6215), .A2(n6214), .A3(n6213), .ZN(n6408) );
  INV_X1 U6922 ( .A(keyinput_255), .ZN(n6403) );
  INV_X1 U6923 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6402) );
  XOR2_X1 U6924 ( .A(DATAI_30_), .B(keyinput_129), .Z(n6218) );
  XOR2_X1 U6925 ( .A(DATAI_31_), .B(keyinput_128), .Z(n6217) );
  XNOR2_X1 U6926 ( .A(DATAI_27_), .B(keyinput_132), .ZN(n6216) );
  AOI21_X1 U6927 ( .B1(n6218), .B2(n6217), .A(n6216), .ZN(n6221) );
  XNOR2_X1 U6928 ( .A(DATAI_28_), .B(keyinput_131), .ZN(n6220) );
  XNOR2_X1 U6929 ( .A(DATAI_29_), .B(keyinput_130), .ZN(n6219) );
  NAND3_X1 U6930 ( .A1(n6221), .A2(n6220), .A3(n6219), .ZN(n6224) );
  XNOR2_X1 U6931 ( .A(DATAI_26_), .B(keyinput_133), .ZN(n6223) );
  XNOR2_X1 U6932 ( .A(DATAI_25_), .B(keyinput_134), .ZN(n6222) );
  AOI21_X1 U6933 ( .B1(n6224), .B2(n6223), .A(n6222), .ZN(n6227) );
  XOR2_X1 U6934 ( .A(DATAI_24_), .B(keyinput_135), .Z(n6226) );
  XNOR2_X1 U6935 ( .A(DATAI_23_), .B(keyinput_136), .ZN(n6225) );
  NOR3_X1 U6936 ( .A1(n6227), .A2(n6226), .A3(n6225), .ZN(n6230) );
  XOR2_X1 U6937 ( .A(DATAI_22_), .B(keyinput_137), .Z(n6229) );
  XNOR2_X1 U6938 ( .A(DATAI_21_), .B(keyinput_138), .ZN(n6228) );
  NOR3_X1 U6939 ( .A1(n6230), .A2(n6229), .A3(n6228), .ZN(n6233) );
  XOR2_X1 U6940 ( .A(DATAI_20_), .B(keyinput_139), .Z(n6232) );
  XNOR2_X1 U6941 ( .A(DATAI_19_), .B(keyinput_140), .ZN(n6231) );
  NOR3_X1 U6942 ( .A1(n6233), .A2(n6232), .A3(n6231), .ZN(n6236) );
  XOR2_X1 U6943 ( .A(keyinput_141), .B(DATAI_18_), .Z(n6235) );
  XOR2_X1 U6944 ( .A(keyinput_142), .B(DATAI_17_), .Z(n6234) );
  OAI21_X1 U6945 ( .B1(n6236), .B2(n6235), .A(n6234), .ZN(n6239) );
  XNOR2_X1 U6946 ( .A(keyinput_143), .B(DATAI_16_), .ZN(n6238) );
  XNOR2_X1 U6947 ( .A(keyinput_144), .B(DATAI_15_), .ZN(n6237) );
  AOI21_X1 U6948 ( .B1(n6239), .B2(n6238), .A(n6237), .ZN(n6242) );
  XOR2_X1 U6949 ( .A(DATAI_14_), .B(keyinput_145), .Z(n6241) );
  XOR2_X1 U6950 ( .A(DATAI_13_), .B(keyinput_146), .Z(n6240) );
  OAI21_X1 U6951 ( .B1(n6242), .B2(n6241), .A(n6240), .ZN(n6249) );
  XNOR2_X1 U6952 ( .A(DATAI_12_), .B(keyinput_147), .ZN(n6248) );
  XOR2_X1 U6953 ( .A(DATAI_11_), .B(keyinput_148), .Z(n6246) );
  XOR2_X1 U6954 ( .A(DATAI_10_), .B(keyinput_149), .Z(n6245) );
  XNOR2_X1 U6955 ( .A(DATAI_8_), .B(keyinput_151), .ZN(n6244) );
  XNOR2_X1 U6956 ( .A(DATAI_9_), .B(keyinput_150), .ZN(n6243) );
  NAND4_X1 U6957 ( .A1(n6246), .A2(n6245), .A3(n6244), .A4(n6243), .ZN(n6247)
         );
  AOI21_X1 U6958 ( .B1(n6249), .B2(n6248), .A(n6247), .ZN(n6263) );
  XOR2_X1 U6959 ( .A(keyinput_156), .B(DATAI_3_), .Z(n6256) );
  OAI22_X1 U6960 ( .A1(keyinput_154), .A2(DATAI_5_), .B1(keyinput_159), .B2(
        DATAI_0_), .ZN(n6255) );
  NOR2_X1 U6961 ( .A1(n6250), .A2(keyinput_157), .ZN(n6254) );
  AOI22_X1 U6962 ( .A1(keyinput_152), .A2(DATAI_7_), .B1(n6250), .B2(
        keyinput_157), .ZN(n6252) );
  AOI22_X1 U6963 ( .A1(DATAI_5_), .A2(keyinput_154), .B1(DATAI_0_), .B2(
        keyinput_159), .ZN(n6251) );
  OAI211_X1 U6964 ( .C1(keyinput_152), .C2(DATAI_7_), .A(n6252), .B(n6251), 
        .ZN(n6253) );
  NOR4_X1 U6965 ( .A1(n6256), .A2(n6255), .A3(n6254), .A4(n6253), .ZN(n6260)
         );
  XNOR2_X1 U6966 ( .A(DATAI_6_), .B(keyinput_153), .ZN(n6259) );
  XNOR2_X1 U6967 ( .A(DATAI_4_), .B(keyinput_155), .ZN(n6258) );
  XNOR2_X1 U6968 ( .A(keyinput_158), .B(DATAI_1_), .ZN(n6257) );
  NAND4_X1 U6969 ( .A1(n6260), .A2(n6259), .A3(n6258), .A4(n6257), .ZN(n6262)
         );
  XNOR2_X1 U6970 ( .A(keyinput_160), .B(MEMORYFETCH_REG_SCAN_IN), .ZN(n6261)
         );
  OAI21_X1 U6971 ( .B1(n6263), .B2(n6262), .A(n6261), .ZN(n6267) );
  XOR2_X1 U6972 ( .A(keyinput_161), .B(NA_N), .Z(n6266) );
  XNOR2_X1 U6973 ( .A(n7634), .B(keyinput_163), .ZN(n6265) );
  XNOR2_X1 U6974 ( .A(keyinput_162), .B(BS16_N), .ZN(n6264) );
  NAND4_X1 U6975 ( .A1(n6267), .A2(n6266), .A3(n6265), .A4(n6264), .ZN(n6269)
         );
  XNOR2_X1 U6976 ( .A(keyinput_164), .B(HOLD), .ZN(n6268) );
  NAND2_X1 U6977 ( .A1(n6269), .A2(n6268), .ZN(n6273) );
  XOR2_X1 U6978 ( .A(keyinput_167), .B(CODEFETCH_REG_SCAN_IN), .Z(n6272) );
  XNOR2_X1 U6979 ( .A(keyinput_166), .B(ADS_N_REG_SCAN_IN), .ZN(n6271) );
  XNOR2_X1 U6980 ( .A(keyinput_165), .B(READREQUEST_REG_SCAN_IN), .ZN(n6270)
         );
  NAND4_X1 U6981 ( .A1(n6273), .A2(n6272), .A3(n6271), .A4(n6270), .ZN(n6276)
         );
  XNOR2_X1 U6982 ( .A(keyinput_168), .B(M_IO_N_REG_SCAN_IN), .ZN(n6275) );
  INV_X1 U6983 ( .A(D_C_N_REG_SCAN_IN), .ZN(n7303) );
  XNOR2_X1 U6984 ( .A(n7303), .B(keyinput_169), .ZN(n6274) );
  AOI21_X1 U6985 ( .B1(n6276), .B2(n6275), .A(n6274), .ZN(n6279) );
  XNOR2_X1 U6986 ( .A(STATEBS16_REG_SCAN_IN), .B(keyinput_171), .ZN(n6278) );
  XNOR2_X1 U6987 ( .A(keyinput_170), .B(REQUESTPENDING_REG_SCAN_IN), .ZN(n6277) );
  NOR3_X1 U6988 ( .A1(n6279), .A2(n6278), .A3(n6277), .ZN(n6282) );
  XOR2_X1 U6989 ( .A(keyinput_172), .B(MORE_REG_SCAN_IN), .Z(n6281) );
  XNOR2_X1 U6990 ( .A(keyinput_173), .B(FLUSH_REG_SCAN_IN), .ZN(n6280) );
  NOR3_X1 U6991 ( .A1(n6282), .A2(n6281), .A3(n6280), .ZN(n6288) );
  XNOR2_X1 U6992 ( .A(keyinput_174), .B(W_R_N_REG_SCAN_IN), .ZN(n6287) );
  XNOR2_X1 U6993 ( .A(keyinput_175), .B(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6285)
         );
  XNOR2_X1 U6994 ( .A(keyinput_177), .B(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6284)
         );
  XNOR2_X1 U6995 ( .A(keyinput_176), .B(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6283)
         );
  NOR3_X1 U6996 ( .A1(n6285), .A2(n6284), .A3(n6283), .ZN(n6286) );
  OAI21_X1 U6997 ( .B1(n6288), .B2(n6287), .A(n6286), .ZN(n6292) );
  XNOR2_X1 U6998 ( .A(n7232), .B(keyinput_178), .ZN(n6291) );
  XOR2_X1 U6999 ( .A(REIP_REG_30__SCAN_IN), .B(keyinput_180), .Z(n6290) );
  XNOR2_X1 U7000 ( .A(REIP_REG_31__SCAN_IN), .B(keyinput_179), .ZN(n6289) );
  AOI211_X1 U7001 ( .C1(n6292), .C2(n6291), .A(n6290), .B(n6289), .ZN(n6300)
         );
  XNOR2_X1 U7002 ( .A(REIP_REG_28__SCAN_IN), .B(keyinput_182), .ZN(n6299) );
  XNOR2_X1 U7003 ( .A(REIP_REG_29__SCAN_IN), .B(keyinput_181), .ZN(n6298) );
  XOR2_X1 U7004 ( .A(REIP_REG_25__SCAN_IN), .B(keyinput_185), .Z(n6296) );
  XNOR2_X1 U7005 ( .A(REIP_REG_24__SCAN_IN), .B(keyinput_186), .ZN(n6295) );
  XNOR2_X1 U7006 ( .A(REIP_REG_26__SCAN_IN), .B(keyinput_184), .ZN(n6294) );
  XNOR2_X1 U7007 ( .A(REIP_REG_27__SCAN_IN), .B(keyinput_183), .ZN(n6293) );
  NAND4_X1 U7008 ( .A1(n6296), .A2(n6295), .A3(n6294), .A4(n6293), .ZN(n6297)
         );
  NOR4_X1 U7009 ( .A1(n6300), .A2(n6299), .A3(n6298), .A4(n6297), .ZN(n6304)
         );
  XOR2_X1 U7010 ( .A(REIP_REG_23__SCAN_IN), .B(keyinput_187), .Z(n6303) );
  XNOR2_X1 U7011 ( .A(REIP_REG_21__SCAN_IN), .B(keyinput_189), .ZN(n6302) );
  XNOR2_X1 U7012 ( .A(REIP_REG_22__SCAN_IN), .B(keyinput_188), .ZN(n6301) );
  OAI211_X1 U7013 ( .C1(n6304), .C2(n6303), .A(n6302), .B(n6301), .ZN(n6307)
         );
  XOR2_X1 U7014 ( .A(REIP_REG_19__SCAN_IN), .B(keyinput_191), .Z(n6306) );
  XNOR2_X1 U7015 ( .A(REIP_REG_20__SCAN_IN), .B(keyinput_190), .ZN(n6305) );
  NAND3_X1 U7016 ( .A1(n6307), .A2(n6306), .A3(n6305), .ZN(n6311) );
  XOR2_X1 U7017 ( .A(REIP_REG_18__SCAN_IN), .B(keyinput_192), .Z(n6310) );
  XNOR2_X1 U7018 ( .A(REIP_REG_16__SCAN_IN), .B(keyinput_194), .ZN(n6309) );
  XNOR2_X1 U7019 ( .A(REIP_REG_17__SCAN_IN), .B(keyinput_193), .ZN(n6308) );
  NAND4_X1 U7020 ( .A1(n6311), .A2(n6310), .A3(n6309), .A4(n6308), .ZN(n6314)
         );
  XOR2_X1 U7021 ( .A(keyinput_196), .B(BE_N_REG_2__SCAN_IN), .Z(n6313) );
  XNOR2_X1 U7022 ( .A(keyinput_195), .B(BE_N_REG_3__SCAN_IN), .ZN(n6312) );
  NAND3_X1 U7023 ( .A1(n6314), .A2(n6313), .A3(n6312), .ZN(n6318) );
  XNOR2_X1 U7024 ( .A(keyinput_197), .B(BE_N_REG_1__SCAN_IN), .ZN(n6317) );
  XNOR2_X1 U7025 ( .A(n7228), .B(keyinput_199), .ZN(n6316) );
  XNOR2_X1 U7026 ( .A(keyinput_198), .B(BE_N_REG_0__SCAN_IN), .ZN(n6315) );
  AOI211_X1 U7027 ( .C1(n6318), .C2(n6317), .A(n6316), .B(n6315), .ZN(n6321)
         );
  XNOR2_X1 U7028 ( .A(n7225), .B(keyinput_200), .ZN(n6320) );
  XNOR2_X1 U7029 ( .A(keyinput_201), .B(ADDRESS_REG_27__SCAN_IN), .ZN(n6319)
         );
  OAI21_X1 U7030 ( .B1(n6321), .B2(n6320), .A(n6319), .ZN(n6324) );
  XNOR2_X1 U7031 ( .A(n7220), .B(keyinput_202), .ZN(n6323) );
  XNOR2_X1 U7032 ( .A(keyinput_203), .B(ADDRESS_REG_25__SCAN_IN), .ZN(n6322)
         );
  AOI21_X1 U7033 ( .B1(n6324), .B2(n6323), .A(n6322), .ZN(n6328) );
  INV_X1 U7034 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n7215) );
  XNOR2_X1 U7035 ( .A(n7215), .B(keyinput_204), .ZN(n6327) );
  XNOR2_X1 U7036 ( .A(keyinput_205), .B(ADDRESS_REG_23__SCAN_IN), .ZN(n6326)
         );
  XNOR2_X1 U7037 ( .A(keyinput_206), .B(ADDRESS_REG_22__SCAN_IN), .ZN(n6325)
         );
  OAI211_X1 U7038 ( .C1(n6328), .C2(n6327), .A(n6326), .B(n6325), .ZN(n6331)
         );
  XOR2_X1 U7039 ( .A(keyinput_207), .B(ADDRESS_REG_21__SCAN_IN), .Z(n6330) );
  XOR2_X1 U7040 ( .A(keyinput_208), .B(ADDRESS_REG_20__SCAN_IN), .Z(n6329) );
  NAND3_X1 U7041 ( .A1(n6331), .A2(n6330), .A3(n6329), .ZN(n6343) );
  INV_X1 U7042 ( .A(keyinput_209), .ZN(n6336) );
  INV_X1 U7043 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n7202) );
  INV_X1 U7044 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n7205) );
  OAI22_X1 U7045 ( .A1(n7202), .A2(keyinput_211), .B1(n7205), .B2(keyinput_209), .ZN(n6334) );
  OAI22_X1 U7046 ( .A1(ADDRESS_REG_16__SCAN_IN), .A2(keyinput_212), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(keyinput_213), .ZN(n6333) );
  OAI22_X1 U7047 ( .A1(n7195), .A2(keyinput_214), .B1(ADDRESS_REG_13__SCAN_IN), 
        .B2(keyinput_215), .ZN(n6332) );
  NOR3_X1 U7048 ( .A1(n6334), .A2(n6333), .A3(n6332), .ZN(n6335) );
  OAI21_X1 U7049 ( .B1(n6336), .B2(ADDRESS_REG_19__SCAN_IN), .A(n6335), .ZN(
        n6340) );
  AOI22_X1 U7050 ( .A1(n7202), .A2(keyinput_211), .B1(keyinput_213), .B2(
        ADDRESS_REG_15__SCAN_IN), .ZN(n6338) );
  AOI22_X1 U7051 ( .A1(n7195), .A2(keyinput_214), .B1(ADDRESS_REG_16__SCAN_IN), 
        .B2(keyinput_212), .ZN(n6337) );
  NAND2_X1 U7052 ( .A1(n6338), .A2(n6337), .ZN(n6339) );
  AOI211_X1 U7053 ( .C1(ADDRESS_REG_13__SCAN_IN), .C2(keyinput_215), .A(n6340), 
        .B(n6339), .ZN(n6342) );
  XNOR2_X1 U7054 ( .A(keyinput_210), .B(ADDRESS_REG_18__SCAN_IN), .ZN(n6341)
         );
  NAND3_X1 U7055 ( .A1(n6343), .A2(n6342), .A3(n6341), .ZN(n6346) );
  XOR2_X1 U7056 ( .A(keyinput_216), .B(ADDRESS_REG_12__SCAN_IN), .Z(n6345) );
  XNOR2_X1 U7057 ( .A(n7189), .B(keyinput_217), .ZN(n6344) );
  AOI21_X1 U7058 ( .B1(n6346), .B2(n6345), .A(n6344), .ZN(n6353) );
  XNOR2_X1 U7059 ( .A(keyinput_218), .B(ADDRESS_REG_10__SCAN_IN), .ZN(n6352)
         );
  INV_X1 U7060 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n7180) );
  XNOR2_X1 U7061 ( .A(n7180), .B(keyinput_222), .ZN(n6350) );
  INV_X1 U7062 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n7186) );
  XNOR2_X1 U7063 ( .A(n7186), .B(keyinput_219), .ZN(n6349) );
  XNOR2_X1 U7064 ( .A(keyinput_220), .B(ADDRESS_REG_8__SCAN_IN), .ZN(n6348) );
  XNOR2_X1 U7065 ( .A(keyinput_221), .B(ADDRESS_REG_7__SCAN_IN), .ZN(n6347) );
  NOR4_X1 U7066 ( .A1(n6350), .A2(n6349), .A3(n6348), .A4(n6347), .ZN(n6351)
         );
  OAI21_X1 U7067 ( .B1(n6353), .B2(n6352), .A(n6351), .ZN(n6356) );
  INV_X1 U7068 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n7178) );
  XNOR2_X1 U7069 ( .A(n7178), .B(keyinput_224), .ZN(n6355) );
  XNOR2_X1 U7070 ( .A(keyinput_223), .B(ADDRESS_REG_5__SCAN_IN), .ZN(n6354) );
  NAND3_X1 U7071 ( .A1(n6356), .A2(n6355), .A3(n6354), .ZN(n6358) );
  XOR2_X1 U7072 ( .A(keyinput_225), .B(ADDRESS_REG_3__SCAN_IN), .Z(n6357) );
  NAND2_X1 U7073 ( .A1(n6358), .A2(n6357), .ZN(n6365) );
  INV_X1 U7074 ( .A(STATE_REG_2__SCAN_IN), .ZN(n7621) );
  INV_X1 U7075 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n7172) );
  OAI22_X1 U7076 ( .A1(n7621), .A2(keyinput_229), .B1(n7172), .B2(keyinput_228), .ZN(n6359) );
  AOI221_X1 U7077 ( .B1(n7621), .B2(keyinput_229), .C1(keyinput_228), .C2(
        n7172), .A(n6359), .ZN(n6364) );
  XOR2_X1 U7078 ( .A(keyinput_227), .B(ADDRESS_REG_1__SCAN_IN), .Z(n6363) );
  OAI22_X1 U7079 ( .A1(n6361), .A2(keyinput_230), .B1(ADDRESS_REG_2__SCAN_IN), 
        .B2(keyinput_226), .ZN(n6360) );
  AOI221_X1 U7080 ( .B1(n6361), .B2(keyinput_230), .C1(keyinput_226), .C2(
        ADDRESS_REG_2__SCAN_IN), .A(n6360), .ZN(n6362) );
  NAND4_X1 U7081 ( .A1(n6365), .A2(n6364), .A3(n6363), .A4(n6362), .ZN(n6371)
         );
  XNOR2_X1 U7082 ( .A(n7619), .B(keyinput_231), .ZN(n6370) );
  XOR2_X1 U7083 ( .A(keyinput_232), .B(DATAWIDTH_REG_0__SCAN_IN), .Z(n6368) );
  INV_X1 U7084 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7610) );
  XNOR2_X1 U7085 ( .A(n7610), .B(keyinput_233), .ZN(n6367) );
  XNOR2_X1 U7086 ( .A(keyinput_234), .B(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6366)
         );
  NAND3_X1 U7087 ( .A1(n6368), .A2(n6367), .A3(n6366), .ZN(n6369) );
  AOI21_X1 U7088 ( .B1(n6371), .B2(n6370), .A(n6369), .ZN(n6378) );
  XOR2_X1 U7089 ( .A(keyinput_235), .B(DATAWIDTH_REG_3__SCAN_IN), .Z(n6377) );
  XNOR2_X1 U7090 ( .A(n7112), .B(keyinput_237), .ZN(n6375) );
  XNOR2_X1 U7091 ( .A(n7111), .B(keyinput_236), .ZN(n6374) );
  XNOR2_X1 U7092 ( .A(n7113), .B(keyinput_238), .ZN(n6373) );
  XNOR2_X1 U7093 ( .A(keyinput_239), .B(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6372)
         );
  NOR4_X1 U7094 ( .A1(n6375), .A2(n6374), .A3(n6373), .A4(n6372), .ZN(n6376)
         );
  OAI21_X1 U7095 ( .B1(n6378), .B2(n6377), .A(n6376), .ZN(n6385) );
  XOR2_X1 U7096 ( .A(keyinput_240), .B(DATAWIDTH_REG_8__SCAN_IN), .Z(n6384) );
  XNOR2_X1 U7097 ( .A(keyinput_244), .B(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6382)
         );
  XNOR2_X1 U7098 ( .A(keyinput_241), .B(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6381)
         );
  XNOR2_X1 U7099 ( .A(keyinput_242), .B(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6380)
         );
  XNOR2_X1 U7100 ( .A(keyinput_243), .B(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6379)
         );
  NAND4_X1 U7101 ( .A1(n6382), .A2(n6381), .A3(n6380), .A4(n6379), .ZN(n6383)
         );
  AOI21_X1 U7102 ( .B1(n6385), .B2(n6384), .A(n6383), .ZN(n6388) );
  XNOR2_X1 U7103 ( .A(keyinput_245), .B(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6387)
         );
  XNOR2_X1 U7104 ( .A(n7119), .B(keyinput_246), .ZN(n6386) );
  OAI21_X1 U7105 ( .B1(n6388), .B2(n6387), .A(n6386), .ZN(n6391) );
  INV_X1 U7106 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n7120) );
  XNOR2_X1 U7107 ( .A(n7120), .B(keyinput_247), .ZN(n6390) );
  XNOR2_X1 U7108 ( .A(n7121), .B(keyinput_248), .ZN(n6389) );
  AOI21_X1 U7109 ( .B1(n6391), .B2(n6390), .A(n6389), .ZN(n6394) );
  INV_X1 U7110 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n7122) );
  XNOR2_X1 U7111 ( .A(n7122), .B(keyinput_249), .ZN(n6393) );
  XNOR2_X1 U7112 ( .A(keyinput_250), .B(DATAWIDTH_REG_18__SCAN_IN), .ZN(n6392)
         );
  OAI21_X1 U7113 ( .B1(n6394), .B2(n6393), .A(n6392), .ZN(n6397) );
  XNOR2_X1 U7114 ( .A(n7124), .B(keyinput_251), .ZN(n6396) );
  INV_X1 U7115 ( .A(DATAWIDTH_REG_20__SCAN_IN), .ZN(n7125) );
  XNOR2_X1 U7116 ( .A(n7125), .B(keyinput_252), .ZN(n6395) );
  AOI21_X1 U7117 ( .B1(n6397), .B2(n6396), .A(n6395), .ZN(n6400) );
  XNOR2_X1 U7118 ( .A(n7126), .B(keyinput_253), .ZN(n6399) );
  XNOR2_X1 U7119 ( .A(keyinput_254), .B(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6398)
         );
  NOR3_X1 U7120 ( .A1(n6400), .A2(n6399), .A3(n6398), .ZN(n6401) );
  AOI21_X1 U7121 ( .B1(n6403), .B2(n6402), .A(n6401), .ZN(n6406) );
  INV_X1 U7122 ( .A(n6406), .ZN(n6404) );
  NOR2_X1 U7123 ( .A1(n6404), .A2(keyinput_255), .ZN(n6405) );
  OAI22_X1 U7124 ( .A1(n6406), .A2(DATAWIDTH_REG_23__SCAN_IN), .B1(
        keyinput_127), .B2(n6405), .ZN(n6407) );
  OAI211_X1 U7125 ( .C1(keyinput_127), .C2(DATAWIDTH_REG_23__SCAN_IN), .A(
        n6408), .B(n6407), .ZN(n6422) );
  NAND2_X1 U7126 ( .A1(n6409), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n6418) );
  OAI22_X1 U7127 ( .A1(n6413), .A2(n6412), .B1(n6411), .B2(n6410), .ZN(n6414)
         );
  AOI21_X1 U7128 ( .B1(n6416), .B2(n6415), .A(n6414), .ZN(n6417) );
  OAI211_X1 U7129 ( .C1(n6420), .C2(n6419), .A(n6418), .B(n6417), .ZN(n6421)
         );
  XNOR2_X1 U7130 ( .A(n6422), .B(n6421), .ZN(U3091) );
  AOI21_X1 U7131 ( .B1(n6425), .B2(n6424), .A(n6423), .ZN(n7364) );
  NAND2_X1 U7132 ( .A1(n7364), .A2(n7298), .ZN(n6429) );
  AND2_X1 U7133 ( .A1(n7370), .A2(REIP_REG_8__SCAN_IN), .ZN(n7360) );
  NOR2_X1 U7134 ( .A1(n7302), .A2(n6426), .ZN(n6427) );
  AOI211_X1 U7135 ( .C1(n7296), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n7360), 
        .B(n6427), .ZN(n6428) );
  OAI211_X1 U7136 ( .C1(n6976), .C2(n6430), .A(n6429), .B(n6428), .ZN(U2978)
         );
  INV_X1 U7137 ( .A(DATAI_11_), .ZN(n6431) );
  INV_X1 U7138 ( .A(EAX_REG_11__SCAN_IN), .ZN(n7679) );
  OAI222_X1 U7139 ( .A1(n6833), .A2(n6431), .B1(n6829), .B2(n7679), .C1(n6831), 
        .C2(n6967), .ZN(U2880) );
  INV_X1 U7140 ( .A(n6433), .ZN(n6434) );
  NOR2_X1 U7141 ( .A1(n6435), .A2(n6434), .ZN(n6436) );
  XNOR2_X1 U7142 ( .A(n6432), .B(n6436), .ZN(n7284) );
  INV_X1 U7143 ( .A(n6472), .ZN(n7101) );
  NOR3_X1 U7144 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6437), .A3(n7101), 
        .ZN(n6445) );
  AOI22_X1 U7145 ( .A1(n6439), .A2(n4903), .B1(n7386), .B2(n6438), .ZN(n6441)
         );
  AOI21_X1 U7146 ( .B1(n7100), .B2(n6441), .A(n6440), .ZN(n6444) );
  INV_X1 U7147 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6442) );
  OAI22_X1 U7148 ( .A1(n7090), .A2(n7480), .B1(n7088), .B2(n6442), .ZN(n6443)
         );
  NOR3_X1 U7149 ( .A1(n6445), .A2(n6444), .A3(n6443), .ZN(n6446) );
  OAI21_X1 U7150 ( .B1(n7284), .B2(n7350), .A(n6446), .ZN(U3012) );
  AOI21_X1 U7151 ( .B1(n6448), .B2(n5851), .A(n6447), .ZN(n6957) );
  INV_X1 U7152 ( .A(n6957), .ZN(n6463) );
  INV_X1 U7153 ( .A(n6955), .ZN(n6456) );
  NAND3_X1 U7154 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_11__SCAN_IN), .A3(
        n6449), .ZN(n6494) );
  INV_X1 U7155 ( .A(REIP_REG_12__SCAN_IN), .ZN(n7190) );
  OAI21_X1 U7156 ( .B1(n5837), .B2(n6451), .A(n6450), .ZN(n6452) );
  AND2_X1 U7157 ( .A1(n6452), .A2(n6484), .ZN(n7387) );
  INV_X1 U7158 ( .A(n7387), .ZN(n6459) );
  OAI22_X1 U7159 ( .A1(n7535), .A2(n6459), .B1(n6458), .B2(n7529), .ZN(n6453)
         );
  AOI211_X1 U7160 ( .C1(n7501), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n7487), 
        .B(n6453), .ZN(n6454) );
  OAI221_X1 U7161 ( .B1(REIP_REG_12__SCAN_IN), .B2(n6494), .C1(n7190), .C2(
        n6495), .A(n6454), .ZN(n6455) );
  AOI21_X1 U7162 ( .B1(n7504), .B2(n6456), .A(n6455), .ZN(n6457) );
  OAI21_X1 U7163 ( .B1(n6463), .B2(n7537), .A(n6457), .ZN(U2815) );
  OAI22_X1 U7164 ( .A1(n3659), .A2(n6459), .B1(n6458), .B2(n7259), .ZN(n6460)
         );
  AOI21_X1 U7165 ( .B1(n6957), .B2(n6793), .A(n6460), .ZN(n6461) );
  INV_X1 U7166 ( .A(n6461), .ZN(U2847) );
  INV_X1 U7167 ( .A(DATAI_12_), .ZN(n6462) );
  INV_X1 U7168 ( .A(EAX_REG_12__SCAN_IN), .ZN(n7683) );
  OAI222_X1 U7169 ( .A1(n6463), .A2(n6831), .B1(n6833), .B2(n6462), .C1(n6829), 
        .C2(n7683), .ZN(U2879) );
  AOI21_X1 U7170 ( .B1(n6466), .B2(n6465), .A(n6464), .ZN(n6473) );
  NAND2_X1 U7171 ( .A1(n6473), .A2(n7298), .ZN(n6470) );
  OAI22_X1 U7172 ( .A1(n7283), .A2(n5826), .B1(n7088), .B2(n7184), .ZN(n6467)
         );
  AOI21_X1 U7173 ( .B1(n7278), .B2(n6468), .A(n6467), .ZN(n6469) );
  OAI211_X1 U7174 ( .C1(n6976), .C2(n6471), .A(n6470), .B(n6469), .ZN(U2977)
         );
  NAND2_X1 U7175 ( .A1(n6474), .A2(n6472), .ZN(n7373) );
  NOR2_X1 U7176 ( .A1(n7362), .A2(n7373), .ZN(n7379) );
  INV_X1 U7177 ( .A(n7379), .ZN(n6480) );
  NAND2_X1 U7178 ( .A1(n6473), .A2(n7419), .ZN(n6479) );
  OAI21_X1 U7179 ( .B1(n7062), .B2(n6474), .A(n7357), .ZN(n7358) );
  AOI21_X1 U7180 ( .B1(n7063), .B2(n7362), .A(n7358), .ZN(n7060) );
  OAI21_X1 U7181 ( .B1(n6475), .B2(n7079), .A(n7060), .ZN(n7376) );
  OAI22_X1 U7182 ( .A1(n7090), .A2(n6476), .B1(n7184), .B2(n7088), .ZN(n6477)
         );
  AOI21_X1 U7183 ( .B1(n7376), .B2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n6477), 
        .ZN(n6478) );
  OAI211_X1 U7184 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6480), .A(n6479), 
        .B(n6478), .ZN(U3009) );
  XOR2_X1 U7185 ( .A(n6482), .B(n6481), .Z(n6949) );
  INV_X1 U7186 ( .A(n6503), .ZN(n6486) );
  NAND2_X1 U7187 ( .A1(n6484), .A2(n6483), .ZN(n6485) );
  NAND2_X1 U7188 ( .A1(n6486), .A2(n6485), .ZN(n7089) );
  OAI22_X1 U7189 ( .A1(n7089), .A2(n3659), .B1(n6487), .B2(n7259), .ZN(n6488)
         );
  AOI21_X1 U7190 ( .B1(n6949), .B2(n6793), .A(n6488), .ZN(n6489) );
  INV_X1 U7191 ( .A(n6489), .ZN(U2846) );
  INV_X1 U7192 ( .A(n6949), .ZN(n6830) );
  INV_X1 U7193 ( .A(n6947), .ZN(n6498) );
  AOI21_X1 U7194 ( .B1(n7501), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n7487), 
        .ZN(n6491) );
  NAND2_X1 U7195 ( .A1(n7519), .A2(EBX_REG_13__SCAN_IN), .ZN(n6490) );
  OAI211_X1 U7196 ( .C1(n7535), .C2(n7089), .A(n6491), .B(n6490), .ZN(n6497)
         );
  INV_X1 U7197 ( .A(REIP_REG_13__SCAN_IN), .ZN(n7191) );
  OAI21_X1 U7198 ( .B1(REIP_REG_13__SCAN_IN), .B2(REIP_REG_12__SCAN_IN), .A(
        n6492), .ZN(n6493) );
  OAI22_X1 U7199 ( .A1(n6495), .A2(n7191), .B1(n6494), .B2(n6493), .ZN(n6496)
         );
  AOI211_X1 U7200 ( .C1(n7504), .C2(n6498), .A(n6497), .B(n6496), .ZN(n6499)
         );
  OAI21_X1 U7201 ( .B1(n6830), .B2(n7537), .A(n6499), .ZN(U2814) );
  OAI21_X1 U7202 ( .B1(n6501), .B2(n6500), .A(n6741), .ZN(n6941) );
  INV_X1 U7203 ( .A(n6937), .ZN(n6511) );
  OR2_X1 U7204 ( .A1(n6503), .A2(n6502), .ZN(n6504) );
  NAND2_X1 U7205 ( .A1(n6745), .A2(n6504), .ZN(n7325) );
  INV_X1 U7206 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6795) );
  OAI22_X1 U7207 ( .A1(n7535), .A2(n7325), .B1(n7529), .B2(n6795), .ZN(n6510)
         );
  NAND3_X1 U7208 ( .A1(n7468), .A2(n6506), .A3(n6505), .ZN(n6508) );
  INV_X1 U7209 ( .A(REIP_REG_14__SCAN_IN), .ZN(n7193) );
  AOI21_X1 U7210 ( .B1(n7468), .B2(n6721), .A(n7466), .ZN(n6743) );
  AOI21_X1 U7211 ( .B1(n7501), .B2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n7487), 
        .ZN(n6507) );
  OAI221_X1 U7212 ( .B1(REIP_REG_14__SCAN_IN), .B2(n6508), .C1(n7193), .C2(
        n6743), .A(n6507), .ZN(n6509) );
  AOI211_X1 U7213 ( .C1(n7504), .C2(n6511), .A(n6510), .B(n6509), .ZN(n6512)
         );
  OAI21_X1 U7214 ( .B1(n6941), .B2(n7537), .A(n6512), .ZN(U2813) );
  AOI21_X1 U7215 ( .B1(n7598), .B2(n6567), .A(n6572), .ZN(n6574) );
  NOR2_X1 U7216 ( .A1(n6572), .A2(n3969), .ZN(n6514) );
  OAI21_X1 U7217 ( .B1(n6514), .B2(n6513), .A(n7598), .ZN(n6517) );
  NAND3_X1 U7218 ( .A1(n7552), .A2(n7548), .A3(n6515), .ZN(n6516) );
  OAI211_X1 U7219 ( .C1(n6574), .C2(n6518), .A(n6517), .B(n6516), .ZN(U3456)
         );
  NAND2_X1 U7220 ( .A1(n4187), .A2(n6842), .ZN(n6841) );
  INV_X1 U7221 ( .A(n6841), .ZN(n6520) );
  XNOR2_X1 U7222 ( .A(n6524), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6538)
         );
  INV_X1 U7223 ( .A(n6558), .ZN(n6526) );
  AOI21_X1 U7224 ( .B1(n6527), .B2(n6525), .A(n6526), .ZN(n6614) );
  NAND2_X1 U7225 ( .A1(n7370), .A2(REIP_REG_28__SCAN_IN), .ZN(n6535) );
  NAND2_X1 U7226 ( .A1(n7296), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6528)
         );
  OAI211_X1 U7227 ( .C1(n6620), .C2(n7302), .A(n6535), .B(n6528), .ZN(n6529)
         );
  AOI21_X1 U7228 ( .B1(n6614), .B2(n7297), .A(n6529), .ZN(n6530) );
  OAI21_X1 U7229 ( .B1(n6538), .B2(n7543), .A(n6530), .ZN(U2958) );
  INV_X1 U7230 ( .A(n6546), .ZN(n6531) );
  OAI21_X1 U7231 ( .B1(n6533), .B2(n6532), .A(n6531), .ZN(n6760) );
  OAI211_X1 U7232 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .A(n6549), .B(n6540), .ZN(n6534) );
  OAI211_X1 U7233 ( .C1(n6760), .C2(n7090), .A(n6535), .B(n6534), .ZN(n6536)
         );
  AOI21_X1 U7234 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n6977), .A(n6536), 
        .ZN(n6537) );
  OAI21_X1 U7235 ( .B1(n6538), .B2(n7350), .A(n6537), .ZN(U2990) );
  OAI21_X1 U7236 ( .B1(n6541), .B2(n6540), .A(n6539), .ZN(n6542) );
  AOI21_X1 U7237 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n4171), .A(n6543), 
        .ZN(n6544) );
  XNOR2_X1 U7238 ( .A(n6545), .B(n6544), .ZN(n6563) );
  XOR2_X1 U7239 ( .A(n6547), .B(n6546), .Z(n6758) );
  INV_X1 U7240 ( .A(n6758), .ZN(n6612) );
  NOR2_X1 U7241 ( .A1(n7088), .A2(n7224), .ZN(n6559) );
  INV_X1 U7242 ( .A(n6559), .ZN(n6551) );
  NAND3_X1 U7243 ( .A1(n6549), .A2(n6548), .A3(n6552), .ZN(n6550) );
  OAI211_X1 U7244 ( .C1(n6553), .C2(n6552), .A(n6551), .B(n6550), .ZN(n6554)
         );
  AOI21_X1 U7245 ( .B1(n6612), .B2(n7418), .A(n6554), .ZN(n6555) );
  OAI21_X1 U7246 ( .B1(n6563), .B2(n7350), .A(n6555), .ZN(U2989) );
  AOI21_X1 U7247 ( .B1(n6558), .B2(n6557), .A(n6556), .ZN(n6606) );
  AOI21_X1 U7248 ( .B1(n7296), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n6559), 
        .ZN(n6560) );
  OAI21_X1 U7249 ( .B1(n6610), .B2(n7302), .A(n6560), .ZN(n6561) );
  AOI21_X1 U7250 ( .B1(n6606), .B2(n7297), .A(n6561), .ZN(n6562) );
  OAI21_X1 U7251 ( .B1(n6563), .B2(n7543), .A(n6562), .ZN(U2957) );
  AND2_X1 U7252 ( .A1(n6565), .A2(n6564), .ZN(n6569) );
  NOR3_X1 U7253 ( .A1(n6567), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n6566), 
        .ZN(n6568) );
  AOI211_X1 U7254 ( .C1(n6570), .C2(n7548), .A(n6569), .B(n6568), .ZN(n6571)
         );
  OAI22_X1 U7255 ( .A1(n6574), .A2(n6573), .B1(n6572), .B2(n6571), .ZN(U3459)
         );
  AOI22_X1 U7256 ( .A1(n7706), .A2(DATAI_30_), .B1(n7709), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n6578) );
  AND2_X1 U7257 ( .A1(n6575), .A2(n4237), .ZN(n6576) );
  NAND2_X1 U7258 ( .A1(n7710), .A2(DATAI_14_), .ZN(n6577) );
  OAI211_X1 U7259 ( .C1(n6581), .C2(n6831), .A(n6578), .B(n6577), .ZN(U2861)
         );
  INV_X1 U7260 ( .A(EBX_REG_30__SCAN_IN), .ZN(n6580) );
  OAI222_X1 U7261 ( .A1(n7256), .A2(n6581), .B1(n6580), .B2(n7259), .C1(n6579), 
        .C2(n3659), .ZN(U2829) );
  OR2_X1 U7262 ( .A1(n6583), .A2(n6582), .ZN(n6585) );
  NOR2_X1 U7263 ( .A1(n6585), .A2(n6584), .ZN(n6592) );
  INV_X1 U7264 ( .A(n6586), .ZN(n6587) );
  NAND2_X1 U7265 ( .A1(n6588), .A2(n6587), .ZN(n6591) );
  NAND2_X1 U7266 ( .A1(n6593), .A2(n6589), .ZN(n6590) );
  OAI211_X1 U7267 ( .C1(n6593), .C2(n6592), .A(n6591), .B(n6590), .ZN(n7573)
         );
  NAND2_X1 U7268 ( .A1(n6594), .A2(n4884), .ZN(n7307) );
  AOI21_X1 U7269 ( .B1(n7307), .B2(n7131), .A(READY_N), .ZN(n7316) );
  OR2_X1 U7270 ( .A1(n6595), .A2(n7316), .ZN(n7570) );
  AND2_X1 U7271 ( .A1(n7570), .A2(n7581), .ZN(n7544) );
  MUX2_X1 U7272 ( .A(MORE_REG_SCAN_IN), .B(n7573), .S(n7544), .Z(U3471) );
  INV_X1 U7273 ( .A(n6797), .ZN(n6605) );
  INV_X1 U7274 ( .A(REIP_REG_31__SCAN_IN), .ZN(n7229) );
  NOR3_X1 U7275 ( .A1(n6597), .A2(n6756), .A3(n6596), .ZN(n6600) );
  NAND3_X1 U7276 ( .A1(REIP_REG_30__SCAN_IN), .A2(REIP_REG_29__SCAN_IN), .A3(
        n7229), .ZN(n6598) );
  NOR2_X1 U7277 ( .A1(n6607), .A2(n6598), .ZN(n6599) );
  AOI211_X1 U7278 ( .C1(PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n7501), .A(n6600), 
        .B(n6599), .ZN(n6601) );
  OAI21_X1 U7279 ( .B1(n6602), .B2(n7229), .A(n6601), .ZN(n6603) );
  AOI21_X1 U7280 ( .B1(n6755), .B2(n7521), .A(n6603), .ZN(n6604) );
  OAI21_X1 U7281 ( .B1(n6605), .B2(n7537), .A(n6604), .ZN(U2796) );
  INV_X1 U7282 ( .A(n6606), .ZN(n6802) );
  MUX2_X1 U7283 ( .A(n6607), .B(n6615), .S(REIP_REG_29__SCAN_IN), .Z(n6609) );
  AOI22_X1 U7284 ( .A1(n7519), .A2(EBX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n7501), .ZN(n6608) );
  OAI211_X1 U7285 ( .C1(n7541), .C2(n6610), .A(n6609), .B(n6608), .ZN(n6611)
         );
  AOI21_X1 U7286 ( .B1(n6612), .B2(n7521), .A(n6611), .ZN(n6613) );
  OAI21_X1 U7287 ( .B1(n6802), .B2(n7537), .A(n6613), .ZN(U2798) );
  INV_X1 U7288 ( .A(n6614), .ZN(n6805) );
  INV_X1 U7289 ( .A(n6760), .ZN(n6622) );
  INV_X1 U7290 ( .A(n6615), .ZN(n6616) );
  OAI21_X1 U7291 ( .B1(REIP_REG_28__SCAN_IN), .B2(n6617), .A(n6616), .ZN(n6619) );
  AOI22_X1 U7292 ( .A1(n7519), .A2(EBX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n7501), .ZN(n6618) );
  OAI211_X1 U7293 ( .C1(n7541), .C2(n6620), .A(n6619), .B(n6618), .ZN(n6621)
         );
  AOI21_X1 U7294 ( .B1(n6622), .B2(n7521), .A(n6621), .ZN(n6623) );
  OAI21_X1 U7295 ( .B1(n6805), .B2(n7537), .A(n6623), .ZN(U2799) );
  XNOR2_X1 U7296 ( .A(n6641), .B(n6624), .ZN(n6979) );
  OAI21_X1 U7297 ( .B1(n6625), .B2(n6626), .A(n6525), .ZN(n6840) );
  INV_X1 U7298 ( .A(n6840), .ZN(n6627) );
  NAND2_X1 U7299 ( .A1(n6627), .A2(n7522), .ZN(n6634) );
  OAI22_X1 U7300 ( .A1(n7531), .A2(n6835), .B1(n7529), .B2(n6762), .ZN(n6632)
         );
  NOR2_X1 U7301 ( .A1(n7457), .A2(n6628), .ZN(n6630) );
  INV_X1 U7302 ( .A(n6644), .ZN(n6629) );
  MUX2_X1 U7303 ( .A(n6630), .B(n6629), .S(REIP_REG_27__SCAN_IN), .Z(n6631) );
  AOI211_X1 U7304 ( .C1(n7504), .C2(n6837), .A(n6632), .B(n6631), .ZN(n6633)
         );
  OAI211_X1 U7305 ( .C1(n6979), .C2(n7535), .A(n6634), .B(n6633), .ZN(U2800)
         );
  INV_X1 U7306 ( .A(n6625), .ZN(n6636) );
  NAND2_X1 U7307 ( .A1(n6638), .A2(n6639), .ZN(n6640) );
  NAND2_X1 U7308 ( .A1(n6641), .A2(n6640), .ZN(n6991) );
  INV_X1 U7309 ( .A(n6991), .ZN(n6648) );
  AOI21_X1 U7310 ( .B1(n7468), .B2(n6642), .A(REIP_REG_26__SCAN_IN), .ZN(n6643) );
  OAI22_X1 U7311 ( .A1(n6644), .A2(n6643), .B1(n6845), .B2(n7531), .ZN(n6647)
         );
  INV_X1 U7312 ( .A(n6849), .ZN(n6645) );
  INV_X1 U7313 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6763) );
  OAI22_X1 U7314 ( .A1(n7541), .A2(n6645), .B1(n7529), .B2(n6763), .ZN(n6646)
         );
  AOI211_X1 U7315 ( .C1(n6648), .C2(n7521), .A(n6647), .B(n6646), .ZN(n6649)
         );
  OAI21_X1 U7316 ( .B1(n6846), .B2(n7537), .A(n6649), .ZN(U2801) );
  INV_X1 U7317 ( .A(n6651), .ZN(n6666) );
  INV_X1 U7318 ( .A(n6635), .ZN(n6652) );
  OAI21_X1 U7319 ( .B1(n3770), .B2(n6666), .A(n6652), .ZN(n6812) );
  INV_X1 U7320 ( .A(n6812), .ZN(n6859) );
  OR2_X1 U7321 ( .A1(n6677), .A2(n6653), .ZN(n6654) );
  NAND2_X1 U7322 ( .A1(n6638), .A2(n6654), .ZN(n6999) );
  INV_X1 U7323 ( .A(n6857), .ZN(n6660) );
  MUX2_X1 U7324 ( .A(n6655), .B(REIP_REG_24__SCAN_IN), .S(REIP_REG_25__SCAN_IN), .Z(n6658) );
  NAND2_X1 U7325 ( .A1(n7519), .A2(EBX_REG_25__SCAN_IN), .ZN(n6657) );
  NAND2_X1 U7326 ( .A1(n7501), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6656)
         );
  OAI211_X1 U7327 ( .C1(n6658), .C2(n7457), .A(n6657), .B(n6656), .ZN(n6659)
         );
  AOI21_X1 U7328 ( .B1(n7504), .B2(n6660), .A(n6659), .ZN(n6662) );
  OAI21_X1 U7329 ( .B1(n6669), .B2(n7457), .A(n7436), .ZN(n7534) );
  NAND2_X1 U7330 ( .A1(n7534), .A2(REIP_REG_25__SCAN_IN), .ZN(n6661) );
  OAI211_X1 U7331 ( .C1(n6999), .C2(n7535), .A(n6662), .B(n6661), .ZN(n6663)
         );
  AOI21_X1 U7332 ( .B1(n6859), .B2(n7522), .A(n6663), .ZN(n6664) );
  INV_X1 U7333 ( .A(n6664), .ZN(U2802) );
  AOI21_X1 U7334 ( .B1(n6667), .B2(n6665), .A(n6666), .ZN(n6874) );
  INV_X1 U7335 ( .A(n6874), .ZN(n6815) );
  NOR2_X1 U7336 ( .A1(REIP_REG_24__SCAN_IN), .A2(n7457), .ZN(n6668) );
  AOI22_X1 U7337 ( .A1(EBX_REG_24__SCAN_IN), .A2(n7519), .B1(n6669), .B2(n6668), .ZN(n6670) );
  OAI21_X1 U7338 ( .B1(n6671), .B2(n7531), .A(n6670), .ZN(n6672) );
  AOI21_X1 U7339 ( .B1(REIP_REG_24__SCAN_IN), .B2(n7534), .A(n6672), .ZN(n6680) );
  INV_X1 U7340 ( .A(n6673), .ZN(n7013) );
  INV_X1 U7341 ( .A(n6674), .ZN(n6675) );
  AOI21_X1 U7342 ( .B1(n7014), .B2(n7013), .A(n6675), .ZN(n6676) );
  OR2_X1 U7343 ( .A1(n6677), .A2(n6676), .ZN(n7004) );
  OAI22_X1 U7344 ( .A1(n7004), .A2(n7535), .B1(n6872), .B2(n7541), .ZN(n6678)
         );
  INV_X1 U7345 ( .A(n6678), .ZN(n6679) );
  OAI211_X1 U7346 ( .C1(n6815), .C2(n7537), .A(n6680), .B(n6679), .ZN(U2803)
         );
  INV_X1 U7347 ( .A(n6682), .ZN(n6683) );
  OAI21_X1 U7348 ( .B1(n6684), .B2(n6681), .A(n6683), .ZN(n6890) );
  INV_X1 U7349 ( .A(n7014), .ZN(n6685) );
  OAI21_X1 U7350 ( .B1(n6686), .B2(n6697), .A(n6685), .ZN(n7028) );
  AOI22_X1 U7351 ( .A1(n7504), .A2(n6893), .B1(n7519), .B2(EBX_REG_22__SCAN_IN), .ZN(n6687) );
  OAI21_X1 U7352 ( .B1(n7028), .B2(n7535), .A(n6687), .ZN(n6692) );
  INV_X1 U7353 ( .A(REIP_REG_21__SCAN_IN), .ZN(n7207) );
  INV_X1 U7354 ( .A(REIP_REG_22__SCAN_IN), .ZN(n7210) );
  INV_X1 U7355 ( .A(n7528), .ZN(n6688) );
  OR2_X1 U7356 ( .A1(n7457), .A2(n6689), .ZN(n7527) );
  AOI211_X1 U7357 ( .C1(n7207), .C2(n7210), .A(n6688), .B(n7527), .ZN(n6691)
         );
  AOI21_X1 U7358 ( .B1(n7468), .B2(n6689), .A(n7466), .ZN(n6712) );
  OAI22_X1 U7359 ( .A1(n6712), .A2(n7210), .B1(n6889), .B2(n7531), .ZN(n6690)
         );
  NOR3_X1 U7360 ( .A1(n6692), .A2(n6691), .A3(n6690), .ZN(n6693) );
  OAI21_X1 U7361 ( .B1(n6890), .B2(n7537), .A(n6693), .ZN(U2805) );
  NOR2_X1 U7362 ( .A1(n3667), .A2(n6694), .ZN(n6695) );
  OR2_X1 U7363 ( .A1(n6681), .A2(n6695), .ZN(n6902) );
  INV_X1 U7364 ( .A(n6902), .ZN(n7702) );
  AOI22_X1 U7365 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n7501), .B1(
        EBX_REG_21__SCAN_IN), .B2(n7519), .ZN(n6696) );
  OAI221_X1 U7366 ( .B1(REIP_REG_21__SCAN_IN), .B2(n7527), .C1(n7207), .C2(
        n6712), .A(n6696), .ZN(n6702) );
  AOI21_X1 U7367 ( .B1(n6698), .B2(n6709), .A(n6697), .ZN(n6699) );
  INV_X1 U7368 ( .A(n6699), .ZN(n7035) );
  OAI22_X1 U7369 ( .A1(n7035), .A2(n7535), .B1(n6700), .B2(n7541), .ZN(n6701)
         );
  AOI211_X1 U7370 ( .C1(n7702), .C2(n7522), .A(n6702), .B(n6701), .ZN(n6703)
         );
  INV_X1 U7371 ( .A(n6703), .ZN(U2806) );
  AND2_X1 U7372 ( .A1(n6704), .A2(n6705), .ZN(n6706) );
  OR2_X1 U7373 ( .A1(n6706), .A2(n3667), .ZN(n6906) );
  NAND2_X1 U7374 ( .A1(n3675), .A2(n6707), .ZN(n6708) );
  NAND2_X1 U7375 ( .A1(n6709), .A2(n6708), .ZN(n7043) );
  OAI22_X1 U7376 ( .A1(n7043), .A2(n7535), .B1(n6905), .B2(n7531), .ZN(n6714)
         );
  AOI21_X1 U7377 ( .B1(n7468), .B2(n6710), .A(REIP_REG_20__SCAN_IN), .ZN(n6711) );
  OAI22_X1 U7378 ( .A1(n6712), .A2(n6711), .B1(n6768), .B2(n7529), .ZN(n6713)
         );
  AOI211_X1 U7379 ( .C1(n7504), .C2(n6909), .A(n6714), .B(n6713), .ZN(n6715)
         );
  OAI21_X1 U7380 ( .B1(n6906), .B2(n7537), .A(n6715), .ZN(U2807) );
  AOI21_X1 U7381 ( .B1(n6718), .B2(n6716), .A(n6717), .ZN(n6918) );
  INV_X1 U7382 ( .A(n6918), .ZN(n6822) );
  OAI21_X1 U7383 ( .B1(n6722), .B2(n7429), .A(n6743), .ZN(n7512) );
  AOI22_X1 U7384 ( .A1(EBX_REG_18__SCAN_IN), .A2(n7519), .B1(
        REIP_REG_18__SCAN_IN), .B2(n7512), .ZN(n6719) );
  OAI211_X1 U7385 ( .C1(n7531), .C2(n6720), .A(n6719), .B(n7514), .ZN(n6727)
         );
  INV_X1 U7386 ( .A(REIP_REG_18__SCAN_IN), .ZN(n7201) );
  NOR2_X1 U7387 ( .A1(n7457), .A2(n6721), .ZN(n6734) );
  AND3_X1 U7388 ( .A1(n7201), .A2(n6722), .A3(n6734), .ZN(n7513) );
  AOI21_X1 U7389 ( .B1(n6723), .B2(n3668), .A(n3718), .ZN(n7417) );
  INV_X1 U7390 ( .A(n7417), .ZN(n6725) );
  INV_X1 U7391 ( .A(n6724), .ZN(n6916) );
  OAI22_X1 U7392 ( .A1(n6725), .A2(n7535), .B1(n6916), .B2(n7541), .ZN(n6726)
         );
  NOR3_X1 U7393 ( .A1(n6727), .A2(n7513), .A3(n6726), .ZN(n6728) );
  OAI21_X1 U7394 ( .B1(n6822), .B2(n7537), .A(n6728), .ZN(U2809) );
  AOI21_X1 U7395 ( .B1(n6731), .B2(n6729), .A(n6730), .ZN(n6924) );
  INV_X1 U7396 ( .A(n6924), .ZN(n6790) );
  INV_X1 U7397 ( .A(n6922), .ZN(n6738) );
  AOI21_X1 U7398 ( .B1(n6732), .B2(n6747), .A(n6785), .ZN(n7404) );
  INV_X1 U7399 ( .A(n7404), .ZN(n6788) );
  AOI21_X1 U7400 ( .B1(n7501), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n7487), 
        .ZN(n6733) );
  OAI21_X1 U7401 ( .B1(n6788), .B2(n7535), .A(n6733), .ZN(n6737) );
  NAND2_X1 U7402 ( .A1(n6734), .A2(n7196), .ZN(n6750) );
  INV_X1 U7403 ( .A(n6734), .ZN(n7510) );
  NOR2_X1 U7404 ( .A1(n7196), .A2(n7510), .ZN(n7506) );
  AOI22_X1 U7405 ( .A1(EBX_REG_16__SCAN_IN), .A2(n7519), .B1(n7506), .B2(n7198), .ZN(n6735) );
  OAI221_X1 U7406 ( .B1(n7198), .B2(n6743), .C1(n7198), .C2(n6750), .A(n6735), 
        .ZN(n6736) );
  AOI211_X1 U7407 ( .C1(n7504), .C2(n6738), .A(n6737), .B(n6736), .ZN(n6739)
         );
  OAI21_X1 U7408 ( .B1(n6790), .B2(n7537), .A(n6739), .ZN(U2811) );
  INV_X1 U7409 ( .A(n6729), .ZN(n6740) );
  AOI21_X1 U7410 ( .B1(n6742), .B2(n6741), .A(n6740), .ZN(n6933) );
  OAI22_X1 U7411 ( .A1(n6791), .A2(n7529), .B1(n7196), .B2(n6743), .ZN(n6753)
         );
  NAND2_X1 U7412 ( .A1(n6745), .A2(n6744), .ZN(n6746) );
  NAND2_X1 U7413 ( .A1(n6747), .A2(n6746), .ZN(n7076) );
  NOR2_X1 U7414 ( .A1(n7535), .A2(n7076), .ZN(n6748) );
  AOI211_X1 U7415 ( .C1(n7501), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n7487), 
        .B(n6748), .ZN(n6749) );
  OAI211_X1 U7416 ( .C1(n7541), .C2(n6751), .A(n6750), .B(n6749), .ZN(n6752)
         );
  AOI211_X1 U7417 ( .C1(n6933), .C2(n7522), .A(n6753), .B(n6752), .ZN(n6754)
         );
  INV_X1 U7418 ( .A(n6754), .ZN(U2812) );
  INV_X1 U7419 ( .A(n6755), .ZN(n6757) );
  OAI22_X1 U7420 ( .A1(n6757), .A2(n3659), .B1(n7259), .B2(n6756), .ZN(U2828)
         );
  OAI222_X1 U7421 ( .A1(n7256), .A2(n6802), .B1(n6759), .B2(n7259), .C1(n6758), 
        .C2(n3659), .ZN(U2830) );
  OAI222_X1 U7422 ( .A1(n7256), .A2(n6805), .B1(n6761), .B2(n7259), .C1(n6760), 
        .C2(n3659), .ZN(U2831) );
  OAI222_X1 U7423 ( .A1(n6840), .A2(n7256), .B1(n6762), .B2(n7259), .C1(n3659), 
        .C2(n6979), .ZN(U2832) );
  OAI222_X1 U7424 ( .A1(n6846), .A2(n7256), .B1(n6763), .B2(n7259), .C1(n6991), 
        .C2(n3659), .ZN(U2833) );
  OAI222_X1 U7425 ( .A1(n6812), .A2(n7256), .B1(n6764), .B2(n7259), .C1(n6999), 
        .C2(n3659), .ZN(U2834) );
  INV_X1 U7426 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6765) );
  OAI222_X1 U7427 ( .A1(n7256), .A2(n6815), .B1(n6765), .B2(n7259), .C1(n7004), 
        .C2(n3659), .ZN(U2835) );
  INV_X1 U7428 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6766) );
  OAI222_X1 U7429 ( .A1(n7256), .A2(n6890), .B1(n6766), .B2(n7259), .C1(n7028), 
        .C2(n3659), .ZN(U2837) );
  OAI222_X1 U7430 ( .A1(n6902), .A2(n7256), .B1(n6767), .B2(n7259), .C1(n3659), 
        .C2(n7035), .ZN(U2838) );
  OAI22_X1 U7431 ( .A1(n7043), .A2(n3659), .B1(n6768), .B2(n7259), .ZN(n6769)
         );
  INV_X1 U7432 ( .A(n6769), .ZN(n6770) );
  OAI21_X1 U7433 ( .B1(n6906), .B2(n7256), .A(n6770), .ZN(U2839) );
  NAND2_X1 U7434 ( .A1(n6772), .A2(n6771), .ZN(n6773) );
  AND2_X1 U7435 ( .A1(n6704), .A2(n6773), .ZN(n7699) );
  INV_X1 U7436 ( .A(n7699), .ZN(n6779) );
  NAND2_X1 U7437 ( .A1(n6775), .A2(n6774), .ZN(n6776) );
  AND2_X1 U7438 ( .A1(n3675), .A2(n6776), .ZN(n7520) );
  INV_X1 U7439 ( .A(n7520), .ZN(n6777) );
  OAI222_X1 U7440 ( .A1(n6779), .A2(n7256), .B1(n6778), .B2(n7259), .C1(n3659), 
        .C2(n6777), .ZN(U2840) );
  AOI22_X1 U7441 ( .A1(n7417), .A2(n6780), .B1(EBX_REG_18__SCAN_IN), .B2(n5152), .ZN(n6781) );
  OAI21_X1 U7442 ( .B1(n6822), .B2(n7256), .A(n6781), .ZN(U2841) );
  OR2_X1 U7443 ( .A1(n6730), .A2(n6782), .ZN(n6783) );
  AND2_X1 U7444 ( .A1(n6716), .A2(n6783), .ZN(n7696) );
  INV_X1 U7445 ( .A(n7696), .ZN(n6787) );
  OAI21_X1 U7446 ( .B1(n6785), .B2(n6784), .A(n3668), .ZN(n7502) );
  OAI222_X1 U7447 ( .A1(n6787), .A2(n7256), .B1(n6786), .B2(n7259), .C1(n3659), 
        .C2(n7502), .ZN(U2842) );
  INV_X1 U7448 ( .A(EBX_REG_16__SCAN_IN), .ZN(n6789) );
  OAI222_X1 U7449 ( .A1(n6790), .A2(n7256), .B1(n6789), .B2(n7259), .C1(n3659), 
        .C2(n6788), .ZN(U2843) );
  OAI22_X1 U7450 ( .A1(n7076), .A2(n3659), .B1(n6791), .B2(n7259), .ZN(n6792)
         );
  AOI21_X1 U7451 ( .B1(n6933), .B2(n6793), .A(n6792), .ZN(n6794) );
  INV_X1 U7452 ( .A(n6794), .ZN(U2844) );
  OAI222_X1 U7453 ( .A1(n7325), .A2(n3659), .B1(n6795), .B2(n7259), .C1(n6941), 
        .C2(n7256), .ZN(U2845) );
  AOI22_X1 U7454 ( .A1(n7706), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n7709), .ZN(n6798) );
  NAND2_X1 U7455 ( .A1(n6799), .A2(n6798), .ZN(U2860) );
  AOI22_X1 U7456 ( .A1(n7706), .A2(DATAI_29_), .B1(n7709), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6801) );
  NAND2_X1 U7457 ( .A1(n7710), .A2(DATAI_13_), .ZN(n6800) );
  OAI211_X1 U7458 ( .C1(n6802), .C2(n6831), .A(n6801), .B(n6800), .ZN(U2862)
         );
  AOI22_X1 U7459 ( .A1(n7706), .A2(DATAI_28_), .B1(n7709), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6804) );
  NAND2_X1 U7460 ( .A1(n7710), .A2(DATAI_12_), .ZN(n6803) );
  OAI211_X1 U7461 ( .C1(n6805), .C2(n6831), .A(n6804), .B(n6803), .ZN(U2863)
         );
  AOI22_X1 U7462 ( .A1(n7706), .A2(DATAI_27_), .B1(n7709), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6807) );
  NAND2_X1 U7463 ( .A1(n7710), .A2(DATAI_11_), .ZN(n6806) );
  OAI211_X1 U7464 ( .C1(n6840), .C2(n6831), .A(n6807), .B(n6806), .ZN(U2864)
         );
  AOI22_X1 U7465 ( .A1(n7706), .A2(DATAI_26_), .B1(n7709), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6809) );
  NAND2_X1 U7466 ( .A1(n7710), .A2(DATAI_10_), .ZN(n6808) );
  OAI211_X1 U7467 ( .C1(n6846), .C2(n6831), .A(n6809), .B(n6808), .ZN(U2865)
         );
  AOI22_X1 U7468 ( .A1(n7706), .A2(DATAI_25_), .B1(n7709), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6811) );
  NAND2_X1 U7469 ( .A1(n7710), .A2(DATAI_9_), .ZN(n6810) );
  OAI211_X1 U7470 ( .C1(n6812), .C2(n6831), .A(n6811), .B(n6810), .ZN(U2866)
         );
  AOI22_X1 U7471 ( .A1(n7706), .A2(DATAI_24_), .B1(n7709), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n6814) );
  NAND2_X1 U7472 ( .A1(n7710), .A2(DATAI_8_), .ZN(n6813) );
  OAI211_X1 U7473 ( .C1(n6815), .C2(n6831), .A(n6814), .B(n6813), .ZN(U2867)
         );
  AOI22_X1 U7474 ( .A1(n7706), .A2(DATAI_22_), .B1(n7709), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6817) );
  NAND2_X1 U7475 ( .A1(n7710), .A2(DATAI_6_), .ZN(n6816) );
  OAI211_X1 U7476 ( .C1(n6890), .C2(n6831), .A(n6817), .B(n6816), .ZN(U2869)
         );
  AOI22_X1 U7477 ( .A1(n7706), .A2(DATAI_20_), .B1(n7709), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6819) );
  NAND2_X1 U7478 ( .A1(n7710), .A2(DATAI_4_), .ZN(n6818) );
  OAI211_X1 U7479 ( .C1(n6906), .C2(n6831), .A(n6819), .B(n6818), .ZN(U2871)
         );
  AOI22_X1 U7480 ( .A1(n7706), .A2(DATAI_18_), .B1(n7709), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6821) );
  NAND2_X1 U7481 ( .A1(n7710), .A2(DATAI_2_), .ZN(n6820) );
  OAI211_X1 U7482 ( .C1(n6822), .C2(n6831), .A(n6821), .B(n6820), .ZN(U2873)
         );
  INV_X1 U7483 ( .A(n7710), .ZN(n6825) );
  NAND2_X1 U7484 ( .A1(n6924), .A2(n7707), .ZN(n6824) );
  AOI22_X1 U7485 ( .A1(n7706), .A2(DATAI_16_), .B1(n7709), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6823) );
  OAI211_X1 U7486 ( .C1(n5141), .C2(n6825), .A(n6824), .B(n6823), .ZN(U2875)
         );
  INV_X1 U7487 ( .A(DATAI_15_), .ZN(n6827) );
  INV_X1 U7488 ( .A(EAX_REG_15__SCAN_IN), .ZN(n7695) );
  INV_X1 U7489 ( .A(n6933), .ZN(n6826) );
  OAI222_X1 U7490 ( .A1(n6833), .A2(n6827), .B1(n6829), .B2(n7695), .C1(n6831), 
        .C2(n6826), .ZN(U2876) );
  INV_X1 U7491 ( .A(DATAI_14_), .ZN(n6828) );
  INV_X1 U7492 ( .A(EAX_REG_14__SCAN_IN), .ZN(n7690) );
  OAI222_X1 U7493 ( .A1(n6833), .A2(n6828), .B1(n6829), .B2(n7690), .C1(n6831), 
        .C2(n6941), .ZN(U2877) );
  INV_X1 U7494 ( .A(DATAI_13_), .ZN(n6832) );
  INV_X1 U7495 ( .A(EAX_REG_13__SCAN_IN), .ZN(n7686) );
  OAI222_X1 U7496 ( .A1(n6833), .A2(n6832), .B1(n6831), .B2(n6830), .C1(n7686), 
        .C2(n6829), .ZN(U2878) );
  NAND3_X1 U7497 ( .A1(n6978), .A2(n6834), .A3(n7298), .ZN(n6839) );
  NAND2_X1 U7498 ( .A1(n7370), .A2(REIP_REG_27__SCAN_IN), .ZN(n6980) );
  OAI21_X1 U7499 ( .B1(n7283), .B2(n6835), .A(n6980), .ZN(n6836) );
  AOI21_X1 U7500 ( .B1(n6837), .B2(n7278), .A(n6836), .ZN(n6838) );
  OAI211_X1 U7501 ( .C1(n6976), .C2(n6840), .A(n6839), .B(n6838), .ZN(U2959)
         );
  OAI21_X1 U7502 ( .B1(n4187), .B2(n6842), .A(n6841), .ZN(n6844) );
  XOR2_X1 U7503 ( .A(n6844), .B(n6843), .Z(n6994) );
  NAND2_X1 U7504 ( .A1(n7370), .A2(REIP_REG_26__SCAN_IN), .ZN(n6990) );
  OAI21_X1 U7505 ( .B1(n7283), .B2(n6845), .A(n6990), .ZN(n6848) );
  NOR2_X1 U7506 ( .A1(n6846), .A2(n6976), .ZN(n6847) );
  AOI211_X1 U7507 ( .C1(n7278), .C2(n6849), .A(n6848), .B(n6847), .ZN(n6850)
         );
  OAI21_X1 U7508 ( .B1(n6994), .B2(n7543), .A(n6850), .ZN(U2960) );
  AOI21_X1 U7509 ( .B1(n6853), .B2(n6855), .A(n6852), .ZN(n6854) );
  AOI21_X1 U7510 ( .B1(n6519), .B2(n6855), .A(n6854), .ZN(n7003) );
  NAND2_X1 U7511 ( .A1(n7370), .A2(REIP_REG_25__SCAN_IN), .ZN(n6998) );
  NAND2_X1 U7512 ( .A1(n7296), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6856)
         );
  OAI211_X1 U7513 ( .C1(n7302), .C2(n6857), .A(n6998), .B(n6856), .ZN(n6858)
         );
  AOI21_X1 U7514 ( .B1(n6859), .B2(n7297), .A(n6858), .ZN(n6860) );
  OAI21_X1 U7515 ( .B1(n7003), .B2(n7543), .A(n6860), .ZN(U2961) );
  INV_X1 U7516 ( .A(n6861), .ZN(n6862) );
  XNOR2_X1 U7517 ( .A(n7066), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n7052)
         );
  NAND2_X1 U7518 ( .A1(n4187), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6864) );
  XNOR2_X1 U7519 ( .A(n7066), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6895)
         );
  NAND2_X1 U7520 ( .A1(n6896), .A2(n6895), .ZN(n7032) );
  NAND2_X1 U7521 ( .A1(n6888), .A2(n6866), .ZN(n6869) );
  NAND4_X1 U7522 ( .A1(n6865), .A2(n4187), .A3(n6867), .A4(n7024), .ZN(n6880)
         );
  NAND2_X1 U7523 ( .A1(n6869), .A2(n6868), .ZN(n6870) );
  XNOR2_X1 U7524 ( .A(n6870), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n7011)
         );
  INV_X1 U7525 ( .A(REIP_REG_24__SCAN_IN), .ZN(n7212) );
  NOR2_X1 U7526 ( .A1(n7088), .A2(n7212), .ZN(n7008) );
  AOI21_X1 U7527 ( .B1(n7296), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n7008), 
        .ZN(n6871) );
  OAI21_X1 U7528 ( .B1(n6872), .B2(n7302), .A(n6871), .ZN(n6873) );
  AOI21_X1 U7529 ( .B1(n6874), .B2(n7297), .A(n6873), .ZN(n6875) );
  OAI21_X1 U7530 ( .B1(n7011), .B2(n7543), .A(n6875), .ZN(U2962) );
  OR2_X1 U7531 ( .A1(n6682), .A2(n6876), .ZN(n6877) );
  NAND2_X1 U7532 ( .A1(n6665), .A2(n6877), .ZN(n7705) );
  INV_X1 U7533 ( .A(n6878), .ZN(n6879) );
  NAND2_X1 U7534 ( .A1(n4171), .A2(n6879), .ZN(n6881) );
  OAI21_X1 U7535 ( .B1(n6882), .B2(n6881), .A(n6880), .ZN(n6883) );
  XNOR2_X1 U7536 ( .A(n6883), .B(n7016), .ZN(n7012) );
  NAND2_X1 U7537 ( .A1(n7012), .A2(n7298), .ZN(n6886) );
  NOR2_X1 U7538 ( .A1(n7088), .A2(n7526), .ZN(n7015) );
  NOR2_X1 U7539 ( .A1(n7302), .A2(n7542), .ZN(n6884) );
  AOI211_X1 U7540 ( .C1(n7296), .C2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n7015), 
        .B(n6884), .ZN(n6885) );
  OAI211_X1 U7541 ( .C1(n6976), .C2(n7705), .A(n6886), .B(n6885), .ZN(U2963)
         );
  XNOR2_X1 U7542 ( .A(n7066), .B(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6887)
         );
  XNOR2_X1 U7543 ( .A(n6888), .B(n6887), .ZN(n7031) );
  NAND2_X1 U7544 ( .A1(n7370), .A2(REIP_REG_22__SCAN_IN), .ZN(n7027) );
  OAI21_X1 U7545 ( .B1(n7283), .B2(n6889), .A(n7027), .ZN(n6892) );
  NOR2_X1 U7546 ( .A1(n6890), .A2(n6976), .ZN(n6891) );
  AOI211_X1 U7547 ( .C1(n7278), .C2(n6893), .A(n6892), .B(n6891), .ZN(n6894)
         );
  OAI21_X1 U7548 ( .B1(n7031), .B2(n7543), .A(n6894), .ZN(U2964) );
  OR2_X1 U7549 ( .A1(n6896), .A2(n6895), .ZN(n7033) );
  NAND3_X1 U7550 ( .A1(n7033), .A2(n7032), .A3(n7298), .ZN(n6901) );
  NAND2_X1 U7551 ( .A1(n7370), .A2(REIP_REG_21__SCAN_IN), .ZN(n7034) );
  OAI21_X1 U7552 ( .B1(n7283), .B2(n6897), .A(n7034), .ZN(n6898) );
  AOI21_X1 U7553 ( .B1(n7278), .B2(n6899), .A(n6898), .ZN(n6900) );
  OAI211_X1 U7554 ( .C1(n6976), .C2(n6902), .A(n6901), .B(n6900), .ZN(U2965)
         );
  NOR2_X1 U7555 ( .A1(n6865), .A2(n7044), .ZN(n6903) );
  MUX2_X1 U7556 ( .A(n6865), .B(n6903), .S(n4171), .Z(n6904) );
  XNOR2_X1 U7557 ( .A(n6904), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n7050)
         );
  NAND2_X1 U7558 ( .A1(n7370), .A2(REIP_REG_20__SCAN_IN), .ZN(n7042) );
  OAI21_X1 U7559 ( .B1(n7283), .B2(n6905), .A(n7042), .ZN(n6908) );
  NOR2_X1 U7560 ( .A1(n6906), .A2(n6976), .ZN(n6907) );
  AOI211_X1 U7561 ( .C1(n7278), .C2(n6909), .A(n6908), .B(n6907), .ZN(n6910)
         );
  OAI21_X1 U7562 ( .B1(n7050), .B2(n7543), .A(n6910), .ZN(U2966) );
  NAND2_X1 U7563 ( .A1(n6911), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6913) );
  AOI21_X1 U7564 ( .B1(n4187), .B2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n6911), 
        .ZN(n7068) );
  NAND2_X1 U7565 ( .A1(n7068), .A2(n7073), .ZN(n6912) );
  MUX2_X1 U7566 ( .A(n6913), .B(n6912), .S(n4187), .Z(n6914) );
  XNOR2_X1 U7567 ( .A(n6914), .B(n7423), .ZN(n7416) );
  AOI22_X1 U7568 ( .A1(n7296), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .B1(n7370), 
        .B2(REIP_REG_18__SCAN_IN), .ZN(n6915) );
  OAI21_X1 U7569 ( .B1(n6916), .B2(n7302), .A(n6915), .ZN(n6917) );
  AOI21_X1 U7570 ( .B1(n6918), .B2(n7297), .A(n6917), .ZN(n6919) );
  OAI21_X1 U7571 ( .B1(n7416), .B2(n7543), .A(n6919), .ZN(U2968) );
  XNOR2_X1 U7572 ( .A(n7066), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6920)
         );
  XNOR2_X1 U7573 ( .A(n3669), .B(n6920), .ZN(n7405) );
  INV_X1 U7574 ( .A(n7405), .ZN(n6926) );
  AOI22_X1 U7575 ( .A1(n7296), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n7370), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n6921) );
  OAI21_X1 U7576 ( .B1(n6922), .B2(n7302), .A(n6921), .ZN(n6923) );
  AOI21_X1 U7577 ( .B1(n6924), .B2(n7297), .A(n6923), .ZN(n6925) );
  OAI21_X1 U7578 ( .B1(n6926), .B2(n7543), .A(n6925), .ZN(U2970) );
  XNOR2_X1 U7579 ( .A(n7066), .B(n7401), .ZN(n6928) );
  XNOR2_X1 U7580 ( .A(n6927), .B(n6928), .ZN(n7087) );
  INV_X1 U7581 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6931) );
  NAND2_X1 U7582 ( .A1(n7278), .A2(n6929), .ZN(n6930) );
  NAND2_X1 U7583 ( .A1(n7370), .A2(REIP_REG_15__SCAN_IN), .ZN(n7075) );
  OAI211_X1 U7584 ( .C1(n7283), .C2(n6931), .A(n6930), .B(n7075), .ZN(n6932)
         );
  AOI21_X1 U7585 ( .B1(n6933), .B2(n7297), .A(n6932), .ZN(n6934) );
  OAI21_X1 U7586 ( .B1(n7087), .B2(n7543), .A(n6934), .ZN(U2971) );
  XNOR2_X1 U7587 ( .A(n7066), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6935)
         );
  XNOR2_X1 U7588 ( .A(n6936), .B(n6935), .ZN(n7329) );
  NAND2_X1 U7589 ( .A1(n7329), .A2(n7298), .ZN(n6940) );
  AND2_X1 U7590 ( .A1(n7370), .A2(REIP_REG_14__SCAN_IN), .ZN(n7326) );
  NOR2_X1 U7591 ( .A1(n7302), .A2(n6937), .ZN(n6938) );
  AOI211_X1 U7592 ( .C1(n7296), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n7326), 
        .B(n6938), .ZN(n6939) );
  OAI211_X1 U7593 ( .C1(n6976), .C2(n6941), .A(n6940), .B(n6939), .ZN(U2972)
         );
  OAI21_X1 U7594 ( .B1(n6944), .B2(n6943), .A(n6942), .ZN(n6945) );
  INV_X1 U7595 ( .A(n6945), .ZN(n7098) );
  AOI22_X1 U7596 ( .A1(n7296), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .B1(n7370), 
        .B2(REIP_REG_13__SCAN_IN), .ZN(n6946) );
  OAI21_X1 U7597 ( .B1(n6947), .B2(n7302), .A(n6946), .ZN(n6948) );
  AOI21_X1 U7598 ( .B1(n6949), .B2(n7297), .A(n6948), .ZN(n6950) );
  OAI21_X1 U7599 ( .B1(n7098), .B2(n7543), .A(n6950), .ZN(U2973) );
  OAI21_X1 U7600 ( .B1(n4172), .B2(n7066), .A(n6951), .ZN(n6953) );
  MUX2_X1 U7601 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .B(n4173), .S(n7066), 
        .Z(n6969) );
  NOR2_X1 U7602 ( .A1(n6970), .A2(n6969), .ZN(n6968) );
  AOI21_X1 U7603 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n4187), .A(n6968), 
        .ZN(n6962) );
  XNOR2_X1 U7604 ( .A(n7066), .B(n4174), .ZN(n6961) );
  NOR2_X1 U7605 ( .A1(n6962), .A2(n6961), .ZN(n6960) );
  AOI21_X1 U7606 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n4187), .A(n6960), 
        .ZN(n6952) );
  XOR2_X1 U7607 ( .A(n6953), .B(n6952), .Z(n7388) );
  INV_X1 U7608 ( .A(n7388), .ZN(n6959) );
  AOI22_X1 U7609 ( .A1(n7296), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .B1(n7370), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n6954) );
  OAI21_X1 U7610 ( .B1(n6955), .B2(n7302), .A(n6954), .ZN(n6956) );
  AOI21_X1 U7611 ( .B1(n6957), .B2(n7297), .A(n6956), .ZN(n6958) );
  OAI21_X1 U7612 ( .B1(n6959), .B2(n7543), .A(n6958), .ZN(U2974) );
  AOI21_X1 U7613 ( .B1(n6962), .B2(n6961), .A(n6960), .ZN(n7397) );
  NAND2_X1 U7614 ( .A1(n7397), .A2(n7298), .ZN(n6966) );
  NAND2_X1 U7615 ( .A1(n7370), .A2(REIP_REG_11__SCAN_IN), .ZN(n7393) );
  OAI21_X1 U7616 ( .B1(n7283), .B2(n5858), .A(n7393), .ZN(n6963) );
  AOI21_X1 U7617 ( .B1(n7278), .B2(n6964), .A(n6963), .ZN(n6965) );
  OAI211_X1 U7618 ( .C1(n6976), .C2(n6967), .A(n6966), .B(n6965), .ZN(U2975)
         );
  AOI21_X1 U7619 ( .B1(n6970), .B2(n6969), .A(n6968), .ZN(n7377) );
  NAND2_X1 U7620 ( .A1(n7377), .A2(n7298), .ZN(n6974) );
  AND2_X1 U7621 ( .A1(n7370), .A2(REIP_REG_10__SCAN_IN), .ZN(n7374) );
  NOR2_X1 U7622 ( .A1(n7302), .A2(n6971), .ZN(n6972) );
  AOI211_X1 U7623 ( .C1(n7296), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n7374), 
        .B(n6972), .ZN(n6973) );
  OAI211_X1 U7624 ( .C1(n6976), .C2(n6975), .A(n6974), .B(n6973), .ZN(U2976)
         );
  INV_X1 U7625 ( .A(n6977), .ZN(n6987) );
  NAND3_X1 U7626 ( .A1(n6978), .A2(n6834), .A3(n7419), .ZN(n6985) );
  INV_X1 U7627 ( .A(n6979), .ZN(n6983) );
  OAI21_X1 U7628 ( .B1(n6981), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n6980), 
        .ZN(n6982) );
  AOI21_X1 U7629 ( .B1(n6983), .B2(n7418), .A(n6982), .ZN(n6984) );
  OAI211_X1 U7630 ( .C1(n6987), .C2(n6986), .A(n6985), .B(n6984), .ZN(U2991)
         );
  INV_X1 U7631 ( .A(n7006), .ZN(n7001) );
  OAI211_X1 U7632 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A(n6996), .B(n6988), .ZN(n6989) );
  OAI211_X1 U7633 ( .C1(n6991), .C2(n7090), .A(n6990), .B(n6989), .ZN(n6992)
         );
  AOI21_X1 U7634 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n7001), .A(n6992), 
        .ZN(n6993) );
  OAI21_X1 U7635 ( .B1(n6994), .B2(n7350), .A(n6993), .ZN(U2992) );
  NAND2_X1 U7636 ( .A1(n6996), .A2(n6995), .ZN(n6997) );
  OAI211_X1 U7637 ( .C1(n6999), .C2(n7090), .A(n6998), .B(n6997), .ZN(n7000)
         );
  AOI21_X1 U7638 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n7001), .A(n7000), 
        .ZN(n7002) );
  OAI21_X1 U7639 ( .B1(n7003), .B2(n7350), .A(n7002), .ZN(U2993) );
  INV_X1 U7640 ( .A(n7004), .ZN(n7009) );
  AOI21_X1 U7641 ( .B1(n7017), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n7005) );
  NOR2_X1 U7642 ( .A1(n7006), .A2(n7005), .ZN(n7007) );
  AOI211_X1 U7643 ( .C1(n7418), .C2(n7009), .A(n7008), .B(n7007), .ZN(n7010)
         );
  OAI21_X1 U7644 ( .B1(n7011), .B2(n7350), .A(n7010), .ZN(U2994) );
  INV_X1 U7645 ( .A(n7012), .ZN(n7022) );
  XNOR2_X1 U7646 ( .A(n7014), .B(n7013), .ZN(n7536) );
  AOI21_X1 U7647 ( .B1(n7017), .B2(n7016), .A(n7015), .ZN(n7018) );
  OAI21_X1 U7648 ( .B1(n7536), .B2(n7090), .A(n7018), .ZN(n7019) );
  AOI21_X1 U7649 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n7020), .A(n7019), 
        .ZN(n7021) );
  OAI21_X1 U7650 ( .B1(n7022), .B2(n7350), .A(n7021), .ZN(U2995) );
  NOR2_X1 U7651 ( .A1(n7056), .A2(n7023), .ZN(n7037) );
  XNOR2_X1 U7652 ( .A(n7024), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n7025)
         );
  NAND2_X1 U7653 ( .A1(n7037), .A2(n7025), .ZN(n7026) );
  OAI211_X1 U7654 ( .C1(n7028), .C2(n7090), .A(n7027), .B(n7026), .ZN(n7029)
         );
  AOI21_X1 U7655 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n7048), .A(n7029), 
        .ZN(n7030) );
  OAI21_X1 U7656 ( .B1(n7031), .B2(n7350), .A(n7030), .ZN(U2996) );
  INV_X1 U7657 ( .A(n7048), .ZN(n7041) );
  NAND3_X1 U7658 ( .A1(n7033), .A2(n7032), .A3(n7419), .ZN(n7039) );
  OAI21_X1 U7659 ( .B1(n7035), .B2(n7090), .A(n7034), .ZN(n7036) );
  AOI21_X1 U7660 ( .B1(n7037), .B2(n7040), .A(n7036), .ZN(n7038) );
  OAI211_X1 U7661 ( .C1(n7041), .C2(n7040), .A(n7039), .B(n7038), .ZN(U2997)
         );
  OAI21_X1 U7662 ( .B1(n7043), .B2(n7090), .A(n7042), .ZN(n7047) );
  NOR2_X1 U7663 ( .A1(n7045), .A2(n7044), .ZN(n7046) );
  AOI211_X1 U7664 ( .C1(INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n7048), .A(n7047), .B(n7046), .ZN(n7049) );
  OAI21_X1 U7665 ( .B1(n7050), .B2(n7350), .A(n7049), .ZN(U2998) );
  OAI21_X1 U7666 ( .B1(n6862), .B2(n7052), .A(n7051), .ZN(n7299) );
  AOI22_X1 U7667 ( .A1(n7520), .A2(n7418), .B1(n7370), .B2(
        REIP_REG_19__SCAN_IN), .ZN(n7055) );
  NAND2_X1 U7668 ( .A1(n7053), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n7054) );
  OAI211_X1 U7669 ( .C1(n7056), .C2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n7055), .B(n7054), .ZN(n7057) );
  AOI21_X1 U7670 ( .B1(n7299), .B2(n7419), .A(n7057), .ZN(n7058) );
  INV_X1 U7671 ( .A(n7058), .ZN(U2999) );
  INV_X1 U7672 ( .A(n7059), .ZN(n7069) );
  OAI21_X1 U7673 ( .B1(n7062), .B2(n7061), .A(n7060), .ZN(n7081) );
  AOI21_X1 U7674 ( .B1(n7063), .B2(n7069), .A(n7081), .ZN(n7064) );
  OAI21_X1 U7675 ( .B1(n7065), .B2(n7079), .A(n7064), .ZN(n7410) );
  INV_X1 U7676 ( .A(n7410), .ZN(n7074) );
  XNOR2_X1 U7677 ( .A(n7066), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n7067)
         );
  XNOR2_X1 U7678 ( .A(n7068), .B(n7067), .ZN(n7292) );
  NAND2_X1 U7679 ( .A1(n7292), .A2(n7419), .ZN(n7072) );
  NOR2_X1 U7680 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n7069), .ZN(n7411)
         );
  OAI22_X1 U7681 ( .A1(n7502), .A2(n7090), .B1(n7088), .B2(n7199), .ZN(n7070)
         );
  AOI21_X1 U7682 ( .B1(n7383), .B2(n7411), .A(n7070), .ZN(n7071) );
  OAI211_X1 U7683 ( .C1(n7074), .C2(n7073), .A(n7072), .B(n7071), .ZN(U3001)
         );
  NOR2_X1 U7684 ( .A1(n7414), .A2(n7400), .ZN(n7085) );
  OAI21_X1 U7685 ( .B1(n7090), .B2(n7076), .A(n7075), .ZN(n7084) );
  INV_X1 U7686 ( .A(n7077), .ZN(n7078) );
  NOR2_X1 U7687 ( .A1(n7079), .A2(n7078), .ZN(n7080) );
  AND2_X1 U7688 ( .A1(n7340), .A2(n7400), .ZN(n7082) );
  NOR2_X1 U7689 ( .A1(n7396), .A2(n7082), .ZN(n7409) );
  NOR2_X1 U7690 ( .A1(n7409), .A2(n7401), .ZN(n7083) );
  AOI211_X1 U7691 ( .C1(n7085), .C2(n7401), .A(n7084), .B(n7083), .ZN(n7086)
         );
  OAI21_X1 U7692 ( .B1(n7087), .B2(n7350), .A(n7086), .ZN(U3003) );
  NOR2_X1 U7693 ( .A1(n7414), .A2(n7385), .ZN(n7093) );
  OAI22_X1 U7694 ( .A1(n7090), .A2(n7089), .B1(n7191), .B2(n7088), .ZN(n7091)
         );
  AOI21_X1 U7695 ( .B1(n7093), .B2(n7092), .A(n7091), .ZN(n7097) );
  INV_X1 U7696 ( .A(n7396), .ZN(n7094) );
  OAI21_X1 U7697 ( .B1(n7095), .B2(n7331), .A(n7094), .ZN(n7328) );
  NAND2_X1 U7698 ( .A1(n7328), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n7096) );
  OAI211_X1 U7699 ( .C1(n7098), .C2(n7350), .A(n7097), .B(n7096), .ZN(U3005)
         );
  INV_X1 U7700 ( .A(n7459), .ZN(n7105) );
  INV_X1 U7701 ( .A(n7099), .ZN(n7104) );
  AOI221_X1 U7702 ( .B1(n7102), .B2(n4111), .C1(n7101), .C2(n4111), .A(n7100), 
        .ZN(n7103) );
  AOI211_X1 U7703 ( .C1(n7418), .C2(n7105), .A(n7104), .B(n7103), .ZN(n7106)
         );
  OAI21_X1 U7704 ( .B1(n7107), .B2(n7350), .A(n7106), .ZN(U3014) );
  INV_X1 U7705 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n7109) );
  NAND2_X1 U7706 ( .A1(STATE_REG_1__SCAN_IN), .A2(n7619), .ZN(n7627) );
  AOI21_X1 U7707 ( .B1(n7621), .B2(STATE_REG_1__SCAN_IN), .A(n7619), .ZN(n7135) );
  INV_X1 U7708 ( .A(n3658), .ZN(n7128) );
  NAND2_X1 U7709 ( .A1(n7621), .A2(n7619), .ZN(n7304) );
  AOI21_X1 U7710 ( .B1(n7108), .B2(n7304), .A(n7128), .ZN(n7607) );
  AOI21_X1 U7711 ( .B1(n7109), .B2(n7128), .A(n7607), .ZN(U3451) );
  NOR2_X1 U7712 ( .A1(n3658), .A2(n7110), .ZN(U3180) );
  AND2_X1 U7713 ( .A1(n7128), .A2(DATAWIDTH_REG_3__SCAN_IN), .ZN(U3179) );
  NOR2_X1 U7714 ( .A1(n3658), .A2(n7111), .ZN(U3178) );
  NOR2_X1 U7715 ( .A1(n3658), .A2(n7112), .ZN(U3177) );
  NOR2_X1 U7716 ( .A1(n3658), .A2(n7113), .ZN(U3176) );
  AND2_X1 U7717 ( .A1(n7128), .A2(DATAWIDTH_REG_7__SCAN_IN), .ZN(U3175) );
  AND2_X1 U7718 ( .A1(n7128), .A2(DATAWIDTH_REG_8__SCAN_IN), .ZN(U3174) );
  INV_X1 U7719 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n7114) );
  NOR2_X1 U7720 ( .A1(n3658), .A2(n7114), .ZN(U3173) );
  INV_X1 U7721 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n7115) );
  NOR2_X1 U7722 ( .A1(n3658), .A2(n7115), .ZN(U3172) );
  INV_X1 U7723 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n7116) );
  NOR2_X1 U7724 ( .A1(n3658), .A2(n7116), .ZN(U3171) );
  INV_X1 U7725 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n7117) );
  NOR2_X1 U7726 ( .A1(n3658), .A2(n7117), .ZN(U3170) );
  INV_X1 U7727 ( .A(DATAWIDTH_REG_13__SCAN_IN), .ZN(n7118) );
  NOR2_X1 U7728 ( .A1(n3658), .A2(n7118), .ZN(U3169) );
  NOR2_X1 U7729 ( .A1(n3658), .A2(n7119), .ZN(U3168) );
  NOR2_X1 U7730 ( .A1(n3658), .A2(n7120), .ZN(U3167) );
  NOR2_X1 U7731 ( .A1(n3658), .A2(n7121), .ZN(U3166) );
  NOR2_X1 U7732 ( .A1(n3658), .A2(n7122), .ZN(U3165) );
  NOR2_X1 U7733 ( .A1(n3658), .A2(n7123), .ZN(U3164) );
  NOR2_X1 U7734 ( .A1(n3658), .A2(n7124), .ZN(U3163) );
  NOR2_X1 U7735 ( .A1(n3658), .A2(n7125), .ZN(U3162) );
  NOR2_X1 U7736 ( .A1(n3658), .A2(n7126), .ZN(U3161) );
  INV_X1 U7737 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n7127) );
  NOR2_X1 U7738 ( .A1(n3658), .A2(n7127), .ZN(U3160) );
  AND2_X1 U7739 ( .A1(n7128), .A2(DATAWIDTH_REG_23__SCAN_IN), .ZN(U3159) );
  AND2_X1 U7740 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n7128), .ZN(U3158) );
  AND2_X1 U7741 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n7128), .ZN(U3157) );
  AND2_X1 U7742 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n7128), .ZN(U3156) );
  AND2_X1 U7743 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n7128), .ZN(U3155) );
  AND2_X1 U7744 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n7128), .ZN(U3154) );
  AND2_X1 U7745 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n7128), .ZN(U3153) );
  AND2_X1 U7746 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n7128), .ZN(U3152) );
  AND2_X1 U7747 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n7128), .ZN(U3151) );
  NOR2_X1 U7748 ( .A1(n7130), .A2(n7129), .ZN(U3019) );
  INV_X2 U7749 ( .A(n7322), .ZN(n7580) );
  AOI21_X1 U7750 ( .B1(n7132), .B2(n7554), .A(n7131), .ZN(n7133) );
  AND2_X1 U7751 ( .A1(n7164), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U7752 ( .A(ADS_N_REG_SCAN_IN), .ZN(n7134) );
  AOI21_X1 U7753 ( .B1(n7135), .B2(n7134), .A(n7309), .ZN(U2789) );
  AOI22_X1 U7754 ( .A1(n7580), .A2(LWORD_REG_0__SCAN_IN), .B1(n7169), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n7136) );
  OAI21_X1 U7755 ( .B1(n7638), .B2(n7152), .A(n7136), .ZN(U2923) );
  AOI22_X1 U7756 ( .A1(n7580), .A2(LWORD_REG_1__SCAN_IN), .B1(n7169), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n7137) );
  OAI21_X1 U7757 ( .B1(n7641), .B2(n7152), .A(n7137), .ZN(U2922) );
  AOI22_X1 U7758 ( .A1(n7580), .A2(LWORD_REG_2__SCAN_IN), .B1(n7169), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n7138) );
  OAI21_X1 U7759 ( .B1(n7645), .B2(n7152), .A(n7138), .ZN(U2921) );
  AOI22_X1 U7760 ( .A1(n7580), .A2(LWORD_REG_3__SCAN_IN), .B1(n7164), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n7139) );
  OAI21_X1 U7761 ( .B1(n7648), .B2(n7152), .A(n7139), .ZN(U2920) );
  AOI22_X1 U7762 ( .A1(n7580), .A2(LWORD_REG_4__SCAN_IN), .B1(n7169), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n7140) );
  OAI21_X1 U7763 ( .B1(n7652), .B2(n7152), .A(n7140), .ZN(U2919) );
  AOI22_X1 U7764 ( .A1(n7580), .A2(LWORD_REG_5__SCAN_IN), .B1(n7164), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n7141) );
  OAI21_X1 U7765 ( .B1(n7656), .B2(n7152), .A(n7141), .ZN(U2918) );
  AOI22_X1 U7766 ( .A1(n7580), .A2(LWORD_REG_6__SCAN_IN), .B1(n7169), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n7142) );
  OAI21_X1 U7767 ( .B1(n7660), .B2(n7152), .A(n7142), .ZN(U2917) );
  AOI22_X1 U7768 ( .A1(n7580), .A2(LWORD_REG_7__SCAN_IN), .B1(n7169), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n7143) );
  OAI21_X1 U7769 ( .B1(n4304), .B2(n7152), .A(n7143), .ZN(U2916) );
  AOI22_X1 U7770 ( .A1(n7580), .A2(LWORD_REG_8__SCAN_IN), .B1(n7169), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n7144) );
  OAI21_X1 U7771 ( .B1(n7668), .B2(n7152), .A(n7144), .ZN(U2915) );
  AOI22_X1 U7772 ( .A1(n7580), .A2(LWORD_REG_9__SCAN_IN), .B1(n7169), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n7145) );
  OAI21_X1 U7773 ( .B1(n7672), .B2(n7152), .A(n7145), .ZN(U2914) );
  AOI22_X1 U7774 ( .A1(n7580), .A2(LWORD_REG_10__SCAN_IN), .B1(n7169), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n7146) );
  OAI21_X1 U7775 ( .B1(n7676), .B2(n7152), .A(n7146), .ZN(U2913) );
  AOI22_X1 U7776 ( .A1(n7580), .A2(LWORD_REG_11__SCAN_IN), .B1(n7169), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n7147) );
  OAI21_X1 U7777 ( .B1(n7679), .B2(n7152), .A(n7147), .ZN(U2912) );
  AOI22_X1 U7778 ( .A1(n7580), .A2(LWORD_REG_12__SCAN_IN), .B1(n7169), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n7148) );
  OAI21_X1 U7779 ( .B1(n7683), .B2(n7152), .A(n7148), .ZN(U2911) );
  AOI22_X1 U7780 ( .A1(n7580), .A2(LWORD_REG_13__SCAN_IN), .B1(n7169), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n7149) );
  OAI21_X1 U7781 ( .B1(n7686), .B2(n7152), .A(n7149), .ZN(U2910) );
  AOI22_X1 U7782 ( .A1(n7580), .A2(LWORD_REG_14__SCAN_IN), .B1(n7169), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n7150) );
  OAI21_X1 U7783 ( .B1(n7690), .B2(n7152), .A(n7150), .ZN(U2909) );
  AOI22_X1 U7784 ( .A1(n7580), .A2(LWORD_REG_15__SCAN_IN), .B1(n7169), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n7151) );
  OAI21_X1 U7785 ( .B1(n7695), .B2(n7152), .A(n7151), .ZN(U2908) );
  INV_X1 U7786 ( .A(EAX_REG_16__SCAN_IN), .ZN(n7636) );
  AOI22_X1 U7787 ( .A1(n7580), .A2(UWORD_REG_0__SCAN_IN), .B1(n7169), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n7154) );
  OAI21_X1 U7788 ( .B1(n7636), .B2(n7171), .A(n7154), .ZN(U2907) );
  AOI22_X1 U7789 ( .A1(n7580), .A2(UWORD_REG_1__SCAN_IN), .B1(n7169), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n7155) );
  OAI21_X1 U7790 ( .B1(n4476), .B2(n7171), .A(n7155), .ZN(U2906) );
  INV_X1 U7791 ( .A(EAX_REG_18__SCAN_IN), .ZN(n7643) );
  AOI22_X1 U7792 ( .A1(n7580), .A2(UWORD_REG_2__SCAN_IN), .B1(n7169), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n7156) );
  OAI21_X1 U7793 ( .B1(n7643), .B2(n7171), .A(n7156), .ZN(U2905) );
  AOI22_X1 U7794 ( .A1(n7580), .A2(UWORD_REG_3__SCAN_IN), .B1(n7164), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n7157) );
  OAI21_X1 U7795 ( .B1(n4511), .B2(n7171), .A(n7157), .ZN(U2904) );
  INV_X1 U7796 ( .A(EAX_REG_20__SCAN_IN), .ZN(n7650) );
  AOI22_X1 U7797 ( .A1(n7580), .A2(UWORD_REG_4__SCAN_IN), .B1(n7164), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n7158) );
  OAI21_X1 U7798 ( .B1(n7650), .B2(n7171), .A(n7158), .ZN(U2903) );
  INV_X1 U7799 ( .A(EAX_REG_21__SCAN_IN), .ZN(n7654) );
  AOI22_X1 U7800 ( .A1(n7580), .A2(UWORD_REG_5__SCAN_IN), .B1(n7164), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n7159) );
  OAI21_X1 U7801 ( .B1(n7654), .B2(n7171), .A(n7159), .ZN(U2902) );
  INV_X1 U7802 ( .A(EAX_REG_22__SCAN_IN), .ZN(n7658) );
  AOI22_X1 U7803 ( .A1(n7580), .A2(UWORD_REG_6__SCAN_IN), .B1(n7164), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n7160) );
  OAI21_X1 U7804 ( .B1(n7658), .B2(n7171), .A(n7160), .ZN(U2901) );
  INV_X1 U7805 ( .A(EAX_REG_23__SCAN_IN), .ZN(n7662) );
  AOI22_X1 U7806 ( .A1(n7580), .A2(UWORD_REG_7__SCAN_IN), .B1(n7164), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n7161) );
  OAI21_X1 U7807 ( .B1(n7662), .B2(n7171), .A(n7161), .ZN(U2900) );
  INV_X1 U7808 ( .A(EAX_REG_24__SCAN_IN), .ZN(n7665) );
  AOI22_X1 U7809 ( .A1(n7580), .A2(UWORD_REG_8__SCAN_IN), .B1(n7164), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n7162) );
  OAI21_X1 U7810 ( .B1(n7665), .B2(n7171), .A(n7162), .ZN(U2899) );
  INV_X1 U7811 ( .A(EAX_REG_25__SCAN_IN), .ZN(n7670) );
  AOI22_X1 U7812 ( .A1(n7580), .A2(UWORD_REG_9__SCAN_IN), .B1(n7164), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n7163) );
  OAI21_X1 U7813 ( .B1(n7670), .B2(n7171), .A(n7163), .ZN(U2898) );
  INV_X1 U7814 ( .A(EAX_REG_26__SCAN_IN), .ZN(n7674) );
  AOI22_X1 U7815 ( .A1(n7580), .A2(UWORD_REG_10__SCAN_IN), .B1(n7164), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n7165) );
  OAI21_X1 U7816 ( .B1(n7674), .B2(n7171), .A(n7165), .ZN(U2897) );
  AOI22_X1 U7817 ( .A1(n7580), .A2(UWORD_REG_11__SCAN_IN), .B1(n7169), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n7166) );
  OAI21_X1 U7818 ( .B1(n4669), .B2(n7171), .A(n7166), .ZN(U2896) );
  INV_X1 U7819 ( .A(EAX_REG_28__SCAN_IN), .ZN(n7681) );
  AOI22_X1 U7820 ( .A1(n7580), .A2(UWORD_REG_12__SCAN_IN), .B1(n7169), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n7167) );
  OAI21_X1 U7821 ( .B1(n7681), .B2(n7171), .A(n7167), .ZN(U2895) );
  AOI22_X1 U7822 ( .A1(n7580), .A2(UWORD_REG_13__SCAN_IN), .B1(n7169), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n7168) );
  OAI21_X1 U7823 ( .B1(n4712), .B2(n7171), .A(n7168), .ZN(U2894) );
  INV_X1 U7824 ( .A(EAX_REG_30__SCAN_IN), .ZN(n7688) );
  AOI22_X1 U7825 ( .A1(n7580), .A2(UWORD_REG_14__SCAN_IN), .B1(n7169), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n7170) );
  OAI21_X1 U7826 ( .B1(n7688), .B2(n7171), .A(n7170), .ZN(U2893) );
  NAND2_X1 U7827 ( .A1(n7309), .A2(n7621), .ZN(n7230) );
  INV_X1 U7828 ( .A(REIP_REG_1__SCAN_IN), .ZN(n7435) );
  NAND2_X1 U7829 ( .A1(STATE_REG_2__SCAN_IN), .A2(n7309), .ZN(n7218) );
  CLKBUF_X1 U7830 ( .A(n7218), .Z(n7226) );
  OAI222_X1 U7831 ( .A1(n7219), .A2(n7434), .B1(n7172), .B2(n7309), .C1(n7435), 
        .C2(n7226), .ZN(U3184) );
  INV_X1 U7832 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n7173) );
  OAI222_X1 U7833 ( .A1(n7230), .A2(n7174), .B1(n7173), .B2(n7309), .C1(n7434), 
        .C2(n7218), .ZN(U3185) );
  INV_X1 U7834 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n7175) );
  OAI222_X1 U7835 ( .A1(n7230), .A2(n7453), .B1(n7175), .B2(n7309), .C1(n7174), 
        .C2(n7226), .ZN(U3186) );
  INV_X1 U7836 ( .A(REIP_REG_5__SCAN_IN), .ZN(n7177) );
  INV_X1 U7837 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n7176) );
  OAI222_X1 U7838 ( .A1(n7230), .A2(n7177), .B1(n7176), .B2(n7309), .C1(n7453), 
        .C2(n7226), .ZN(U3187) );
  OAI222_X1 U7839 ( .A1(n7230), .A2(n6442), .B1(n7178), .B2(n7309), .C1(n7177), 
        .C2(n7226), .ZN(U3188) );
  INV_X1 U7840 ( .A(REIP_REG_7__SCAN_IN), .ZN(n7494) );
  INV_X1 U7841 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n7179) );
  OAI222_X1 U7842 ( .A1(n7230), .A2(n7494), .B1(n7179), .B2(n7309), .C1(n6442), 
        .C2(n7226), .ZN(U3189) );
  OAI222_X1 U7843 ( .A1(n7219), .A2(n7181), .B1(n7180), .B2(n7309), .C1(n7494), 
        .C2(n7218), .ZN(U3190) );
  INV_X1 U7844 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n7182) );
  OAI222_X1 U7845 ( .A1(n7219), .A2(n7184), .B1(n7182), .B2(n7309), .C1(n7181), 
        .C2(n7226), .ZN(U3191) );
  INV_X1 U7846 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n7183) );
  INV_X1 U7847 ( .A(REIP_REG_10__SCAN_IN), .ZN(n7185) );
  OAI222_X1 U7848 ( .A1(n7226), .A2(n7184), .B1(n7183), .B2(n7309), .C1(n7185), 
        .C2(n7219), .ZN(U3192) );
  OAI222_X1 U7849 ( .A1(n7219), .A2(n7188), .B1(n7186), .B2(n7309), .C1(n7185), 
        .C2(n7218), .ZN(U3193) );
  INV_X1 U7850 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n7187) );
  OAI222_X1 U7851 ( .A1(n7226), .A2(n7188), .B1(n7187), .B2(n7309), .C1(n7190), 
        .C2(n7219), .ZN(U3194) );
  OAI222_X1 U7852 ( .A1(n7218), .A2(n7190), .B1(n7189), .B2(n7309), .C1(n7191), 
        .C2(n7219), .ZN(U3195) );
  INV_X1 U7853 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n7192) );
  OAI222_X1 U7854 ( .A1(n7219), .A2(n7193), .B1(n7192), .B2(n7309), .C1(n7191), 
        .C2(n7226), .ZN(U3196) );
  OAI222_X1 U7855 ( .A1(n7219), .A2(n7196), .B1(n7194), .B2(n7309), .C1(n7193), 
        .C2(n7226), .ZN(U3197) );
  OAI222_X1 U7856 ( .A1(n7218), .A2(n7196), .B1(n7195), .B2(n7309), .C1(n7198), 
        .C2(n7219), .ZN(U3198) );
  INV_X1 U7857 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n7197) );
  OAI222_X1 U7858 ( .A1(n7218), .A2(n7198), .B1(n7197), .B2(n7309), .C1(n7199), 
        .C2(n7219), .ZN(U3199) );
  INV_X1 U7859 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n7200) );
  OAI222_X1 U7860 ( .A1(n7219), .A2(n7201), .B1(n7200), .B2(n7309), .C1(n7199), 
        .C2(n7226), .ZN(U3200) );
  OAI222_X1 U7861 ( .A1(n7230), .A2(n7203), .B1(n7202), .B2(n7309), .C1(n7201), 
        .C2(n7226), .ZN(U3201) );
  INV_X1 U7862 ( .A(REIP_REG_20__SCAN_IN), .ZN(n7206) );
  INV_X1 U7863 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n7204) );
  OAI222_X1 U7864 ( .A1(n7230), .A2(n7206), .B1(n7204), .B2(n7309), .C1(n7203), 
        .C2(n7226), .ZN(U3202) );
  OAI222_X1 U7865 ( .A1(n7218), .A2(n7206), .B1(n7205), .B2(n7309), .C1(n7207), 
        .C2(n7219), .ZN(U3203) );
  INV_X1 U7866 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n7208) );
  OAI222_X1 U7867 ( .A1(n7230), .A2(n7210), .B1(n7208), .B2(n7309), .C1(n7207), 
        .C2(n7226), .ZN(U3204) );
  INV_X1 U7868 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n7209) );
  OAI222_X1 U7869 ( .A1(n7218), .A2(n7210), .B1(n7209), .B2(n7309), .C1(n7526), 
        .C2(n7219), .ZN(U3205) );
  INV_X1 U7870 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n7211) );
  OAI222_X1 U7871 ( .A1(n7218), .A2(n7526), .B1(n7211), .B2(n7309), .C1(n7212), 
        .C2(n7219), .ZN(U3206) );
  INV_X1 U7872 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n7213) );
  OAI222_X1 U7873 ( .A1(n7230), .A2(n7214), .B1(n7213), .B2(n7309), .C1(n7212), 
        .C2(n7226), .ZN(U3207) );
  INV_X1 U7874 ( .A(REIP_REG_26__SCAN_IN), .ZN(n7217) );
  OAI222_X1 U7875 ( .A1(n7219), .A2(n7217), .B1(n7215), .B2(n7309), .C1(n7214), 
        .C2(n7226), .ZN(U3208) );
  INV_X1 U7876 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n7216) );
  OAI222_X1 U7877 ( .A1(n7218), .A2(n7217), .B1(n7216), .B2(n7309), .C1(n7221), 
        .C2(n7219), .ZN(U3209) );
  OAI222_X1 U7878 ( .A1(n7226), .A2(n7221), .B1(n7220), .B2(n7309), .C1(n7222), 
        .C2(n7219), .ZN(U3210) );
  INV_X1 U7879 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n7223) );
  OAI222_X1 U7880 ( .A1(n7230), .A2(n7224), .B1(n7223), .B2(n7309), .C1(n7222), 
        .C2(n7226), .ZN(U3211) );
  OAI222_X1 U7881 ( .A1(n7230), .A2(n7227), .B1(n7225), .B2(n7309), .C1(n7224), 
        .C2(n7226), .ZN(U3212) );
  OAI222_X1 U7882 ( .A1(n7230), .A2(n7229), .B1(n7228), .B2(n7309), .C1(n7227), 
        .C2(n7226), .ZN(U3213) );
  AOI22_X1 U7883 ( .A1(n7309), .A2(n7232), .B1(n7231), .B2(n7627), .ZN(U3445)
         );
  AOI221_X1 U7884 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(REIP_REG_1__SCAN_IN), 
        .C1(REIP_REG_0__SCAN_IN), .C2(REIP_REG_1__SCAN_IN), .A(
        DATAWIDTH_REG_1__SCAN_IN), .ZN(n7243) );
  NOR4_X1 U7885 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(
        DATAWIDTH_REG_30__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_28__SCAN_IN), .ZN(n7236) );
  NOR4_X1 U7886 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n7235) );
  NOR4_X1 U7887 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(DATAWIDTH_REG_3__SCAN_IN), 
        .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_23__SCAN_IN), .ZN(
        n7234) );
  NOR4_X1 U7888 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_26__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_24__SCAN_IN), .ZN(n7233) );
  NAND4_X1 U7889 ( .A1(n7236), .A2(n7235), .A3(n7234), .A4(n7233), .ZN(n7242)
         );
  NOR4_X1 U7890 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), .A3(DATAWIDTH_REG_5__SCAN_IN), .A4(DATAWIDTH_REG_9__SCAN_IN), .ZN(n7240) );
  AOI211_X1 U7891 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_2__SCAN_IN), .B(
        DATAWIDTH_REG_4__SCAN_IN), .ZN(n7239) );
  NOR4_X1 U7892 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_17__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n7238) );
  NOR4_X1 U7893 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n7237) );
  NAND4_X1 U7894 ( .A1(n7240), .A2(n7239), .A3(n7238), .A4(n7237), .ZN(n7241)
         );
  NOR2_X1 U7895 ( .A1(n7242), .A2(n7241), .ZN(n7255) );
  MUX2_X1 U7896 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(n7243), .S(n7255), .Z(
        U2795) );
  INV_X1 U7897 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n7247) );
  INV_X1 U7898 ( .A(BE_N_REG_2__SCAN_IN), .ZN(n7244) );
  AOI22_X1 U7899 ( .A1(n7309), .A2(n7247), .B1(n7244), .B2(n7627), .ZN(U3446)
         );
  AOI21_X1 U7900 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7245) );
  OAI221_X1 U7901 ( .B1(REIP_REG_1__SCAN_IN), .B2(n7245), .C1(n7435), .C2(
        REIP_REG_0__SCAN_IN), .A(n7255), .ZN(n7246) );
  OAI21_X1 U7902 ( .B1(n7255), .B2(n7247), .A(n7246), .ZN(U3468) );
  INV_X1 U7903 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n7251) );
  AOI22_X1 U7904 ( .A1(n7309), .A2(n7251), .B1(n7248), .B2(n7627), .ZN(U3447)
         );
  NOR3_X1 U7905 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(REIP_REG_0__SCAN_IN), .ZN(n7249) );
  OAI21_X1 U7906 ( .B1(REIP_REG_1__SCAN_IN), .B2(n7249), .A(n7255), .ZN(n7250)
         );
  OAI21_X1 U7907 ( .B1(n7255), .B2(n7251), .A(n7250), .ZN(U2794) );
  INV_X1 U7908 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n7254) );
  INV_X1 U7909 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n7252) );
  AOI22_X1 U7910 ( .A1(n7309), .A2(n7254), .B1(n7252), .B2(n7627), .ZN(U3448)
         );
  OAI21_X1 U7911 ( .B1(REIP_REG_0__SCAN_IN), .B2(REIP_REG_1__SCAN_IN), .A(
        n7255), .ZN(n7253) );
  OAI21_X1 U7912 ( .B1(n7255), .B2(n7254), .A(n7253), .ZN(U3469) );
  OAI22_X1 U7913 ( .A1(n7705), .A2(n7256), .B1(n7536), .B2(n3659), .ZN(n7257)
         );
  INV_X1 U7914 ( .A(n7257), .ZN(n7258) );
  OAI21_X1 U7915 ( .B1(n7259), .B2(n7530), .A(n7258), .ZN(U2836) );
  AOI22_X1 U7916 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n7296), .B1(n7370), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n7266) );
  NAND2_X1 U7917 ( .A1(n7261), .A2(n7260), .ZN(n7262) );
  XOR2_X1 U7918 ( .A(n7263), .B(n7262), .Z(n7339) );
  AOI22_X1 U7919 ( .A1(n7339), .A2(n7298), .B1(n7297), .B2(n7264), .ZN(n7265)
         );
  OAI211_X1 U7920 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n7302), .A(n7266), 
        .B(n7265), .ZN(U2985) );
  AOI22_X1 U7921 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n7296), .B1(n7370), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n7274) );
  NAND2_X1 U7922 ( .A1(n7268), .A2(n7267), .ZN(n7270) );
  XNOR2_X1 U7923 ( .A(n7270), .B(n7269), .ZN(n7351) );
  INV_X1 U7924 ( .A(n7351), .ZN(n7272) );
  AOI22_X1 U7925 ( .A1(n7272), .A2(n7298), .B1(n7271), .B2(n7297), .ZN(n7273)
         );
  OAI211_X1 U7926 ( .C1(n7302), .C2(n7275), .A(n7274), .B(n7273), .ZN(U2984)
         );
  INV_X1 U7927 ( .A(n7276), .ZN(n7279) );
  INV_X1 U7928 ( .A(n7277), .ZN(n7473) );
  AOI222_X1 U7929 ( .A1(n7279), .A2(n7298), .B1(n7297), .B2(n7475), .C1(n7473), 
        .C2(n7278), .ZN(n7281) );
  OAI211_X1 U7930 ( .C1(n7283), .C2(n7282), .A(n7281), .B(n7280), .ZN(U2981)
         );
  AOI22_X1 U7931 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n7296), .B1(n7370), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n7287) );
  INV_X1 U7932 ( .A(n7284), .ZN(n7285) );
  AOI22_X1 U7933 ( .A1(n7285), .A2(n7298), .B1(n7297), .B2(n7484), .ZN(n7286)
         );
  OAI211_X1 U7934 ( .C1(n7302), .C2(n7486), .A(n7287), .B(n7286), .ZN(U2980)
         );
  AOI22_X1 U7935 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n7296), .B1(n7370), 
        .B2(REIP_REG_7__SCAN_IN), .ZN(n7291) );
  AOI21_X1 U7936 ( .B1(n7289), .B2(n7288), .A(n3744), .ZN(n7368) );
  AOI22_X1 U7937 ( .A1(n7368), .A2(n7298), .B1(n7297), .B2(n7498), .ZN(n7290)
         );
  OAI211_X1 U7938 ( .C1(n7302), .C2(n7500), .A(n7291), .B(n7290), .ZN(U2979)
         );
  AOI22_X1 U7939 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n7296), .B1(n7370), 
        .B2(REIP_REG_17__SCAN_IN), .ZN(n7294) );
  AOI22_X1 U7940 ( .A1(n7292), .A2(n7298), .B1(n7297), .B2(n7696), .ZN(n7293)
         );
  OAI211_X1 U7941 ( .C1(n7302), .C2(n7295), .A(n7294), .B(n7293), .ZN(U2969)
         );
  AOI22_X1 U7942 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n7296), .B1(n7370), 
        .B2(REIP_REG_19__SCAN_IN), .ZN(n7301) );
  AOI22_X1 U7943 ( .A1(n7299), .A2(n7298), .B1(n7297), .B2(n7699), .ZN(n7300)
         );
  OAI211_X1 U7944 ( .C1(n7302), .C2(n7525), .A(n7301), .B(n7300), .ZN(U2967)
         );
  OAI222_X1 U7945 ( .A1(n7309), .A2(n7304), .B1(n7309), .B2(n7303), .C1(
        CODEFETCH_REG_SCAN_IN), .C2(n7627), .ZN(U2791) );
  OAI21_X1 U7946 ( .B1(n7305), .B2(READREQUEST_REG_SCAN_IN), .A(n7320), .ZN(
        n7306) );
  OAI21_X1 U7947 ( .B1(n7320), .B2(n7307), .A(n7306), .ZN(U3474) );
  AOI22_X1 U7948 ( .A1(n7309), .A2(READREQUEST_REG_SCAN_IN), .B1(n7308), .B2(
        n7627), .ZN(U3470) );
  NOR2_X1 U7949 ( .A1(n7621), .A2(n7310), .ZN(n7612) );
  NAND2_X1 U7950 ( .A1(STATE_REG_0__SCAN_IN), .A2(REQUESTPENDING_REG_SCAN_IN), 
        .ZN(n7622) );
  NAND2_X1 U7951 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n7618) );
  AOI21_X1 U7952 ( .B1(READY_N), .B2(STATE_REG_1__SCAN_IN), .A(n7311), .ZN(
        n7312) );
  OAI221_X1 U7953 ( .B1(n7612), .B2(n7622), .C1(n7612), .C2(n7618), .A(n7312), 
        .ZN(U3182) );
  NAND2_X1 U7954 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .ZN(n7591) );
  OAI21_X1 U7955 ( .B1(n7591), .B2(READY_N), .A(n7584), .ZN(n7313) );
  INV_X1 U7956 ( .A(n7313), .ZN(n7315) );
  OAI21_X1 U7957 ( .B1(n7592), .B2(n7315), .A(n7314), .ZN(U3150) );
  INV_X1 U7958 ( .A(n7316), .ZN(n7317) );
  AOI211_X1 U7959 ( .C1(n4054), .C2(n7608), .A(n7584), .B(n7317), .ZN(n7319)
         );
  OAI21_X1 U7960 ( .B1(n7319), .B2(n7318), .A(n7596), .ZN(n7324) );
  OAI211_X1 U7961 ( .C1(READY_N), .C2(n7322), .A(n7321), .B(n7320), .ZN(n7323)
         );
  MUX2_X1 U7962 ( .A(REQUESTPENDING_REG_SCAN_IN), .B(n7324), .S(n7323), .Z(
        U3472) );
  INV_X1 U7963 ( .A(n7325), .ZN(n7327) );
  AOI21_X1 U7964 ( .B1(n7418), .B2(n7327), .A(n7326), .ZN(n7334) );
  AOI22_X1 U7965 ( .A1(n7329), .A2(n7419), .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n7328), .ZN(n7333) );
  NAND3_X1 U7966 ( .A1(n7331), .A2(n7330), .A3(n7383), .ZN(n7332) );
  NAND3_X1 U7967 ( .A1(n7334), .A2(n7333), .A3(n7332), .ZN(U3004) );
  AOI22_X1 U7968 ( .A1(n7418), .A2(n7335), .B1(n7370), .B2(REIP_REG_1__SCAN_IN), .ZN(n7344) );
  OAI21_X1 U7969 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n7337), .A(n7336), 
        .ZN(n7338) );
  AOI22_X1 U7970 ( .A1(n7419), .A2(n7339), .B1(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .B2(n7338), .ZN(n7343) );
  NAND3_X1 U7971 ( .A1(n4078), .A2(n7341), .A3(n7340), .ZN(n7342) );
  NAND3_X1 U7972 ( .A1(n7344), .A2(n7343), .A3(n7342), .ZN(U3017) );
  NAND2_X1 U7973 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n7346) );
  OAI21_X1 U7974 ( .B1(n7349), .B2(n7346), .A(n7345), .ZN(n7348) );
  AOI222_X1 U7975 ( .A1(n7348), .A2(n7386), .B1(n7418), .B2(n7347), .C1(
        REIP_REG_2__SCAN_IN), .C2(n7370), .ZN(n7356) );
  NAND2_X1 U7976 ( .A1(n7349), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n7352)
         );
  OAI22_X1 U7977 ( .A1(n7353), .A2(n7352), .B1(n7351), .B2(n7350), .ZN(n7354)
         );
  INV_X1 U7978 ( .A(n7354), .ZN(n7355) );
  OAI211_X1 U7979 ( .C1(n7357), .C2(n7349), .A(n7356), .B(n7355), .ZN(U3016)
         );
  AOI21_X1 U7980 ( .B1(n7386), .B2(n7359), .A(n7358), .ZN(n7372) );
  INV_X1 U7981 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n7367) );
  AOI21_X1 U7982 ( .B1(n7418), .B2(n7361), .A(n7360), .ZN(n7366) );
  AOI21_X1 U7983 ( .B1(n7367), .B2(n4809), .A(n7373), .ZN(n7363) );
  AOI22_X1 U7984 ( .A1(n7364), .A2(n7419), .B1(n7363), .B2(n7362), .ZN(n7365)
         );
  OAI211_X1 U7985 ( .C1(n7372), .C2(n7367), .A(n7366), .B(n7365), .ZN(U3010)
         );
  AOI222_X1 U7986 ( .A1(REIP_REG_7__SCAN_IN), .A2(n7370), .B1(n7418), .B2(
        n7369), .C1(n7419), .C2(n7368), .ZN(n7371) );
  OAI221_X1 U7987 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n7373), .C1(n4809), .C2(n7372), .A(n7371), .ZN(U3011) );
  AOI21_X1 U7988 ( .B1(n7418), .B2(n7375), .A(n7374), .ZN(n7382) );
  AOI22_X1 U7989 ( .A1(n7377), .A2(n7419), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n7376), .ZN(n7381) );
  OAI211_X1 U7990 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A(n7379), .B(n7378), .ZN(n7380) );
  NAND3_X1 U7991 ( .A1(n7382), .A2(n7381), .A3(n7380), .ZN(U3008) );
  AOI21_X1 U7992 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n7383), .A(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n7392) );
  INV_X1 U7993 ( .A(n7384), .ZN(n7412) );
  AOI221_X1 U7994 ( .B1(n7386), .B2(n7385), .C1(n7412), .C2(n7385), .A(n7396), 
        .ZN(n7391) );
  AOI22_X1 U7995 ( .A1(n7388), .A2(n7419), .B1(n7418), .B2(n7387), .ZN(n7390)
         );
  NAND2_X1 U7996 ( .A1(n7370), .A2(REIP_REG_12__SCAN_IN), .ZN(n7389) );
  OAI211_X1 U7997 ( .C1(n7392), .C2(n7391), .A(n7390), .B(n7389), .ZN(U3006)
         );
  INV_X1 U7998 ( .A(n7393), .ZN(n7394) );
  AOI21_X1 U7999 ( .B1(n7418), .B2(n7395), .A(n7394), .ZN(n7399) );
  AOI22_X1 U8000 ( .A1(n7397), .A2(n7419), .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n7396), .ZN(n7398) );
  OAI211_X1 U8001 ( .C1(INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n7414), .A(n7399), .B(n7398), .ZN(U3007) );
  AOI211_X1 U8002 ( .C1(n7408), .C2(n7401), .A(n7414), .B(n7400), .ZN(n7403)
         );
  NAND2_X1 U8003 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n7402) );
  AOI22_X1 U8004 ( .A1(n7370), .A2(REIP_REG_16__SCAN_IN), .B1(n7403), .B2(
        n7402), .ZN(n7407) );
  AOI22_X1 U8005 ( .A1(n7405), .A2(n7419), .B1(n7418), .B2(n7404), .ZN(n7406)
         );
  OAI211_X1 U8006 ( .C1(n7409), .C2(n7408), .A(n7407), .B(n7406), .ZN(U3002)
         );
  AOI21_X1 U8007 ( .B1(n7412), .B2(n7411), .A(n7410), .ZN(n7424) );
  NOR3_X1 U8008 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n7414), .A3(n7413), 
        .ZN(n7415) );
  AOI21_X1 U8009 ( .B1(REIP_REG_18__SCAN_IN), .B2(n7370), .A(n7415), .ZN(n7422) );
  INV_X1 U8010 ( .A(n7416), .ZN(n7420) );
  AOI22_X1 U8011 ( .A1(n7420), .A2(n7419), .B1(n7418), .B2(n7417), .ZN(n7421)
         );
  OAI211_X1 U8012 ( .C1(n7424), .C2(n7423), .A(n7422), .B(n7421), .ZN(U3000)
         );
  INV_X1 U8013 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n7433) );
  OAI22_X1 U8014 ( .A1(n7535), .A2(n7426), .B1(n7425), .B2(n7452), .ZN(n7427)
         );
  AOI21_X1 U8015 ( .B1(n7519), .B2(EBX_REG_0__SCAN_IN), .A(n7427), .ZN(n7428)
         );
  OAI21_X1 U8016 ( .B1(n7429), .B2(n4999), .A(n7428), .ZN(n7430) );
  AOI21_X1 U8017 ( .B1(n7431), .B2(n7474), .A(n7430), .ZN(n7432) );
  OAI221_X1 U8018 ( .B1(n7433), .B2(n7531), .C1(n7433), .C2(n7541), .A(n7432), 
        .ZN(U2827) );
  NOR2_X1 U8019 ( .A1(n7435), .A2(n7434), .ZN(n7437) );
  AOI21_X1 U8020 ( .B1(n7437), .B2(n7436), .A(REIP_REG_3__SCAN_IN), .ZN(n7445)
         );
  AOI21_X1 U8021 ( .B1(n7468), .B2(n7456), .A(n7466), .ZN(n7454) );
  OAI22_X1 U8022 ( .A1(n7439), .A2(n7529), .B1(n7452), .B2(n7438), .ZN(n7440)
         );
  INV_X1 U8023 ( .A(n7440), .ZN(n7444) );
  INV_X1 U8024 ( .A(n7441), .ZN(n7442) );
  AOI22_X1 U8025 ( .A1(n7521), .A2(n7442), .B1(PHYADDRPOINTER_REG_3__SCAN_IN), 
        .B2(n7501), .ZN(n7443) );
  OAI211_X1 U8026 ( .C1(n7445), .C2(n7454), .A(n7444), .B(n7443), .ZN(n7446)
         );
  INV_X1 U8027 ( .A(n7446), .ZN(n7451) );
  INV_X1 U8028 ( .A(n7447), .ZN(n7448) );
  AOI22_X1 U8029 ( .A1(n7449), .A2(n7474), .B1(n7504), .B2(n7448), .ZN(n7450)
         );
  NAND2_X1 U8030 ( .A1(n7451), .A2(n7450), .ZN(U2824) );
  OAI22_X1 U8031 ( .A1(n7454), .A2(n7453), .B1(n7545), .B2(n7452), .ZN(n7455)
         );
  AOI211_X1 U8032 ( .C1(n7501), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n7487), 
        .B(n7455), .ZN(n7464) );
  NOR3_X1 U8033 ( .A1(n7457), .A2(REIP_REG_4__SCAN_IN), .A3(n7456), .ZN(n7461)
         );
  OAI22_X1 U8034 ( .A1(n7535), .A2(n7459), .B1(n7529), .B2(n7458), .ZN(n7460)
         );
  AOI211_X1 U8035 ( .C1(n7474), .C2(n7462), .A(n7461), .B(n7460), .ZN(n7463)
         );
  OAI211_X1 U8036 ( .C1(n7465), .C2(n7541), .A(n7464), .B(n7463), .ZN(U2823)
         );
  AOI21_X1 U8037 ( .B1(n7468), .B2(n7467), .A(n7466), .ZN(n7495) );
  AOI21_X1 U8038 ( .B1(n7469), .B2(n7468), .A(REIP_REG_5__SCAN_IN), .ZN(n7478)
         );
  OAI22_X1 U8039 ( .A1(n7535), .A2(n7471), .B1(n7470), .B2(n7529), .ZN(n7472)
         );
  AOI211_X1 U8040 ( .C1(n7501), .C2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n7487), 
        .B(n7472), .ZN(n7477) );
  AOI22_X1 U8041 ( .A1(n7475), .A2(n7474), .B1(n7504), .B2(n7473), .ZN(n7476)
         );
  OAI211_X1 U8042 ( .C1(n7495), .C2(n7478), .A(n7477), .B(n7476), .ZN(U2822)
         );
  OAI22_X1 U8043 ( .A1(n7535), .A2(n7480), .B1(n7479), .B2(n7531), .ZN(n7481)
         );
  AOI211_X1 U8044 ( .C1(n7519), .C2(EBX_REG_6__SCAN_IN), .A(n7487), .B(n7481), 
        .ZN(n7482) );
  OAI221_X1 U8045 ( .B1(REIP_REG_6__SCAN_IN), .B2(n7493), .C1(n6442), .C2(
        n7495), .A(n7482), .ZN(n7483) );
  AOI21_X1 U8046 ( .B1(n7522), .B2(n7484), .A(n7483), .ZN(n7485) );
  OAI21_X1 U8047 ( .B1(n7486), .B2(n7541), .A(n7485), .ZN(U2821) );
  AOI21_X1 U8048 ( .B1(n7501), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n7487), 
        .ZN(n7489) );
  NAND2_X1 U8049 ( .A1(n7519), .A2(EBX_REG_7__SCAN_IN), .ZN(n7488) );
  OAI211_X1 U8050 ( .C1(n7535), .C2(n7490), .A(n7489), .B(n7488), .ZN(n7497)
         );
  OAI21_X1 U8051 ( .B1(REIP_REG_6__SCAN_IN), .B2(REIP_REG_7__SCAN_IN), .A(
        n7491), .ZN(n7492) );
  OAI22_X1 U8052 ( .A1(n7495), .A2(n7494), .B1(n7493), .B2(n7492), .ZN(n7496)
         );
  AOI211_X1 U8053 ( .C1(n7498), .C2(n7522), .A(n7497), .B(n7496), .ZN(n7499)
         );
  OAI21_X1 U8054 ( .B1(n7500), .B2(n7541), .A(n7499), .ZN(U2820) );
  AOI22_X1 U8055 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n7501), .B1(
        EBX_REG_17__SCAN_IN), .B2(n7519), .ZN(n7509) );
  INV_X1 U8056 ( .A(n7502), .ZN(n7503) );
  AOI222_X1 U8057 ( .A1(n7696), .A2(n7522), .B1(n7505), .B2(n7504), .C1(n7521), 
        .C2(n7503), .ZN(n7508) );
  OAI221_X1 U8058 ( .B1(REIP_REG_17__SCAN_IN), .B2(REIP_REG_16__SCAN_IN), .C1(
        REIP_REG_17__SCAN_IN), .C2(n7506), .A(n7512), .ZN(n7507) );
  NAND4_X1 U8059 ( .A1(n7509), .A2(n7508), .A3(n7514), .A4(n7507), .ZN(U2810)
         );
  NOR3_X1 U8060 ( .A1(REIP_REG_19__SCAN_IN), .A2(n7511), .A3(n7510), .ZN(n7518) );
  INV_X1 U8061 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n7516) );
  OAI21_X1 U8062 ( .B1(n7513), .B2(n7512), .A(REIP_REG_19__SCAN_IN), .ZN(n7515) );
  OAI211_X1 U8063 ( .C1(n7531), .C2(n7516), .A(n7515), .B(n7514), .ZN(n7517)
         );
  AOI211_X1 U8064 ( .C1(n7519), .C2(EBX_REG_19__SCAN_IN), .A(n7518), .B(n7517), 
        .ZN(n7524) );
  AOI22_X1 U8065 ( .A1(n7699), .A2(n7522), .B1(n7521), .B2(n7520), .ZN(n7523)
         );
  OAI211_X1 U8066 ( .C1(n7525), .C2(n7541), .A(n7524), .B(n7523), .ZN(U2808)
         );
  OAI21_X1 U8067 ( .B1(n7528), .B2(n7527), .A(n7526), .ZN(n7533) );
  OAI22_X1 U8068 ( .A1(n4565), .A2(n7531), .B1(n7530), .B2(n7529), .ZN(n7532)
         );
  AOI21_X1 U8069 ( .B1(n7534), .B2(n7533), .A(n7532), .ZN(n7540) );
  OAI22_X1 U8070 ( .A1(n7705), .A2(n7537), .B1(n7536), .B2(n7535), .ZN(n7538)
         );
  INV_X1 U8071 ( .A(n7538), .ZN(n7539) );
  OAI211_X1 U8072 ( .C1(n7542), .C2(n7541), .A(n7540), .B(n7539), .ZN(U2804)
         );
  OAI21_X1 U8073 ( .B1(n7544), .B2(n7571), .A(n7543), .ZN(U2793) );
  INV_X1 U8074 ( .A(n4783), .ZN(n7547) );
  INV_X1 U8075 ( .A(n7545), .ZN(n7546) );
  NAND4_X1 U8076 ( .A1(n7549), .A2(n7548), .A3(n7547), .A4(n7546), .ZN(n7550)
         );
  OAI21_X1 U8077 ( .B1(n7552), .B2(n7551), .A(n7550), .ZN(U3455) );
  INV_X1 U8078 ( .A(n7553), .ZN(n7583) );
  INV_X1 U8079 ( .A(n7554), .ZN(n7630) );
  INV_X1 U8080 ( .A(n7555), .ZN(n7564) );
  NOR3_X1 U8081 ( .A1(n7557), .A2(n3937), .A3(n7556), .ZN(n7558) );
  NAND2_X1 U8082 ( .A1(n7558), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n7562) );
  OAI22_X1 U8083 ( .A1(n7560), .A2(n7559), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n7558), .ZN(n7561) );
  NAND2_X1 U8084 ( .A1(n7562), .A2(n7561), .ZN(n7563) );
  AOI222_X1 U8085 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n7564), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n7563), .C1(n7564), .C2(n7563), 
        .ZN(n7567) );
  INV_X1 U8086 ( .A(n7567), .ZN(n7569) );
  OAI21_X1 U8087 ( .B1(n7567), .B2(n7566), .A(n7565), .ZN(n7568) );
  OAI21_X1 U8088 ( .B1(n7569), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n7568), 
        .ZN(n7579) );
  INV_X1 U8089 ( .A(MORE_REG_SCAN_IN), .ZN(n7572) );
  AOI21_X1 U8090 ( .B1(n7572), .B2(n7571), .A(n7570), .ZN(n7574) );
  OR4_X1 U8091 ( .A1(n7576), .A2(n7575), .A3(n7574), .A4(n7573), .ZN(n7577) );
  AOI211_X1 U8092 ( .C1(n7579), .C2(n7130), .A(n7578), .B(n7577), .ZN(n7606)
         );
  AOI22_X1 U8093 ( .A1(n7606), .A2(n7581), .B1(READY_N), .B2(n7580), .ZN(n7582) );
  AOI21_X1 U8094 ( .B1(READY_N), .B2(n7584), .A(n7597), .ZN(n7595) );
  OAI21_X1 U8095 ( .B1(READY_N), .B2(n7585), .A(n7605), .ZN(n7588) );
  NAND2_X1 U8096 ( .A1(n7597), .A2(n7586), .ZN(n7587) );
  OAI21_X1 U8097 ( .B1(n7588), .B2(n7597), .A(n7587), .ZN(n7590) );
  OAI211_X1 U8098 ( .C1(n7595), .C2(n7591), .A(n7590), .B(n7589), .ZN(U3149)
         );
  AOI211_X1 U8099 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n7597), .A(n7593), .B(
        n7592), .ZN(n7594) );
  INV_X1 U8100 ( .A(n7594), .ZN(U3453) );
  NAND2_X1 U8101 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n7595), .ZN(n7601) );
  INV_X1 U8102 ( .A(n7596), .ZN(n7599) );
  AOI21_X1 U8103 ( .B1(n7599), .B2(n7598), .A(n7597), .ZN(n7600) );
  OAI22_X1 U8104 ( .A1(n7602), .A2(n7601), .B1(n7600), .B2(
        STATE2_REG_0__SCAN_IN), .ZN(n7604) );
  OAI211_X1 U8105 ( .C1(n7606), .C2(n7605), .A(n7604), .B(n7603), .ZN(U3148)
         );
  INV_X1 U8106 ( .A(n7607), .ZN(n7609) );
  OAI21_X1 U8107 ( .B1(n3658), .B2(n7608), .A(n7609), .ZN(U2792) );
  OAI21_X1 U8108 ( .B1(n3658), .B2(n7610), .A(n7609), .ZN(U3452) );
  AOI21_X1 U8109 ( .B1(READY_N), .B2(STATE_REG_1__SCAN_IN), .A(n7612), .ZN(
        n7613) );
  INV_X1 U8110 ( .A(n7613), .ZN(n7615) );
  INV_X1 U8111 ( .A(NA_N), .ZN(n7614) );
  AOI221_X1 U8112 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n7614), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n7625) );
  AOI21_X1 U8113 ( .B1(n7616), .B2(n7615), .A(n7625), .ZN(n7617) );
  OAI221_X1 U8114 ( .B1(n7309), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n7309), 
        .C2(n7618), .A(n7617), .ZN(U3181) );
  AOI221_X1 U8115 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n7634), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7620) );
  AOI221_X1 U8116 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n7620), .C2(HOLD), .A(n7619), .ZN(n7626) );
  OAI21_X1 U8117 ( .B1(NA_N), .B2(n7622), .A(n7621), .ZN(n7623) );
  NAND3_X1 U8118 ( .A1(READY_N), .A2(n7623), .A3(STATE_REG_1__SCAN_IN), .ZN(
        n7624) );
  OAI21_X1 U8119 ( .B1(n7626), .B2(n7625), .A(n7624), .ZN(U3183) );
  AOI22_X1 U8120 ( .A1(n7309), .A2(n7629), .B1(n7628), .B2(n7627), .ZN(U3473)
         );
  AOI22_X1 U8121 ( .A1(DATAI_0_), .A2(n7692), .B1(UWORD_REG_0__SCAN_IN), .B2(
        n7691), .ZN(n7635) );
  OAI21_X1 U8122 ( .B1(n7636), .B2(n7694), .A(n7635), .ZN(U2924) );
  AOI22_X1 U8123 ( .A1(DATAI_0_), .A2(n7692), .B1(LWORD_REG_0__SCAN_IN), .B2(
        n7691), .ZN(n7637) );
  OAI21_X1 U8124 ( .B1(n7638), .B2(n7694), .A(n7637), .ZN(U2939) );
  AOI22_X1 U8125 ( .A1(DATAI_1_), .A2(n7692), .B1(UWORD_REG_1__SCAN_IN), .B2(
        n7691), .ZN(n7639) );
  OAI21_X1 U8126 ( .B1(n4476), .B2(n7694), .A(n7639), .ZN(U2925) );
  AOI22_X1 U8127 ( .A1(DATAI_1_), .A2(n7692), .B1(LWORD_REG_1__SCAN_IN), .B2(
        n7691), .ZN(n7640) );
  OAI21_X1 U8128 ( .B1(n7641), .B2(n7694), .A(n7640), .ZN(U2940) );
  AOI22_X1 U8129 ( .A1(DATAI_2_), .A2(n7692), .B1(UWORD_REG_2__SCAN_IN), .B2(
        n7691), .ZN(n7642) );
  OAI21_X1 U8130 ( .B1(n7643), .B2(n7694), .A(n7642), .ZN(U2926) );
  AOI22_X1 U8131 ( .A1(DATAI_2_), .A2(n7692), .B1(LWORD_REG_2__SCAN_IN), .B2(
        n7691), .ZN(n7644) );
  OAI21_X1 U8132 ( .B1(n7645), .B2(n7694), .A(n7644), .ZN(U2941) );
  AOI22_X1 U8133 ( .A1(DATAI_3_), .A2(n7692), .B1(UWORD_REG_3__SCAN_IN), .B2(
        n7691), .ZN(n7646) );
  OAI21_X1 U8134 ( .B1(n4511), .B2(n7694), .A(n7646), .ZN(U2927) );
  AOI22_X1 U8135 ( .A1(DATAI_3_), .A2(n7692), .B1(LWORD_REG_3__SCAN_IN), .B2(
        n7691), .ZN(n7647) );
  OAI21_X1 U8136 ( .B1(n7648), .B2(n7694), .A(n7647), .ZN(U2942) );
  AOI22_X1 U8137 ( .A1(DATAI_4_), .A2(n7692), .B1(UWORD_REG_4__SCAN_IN), .B2(
        n7666), .ZN(n7649) );
  OAI21_X1 U8138 ( .B1(n7650), .B2(n7694), .A(n7649), .ZN(U2928) );
  AOI22_X1 U8139 ( .A1(DATAI_4_), .A2(n7692), .B1(LWORD_REG_4__SCAN_IN), .B2(
        n7666), .ZN(n7651) );
  OAI21_X1 U8140 ( .B1(n7652), .B2(n7694), .A(n7651), .ZN(U2943) );
  AOI22_X1 U8141 ( .A1(DATAI_5_), .A2(n7692), .B1(UWORD_REG_5__SCAN_IN), .B2(
        n7666), .ZN(n7653) );
  OAI21_X1 U8142 ( .B1(n7654), .B2(n7694), .A(n7653), .ZN(U2929) );
  AOI22_X1 U8143 ( .A1(DATAI_5_), .A2(n7692), .B1(LWORD_REG_5__SCAN_IN), .B2(
        n7666), .ZN(n7655) );
  OAI21_X1 U8144 ( .B1(n7656), .B2(n7694), .A(n7655), .ZN(U2944) );
  AOI22_X1 U8145 ( .A1(DATAI_6_), .A2(n7692), .B1(UWORD_REG_6__SCAN_IN), .B2(
        n7666), .ZN(n7657) );
  OAI21_X1 U8146 ( .B1(n7658), .B2(n7694), .A(n7657), .ZN(U2930) );
  AOI22_X1 U8147 ( .A1(DATAI_6_), .A2(n7692), .B1(LWORD_REG_6__SCAN_IN), .B2(
        n7666), .ZN(n7659) );
  OAI21_X1 U8148 ( .B1(n7660), .B2(n7694), .A(n7659), .ZN(U2945) );
  AOI22_X1 U8149 ( .A1(DATAI_7_), .A2(n7692), .B1(UWORD_REG_7__SCAN_IN), .B2(
        n7666), .ZN(n7661) );
  OAI21_X1 U8150 ( .B1(n7662), .B2(n7694), .A(n7661), .ZN(U2931) );
  AOI22_X1 U8151 ( .A1(DATAI_7_), .A2(n7692), .B1(LWORD_REG_7__SCAN_IN), .B2(
        n7666), .ZN(n7663) );
  OAI21_X1 U8152 ( .B1(n4304), .B2(n7694), .A(n7663), .ZN(U2946) );
  AOI22_X1 U8153 ( .A1(DATAI_8_), .A2(n7692), .B1(UWORD_REG_8__SCAN_IN), .B2(
        n7666), .ZN(n7664) );
  OAI21_X1 U8154 ( .B1(n7665), .B2(n7694), .A(n7664), .ZN(U2932) );
  AOI22_X1 U8155 ( .A1(DATAI_8_), .A2(n7692), .B1(LWORD_REG_8__SCAN_IN), .B2(
        n7666), .ZN(n7667) );
  OAI21_X1 U8156 ( .B1(n7668), .B2(n7694), .A(n7667), .ZN(U2947) );
  AOI22_X1 U8157 ( .A1(DATAI_9_), .A2(n7692), .B1(UWORD_REG_9__SCAN_IN), .B2(
        n7691), .ZN(n7669) );
  OAI21_X1 U8158 ( .B1(n7670), .B2(n7694), .A(n7669), .ZN(U2933) );
  AOI22_X1 U8159 ( .A1(DATAI_9_), .A2(n7692), .B1(LWORD_REG_9__SCAN_IN), .B2(
        n7691), .ZN(n7671) );
  OAI21_X1 U8160 ( .B1(n7672), .B2(n7694), .A(n7671), .ZN(U2948) );
  AOI22_X1 U8161 ( .A1(DATAI_10_), .A2(n7692), .B1(UWORD_REG_10__SCAN_IN), 
        .B2(n7691), .ZN(n7673) );
  OAI21_X1 U8162 ( .B1(n7674), .B2(n7694), .A(n7673), .ZN(U2934) );
  AOI22_X1 U8163 ( .A1(DATAI_10_), .A2(n7692), .B1(LWORD_REG_10__SCAN_IN), 
        .B2(n7691), .ZN(n7675) );
  OAI21_X1 U8164 ( .B1(n7676), .B2(n7694), .A(n7675), .ZN(U2949) );
  AOI22_X1 U8165 ( .A1(DATAI_11_), .A2(n7692), .B1(UWORD_REG_11__SCAN_IN), 
        .B2(n7691), .ZN(n7677) );
  OAI21_X1 U8166 ( .B1(n4669), .B2(n7694), .A(n7677), .ZN(U2935) );
  AOI22_X1 U8167 ( .A1(DATAI_11_), .A2(n7692), .B1(LWORD_REG_11__SCAN_IN), 
        .B2(n7691), .ZN(n7678) );
  OAI21_X1 U8168 ( .B1(n7679), .B2(n7694), .A(n7678), .ZN(U2950) );
  AOI22_X1 U8169 ( .A1(DATAI_12_), .A2(n7692), .B1(UWORD_REG_12__SCAN_IN), 
        .B2(n7691), .ZN(n7680) );
  OAI21_X1 U8170 ( .B1(n7681), .B2(n7694), .A(n7680), .ZN(U2936) );
  AOI22_X1 U8171 ( .A1(DATAI_12_), .A2(n7692), .B1(LWORD_REG_12__SCAN_IN), 
        .B2(n7691), .ZN(n7682) );
  OAI21_X1 U8172 ( .B1(n7683), .B2(n7694), .A(n7682), .ZN(U2951) );
  AOI22_X1 U8173 ( .A1(DATAI_13_), .A2(n7692), .B1(UWORD_REG_13__SCAN_IN), 
        .B2(n7691), .ZN(n7684) );
  OAI21_X1 U8174 ( .B1(n4712), .B2(n7694), .A(n7684), .ZN(U2937) );
  AOI22_X1 U8175 ( .A1(DATAI_13_), .A2(n7692), .B1(LWORD_REG_13__SCAN_IN), 
        .B2(n7691), .ZN(n7685) );
  OAI21_X1 U8176 ( .B1(n7686), .B2(n7694), .A(n7685), .ZN(U2952) );
  AOI22_X1 U8177 ( .A1(DATAI_14_), .A2(n7692), .B1(UWORD_REG_14__SCAN_IN), 
        .B2(n7691), .ZN(n7687) );
  OAI21_X1 U8178 ( .B1(n7688), .B2(n7694), .A(n7687), .ZN(U2938) );
  AOI22_X1 U8179 ( .A1(DATAI_14_), .A2(n7692), .B1(LWORD_REG_14__SCAN_IN), 
        .B2(n7691), .ZN(n7689) );
  OAI21_X1 U8180 ( .B1(n7690), .B2(n7694), .A(n7689), .ZN(U2953) );
  AOI22_X1 U8181 ( .A1(DATAI_15_), .A2(n7692), .B1(LWORD_REG_15__SCAN_IN), 
        .B2(n7691), .ZN(n7693) );
  OAI21_X1 U8182 ( .B1(n7695), .B2(n7694), .A(n7693), .ZN(U2954) );
  AOI22_X1 U8183 ( .A1(n7696), .A2(n7707), .B1(n7706), .B2(DATAI_17_), .ZN(
        n7698) );
  AOI22_X1 U8184 ( .A1(n7710), .A2(DATAI_1_), .B1(n7709), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n7697) );
  NAND2_X1 U8185 ( .A1(n7698), .A2(n7697), .ZN(U2874) );
  AOI22_X1 U8186 ( .A1(n7699), .A2(n7707), .B1(n7706), .B2(DATAI_19_), .ZN(
        n7701) );
  AOI22_X1 U8187 ( .A1(n7710), .A2(DATAI_3_), .B1(n7709), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n7700) );
  NAND2_X1 U8188 ( .A1(n7701), .A2(n7700), .ZN(U2872) );
  AOI22_X1 U8189 ( .A1(n7702), .A2(n7707), .B1(n7706), .B2(DATAI_21_), .ZN(
        n7704) );
  AOI22_X1 U8190 ( .A1(n7710), .A2(DATAI_5_), .B1(n7709), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n7703) );
  NAND2_X1 U8191 ( .A1(n7704), .A2(n7703), .ZN(U2870) );
  INV_X1 U8192 ( .A(n7705), .ZN(n7708) );
  AOI22_X1 U8193 ( .A1(n7708), .A2(n7707), .B1(n7706), .B2(DATAI_23_), .ZN(
        n7712) );
  AOI22_X1 U8194 ( .A1(n7710), .A2(DATAI_7_), .B1(n7709), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n7711) );
  NAND2_X1 U8195 ( .A1(n7712), .A2(n7711), .ZN(U2868) );
  CLKBUF_X1 U3715 ( .A(n3928), .Z(n5094) );
  CLKBUF_X1 U3774 ( .A(n7164), .Z(n7169) );
endmodule

