

module b22_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16363, n16364, n16365, n16366,
         n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
         n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
         n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
         n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
         n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
         n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
         n16415, n16416, n16417, n16418, n16419, n16423;

  INV_X1 U7522 ( .A(n13341), .ZN(n13411) );
  BUF_X2 U7523 ( .A(n13038), .Z(n8633) );
  CLKBUF_X2 U7524 ( .A(n9732), .Z(n13386) );
  INV_X1 U7525 ( .A(n13378), .ZN(n9659) );
  AND4_X1 U7526 ( .A1(n8818), .A2(n8817), .A3(n8816), .A4(n8815), .ZN(n16104)
         );
  AND2_X1 U7527 ( .A1(n14680), .A2(n12848), .ZN(n9732) );
  INV_X2 U7528 ( .A(n12551), .ZN(n12682) );
  NAND2_X1 U7529 ( .A1(n12540), .A2(n16039), .ZN(n12547) );
  NAND2_X1 U7530 ( .A1(n10860), .A2(n15095), .ZN(n12553) );
  AND2_X2 U7531 ( .A1(n10080), .A2(n10081), .ZN(n12526) );
  INV_X1 U7532 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n15627) );
  INV_X4 U7533 ( .A(n14549), .ZN(n16405) );
  INV_X1 U7535 ( .A(n16423), .ZN(n7422) );
  INV_X1 U7536 ( .A(n8012), .ZN(n12494) );
  INV_X1 U7537 ( .A(n10228), .ZN(n11234) );
  AND2_X1 U7538 ( .A1(n9344), .A2(n8323), .ZN(n7664) );
  OR2_X1 U7539 ( .A1(n9578), .A2(n7582), .ZN(n7734) );
  INV_X1 U7540 ( .A(n12518), .ZN(n12203) );
  CLKBUF_X2 U7541 ( .A(n11234), .Z(n8541) );
  AND2_X1 U7542 ( .A1(n10080), .A2(n12308), .ZN(n12685) );
  INV_X1 U7543 ( .A(n12316), .ZN(n12398) );
  AND2_X1 U7544 ( .A1(n7663), .A2(n7661), .ZN(n7660) );
  INV_X1 U7546 ( .A(n10763), .ZN(n12836) );
  INV_X1 U7547 ( .A(n8825), .ZN(n7738) );
  XNOR2_X1 U7548 ( .A(n8367), .B(n12849), .ZN(n9271) );
  INV_X1 U7549 ( .A(n9419), .ZN(n12709) );
  AND2_X1 U7550 ( .A1(n7736), .A2(n7735), .ZN(n15812) );
  INV_X1 U7551 ( .A(n11830), .ZN(n13109) );
  NAND3_X1 U7552 ( .A1(n8090), .A2(n7642), .A3(n7641), .ZN(n16079) );
  NAND2_X1 U7553 ( .A1(n7655), .A2(n10012), .ZN(n13078) );
  OAI21_X1 U7554 ( .B1(n9271), .B2(n16107), .A(n9270), .ZN(n13743) );
  NAND2_X1 U7555 ( .A1(n14113), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8800) );
  OAI21_X1 U7556 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n10797), .A(n10643), .ZN(
        n10644) );
  INV_X1 U7557 ( .A(n9660), .ZN(n14301) );
  INV_X1 U7558 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9344) );
  NAND2_X1 U7559 ( .A1(n11830), .A2(n10095), .ZN(n13321) );
  AND2_X1 U7560 ( .A1(n12316), .A2(n10095), .ZN(n7423) );
  NAND2_X2 U7561 ( .A1(n15971), .A2(n13643), .ZN(n13644) );
  OR2_X2 U7562 ( .A1(n10696), .A2(n10695), .ZN(n8282) );
  OAI211_X1 U7563 ( .C1(n8873), .C2(n9474), .A(n8858), .B(n8857), .ZN(n12881)
         );
  OR2_X2 U7565 ( .A1(n13260), .A2(n7859), .ZN(n7850) );
  OAI21_X2 U7566 ( .B1(n9890), .B2(n9823), .A(n9662), .ZN(n9663) );
  INV_X4 U7567 ( .A(n8874), .ZN(n9092) );
  AOI21_X2 U7568 ( .B1(n14950), .B2(n14949), .A(n8032), .ZN(n14934) );
  CLKBUF_X2 U7569 ( .A(n13420), .Z(n7424) );
  OAI21_X2 U7570 ( .B1(n9503), .B2(n8161), .A(n9506), .ZN(n9515) );
  AOI21_X2 U7571 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n14288), .A(n14282), .ZN(
        n14295) );
  NAND2_X2 U7572 ( .A1(n13884), .A2(n9248), .ZN(n13872) );
  NAND2_X2 U7573 ( .A1(n8005), .A2(n11782), .ZN(n12616) );
  AOI21_X2 U7574 ( .B1(n10703), .B2(n10702), .A(n10701), .ZN(n10954) );
  XNOR2_X2 U7575 ( .A(n8800), .B(n8799), .ZN(n13465) );
  CLKBUF_X1 U7576 ( .A(n12685), .Z(n7425) );
  BUF_X4 U7578 ( .A(n12685), .Z(n7427) );
  NOR2_X2 U7579 ( .A1(n10560), .A2(n7474), .ZN(n10691) );
  NOR2_X2 U7580 ( .A1(n10503), .A2(n10502), .ZN(n10560) );
  OAI211_X2 U7581 ( .C1(n8874), .C2(n9457), .A(n8824), .B(n8823), .ZN(n8825)
         );
  OAI21_X2 U7582 ( .B1(n10954), .B2(n10953), .A(n10952), .ZN(n11115) );
  NAND2_X2 U7583 ( .A1(n10399), .A2(n10398), .ZN(n16246) );
  INV_X1 U7584 ( .A(n12992), .ZN(n9130) );
  AOI22_X2 U7585 ( .A1(n10492), .A2(n10491), .B1(n10497), .B2(n10490), .ZN(
        n10566) );
  OAI22_X2 U7586 ( .A1(n10469), .A2(n10468), .B1(n10292), .B2(n10485), .ZN(
        n10492) );
  NAND2_X4 U7587 ( .A1(n10155), .A2(n12183), .ZN(n12483) );
  XNOR2_X2 U7588 ( .A(n9400), .B(n9401), .ZN(n15786) );
  AOI21_X1 U7589 ( .B1(n7773), .B2(n14529), .A(n8039), .ZN(n14565) );
  NAND2_X1 U7590 ( .A1(n15008), .A2(n15007), .ZN(n15006) );
  NOR2_X1 U7591 ( .A1(n13711), .A2(n13710), .ZN(n13715) );
  OR2_X1 U7592 ( .A1(n9166), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9178) );
  NAND2_X1 U7593 ( .A1(n9786), .A2(n9785), .ZN(n13146) );
  NAND2_X2 U7594 ( .A1(n12868), .A2(n12866), .ZN(n16050) );
  NAND2_X1 U7595 ( .A1(n9731), .A2(n9730), .ZN(n16169) );
  INV_X1 U7596 ( .A(n14224), .ZN(n16127) );
  INV_X2 U7597 ( .A(n16104), .ZN(n7428) );
  CLKBUF_X2 U7598 ( .A(n9789), .Z(n11931) );
  AND2_X1 U7599 ( .A1(n7734), .A2(n7733), .ZN(n9590) );
  NAND2_X1 U7600 ( .A1(n7430), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8269) );
  INV_X2 U7601 ( .A(n12016), .ZN(n12686) );
  AOI21_X1 U7602 ( .B1(n9408), .B2(n7907), .A(n7532), .ZN(n7906) );
  NAND2_X1 U7603 ( .A1(n9546), .A2(n9635), .ZN(n14314) );
  NAND2_X1 U7604 ( .A1(n9419), .A2(P3_U3151), .ZN(n14119) );
  INV_X2 U7605 ( .A(n9419), .ZN(n12298) );
  NAND4_X1 U7606 ( .A1(n7660), .A2(n7662), .A3(n7489), .A4(n7659), .ZN(n10012)
         );
  INV_X2 U7607 ( .A(n9360), .ZN(n9419) );
  AND4_X1 U7608 ( .A1(n9532), .A2(n9531), .A3(n9530), .A4(n9529), .ZN(n9537)
         );
  INV_X2 U7609 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  AOI21_X1 U7610 ( .B1(n8211), .B2(n8210), .A(n8209), .ZN(n8249) );
  NAND2_X1 U7611 ( .A1(n13972), .A2(n13971), .ZN(n14038) );
  XNOR2_X1 U7612 ( .A(n13024), .B(n12849), .ZN(n8036) );
  AND2_X1 U7613 ( .A1(n13779), .A2(n13778), .ZN(n14041) );
  NAND2_X1 U7614 ( .A1(n13760), .A2(n12970), .ZN(n13024) );
  XNOR2_X1 U7615 ( .A(n13784), .B(n13785), .ZN(n14051) );
  AND2_X1 U7616 ( .A1(n13756), .A2(n13755), .ZN(n13972) );
  NAND2_X1 U7617 ( .A1(n8207), .A2(n9257), .ZN(n13784) );
  NAND2_X1 U7618 ( .A1(n8017), .A2(n7593), .ZN(n7985) );
  OAI211_X1 U7619 ( .C1(n14566), .C2(n16262), .A(n14565), .B(n14564), .ZN(
        n14646) );
  AND2_X1 U7620 ( .A1(n8068), .A2(n8067), .ZN(n14571) );
  OR2_X1 U7621 ( .A1(n14565), .A2(n16405), .ZN(n8616) );
  NAND2_X1 U7622 ( .A1(n13796), .A2(n8205), .ZN(n8203) );
  NAND2_X1 U7623 ( .A1(n7638), .A2(n12853), .ZN(n13796) );
  NAND2_X1 U7624 ( .A1(n14778), .A2(n14777), .ZN(n14776) );
  NOR2_X1 U7625 ( .A1(n14366), .A2(n14358), .ZN(n14360) );
  NAND3_X1 U7626 ( .A1(n8588), .A2(n8587), .A3(n8589), .ZN(n8585) );
  NOR2_X1 U7627 ( .A1(n13715), .A2(n7979), .ZN(n13716) );
  OAI21_X1 U7628 ( .B1(n13833), .B2(n12962), .A(n12957), .ZN(n13826) );
  NAND2_X1 U7629 ( .A1(n14406), .A2(n7510), .ZN(n8588) );
  AOI21_X1 U7630 ( .B1(n14423), .B2(n14420), .A(n7475), .ZN(n14406) );
  NAND2_X1 U7631 ( .A1(n14351), .A2(n7485), .ZN(n14423) );
  NAND2_X1 U7632 ( .A1(n8066), .A2(n8596), .ZN(n14435) );
  NAND2_X1 U7633 ( .A1(n7652), .A2(n7651), .ZN(n12362) );
  NAND2_X1 U7634 ( .A1(n12274), .A2(n12273), .ZN(n14125) );
  NAND2_X1 U7635 ( .A1(n7654), .A2(n7653), .ZN(n11981) );
  NAND2_X1 U7636 ( .A1(n8197), .A2(n8196), .ZN(n13921) );
  AND2_X1 U7637 ( .A1(n8470), .A2(n8472), .ZN(n12147) );
  NAND2_X1 U7638 ( .A1(n11735), .A2(n11878), .ZN(n11974) );
  OR2_X1 U7639 ( .A1(n13654), .A2(n13655), .ZN(n8284) );
  NAND2_X1 U7640 ( .A1(n11334), .A2(n11333), .ZN(n13202) );
  NOR2_X1 U7641 ( .A1(n9178), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9195) );
  OR2_X1 U7642 ( .A1(n11462), .A2(n11461), .ZN(n13636) );
  AND2_X1 U7643 ( .A1(n8282), .A2(n8281), .ZN(n11109) );
  NOR2_X1 U7644 ( .A1(n11460), .A2(n11459), .ZN(n11462) );
  OR2_X1 U7645 ( .A1(n10713), .A2(n10712), .ZN(n8442) );
  NAND2_X1 U7646 ( .A1(n11548), .A2(n11547), .ZN(n12601) );
  INV_X1 U7647 ( .A(n12731), .ZN(n7429) );
  NAND2_X1 U7648 ( .A1(n8091), .A2(n11364), .ZN(n12592) );
  OAI21_X1 U7649 ( .B1(n14520), .B2(n10417), .A(n14549), .ZN(n14497) );
  OR2_X1 U7650 ( .A1(n9229), .A2(n13004), .ZN(n11414) );
  AND2_X1 U7651 ( .A1(n12901), .A2(n12902), .ZN(n13000) );
  AND2_X1 U7652 ( .A1(n12877), .A2(n12870), .ZN(n13001) );
  NAND2_X1 U7653 ( .A1(n12887), .A2(n12886), .ZN(n9223) );
  NAND2_X1 U7654 ( .A1(n7998), .A2(n9722), .ZN(n14224) );
  NAND2_X1 U7655 ( .A1(n7906), .A2(n7905), .ZN(n9424) );
  AND3_X1 U7656 ( .A1(n8893), .A2(n8892), .A3(n8891), .ZN(n16215) );
  NAND2_X2 U7657 ( .A1(n9642), .A2(n7971), .ZN(n14266) );
  NAND4_X1 U7658 ( .A1(n8885), .A2(n8884), .A3(n8883), .A4(n8882), .ZN(n13618)
         );
  NAND4_X1 U7659 ( .A1(n8809), .A2(n7639), .A3(n8215), .A4(n8810), .ZN(n13624)
         );
  AND4_X1 U7660 ( .A1(n8841), .A2(n8840), .A3(n8839), .A4(n8838), .ZN(n16102)
         );
  AOI21_X1 U7661 ( .B1(P3_REG2_REG_4__SCAN_IN), .B2(n10485), .A(n10482), .ZN(
        n10505) );
  AND4_X1 U7662 ( .A1(n8831), .A2(n8830), .A3(n8829), .A4(n8828), .ZN(n16052)
         );
  AND4_X1 U7663 ( .A1(n8868), .A2(n8867), .A3(n8866), .A4(n8865), .ZN(n11306)
         );
  NAND2_X1 U7664 ( .A1(n9209), .A2(n9272), .ZN(n10454) );
  NAND2_X2 U7665 ( .A1(n7470), .A2(n8269), .ZN(n14547) );
  NAND4_X1 U7666 ( .A1(n9668), .A2(n9667), .A3(n9666), .A4(n9665), .ZN(n14265)
         );
  NAND2_X1 U7667 ( .A1(n9214), .A2(n9213), .ZN(n10314) );
  INV_X2 U7668 ( .A(n13321), .ZN(n9720) );
  NAND2_X2 U7669 ( .A1(n8804), .A2(n14120), .ZN(n12992) );
  NAND2_X2 U7670 ( .A1(n8398), .A2(n9419), .ZN(n8873) );
  NAND2_X1 U7671 ( .A1(n9356), .A2(n15253), .ZN(n10157) );
  CLKBUF_X1 U7672 ( .A(n13378), .Z(n8004) );
  INV_X1 U7673 ( .A(n13378), .ZN(n7430) );
  INV_X4 U7674 ( .A(n13038), .ZN(n8634) );
  OAI21_X1 U7675 ( .B1(n10095), .B2(n8047), .A(n8046), .ZN(n9387) );
  XNOR2_X1 U7676 ( .A(n8190), .B(n8802), .ZN(n14120) );
  NAND2_X1 U7677 ( .A1(n9348), .A2(n10106), .ZN(n16039) );
  XNOR2_X1 U7678 ( .A(n10013), .B(n15237), .ZN(n15243) );
  BUF_X1 U7679 ( .A(n12709), .Z(n8006) );
  INV_X1 U7680 ( .A(n9362), .ZN(n9366) );
  NAND2_X2 U7681 ( .A1(n10095), .A2(P3_U3151), .ZN(n13462) );
  NAND2_X1 U7682 ( .A1(n7752), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7751) );
  MUX2_X1 U7683 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9545), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n9546) );
  XNOR2_X1 U7684 ( .A(n9840), .B(P1_IR_REG_21__SCAN_IN), .ZN(n12540) );
  XNOR2_X1 U7685 ( .A(n9544), .B(P2_IR_REG_21__SCAN_IN), .ZN(n13350) );
  NAND2_X1 U7686 ( .A1(n8801), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8190) );
  NAND2_X1 U7687 ( .A1(n10095), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8046) );
  NAND2_X1 U7688 ( .A1(n10109), .A2(n10108), .ZN(n12752) );
  NAND2_X1 U7689 ( .A1(n10012), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8181) );
  XNOR2_X1 U7690 ( .A(n9843), .B(P1_IR_REG_22__SCAN_IN), .ZN(n15263) );
  NAND2_X1 U7691 ( .A1(n7686), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10013) );
  NAND2_X1 U7692 ( .A1(n9635), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9540) );
  OAI21_X1 U7693 ( .B1(n9360), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n7993), .ZN(
        n9362) );
  OR2_X1 U7694 ( .A1(n10319), .A2(n8813), .ZN(n10317) );
  AND3_X1 U7695 ( .A1(n8561), .A2(n9410), .A3(n9346), .ZN(n10104) );
  XNOR2_X1 U7696 ( .A(n9405), .B(n9404), .ZN(n9723) );
  AND2_X1 U7697 ( .A1(n8871), .A2(n8781), .ZN(n7629) );
  XNOR2_X1 U7698 ( .A(n7835), .B(n8856), .ZN(n10485) );
  AND2_X1 U7699 ( .A1(n9346), .A2(n9410), .ZN(n10526) );
  NOR2_X1 U7700 ( .A1(n9334), .A2(n8056), .ZN(n9543) );
  NAND2_X1 U7701 ( .A1(n8159), .A2(n8157), .ZN(n9360) );
  NAND2_X1 U7702 ( .A1(n8430), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8834) );
  NOR2_X1 U7703 ( .A1(n8786), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n8653) );
  OR2_X1 U7704 ( .A1(n8879), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8894) );
  AND2_X1 U7705 ( .A1(n8777), .A2(n8214), .ZN(n7630) );
  AND4_X1 U7706 ( .A1(n8780), .A2(n8779), .A3(n8981), .A4(n8778), .ZN(n8781)
         );
  AND2_X1 U7707 ( .A1(n8651), .A2(n8788), .ZN(n7750) );
  AND4_X1 U7708 ( .A1(n9329), .A2(n9328), .A3(n9327), .A4(n9326), .ZN(n9332)
         );
  AND3_X1 U7709 ( .A1(n7650), .A2(n7649), .A3(n7648), .ZN(n7662) );
  AND4_X1 U7710 ( .A1(n9524), .A2(n9345), .A3(n9523), .A4(n15648), .ZN(n7663)
         );
  NAND3_X1 U7711 ( .A1(n8391), .A2(n8390), .A3(n8774), .ZN(n8844) );
  AND4_X1 U7712 ( .A1(n8776), .A2(n8889), .A3(n8888), .A4(n8922), .ZN(n8777)
         );
  AND2_X1 U7713 ( .A1(n9403), .A2(n9404), .ZN(n9396) );
  AND3_X1 U7714 ( .A1(n9331), .A2(n9330), .A3(n9427), .ZN(n9494) );
  INV_X1 U7715 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n15649) );
  INV_X1 U7716 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9534) );
  INV_X1 U7717 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9535) );
  INV_X1 U7718 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9529) );
  INV_X1 U7719 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9523) );
  INV_X1 U7720 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n9533) );
  NOR2_X1 U7721 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n9328) );
  NOR2_X1 U7722 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n7650) );
  INV_X1 U7723 ( .A(P2_RD_REG_SCAN_IN), .ZN(n8796) );
  NOR2_X1 U7724 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n7649) );
  NOR2_X1 U7725 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n7648) );
  NOR2_X1 U7726 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n8780) );
  NOR2_X1 U7727 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n8779) );
  INV_X1 U7728 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9427) );
  INV_X1 U7729 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8390) );
  INV_X1 U7730 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8774) );
  NOR2_X1 U7731 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n8784) );
  INV_X1 U7732 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8889) );
  INV_X1 U7733 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8888) );
  NOR2_X1 U7734 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n9331) );
  NOR2_X1 U7735 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n9330) );
  INV_X4 U7736 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7737 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9205) );
  INV_X1 U7738 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8922) );
  NOR2_X1 U7739 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n9327) );
  INV_X1 U7740 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n15650) );
  NOR2_X1 U7741 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n8776) );
  NOR2_X1 U7742 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n9326) );
  INV_X1 U7743 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8981) );
  AOI21_X2 U7744 ( .B1(n14339), .B2(n14338), .A(n14337), .ZN(n14528) );
  NAND2_X1 U7745 ( .A1(n7784), .A2(n11925), .ZN(n14339) );
  NOR2_X1 U7746 ( .A1(n15946), .A2(n15947), .ZN(n15945) );
  NAND2_X1 U7747 ( .A1(n7749), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9405) );
  NOR2_X2 U7748 ( .A1(n12049), .A2(n14336), .ZN(n8277) );
  BUF_X4 U7749 ( .A(n14534), .Z(n7431) );
  NAND2_X1 U7750 ( .A1(n9809), .A2(n10793), .ZN(n14534) );
  NOR2_X2 U7751 ( .A1(n14508), .A2(n14609), .ZN(n14490) );
  INV_X1 U7753 ( .A(n7423), .ZN(n7432) );
  INV_X2 U7754 ( .A(n7423), .ZN(n7433) );
  NOR2_X2 U7755 ( .A1(n13183), .A2(n10813), .ZN(n11282) );
  NAND2_X1 U7756 ( .A1(n11830), .A2(n9419), .ZN(n13378) );
  INV_X1 U7757 ( .A(n13321), .ZN(n7434) );
  OR2_X1 U7758 ( .A1(n13482), .A2(n13838), .ZN(n12861) );
  NOR2_X1 U7759 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n9845) );
  CLKBUF_X1 U7760 ( .A(n9041), .Z(n9086) );
  INV_X1 U7761 ( .A(n13465), .ZN(n8804) );
  NOR2_X1 U7762 ( .A1(n7595), .A2(n7746), .ZN(n7745) );
  INV_X1 U7763 ( .A(n9250), .ZN(n7746) );
  AND2_X1 U7764 ( .A1(n8653), .A2(n8787), .ZN(n8652) );
  INV_X1 U7765 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8787) );
  INV_X1 U7766 ( .A(n12848), .ZN(n9638) );
  NAND2_X1 U7767 ( .A1(n8305), .A2(n8308), .ZN(n8301) );
  NAND2_X1 U7768 ( .A1(n14401), .A2(n14355), .ZN(n8309) );
  NAND2_X1 U7769 ( .A1(n12490), .A2(n12489), .ZN(n8549) );
  OAI21_X1 U7770 ( .B1(n9515), .B2(n7762), .A(n7759), .ZN(n10522) );
  AND2_X1 U7771 ( .A1(n7760), .A2(n8141), .ZN(n7759) );
  AOI21_X1 U7772 ( .B1(n8144), .B2(n8146), .A(n8142), .ZN(n8141) );
  NAND2_X1 U7773 ( .A1(n7761), .A2(n7911), .ZN(n7760) );
  NAND2_X1 U7774 ( .A1(n7829), .A2(n7828), .ZN(n8440) );
  INV_X1 U7775 ( .A(n10510), .ZN(n7828) );
  INV_X1 U7776 ( .A(n10511), .ZN(n7829) );
  NAND2_X1 U7777 ( .A1(n9115), .A2(n12956), .ZN(n13833) );
  NAND2_X1 U7778 ( .A1(n13812), .A2(n13813), .ZN(n7638) );
  NAND2_X1 U7779 ( .A1(n8399), .A2(n8634), .ZN(n8398) );
  NAND2_X1 U7780 ( .A1(n9284), .A2(n9285), .ZN(n9500) );
  NOR2_X1 U7781 ( .A1(n13435), .A2(n8612), .ZN(n8611) );
  INV_X1 U7782 ( .A(n11250), .ZN(n8612) );
  NAND2_X1 U7783 ( .A1(n14943), .A2(n13075), .ZN(n14926) );
  NAND2_X2 U7784 ( .A1(n15245), .A2(n13078), .ZN(n12316) );
  INV_X2 U7785 ( .A(n9419), .ZN(n10095) );
  NAND2_X1 U7786 ( .A1(n13162), .A2(n13163), .ZN(n8701) );
  NAND2_X1 U7787 ( .A1(n12627), .A2(n12624), .ZN(n7918) );
  NAND2_X1 U7788 ( .A1(n7467), .A2(n13214), .ZN(n8097) );
  INV_X1 U7789 ( .A(n8112), .ZN(n8114) );
  NAND2_X1 U7790 ( .A1(n13239), .A2(n13238), .ZN(n8710) );
  INV_X1 U7791 ( .A(n12658), .ZN(n7925) );
  NAND2_X1 U7792 ( .A1(n13304), .A2(n8683), .ZN(n8682) );
  NOR2_X1 U7793 ( .A1(n11354), .A2(n8340), .ZN(n8339) );
  INV_X1 U7794 ( .A(n11051), .ZN(n8340) );
  NAND2_X1 U7795 ( .A1(n14860), .A2(n16090), .ZN(n12555) );
  NAND2_X1 U7796 ( .A1(n10958), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8441) );
  NAND2_X1 U7797 ( .A1(n11669), .A2(n13000), .ZN(n7632) );
  INV_X1 U7798 ( .A(n9257), .ZN(n8206) );
  AOI21_X1 U7799 ( .B1(n8374), .B2(n8372), .A(n7517), .ZN(n8371) );
  AND2_X1 U7800 ( .A1(n13801), .A2(n9165), .ZN(n8259) );
  AND2_X1 U7801 ( .A1(n9258), .A2(n9257), .ZN(n13797) );
  AND2_X1 U7802 ( .A1(n7567), .A2(n8651), .ZN(n7870) );
  NAND2_X1 U7803 ( .A1(n13403), .A2(n13395), .ZN(n13407) );
  INV_X1 U7804 ( .A(n13416), .ZN(n8129) );
  AND2_X1 U7805 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(n13367), .ZN(n13381) );
  AND2_X1 U7806 ( .A1(n8585), .A2(n8583), .ZN(n14366) );
  NOR2_X1 U7807 ( .A1(n14368), .A2(n8584), .ZN(n8583) );
  INV_X1 U7808 ( .A(n8586), .ZN(n8584) );
  AOI21_X1 U7809 ( .B1(n8299), .B2(n8301), .A(n8298), .ZN(n8297) );
  OR2_X1 U7810 ( .A1(n8303), .A2(n8300), .ZN(n8299) );
  INV_X1 U7811 ( .A(n8308), .ZN(n8300) );
  AND2_X1 U7812 ( .A1(n8304), .A2(n14384), .ZN(n8303) );
  NAND2_X1 U7813 ( .A1(n8305), .A2(n8307), .ZN(n8304) );
  NOR2_X1 U7814 ( .A1(n8610), .A2(n8599), .ZN(n8598) );
  AND2_X1 U7815 ( .A1(n14599), .A2(n14350), .ZN(n8610) );
  INV_X1 U7816 ( .A(n8601), .ZN(n8599) );
  NAND2_X1 U7817 ( .A1(n14599), .A2(n14437), .ZN(n8321) );
  XNOR2_X1 U7818 ( .A(n14547), .B(n14266), .ZN(n13420) );
  INV_X1 U7819 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n9538) );
  NAND2_X1 U7820 ( .A1(n14849), .A2(n8541), .ZN(n12117) );
  OR2_X1 U7821 ( .A1(n9851), .A2(n8169), .ZN(n8168) );
  NOR2_X1 U7822 ( .A1(n7665), .A2(n9850), .ZN(n9851) );
  NAND2_X1 U7823 ( .A1(n15006), .A2(n8354), .ZN(n8353) );
  NOR2_X1 U7824 ( .A1(n14984), .A2(n8355), .ZN(n8354) );
  INV_X1 U7825 ( .A(n13069), .ZN(n8355) );
  NOR2_X1 U7826 ( .A1(n12739), .A2(n8672), .ZN(n8671) );
  INV_X1 U7827 ( .A(n12006), .ZN(n8672) );
  NAND2_X1 U7828 ( .A1(n16079), .A2(n10123), .ZN(n12552) );
  NAND2_X1 U7829 ( .A1(n12555), .A2(n12552), .ZN(n8087) );
  INV_X1 U7830 ( .A(n15108), .ZN(n13076) );
  NAND2_X1 U7831 ( .A1(n10791), .A2(n10790), .ZN(n10912) );
  AND2_X1 U7832 ( .A1(n8721), .A2(n15658), .ZN(n8561) );
  AND2_X1 U7833 ( .A1(n10523), .A2(n10247), .ZN(n10521) );
  INV_X1 U7834 ( .A(n9504), .ZN(n8161) );
  XNOR2_X1 U7835 ( .A(n9505), .B(SI_9_), .ZN(n9503) );
  INV_X1 U7836 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n15730) );
  OAI21_X1 U7837 ( .B1(n15679), .B2(n15710), .A(n15707), .ZN(n15731) );
  NAND2_X1 U7838 ( .A1(n10458), .A2(n16104), .ZN(n8631) );
  INV_X1 U7839 ( .A(n9086), .ZN(n9201) );
  AND4_X1 U7840 ( .A1(n8917), .A2(n8916), .A3(n8915), .A4(n8914), .ZN(n11860)
         );
  NAND2_X1 U7841 ( .A1(n8803), .A2(n13465), .ZN(n12988) );
  NAND2_X1 U7842 ( .A1(n8804), .A2(n8803), .ZN(n9041) );
  INV_X1 U7843 ( .A(n14120), .ZN(n8803) );
  INV_X1 U7844 ( .A(n8438), .ZN(n10707) );
  OR2_X1 U7845 ( .A1(n8432), .A2(n13655), .ZN(n7822) );
  NOR2_X1 U7846 ( .A1(n7824), .A2(n11466), .ZN(n7823) );
  INV_X1 U7847 ( .A(n8431), .ZN(n7824) );
  NAND2_X1 U7848 ( .A1(n16294), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8431) );
  NAND2_X1 U7849 ( .A1(n13751), .A2(n8368), .ZN(n8367) );
  NAND2_X1 U7850 ( .A1(n9222), .A2(n8369), .ZN(n8368) );
  INV_X1 U7851 ( .A(n13776), .ZN(n8369) );
  AND2_X1 U7852 ( .A1(n9195), .A2(n9194), .ZN(n13744) );
  NAND2_X1 U7853 ( .A1(n7744), .A2(n7743), .ZN(n9253) );
  AND2_X1 U7854 ( .A1(n8723), .A2(n12817), .ZN(n7743) );
  AOI21_X1 U7855 ( .B1(n13910), .B2(n7728), .A(n7516), .ZN(n7727) );
  INV_X1 U7856 ( .A(n9245), .ZN(n7728) );
  NAND2_X1 U7857 ( .A1(n9031), .A2(n12932), .ZN(n13909) );
  INV_X1 U7858 ( .A(n8396), .ZN(n8395) );
  OAI22_X1 U7859 ( .A1(n9235), .A2(n8397), .B1(n16273), .B2(n12031), .ZN(n8396) );
  NAND2_X1 U7860 ( .A1(n16053), .A2(n9226), .ZN(n16098) );
  NAND2_X1 U7861 ( .A1(n8203), .A2(n8202), .ZN(n13768) );
  AND2_X1 U7862 ( .A1(n13771), .A2(n8204), .ZN(n8202) );
  INV_X1 U7863 ( .A(n7626), .ZN(n7625) );
  OAI21_X1 U7864 ( .B1(n8191), .B2(n13858), .A(n12952), .ZN(n7626) );
  NAND2_X1 U7865 ( .A1(n12850), .A2(n8258), .ZN(n13785) );
  OR2_X1 U7866 ( .A1(n13814), .A2(n9256), .ZN(n8377) );
  NAND2_X1 U7867 ( .A1(n9135), .A2(n12861), .ZN(n13812) );
  NAND2_X1 U7868 ( .A1(n13826), .A2(n9134), .ZN(n9135) );
  NAND2_X1 U7870 ( .A1(n16051), .A2(n12868), .ZN(n8213) );
  NAND2_X1 U7871 ( .A1(n7462), .A2(n8652), .ZN(n8400) );
  NAND2_X1 U7872 ( .A1(n9164), .A2(n8768), .ZN(n9175) );
  XNOR2_X1 U7873 ( .A(n9275), .B(P3_IR_REG_26__SCAN_IN), .ZN(n9285) );
  NAND3_X1 U7874 ( .A1(n8227), .A2(n7694), .A3(n8758), .ZN(n9105) );
  INV_X1 U7875 ( .A(n9102), .ZN(n7694) );
  NAND2_X1 U7876 ( .A1(n9077), .A2(n9076), .ZN(n8756) );
  INV_X1 U7877 ( .A(n7709), .ZN(n7708) );
  NAND2_X1 U7878 ( .A1(n14122), .A2(n14123), .ZN(n8469) );
  INV_X1 U7879 ( .A(n14206), .ZN(n8460) );
  OAI21_X1 U7880 ( .B1(n8482), .B2(n8474), .A(n8481), .ZN(n8473) );
  NAND2_X1 U7881 ( .A1(n8512), .A2(n8511), .ZN(n11688) );
  AND2_X1 U7882 ( .A1(n11517), .A2(n11514), .ZN(n8511) );
  NOR2_X1 U7883 ( .A1(n11818), .A2(n8479), .ZN(n8478) );
  INV_X1 U7884 ( .A(n11814), .ZN(n8479) );
  AND4_X1 U7885 ( .A1(n13330), .A2(n13329), .A3(n13328), .A4(n13327), .ZN(
        n14355) );
  AND2_X1 U7886 ( .A1(n13107), .A2(n13106), .ZN(n14345) );
  AND2_X1 U7887 ( .A1(n9639), .A2(n12848), .ZN(n9744) );
  AND2_X1 U7888 ( .A1(n10397), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7737) );
  XNOR2_X1 U7889 ( .A(n14633), .B(n14251), .ZN(n13442) );
  NOR2_X1 U7890 ( .A1(n11270), .A2(n11269), .ZN(n7800) );
  NOR2_X1 U7891 ( .A1(n13434), .A2(n7789), .ZN(n7788) );
  INV_X1 U7892 ( .A(n11248), .ZN(n7789) );
  NAND2_X1 U7893 ( .A1(n10553), .A2(n7443), .ZN(n7808) );
  NAND2_X1 U7894 ( .A1(n7443), .A2(n13429), .ZN(n7807) );
  INV_X1 U7895 ( .A(n7614), .ZN(n7615) );
  XNOR2_X1 U7896 ( .A(n9637), .B(P2_IR_REG_30__SCAN_IN), .ZN(n9639) );
  NAND2_X1 U7897 ( .A1(n9636), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9637) );
  INV_X1 U7898 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9404) );
  INV_X1 U7899 ( .A(n14795), .ZN(n7646) );
  NAND2_X1 U7900 ( .A1(n12123), .A2(n12122), .ZN(n12124) );
  NAND2_X1 U7901 ( .A1(n12124), .A2(n12125), .ZN(n12200) );
  INV_X1 U7902 ( .A(n8554), .ZN(n8553) );
  OAI21_X1 U7903 ( .B1(n14748), .B2(n8555), .A(n14758), .ZN(n8554) );
  NAND2_X1 U7904 ( .A1(n14835), .A2(n11234), .ZN(n12484) );
  AND4_X1 U7905 ( .A1(n10118), .A2(n10117), .A3(n10116), .A4(n10115), .ZN(
        n12561) );
  NAND2_X1 U7906 ( .A1(n14992), .A2(n14837), .ZN(n8356) );
  NOR2_X1 U7907 ( .A1(n14980), .A2(n8082), .ZN(n8081) );
  INV_X1 U7908 ( .A(n13053), .ZN(n8082) );
  NAND2_X1 U7909 ( .A1(n15014), .A2(n15013), .ZN(n13052) );
  NAND2_X1 U7910 ( .A1(n13052), .A2(n8665), .ZN(n14998) );
  NOR2_X1 U7911 ( .A1(n15007), .A2(n8666), .ZN(n8665) );
  INV_X1 U7912 ( .A(n13051), .ZN(n8666) );
  AOI21_X1 U7913 ( .B1(n15025), .B2(n8328), .A(n7514), .ZN(n8327) );
  INV_X1 U7914 ( .A(n13066), .ZN(n8328) );
  NAND2_X1 U7915 ( .A1(n8357), .A2(n8358), .ZN(n15041) );
  AOI21_X1 U7916 ( .B1(n8359), .B2(n15076), .A(n7481), .ZN(n8358) );
  NAND2_X1 U7917 ( .A1(n12005), .A2(n12738), .ZN(n12007) );
  OAI21_X1 U7918 ( .B1(n11394), .B2(n7680), .A(n7518), .ZN(n11598) );
  INV_X1 U7919 ( .A(n8656), .ZN(n7680) );
  NAND2_X1 U7920 ( .A1(n7679), .A2(n8656), .ZN(n7678) );
  OAI21_X1 U7921 ( .B1(n11097), .B2(n7676), .A(n7453), .ZN(n10984) );
  NAND2_X1 U7922 ( .A1(n14857), .A2(n12544), .ZN(n7675) );
  INV_X1 U7923 ( .A(n11097), .ZN(n7673) );
  NAND2_X1 U7924 ( .A1(n7674), .A2(n12544), .ZN(n10868) );
  AND2_X1 U7925 ( .A1(n16158), .A2(n16369), .ZN(n16190) );
  NAND2_X1 U7926 ( .A1(n12505), .A2(n12307), .ZN(n12692) );
  NAND2_X1 U7927 ( .A1(n7975), .A2(n7974), .ZN(n10015) );
  NAND2_X1 U7928 ( .A1(n7976), .A2(n8169), .ZN(n7974) );
  NAND2_X1 U7929 ( .A1(n10014), .A2(n7973), .ZN(n7975) );
  NAND2_X1 U7930 ( .A1(n12297), .A2(n8428), .ZN(n12474) );
  AND2_X1 U7931 ( .A1(n8429), .A2(n12296), .ZN(n8428) );
  INV_X1 U7932 ( .A(n12471), .ZN(n8429) );
  OAI21_X1 U7933 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n15694), .A(n15693), .ZN(
        n15754) );
  OAI21_X1 U7934 ( .B1(n13471), .B2(n13595), .A(n13470), .ZN(n8063) );
  NAND3_X1 U7935 ( .A1(n7884), .A2(n7885), .A3(n8057), .ZN(n11303) );
  OR2_X1 U7936 ( .A1(n11392), .A2(n8873), .ZN(n9152) );
  NAND2_X1 U7937 ( .A1(n13380), .A2(n13379), .ZN(n14569) );
  NOR2_X1 U7938 ( .A1(n7497), .A2(n8496), .ZN(n7611) );
  NAND2_X1 U7939 ( .A1(n8498), .A2(n8497), .ZN(n8496) );
  INV_X1 U7940 ( .A(n9825), .ZN(n8498) );
  INV_X1 U7941 ( .A(n14401), .ZN(n14580) );
  NAND2_X1 U7942 ( .A1(n12426), .A2(n12425), .ZN(n15147) );
  NAND2_X1 U7943 ( .A1(n12509), .A2(n12508), .ZN(n15115) );
  NAND2_X1 U7944 ( .A1(n14922), .A2(n7687), .ZN(n15116) );
  OAI21_X1 U7945 ( .B1(n14939), .B2(n8718), .A(n14933), .ZN(n7687) );
  NAND2_X1 U7946 ( .A1(n8663), .A2(n8662), .ZN(n14922) );
  INV_X1 U7947 ( .A(n14939), .ZN(n8663) );
  AND2_X1 U7948 ( .A1(n7958), .A2(n7957), .ZN(n15876) );
  NAND2_X1 U7949 ( .A1(n12574), .A2(n12573), .ZN(n12579) );
  NAND2_X1 U7950 ( .A1(n8535), .A2(n12582), .ZN(n8534) );
  NAND2_X1 U7951 ( .A1(n13360), .A2(n14268), .ZN(n7798) );
  NAND2_X1 U7952 ( .A1(n14268), .A2(n13349), .ZN(n13118) );
  OAI21_X1 U7953 ( .B1(n8094), .B2(n13147), .A(n7529), .ZN(n8093) );
  NAND2_X1 U7954 ( .A1(n7565), .A2(n13158), .ZN(n7862) );
  INV_X1 U7955 ( .A(n13158), .ZN(n7864) );
  INV_X1 U7956 ( .A(n7565), .ZN(n7865) );
  NAND2_X1 U7957 ( .A1(n13180), .A2(n13179), .ZN(n8100) );
  INV_X1 U7958 ( .A(n13180), .ZN(n8101) );
  AND2_X1 U7959 ( .A1(n12626), .A2(n7920), .ZN(n7919) );
  INV_X1 U7960 ( .A(n12624), .ZN(n7920) );
  NAND2_X1 U7961 ( .A1(n8532), .A2(n12622), .ZN(n8531) );
  INV_X1 U7962 ( .A(n12623), .ZN(n8532) );
  NOR2_X1 U7963 ( .A1(n7464), .A2(n8120), .ZN(n8119) );
  AOI21_X1 U7964 ( .B1(n13192), .B2(n13191), .A(n13190), .ZN(n13194) );
  AND2_X1 U7965 ( .A1(n13207), .A2(n13206), .ZN(n8699) );
  NAND2_X1 U7966 ( .A1(n12632), .A2(n8526), .ZN(n8525) );
  NAND2_X1 U7967 ( .A1(n12634), .A2(n7936), .ZN(n7935) );
  AND2_X1 U7968 ( .A1(n7483), .A2(n7933), .ZN(n7932) );
  AND2_X1 U7969 ( .A1(n7937), .A2(n7935), .ZN(n7933) );
  NOR2_X1 U7970 ( .A1(n12634), .A2(n7936), .ZN(n7937) );
  INV_X1 U7971 ( .A(n13219), .ZN(n8095) );
  AND2_X1 U7972 ( .A1(n8710), .A2(n8709), .ZN(n8707) );
  AOI21_X1 U7973 ( .B1(n8708), .B2(n8705), .A(n8704), .ZN(n8703) );
  INV_X1 U7974 ( .A(n13241), .ZN(n8704) );
  INV_X1 U7975 ( .A(n8710), .ZN(n8705) );
  AND2_X1 U7976 ( .A1(n13237), .A2(n8712), .ZN(n8711) );
  OAI22_X1 U7977 ( .A1(n14493), .A2(n13341), .B1(n14345), .B2(n13360), .ZN(
        n13242) );
  NAND2_X1 U7978 ( .A1(n7922), .A2(n7921), .ZN(n12667) );
  AOI21_X1 U7979 ( .B1(n7923), .B2(n7588), .A(n7437), .ZN(n7921) );
  INV_X1 U7980 ( .A(n7757), .ZN(n7756) );
  OAI21_X1 U7981 ( .B1(n9464), .B2(n7758), .A(n9484), .ZN(n7757) );
  INV_X1 U7982 ( .A(n9467), .ZN(n7758) );
  NAND2_X1 U7983 ( .A1(n11412), .A2(n9223), .ZN(n9229) );
  NAND2_X1 U7984 ( .A1(n8104), .A2(n8105), .ZN(n8103) );
  AND2_X1 U7985 ( .A1(n8111), .A2(n7562), .ZN(n8104) );
  NAND2_X1 U7986 ( .A1(n7850), .A2(n13261), .ZN(n8105) );
  INV_X1 U7987 ( .A(n8107), .ZN(n8106) );
  OAI21_X1 U7988 ( .B1(n13290), .B2(n8108), .A(n13289), .ZN(n8107) );
  NAND2_X1 U7989 ( .A1(n8110), .A2(n7449), .ZN(n8108) );
  AND2_X1 U7990 ( .A1(n7852), .A2(n8110), .ZN(n7851) );
  INV_X1 U7991 ( .A(n13303), .ZN(n8683) );
  INV_X1 U7992 ( .A(n11946), .ZN(n8296) );
  INV_X1 U7993 ( .A(n12300), .ZN(n8427) );
  AOI21_X1 U7994 ( .B1(n8135), .B2(n8140), .A(n8133), .ZN(n8132) );
  OR2_X1 U7995 ( .A1(n10912), .A2(n8134), .ZN(n8131) );
  INV_X1 U7996 ( .A(n11320), .ZN(n8133) );
  AND2_X1 U7997 ( .A1(n8151), .A2(n10783), .ZN(n8150) );
  NAND2_X1 U7998 ( .A1(n10776), .A2(n8152), .ZN(n8151) );
  NAND2_X1 U7999 ( .A1(n10522), .A2(n10521), .ZN(n10524) );
  NAND2_X1 U8000 ( .A1(n7910), .A2(n7912), .ZN(n7763) );
  NAND2_X1 U8001 ( .A1(n15669), .A2(n8576), .ZN(n15670) );
  NAND2_X1 U8002 ( .A1(n8577), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n8576) );
  INV_X1 U8003 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n8577) );
  OAI21_X1 U8004 ( .B1(n13501), .B2(n13498), .A(n13497), .ZN(n12819) );
  OAI21_X1 U8005 ( .B1(n12795), .B2(n8648), .A(n12802), .ZN(n8647) );
  NAND2_X1 U8006 ( .A1(n8649), .A2(n7499), .ZN(n7886) );
  INV_X1 U8007 ( .A(n12157), .ZN(n7887) );
  NAND2_X1 U8008 ( .A1(n8027), .A2(n8026), .ZN(n7819) );
  NAND2_X1 U8009 ( .A1(n13676), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8026) );
  OR2_X1 U8010 ( .A1(n14068), .A2(n13848), .ZN(n12957) );
  INV_X1 U8011 ( .A(n13797), .ZN(n13795) );
  INV_X1 U8012 ( .A(n13862), .ZN(n13837) );
  INV_X1 U8013 ( .A(n8194), .ZN(n8193) );
  OAI21_X1 U8014 ( .B1(n13893), .B2(n8195), .A(n13876), .ZN(n8194) );
  NAND2_X1 U8015 ( .A1(n13621), .A2(n8848), .ZN(n12870) );
  NAND2_X1 U8016 ( .A1(n9125), .A2(n9124), .ZN(n7720) );
  AND2_X1 U8017 ( .A1(n9210), .A2(n9204), .ZN(n9207) );
  INV_X1 U8018 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9204) );
  NAND2_X1 U8019 ( .A1(n8238), .A2(n8243), .ZN(n8237) );
  AND2_X1 U8020 ( .A1(n8238), .A2(n8242), .ZN(n8236) );
  OAI21_X1 U8021 ( .B1(n8965), .B2(n7714), .A(n7712), .ZN(n7715) );
  INV_X1 U8022 ( .A(n7713), .ZN(n7712) );
  INV_X1 U8023 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n8735) );
  INV_X1 U8024 ( .A(n8734), .ZN(n8233) );
  INV_X1 U8025 ( .A(n8232), .ZN(n8231) );
  OAI21_X1 U8026 ( .B1(n8901), .B2(n8233), .A(n8918), .ZN(n8232) );
  INV_X1 U8027 ( .A(n10027), .ZN(n8508) );
  INV_X1 U8028 ( .A(n8510), .ZN(n8509) );
  INV_X1 U8029 ( .A(n10615), .ZN(n8506) );
  INV_X1 U8030 ( .A(n14186), .ZN(n8455) );
  NOR2_X1 U8031 ( .A1(n14563), .A2(n8275), .ZN(n8274) );
  INV_X1 U8032 ( .A(n8276), .ZN(n8275) );
  NOR2_X1 U8033 ( .A1(n14446), .A2(n14427), .ZN(n8264) );
  NAND2_X1 U8034 ( .A1(n14463), .A2(n14437), .ZN(n8609) );
  XNOR2_X1 U8035 ( .A(n14446), .B(n14456), .ZN(n8312) );
  INV_X1 U8036 ( .A(n11948), .ZN(n8295) );
  NAND2_X1 U8037 ( .A1(n11828), .A2(n7814), .ZN(n7813) );
  OR2_X1 U8038 ( .A1(n11826), .A2(n13439), .ZN(n11828) );
  NOR2_X1 U8039 ( .A1(n7782), .A2(n7779), .ZN(n7778) );
  INV_X1 U8040 ( .A(n13436), .ZN(n7779) );
  NAND2_X1 U8041 ( .A1(n8293), .A2(n7457), .ZN(n8292) );
  AOI21_X1 U8042 ( .B1(n13429), .B2(n8594), .A(n7527), .ZN(n8593) );
  INV_X1 U8043 ( .A(n10537), .ZN(n8594) );
  NAND2_X1 U8044 ( .A1(n10536), .A2(n8592), .ZN(n7787) );
  AND2_X1 U8045 ( .A1(n13429), .A2(n10535), .ZN(n8592) );
  INV_X1 U8046 ( .A(n8056), .ZN(n7613) );
  NOR2_X1 U8047 ( .A1(n9415), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n9495) );
  NAND2_X1 U8048 ( .A1(n14845), .A2(n8541), .ZN(n12379) );
  NAND2_X1 U8049 ( .A1(n14852), .A2(n8541), .ZN(n11726) );
  NAND2_X1 U8050 ( .A1(n14848), .A2(n8541), .ZN(n12201) );
  NAND2_X1 U8051 ( .A1(n10157), .A2(n12547), .ZN(n11965) );
  AND2_X1 U8052 ( .A1(n15076), .A2(n13044), .ZN(n8677) );
  INV_X1 U8053 ( .A(n11578), .ZN(n8350) );
  AOI21_X1 U8054 ( .B1(n8339), .B2(n8337), .A(n7543), .ZN(n8336) );
  INV_X1 U8055 ( .A(n8339), .ZN(n8338) );
  NAND2_X1 U8056 ( .A1(n7544), .A2(n12553), .ZN(n8331) );
  NOR2_X1 U8057 ( .A1(n14862), .A2(n16031), .ZN(n12546) );
  NAND2_X1 U8058 ( .A1(n8187), .A2(n10859), .ZN(n16144) );
  NOR2_X1 U8059 ( .A1(n9850), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n7658) );
  NOR2_X1 U8060 ( .A1(n12697), .A2(n8413), .ZN(n8412) );
  INV_X1 U8061 ( .A(n12695), .ZN(n8413) );
  NAND2_X1 U8062 ( .A1(n12507), .A2(n12506), .ZN(n12505) );
  INV_X1 U8063 ( .A(n7970), .ZN(n7968) );
  OAI21_X1 U8064 ( .B1(n10524), .B2(n10775), .A(n8150), .ZN(n11002) );
  NAND2_X1 U8065 ( .A1(n8143), .A2(n9770), .ZN(n9867) );
  OAI21_X1 U8066 ( .B1(n9515), .B2(n7912), .A(n7910), .ZN(n9769) );
  INV_X1 U8067 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9524) );
  INV_X1 U8068 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n15635) );
  OR2_X1 U8069 ( .A1(n9468), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9526) );
  AOI21_X1 U8070 ( .B1(n9445), .B2(n8080), .A(n7531), .ZN(n8078) );
  NAND2_X1 U8071 ( .A1(n9381), .A2(n9380), .ZN(n9386) );
  XNOR2_X1 U8072 ( .A(n15672), .B(n15673), .ZN(n15723) );
  OAI21_X1 U8073 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(n15678), .A(n15677), .ZN(
        n15710) );
  NAND2_X1 U8074 ( .A1(n15684), .A2(n15683), .ZN(n15741) );
  OR2_X1 U8075 ( .A1(n15738), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n15683) );
  OAI21_X1 U8076 ( .B1(n15686), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n15685), .ZN(
        n15688) );
  OR2_X1 U8077 ( .A1(n15740), .A2(n15741), .ZN(n15685) );
  NAND2_X1 U8078 ( .A1(n15894), .A2(n15893), .ZN(n8564) );
  NAND2_X1 U8079 ( .A1(n13466), .A2(n12835), .ZN(n7901) );
  INV_X1 U8080 ( .A(n11859), .ZN(n8644) );
  INV_X1 U8081 ( .A(n11853), .ZN(n8641) );
  NAND2_X1 U8082 ( .A1(n16057), .A2(n16055), .ZN(n16051) );
  AND2_X1 U8083 ( .A1(n13490), .A2(n8635), .ZN(n7893) );
  NAND2_X1 U8084 ( .A1(n8627), .A2(n7428), .ZN(n8630) );
  AND2_X1 U8085 ( .A1(n12805), .A2(n13525), .ZN(n8024) );
  OR2_X1 U8086 ( .A1(n13579), .A2(n13580), .ZN(n7894) );
  AND2_X1 U8087 ( .A1(n7877), .A2(n7875), .ZN(n13585) );
  NAND2_X1 U8088 ( .A1(n7876), .A2(n12833), .ZN(n7875) );
  INV_X1 U8089 ( .A(n13507), .ZN(n7876) );
  OAI211_X1 U8090 ( .C1(n12975), .C2(n12960), .A(n7705), .B(n13017), .ZN(n7704) );
  NAND2_X1 U8091 ( .A1(n7540), .A2(n12960), .ZN(n7705) );
  AND4_X1 U8092 ( .A1(n9062), .A2(n9061), .A3(n9060), .A4(n9059), .ZN(n12807)
         );
  OR2_X1 U8093 ( .A1(n12988), .A2(n8813), .ZN(n8817) );
  OR2_X1 U8094 ( .A1(n9041), .A2(n16070), .ZN(n8815) );
  NAND2_X1 U8095 ( .A1(n10327), .A2(n10064), .ZN(n10065) );
  XNOR2_X1 U8096 ( .A(n10498), .B(n10497), .ZN(n10297) );
  NOR2_X1 U8097 ( .A1(n10506), .A2(n7525), .ZN(n10511) );
  OR2_X1 U8098 ( .A1(n8903), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n8920) );
  NOR2_X1 U8099 ( .A1(n10574), .A2(n8896), .ZN(n10709) );
  AND2_X1 U8100 ( .A1(n7834), .A2(n7484), .ZN(n11124) );
  AND2_X1 U8101 ( .A1(n8442), .A2(n8441), .ZN(n11120) );
  NAND2_X1 U8102 ( .A1(n10958), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8281) );
  NOR2_X1 U8103 ( .A1(n11454), .A2(n7576), .ZN(n13654) );
  NOR2_X1 U8104 ( .A1(n7826), .A2(n11995), .ZN(n7821) );
  NOR2_X1 U8105 ( .A1(n13647), .A2(n13646), .ZN(n7978) );
  NAND2_X1 U8106 ( .A1(n7819), .A2(n7818), .ZN(n8447) );
  NAND2_X1 U8107 ( .A1(n8016), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8448) );
  AND2_X1 U8108 ( .A1(n12946), .A2(n12947), .ZN(n13876) );
  NAND2_X1 U8109 ( .A1(n13894), .A2(n13893), .ZN(n13892) );
  AND4_X1 U8110 ( .A1(n9075), .A2(n9074), .A3(n9073), .A4(n9072), .ZN(n13900)
         );
  AOI21_X1 U8111 ( .B1(n8198), .B2(n8201), .A(n7597), .ZN(n8196) );
  INV_X1 U8112 ( .A(n12920), .ZN(n8201) );
  NOR2_X1 U8113 ( .A1(n8384), .A2(n16312), .ZN(n8385) );
  NAND2_X1 U8114 ( .A1(n16312), .A2(n8384), .ZN(n8383) );
  NAND2_X1 U8115 ( .A1(n8392), .A2(n8393), .ZN(n7723) );
  NAND2_X1 U8116 ( .A1(n7479), .A2(n9237), .ZN(n8397) );
  NAND2_X1 U8117 ( .A1(n7633), .A2(n12907), .ZN(n12027) );
  NAND2_X1 U8118 ( .A1(n7632), .A2(n7490), .ZN(n7633) );
  INV_X1 U8119 ( .A(n12901), .ZN(n7631) );
  NAND2_X1 U8120 ( .A1(n7632), .A2(n12901), .ZN(n11803) );
  AOI21_X1 U8121 ( .B1(n13006), .B2(n7622), .A(n7621), .ZN(n7620) );
  INV_X1 U8122 ( .A(n12886), .ZN(n7622) );
  INV_X1 U8123 ( .A(n12891), .ZN(n7621) );
  NAND2_X1 U8124 ( .A1(n16098), .A2(n16099), .ZN(n8386) );
  OR2_X1 U8125 ( .A1(n9041), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8838) );
  AOI21_X1 U8126 ( .B1(n8205), .B2(n9160), .A(n12852), .ZN(n8204) );
  NAND2_X1 U8127 ( .A1(n13814), .A2(n8375), .ZN(n8370) );
  AOI21_X1 U8128 ( .B1(n8375), .B2(n9256), .A(n7513), .ZN(n8374) );
  NOR2_X1 U8129 ( .A1(n13797), .A2(n8376), .ZN(n8375) );
  INV_X1 U8130 ( .A(n8378), .ZN(n8376) );
  NAND2_X1 U8131 ( .A1(n8377), .A2(n8378), .ZN(n13798) );
  NAND2_X1 U8132 ( .A1(n7744), .A2(n12817), .ZN(n13835) );
  OR2_X1 U8133 ( .A1(n12961), .A2(n12962), .ZN(n13834) );
  AOI21_X1 U8134 ( .B1(n8193), .B2(n8195), .A(n8192), .ZN(n8191) );
  INV_X1 U8135 ( .A(n12947), .ZN(n8192) );
  NAND2_X1 U8136 ( .A1(n13894), .A2(n8193), .ZN(n7627) );
  INV_X1 U8137 ( .A(n16107), .ZN(n16054) );
  AND2_X1 U8138 ( .A1(n9007), .A2(n9006), .ZN(n9242) );
  INV_X1 U8139 ( .A(n12156), .ZN(n14031) );
  INV_X1 U8140 ( .A(n13615), .ZN(n12031) );
  NAND2_X1 U8141 ( .A1(n10462), .A2(n12974), .ZN(n16103) );
  NAND2_X1 U8142 ( .A1(n9236), .A2(n9235), .ZN(n11673) );
  AND2_X1 U8143 ( .A1(n9220), .A2(n9302), .ZN(n16178) );
  NAND2_X1 U8144 ( .A1(n8985), .A2(n8065), .ZN(n8823) );
  NAND2_X1 U8145 ( .A1(n9289), .A2(n9288), .ZN(n10457) );
  OR2_X1 U8146 ( .A1(n9500), .A2(P3_D_REG_0__SCAN_IN), .ZN(n9289) );
  OAI22_X1 U8147 ( .A1(n12977), .A2(n12976), .B1(P2_DATAO_REG_29__SCAN_IN), 
        .B2(n13364), .ZN(n12979) );
  NAND2_X1 U8148 ( .A1(n9150), .A2(n8766), .ZN(n9162) );
  OAI21_X1 U8149 ( .B1(n9136), .B2(n13294), .A(n8216), .ZN(n9148) );
  NAND2_X1 U8150 ( .A1(n9105), .A2(n8760), .ZN(n9117) );
  NAND2_X1 U8151 ( .A1(n8225), .A2(n13096), .ZN(n8224) );
  NOR2_X1 U8152 ( .A1(n8223), .A2(n7603), .ZN(n8222) );
  NAND2_X1 U8153 ( .A1(n8756), .A2(n8755), .ZN(n8757) );
  INV_X1 U8154 ( .A(n9207), .ZN(n9213) );
  AND2_X1 U8155 ( .A1(n9203), .A2(n9202), .ZN(n9210) );
  NAND2_X1 U8156 ( .A1(n8226), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8225) );
  INV_X1 U8157 ( .A(n8755), .ZN(n8226) );
  NAND2_X1 U8158 ( .A1(n8754), .A2(n8753), .ZN(n9077) );
  NAND2_X1 U8159 ( .A1(n9065), .A2(n8752), .ZN(n8754) );
  NOR2_X1 U8160 ( .A1(n9066), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n9203) );
  OAI21_X1 U8161 ( .B1(n9033), .B2(n7698), .A(n7695), .ZN(n9065) );
  AOI21_X1 U8162 ( .B1(n7699), .B2(n7697), .A(n7696), .ZN(n7695) );
  INV_X1 U8163 ( .A(n7699), .ZN(n7698) );
  INV_X1 U8164 ( .A(n8751), .ZN(n7696) );
  INV_X1 U8165 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8778) );
  NAND2_X1 U8166 ( .A1(n8744), .A2(n8745), .ZN(n8990) );
  AND2_X1 U8167 ( .A1(n8239), .A2(n8244), .ZN(n8238) );
  NAND2_X1 U8168 ( .A1(n8245), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n8244) );
  NAND2_X1 U8169 ( .A1(n7575), .A2(n8240), .ZN(n8239) );
  INV_X1 U8170 ( .A(n8742), .ZN(n8245) );
  INV_X1 U8171 ( .A(n7575), .ZN(n8243) );
  NAND2_X1 U8172 ( .A1(n7711), .A2(n8741), .ZN(n8978) );
  NAND2_X1 U8173 ( .A1(n8965), .A2(n8964), .ZN(n7711) );
  INV_X1 U8174 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n8736) );
  XNOR2_X1 U8175 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n8918) );
  NAND2_X1 U8176 ( .A1(n8733), .A2(n8732), .ZN(n8902) );
  NAND2_X1 U8177 ( .A1(n8217), .A2(n7451), .ZN(n8733) );
  XNOR2_X1 U8178 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n8901) );
  NAND2_X1 U8179 ( .A1(n8856), .A2(n8775), .ZN(n8389) );
  XNOR2_X1 U8180 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8854) );
  XNOR2_X1 U8181 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8842) );
  AND2_X1 U8182 ( .A1(n9631), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8820) );
  XNOR2_X1 U8183 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8821) );
  NAND2_X1 U8184 ( .A1(n8821), .A2(n8820), .ZN(n8819) );
  NOR2_X1 U8185 ( .A1(n10404), .A2(n10400), .ZN(n8510) );
  INV_X1 U8186 ( .A(n14173), .ZN(n8490) );
  INV_X1 U8187 ( .A(n14174), .ZN(n8491) );
  AOI21_X1 U8188 ( .B1(n8459), .B2(n8463), .A(n7435), .ZN(n8457) );
  INV_X1 U8189 ( .A(n14200), .ZN(n7619) );
  NAND2_X1 U8190 ( .A1(n12147), .A2(n12148), .ZN(n12236) );
  NAND2_X1 U8191 ( .A1(n8450), .A2(n14136), .ZN(n8449) );
  NAND2_X1 U8192 ( .A1(n8465), .A2(n8468), .ZN(n8464) );
  NAND2_X1 U8193 ( .A1(n14124), .A2(n8469), .ZN(n8467) );
  NAND2_X1 U8194 ( .A1(n11141), .A2(n11142), .ZN(n11506) );
  NAND2_X1 U8195 ( .A1(n12237), .A2(n12238), .ZN(n12274) );
  AND2_X1 U8196 ( .A1(n10202), .A2(n9634), .ZN(n14195) );
  AOI21_X1 U8197 ( .B1(n8478), .B2(n11815), .A(n11957), .ZN(n8477) );
  AND2_X1 U8198 ( .A1(n13090), .A2(n13350), .ZN(n9670) );
  NAND2_X1 U8199 ( .A1(n8415), .A2(n8129), .ZN(n8127) );
  NAND2_X1 U8200 ( .A1(n8421), .A2(n8420), .ZN(n8419) );
  AOI21_X1 U8201 ( .B1(n13403), .B2(n8418), .A(n8417), .ZN(n8416) );
  OAI22_X1 U8202 ( .A1(n8713), .A2(n13317), .B1(n13332), .B2(n13331), .ZN(
        n8130) );
  OR2_X1 U8203 ( .A1(n13320), .A2(n8714), .ZN(n8713) );
  INV_X1 U8204 ( .A(n13461), .ZN(n8122) );
  INV_X1 U8205 ( .A(n9567), .ZN(n7733) );
  INV_X1 U8206 ( .A(n15814), .ZN(n7735) );
  XNOR2_X1 U8207 ( .A(n12216), .B(n15836), .ZN(n15833) );
  NOR2_X1 U8208 ( .A1(n12215), .A2(n7748), .ZN(n12216) );
  AND2_X1 U8209 ( .A1(n12221), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7748) );
  NOR2_X1 U8210 ( .A1(n15833), .A2(n15832), .ZN(n15831) );
  NAND2_X1 U8211 ( .A1(n8299), .A2(n8154), .ZN(n8153) );
  AOI21_X1 U8212 ( .B1(n14405), .B2(n8155), .A(n14368), .ZN(n8154) );
  NOR2_X1 U8213 ( .A1(n8301), .A2(n8156), .ZN(n8155) );
  INV_X1 U8214 ( .A(n14407), .ZN(n8156) );
  NAND2_X1 U8215 ( .A1(n14367), .A2(n14368), .ZN(n8069) );
  NAND2_X1 U8216 ( .A1(n8585), .A2(n8586), .ZN(n14367) );
  INV_X1 U8217 ( .A(n14366), .ZN(n8070) );
  NAND2_X1 U8218 ( .A1(n7436), .A2(n7804), .ZN(n7803) );
  INV_X1 U8219 ( .A(n8297), .ZN(n7805) );
  NAND2_X1 U8220 ( .A1(n8590), .A2(n7476), .ZN(n8589) );
  NAND2_X1 U8221 ( .A1(n14393), .A2(n8591), .ZN(n8590) );
  NAND2_X1 U8222 ( .A1(n14653), .A2(n13315), .ZN(n8310) );
  AOI22_X1 U8223 ( .A1(n14421), .A2(n14422), .B1(n14427), .B2(n14440), .ZN(
        n14405) );
  NAND2_X1 U8224 ( .A1(n14405), .A2(n14407), .ZN(n14404) );
  OR2_X1 U8225 ( .A1(n14446), .A2(n14456), .ZN(n8055) );
  OR2_X1 U8226 ( .A1(n8318), .A2(n8315), .ZN(n8314) );
  INV_X1 U8227 ( .A(n8321), .ZN(n8315) );
  AND2_X1 U8228 ( .A1(n14464), .A2(n8319), .ZN(n8318) );
  NAND2_X1 U8229 ( .A1(n8320), .A2(n7439), .ZN(n8319) );
  NAND2_X1 U8230 ( .A1(n8321), .A2(n7439), .ZN(n8316) );
  INV_X1 U8231 ( .A(n8312), .ZN(n14436) );
  NAND2_X1 U8232 ( .A1(n14476), .A2(n14487), .ZN(n8322) );
  AOI21_X1 U8233 ( .B1(n8604), .B2(n14346), .A(n8602), .ZN(n8601) );
  INV_X1 U8234 ( .A(n14348), .ZN(n8602) );
  AOI21_X1 U8235 ( .B1(n14482), .B2(n14328), .A(n7594), .ZN(n14478) );
  NOR2_X1 U8236 ( .A1(n14609), .A2(n14345), .ZN(n8605) );
  NAND2_X1 U8237 ( .A1(n8608), .A2(n8607), .ZN(n8606) );
  INV_X1 U8238 ( .A(n14483), .ZN(n8608) );
  NAND2_X1 U8239 ( .A1(n14504), .A2(n8003), .ZN(n14482) );
  NAND2_X1 U8240 ( .A1(n14667), .A2(n14524), .ZN(n8003) );
  AOI21_X1 U8241 ( .B1(n14528), .B2(n14342), .A(n14341), .ZN(n14498) );
  NAND2_X1 U8242 ( .A1(n7812), .A2(n7814), .ZN(n12043) );
  OR2_X1 U8243 ( .A1(n11828), .A2(n7816), .ZN(n7812) );
  NAND2_X1 U8244 ( .A1(n11828), .A2(n11827), .ZN(n11834) );
  NAND2_X1 U8245 ( .A1(n11834), .A2(n13441), .ZN(n11947) );
  NAND2_X1 U8246 ( .A1(n11762), .A2(n13436), .ZN(n7783) );
  OR2_X1 U8247 ( .A1(n11274), .A2(n11267), .ZN(n11275) );
  NAND2_X1 U8248 ( .A1(n11247), .A2(n11246), .ZN(n7790) );
  AOI21_X1 U8249 ( .B1(n10586), .B2(n7811), .A(n7508), .ZN(n7810) );
  INV_X1 U8250 ( .A(n10552), .ZN(n7811) );
  NAND2_X1 U8251 ( .A1(n10536), .A2(n10535), .ZN(n8595) );
  AND2_X1 U8252 ( .A1(n9901), .A2(n9906), .ZN(n13423) );
  NAND2_X1 U8253 ( .A1(n7424), .A2(n9891), .ZN(n10659) );
  INV_X1 U8254 ( .A(n14438), .ZN(n14521) );
  INV_X1 U8255 ( .A(n13423), .ZN(n10660) );
  NAND2_X1 U8256 ( .A1(n13343), .A2(n13342), .ZN(n14311) );
  NAND2_X1 U8257 ( .A1(n11924), .A2(n11923), .ZN(n14633) );
  NAND2_X1 U8258 ( .A1(n10799), .A2(n10798), .ZN(n13183) );
  NAND2_X1 U8259 ( .A1(n10555), .A2(n10554), .ZN(n16269) );
  INV_X1 U8260 ( .A(n8691), .ZN(n8689) );
  INV_X1 U8261 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n9335) );
  OR2_X1 U8262 ( .A1(n9541), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n9542) );
  NAND2_X1 U8263 ( .A1(n9625), .A2(n9624), .ZN(n13421) );
  NOR2_X1 U8264 ( .A1(n9620), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n7841) );
  INV_X1 U8265 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n9627) );
  NOR2_X2 U8266 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n9403) );
  AND2_X1 U8267 ( .A1(n10734), .A2(n10732), .ZN(n8015) );
  INV_X1 U8268 ( .A(n12483), .ZN(n12520) );
  NAND2_X1 U8269 ( .A1(n14776), .A2(n7455), .ZN(n8017) );
  INV_X1 U8270 ( .A(n14731), .ZN(n7965) );
  NAND2_X1 U8271 ( .A1(n14815), .A2(n14819), .ZN(n14747) );
  NAND2_X1 U8272 ( .A1(n14747), .A2(n14748), .ZN(n14746) );
  NAND2_X1 U8273 ( .A1(n14837), .A2(n8541), .ZN(n12449) );
  NAND2_X1 U8274 ( .A1(n12200), .A2(n12199), .ZN(n12207) );
  NAND2_X1 U8275 ( .A1(n7985), .A2(n7984), .ZN(n7647) );
  INV_X1 U8276 ( .A(n14784), .ZN(n7984) );
  NAND2_X1 U8277 ( .A1(n11981), .A2(n8558), .ZN(n12123) );
  AND2_X1 U8278 ( .A1(n11982), .A2(n11980), .ZN(n8558) );
  OR2_X1 U8279 ( .A1(n12470), .A2(n12469), .ZN(n8550) );
  NAND2_X1 U8280 ( .A1(n14846), .A2(n8541), .ZN(n12372) );
  NAND2_X1 U8281 ( .A1(n12362), .A2(n8560), .ZN(n14706) );
  AND2_X1 U8282 ( .A1(n14707), .A2(n12361), .ZN(n8560) );
  NAND2_X1 U8283 ( .A1(n14706), .A2(n8559), .ZN(n14817) );
  AND2_X1 U8284 ( .A1(n12377), .A2(n12371), .ZN(n8559) );
  NAND2_X1 U8285 ( .A1(n14817), .A2(n14816), .ZN(n14815) );
  AND4_X1 U8286 ( .A1(n11559), .A2(n11558), .A3(n11557), .A4(n11556), .ZN(
        n12606) );
  AND2_X1 U8287 ( .A1(n10083), .A2(n10082), .ZN(n10084) );
  NAND2_X1 U8288 ( .A1(n12526), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n10091) );
  NAND2_X1 U8289 ( .A1(n8540), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8170) );
  NAND2_X1 U8290 ( .A1(n8168), .A2(n8167), .ZN(n8166) );
  NAND2_X1 U8291 ( .A1(n12701), .A2(n12700), .ZN(n14911) );
  AND2_X1 U8292 ( .A1(n12525), .A2(n12513), .ZN(n14927) );
  AND2_X1 U8293 ( .A1(n14970), .A2(n8356), .ZN(n8352) );
  INV_X1 U8294 ( .A(n15138), .ZN(n14992) );
  NAND2_X1 U8295 ( .A1(n15006), .A2(n13069), .ZN(n14985) );
  NAND2_X1 U8296 ( .A1(n15039), .A2(n8674), .ZN(n15027) );
  AND2_X1 U8297 ( .A1(n15028), .A2(n13049), .ZN(n8674) );
  OAI21_X1 U8298 ( .B1(n13045), .B2(n7685), .A(n7683), .ZN(n13048) );
  AND2_X1 U8299 ( .A1(n7684), .A2(n15056), .ZN(n7683) );
  OR2_X1 U8300 ( .A1(n8677), .A2(n7685), .ZN(n7684) );
  INV_X1 U8301 ( .A(n13046), .ZN(n7685) );
  NAND2_X1 U8302 ( .A1(n13045), .A2(n8677), .ZN(n15071) );
  NAND2_X1 U8303 ( .A1(n8362), .A2(n8361), .ZN(n15073) );
  INV_X1 U8304 ( .A(n15075), .ZN(n8362) );
  OAI21_X1 U8305 ( .B1(n12252), .B2(n12743), .A(n12253), .ZN(n12255) );
  NAND2_X1 U8306 ( .A1(n12247), .A2(n8678), .ZN(n13045) );
  NOR2_X1 U8307 ( .A1(n12254), .A2(n8679), .ZN(n8678) );
  INV_X1 U8308 ( .A(n12246), .ZN(n8679) );
  OAI21_X1 U8309 ( .B1(n12007), .B2(n8670), .A(n7681), .ZN(n12245) );
  INV_X1 U8310 ( .A(n7682), .ZN(n7681) );
  OAI21_X1 U8311 ( .B1(n8671), .B2(n8670), .A(n12173), .ZN(n7682) );
  NAND2_X1 U8312 ( .A1(n12007), .A2(n8671), .ZN(n12080) );
  NAND2_X1 U8313 ( .A1(n12004), .A2(n12003), .ZN(n14705) );
  INV_X1 U8314 ( .A(n12738), .ZN(n11783) );
  NAND2_X1 U8315 ( .A1(n11784), .A2(n11783), .ZN(n12001) );
  NAND2_X1 U8316 ( .A1(n11788), .A2(n11787), .ZN(n12005) );
  NAND2_X1 U8317 ( .A1(n11598), .A2(n11549), .ZN(n16320) );
  NOR2_X1 U8318 ( .A1(n8658), .A2(n12731), .ZN(n8654) );
  AOI21_X1 U8320 ( .B1(n12733), .B2(n8657), .A(n7511), .ZN(n8656) );
  INV_X1 U8321 ( .A(n11374), .ZN(n8657) );
  NAND2_X1 U8322 ( .A1(n11373), .A2(n11372), .ZN(n11394) );
  NAND2_X1 U8323 ( .A1(n11394), .A2(n7429), .ZN(n11396) );
  NAND2_X1 U8324 ( .A1(n11049), .A2(n12728), .ZN(n8341) );
  AND2_X1 U8325 ( .A1(n10859), .A2(n16162), .ZN(n7657) );
  NAND2_X1 U8326 ( .A1(n10864), .A2(n10863), .ZN(n11097) );
  NAND2_X1 U8327 ( .A1(n12353), .A2(n12352), .ZN(n15184) );
  INV_X1 U8328 ( .A(n16194), .ZN(n16379) );
  INV_X1 U8329 ( .A(n16158), .ZN(n16372) );
  AND2_X1 U8330 ( .A1(n11553), .A2(n11552), .ZN(n16324) );
  AND2_X1 U8331 ( .A1(n9695), .A2(n9694), .ZN(n10144) );
  INV_X1 U8332 ( .A(n8412), .ZN(n8411) );
  AOI21_X1 U8333 ( .B1(n8412), .B2(n8410), .A(n8409), .ZN(n8408) );
  INV_X1 U8334 ( .A(n12707), .ZN(n8409) );
  INV_X1 U8335 ( .A(n12691), .ZN(n8410) );
  NAND2_X1 U8336 ( .A1(n10104), .A2(n7969), .ZN(n9354) );
  NOR2_X1 U8337 ( .A1(n7507), .A2(n7970), .ZN(n7969) );
  INV_X1 U8338 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8542) );
  OR2_X1 U8339 ( .A1(n12457), .A2(n12456), .ZN(n12297) );
  NAND2_X1 U8340 ( .A1(n11718), .A2(n11717), .ZN(n12293) );
  NOR2_X1 U8341 ( .A1(n10914), .A2(n8136), .ZN(n8135) );
  INV_X1 U8342 ( .A(n8138), .ZN(n8136) );
  NAND2_X1 U8343 ( .A1(n10912), .A2(n8139), .ZN(n8137) );
  NAND2_X1 U8344 ( .A1(n10911), .A2(n15280), .ZN(n8138) );
  OR2_X1 U8345 ( .A1(n10528), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n10757) );
  AND2_X1 U8346 ( .A1(n9875), .A2(n9774), .ZN(n11781) );
  XNOR2_X1 U8347 ( .A(n9867), .B(n9865), .ZN(n11780) );
  XNOR2_X1 U8348 ( .A(n9503), .B(n9504), .ZN(n11362) );
  NAND2_X1 U8349 ( .A1(n9424), .A2(n9423), .ZN(n8079) );
  NOR2_X1 U8350 ( .A1(n15715), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n15717) );
  XNOR2_X1 U8351 ( .A(n15723), .B(n15674), .ZN(n15724) );
  NAND2_X1 U8352 ( .A1(n8573), .A2(n15726), .ZN(n15727) );
  NAND2_X1 U8353 ( .A1(n8570), .A2(n15735), .ZN(n15736) );
  NAND2_X1 U8354 ( .A1(n15917), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n8570) );
  OR2_X1 U8355 ( .A1(n15869), .A2(n15868), .ZN(n7960) );
  AOI21_X1 U8356 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n15692), .A(n15691), .ZN(
        n15750) );
  NOR2_X1 U8357 ( .A1(n15746), .A2(n15745), .ZN(n15691) );
  AOI22_X1 U8358 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(n15928), .B1(n15754), 
        .B2(n15696), .ZN(n15757) );
  NOR2_X1 U8359 ( .A1(n15897), .A2(n15766), .ZN(n15770) );
  NAND2_X1 U8360 ( .A1(n15774), .A2(n15902), .ZN(n8567) );
  INV_X1 U8361 ( .A(n11294), .ZN(n9281) );
  NOR2_X1 U8362 ( .A1(n7898), .A2(n13608), .ZN(n7896) );
  NOR2_X1 U8363 ( .A1(n7899), .A2(n7902), .ZN(n7898) );
  NOR2_X1 U8364 ( .A1(n13466), .A2(n12835), .ZN(n7902) );
  INV_X1 U8365 ( .A(n7901), .ZN(n7899) );
  NAND2_X1 U8366 ( .A1(n7901), .A2(n8626), .ZN(n7900) );
  NAND2_X1 U8367 ( .A1(n13585), .A2(n13586), .ZN(n13584) );
  NAND2_X1 U8368 ( .A1(n8631), .A2(n8630), .ZN(n10461) );
  AND3_X1 U8369 ( .A1(n9133), .A2(n9132), .A3(n9131), .ZN(n13838) );
  AND2_X1 U8370 ( .A1(n11304), .A2(n11302), .ZN(n7883) );
  NAND2_X1 U8371 ( .A1(n7623), .A2(n13032), .ZN(n8212) );
  NAND2_X1 U8372 ( .A1(n7624), .A2(n7503), .ZN(n7623) );
  OAI211_X1 U8373 ( .C1(n7704), .C2(n8254), .A(n8251), .B(n7703), .ZN(n7702)
         );
  INV_X1 U8374 ( .A(n8255), .ZN(n8254) );
  AND2_X1 U8375 ( .A1(n8252), .A2(n8256), .ZN(n8251) );
  NAND2_X1 U8376 ( .A1(n7704), .A2(n8246), .ZN(n7703) );
  INV_X1 U8377 ( .A(n8256), .ZN(n8250) );
  AOI21_X1 U8378 ( .B1(n13761), .B2(n9201), .A(n9200), .ZN(n13776) );
  OR2_X1 U8379 ( .A1(n12992), .A2(n8388), .ZN(n7639) );
  OR2_X1 U8380 ( .A1(n11455), .A2(n16317), .ZN(n8285) );
  INV_X1 U8381 ( .A(n8279), .ZN(n15985) );
  OR2_X1 U8382 ( .A1(n15979), .A2(n15980), .ZN(n8436) );
  OR2_X1 U8383 ( .A1(n8447), .A2(n13694), .ZN(n8444) );
  OR2_X1 U8384 ( .A1(n13677), .A2(n8445), .ZN(n8443) );
  NAND2_X1 U8385 ( .A1(n8446), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8445) );
  INV_X1 U8386 ( .A(n13694), .ZN(n8446) );
  NOR2_X1 U8387 ( .A1(n13712), .A2(n8287), .ZN(n8286) );
  AND2_X1 U8388 ( .A1(n13713), .A2(n13721), .ZN(n8287) );
  OAI21_X1 U8389 ( .B1(n13715), .B2(n8289), .A(n15931), .ZN(n8288) );
  AND2_X1 U8390 ( .A1(n13711), .A2(n13710), .ZN(n8289) );
  AND2_X1 U8391 ( .A1(n8448), .A2(n8447), .ZN(n13695) );
  XNOR2_X1 U8392 ( .A(n8060), .B(n8059), .ZN(n13731) );
  INV_X1 U8393 ( .A(n13725), .ZN(n8059) );
  NAND2_X1 U8394 ( .A1(n8443), .A2(n7817), .ZN(n8060) );
  AND2_X1 U8395 ( .A1(n8444), .A2(n7610), .ZN(n7817) );
  AND2_X1 U8396 ( .A1(n9956), .A2(n9955), .ZN(n15966) );
  OAI21_X1 U8397 ( .B1(n15984), .B2(n13733), .A(n8050), .ZN(n8049) );
  INV_X1 U8398 ( .A(n13730), .ZN(n8050) );
  NAND2_X1 U8399 ( .A1(n9038), .A2(n9037), .ZN(n13918) );
  NOR2_X1 U8400 ( .A1(n8036), .A2(n14018), .ZN(n8035) );
  NAND2_X1 U8401 ( .A1(n9177), .A2(n9176), .ZN(n14042) );
  NAND2_X1 U8402 ( .A1(n8208), .A2(n9258), .ZN(n8207) );
  INV_X1 U8403 ( .A(n13796), .ZN(n8208) );
  NAND2_X1 U8404 ( .A1(n9107), .A2(n9106), .ZN(n14074) );
  NAND2_X1 U8405 ( .A1(n9094), .A2(n9093), .ZN(n14080) );
  NAND2_X1 U8406 ( .A1(n9056), .A2(n9055), .ZN(n14089) );
  NAND2_X1 U8407 ( .A1(n8791), .A2(n7506), .ZN(n14113) );
  INV_X1 U8408 ( .A(n8400), .ZN(n8791) );
  INV_X1 U8409 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n14112) );
  NAND2_X1 U8410 ( .A1(n8801), .A2(n8792), .ZN(n13037) );
  NAND2_X1 U8411 ( .A1(n9162), .A2(n9161), .ZN(n9164) );
  INV_X1 U8412 ( .A(SI_20_), .ZN(n15280) );
  INV_X1 U8413 ( .A(n14437), .ZN(n14350) );
  OR2_X1 U8414 ( .A1(n14179), .A2(n7473), .ZN(n8489) );
  AND2_X1 U8415 ( .A1(n8486), .A2(n14232), .ZN(n8485) );
  INV_X1 U8416 ( .A(n8487), .ZN(n8486) );
  OAI21_X1 U8417 ( .B1(n8489), .B2(n8492), .A(n8488), .ZN(n8487) );
  NAND2_X1 U8418 ( .A1(n14179), .A2(n7473), .ZN(n8488) );
  OR2_X1 U8419 ( .A1(n14240), .A2(n14241), .ZN(n14238) );
  NAND2_X1 U8420 ( .A1(n8500), .A2(n8499), .ZN(n9826) );
  INV_X1 U8421 ( .A(n8501), .ZN(n8499) );
  INV_X1 U8422 ( .A(n14493), .ZN(n14609) );
  NAND2_X1 U8423 ( .A1(n11688), .A2(n7616), .ZN(n11816) );
  OR2_X1 U8424 ( .A1(n11689), .A2(n11690), .ZN(n7616) );
  NAND2_X1 U8425 ( .A1(n13265), .A2(n13264), .ZN(n14599) );
  OR2_X1 U8426 ( .A1(n13262), .A2(n13321), .ZN(n13265) );
  OR2_X1 U8427 ( .A1(n13378), .A2(n9721), .ZN(n9722) );
  NOR2_X1 U8428 ( .A1(n7611), .A2(n7519), .ZN(n10028) );
  NAND2_X1 U8429 ( .A1(n10028), .A2(n10027), .ZN(n10402) );
  AND3_X1 U8430 ( .A1(n11842), .A2(n11841), .A3(n11840), .ZN(n13226) );
  NAND2_X1 U8431 ( .A1(n11833), .A2(n11832), .ZN(n13221) );
  OAI21_X1 U8432 ( .B1(n8130), .B2(n8124), .A(n8121), .ZN(n8688) );
  INV_X1 U8433 ( .A(n8125), .ZN(n8124) );
  AOI21_X1 U8434 ( .B1(n8125), .B2(n8123), .A(n8122), .ZN(n8121) );
  AND2_X1 U8435 ( .A1(n8127), .A2(n7609), .ZN(n8125) );
  INV_X1 U8436 ( .A(n14355), .ZN(n14330) );
  INV_X1 U8437 ( .A(n13215), .ZN(n14253) );
  AND3_X1 U8438 ( .A1(n9641), .A2(n9643), .A3(n9640), .ZN(n7971) );
  NOR2_X1 U8439 ( .A1(n9580), .A2(n9579), .ZN(n9578) );
  NOR2_X1 U8440 ( .A1(n11643), .A2(n11642), .ZN(n12215) );
  AOI21_X1 U8441 ( .B1(n14562), .B2(n16306), .A(n14364), .ZN(n8615) );
  XNOR2_X1 U8442 ( .A(n14331), .B(n14359), .ZN(n14566) );
  INV_X1 U8443 ( .A(n8617), .ZN(n8039) );
  XNOR2_X1 U8444 ( .A(n14360), .B(n14359), .ZN(n7773) );
  AOI21_X1 U8445 ( .B1(n14363), .B2(n14438), .A(n8618), .ZN(n8617) );
  AND2_X1 U8446 ( .A1(n13323), .A2(n13322), .ZN(n14401) );
  NAND2_X1 U8447 ( .A1(n11927), .A2(n11926), .ZN(n14336) );
  OAI21_X1 U8448 ( .B1(n16350), .B2(n7457), .A(n8293), .ZN(n11905) );
  NAND2_X1 U8449 ( .A1(n11245), .A2(n11244), .ZN(n13197) );
  NAND2_X1 U8450 ( .A1(n11136), .A2(n11135), .ZN(n16304) );
  NAND2_X1 U8451 ( .A1(n10582), .A2(n10586), .ZN(n10581) );
  NAND2_X1 U8452 ( .A1(n10553), .A2(n10552), .ZN(n10582) );
  NAND2_X1 U8453 ( .A1(n15784), .A2(n9629), .ZN(n14510) );
  AND2_X2 U8454 ( .A1(n9897), .A2(n9896), .ZN(n16358) );
  NOR2_X1 U8455 ( .A1(n8691), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n8690) );
  AND2_X1 U8456 ( .A1(n9698), .A2(n9700), .ZN(n9356) );
  INV_X1 U8457 ( .A(n8176), .ZN(n8175) );
  AND2_X1 U8458 ( .A1(n8174), .A2(n8547), .ZN(n8173) );
  NAND2_X1 U8459 ( .A1(n8176), .A2(n8179), .ZN(n8174) );
  OAI21_X1 U8460 ( .B1(n14756), .B2(n7646), .A(n7536), .ZN(n14721) );
  OR2_X1 U8461 ( .A1(n12396), .A2(n12397), .ZN(n8163) );
  OR2_X1 U8462 ( .A1(n14760), .A2(n7646), .ZN(n7645) );
  NAND2_X1 U8463 ( .A1(n12401), .A2(n12400), .ZN(n15174) );
  OAI21_X1 U8464 ( .B1(n14738), .B2(n8543), .A(n8544), .ZN(n7966) );
  AOI21_X1 U8465 ( .B1(n7524), .B2(n8547), .A(n8545), .ZN(n8544) );
  NAND2_X1 U8466 ( .A1(n7548), .A2(n8180), .ZN(n8543) );
  NOR2_X1 U8467 ( .A1(n12504), .A2(n12503), .ZN(n8545) );
  NAND2_X1 U8468 ( .A1(n12327), .A2(n12326), .ZN(n15159) );
  AOI21_X1 U8469 ( .B1(n14768), .B2(n14769), .A(n7440), .ZN(n14738) );
  INV_X1 U8470 ( .A(n15049), .ZN(n15169) );
  OR2_X1 U8471 ( .A1(n15255), .A2(n8724), .ZN(n12476) );
  NAND2_X1 U8472 ( .A1(n8551), .A2(n8550), .ZN(n14805) );
  OAI21_X1 U8473 ( .B1(n14768), .B2(n7440), .A(n8178), .ZN(n8551) );
  INV_X1 U8474 ( .A(n12606), .ZN(n14850) );
  NAND4_X1 U8475 ( .A1(n10877), .A2(n10876), .A3(n10875), .A4(n10874), .ZN(
        n14856) );
  AND2_X1 U8476 ( .A1(n12539), .A2(n12538), .ZN(n15108) );
  XNOR2_X1 U8477 ( .A(n13074), .B(n13056), .ZN(n15111) );
  OR2_X1 U8478 ( .A1(n15115), .A2(n14699), .ZN(n13072) );
  AOI21_X1 U8479 ( .B1(n14940), .B2(n8662), .A(n8660), .ZN(n8659) );
  OAI21_X1 U8480 ( .B1(n7465), .B2(n8661), .A(n13055), .ZN(n8660) );
  OR2_X1 U8481 ( .A1(n14983), .A2(n14982), .ZN(n15142) );
  NAND2_X1 U8482 ( .A1(n14998), .A2(n13053), .ZN(n14981) );
  NOR2_X1 U8483 ( .A1(n15114), .A2(n7581), .ZN(n8089) );
  INV_X1 U8484 ( .A(n15113), .ZN(n8366) );
  OR2_X1 U8485 ( .A1(n7951), .A2(n15717), .ZN(n7950) );
  AND2_X1 U8486 ( .A1(n15715), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n7951) );
  AOI21_X1 U8487 ( .B1(n7468), .B2(n7955), .A(n15744), .ZN(n15874) );
  NAND2_X1 U8488 ( .A1(n7468), .A2(n7954), .ZN(n8575) );
  NOR2_X1 U8489 ( .A1(n15870), .A2(n7956), .ZN(n7954) );
  INV_X1 U8490 ( .A(n15744), .ZN(n7956) );
  AOI21_X1 U8491 ( .B1(n15748), .B2(n15747), .A(n15876), .ZN(n15881) );
  AND2_X1 U8492 ( .A1(n7964), .A2(n7963), .ZN(n15890) );
  NAND2_X1 U8493 ( .A1(n15755), .A2(n15756), .ZN(n7963) );
  NAND2_X1 U8494 ( .A1(n8567), .A2(n8568), .ZN(n7942) );
  NAND2_X1 U8495 ( .A1(n15771), .A2(n15772), .ZN(n15773) );
  INV_X1 U8496 ( .A(n15908), .ZN(n7945) );
  NAND2_X1 U8497 ( .A1(n7940), .A2(n7939), .ZN(n15909) );
  NAND2_X1 U8498 ( .A1(n15771), .A2(n7941), .ZN(n7940) );
  NAND2_X1 U8499 ( .A1(n8567), .A2(n8568), .ZN(n7939) );
  NOR2_X1 U8500 ( .A1(n8566), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n7941) );
  OR2_X1 U8501 ( .A1(n12553), .A2(n12551), .ZN(n7989) );
  AOI21_X1 U8502 ( .B1(n12564), .B2(n12563), .A(n12726), .ZN(n7996) );
  NAND2_X1 U8503 ( .A1(n7991), .A2(n12581), .ZN(n7990) );
  INV_X1 U8504 ( .A(n12582), .ZN(n7991) );
  OAI211_X1 U8505 ( .C1(n13122), .C2(n14268), .A(n13121), .B(n7798), .ZN(
        n13123) );
  AND2_X1 U8506 ( .A1(n13126), .A2(n13125), .ZN(n13131) );
  AND2_X1 U8507 ( .A1(n13113), .A2(n13112), .ZN(n13136) );
  MUX2_X1 U8508 ( .A(n14850), .B(n16338), .S(n12551), .Z(n12608) );
  AND2_X1 U8509 ( .A1(n8700), .A2(n7863), .ZN(n7860) );
  OR2_X1 U8510 ( .A1(n13162), .A2(n13163), .ZN(n8700) );
  NOR2_X1 U8511 ( .A1(n8520), .A2(n8519), .ZN(n8518) );
  NOR2_X1 U8512 ( .A1(n8520), .A2(n12605), .ZN(n8517) );
  AND2_X1 U8513 ( .A1(n13187), .A2(n8100), .ZN(n8099) );
  NOR2_X1 U8514 ( .A1(n7500), .A2(n7845), .ZN(n7844) );
  INV_X1 U8515 ( .A(n13186), .ZN(n7845) );
  NAND2_X1 U8516 ( .A1(n8533), .A2(n12623), .ZN(n8530) );
  INV_X1 U8517 ( .A(n12622), .ZN(n8533) );
  NAND2_X1 U8518 ( .A1(n7846), .A2(n7843), .ZN(n13192) );
  NAND2_X1 U8519 ( .A1(n7848), .A2(n7847), .ZN(n7846) );
  NAND2_X1 U8520 ( .A1(n8098), .A2(n7844), .ZN(n7843) );
  NOR2_X1 U8521 ( .A1(n13187), .A2(n7542), .ZN(n7847) );
  NAND2_X1 U8522 ( .A1(n7916), .A2(n7918), .ZN(n12630) );
  AND2_X1 U8523 ( .A1(n12631), .A2(n7917), .ZN(n7914) );
  NAND2_X1 U8524 ( .A1(n7919), .A2(n7918), .ZN(n7917) );
  INV_X1 U8525 ( .A(n12633), .ZN(n8526) );
  NOR2_X1 U8526 ( .A1(n7868), .A2(n8698), .ZN(n7867) );
  AND2_X1 U8527 ( .A1(n8119), .A2(n8118), .ZN(n7868) );
  NAND2_X1 U8528 ( .A1(n8697), .A2(n8699), .ZN(n8696) );
  OAI21_X1 U8529 ( .B1(n8699), .B2(n8113), .A(n8697), .ZN(n8112) );
  NAND2_X1 U8530 ( .A1(n8118), .A2(n8119), .ZN(n8113) );
  NOR2_X1 U8531 ( .A1(n8699), .A2(n8117), .ZN(n8116) );
  NOR2_X1 U8532 ( .A1(n7438), .A2(n7932), .ZN(n7931) );
  NAND2_X1 U8533 ( .A1(n13224), .A2(n13225), .ZN(n8694) );
  AOI21_X1 U8534 ( .B1(n13220), .B2(n13219), .A(n13218), .ZN(n8693) );
  INV_X1 U8535 ( .A(n12650), .ZN(n8019) );
  INV_X1 U8536 ( .A(n12653), .ZN(n7930) );
  AND2_X1 U8537 ( .A1(n12653), .A2(n7929), .ZN(n7928) );
  NAND2_X1 U8538 ( .A1(n7836), .A2(n8702), .ZN(n13243) );
  INV_X1 U8539 ( .A(n8708), .ZN(n8706) );
  NOR2_X1 U8540 ( .A1(n7509), .A2(n7924), .ZN(n7923) );
  NOR2_X1 U8541 ( .A1(n7925), .A2(n12660), .ZN(n7924) );
  NOR2_X1 U8542 ( .A1(n13785), .A2(n13795), .ZN(n12854) );
  NAND2_X1 U8543 ( .A1(n7857), .A2(n7856), .ZN(n7855) );
  OR2_X1 U8544 ( .A1(n7449), .A2(n7858), .ZN(n7857) );
  OR2_X1 U8545 ( .A1(n7449), .A2(n13259), .ZN(n7856) );
  OR2_X1 U8546 ( .A1(n7449), .A2(n7853), .ZN(n7852) );
  INV_X1 U8547 ( .A(n8135), .ZN(n8134) );
  INV_X1 U8548 ( .A(n10523), .ZN(n8152) );
  NOR2_X1 U8549 ( .A1(n10241), .A2(n8425), .ZN(n8424) );
  INV_X1 U8550 ( .A(n9870), .ZN(n8425) );
  INV_X1 U8551 ( .A(n9239), .ZN(n7726) );
  INV_X1 U8552 ( .A(n7725), .ZN(n7724) );
  OAI21_X1 U8553 ( .B1(n8393), .B2(n7726), .A(n8383), .ZN(n7725) );
  INV_X1 U8554 ( .A(n8375), .ZN(n8372) );
  INV_X1 U8555 ( .A(n8374), .ZN(n8373) );
  INV_X1 U8556 ( .A(n8741), .ZN(n7714) );
  OAI21_X1 U8557 ( .B1(n8964), .B2(n7714), .A(n8977), .ZN(n7713) );
  INV_X1 U8558 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9714) );
  INV_X1 U8559 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9518) );
  NAND2_X1 U8560 ( .A1(n14574), .A2(n14356), .ZN(n8308) );
  NOR2_X1 U8561 ( .A1(n11827), .A2(n7816), .ZN(n7815) );
  NOR2_X1 U8562 ( .A1(n14569), .A2(n14574), .ZN(n8276) );
  NOR2_X2 U8563 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n9532) );
  AOI21_X1 U8564 ( .B1(n10524), .B2(n8150), .A(n8148), .ZN(n8147) );
  NAND2_X1 U8565 ( .A1(n8149), .A2(n10785), .ZN(n8148) );
  NAND2_X1 U8566 ( .A1(n8150), .A2(n10775), .ZN(n8149) );
  INV_X1 U8567 ( .A(SI_17_), .ZN(n15477) );
  INV_X1 U8568 ( .A(n8422), .ZN(n8142) );
  AOI21_X1 U8569 ( .B1(n8424), .B2(n9866), .A(n8423), .ZN(n8422) );
  INV_X1 U8570 ( .A(n10243), .ZN(n8423) );
  INV_X1 U8571 ( .A(n8145), .ZN(n8144) );
  OAI21_X1 U8572 ( .B1(n8722), .B2(n8146), .A(n8424), .ZN(n8145) );
  INV_X1 U8573 ( .A(n9770), .ZN(n8146) );
  NAND2_X1 U8574 ( .A1(n10245), .A2(n10244), .ZN(n10523) );
  NAND2_X1 U8575 ( .A1(n9872), .A2(n9871), .ZN(n10243) );
  INV_X1 U8576 ( .A(n9711), .ZN(n7913) );
  NAND2_X1 U8577 ( .A1(n7754), .A2(n7753), .ZN(n9505) );
  AOI21_X1 U8578 ( .B1(n7756), .B2(n7758), .A(n7530), .ZN(n7753) );
  AOI21_X1 U8579 ( .B1(n9422), .B2(n9426), .A(n9444), .ZN(n8076) );
  INV_X1 U8580 ( .A(n9426), .ZN(n8080) );
  INV_X1 U8581 ( .A(n9388), .ZN(n7907) );
  OAI21_X1 U8582 ( .B1(n15714), .B2(P1_ADDR_REG_2__SCAN_IN), .A(n15671), .ZN(
        n15672) );
  INV_X1 U8583 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n15678) );
  NOR2_X1 U8584 ( .A1(n13566), .A2(n12821), .ZN(n12823) );
  XNOR2_X1 U8585 ( .A(n8825), .B(n10763), .ZN(n10458) );
  NOR2_X1 U8586 ( .A1(n8073), .A2(n8072), .ZN(n8071) );
  NOR2_X1 U8587 ( .A1(n13597), .A2(n13519), .ZN(n8072) );
  INV_X1 U8588 ( .A(n13514), .ZN(n8073) );
  NOR2_X1 U8589 ( .A1(n7879), .A2(n13508), .ZN(n7878) );
  INV_X1 U8590 ( .A(n12833), .ZN(n7879) );
  MUX2_X1 U8591 ( .A(n12858), .B(n12857), .S(n12974), .Z(n12968) );
  NAND2_X1 U8592 ( .A1(n8440), .A2(n8439), .ZN(n8438) );
  NAND2_X1 U8593 ( .A1(n10573), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8439) );
  OR2_X1 U8594 ( .A1(n8441), .A2(n11121), .ZN(n7833) );
  OR2_X1 U8595 ( .A1(n8442), .A2(n11121), .ZN(n7831) );
  NAND2_X1 U8596 ( .A1(n8442), .A2(n7832), .ZN(n7830) );
  AND2_X1 U8597 ( .A1(n11121), .A2(n8441), .ZN(n7832) );
  AOI21_X1 U8598 ( .B1(n8284), .B2(n16317), .A(n15924), .ZN(n8283) );
  NOR2_X1 U8599 ( .A1(n15962), .A2(n8280), .ZN(n13663) );
  AND2_X1 U8600 ( .A1(n15958), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8280) );
  INV_X1 U8601 ( .A(n13706), .ZN(n7818) );
  XNOR2_X1 U8602 ( .A(n13721), .B(n13698), .ZN(n13700) );
  AND2_X1 U8603 ( .A1(n9188), .A2(n9187), .ZN(n12855) );
  AND2_X1 U8604 ( .A1(n12927), .A2(n8199), .ZN(n8198) );
  NAND2_X1 U8605 ( .A1(n8200), .A2(n12920), .ZN(n8199) );
  NAND2_X1 U8606 ( .A1(n7724), .A2(n7726), .ZN(n7721) );
  INV_X1 U8607 ( .A(n9229), .ZN(n9230) );
  NAND2_X1 U8608 ( .A1(n8380), .A2(n8379), .ZN(n8378) );
  OR2_X1 U8609 ( .A1(n14058), .A2(n8379), .ZN(n12853) );
  NAND2_X1 U8610 ( .A1(n12108), .A2(n13010), .ZN(n12110) );
  INV_X1 U8611 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8788) );
  INV_X1 U8612 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8651) );
  INV_X1 U8613 ( .A(n8225), .ZN(n8223) );
  NOR2_X1 U8614 ( .A1(n9048), .A2(n7700), .ZN(n7699) );
  INV_X1 U8615 ( .A(n8749), .ZN(n7700) );
  OAI21_X1 U8616 ( .B1(n8989), .B2(n7710), .A(n9017), .ZN(n7709) );
  INV_X1 U8617 ( .A(n8977), .ZN(n8240) );
  NAND2_X1 U8618 ( .A1(n7689), .A2(n8726), .ZN(n7691) );
  AND2_X1 U8619 ( .A1(n8726), .A2(n8725), .ZN(n7688) );
  NAND2_X1 U8620 ( .A1(n8391), .A2(n8390), .ZN(n8430) );
  NAND2_X1 U8621 ( .A1(n8477), .A2(n8475), .ZN(n8474) );
  INV_X1 U8622 ( .A(n8478), .ZN(n8475) );
  NAND2_X1 U8623 ( .A1(n12144), .A2(n12145), .ZN(n8481) );
  NAND2_X1 U8624 ( .A1(n12146), .A2(n8477), .ZN(n8476) );
  INV_X1 U8625 ( .A(n9739), .ZN(n8502) );
  NAND2_X1 U8626 ( .A1(n13449), .A2(n13404), .ZN(n8418) );
  AND2_X1 U8627 ( .A1(n13408), .A2(n13409), .ZN(n8417) );
  INV_X1 U8628 ( .A(n13406), .ZN(n8421) );
  INV_X1 U8629 ( .A(n13405), .ZN(n8420) );
  AND2_X1 U8630 ( .A1(n13332), .A2(n13331), .ZN(n8714) );
  OAI21_X1 U8631 ( .B1(n8681), .B2(n7466), .A(n8680), .ZN(n13319) );
  OR2_X1 U8632 ( .A1(n8683), .A2(n13304), .ZN(n8680) );
  OR2_X1 U8633 ( .A1(n14569), .A2(n14152), .ZN(n14357) );
  NAND2_X1 U8634 ( .A1(n14574), .A2(n14180), .ZN(n8586) );
  INV_X1 U8635 ( .A(n14384), .ZN(n8587) );
  OR2_X1 U8636 ( .A1(n13281), .A2(n14159), .ZN(n13298) );
  INV_X1 U8637 ( .A(n8322), .ZN(n8320) );
  NOR2_X1 U8638 ( .A1(n7521), .A2(n7786), .ZN(n7785) );
  INV_X1 U8639 ( .A(n8593), .ZN(n7786) );
  AND2_X1 U8640 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9790) );
  OR2_X1 U8641 ( .A1(n13202), .A2(n11347), .ZN(n11907) );
  OR2_X1 U8642 ( .A1(n11263), .A2(n13197), .ZN(n11347) );
  OR3_X1 U8643 ( .A1(n14688), .A2(n14690), .A3(n11721), .ZN(n9600) );
  INV_X1 U8644 ( .A(n9532), .ZN(n9620) );
  INV_X1 U8645 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9395) );
  AND2_X1 U8646 ( .A1(n8549), .A2(n8550), .ZN(n8548) );
  NAND2_X1 U8647 ( .A1(n14855), .A2(n8541), .ZN(n11164) );
  NAND2_X1 U8648 ( .A1(n14847), .A2(n8541), .ZN(n12363) );
  NAND2_X1 U8649 ( .A1(n8537), .A2(n12672), .ZN(n8536) );
  INV_X1 U8650 ( .A(n15243), .ZN(n10080) );
  AND2_X1 U8651 ( .A1(n8169), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n8167) );
  AND2_X1 U8652 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n12510), .ZN(n12511) );
  NOR2_X1 U8653 ( .A1(n14812), .A2(n8186), .ZN(n8184) );
  OR2_X1 U8654 ( .A1(n15015), .A2(n15147), .ZN(n7669) );
  NOR2_X1 U8655 ( .A1(n15043), .A2(n15159), .ZN(n8183) );
  INV_X1 U8656 ( .A(n13062), .ZN(n8360) );
  AND2_X1 U8657 ( .A1(n12258), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n12402) );
  INV_X1 U8658 ( .A(n8654), .ZN(n7679) );
  OR2_X1 U8659 ( .A1(n11054), .A2(n11053), .ZN(n11366) );
  INV_X1 U8660 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n10883) );
  NAND2_X1 U8661 ( .A1(n10984), .A2(n10878), .ZN(n10890) );
  INV_X1 U8662 ( .A(n14835), .ZN(n14698) );
  INV_X1 U8663 ( .A(n16162), .ZN(n16143) );
  INV_X1 U8664 ( .A(n10087), .ZN(n7643) );
  NOR2_X1 U8665 ( .A1(n7976), .A2(n8169), .ZN(n7973) );
  INV_X1 U8666 ( .A(n7665), .ZN(n7659) );
  INV_X1 U8667 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9844) );
  INV_X1 U8668 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8668) );
  INV_X1 U8669 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9345) );
  NAND2_X1 U8670 ( .A1(n12303), .A2(n12302), .ZN(n12507) );
  NOR2_X1 U8671 ( .A1(n12301), .A2(n8427), .ZN(n8426) );
  NAND2_X1 U8672 ( .A1(n7549), .A2(n9347), .ZN(n7970) );
  NAND2_X1 U8673 ( .A1(n8403), .A2(n8405), .ZN(n8404) );
  INV_X1 U8674 ( .A(SI_22_), .ZN(n8405) );
  NAND2_X1 U8675 ( .A1(n11322), .A2(SI_22_), .ZN(n8407) );
  INV_X1 U8676 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n15708) );
  AOI22_X1 U8677 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n15730), .B1(n15680), .B2(
        n15731), .ZN(n15681) );
  INV_X1 U8678 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n15639) );
  NOR2_X1 U8679 ( .A1(n12825), .A2(n12824), .ZN(n13483) );
  AND2_X1 U8680 ( .A1(n12823), .A2(n12822), .ZN(n12824) );
  XNOR2_X1 U8681 ( .A(n11329), .B(n10763), .ZN(n11027) );
  AOI21_X1 U8682 ( .B1(n13466), .B2(n12835), .A(n12838), .ZN(n8625) );
  INV_X1 U8683 ( .A(n8625), .ZN(n8623) );
  INV_X1 U8684 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n10705) );
  NAND2_X1 U8685 ( .A1(n12158), .A2(n12157), .ZN(n7890) );
  AND2_X1 U8686 ( .A1(n12833), .A2(n12832), .ZN(n13507) );
  INV_X1 U8687 ( .A(n13620), .ZN(n11209) );
  INV_X1 U8688 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n15531) );
  NAND2_X1 U8689 ( .A1(n12825), .A2(n7882), .ZN(n7881) );
  NAND2_X1 U8690 ( .A1(n13483), .A2(n13838), .ZN(n13539) );
  NAND2_X1 U8691 ( .A1(n11030), .A2(n8637), .ZN(n11205) );
  INV_X1 U8692 ( .A(n11029), .ZN(n8638) );
  NAND2_X1 U8693 ( .A1(n8645), .A2(n8642), .ZN(n11896) );
  NAND2_X1 U8694 ( .A1(n11854), .A2(n11853), .ZN(n8645) );
  NAND2_X1 U8695 ( .A1(n7890), .A2(n7459), .ZN(n13557) );
  NAND2_X1 U8696 ( .A1(n7873), .A2(n7872), .ZN(n7871) );
  INV_X1 U8697 ( .A(n13944), .ZN(n13519) );
  OAI21_X1 U8698 ( .B1(n12158), .B2(n7888), .A(n7537), .ZN(n13515) );
  NAND2_X1 U8699 ( .A1(n8649), .A2(n7459), .ZN(n7888) );
  INV_X1 U8700 ( .A(n8647), .ZN(n8646) );
  NAND2_X1 U8701 ( .A1(n13024), .A2(n13023), .ZN(n7624) );
  NOR2_X1 U8702 ( .A1(n13020), .A2(n12996), .ZN(n8246) );
  AOI21_X1 U8703 ( .B1(n8255), .B2(n13020), .A(n8253), .ZN(n8252) );
  NOR2_X1 U8704 ( .A1(n13027), .A2(n12996), .ZN(n8253) );
  AND2_X1 U8705 ( .A1(n13027), .A2(n13036), .ZN(n8255) );
  OR2_X1 U8706 ( .A1(n13042), .A2(n13041), .ZN(n8256) );
  OR2_X1 U8707 ( .A1(n10272), .A2(n10271), .ZN(n10273) );
  AND2_X1 U8708 ( .A1(n10265), .A2(n10478), .ZN(n10266) );
  OR2_X1 U8709 ( .A1(n10264), .A2(n10271), .ZN(n10265) );
  NAND2_X1 U8710 ( .A1(n10274), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n10474) );
  NAND2_X1 U8711 ( .A1(n10266), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n10480) );
  XNOR2_X1 U8712 ( .A(n8438), .B(n10562), .ZN(n10574) );
  INV_X1 U8713 ( .A(n8432), .ZN(n11456) );
  XNOR2_X1 U8714 ( .A(n13658), .B(n15944), .ZN(n15946) );
  NOR2_X1 U8715 ( .A1(n13697), .A2(n13696), .ZN(n13720) );
  NAND2_X1 U8716 ( .A1(n12969), .A2(n12970), .ZN(n13752) );
  NOR2_X1 U8717 ( .A1(n13769), .A2(n7463), .ZN(n13753) );
  NOR2_X1 U8718 ( .A1(n9139), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9154) );
  NAND2_X1 U8719 ( .A1(n12861), .A2(n12862), .ZN(n13825) );
  NAND2_X1 U8720 ( .A1(n9109), .A2(n9108), .ZN(n9120) );
  AND2_X1 U8721 ( .A1(n9095), .A2(n15346), .ZN(n9109) );
  NOR2_X1 U8722 ( .A1(n9084), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9095) );
  NAND2_X1 U8723 ( .A1(n9057), .A2(n15531), .ZN(n9071) );
  AOI21_X1 U8724 ( .B1(n9247), .B2(n9246), .A(n7454), .ZN(n13886) );
  NAND2_X1 U8725 ( .A1(n13886), .A2(n13885), .ZN(n13884) );
  AND4_X1 U8726 ( .A1(n9045), .A2(n9044), .A3(n9043), .A4(n9042), .ZN(n13899)
         );
  AND2_X1 U8727 ( .A1(n9039), .A2(n13518), .ZN(n9057) );
  NAND2_X1 U8728 ( .A1(n13925), .A2(n9245), .ZN(n13911) );
  NOR2_X1 U8729 ( .A1(n9025), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9039) );
  AND2_X1 U8730 ( .A1(n12925), .A2(n9015), .ZN(n13948) );
  NAND2_X1 U8731 ( .A1(n12110), .A2(n12920), .ZN(n13962) );
  OR2_X1 U8732 ( .A1(n13947), .A2(n12793), .ZN(n13961) );
  OR2_X1 U8733 ( .A1(n8958), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8971) );
  NOR2_X1 U8734 ( .A1(n8971), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9008) );
  INV_X1 U8735 ( .A(n13612), .ZN(n13959) );
  AND2_X1 U8736 ( .A1(n12917), .A2(n12916), .ZN(n13008) );
  INV_X1 U8737 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n15536) );
  NAND2_X1 U8738 ( .A1(n8927), .A2(n15536), .ZN(n8944) );
  NOR2_X1 U8739 ( .A1(n8894), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8910) );
  NOR2_X1 U8740 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8862) );
  INV_X1 U8741 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n15338) );
  NAND2_X1 U8742 ( .A1(n7636), .A2(n13001), .ZN(n7635) );
  NAND2_X1 U8743 ( .A1(n8213), .A2(n12866), .ZN(n16100) );
  NAND2_X1 U8744 ( .A1(n16050), .A2(n9225), .ZN(n16053) );
  INV_X1 U8745 ( .A(n13624), .ZN(n16057) );
  NAND2_X1 U8746 ( .A1(n13809), .A2(n13543), .ZN(n9257) );
  NOR2_X1 U8747 ( .A1(n8262), .A2(n8873), .ZN(n8261) );
  AND2_X1 U8748 ( .A1(n12853), .A2(n12859), .ZN(n13813) );
  NAND2_X1 U8749 ( .A1(n9127), .A2(n9126), .ZN(n13482) );
  NAND2_X1 U8750 ( .A1(n9251), .A2(n9250), .ZN(n13849) );
  AND2_X1 U8751 ( .A1(n12955), .A2(n12956), .ZN(n13850) );
  AND4_X1 U8752 ( .A1(n9101), .A2(n9100), .A3(n9099), .A4(n9098), .ZN(n13847)
         );
  AND2_X1 U8753 ( .A1(n9261), .A2(n12974), .ZN(n13943) );
  INV_X1 U8754 ( .A(n16103), .ZN(n13941) );
  NAND2_X1 U8755 ( .A1(n9083), .A2(n9082), .ZN(n14001) );
  NAND2_X1 U8756 ( .A1(n11312), .A2(n12894), .ZN(n8908) );
  AND2_X1 U8757 ( .A1(n14109), .A2(n10332), .ZN(n10349) );
  AND2_X1 U8758 ( .A1(n9221), .A2(n10454), .ZN(n16200) );
  INV_X1 U8759 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8790) );
  NOR2_X1 U8760 ( .A1(n8772), .A2(n8040), .ZN(n12977) );
  AND2_X1 U8761 ( .A1(n15247), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8040) );
  MUX2_X1 U8762 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8789), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n8792) );
  NAND2_X1 U8763 ( .A1(n7462), .A2(n7628), .ZN(n8801) );
  AND2_X1 U8764 ( .A1(n8652), .A2(n8790), .ZN(n7628) );
  OAI21_X1 U8765 ( .B1(n9117), .B2(n9116), .A(n8761), .ZN(n9125) );
  XNOR2_X1 U8766 ( .A(n9274), .B(n9273), .ZN(n10331) );
  INV_X1 U8767 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9273) );
  OAI21_X1 U8768 ( .B1(n9272), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9274) );
  NAND2_X1 U8769 ( .A1(n9207), .A2(n9205), .ZN(n9272) );
  OR2_X1 U8770 ( .A1(n8979), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n8980) );
  NOR2_X1 U8771 ( .A1(n8980), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n9002) );
  NAND2_X1 U8772 ( .A1(n8740), .A2(n8739), .ZN(n8965) );
  INV_X1 U8773 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8966) );
  AOI21_X1 U8774 ( .B1(n8231), .B2(n8233), .A(n7539), .ZN(n8229) );
  XNOR2_X1 U8775 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n8938) );
  AOI21_X1 U8776 ( .B1(n8219), .B2(n8869), .A(n7538), .ZN(n8218) );
  INV_X1 U8777 ( .A(n8730), .ZN(n8219) );
  NAND2_X1 U8778 ( .A1(n8855), .A2(n7716), .ZN(n8217) );
  NOR2_X1 U8779 ( .A1(n7718), .A2(n7717), .ZN(n7716) );
  INV_X1 U8780 ( .A(n8854), .ZN(n7717) );
  INV_X1 U8781 ( .A(n8869), .ZN(n7718) );
  NAND2_X1 U8782 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n8278) );
  OR2_X1 U8783 ( .A1(n11816), .A2(n11815), .ZN(n8480) );
  NOR2_X1 U8784 ( .A1(n14175), .A2(n8493), .ZN(n8492) );
  INV_X1 U8785 ( .A(n14150), .ZN(n8493) );
  AOI21_X1 U8786 ( .B1(n8507), .B2(n8509), .A(n8506), .ZN(n8505) );
  NOR2_X1 U8787 ( .A1(n10030), .A2(n10029), .ZN(n10405) );
  AND2_X1 U8788 ( .A1(n7431), .A2(n14266), .ZN(n9725) );
  NAND2_X1 U8789 ( .A1(n8501), .A2(n9824), .ZN(n8497) );
  NAND2_X1 U8790 ( .A1(n12236), .A2(n12235), .ZN(n12237) );
  NAND2_X1 U8791 ( .A1(n9787), .A2(n9781), .ZN(n8501) );
  NAND2_X1 U8792 ( .A1(n8503), .A2(n8502), .ZN(n8500) );
  AND2_X1 U8793 ( .A1(n13100), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n13268) );
  NAND2_X1 U8794 ( .A1(n8459), .A2(n14186), .ZN(n8456) );
  OAI21_X1 U8795 ( .B1(n8457), .B2(n8455), .A(n7528), .ZN(n8454) );
  OR2_X1 U8796 ( .A1(n11507), .A2(n11508), .ZN(n8514) );
  AND2_X1 U8797 ( .A1(n11144), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n11253) );
  AND2_X1 U8798 ( .A1(n9790), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9828) );
  AND2_X1 U8799 ( .A1(n13396), .A2(n8129), .ZN(n8128) );
  INV_X1 U8800 ( .A(n8128), .ZN(n8123) );
  AND3_X1 U8801 ( .A1(n15789), .A2(P2_IR_REG_0__SCAN_IN), .A3(
        P2_REG1_REG_0__SCAN_IN), .ZN(n15790) );
  OAI21_X1 U8802 ( .B1(n15786), .B2(n9551), .A(n8041), .ZN(n15794) );
  NAND2_X1 U8803 ( .A1(n15786), .A2(n9551), .ZN(n8041) );
  AOI21_X1 U8804 ( .B1(n9562), .B2(P2_REG1_REG_1__SCAN_IN), .A(n15790), .ZN(
        n15803) );
  AOI21_X1 U8805 ( .B1(n10397), .B2(P2_REG2_REG_7__SCAN_IN), .A(n10183), .ZN(
        n15819) );
  AOI21_X1 U8806 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n11134), .A(n10842), .ZN(
        n10845) );
  NOR2_X1 U8807 ( .A1(n10845), .A2(n10844), .ZN(n11070) );
  NOR2_X1 U8808 ( .A1(n11070), .A2(n8008), .ZN(n11073) );
  AND2_X1 U8809 ( .A1(n11243), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8008) );
  NAND2_X1 U8810 ( .A1(n11073), .A2(n11072), .ZN(n11425) );
  AOI21_X1 U8811 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n11691), .A(n11632), .ZN(
        n11636) );
  OR2_X1 U8812 ( .A1(n14287), .A2(n7732), .ZN(n7731) );
  AND2_X1 U8813 ( .A1(n14288), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7732) );
  NAND2_X1 U8814 ( .A1(n9619), .A2(n9618), .ZN(n7842) );
  AND2_X1 U8815 ( .A1(n7731), .A2(n14286), .ZN(n14298) );
  NOR2_X1 U8816 ( .A1(n8273), .A2(n14310), .ZN(n8272) );
  INV_X1 U8817 ( .A(n8274), .ZN(n8273) );
  AND2_X1 U8818 ( .A1(n14361), .A2(n14362), .ZN(n8618) );
  NAND2_X1 U8819 ( .A1(n7806), .A2(n8297), .ZN(n14365) );
  AND2_X1 U8820 ( .A1(n14401), .A2(n14411), .ZN(n14396) );
  AND2_X1 U8821 ( .A1(n8263), .A2(n8264), .ZN(n14411) );
  NOR3_X1 U8822 ( .A1(n14473), .A2(n14599), .A3(n14412), .ZN(n8263) );
  NAND2_X1 U8823 ( .A1(n7797), .A2(n8311), .ZN(n14421) );
  AOI21_X1 U8824 ( .B1(n7442), .B2(n8316), .A(n7546), .ZN(n8311) );
  NAND2_X1 U8825 ( .A1(n14478), .A2(n7442), .ZN(n7797) );
  OR2_X1 U8826 ( .A1(n8597), .A2(n8598), .ZN(n8596) );
  INV_X1 U8827 ( .A(n8609), .ZN(n8597) );
  NAND2_X1 U8828 ( .A1(n7764), .A2(n14325), .ZN(n14517) );
  NAND2_X1 U8829 ( .A1(n12040), .A2(n13442), .ZN(n7784) );
  AND2_X1 U8830 ( .A1(n11943), .A2(n11942), .ZN(n14326) );
  INV_X1 U8831 ( .A(n8277), .ZN(n14535) );
  NAND2_X1 U8832 ( .A1(n12048), .A2(n13227), .ZN(n12049) );
  AND3_X1 U8833 ( .A1(n11704), .A2(n11703), .A3(n11702), .ZN(n13215) );
  OR2_X1 U8834 ( .A1(n11698), .A2(n11819), .ZN(n11765) );
  OR2_X1 U8835 ( .A1(n11338), .A2(n11705), .ZN(n11698) );
  AOI21_X1 U8836 ( .B1(n13437), .B2(n7781), .A(n7482), .ZN(n7780) );
  INV_X1 U8837 ( .A(n11763), .ZN(n7781) );
  NAND2_X1 U8838 ( .A1(n7799), .A2(n11774), .ZN(n11826) );
  OAI21_X1 U8839 ( .B1(n7800), .B2(n8294), .A(n7526), .ZN(n7799) );
  NAND2_X1 U8840 ( .A1(n11275), .A2(n11268), .ZN(n11270) );
  OAI21_X1 U8841 ( .B1(n16269), .B2(n11246), .A(n8290), .ZN(n11274) );
  AOI21_X1 U8842 ( .B1(n13433), .B2(n8291), .A(n7492), .ZN(n8290) );
  INV_X1 U8843 ( .A(n10808), .ZN(n8291) );
  NOR2_X1 U8844 ( .A1(n10800), .A2(n11151), .ZN(n11144) );
  OR2_X1 U8845 ( .A1(n10542), .A2(n10925), .ZN(n10800) );
  NAND2_X1 U8846 ( .A1(n8271), .A2(n8270), .ZN(n10813) );
  NAND2_X1 U8847 ( .A1(n7787), .A2(n8593), .ZN(n10679) );
  NAND2_X1 U8848 ( .A1(n10427), .A2(n9904), .ZN(n9905) );
  XNOR2_X1 U8849 ( .A(n13146), .B(n10218), .ZN(n13425) );
  NAND2_X1 U8850 ( .A1(n10656), .A2(n9903), .ZN(n10428) );
  INV_X1 U8851 ( .A(n10431), .ZN(n13424) );
  NAND2_X1 U8852 ( .A1(n10428), .A2(n13424), .ZN(n10427) );
  AOI22_X1 U8853 ( .A1(n10659), .A2(n7775), .B1(n9906), .B2(n7774), .ZN(n10432) );
  AND2_X1 U8854 ( .A1(n10658), .A2(n9906), .ZN(n7775) );
  INV_X1 U8855 ( .A(n9901), .ZN(n7774) );
  XNOR2_X1 U8856 ( .A(n14264), .B(n16169), .ZN(n10431) );
  NAND2_X1 U8857 ( .A1(n10432), .A2(n10431), .ZN(n10430) );
  AND2_X1 U8858 ( .A1(n9670), .A2(n9669), .ZN(n14438) );
  NAND2_X1 U8859 ( .A1(n10657), .A2(n10660), .ZN(n10656) );
  AND2_X1 U8860 ( .A1(n10283), .A2(n13121), .ZN(n10666) );
  NOR2_X1 U8861 ( .A1(n13090), .A2(n13350), .ZN(n9809) );
  NOR2_X1 U8862 ( .A1(n10087), .A2(n9419), .ZN(n7791) );
  INV_X1 U8863 ( .A(n16353), .ZN(n16170) );
  NAND2_X1 U8864 ( .A1(n9538), .A2(n9539), .ZN(n8691) );
  NAND2_X1 U8865 ( .A1(n7613), .A2(n7472), .ZN(n7614) );
  AND2_X1 U8866 ( .A1(n7472), .A2(n9538), .ZN(n7612) );
  NAND2_X1 U8867 ( .A1(n9336), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9338) );
  NAND2_X1 U8868 ( .A1(n9338), .A2(n9534), .ZN(n9340) );
  XNOR2_X1 U8869 ( .A(n9342), .B(n9535), .ZN(n11530) );
  NAND3_X1 U8870 ( .A1(n8404), .A2(n8406), .A3(n8407), .ZN(n11527) );
  INV_X1 U8871 ( .A(n11324), .ZN(n8406) );
  OR2_X1 U8872 ( .A1(n9674), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n9754) );
  OR2_X1 U8873 ( .A1(n9476), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n9492) );
  OR2_X1 U8874 ( .A1(n9450), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n9476) );
  NAND2_X1 U8875 ( .A1(n14854), .A2(n8541), .ZN(n11231) );
  AND2_X1 U8876 ( .A1(n8177), .A2(n8548), .ZN(n8176) );
  NAND2_X1 U8877 ( .A1(n8178), .A2(n7440), .ZN(n8177) );
  NOR2_X1 U8878 ( .A1(n11366), .A2(n11365), .ZN(n11376) );
  NAND2_X1 U8879 ( .A1(n10728), .A2(n10727), .ZN(n10733) );
  INV_X1 U8880 ( .A(n14697), .ZN(n8546) );
  NAND2_X1 U8881 ( .A1(n7574), .A2(n8549), .ZN(n8547) );
  NAND2_X1 U8882 ( .A1(n14853), .A2(n8541), .ZN(n11479) );
  NAND2_X1 U8883 ( .A1(n11488), .A2(n8556), .ZN(n11725) );
  NOR2_X1 U8884 ( .A1(n11491), .A2(n8557), .ZN(n8556) );
  INV_X1 U8885 ( .A(n11487), .ZN(n8557) );
  NAND2_X1 U8886 ( .A1(n12416), .A2(n8165), .ZN(n8164) );
  INV_X1 U8887 ( .A(n12417), .ZN(n8165) );
  NAND2_X1 U8888 ( .A1(n14836), .A2(n8541), .ZN(n12466) );
  NOR2_X1 U8889 ( .A1(n12185), .A2(n12184), .ZN(n12258) );
  OR2_X1 U8890 ( .A1(n12083), .A2(n12082), .ZN(n12185) );
  CLKBUF_X1 U8891 ( .A(n11965), .Z(n8012) );
  AND2_X1 U8892 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n10873) );
  OR2_X1 U8893 ( .A1(n11583), .A2(n11582), .ZN(n11790) );
  NOR2_X1 U8894 ( .A1(n12340), .A2(n14733), .ZN(n12328) );
  INV_X1 U8895 ( .A(n11975), .ZN(n7653) );
  INV_X1 U8896 ( .A(n11974), .ZN(n7654) );
  OAI22_X1 U8897 ( .A1(n10123), .A2(n10228), .B1(n16090), .B2(n11965), .ZN(
        n8171) );
  NOR2_X1 U8898 ( .A1(n11790), .A2(n11789), .ZN(n12013) );
  INV_X1 U8899 ( .A(n15263), .ZN(n12784) );
  NAND2_X1 U8900 ( .A1(n14918), .A2(n15105), .ZN(n14917) );
  INV_X1 U8901 ( .A(n14949), .ZN(n8661) );
  INV_X1 U8902 ( .A(n8718), .ZN(n8664) );
  AND2_X1 U8903 ( .A1(n15119), .A2(n13071), .ZN(n8032) );
  INV_X1 U8904 ( .A(n7465), .ZN(n8662) );
  NOR2_X1 U8905 ( .A1(n14940), .A2(n14949), .ZN(n14939) );
  OAI21_X1 U8906 ( .B1(n14698), .B2(n15126), .A(n14954), .ZN(n14940) );
  NAND2_X1 U8907 ( .A1(n15000), .A2(n8184), .ZN(n14958) );
  NAND2_X1 U8908 ( .A1(n14956), .A2(n14955), .ZN(n14954) );
  NAND2_X1 U8909 ( .A1(n14969), .A2(n8720), .ZN(n14953) );
  NAND2_X1 U8910 ( .A1(n15000), .A2(n14992), .ZN(n14991) );
  INV_X1 U8911 ( .A(n12461), .ZN(n12460) );
  NAND2_X1 U8912 ( .A1(n13068), .A2(n13067), .ZN(n15008) );
  AND2_X1 U8913 ( .A1(n15011), .A2(n8327), .ZN(n8324) );
  NAND2_X1 U8914 ( .A1(n8183), .A2(n15021), .ZN(n15015) );
  NAND2_X1 U8915 ( .A1(n15027), .A2(n13050), .ZN(n15014) );
  INV_X1 U8916 ( .A(n8183), .ZN(n15029) );
  NAND2_X1 U8917 ( .A1(n15061), .A2(n15169), .ZN(n15043) );
  NAND2_X1 U8918 ( .A1(n13048), .A2(n7491), .ZN(n15039) );
  OR2_X1 U8919 ( .A1(n15081), .A2(n15184), .ZN(n15079) );
  NOR2_X2 U8920 ( .A1(n15079), .A2(n15174), .ZN(n15061) );
  NAND2_X1 U8921 ( .A1(n12245), .A2(n12743), .ZN(n12247) );
  NAND2_X1 U8922 ( .A1(n12081), .A2(n15206), .ZN(n12182) );
  NAND2_X1 U8923 ( .A1(n7672), .A2(n7671), .ZN(n12010) );
  NOR2_X1 U8924 ( .A1(n14705), .A2(n12010), .ZN(n12081) );
  NOR2_X1 U8925 ( .A1(n11580), .A2(n8350), .ZN(n8349) );
  OR2_X1 U8926 ( .A1(n11567), .A2(n11566), .ZN(n11583) );
  AND2_X1 U8927 ( .A1(n11376), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11554) );
  NAND2_X1 U8928 ( .A1(n11554), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n11567) );
  NAND2_X1 U8929 ( .A1(n11398), .A2(n11399), .ZN(n11397) );
  NAND2_X1 U8930 ( .A1(n8335), .A2(n8336), .ZN(n11400) );
  OR2_X1 U8931 ( .A1(n11049), .A2(n8338), .ZN(n8335) );
  AND2_X1 U8932 ( .A1(n11062), .A2(n8342), .ZN(n11398) );
  NAND2_X1 U8933 ( .A1(n7670), .A2(n16208), .ZN(n10991) );
  INV_X1 U8934 ( .A(n11101), .ZN(n7670) );
  NOR2_X1 U8935 ( .A1(n10991), .A2(n12575), .ZN(n11062) );
  NAND2_X1 U8936 ( .A1(n16141), .A2(n16189), .ZN(n11101) );
  INV_X1 U8937 ( .A(n8331), .ZN(n8332) );
  NAND2_X1 U8938 ( .A1(n12556), .A2(n12553), .ZN(n10857) );
  NAND2_X1 U8939 ( .A1(n8086), .A2(n8087), .ZN(n8085) );
  INV_X1 U8940 ( .A(n16071), .ZN(n8086) );
  INV_X1 U8941 ( .A(n14785), .ZN(n14806) );
  INV_X1 U8942 ( .A(n10857), .ZN(n12725) );
  INV_X1 U8943 ( .A(n8087), .ZN(n16073) );
  INV_X1 U8944 ( .A(n12752), .ZN(n16038) );
  INV_X1 U8945 ( .A(n16142), .ZN(n16322) );
  NAND2_X1 U8946 ( .A1(n11565), .A2(n11564), .ZN(n16365) );
  NOR2_X1 U8947 ( .A1(n10150), .A2(n10145), .ZN(n10855) );
  AND2_X1 U8948 ( .A1(n12708), .A2(n12699), .ZN(n14681) );
  NAND2_X1 U8949 ( .A1(n8414), .A2(n8412), .ZN(n12708) );
  NAND2_X1 U8950 ( .A1(n8414), .A2(n12695), .ZN(n12698) );
  XNOR2_X1 U8951 ( .A(n12692), .B(n12691), .ZN(n13363) );
  OAI21_X1 U8952 ( .B1(n12507), .B2(n12506), .A(n12505), .ZN(n14683) );
  XNOR2_X1 U8953 ( .A(n7972), .B(P1_IR_REG_25__SCAN_IN), .ZN(n9700) );
  NAND2_X1 U8954 ( .A1(n9354), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7972) );
  NAND2_X1 U8955 ( .A1(n9350), .A2(n9349), .ZN(n9352) );
  INV_X1 U8956 ( .A(n9350), .ZN(n9357) );
  NAND2_X1 U8957 ( .A1(n8407), .A2(n8404), .ZN(n12314) );
  XNOR2_X1 U8958 ( .A(n11008), .B(n11007), .ZN(n13108) );
  XNOR2_X1 U8959 ( .A(n9769), .B(n8722), .ZN(n11562) );
  OR2_X1 U8960 ( .A1(n9526), .A2(n9525), .ZN(n9718) );
  NAND2_X1 U8961 ( .A1(n7909), .A2(n9517), .ZN(n9712) );
  NAND2_X1 U8962 ( .A1(n7755), .A2(n9467), .ZN(n9485) );
  NAND2_X1 U8963 ( .A1(n9465), .A2(n9464), .ZN(n7755) );
  OR2_X1 U8964 ( .A1(n9412), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n9432) );
  NAND2_X1 U8965 ( .A1(n8667), .A2(n9344), .ZN(n9389) );
  INV_X1 U8966 ( .A(n9382), .ZN(n8667) );
  NAND2_X1 U8967 ( .A1(n7908), .A2(n9388), .ZN(n8401) );
  NAND2_X1 U8968 ( .A1(n9370), .A2(n15627), .ZN(n9382) );
  AND2_X1 U8969 ( .A1(n8323), .A2(n15622), .ZN(n9370) );
  NAND2_X1 U8970 ( .A1(n9360), .A2(n9631), .ZN(n7988) );
  INV_X1 U8971 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n15715) );
  XNOR2_X1 U8972 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n15716) );
  NAND2_X1 U8973 ( .A1(n7938), .A2(n15729), .ZN(n15733) );
  NAND2_X1 U8974 ( .A1(n15867), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n7938) );
  NAND2_X1 U8975 ( .A1(n15690), .A2(n15689), .ZN(n15745) );
  NAND2_X1 U8976 ( .A1(n7953), .A2(n7952), .ZN(n7958) );
  NAND2_X1 U8977 ( .A1(n8575), .A2(n8574), .ZN(n7952) );
  INV_X1 U8978 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n8574) );
  AOI22_X1 U8979 ( .A1(n15757), .A2(n15697), .B1(P3_ADDR_REG_13__SCAN_IN), 
        .B2(n15758), .ZN(n15761) );
  NAND2_X1 U8980 ( .A1(n13558), .A2(n12798), .ZN(n13472) );
  OAI21_X1 U8981 ( .B1(n11854), .B2(n8643), .A(n8639), .ZN(n12099) );
  AND2_X1 U8982 ( .A1(n8640), .A2(n11895), .ZN(n8639) );
  NAND2_X1 U8983 ( .A1(n8642), .A2(n8641), .ZN(n8640) );
  NAND2_X1 U8984 ( .A1(n7894), .A2(n7893), .ZN(n13489) );
  AND2_X1 U8985 ( .A1(n7894), .A2(n8635), .ZN(n13491) );
  INV_X1 U8986 ( .A(n10461), .ZN(n8629) );
  NAND2_X1 U8987 ( .A1(n7890), .A2(n12161), .ZN(n12163) );
  NAND2_X1 U8988 ( .A1(n11204), .A2(n11205), .ZN(n11206) );
  NAND2_X1 U8989 ( .A1(n11030), .A2(n11029), .ZN(n11036) );
  NAND2_X1 U8990 ( .A1(n8645), .A2(n11856), .ZN(n11858) );
  INV_X1 U8991 ( .A(n13887), .ZN(n13574) );
  NAND2_X1 U8992 ( .A1(n7892), .A2(n7891), .ZN(n13550) );
  AOI21_X1 U8993 ( .B1(n7893), .B2(n13580), .A(n7541), .ZN(n7891) );
  NAND2_X1 U8994 ( .A1(n13579), .A2(n7893), .ZN(n7892) );
  NAND2_X1 U8995 ( .A1(n13557), .A2(n12795), .ZN(n13558) );
  AND3_X1 U8996 ( .A1(n7871), .A2(n12820), .A3(n13848), .ZN(n13566) );
  NAND2_X1 U8997 ( .A1(n7871), .A2(n12820), .ZN(n13567) );
  NAND2_X1 U8998 ( .A1(n10626), .A2(n10627), .ZN(n10766) );
  OR2_X1 U8999 ( .A1(n10350), .A2(n11091), .ZN(n13595) );
  NOR2_X1 U9000 ( .A1(n10347), .A2(n10462), .ZN(n13602) );
  INV_X1 U9001 ( .A(n13033), .ZN(n8210) );
  INV_X1 U9002 ( .A(n13847), .ZN(n13874) );
  INV_X1 U9003 ( .A(n13900), .ZN(n13873) );
  INV_X1 U9004 ( .A(n12807), .ZN(n13913) );
  INV_X1 U9005 ( .A(n13899), .ZN(n13928) );
  OR2_X1 U9006 ( .A1(n10322), .A2(n8814), .ZN(n10324) );
  INV_X1 U9007 ( .A(n8440), .ZN(n10572) );
  INV_X1 U9008 ( .A(n8442), .ZN(n10957) );
  INV_X1 U9009 ( .A(n8282), .ZN(n10945) );
  AND2_X1 U9010 ( .A1(n8285), .A2(n8284), .ZN(n15925) );
  AND2_X1 U9011 ( .A1(n7446), .A2(n7827), .ZN(n15923) );
  INV_X1 U9012 ( .A(n13631), .ZN(n8435) );
  OAI21_X1 U9013 ( .B1(n15979), .B2(n8434), .A(n8433), .ZN(n13675) );
  NAND2_X1 U9014 ( .A1(n8437), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8434) );
  INV_X1 U9015 ( .A(n13633), .ZN(n8437) );
  AND2_X1 U9016 ( .A1(n12986), .A2(n12985), .ZN(n13739) );
  INV_X1 U9017 ( .A(n8036), .ZN(n13748) );
  OR2_X1 U9018 ( .A1(n13744), .A2(n9196), .ZN(n13761) );
  NAND2_X1 U9019 ( .A1(n13892), .A2(n12942), .ZN(n13877) );
  NAND2_X1 U9020 ( .A1(n9070), .A2(n9069), .ZN(n14005) );
  OR2_X1 U9021 ( .A1(n11991), .A2(n8385), .ZN(n8381) );
  AND3_X1 U9022 ( .A1(n8988), .A2(n8987), .A3(n8986), .ZN(n12156) );
  OAI21_X1 U9023 ( .B1(n9236), .B2(n8397), .A(n8395), .ZN(n12030) );
  NAND2_X1 U9024 ( .A1(n11673), .A2(n9237), .ZN(n11804) );
  NAND2_X1 U9025 ( .A1(n8877), .A2(n12886), .ZN(n11533) );
  OR2_X1 U9026 ( .A1(n11094), .A2(n16115), .ZN(n13963) );
  AND2_X1 U9027 ( .A1(n16121), .A2(n11214), .ZN(n13967) );
  OR2_X1 U9028 ( .A1(n11091), .A2(n11093), .ZN(n16113) );
  INV_X1 U9029 ( .A(n16113), .ZN(n13868) );
  NAND2_X1 U9030 ( .A1(n8203), .A2(n8204), .ZN(n13766) );
  INV_X1 U9031 ( .A(n13739), .ZN(n16416) );
  OAI21_X1 U9032 ( .B1(n13464), .B2(n8873), .A(n12978), .ZN(n16409) );
  NAND2_X1 U9033 ( .A1(n16415), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n7741) );
  NAND2_X1 U9034 ( .A1(n8260), .A2(n9165), .ZN(n14048) );
  NAND2_X1 U9035 ( .A1(n8370), .A2(n8374), .ZN(n13786) );
  NAND2_X1 U9036 ( .A1(n8375), .A2(n8377), .ZN(n13800) );
  NAND2_X1 U9037 ( .A1(n9119), .A2(n9118), .ZN(n14068) );
  AND2_X1 U9038 ( .A1(n13841), .A2(n13840), .ZN(n14066) );
  NAND2_X1 U9039 ( .A1(n7627), .A2(n8191), .ZN(n13859) );
  OR2_X1 U9040 ( .A1(n14016), .A2(n14015), .ZN(n14090) );
  NAND2_X1 U9041 ( .A1(n8995), .A2(n8994), .ZN(n14097) );
  INV_X1 U9042 ( .A(n9242), .ZN(n14101) );
  NAND2_X1 U9043 ( .A1(n7637), .A2(n12875), .ZN(n11297) );
  AND2_X1 U9044 ( .A1(n9287), .A2(n9286), .ZN(n14108) );
  OR2_X1 U9045 ( .A1(n9500), .A2(P3_D_REG_1__SCAN_IN), .ZN(n9287) );
  INV_X1 U9046 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n8799) );
  XNOR2_X1 U9047 ( .A(n9175), .B(n9174), .ZN(n11869) );
  OR2_X1 U9048 ( .A1(n9148), .A2(n9147), .ZN(n9149) );
  NAND2_X1 U9049 ( .A1(n9277), .A2(n9278), .ZN(n11294) );
  NAND2_X1 U9050 ( .A1(n8227), .A2(n8758), .ZN(n9103) );
  MUX2_X1 U9051 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9212), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n9214) );
  OAI211_X1 U9052 ( .C1(n8756), .C2(n13096), .A(n8225), .B(n8221), .ZN(n9091)
         );
  NAND2_X1 U9053 ( .A1(n8756), .A2(n7603), .ZN(n8221) );
  INV_X1 U9054 ( .A(SI_19_), .ZN(n15473) );
  INV_X1 U9055 ( .A(SI_18_), .ZN(n11001) );
  NAND2_X1 U9056 ( .A1(n7701), .A2(n8749), .ZN(n9050) );
  NAND2_X1 U9057 ( .A1(n9033), .A2(n9032), .ZN(n7701) );
  NAND2_X1 U9058 ( .A1(n8781), .A2(n8935), .ZN(n9034) );
  NAND2_X1 U9059 ( .A1(n7707), .A2(n8746), .ZN(n9018) );
  NAND2_X1 U9060 ( .A1(n8990), .A2(n8989), .ZN(n7707) );
  INV_X1 U9061 ( .A(SI_15_), .ZN(n10244) );
  INV_X1 U9062 ( .A(SI_14_), .ZN(n9871) );
  OAI211_X1 U9063 ( .C1(n8978), .C2(n8243), .A(n8235), .B(n8238), .ZN(n9001)
         );
  NAND2_X1 U9064 ( .A1(n8978), .A2(n8241), .ZN(n8235) );
  INV_X1 U9065 ( .A(SI_12_), .ZN(n15485) );
  NAND2_X1 U9066 ( .A1(n8924), .A2(n8933), .ZN(n10958) );
  NAND2_X1 U9067 ( .A1(n8230), .A2(n8734), .ZN(n8919) );
  NAND2_X1 U9068 ( .A1(n8902), .A2(n8901), .ZN(n8230) );
  NAND2_X1 U9069 ( .A1(n8731), .A2(n8730), .ZN(n8870) );
  NAND2_X1 U9070 ( .A1(n8855), .A2(n8854), .ZN(n8731) );
  XNOR2_X1 U9071 ( .A(n8872), .B(P3_IR_REG_5__SCAN_IN), .ZN(n10497) );
  OAI21_X1 U9072 ( .B1(n8844), .B2(P3_IR_REG_3__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7835) );
  OAI211_X1 U9073 ( .C1(n8819), .C2(n7689), .A(n8726), .B(n7690), .ZN(n8843)
         );
  NAND2_X1 U9074 ( .A1(n7693), .A2(n8832), .ZN(n7690) );
  INV_X1 U9075 ( .A(n8725), .ZN(n7693) );
  NAND2_X1 U9076 ( .A1(n8819), .A2(n8725), .ZN(n8833) );
  CLKBUF_X1 U9077 ( .A(n10327), .Z(n8065) );
  AND2_X1 U9078 ( .A1(n8480), .A2(n8478), .ZN(n11958) );
  NAND2_X1 U9079 ( .A1(n8480), .A2(n11814), .ZN(n11817) );
  NAND2_X1 U9080 ( .A1(n13278), .A2(n9720), .ZN(n8162) );
  INV_X1 U9081 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n11151) );
  INV_X1 U9082 ( .A(n8500), .ZN(n9783) );
  NAND2_X1 U9083 ( .A1(n8466), .A2(n8469), .ZN(n14166) );
  OR2_X1 U9084 ( .A1(n14125), .A2(n14124), .ZN(n8466) );
  XNOR2_X1 U9085 ( .A(n9724), .B(n9725), .ZN(n9664) );
  NAND2_X1 U9086 ( .A1(n8452), .A2(n8457), .ZN(n14187) );
  OR2_X1 U9087 ( .A1(n14125), .A2(n8458), .ZN(n8452) );
  AND2_X1 U9088 ( .A1(n8512), .A2(n11514), .ZN(n11518) );
  INV_X1 U9089 ( .A(n7618), .ZN(n7617) );
  OAI21_X1 U9090 ( .B1(n8449), .B2(n7619), .A(n14141), .ZN(n7618) );
  NAND2_X1 U9091 ( .A1(n8451), .A2(n8449), .ZN(n14201) );
  NAND2_X1 U9092 ( .A1(n8461), .A2(n8464), .ZN(n14207) );
  NAND2_X1 U9093 ( .A1(n14125), .A2(n8462), .ZN(n8461) );
  INV_X1 U9094 ( .A(n8512), .ZN(n11515) );
  NAND2_X1 U9095 ( .A1(n11816), .A2(n8478), .ZN(n8471) );
  AND2_X1 U9096 ( .A1(n13417), .A2(n13455), .ZN(n8687) );
  NAND4_X1 U9097 ( .A1(n9748), .A2(n9747), .A3(n9746), .A4(n9745), .ZN(n14263)
         );
  AOI21_X1 U9098 ( .B1(n9562), .B2(P2_REG2_REG_1__SCAN_IN), .A(n15793), .ZN(
        n15806) );
  AOI21_X1 U9099 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n15809), .A(n15801), .ZN(
        n9684) );
  AOI21_X1 U9100 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n9729), .A(n9682), .ZN(
        n9580) );
  AOI21_X1 U9101 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n9729), .A(n9685), .ZN(
        n9577) );
  INV_X1 U9102 ( .A(n7734), .ZN(n9568) );
  NOR2_X1 U9103 ( .A1(n9590), .A2(n7578), .ZN(n9593) );
  AOI21_X1 U9104 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n9817), .A(n9587), .ZN(
        n9589) );
  AOI21_X1 U9105 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n10022), .A(n9761), .ZN(
        n9764) );
  INV_X1 U9106 ( .A(n7736), .ZN(n15815) );
  NOR2_X1 U9107 ( .A1(n15812), .A2(n8009), .ZN(n10196) );
  AND2_X1 U9108 ( .A1(n15822), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8009) );
  NAND2_X1 U9109 ( .A1(n10196), .A2(n10195), .ZN(n10647) );
  AOI21_X1 U9110 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n11134), .A(n10834), .ZN(
        n10838) );
  NAND2_X1 U9111 ( .A1(n11425), .A2(n7747), .ZN(n11426) );
  OR2_X1 U9112 ( .A1(n11431), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7747) );
  NOR2_X1 U9113 ( .A1(n11640), .A2(n8007), .ZN(n11643) );
  AND2_X1 U9114 ( .A1(n11691), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8007) );
  NOR2_X1 U9115 ( .A1(n12223), .A2(n15826), .ZN(n12226) );
  NOR2_X1 U9116 ( .A1(n15831), .A2(n12217), .ZN(n12219) );
  NOR2_X1 U9117 ( .A1(n14298), .A2(n7730), .ZN(n14289) );
  NOR2_X1 U9118 ( .A1(n7731), .A2(n14286), .ZN(n7730) );
  NAND2_X1 U9119 ( .A1(n14289), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n14300) );
  OR2_X1 U9120 ( .A1(n9566), .A2(n14314), .ZN(n15817) );
  AOI21_X1 U9121 ( .B1(n14296), .B2(n11940), .A(n8044), .ZN(n8043) );
  INV_X1 U9122 ( .A(n14297), .ZN(n8042) );
  AND2_X1 U9123 ( .A1(n13385), .A2(n13384), .ZN(n14371) );
  NAND2_X1 U9124 ( .A1(n14365), .A2(n8153), .ZN(n14567) );
  AOI21_X1 U9125 ( .B1(n7803), .B2(n7802), .A(n7801), .ZN(n8067) );
  NOR2_X1 U9126 ( .A1(n8153), .A2(n12045), .ZN(n7801) );
  NAND2_X1 U9127 ( .A1(n8588), .A2(n8589), .ZN(n14385) );
  NAND2_X1 U9128 ( .A1(n8302), .A2(n8305), .ZN(n14377) );
  NAND2_X1 U9129 ( .A1(n14404), .A2(n8306), .ZN(n8302) );
  OAI21_X1 U9130 ( .B1(n14406), .B2(n14407), .A(n7444), .ZN(n14392) );
  NAND2_X1 U9131 ( .A1(n14404), .A2(n8310), .ZN(n14391) );
  NAND2_X1 U9132 ( .A1(n8313), .A2(n8314), .ZN(n14434) );
  OR2_X1 U9133 ( .A1(n14478), .A2(n8316), .ZN(n8313) );
  NAND2_X1 U9134 ( .A1(n8317), .A2(n7439), .ZN(n14465) );
  NAND2_X1 U9135 ( .A1(n14478), .A2(n8322), .ZN(n8317) );
  NAND2_X1 U9136 ( .A1(n8600), .A2(n8601), .ZN(n14454) );
  NAND2_X1 U9137 ( .A1(n8606), .A2(n8603), .ZN(n14469) );
  INV_X1 U9138 ( .A(n8605), .ZN(n8603) );
  AND2_X1 U9139 ( .A1(n13098), .A2(n13097), .ZN(n14493) );
  NAND2_X1 U9140 ( .A1(n12043), .A2(n11948), .ZN(n14323) );
  NAND2_X1 U9141 ( .A1(n11947), .A2(n11946), .ZN(n12041) );
  INV_X1 U9142 ( .A(n14633), .ZN(n13227) );
  NAND2_X1 U9143 ( .A1(n7783), .A2(n11763), .ZN(n11908) );
  NAND2_X1 U9144 ( .A1(n16350), .A2(n11345), .ZN(n11772) );
  INV_X1 U9145 ( .A(n7800), .ZN(n16350) );
  NAND2_X1 U9146 ( .A1(n11277), .A2(n11250), .ZN(n11252) );
  NAND2_X1 U9147 ( .A1(n7790), .A2(n11248), .ZN(n11279) );
  NAND2_X1 U9148 ( .A1(n10809), .A2(n13433), .ZN(n11266) );
  NAND2_X1 U9149 ( .A1(n16269), .A2(n10808), .ZN(n10809) );
  NAND2_X1 U9150 ( .A1(n7809), .A2(n7810), .ZN(n10673) );
  OR2_X1 U9151 ( .A1(n10553), .A2(n13429), .ZN(n7809) );
  NAND2_X1 U9152 ( .A1(n8595), .A2(n10537), .ZN(n10587) );
  INV_X1 U9153 ( .A(n16169), .ZN(n10436) );
  NAND2_X1 U9154 ( .A1(n7776), .A2(n13423), .ZN(n10662) );
  INV_X1 U9155 ( .A(n14510), .ZN(n16394) );
  INV_X1 U9156 ( .A(n13216), .ZN(n13217) );
  NAND2_X2 U9157 ( .A1(n10024), .A2(n10023), .ZN(n16223) );
  INV_X1 U9158 ( .A(n14311), .ZN(n14641) );
  OAI211_X1 U9159 ( .C1(n16262), .C2(n14581), .A(n8002), .B(n8000), .ZN(n14649) );
  NOR2_X1 U9160 ( .A1(n14579), .A2(n8001), .ZN(n8000) );
  INV_X1 U9161 ( .A(n14578), .ZN(n8002) );
  AND2_X1 U9162 ( .A1(n14580), .A2(n16170), .ZN(n8001) );
  INV_X1 U9163 ( .A(n14336), .ZN(n14674) );
  INV_X1 U9164 ( .A(n14547), .ZN(n10283) );
  AND2_X1 U9165 ( .A1(n9645), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15784) );
  OR2_X1 U9166 ( .A1(n9616), .A2(n9615), .ZN(n15783) );
  INV_X1 U9167 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n14676) );
  NAND2_X1 U9168 ( .A1(n9636), .A2(n7794), .ZN(n12848) );
  AOI21_X1 U9169 ( .B1(n7796), .B2(n7495), .A(n7795), .ZN(n7794) );
  NOR2_X1 U9170 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n7795) );
  XNOR2_X1 U9171 ( .A(n9337), .B(n9533), .ZN(n14688) );
  NAND2_X1 U9172 ( .A1(n9340), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9337) );
  NAND2_X1 U9173 ( .A1(n9340), .A2(n9339), .ZN(n14690) );
  OR2_X1 U9174 ( .A1(n9338), .A2(n9534), .ZN(n9339) );
  AOI21_X1 U9175 ( .B1(n9541), .B2(n7498), .A(n8495), .ZN(n8494) );
  NOR2_X1 U9176 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n8495) );
  INV_X1 U9177 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n13263) );
  INV_X1 U9178 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10830) );
  INV_X1 U9179 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10761) );
  NAND2_X1 U9180 ( .A1(n8056), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10608) );
  INV_X1 U9181 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9882) );
  INV_X1 U9182 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9780) );
  INV_X1 U9183 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9757) );
  INV_X1 U9184 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9678) );
  INV_X1 U9185 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9430) );
  INV_X1 U9186 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9418) );
  INV_X1 U9187 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9399) );
  NOR2_X1 U9188 ( .A1(n10095), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14685) );
  INV_X1 U9189 ( .A(n9403), .ZN(n7749) );
  OR2_X1 U9190 ( .A1(n10175), .A2(P1_U3086), .ZN(n9696) );
  NAND2_X1 U9191 ( .A1(n10733), .A2(n10732), .ZN(n10736) );
  NAND2_X1 U9192 ( .A1(n11488), .A2(n11487), .ZN(n11490) );
  INV_X1 U9193 ( .A(n8017), .ZN(n14729) );
  NAND2_X1 U9194 ( .A1(n14776), .A2(n8164), .ZN(n14730) );
  NAND2_X1 U9195 ( .A1(n11015), .A2(n11014), .ZN(n7640) );
  NAND2_X1 U9196 ( .A1(n14746), .A2(n12385), .ZN(n14757) );
  OR2_X1 U9197 ( .A1(n12440), .A2(n12439), .ZN(n7967) );
  NAND2_X1 U9198 ( .A1(n12442), .A2(n12441), .ZN(n15138) );
  NAND2_X1 U9199 ( .A1(n11362), .A2(n12491), .ZN(n8091) );
  AOI21_X1 U9200 ( .B1(n14721), .B2(n14722), .A(n7577), .ZN(n14778) );
  INV_X1 U9201 ( .A(n12208), .ZN(n7651) );
  INV_X1 U9202 ( .A(n12207), .ZN(n7652) );
  INV_X1 U9203 ( .A(n7647), .ZN(n14783) );
  INV_X1 U9204 ( .A(n7985), .ZN(n8051) );
  NAND2_X1 U9205 ( .A1(n11981), .A2(n11980), .ZN(n11984) );
  NAND2_X1 U9206 ( .A1(n7644), .A2(n10101), .ZN(n8524) );
  INV_X1 U9207 ( .A(n8523), .ZN(n8522) );
  AND2_X1 U9208 ( .A1(n10738), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14811) );
  NAND2_X1 U9209 ( .A1(n14794), .A2(n14795), .ZN(n14793) );
  NAND2_X1 U9210 ( .A1(n14756), .A2(n14760), .ZN(n14794) );
  NAND2_X1 U9211 ( .A1(n12078), .A2(n12077), .ZN(n14827) );
  NAND2_X1 U9212 ( .A1(n7903), .A2(n7904), .ZN(n12792) );
  NAND2_X1 U9213 ( .A1(n12684), .A2(n12683), .ZN(n7904) );
  OR2_X1 U9214 ( .A1(n12769), .A2(n12770), .ZN(n8022) );
  INV_X1 U9215 ( .A(n12561), .ZN(n14858) );
  AND2_X1 U9216 ( .A1(n10100), .A2(n10098), .ZN(n7983) );
  AND3_X1 U9217 ( .A1(n10091), .A2(n10093), .A3(n10090), .ZN(n7986) );
  INV_X1 U9218 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n15694) );
  XNOR2_X1 U9219 ( .A(n9876), .B(P1_IR_REG_14__SCAN_IN), .ZN(n14901) );
  NAND2_X1 U9220 ( .A1(n7668), .A2(n16322), .ZN(n15102) );
  XNOR2_X1 U9221 ( .A(n14917), .B(n8182), .ZN(n7668) );
  INV_X1 U9222 ( .A(n14911), .ZN(n15105) );
  AND2_X1 U9223 ( .A1(n8351), .A2(n8356), .ZN(n14971) );
  AND2_X1 U9224 ( .A1(n8083), .A2(n7471), .ZN(n14968) );
  INV_X1 U9225 ( .A(n8351), .ZN(n14989) );
  NAND2_X1 U9226 ( .A1(n8325), .A2(n8327), .ZN(n15012) );
  NAND2_X1 U9227 ( .A1(n15040), .A2(n13066), .ZN(n15026) );
  NAND2_X1 U9228 ( .A1(n12338), .A2(n12337), .ZN(n15049) );
  NAND2_X1 U9229 ( .A1(n15071), .A2(n13046), .ZN(n15057) );
  NAND2_X1 U9230 ( .A1(n15073), .A2(n13062), .ZN(n15055) );
  NAND2_X1 U9231 ( .A1(n12178), .A2(n12177), .ZN(n14745) );
  NAND2_X1 U9232 ( .A1(n12080), .A2(n8669), .ZN(n12174) );
  NAND2_X1 U9233 ( .A1(n12007), .A2(n12006), .ZN(n12009) );
  NAND2_X1 U9234 ( .A1(n12001), .A2(n12000), .ZN(n12074) );
  INV_X1 U9235 ( .A(n15054), .ZN(n15058) );
  NAND2_X1 U9236 ( .A1(n11780), .A2(n12491), .ZN(n8005) );
  NAND2_X1 U9237 ( .A1(n11579), .A2(n11578), .ZN(n16326) );
  INV_X1 U9238 ( .A(n16324), .ZN(n16338) );
  NAND2_X1 U9239 ( .A1(n7677), .A2(n8656), .ZN(n11599) );
  NAND2_X1 U9240 ( .A1(n11394), .A2(n8654), .ZN(n7677) );
  NAND2_X1 U9241 ( .A1(n11375), .A2(n12733), .ZN(n11544) );
  NAND2_X1 U9242 ( .A1(n11396), .A2(n11374), .ZN(n11375) );
  INV_X1 U9243 ( .A(n16341), .ZN(n15051) );
  NAND2_X1 U9244 ( .A1(n8341), .A2(n11051), .ZN(n11355) );
  NAND2_X1 U9245 ( .A1(n7673), .A2(n14857), .ZN(n8088) );
  NAND2_X1 U9246 ( .A1(n10168), .A2(n10167), .ZN(n16161) );
  INV_X1 U9247 ( .A(n16163), .ZN(n16337) );
  NAND2_X1 U9248 ( .A1(n16086), .A2(n10936), .ZN(n16163) );
  AND2_X1 U9249 ( .A1(n16159), .A2(n12752), .ZN(n16341) );
  NAND2_X1 U9250 ( .A1(n15102), .A2(n7666), .ZN(n15218) );
  INV_X1 U9251 ( .A(n7667), .ZN(n7666) );
  OAI21_X1 U9252 ( .B1(n8182), .B2(n16378), .A(n15103), .ZN(n7667) );
  NOR2_X1 U9253 ( .A1(n15110), .A2(n15109), .ZN(n8033) );
  NAND2_X1 U9254 ( .A1(n15111), .A2(n16194), .ZN(n8034) );
  INV_X1 U9255 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n15237) );
  INV_X1 U9256 ( .A(n7686), .ZN(n15238) );
  XNOR2_X1 U9257 ( .A(n12712), .B(n12711), .ZN(n15236) );
  OAI21_X1 U9258 ( .B1(n12692), .B2(n8411), .A(n8408), .ZN(n12712) );
  XNOR2_X1 U9259 ( .A(n12312), .B(n12311), .ZN(n15249) );
  NAND2_X1 U9260 ( .A1(n12474), .A2(n12300), .ZN(n12312) );
  XNOR2_X1 U9261 ( .A(n9355), .B(P1_IR_REG_26__SCAN_IN), .ZN(n15253) );
  OAI21_X1 U9262 ( .B1(n9354), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9355) );
  NAND2_X1 U9263 ( .A1(n12297), .A2(n12296), .ZN(n12472) );
  INV_X1 U9264 ( .A(n12540), .ZN(n10944) );
  NAND2_X1 U9265 ( .A1(n8137), .A2(n8135), .ZN(n11321) );
  NAND2_X1 U9266 ( .A1(n8137), .A2(n8138), .ZN(n10915) );
  INV_X1 U9267 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n12336) );
  INV_X1 U9268 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10250) );
  INV_X1 U9269 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9877) );
  INV_X1 U9270 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9509) );
  INV_X1 U9271 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9449) );
  INV_X1 U9272 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9437) );
  NAND2_X1 U9273 ( .A1(n7441), .A2(n15919), .ZN(n15918) );
  INV_X1 U9274 ( .A(n7949), .ZN(n15865) );
  XNOR2_X1 U9275 ( .A(n15727), .B(n8572), .ZN(n15867) );
  INV_X1 U9276 ( .A(n15728), .ZN(n8572) );
  XNOR2_X1 U9277 ( .A(n15733), .B(n8571), .ZN(n15917) );
  INV_X1 U9278 ( .A(n15734), .ZN(n8571) );
  AND2_X1 U9279 ( .A1(n7960), .A2(n7460), .ZN(n15743) );
  AND2_X1 U9280 ( .A1(n7960), .A2(n7959), .ZN(n15871) );
  AND2_X1 U9281 ( .A1(n7460), .A2(n15742), .ZN(n7959) );
  INV_X1 U9282 ( .A(n7958), .ZN(n15878) );
  AOI21_X1 U9283 ( .B1(n15752), .B2(n15751), .A(n15880), .ZN(n15886) );
  NAND2_X1 U9284 ( .A1(n7962), .A2(n7961), .ZN(n15894) );
  NAND2_X1 U9285 ( .A1(n15889), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7961) );
  NAND2_X1 U9286 ( .A1(n15890), .A2(n7448), .ZN(n7962) );
  NOR2_X1 U9287 ( .A1(n15764), .A2(n15765), .ZN(n15896) );
  NAND2_X1 U9288 ( .A1(n15910), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n8582) );
  NAND2_X1 U9289 ( .A1(n7945), .A2(n8566), .ZN(n7943) );
  INV_X1 U9290 ( .A(n8567), .ZN(n7948) );
  INV_X1 U9291 ( .A(n15916), .ZN(n8580) );
  INV_X1 U9292 ( .A(n8063), .ZN(n8062) );
  NAND2_X1 U9293 ( .A1(n7900), .A2(n13587), .ZN(n7897) );
  NAND2_X1 U9294 ( .A1(n13584), .A2(n7896), .ZN(n7895) );
  AND2_X1 U9295 ( .A1(n11303), .A2(n11302), .ZN(n11305) );
  NOR2_X1 U9296 ( .A1(n8250), .A2(n9947), .ZN(n8247) );
  INV_X1 U9297 ( .A(n7702), .ZN(n8248) );
  INV_X1 U9298 ( .A(n8436), .ZN(n15978) );
  OAI21_X1 U9299 ( .B1(n13714), .B2(n15999), .A(n7523), .ZN(P3_U3200) );
  AOI21_X1 U9300 ( .B1(n13731), .B2(n15966), .A(n8049), .ZN(n8048) );
  NAND2_X1 U9301 ( .A1(n9309), .A2(n8054), .ZN(n8053) );
  INV_X1 U9302 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n8054) );
  NOR2_X1 U9303 ( .A1(n7583), .A2(n8029), .ZN(n8028) );
  NOR2_X1 U9304 ( .A1(n16410), .A2(n9324), .ZN(n8029) );
  NAND2_X1 U9305 ( .A1(n7742), .A2(n7739), .ZN(P3_U3455) );
  INV_X1 U9306 ( .A(n7740), .ZN(n7739) );
  NAND2_X1 U9307 ( .A1(n14038), .A2(n16410), .ZN(n7742) );
  OAI21_X1 U9308 ( .B1(n14039), .B2(n14102), .A(n7741), .ZN(n7740) );
  NAND2_X1 U9309 ( .A1(n9164), .A2(n9163), .ZN(n11595) );
  NAND2_X1 U9310 ( .A1(n10402), .A2(n10401), .ZN(n10403) );
  NAND2_X1 U9311 ( .A1(n8485), .A2(n8489), .ZN(n8484) );
  OAI21_X1 U9312 ( .B1(n9827), .B2(n7611), .A(n14232), .ZN(n9838) );
  INV_X1 U9313 ( .A(n8688), .ZN(n8684) );
  NAND2_X1 U9314 ( .A1(n13454), .A2(n8687), .ZN(n8685) );
  NAND2_X1 U9315 ( .A1(n8616), .A2(n8613), .ZN(P2_U3236) );
  INV_X1 U9316 ( .A(n8614), .ZN(n8613) );
  OAI21_X1 U9317 ( .B1(n14566), .B2(n14497), .A(n8615), .ZN(n8614) );
  NAND2_X1 U9318 ( .A1(n7772), .A2(n7770), .ZN(P2_U3528) );
  OR2_X1 U9319 ( .A1(n16358), .A2(n7771), .ZN(n7770) );
  NAND2_X1 U9320 ( .A1(n14646), .A2(n16358), .ZN(n7772) );
  INV_X1 U9321 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n7771) );
  NAND2_X1 U9322 ( .A1(n7769), .A2(n7767), .ZN(P2_U3496) );
  INV_X1 U9323 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n7768) );
  XNOR2_X1 U9324 ( .A(n7966), .B(n12523), .ZN(n12536) );
  OAI21_X1 U9325 ( .B1(n8052), .B2(n14829), .A(n7592), .ZN(P1_U3240) );
  XNOR2_X1 U9326 ( .A(n14805), .B(n7574), .ZN(n8052) );
  OR2_X1 U9327 ( .A1(n16391), .A2(n8364), .ZN(n8363) );
  INV_X1 U9328 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n8364) );
  INV_X1 U9329 ( .A(n7950), .ZN(n15859) );
  INV_X1 U9330 ( .A(n8575), .ZN(n15873) );
  NOR2_X1 U9331 ( .A1(n15890), .A2(n15889), .ZN(n15888) );
  NAND2_X1 U9332 ( .A1(n15773), .A2(n15774), .ZN(n8569) );
  AND2_X1 U9333 ( .A1(n7947), .A2(n7946), .ZN(n15907) );
  NAND2_X1 U9334 ( .A1(n15909), .A2(n15908), .ZN(n7946) );
  OAI211_X1 U9335 ( .C1(n15773), .C2(n8566), .A(n7942), .B(n7945), .ZN(n7947)
         );
  XNOR2_X1 U9336 ( .A(n8581), .B(n8578), .ZN(SUB_1596_U4) );
  XNOR2_X1 U9337 ( .A(n8580), .B(n8579), .ZN(n8578) );
  NAND2_X1 U9338 ( .A1(n7545), .A2(n8582), .ZN(n8581) );
  XNOR2_X1 U9339 ( .A(n15911), .B(n8402), .ZN(n8579) );
  NAND2_X1 U9340 ( .A1(n8038), .A2(n8037), .ZN(n9258) );
  INV_X2 U9341 ( .A(n12543), .ZN(n12551) );
  AND2_X1 U9342 ( .A1(n14129), .A2(n14130), .ZN(n7435) );
  OR2_X1 U9343 ( .A1(n12045), .A2(n7805), .ZN(n7436) );
  AND2_X1 U9344 ( .A1(n12661), .A2(n8528), .ZN(n7437) );
  AND2_X1 U9345 ( .A1(n12637), .A2(n12639), .ZN(n7438) );
  OR2_X1 U9346 ( .A1(n14476), .A2(n14487), .ZN(n7439) );
  INV_X1 U9347 ( .A(n7431), .ZN(n14147) );
  XNOR2_X1 U9348 ( .A(n16365), .B(n14849), .ZN(n12736) );
  AND2_X1 U9349 ( .A1(n12455), .A2(n12454), .ZN(n7440) );
  INV_X1 U9350 ( .A(n13613), .ZN(n8384) );
  INV_X1 U9351 ( .A(n12728), .ZN(n8337) );
  AND2_X1 U9352 ( .A1(n7950), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n7441) );
  NAND2_X1 U9353 ( .A1(n14998), .A2(n8081), .ZN(n8083) );
  INV_X2 U9354 ( .A(n13360), .ZN(n13341) );
  INV_X1 U9355 ( .A(n16240), .ZN(n8342) );
  AND2_X1 U9356 ( .A1(n8314), .A2(n8312), .ZN(n7442) );
  AND2_X1 U9357 ( .A1(n13296), .A2(n13295), .ZN(n14657) );
  AND2_X1 U9358 ( .A1(n7810), .A2(n10672), .ZN(n7443) );
  AOI21_X1 U9359 ( .B1(n13808), .B2(n9201), .A(n9159), .ZN(n13543) );
  INV_X1 U9360 ( .A(n13543), .ZN(n8037) );
  OR2_X1 U9361 ( .A1(n14653), .A2(n14354), .ZN(n7444) );
  INV_X1 U9362 ( .A(n8649), .ZN(n8648) );
  AND2_X1 U9363 ( .A1(n8650), .A2(n12798), .ZN(n8649) );
  INV_X1 U9364 ( .A(n14476), .ZN(n14603) );
  AND2_X1 U9365 ( .A1(n13251), .A2(n13250), .ZN(n14476) );
  AND2_X1 U9366 ( .A1(n7647), .A2(n7596), .ZN(n7445) );
  OR2_X1 U9367 ( .A1(n13655), .A2(n7560), .ZN(n7446) );
  INV_X1 U9368 ( .A(n13421), .ZN(n10793) );
  INV_X1 U9369 ( .A(n10859), .ZN(n15095) );
  INV_X1 U9370 ( .A(n14667), .ZN(n14505) );
  AND2_X1 U9371 ( .A1(n13111), .A2(n13110), .ZN(n14667) );
  AND3_X1 U9372 ( .A1(n13771), .A2(n12854), .A3(n8257), .ZN(n7447) );
  OR2_X1 U9373 ( .A1(n15889), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7448) );
  AND2_X1 U9374 ( .A1(n13277), .A2(n13276), .ZN(n7449) );
  XNOR2_X1 U9375 ( .A(n7819), .B(n7818), .ZN(n13677) );
  INV_X1 U9376 ( .A(n13677), .ZN(n8016) );
  AND4_X1 U9377 ( .A1(n13018), .A2(n7579), .A3(n13017), .A4(n13027), .ZN(n7450) );
  NAND2_X1 U9378 ( .A1(n9146), .A2(n9145), .ZN(n13610) );
  INV_X1 U9379 ( .A(n13610), .ZN(n8379) );
  AND2_X1 U9380 ( .A1(n8218), .A2(n7501), .ZN(n7451) );
  INV_X1 U9381 ( .A(n14812), .ZN(n15126) );
  NAND2_X1 U9382 ( .A1(n12476), .A2(n12475), .ZN(n14812) );
  AND2_X1 U9383 ( .A1(n13335), .A2(n13334), .ZN(n14383) );
  INV_X1 U9384 ( .A(n14383), .ZN(n14574) );
  AND2_X1 U9385 ( .A1(n7659), .A2(n7658), .ZN(n7452) );
  AND2_X1 U9386 ( .A1(n8675), .A2(n7675), .ZN(n7453) );
  AND2_X1 U9387 ( .A1(n14048), .A2(n13775), .ZN(n12851) );
  INV_X1 U9388 ( .A(n12851), .ZN(n8258) );
  INV_X1 U9389 ( .A(n8294), .ZN(n8293) );
  OAI21_X1 U9390 ( .B1(n7457), .B2(n11345), .A(n11773), .ZN(n8294) );
  NAND2_X1 U9391 ( .A1(n12493), .A2(n12492), .ZN(n15119) );
  OAI22_X1 U9392 ( .A1(n14657), .A2(n13341), .B1(n14353), .B2(n13411), .ZN(
        n13304) );
  NAND2_X1 U9393 ( .A1(n12459), .A2(n12458), .ZN(n14972) );
  INV_X1 U9394 ( .A(n14972), .ZN(n15132) );
  INV_X1 U9395 ( .A(n12662), .ZN(n8528) );
  INV_X1 U9396 ( .A(n13259), .ZN(n7859) );
  NOR2_X1 U9397 ( .A1(n14089), .A2(n12807), .ZN(n7454) );
  AND2_X1 U9398 ( .A1(n7965), .A2(n8164), .ZN(n7455) );
  AND2_X1 U9399 ( .A1(n7833), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7456) );
  NOR2_X1 U9400 ( .A1(n13202), .A2(n14255), .ZN(n7457) );
  INV_X1 U9401 ( .A(n13910), .ZN(n7729) );
  INV_X1 U9402 ( .A(n13011), .ZN(n8394) );
  INV_X1 U9403 ( .A(n13437), .ZN(n7782) );
  AND2_X1 U9404 ( .A1(n14396), .A2(n8274), .ZN(n7458) );
  AND2_X1 U9405 ( .A1(n12161), .A2(n7889), .ZN(n7459) );
  AND2_X1 U9406 ( .A1(n8871), .A2(n8777), .ZN(n8935) );
  INV_X1 U9407 ( .A(n8658), .ZN(n12733) );
  XNOR2_X1 U9408 ( .A(n12592), .B(n14852), .ZN(n8658) );
  NAND2_X1 U9409 ( .A1(n12871), .A2(n12875), .ZN(n16099) );
  OR2_X1 U9410 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n15736), .ZN(n7460) );
  AND2_X1 U9411 ( .A1(n15000), .A2(n8185), .ZN(n7461) );
  INV_X1 U9412 ( .A(n10114), .ZN(n12016) );
  AND2_X1 U9413 ( .A1(n15243), .A2(n12308), .ZN(n10114) );
  AND4_X1 U9414 ( .A1(n7630), .A2(n7870), .A3(n8781), .A4(n8871), .ZN(n7462)
         );
  AOI22_X1 U9415 ( .A1(n8703), .A2(n8706), .B1(n8707), .B2(n8711), .ZN(n8702)
         );
  NAND2_X1 U9416 ( .A1(n7913), .A2(n9517), .ZN(n7912) );
  INV_X1 U9417 ( .A(n8670), .ZN(n8669) );
  NAND2_X1 U9418 ( .A1(n8673), .A2(n12079), .ZN(n8670) );
  NOR2_X1 U9419 ( .A1(n14042), .A2(n13787), .ZN(n7463) );
  AND2_X1 U9420 ( .A1(n13196), .A2(n13195), .ZN(n7464) );
  NAND2_X1 U9421 ( .A1(n14923), .A2(n8664), .ZN(n7465) );
  AND2_X1 U9422 ( .A1(n8103), .A2(n8106), .ZN(n7466) );
  OAI21_X1 U9423 ( .B1(n10457), .B2(n13034), .A(n10456), .ZN(n10763) );
  XNOR2_X1 U9424 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8832) );
  INV_X1 U9425 ( .A(n8832), .ZN(n7689) );
  AND2_X1 U9426 ( .A1(n8115), .A2(n8114), .ZN(n7467) );
  OR2_X1 U9427 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n15871), .ZN(n7468) );
  OAI21_X1 U9428 ( .B1(n14125), .B2(n8456), .A(n8453), .ZN(n8061) );
  NAND3_X1 U9429 ( .A1(n9051), .A2(n8652), .A3(n8651), .ZN(n7469) );
  AND2_X1 U9430 ( .A1(n7793), .A2(n7792), .ZN(n7470) );
  NAND2_X1 U9431 ( .A1(n14992), .A2(n14714), .ZN(n7471) );
  AND2_X1 U9432 ( .A1(n9537), .A2(n9536), .ZN(n7472) );
  AND2_X1 U9433 ( .A1(n8491), .A2(n8490), .ZN(n7473) );
  AND2_X1 U9434 ( .A1(n10573), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7474) );
  INV_X1 U9435 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9852) );
  AND2_X1 U9436 ( .A1(n14427), .A2(n14353), .ZN(n7475) );
  NAND2_X1 U9437 ( .A1(n14580), .A2(n14355), .ZN(n7476) );
  INV_X1 U9438 ( .A(n14264), .ZN(n8013) );
  INV_X1 U9439 ( .A(n14446), .ZN(n8265) );
  NAND2_X1 U9440 ( .A1(n8162), .A2(n13280), .ZN(n14446) );
  NAND2_X1 U9441 ( .A1(n7880), .A2(n7881), .ZN(n13541) );
  INV_X1 U9442 ( .A(n13441), .ZN(n7816) );
  XOR2_X1 U9443 ( .A(n15704), .B(n15902), .Z(n7477) );
  AND2_X1 U9444 ( .A1(n13612), .A2(n12156), .ZN(n7478) );
  INV_X1 U9445 ( .A(n13771), .ZN(n13765) );
  XNOR2_X1 U9446 ( .A(n14042), .B(n13787), .ZN(n13771) );
  OR2_X1 U9447 ( .A1(n13615), .A2(n11863), .ZN(n7479) );
  INV_X4 U9448 ( .A(n8873), .ZN(n8822) );
  AND3_X1 U9449 ( .A1(n15627), .A2(n8668), .A3(n15622), .ZN(n7480) );
  NAND4_X1 U9450 ( .A1(n10744), .A2(n10743), .A3(n10742), .A4(n10741), .ZN(
        n14857) );
  AND2_X1 U9451 ( .A1(n15174), .A2(n13063), .ZN(n7481) );
  AND2_X1 U9452 ( .A1(n16392), .A2(n11764), .ZN(n7482) );
  OR2_X1 U9453 ( .A1(n12639), .A2(n12637), .ZN(n7483) );
  OR2_X1 U9454 ( .A1(n11121), .A2(n11120), .ZN(n7484) );
  OR2_X1 U9455 ( .A1(n8265), .A2(n14352), .ZN(n7485) );
  AND3_X1 U9456 ( .A1(n9652), .A2(n9653), .A3(n9651), .ZN(n7486) );
  NOR2_X1 U9457 ( .A1(n11510), .A2(n8513), .ZN(n7487) );
  INV_X1 U9458 ( .A(n13179), .ZN(n8102) );
  AND2_X1 U9459 ( .A1(n13026), .A2(n13028), .ZN(n7488) );
  AND3_X1 U9460 ( .A1(n7480), .A2(n7664), .A3(n8540), .ZN(n7489) );
  NOR2_X1 U9461 ( .A1(n12905), .A2(n7631), .ZN(n7490) );
  AND2_X1 U9462 ( .A1(n13047), .A2(n15042), .ZN(n7491) );
  AND2_X1 U9463 ( .A1(n13183), .A2(n14258), .ZN(n7492) );
  AND2_X1 U9464 ( .A1(n7874), .A2(n13507), .ZN(n7493) );
  NAND2_X1 U9465 ( .A1(n13366), .A2(n13365), .ZN(n14563) );
  INV_X1 U9466 ( .A(n7911), .ZN(n7910) );
  OAI21_X1 U9467 ( .B1(n7912), .B2(n9514), .A(n9713), .ZN(n7911) );
  INV_X1 U9468 ( .A(n8179), .ZN(n8178) );
  OAI21_X1 U9469 ( .B1(n14769), .B2(n7440), .A(n8180), .ZN(n8179) );
  INV_X1 U9470 ( .A(n8267), .ZN(n14444) );
  NAND2_X1 U9471 ( .A1(n8268), .A2(n8265), .ZN(n8267) );
  INV_X1 U9472 ( .A(n8266), .ZN(n14426) );
  NAND2_X1 U9473 ( .A1(n8264), .A2(n8268), .ZN(n8266) );
  AND2_X1 U9474 ( .A1(n12629), .A2(n12628), .ZN(n7494) );
  INV_X1 U9475 ( .A(n12888), .ZN(n13006) );
  XNOR2_X1 U9476 ( .A(n13618), .B(n16215), .ZN(n12888) );
  AND2_X1 U9477 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n7495) );
  NOR2_X1 U9478 ( .A1(n12851), .A2(n8206), .ZN(n8205) );
  AND2_X1 U9479 ( .A1(n8502), .A2(n9824), .ZN(n7496) );
  AND2_X1 U9480 ( .A1(n8503), .A2(n7496), .ZN(n7497) );
  INV_X1 U9481 ( .A(n8568), .ZN(n8566) );
  NAND2_X1 U9482 ( .A1(n15901), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n8568) );
  AND2_X1 U9483 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n7498) );
  AND2_X1 U9484 ( .A1(n7459), .A2(n7887), .ZN(n7499) );
  AND2_X1 U9485 ( .A1(n7542), .A2(n13187), .ZN(n7500) );
  NAND2_X1 U9486 ( .A1(n9430), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7501) );
  INV_X1 U9487 ( .A(n8463), .ZN(n8462) );
  NAND2_X1 U9488 ( .A1(n8468), .A2(n8469), .ZN(n8463) );
  OR2_X1 U9489 ( .A1(n13019), .A2(n13752), .ZN(n7502) );
  AND2_X1 U9490 ( .A1(n13027), .A2(n7488), .ZN(n7503) );
  AND2_X1 U9491 ( .A1(n8436), .A2(n8435), .ZN(n7504) );
  INV_X1 U9492 ( .A(n15076), .ZN(n8361) );
  OR2_X1 U9493 ( .A1(n13442), .A2(n8296), .ZN(n7505) );
  AND2_X1 U9494 ( .A1(n8790), .A2(n8802), .ZN(n7506) );
  INV_X1 U9495 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7976) );
  INV_X1 U9496 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8169) );
  INV_X1 U9497 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8793) );
  INV_X1 U9498 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8802) );
  INV_X1 U9499 ( .A(n12581), .ZN(n8535) );
  INV_X1 U9500 ( .A(n14368), .ZN(n8298) );
  INV_X1 U9501 ( .A(n12146), .ZN(n8482) );
  NAND2_X1 U9502 ( .A1(n9349), .A2(n8542), .ZN(n7507) );
  INV_X1 U9503 ( .A(n14310), .ZN(n14645) );
  NAND2_X1 U9504 ( .A1(n13348), .A2(n13347), .ZN(n14310) );
  NOR2_X1 U9505 ( .A1(n16223), .A2(n14261), .ZN(n7508) );
  NOR2_X1 U9506 ( .A1(n8528), .A2(n12661), .ZN(n7509) );
  AND2_X1 U9507 ( .A1(n7476), .A2(n7444), .ZN(n7510) );
  NOR2_X1 U9508 ( .A1(n12592), .A2(n14852), .ZN(n7511) );
  NOR2_X1 U9509 ( .A1(n12655), .A2(n12657), .ZN(n7512) );
  AND2_X1 U9510 ( .A1(n13809), .A2(n8037), .ZN(n7513) );
  NOR2_X1 U9511 ( .A1(n15159), .A2(n14786), .ZN(n7514) );
  NOR2_X1 U9512 ( .A1(n14705), .A2(n12366), .ZN(n7515) );
  INV_X1 U9513 ( .A(n8698), .ZN(n8697) );
  NOR2_X1 U9514 ( .A1(n13207), .A2(n13206), .ZN(n8698) );
  NOR2_X1 U9515 ( .A1(n13918), .A2(n13928), .ZN(n7516) );
  NOR2_X1 U9516 ( .A1(n14048), .A2(n13801), .ZN(n7517) );
  INV_X1 U9517 ( .A(n8307), .ZN(n8306) );
  NAND2_X1 U9518 ( .A1(n8309), .A2(n8310), .ZN(n8307) );
  AND2_X1 U9519 ( .A1(n11600), .A2(n7678), .ZN(n7518) );
  AND2_X1 U9520 ( .A1(n10021), .A2(n10020), .ZN(n7519) );
  INV_X1 U9521 ( .A(n11204), .ZN(n8636) );
  NAND2_X1 U9522 ( .A1(n8492), .A2(n14179), .ZN(n7520) );
  AND2_X1 U9523 ( .A1(n16246), .A2(n13167), .ZN(n7521) );
  OR2_X1 U9524 ( .A1(n12620), .A2(n12619), .ZN(n7522) );
  AND2_X1 U9525 ( .A1(n8288), .A2(n8286), .ZN(n7523) );
  NOR2_X1 U9526 ( .A1(n14697), .A2(n8548), .ZN(n7524) );
  NAND2_X1 U9527 ( .A1(n12316), .A2(n9419), .ZN(n8724) );
  INV_X1 U9528 ( .A(n8724), .ZN(n7644) );
  AND2_X1 U9529 ( .A1(n10507), .A2(n10508), .ZN(n7525) );
  AND2_X1 U9530 ( .A1(n7782), .A2(n8292), .ZN(n7526) );
  XNOR2_X1 U9531 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8869) );
  AND2_X1 U9532 ( .A1(n16223), .A2(n10674), .ZN(n7527) );
  NAND2_X1 U9533 ( .A1(n14132), .A2(n14133), .ZN(n7528) );
  NAND2_X1 U9534 ( .A1(n13148), .A2(n13149), .ZN(n7529) );
  INV_X1 U9535 ( .A(n8186), .ZN(n8185) );
  NAND2_X1 U9536 ( .A1(n14992), .A2(n15132), .ZN(n8186) );
  AND2_X1 U9537 ( .A1(n9486), .A2(SI_8_), .ZN(n7530) );
  AND2_X1 U9538 ( .A1(n9447), .A2(SI_6_), .ZN(n7531) );
  AND2_X1 U9539 ( .A1(n9409), .A2(SI_4_), .ZN(n7532) );
  AND2_X1 U9540 ( .A1(n14580), .A2(n14330), .ZN(n7533) );
  INV_X1 U9541 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n9618) );
  INV_X1 U9542 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8782) );
  INV_X1 U9543 ( .A(n8643), .ZN(n8642) );
  NAND2_X1 U9544 ( .A1(n8644), .A2(n11856), .ZN(n8643) );
  NAND2_X1 U9545 ( .A1(n8184), .A2(n14947), .ZN(n7534) );
  OR2_X1 U9546 ( .A1(n12579), .A2(n12578), .ZN(n7535) );
  AND2_X1 U9547 ( .A1(n7645), .A2(n8163), .ZN(n7536) );
  AND2_X1 U9548 ( .A1(n8646), .A2(n7886), .ZN(n7537) );
  AND2_X1 U9549 ( .A1(n9418), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7538) );
  AND2_X1 U9550 ( .A1(n8735), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7539) );
  AND2_X1 U9551 ( .A1(n12973), .A2(n13023), .ZN(n7540) );
  INV_X1 U9552 ( .A(n7762), .ZN(n7761) );
  NAND2_X1 U9553 ( .A1(n7763), .A2(n8144), .ZN(n7762) );
  NAND2_X1 U9554 ( .A1(n9172), .A2(n9171), .ZN(n13801) );
  INV_X1 U9555 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8775) );
  NOR2_X1 U9556 ( .A1(n12813), .A2(n13887), .ZN(n7541) );
  AND2_X1 U9557 ( .A1(n8101), .A2(n8102), .ZN(n7542) );
  AND2_X1 U9558 ( .A1(n14854), .A2(n8342), .ZN(n7543) );
  NAND2_X1 U9559 ( .A1(n12561), .A2(n16143), .ZN(n7544) );
  AND2_X1 U9560 ( .A1(n7944), .A2(n7943), .ZN(n7545) );
  AND2_X1 U9561 ( .A1(n13306), .A2(n13305), .ZN(n14653) );
  INV_X1 U9562 ( .A(n14653), .ZN(n14412) );
  INV_X1 U9563 ( .A(n9222), .ZN(n14039) );
  NAND2_X1 U9564 ( .A1(n9193), .A2(n9192), .ZN(n9222) );
  NOR2_X1 U9565 ( .A1(n8265), .A2(n14456), .ZN(n7546) );
  INV_X1 U9566 ( .A(n13466), .ZN(n8626) );
  AOI21_X1 U9567 ( .B1(n12837), .B2(n13787), .A(n12838), .ZN(n13466) );
  OAI21_X1 U9568 ( .B1(n13407), .B2(n8419), .A(n8416), .ZN(n8415) );
  OR2_X1 U9569 ( .A1(n13728), .A2(n15991), .ZN(n7547) );
  AND2_X1 U9570 ( .A1(n8546), .A2(n8547), .ZN(n7548) );
  INV_X1 U9571 ( .A(n8118), .ZN(n8117) );
  NAND2_X1 U9572 ( .A1(n7464), .A2(n8120), .ZN(n8118) );
  NAND2_X1 U9573 ( .A1(n8260), .A2(n8259), .ZN(n12850) );
  NAND2_X1 U9574 ( .A1(n7533), .A2(n8309), .ZN(n8305) );
  NOR2_X1 U9575 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n7549) );
  INV_X1 U9576 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8540) );
  INV_X1 U9577 ( .A(n8459), .ZN(n8458) );
  AND2_X1 U9578 ( .A1(n8464), .A2(n8460), .ZN(n8459) );
  NAND2_X1 U9579 ( .A1(n7613), .A2(n7612), .ZN(n9635) );
  NAND2_X1 U9580 ( .A1(n9542), .A2(n8494), .ZN(n13093) );
  INV_X1 U9581 ( .A(n13093), .ZN(n13090) );
  OR2_X1 U9582 ( .A1(n13224), .A2(n13225), .ZN(n7550) );
  OR2_X1 U9583 ( .A1(n15126), .A2(n14835), .ZN(n7551) );
  OR2_X1 U9584 ( .A1(n13662), .A2(n13663), .ZN(n7552) );
  OR2_X1 U9585 ( .A1(n15725), .A2(n15724), .ZN(n7553) );
  AND2_X1 U9586 ( .A1(n11765), .A2(n11959), .ZN(n7554) );
  OR2_X1 U9587 ( .A1(n8703), .A2(n8707), .ZN(n7555) );
  AND2_X1 U9588 ( .A1(n12615), .A2(n12614), .ZN(n7556) );
  AND2_X1 U9589 ( .A1(n12932), .A2(n12933), .ZN(n13922) );
  AND2_X1 U9590 ( .A1(n12552), .A2(n12543), .ZN(n7557) );
  AND2_X1 U9591 ( .A1(n8299), .A2(n7804), .ZN(n7558) );
  AND2_X1 U9592 ( .A1(n10971), .A2(n10973), .ZN(n7559) );
  NOR2_X1 U9593 ( .A1(n15056), .A2(n8360), .ZN(n8359) );
  AND2_X1 U9594 ( .A1(n8432), .A2(n8431), .ZN(n7560) );
  AND2_X1 U9595 ( .A1(n14967), .A2(n7471), .ZN(n7561) );
  INV_X1 U9596 ( .A(n12385), .ZN(n8555) );
  NOR2_X1 U9597 ( .A1(n13290), .A2(n8109), .ZN(n7562) );
  AND2_X1 U9598 ( .A1(n12814), .A2(n13847), .ZN(n7563) );
  OR2_X1 U9599 ( .A1(n12684), .A2(n12683), .ZN(n7564) );
  OR2_X1 U9600 ( .A1(n13277), .A2(n13276), .ZN(n8110) );
  INV_X1 U9601 ( .A(n8110), .ZN(n8109) );
  AND2_X1 U9602 ( .A1(n13154), .A2(n13153), .ZN(n7565) );
  AND2_X1 U9603 ( .A1(n8485), .A2(n7520), .ZN(n7566) );
  AND2_X1 U9604 ( .A1(n8788), .A2(n8793), .ZN(n7567) );
  NAND2_X1 U9605 ( .A1(n8527), .A2(n12633), .ZN(n7568) );
  INV_X1 U9606 ( .A(n15028), .ZN(n15025) );
  AND2_X1 U9607 ( .A1(n8604), .A2(n8609), .ZN(n7569) );
  AND2_X1 U9608 ( .A1(n9852), .A2(n7976), .ZN(n7570) );
  INV_X1 U9609 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n15658) );
  NOR2_X1 U9610 ( .A1(n14338), .A2(n8295), .ZN(n7571) );
  INV_X1 U9611 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9631) );
  OR2_X1 U9612 ( .A1(n8626), .A2(n8624), .ZN(n7572) );
  AND2_X1 U9613 ( .A1(n8696), .A2(n13213), .ZN(n7573) );
  NAND2_X1 U9614 ( .A1(n9152), .A2(n9151), .ZN(n13809) );
  INV_X1 U9615 ( .A(n13809), .ZN(n8038) );
  INV_X1 U9616 ( .A(n13611), .ZN(n13848) );
  NAND2_X1 U9617 ( .A1(n11506), .A2(n7487), .ZN(n8512) );
  XNOR2_X1 U9618 ( .A(n12570), .B(n14856), .ZN(n12566) );
  INV_X1 U9619 ( .A(n12566), .ZN(n8675) );
  NAND2_X1 U9620 ( .A1(n7723), .A2(n9239), .ZN(n11991) );
  INV_X1 U9621 ( .A(n14369), .ZN(n7804) );
  INV_X1 U9622 ( .A(n14739), .ZN(n8180) );
  NAND2_X1 U9623 ( .A1(n8172), .A2(n12378), .ZN(n14819) );
  XNOR2_X1 U9624 ( .A(n12488), .B(n12487), .ZN(n7574) );
  INV_X1 U9625 ( .A(n9744), .ZN(n9829) );
  NOR2_X1 U9626 ( .A1(n16321), .A2(n16365), .ZN(n7672) );
  AND2_X1 U9627 ( .A1(n8742), .A2(n9775), .ZN(n7575) );
  AND2_X1 U9628 ( .A1(n16294), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7576) );
  AND2_X1 U9629 ( .A1(n12415), .A2(n12414), .ZN(n7577) );
  INV_X1 U9630 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n8387) );
  INV_X1 U9631 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n8388) );
  INV_X1 U9632 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n8047) );
  AND2_X1 U9633 ( .A1(n9817), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7578) );
  INV_X1 U9634 ( .A(n10959), .ZN(n11121) );
  NAND2_X1 U9635 ( .A1(n8381), .A2(n8383), .ZN(n12111) );
  OAI21_X1 U9636 ( .B1(n13925), .B2(n7729), .A(n7727), .ZN(n13897) );
  NOR4_X1 U9637 ( .A1(n13825), .A2(n13858), .A3(n13834), .A4(n13016), .ZN(
        n7579) );
  INV_X1 U9638 ( .A(n12942), .ZN(n8195) );
  AND2_X1 U9639 ( .A1(n8471), .A2(n8477), .ZN(n7580) );
  NAND2_X1 U9640 ( .A1(n12714), .A2(n12713), .ZN(n15101) );
  INV_X1 U9641 ( .A(n15101), .ZN(n8182) );
  AND2_X1 U9642 ( .A1(n15115), .A2(n16366), .ZN(n7581) );
  AND2_X1 U9643 ( .A1(n9784), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7582) );
  INV_X1 U9644 ( .A(n12636), .ZN(n7936) );
  AND2_X1 U9645 ( .A1(n9310), .A2(n9325), .ZN(n7583) );
  AND2_X1 U9646 ( .A1(n13048), .A2(n13047), .ZN(n7584) );
  AND2_X1 U9647 ( .A1(n15264), .A2(n12316), .ZN(n15155) );
  INV_X1 U9648 ( .A(n15155), .ZN(n15021) );
  INV_X1 U9649 ( .A(n14346), .ZN(n8607) );
  AND2_X1 U9650 ( .A1(n12287), .A2(n12286), .ZN(n14524) );
  AND2_X1 U9651 ( .A1(n13045), .A2(n13044), .ZN(n7585) );
  AND2_X1 U9652 ( .A1(n12920), .A2(n12921), .ZN(n13010) );
  INV_X1 U9653 ( .A(n13010), .ZN(n8200) );
  INV_X1 U9654 ( .A(n8140), .ZN(n8139) );
  NOR2_X1 U9655 ( .A1(n10911), .A2(n15280), .ZN(n8140) );
  AND2_X1 U9656 ( .A1(n12080), .A2(n12079), .ZN(n7586) );
  AND2_X1 U9657 ( .A1(n15039), .A2(n13049), .ZN(n7587) );
  AND2_X1 U9658 ( .A1(n12660), .A2(n7925), .ZN(n7588) );
  AND2_X1 U9659 ( .A1(n12247), .A2(n12246), .ZN(n7589) );
  INV_X1 U9660 ( .A(n13315), .ZN(n14354) );
  AND2_X1 U9661 ( .A1(n13314), .A2(n13313), .ZN(n13315) );
  AND2_X1 U9662 ( .A1(n13052), .A2(n13051), .ZN(n7590) );
  INV_X1 U9663 ( .A(n12673), .ZN(n8537) );
  INV_X1 U9664 ( .A(n8189), .ZN(n12257) );
  NOR2_X1 U9665 ( .A1(n12182), .A2(n14745), .ZN(n8189) );
  INV_X1 U9666 ( .A(n7826), .ZN(n7825) );
  NOR2_X1 U9667 ( .A1(n8431), .A2(n13655), .ZN(n7826) );
  AND2_X1 U9668 ( .A1(n8348), .A2(n11581), .ZN(n7591) );
  AND2_X1 U9669 ( .A1(n14813), .A2(n14814), .ZN(n7592) );
  NAND2_X1 U9670 ( .A1(n12418), .A2(n12419), .ZN(n7593) );
  AND2_X1 U9671 ( .A1(n14493), .A2(n14345), .ZN(n7594) );
  AND2_X1 U9672 ( .A1(n14074), .A2(n13862), .ZN(n7595) );
  NAND2_X1 U9673 ( .A1(n12422), .A2(n12423), .ZN(n7596) );
  INV_X1 U9674 ( .A(n12859), .ZN(n8257) );
  INV_X1 U9675 ( .A(n12654), .ZN(n7929) );
  NAND2_X1 U9676 ( .A1(n9016), .A2(n12925), .ZN(n7597) );
  INV_X1 U9677 ( .A(n14619), .ZN(n14536) );
  AND2_X1 U9678 ( .A1(n12276), .A2(n12275), .ZN(n14619) );
  AND2_X1 U9679 ( .A1(n12534), .A2(n12535), .ZN(n7598) );
  AND2_X1 U9680 ( .A1(n7882), .A2(n13838), .ZN(n7599) );
  INV_X1 U9681 ( .A(n8746), .ZN(n7710) );
  OR2_X1 U9682 ( .A1(n8537), .A2(n12672), .ZN(n7600) );
  AND2_X1 U9683 ( .A1(n12362), .A2(n12361), .ZN(n7601) );
  NAND2_X1 U9684 ( .A1(n9051), .A2(n8782), .ZN(n9066) );
  INV_X1 U9685 ( .A(n8242), .ZN(n8241) );
  NAND2_X1 U9686 ( .A1(n8977), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n8242) );
  NAND2_X1 U9687 ( .A1(n12811), .A2(n13873), .ZN(n8635) );
  NAND2_X1 U9688 ( .A1(n12654), .A2(n7930), .ZN(n7602) );
  INV_X1 U9689 ( .A(n12616), .ZN(n7671) );
  INV_X1 U9690 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n13096) );
  INV_X1 U9691 ( .A(n12740), .ZN(n8673) );
  AND2_X1 U9692 ( .A1(n9956), .A2(n8634), .ZN(n15931) );
  INV_X1 U9693 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8214) );
  INV_X1 U9694 ( .A(n9032), .ZN(n7697) );
  AND2_X1 U9695 ( .A1(n8755), .A2(n13096), .ZN(n7603) );
  NAND2_X1 U9696 ( .A1(n8386), .A2(n9227), .ZN(n11295) );
  NAND2_X1 U9697 ( .A1(n7790), .A2(n7788), .ZN(n11277) );
  NAND2_X1 U9698 ( .A1(n12251), .A2(n12250), .ZN(n15190) );
  INV_X1 U9699 ( .A(n15190), .ZN(n8188) );
  INV_X1 U9700 ( .A(n13608), .ZN(n13587) );
  NAND2_X1 U9701 ( .A1(n10344), .A2(n10349), .ZN(n13608) );
  NAND2_X1 U9702 ( .A1(n9138), .A2(n9137), .ZN(n14058) );
  AND2_X1 U9703 ( .A1(n10402), .A2(n8510), .ZN(n7604) );
  NOR2_X1 U9704 ( .A1(n9783), .A2(n9782), .ZN(n7605) );
  INV_X1 U9705 ( .A(n8271), .ZN(n10683) );
  AND2_X1 U9706 ( .A1(n13558), .A2(n8649), .ZN(n7606) );
  INV_X1 U9707 ( .A(n13178), .ZN(n8270) );
  INV_X1 U9708 ( .A(n14486), .ZN(n14529) );
  XNOR2_X1 U9709 ( .A(n9035), .B(n8214), .ZN(n13676) );
  AND2_X1 U9710 ( .A1(n12863), .A2(n13040), .ZN(n12974) );
  INV_X1 U9711 ( .A(n12974), .ZN(n12960) );
  NAND2_X1 U9712 ( .A1(n16178), .A2(n16274), .ZN(n16316) );
  INV_X2 U9713 ( .A(n16415), .ZN(n16410) );
  NAND2_X1 U9714 ( .A1(n16090), .A2(n16031), .ZN(n16077) );
  AND2_X1 U9715 ( .A1(n8632), .A2(n8629), .ZN(n7607) );
  INV_X1 U9716 ( .A(n16348), .ZN(n16262) );
  INV_X1 U9717 ( .A(n9885), .ZN(n13099) );
  OR2_X1 U9718 ( .A1(n7849), .A2(n13090), .ZN(n9885) );
  AND2_X1 U9719 ( .A1(n8762), .A2(n7719), .ZN(n7608) );
  AND2_X1 U9720 ( .A1(n10314), .A2(n13021), .ZN(n13036) );
  XNOR2_X1 U9721 ( .A(n9079), .B(n9202), .ZN(n13733) );
  INV_X1 U9722 ( .A(n13721), .ZN(n13719) );
  OR2_X1 U9723 ( .A1(n13421), .A2(n9660), .ZN(n7849) );
  AND2_X1 U9724 ( .A1(n13455), .A2(n13418), .ZN(n7609) );
  OR2_X1 U9725 ( .A1(n13721), .A2(n13890), .ZN(n7610) );
  INV_X1 U9726 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8795) );
  NAND2_X1 U9727 ( .A1(n9897), .A2(n15783), .ZN(n16359) );
  NAND2_X1 U9728 ( .A1(n14646), .A2(n14668), .ZN(n7769) );
  OR2_X1 U9729 ( .A1(n14668), .A2(n7768), .ZN(n7767) );
  INV_X2 U9730 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n8391) );
  NAND2_X1 U9731 ( .A1(n7615), .A2(n8690), .ZN(n9636) );
  NAND2_X1 U9732 ( .A1(n7614), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9545) );
  NAND2_X1 U9733 ( .A1(n7615), .A2(n8689), .ZN(n7796) );
  OAI21_X2 U9734 ( .B1(n8451), .B2(n7619), .A(n7617), .ZN(n14194) );
  NAND2_X1 U9735 ( .A1(n14194), .A2(n14193), .ZN(n14146) );
  NAND2_X2 U9736 ( .A1(n9547), .A2(n14314), .ZN(n11830) );
  XNOR2_X2 U9737 ( .A(n9540), .B(n9539), .ZN(n9547) );
  OAI21_X2 U9738 ( .B1(n8877), .B2(n12888), .A(n7620), .ZN(n11312) );
  OAI21_X2 U9739 ( .B1(n7627), .B2(n13858), .A(n7625), .ZN(n13846) );
  AND2_X2 U9740 ( .A1(n7629), .A2(n7630), .ZN(n9051) );
  INV_X1 U9741 ( .A(n12027), .ZN(n8956) );
  NAND2_X1 U9742 ( .A1(n7634), .A2(n12875), .ZN(n7636) );
  NAND3_X1 U9743 ( .A1(n8213), .A2(n12866), .A3(n12871), .ZN(n7634) );
  NAND2_X1 U9744 ( .A1(n7635), .A2(n12877), .ZN(n11215) );
  NAND4_X1 U9745 ( .A1(n8213), .A2(n12875), .A3(n12866), .A4(n12871), .ZN(
        n7637) );
  NAND2_X1 U9746 ( .A1(n7640), .A2(n11171), .ZN(n11175) );
  XNOR2_X1 U9747 ( .A(n7640), .B(n11018), .ZN(n11025) );
  INV_X2 U9748 ( .A(n16079), .ZN(n16090) );
  NAND2_X1 U9749 ( .A1(n7423), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7641) );
  NAND2_X1 U9750 ( .A1(n7644), .A2(n7643), .ZN(n7642) );
  NAND3_X1 U9751 ( .A1(n8166), .A2(n8170), .A3(n7656), .ZN(n7655) );
  NAND4_X1 U9752 ( .A1(n8168), .A2(n9346), .A3(n9410), .A4(
        P1_IR_REG_27__SCAN_IN), .ZN(n7656) );
  AND2_X2 U9753 ( .A1(n8187), .A2(n7657), .ZN(n16141) );
  AND3_X2 U9754 ( .A1(n10725), .A2(n10723), .A3(n10724), .ZN(n16162) );
  AND2_X2 U9755 ( .A1(n8522), .A2(n8524), .ZN(n10859) );
  INV_X1 U9756 ( .A(n9850), .ZN(n7661) );
  AND2_X2 U9757 ( .A1(n7480), .A2(n7664), .ZN(n9410) );
  AND2_X2 U9758 ( .A1(n7662), .A2(n7663), .ZN(n9346) );
  NAND4_X1 U9759 ( .A1(n9846), .A2(n9848), .A3(n9849), .A4(n9847), .ZN(n7665)
         );
  NAND2_X1 U9760 ( .A1(n8189), .A2(n8188), .ZN(n15081) );
  INV_X2 U9761 ( .A(n7669), .ZN(n15000) );
  NOR2_X2 U9762 ( .A1(n7669), .A2(n7534), .ZN(n14943) );
  NAND2_X1 U9763 ( .A1(n11097), .A2(n12542), .ZN(n7674) );
  NOR2_X1 U9764 ( .A1(n14857), .A2(n12544), .ZN(n7676) );
  INV_X1 U9765 ( .A(n10123), .ZN(n14860) );
  NAND3_X1 U9766 ( .A1(n10526), .A2(n7452), .A3(n9852), .ZN(n10014) );
  NAND3_X1 U9767 ( .A1(n10526), .A2(n7452), .A3(n7570), .ZN(n7686) );
  NAND2_X1 U9768 ( .A1(n7688), .A2(n8819), .ZN(n7692) );
  NAND3_X1 U9769 ( .A1(n7692), .A2(n8842), .A3(n7691), .ZN(n8729) );
  NAND3_X1 U9770 ( .A1(n8744), .A2(n8746), .A3(n8745), .ZN(n7706) );
  NAND2_X1 U9771 ( .A1(n7706), .A2(n7708), .ZN(n8748) );
  NAND2_X1 U9772 ( .A1(n7715), .A2(n8742), .ZN(n8743) );
  NAND2_X1 U9773 ( .A1(n7720), .A2(n8762), .ZN(n8763) );
  NAND2_X1 U9774 ( .A1(n8764), .A2(n8216), .ZN(n9136) );
  NAND2_X1 U9775 ( .A1(n7720), .A2(n7608), .ZN(n8216) );
  INV_X1 U9776 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7719) );
  NAND2_X1 U9777 ( .A1(n8392), .A2(n7724), .ZN(n7722) );
  NAND3_X1 U9778 ( .A1(n7722), .A2(n7721), .A3(n8382), .ZN(n9241) );
  INV_X1 U9779 ( .A(n13897), .ZN(n9247) );
  OR2_X2 U9780 ( .A1(n10192), .A2(n7737), .ZN(n7736) );
  NAND2_X2 U9781 ( .A1(n7428), .A2(n7738), .ZN(n12866) );
  NAND2_X1 U9782 ( .A1(n9251), .A2(n7745), .ZN(n7744) );
  NAND3_X1 U9783 ( .A1(n9051), .A2(n8652), .A3(n7750), .ZN(n7752) );
  XNOR2_X2 U9784 ( .A(n7751), .B(P3_IR_REG_27__SCAN_IN), .ZN(n13038) );
  NAND2_X1 U9785 ( .A1(n9465), .A2(n7756), .ZN(n7754) );
  NOR2_X1 U9786 ( .A1(n7505), .A2(n7815), .ZN(n7814) );
  NAND3_X1 U9787 ( .A1(n7813), .A2(n7571), .A3(n7765), .ZN(n7764) );
  OR2_X1 U9788 ( .A1(n7505), .A2(n7766), .ZN(n7765) );
  OR2_X1 U9789 ( .A1(n7815), .A2(n13441), .ZN(n7766) );
  NAND2_X1 U9790 ( .A1(n10659), .A2(n10658), .ZN(n7776) );
  NAND2_X1 U9791 ( .A1(n11762), .A2(n7778), .ZN(n7777) );
  NAND2_X1 U9792 ( .A1(n7777), .A2(n7780), .ZN(n11836) );
  NAND2_X1 U9793 ( .A1(n7787), .A2(n7785), .ZN(n10677) );
  NAND2_X1 U9794 ( .A1(n11830), .A2(n7791), .ZN(n7792) );
  NAND3_X1 U9795 ( .A1(n9547), .A2(n14314), .A3(n9562), .ZN(n7793) );
  NAND2_X2 U9796 ( .A1(n9654), .A2(n7486), .ZN(n14268) );
  NAND2_X1 U9797 ( .A1(n14404), .A2(n7558), .ZN(n7802) );
  NAND2_X1 U9798 ( .A1(n14404), .A2(n8299), .ZN(n7806) );
  NAND3_X1 U9799 ( .A1(n7808), .A2(n7807), .A3(n10671), .ZN(n10555) );
  NAND3_X1 U9800 ( .A1(n7822), .A2(n7821), .A3(n7820), .ZN(n7827) );
  NAND2_X1 U9801 ( .A1(n8432), .A2(n7823), .ZN(n7820) );
  NAND3_X1 U9802 ( .A1(n7822), .A2(n7825), .A3(n7820), .ZN(n11457) );
  INV_X1 U9803 ( .A(n7827), .ZN(n13625) );
  NAND3_X1 U9804 ( .A1(n7831), .A2(n7833), .A3(n7830), .ZN(n10960) );
  NAND3_X1 U9805 ( .A1(n7831), .A2(n7456), .A3(n7830), .ZN(n7834) );
  INV_X1 U9806 ( .A(n7834), .ZN(n11122) );
  NAND2_X1 U9807 ( .A1(n7837), .A2(n7555), .ZN(n7836) );
  NAND2_X1 U9808 ( .A1(n7839), .A2(n7838), .ZN(n7837) );
  NAND2_X1 U9809 ( .A1(n13236), .A2(n13235), .ZN(n7838) );
  OAI21_X1 U9810 ( .B1(n13236), .B2(n13235), .A(n13234), .ZN(n7839) );
  NAND2_X1 U9811 ( .A1(n9619), .A2(n7841), .ZN(n7840) );
  NAND2_X1 U9812 ( .A1(n7840), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9628) );
  NAND2_X1 U9813 ( .A1(n7842), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10827) );
  NAND3_X1 U9814 ( .A1(n13175), .A2(n8100), .A3(n13174), .ZN(n7848) );
  NAND4_X2 U9815 ( .A1(n10793), .A2(n13350), .A3(n13093), .A4(n14301), .ZN(
        n13349) );
  INV_X1 U9816 ( .A(n7849), .ZN(n13091) );
  NAND2_X1 U9817 ( .A1(n13260), .A2(n7859), .ZN(n8111) );
  NAND2_X1 U9818 ( .A1(n7854), .A2(n7851), .ZN(n13291) );
  NAND2_X1 U9819 ( .A1(n7859), .A2(n13261), .ZN(n7853) );
  NAND2_X1 U9820 ( .A1(n13260), .A2(n7855), .ZN(n7854) );
  INV_X1 U9821 ( .A(n13261), .ZN(n7858) );
  NAND2_X1 U9822 ( .A1(n7861), .A2(n7860), .ZN(n13170) );
  NAND3_X1 U9823 ( .A1(n13159), .A2(n7862), .A3(n8701), .ZN(n7861) );
  NAND3_X1 U9824 ( .A1(n8701), .A2(n7865), .A3(n7864), .ZN(n7863) );
  NAND2_X1 U9825 ( .A1(n13199), .A2(n8118), .ZN(n7866) );
  NAND2_X1 U9826 ( .A1(n7866), .A2(n7867), .ZN(n7869) );
  NAND2_X1 U9827 ( .A1(n7869), .A2(n7573), .ZN(n13212) );
  INV_X1 U9828 ( .A(n12818), .ZN(n7872) );
  INV_X1 U9829 ( .A(n12819), .ZN(n7873) );
  NAND2_X1 U9830 ( .A1(n13483), .A2(n7599), .ZN(n7880) );
  NAND3_X1 U9831 ( .A1(n7880), .A2(n7881), .A3(n12829), .ZN(n7874) );
  NAND3_X1 U9832 ( .A1(n7880), .A2(n7881), .A3(n7878), .ZN(n7877) );
  INV_X1 U9833 ( .A(n13537), .ZN(n7882) );
  NAND2_X1 U9834 ( .A1(n11303), .A2(n7883), .ZN(n11613) );
  INV_X1 U9835 ( .A(n8058), .ZN(n7884) );
  NAND3_X1 U9836 ( .A1(n11204), .A2(n10765), .A3(n10766), .ZN(n7885) );
  NAND2_X1 U9837 ( .A1(n10765), .A2(n10766), .ZN(n11030) );
  INV_X1 U9838 ( .A(n12164), .ZN(n7889) );
  INV_X1 U9839 ( .A(n7894), .ZN(n13578) );
  OAI211_X1 U9840 ( .C1(n13584), .C2(n7897), .A(n7895), .B(n8062), .ZN(
        P3_U3154) );
  NAND2_X1 U9841 ( .A1(n12792), .A2(n8022), .ZN(n8021) );
  NAND3_X1 U9842 ( .A1(n12681), .A2(n7564), .A3(n12680), .ZN(n7903) );
  NAND2_X1 U9843 ( .A1(n9386), .A2(n9385), .ZN(n7908) );
  NAND3_X1 U9844 ( .A1(n9386), .A2(n9385), .A3(n9408), .ZN(n7905) );
  NAND2_X1 U9845 ( .A1(n9515), .A2(n9514), .ZN(n7909) );
  NAND2_X1 U9846 ( .A1(n12625), .A2(n7918), .ZN(n7915) );
  OR2_X1 U9847 ( .A1(n12625), .A2(n7919), .ZN(n7916) );
  NAND2_X1 U9848 ( .A1(n7915), .A2(n7914), .ZN(n12629) );
  NAND2_X1 U9849 ( .A1(n12659), .A2(n7923), .ZN(n7922) );
  NAND3_X1 U9850 ( .A1(n12652), .A2(n8018), .A3(n7602), .ZN(n7926) );
  NAND2_X1 U9851 ( .A1(n7926), .A2(n7927), .ZN(n8538) );
  NOR2_X1 U9852 ( .A1(n7512), .A2(n7928), .ZN(n7927) );
  NAND2_X1 U9853 ( .A1(n7934), .A2(n7931), .ZN(n12642) );
  NAND3_X1 U9854 ( .A1(n12635), .A2(n7935), .A3(n7483), .ZN(n7934) );
  NAND3_X1 U9855 ( .A1(n7948), .A2(n7945), .A3(n15773), .ZN(n7944) );
  OAI21_X1 U9856 ( .B1(n15863), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n7553), .ZN(
        n7949) );
  XNOR2_X1 U9857 ( .A(n15725), .B(n15724), .ZN(n15863) );
  NAND2_X1 U9858 ( .A1(n15865), .A2(n15866), .ZN(n8573) );
  INV_X1 U9859 ( .A(n15874), .ZN(n7953) );
  INV_X1 U9860 ( .A(n15870), .ZN(n7955) );
  INV_X1 U9861 ( .A(n15877), .ZN(n7957) );
  XNOR2_X1 U9862 ( .A(n15736), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15869) );
  INV_X1 U9863 ( .A(n15884), .ZN(n7964) );
  OAI21_X2 U9864 ( .B1(n7445), .B2(n14713), .A(n7967), .ZN(n14768) );
  AND2_X1 U9865 ( .A1(n10104), .A2(n7968), .ZN(n9350) );
  NAND2_X1 U9866 ( .A1(n10104), .A2(n9347), .ZN(n9348) );
  NAND2_X1 U9867 ( .A1(n8277), .A2(n14619), .ZN(n14537) );
  NOR2_X2 U9868 ( .A1(n10434), .A2(n13146), .ZN(n10214) );
  NOR2_X2 U9869 ( .A1(n16392), .A2(n11907), .ZN(n11906) );
  NAND2_X1 U9870 ( .A1(n11262), .A2(n11282), .ZN(n11263) );
  AOI211_X2 U9871 ( .C1(n14563), .C2(n14332), .A(n14445), .B(n7458), .ZN(
        n14562) );
  NAND2_X1 U9872 ( .A1(n9909), .A2(n9908), .ZN(n10217) );
  OAI21_X1 U9873 ( .B1(n11836), .B2(n11835), .A(n11837), .ZN(n11920) );
  NAND2_X1 U9874 ( .A1(n11337), .A2(n11336), .ZN(n11762) );
  OAI22_X1 U9875 ( .A1(n14498), .A2(n14501), .B1(n14667), .B2(n14343), .ZN(
        n14483) );
  AND3_X2 U9876 ( .A1(n10084), .A2(n10086), .A3(n10085), .ZN(n10123) );
  NAND2_X1 U9877 ( .A1(n10796), .A2(n10795), .ZN(n11247) );
  NAND2_X1 U9878 ( .A1(n10217), .A2(n10216), .ZN(n10536) );
  AND2_X2 U9879 ( .A1(n15243), .A2(n10081), .ZN(n10089) );
  INV_X1 U9880 ( .A(n10737), .ZN(n10734) );
  NAND2_X1 U9881 ( .A1(n11238), .A2(n11237), .ZN(n11488) );
  OAI21_X1 U9882 ( .B1(n12630), .B2(n12631), .A(n7568), .ZN(n7994) );
  INV_X1 U9883 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n8402) );
  NAND2_X1 U9884 ( .A1(n12736), .A2(n12607), .ZN(n8520) );
  OAI21_X1 U9885 ( .B1(n7494), .B2(n7994), .A(n8525), .ZN(n12635) );
  NAND3_X1 U9886 ( .A1(n8516), .A2(n8515), .A3(n7556), .ZN(n12620) );
  NAND2_X1 U9887 ( .A1(n10890), .A2(n8337), .ZN(n11044) );
  INV_X1 U9888 ( .A(n10081), .ZN(n12308) );
  NAND2_X1 U9889 ( .A1(n7977), .A2(n8517), .ZN(n8515) );
  INV_X1 U9890 ( .A(n12604), .ZN(n7977) );
  NAND2_X1 U9891 ( .A1(n12600), .A2(n12599), .ZN(n12604) );
  NAND2_X1 U9892 ( .A1(n8083), .A2(n7561), .ZN(n14966) );
  NAND2_X1 U9893 ( .A1(n8084), .A2(n10861), .ZN(n16136) );
  NAND2_X1 U9894 ( .A1(n15221), .A2(n16391), .ZN(n8365) );
  NAND2_X1 U9895 ( .A1(n10733), .A2(n8015), .ZN(n10972) );
  NAND2_X1 U9896 ( .A1(n10975), .A2(n10974), .ZN(n11014) );
  NAND2_X1 U9897 ( .A1(n11234), .A2(n14862), .ZN(n10162) );
  NAND2_X1 U9898 ( .A1(n7986), .A2(n10092), .ZN(n14862) );
  XNOR2_X1 U9899 ( .A(n10231), .B(n10229), .ZN(n10305) );
  INV_X1 U9900 ( .A(n8061), .ZN(n14134) );
  INV_X1 U9901 ( .A(n8454), .ZN(n8453) );
  NAND2_X1 U9902 ( .A1(n14165), .A2(n8467), .ZN(n8465) );
  NOR2_X2 U9903 ( .A1(n13673), .A2(n7978), .ZN(n13705) );
  NOR2_X2 U9904 ( .A1(n13666), .A2(n13665), .ZN(n13673) );
  NOR2_X1 U9905 ( .A1(n13721), .A2(n13709), .ZN(n7979) );
  NAND2_X1 U9906 ( .A1(n7980), .A2(n13657), .ZN(n13658) );
  NAND2_X1 U9907 ( .A1(n8064), .A2(n8283), .ZN(n7980) );
  NOR2_X1 U9908 ( .A1(n10946), .A2(n16278), .ZN(n11110) );
  NOR2_X1 U9909 ( .A1(n16236), .A2(n10561), .ZN(n10692) );
  NOR2_X1 U9910 ( .A1(n11113), .A2(n11112), .ZN(n11454) );
  NAND3_X1 U9911 ( .A1(n12968), .A2(n7981), .A3(n13757), .ZN(n12972) );
  NAND3_X1 U9912 ( .A1(n12967), .A2(n12965), .A3(n12966), .ZN(n7981) );
  AND2_X1 U9913 ( .A1(n7450), .A2(n7982), .ZN(n13022) );
  NOR2_X1 U9914 ( .A1(n13020), .A2(n7502), .ZN(n7982) );
  NAND2_X1 U9915 ( .A1(n12979), .A2(n12980), .ZN(n12981) );
  NOR2_X1 U9916 ( .A1(n13035), .A2(n13034), .ZN(n8209) );
  NAND2_X1 U9917 ( .A1(n10972), .A2(n7559), .ZN(n11013) );
  INV_X1 U9918 ( .A(n14859), .ZN(n10860) );
  NAND3_X1 U9919 ( .A1(n10099), .A2(n8521), .A3(n7983), .ZN(n14859) );
  NAND2_X1 U9920 ( .A1(n11175), .A2(n11174), .ZN(n11228) );
  NAND2_X1 U9921 ( .A1(n11230), .A2(n11229), .ZN(n11238) );
  NAND2_X1 U9922 ( .A1(n7987), .A2(n10232), .ZN(n10728) );
  NAND2_X1 U9923 ( .A1(n10305), .A2(n10306), .ZN(n7987) );
  OAI211_X1 U9924 ( .C1(n15116), .C2(n16190), .A(n8089), .B(n8366), .ZN(n15221) );
  NAND2_X2 U9925 ( .A1(n10157), .A2(n10933), .ZN(n10228) );
  OAI22_X1 U9926 ( .A1(n10860), .A2(n10228), .B1(n11965), .B2(n10859), .ZN(
        n10233) );
  OAI211_X1 U9927 ( .C1(n9360), .C2(P2_DATAO_REG_0__SCAN_IN), .A(n7988), .B(
        SI_0_), .ZN(n9377) );
  NAND3_X1 U9928 ( .A1(n7535), .A2(n12580), .A3(n8534), .ZN(n7992) );
  INV_X1 U9929 ( .A(n10089), .ZN(n12018) );
  NAND4_X1 U9930 ( .A1(n12558), .A2(n12557), .A3(n12559), .A4(n7989), .ZN(
        n12560) );
  NAND2_X1 U9931 ( .A1(n7992), .A2(n7990), .ZN(n12586) );
  NAND2_X1 U9932 ( .A1(n9360), .A2(n9402), .ZN(n7993) );
  OAI21_X1 U9933 ( .B1(n9867), .B2(n9866), .A(n9870), .ZN(n10242) );
  NAND2_X1 U9934 ( .A1(n8020), .A2(n8019), .ZN(n8018) );
  OAI21_X1 U9935 ( .B1(n8636), .B2(n11029), .A(n11207), .ZN(n8058) );
  NAND2_X1 U9936 ( .A1(n8023), .A2(n13526), .ZN(n13529) );
  INV_X2 U9937 ( .A(n12988), .ZN(n9263) );
  NAND2_X1 U9938 ( .A1(n12545), .A2(n7995), .ZN(n12550) );
  NAND2_X1 U9939 ( .A1(n12553), .A2(n7557), .ZN(n7995) );
  NAND2_X1 U9940 ( .A1(n7997), .A2(n7996), .ZN(n8010) );
  OAI21_X1 U9941 ( .B1(n12564), .B2(n12563), .A(n12562), .ZN(n7997) );
  NAND2_X1 U9942 ( .A1(n12647), .A2(n12646), .ZN(n12651) );
  INV_X1 U9943 ( .A(n12651), .ZN(n8020) );
  NAND2_X1 U9944 ( .A1(n8630), .A2(n8632), .ZN(n8628) );
  NAND2_X1 U9945 ( .A1(n11613), .A2(n11612), .ZN(n11624) );
  NAND2_X1 U9946 ( .A1(n8074), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9276) );
  AND2_X2 U9947 ( .A1(n8279), .A2(n7552), .ZN(n13666) );
  XNOR2_X1 U9948 ( .A(n13663), .B(n13662), .ZN(n15986) );
  NAND2_X1 U9949 ( .A1(n13753), .A2(n13752), .ZN(n13751) );
  INV_X1 U9950 ( .A(n11671), .ZN(n9236) );
  NAND2_X1 U9951 ( .A1(n13940), .A2(n13939), .ZN(n13938) );
  OAI21_X1 U9952 ( .B1(n9323), .B2(n9309), .A(n9314), .ZN(P3_U3488) );
  OAI21_X1 U9953 ( .B1(n9323), .B2(n16415), .A(n8028), .ZN(P3_U3456) );
  AOI21_X1 U9954 ( .B1(n7434), .B2(n10101), .A(n7999), .ZN(n7998) );
  NOR2_X1 U9955 ( .A1(n11830), .A2(n9723), .ZN(n7999) );
  NAND2_X1 U9956 ( .A1(n8158), .A2(n8402), .ZN(n8157) );
  NAND2_X1 U9957 ( .A1(n11277), .A2(n8611), .ZN(n11337) );
  NAND2_X1 U9958 ( .A1(n10677), .A2(n10675), .ZN(n10540) );
  NAND2_X1 U9959 ( .A1(n8079), .A2(n9426), .ZN(n9446) );
  NAND3_X1 U9960 ( .A1(n9369), .A2(n9368), .A3(n9367), .ZN(n9375) );
  OR2_X1 U9961 ( .A1(n13194), .A2(n13193), .ZN(n13199) );
  NAND2_X1 U9962 ( .A1(n8130), .A2(n8128), .ZN(n8126) );
  NAND2_X1 U9963 ( .A1(n13292), .A2(n8682), .ZN(n8681) );
  OAI21_X1 U9964 ( .B1(n8693), .B2(n8692), .A(n8694), .ZN(n13230) );
  AOI21_X1 U9965 ( .B1(n8094), .B2(n13147), .A(n13143), .ZN(n8092) );
  NAND3_X2 U9966 ( .A1(n9332), .A2(n9494), .A3(n9396), .ZN(n8056) );
  AOI21_X1 U9967 ( .B1(n13233), .B2(n13232), .A(n13231), .ZN(n13236) );
  INV_X1 U9968 ( .A(n12000), .ZN(n8347) );
  INV_X1 U9969 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8794) );
  NAND2_X1 U9970 ( .A1(n8126), .A2(n8127), .ZN(n13454) );
  INV_X1 U9971 ( .A(n13243), .ZN(n13246) );
  NAND2_X1 U9972 ( .A1(n13140), .A2(n13139), .ZN(n8094) );
  OAI211_X1 U9973 ( .C1(n15112), .C2(n16190), .A(n8034), .B(n8033), .ZN(n15220) );
  NAND2_X1 U9974 ( .A1(n8695), .A2(n7550), .ZN(n8692) );
  NAND2_X1 U9975 ( .A1(n8325), .A2(n8324), .ZN(n13068) );
  OAI21_X1 U9976 ( .B1(n8093), .B2(n8092), .A(n13152), .ZN(n13159) );
  NAND2_X1 U9977 ( .A1(n13212), .A2(n13211), .ZN(n8096) );
  NAND2_X1 U9978 ( .A1(n8010), .A2(n8030), .ZN(n12574) );
  NAND2_X1 U9979 ( .A1(n12560), .A2(n8011), .ZN(n12564) );
  NAND2_X1 U9980 ( .A1(n12549), .A2(n12550), .ZN(n8011) );
  NAND2_X1 U9981 ( .A1(n11725), .A2(n11724), .ZN(n11880) );
  NAND2_X1 U9982 ( .A1(n14435), .A2(n8055), .ZN(n14351) );
  NAND3_X1 U9983 ( .A1(n14815), .A2(n14819), .A3(n12385), .ZN(n8552) );
  NAND2_X1 U9984 ( .A1(n10089), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8521) );
  NAND2_X1 U9985 ( .A1(n14483), .A2(n7569), .ZN(n8066) );
  NAND2_X1 U9986 ( .A1(n12806), .A2(n8024), .ZN(n8023) );
  INV_X1 U9987 ( .A(n9282), .ZN(n11393) );
  INV_X1 U9988 ( .A(n10458), .ZN(n8627) );
  NAND2_X2 U9989 ( .A1(n9949), .A2(n10095), .ZN(n8874) );
  NAND2_X4 U9990 ( .A1(n13037), .A2(n8634), .ZN(n9949) );
  NAND4_X2 U9991 ( .A1(n8853), .A2(n8852), .A3(n8851), .A4(n8850), .ZN(n13620)
         );
  AND2_X1 U9992 ( .A1(n8014), .A2(n10227), .ZN(n10306) );
  NAND2_X1 U9993 ( .A1(n10226), .A2(n12203), .ZN(n8014) );
  INV_X1 U9994 ( .A(n13675), .ZN(n8027) );
  NAND2_X1 U9995 ( .A1(n9051), .A2(n8652), .ZN(n9278) );
  NAND2_X1 U9996 ( .A1(n11617), .A2(n11616), .ZN(n11854) );
  AOI21_X1 U9997 ( .B1(n13550), .B2(n12815), .A(n7563), .ZN(n13501) );
  NOR2_X1 U9998 ( .A1(n10293), .A2(n8864), .ZN(n10506) );
  AOI21_X1 U9999 ( .B1(P3_REG2_REG_14__SCAN_IN), .B2(n15958), .A(n15969), .ZN(
        n13630) );
  NOR2_X1 U10000 ( .A1(n13628), .A2(n15940), .ZN(n15968) );
  OAI211_X1 U10001 ( .C1(n12792), .C2(n12791), .A(n8021), .B(n12790), .ZN(
        P1_U3242) );
  NAND2_X1 U10002 ( .A1(n8326), .A2(n15025), .ZN(n8325) );
  NAND2_X1 U10003 ( .A1(n14936), .A2(n14935), .ZN(n15113) );
  NAND2_X1 U10004 ( .A1(n13070), .A2(n7551), .ZN(n14950) );
  NAND2_X1 U10005 ( .A1(n7591), .A2(n12736), .ZN(n11779) );
  NAND3_X1 U10006 ( .A1(n8386), .A2(n9227), .A3(n9228), .ZN(n11217) );
  NAND2_X1 U10007 ( .A1(n8552), .A2(n8553), .ZN(n14756) );
  OAI21_X1 U10008 ( .B1(n12536), .B2(n14829), .A(n7598), .ZN(P1_U3220) );
  NOR2_X2 U10009 ( .A1(n8844), .A2(n8389), .ZN(n8871) );
  NAND2_X1 U10010 ( .A1(n14706), .A2(n12371), .ZN(n8172) );
  NAND2_X1 U10011 ( .A1(n8085), .A2(n10124), .ZN(n10858) );
  NAND2_X1 U10012 ( .A1(n8365), .A2(n8363), .ZN(P1_U3524) );
  NAND2_X1 U10013 ( .A1(n8444), .A2(n8443), .ZN(n13718) );
  INV_X1 U10014 ( .A(n8031), .ZN(n8030) );
  OAI21_X1 U10015 ( .B1(n12568), .B2(n12567), .A(n12566), .ZN(n8031) );
  NAND2_X1 U10016 ( .A1(n12667), .A2(n12663), .ZN(n12666) );
  AOI21_X1 U10017 ( .B1(n8248), .B2(n8249), .A(n8247), .ZN(P3_U3296) );
  INV_X1 U10018 ( .A(n15040), .ZN(n8326) );
  NAND2_X1 U10019 ( .A1(n12181), .A2(n12180), .ZN(n12252) );
  NAND2_X1 U10020 ( .A1(n9148), .A2(n9147), .ZN(n9150) );
  NAND2_X1 U10021 ( .A1(n8353), .A2(n8352), .ZN(n14969) );
  NAND2_X1 U10022 ( .A1(n8748), .A2(n8747), .ZN(n9033) );
  INV_X1 U10023 ( .A(n8346), .ZN(n8345) );
  NAND2_X1 U10024 ( .A1(n12255), .A2(n12254), .ZN(n13060) );
  NAND2_X1 U10025 ( .A1(n8344), .A2(n8343), .ZN(n12179) );
  NOR2_X1 U10026 ( .A1(n8035), .A2(n13743), .ZN(n9323) );
  NAND2_X1 U10027 ( .A1(n8729), .A2(n8728), .ZN(n8855) );
  NAND2_X1 U10028 ( .A1(n8228), .A2(n8229), .ZN(n8940) );
  NAND2_X1 U10029 ( .A1(n10857), .A2(n10858), .ZN(n8084) );
  NAND2_X1 U10030 ( .A1(n12819), .A2(n12818), .ZN(n12820) );
  NAND2_X1 U10031 ( .A1(n9051), .A2(n8653), .ZN(n8074) );
  NAND2_X1 U10032 ( .A1(n13529), .A2(n12809), .ZN(n13579) );
  NAND2_X1 U10033 ( .A1(n11204), .A2(n11035), .ZN(n8057) );
  NAND2_X1 U10034 ( .A1(n8978), .A2(n8236), .ZN(n8234) );
  AOI21_X2 U10035 ( .B1(n14273), .B2(P2_REG2_REG_16__SCAN_IN), .A(n14272), 
        .ZN(n14275) );
  XNOR2_X1 U10036 ( .A(n8043), .B(n8042), .ZN(n14309) );
  AND2_X1 U10037 ( .A1(n14295), .A2(n14294), .ZN(n8044) );
  NAND2_X1 U10038 ( .A1(n8160), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n8159) );
  NAND2_X1 U10039 ( .A1(n8045), .A2(n8536), .ZN(n12676) );
  NAND3_X1 U10040 ( .A1(n12671), .A2(n12670), .A3(n7600), .ZN(n8045) );
  NAND2_X1 U10041 ( .A1(n15973), .A2(n15972), .ZN(n15971) );
  NOR2_X2 U10042 ( .A1(n15989), .A2(n15990), .ZN(n15988) );
  NAND3_X1 U10043 ( .A1(n13732), .A2(n8048), .A3(n7547), .ZN(P3_U3201) );
  NAND2_X1 U10044 ( .A1(n8562), .A2(n8565), .ZN(n15764) );
  NAND2_X1 U10045 ( .A1(n8738), .A2(n8737), .ZN(n8952) );
  OAI21_X1 U10046 ( .B1(n14038), .B2(n9309), .A(n8053), .ZN(n13973) );
  OAI21_X1 U10047 ( .B1(n13814), .B2(n8373), .A(n8371), .ZN(n9260) );
  OAI211_X1 U10048 ( .C1(n13753), .C2(n13752), .A(n13751), .B(n16054), .ZN(
        n13756) );
  OR2_X1 U10049 ( .A1(n10540), .A2(n10554), .ZN(n10796) );
  NAND2_X1 U10050 ( .A1(n13515), .A2(n8071), .ZN(n12806) );
  NAND2_X1 U10051 ( .A1(n13626), .A2(n13638), .ZN(n13627) );
  XNOR2_X1 U10052 ( .A(n13627), .B(n15944), .ZN(n15941) );
  NAND2_X1 U10053 ( .A1(n13631), .A2(n8437), .ZN(n8433) );
  XNOR2_X2 U10054 ( .A(n8834), .B(P3_IR_REG_2__SCAN_IN), .ZN(n10076) );
  NOR2_X1 U10055 ( .A1(n15923), .A2(n15922), .ZN(n15921) );
  INV_X1 U10057 ( .A(n8473), .ZN(n8472) );
  XNOR2_X2 U10058 ( .A(n11109), .B(n11121), .ZN(n10946) );
  NAND2_X1 U10059 ( .A1(n11455), .A2(n8284), .ZN(n8064) );
  NOR2_X2 U10060 ( .A1(n13707), .A2(n13708), .ZN(n13711) );
  NOR2_X2 U10061 ( .A1(n13674), .A2(n14011), .ZN(n13707) );
  NOR2_X1 U10062 ( .A1(n10692), .A2(n10693), .ZN(n10696) );
  NAND2_X1 U10063 ( .A1(n11920), .A2(n7816), .ZN(n11922) );
  NAND3_X1 U10064 ( .A1(n8070), .A2(n8069), .A3(n14529), .ZN(n8068) );
  NOR2_X1 U10065 ( .A1(n10709), .A2(n10710), .ZN(n10713) );
  AOI21_X1 U10066 ( .B1(n13956), .B2(n12797), .A(n8717), .ZN(n13940) );
  OAI22_X1 U10067 ( .A1(n13872), .A2(n9249), .B1(n13878), .B2(n13574), .ZN(
        n13861) );
  NAND4_X1 U10068 ( .A1(n8785), .A2(n8784), .A3(n8783), .A4(n9205), .ZN(n8786)
         );
  AOI21_X1 U10069 ( .B1(n8075), .B2(n15835), .A(n14307), .ZN(n14308) );
  XNOR2_X1 U10070 ( .A(n14303), .B(n14302), .ZN(n8075) );
  NAND2_X1 U10071 ( .A1(n9424), .A2(n8076), .ZN(n8077) );
  NAND2_X1 U10072 ( .A1(n8077), .A2(n8078), .ZN(n9465) );
  INV_X1 U10073 ( .A(n8083), .ZN(n14982) );
  NAND2_X1 U10074 ( .A1(n10868), .A2(n8088), .ZN(n8676) );
  OR2_X1 U10075 ( .A1(n12316), .A2(n14867), .ZN(n8090) );
  NAND2_X1 U10076 ( .A1(n8097), .A2(n8096), .ZN(n13220) );
  NAND3_X1 U10077 ( .A1(n8097), .A2(n8096), .A3(n8095), .ZN(n8695) );
  NAND3_X1 U10078 ( .A1(n13175), .A2(n13174), .A3(n8099), .ZN(n8098) );
  NAND2_X1 U10079 ( .A1(n13199), .A2(n8116), .ZN(n8115) );
  INV_X1 U10080 ( .A(n13198), .ZN(n8120) );
  NAND2_X1 U10081 ( .A1(n8131), .A2(n8132), .ZN(n11322) );
  NAND2_X1 U10082 ( .A1(n9769), .A2(n8722), .ZN(n8143) );
  INV_X1 U10083 ( .A(n8147), .ZN(n10791) );
  NAND2_X1 U10084 ( .A1(n10524), .A2(n10523), .ZN(n10777) );
  NAND3_X1 U10085 ( .A1(n8796), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n8158) );
  NAND3_X1 U10086 ( .A1(n8795), .A2(n16002), .A3(n8794), .ZN(n8160) );
  XNOR2_X1 U10087 ( .A(n8171), .B(n12203), .ZN(n10231) );
  NAND2_X1 U10088 ( .A1(n10972), .A2(n10971), .ZN(n10975) );
  OAI21_X1 U10089 ( .B1(n14768), .B2(n8175), .A(n8173), .ZN(n14696) );
  XNOR2_X2 U10090 ( .A(n8181), .B(n9852), .ZN(n15245) );
  NOR2_X2 U10091 ( .A1(n14926), .A2(n13076), .ZN(n14918) );
  INV_X1 U10092 ( .A(n16077), .ZN(n8187) );
  NOR2_X2 U10093 ( .A1(n11603), .A2(n12601), .ZN(n16323) );
  OR2_X2 U10094 ( .A1(n11397), .A2(n12592), .ZN(n11603) );
  NAND2_X1 U10095 ( .A1(n12108), .A2(n8198), .ZN(n8197) );
  XNOR2_X1 U10096 ( .A(n8212), .B(n13021), .ZN(n8211) );
  NAND2_X1 U10097 ( .A1(n13622), .A2(n16116), .ZN(n12871) );
  NAND3_X1 U10098 ( .A1(n13465), .A2(n8803), .A3(P3_REG1_REG_0__SCAN_IN), .ZN(
        n8215) );
  NAND2_X1 U10099 ( .A1(n8217), .A2(n8218), .ZN(n8887) );
  NAND2_X1 U10100 ( .A1(n8756), .A2(n8222), .ZN(n8220) );
  OAI211_X1 U10101 ( .C1(n8756), .C2(n8224), .A(n8220), .B(
        P2_DATAO_REG_20__SCAN_IN), .ZN(n8227) );
  NAND2_X1 U10102 ( .A1(n8902), .A2(n8231), .ZN(n8228) );
  OAI211_X1 U10103 ( .C1(n8978), .C2(n8237), .A(n8234), .B(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n8745) );
  INV_X1 U10104 ( .A(n9164), .ZN(n8262) );
  NAND2_X1 U10105 ( .A1(n8261), .A2(n9163), .ZN(n8260) );
  NOR2_X1 U10106 ( .A1(n14473), .A2(n14599), .ZN(n8268) );
  INV_X1 U10107 ( .A(n8268), .ZN(n14457) );
  NOR2_X2 U10108 ( .A1(n10684), .A2(n16246), .ZN(n8271) );
  AND2_X1 U10109 ( .A1(n14396), .A2(n8276), .ZN(n14370) );
  NAND2_X1 U10110 ( .A1(n14396), .A2(n8272), .ZN(n14319) );
  NAND2_X1 U10111 ( .A1(n14396), .A2(n14383), .ZN(n14378) );
  NOR2_X2 U10112 ( .A1(n11846), .A2(n13221), .ZN(n12048) );
  XNOR2_X1 U10113 ( .A(n8278), .B(P3_IR_REG_1__SCAN_IN), .ZN(n10327) );
  OR2_X2 U10114 ( .A1(n15986), .A2(n15987), .ZN(n8279) );
  XNOR2_X1 U10115 ( .A(n13654), .B(n13655), .ZN(n11455) );
  INV_X1 U10116 ( .A(n8285), .ZN(n13656) );
  INV_X1 U10117 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n8323) );
  NAND2_X1 U10118 ( .A1(n8329), .A2(n12553), .ZN(n16138) );
  NAND2_X1 U10119 ( .A1(n10891), .A2(n12725), .ZN(n8329) );
  OAI211_X1 U10120 ( .C1(n10891), .C2(n8331), .A(n8330), .B(n10892), .ZN(
        n11106) );
  NAND2_X1 U10121 ( .A1(n10857), .A2(n8332), .ZN(n8330) );
  NAND2_X1 U10122 ( .A1(n10097), .A2(n12552), .ZN(n10891) );
  NAND2_X1 U10123 ( .A1(n8334), .A2(n8333), .ZN(n11361) );
  AOI21_X1 U10124 ( .B1(n8336), .B2(n8338), .A(n7429), .ZN(n8333) );
  NAND2_X1 U10125 ( .A1(n11049), .A2(n8336), .ZN(n8334) );
  NAND2_X1 U10126 ( .A1(n11784), .A2(n8345), .ZN(n8344) );
  AOI21_X1 U10127 ( .B1(n8345), .B2(n8347), .A(n7515), .ZN(n8343) );
  OAI21_X1 U10128 ( .B1(n11783), .B2(n8347), .A(n12073), .ZN(n8346) );
  NAND2_X1 U10129 ( .A1(n11579), .A2(n8349), .ZN(n8348) );
  CLKBUF_X1 U10130 ( .A(n8353), .Z(n8351) );
  NAND2_X1 U10131 ( .A1(n15075), .A2(n8359), .ZN(n8357) );
  OR2_X2 U10132 ( .A1(n13923), .A2(n13922), .ZN(n13925) );
  INV_X1 U10133 ( .A(n14058), .ZN(n8380) );
  AOI21_X1 U10134 ( .B1(n8385), .B2(n8383), .A(n7478), .ZN(n8382) );
  OR2_X1 U10135 ( .A1(n8430), .A2(n8387), .ZN(n10066) );
  OR2_X1 U10136 ( .A1(n8430), .A2(n8388), .ZN(n10061) );
  NAND2_X1 U10137 ( .A1(n9236), .A2(n8395), .ZN(n8392) );
  AOI21_X1 U10138 ( .B1(n8395), .B2(n8397), .A(n8394), .ZN(n8393) );
  NAND2_X1 U10139 ( .A1(n8792), .A2(n8801), .ZN(n8399) );
  NAND2_X1 U10140 ( .A1(n8400), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8789) );
  NOR2_X1 U10141 ( .A1(n13772), .A2(n13771), .ZN(n13769) );
  NAND2_X1 U10142 ( .A1(n9253), .A2(n9252), .ZN(n13823) );
  NAND2_X1 U10143 ( .A1(n13060), .A2(n13059), .ZN(n15075) );
  NAND2_X1 U10144 ( .A1(n11314), .A2(n13005), .ZN(n11313) );
  NOR2_X1 U10145 ( .A1(n8876), .A2(n8875), .ZN(n16199) );
  NAND2_X1 U10146 ( .A1(n9047), .A2(n9046), .ZN(n13902) );
  NAND2_X1 U10147 ( .A1(n12029), .A2(n8957), .ZN(n11994) );
  NAND2_X2 U10148 ( .A1(n9255), .A2(n9254), .ZN(n13814) );
  INV_X1 U10149 ( .A(n13001), .ZN(n9228) );
  NOR2_X2 U10150 ( .A1(n8847), .A2(n8846), .ZN(n11329) );
  NAND2_X1 U10151 ( .A1(n14932), .A2(n13072), .ZN(n13074) );
  NAND2_X1 U10152 ( .A1(n8822), .A2(n9455), .ZN(n8824) );
  XNOR2_X1 U10153 ( .A(n8401), .B(n9407), .ZN(n10865) );
  INV_X1 U10154 ( .A(n11322), .ZN(n8403) );
  NAND2_X1 U10155 ( .A1(n11527), .A2(n8407), .ZN(n11712) );
  NAND2_X1 U10156 ( .A1(n12692), .A2(n12691), .ZN(n8414) );
  NAND2_X1 U10157 ( .A1(n12474), .A2(n8426), .ZN(n12303) );
  OR2_X2 U10158 ( .A1(n11124), .A2(n11123), .ZN(n8432) );
  XNOR2_X1 U10159 ( .A(n13630), .B(n13662), .ZN(n15979) );
  INV_X1 U10160 ( .A(n8448), .ZN(n13692) );
  INV_X1 U10161 ( .A(n14137), .ZN(n8450) );
  NAND2_X1 U10162 ( .A1(n14158), .A2(n14157), .ZN(n8451) );
  NAND2_X1 U10163 ( .A1(n14127), .A2(n14128), .ZN(n8468) );
  OR2_X1 U10164 ( .A1(n8476), .A2(n11816), .ZN(n8470) );
  NAND2_X1 U10165 ( .A1(n14238), .A2(n7566), .ZN(n8483) );
  OAI211_X1 U10166 ( .C1(n14238), .C2(n8484), .A(n8483), .B(n14185), .ZN(
        P2_U3192) );
  NAND2_X1 U10167 ( .A1(n14238), .A2(n14150), .ZN(n14176) );
  INV_X1 U10168 ( .A(n9740), .ZN(n8503) );
  NAND2_X1 U10169 ( .A1(n8504), .A2(n8505), .ZN(n10918) );
  NAND2_X1 U10170 ( .A1(n10028), .A2(n8507), .ZN(n8504) );
  AOI21_X1 U10171 ( .B1(n8510), .B2(n8508), .A(n10616), .ZN(n8507) );
  NAND2_X1 U10172 ( .A1(n11506), .A2(n8514), .ZN(n11509) );
  INV_X1 U10173 ( .A(n8514), .ZN(n8513) );
  NAND2_X1 U10174 ( .A1(n12603), .A2(n8518), .ZN(n8516) );
  INV_X1 U10175 ( .A(n12602), .ZN(n8519) );
  NAND2_X1 U10176 ( .A1(n14859), .A2(n10859), .ZN(n12556) );
  OAI22_X1 U10177 ( .A1(n7432), .A2(n10102), .B1(n12316), .B2(n10103), .ZN(
        n8523) );
  INV_X1 U10178 ( .A(n12632), .ZN(n8527) );
  NAND2_X1 U10179 ( .A1(n12642), .A2(n12643), .ZN(n12641) );
  NAND3_X1 U10180 ( .A1(n12621), .A2(n7522), .A3(n8530), .ZN(n8529) );
  NAND2_X1 U10181 ( .A1(n8529), .A2(n8531), .ZN(n12625) );
  NAND2_X1 U10182 ( .A1(n8538), .A2(n8539), .ZN(n12659) );
  NAND2_X1 U10183 ( .A1(n12657), .A2(n12655), .ZN(n8539) );
  NAND3_X1 U10184 ( .A1(n9346), .A2(n9410), .A3(n8721), .ZN(n10821) );
  NOR2_X1 U10185 ( .A1(n15896), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n15766) );
  NAND2_X1 U10186 ( .A1(n8564), .A2(n8563), .ZN(n8562) );
  INV_X1 U10187 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8563) );
  INV_X1 U10188 ( .A(n15892), .ZN(n8565) );
  XNOR2_X1 U10189 ( .A(n8569), .B(n7477), .ZN(SUB_1596_U63) );
  NAND2_X1 U10190 ( .A1(n14407), .A2(n7444), .ZN(n8591) );
  NOR2_X1 U10191 ( .A1(n14349), .A2(n8605), .ZN(n8604) );
  NAND2_X1 U10192 ( .A1(n14483), .A2(n8604), .ZN(n8600) );
  OAI211_X1 U10193 ( .C1(n13584), .C2(n7572), .A(n8621), .B(n8619), .ZN(n12846) );
  OAI22_X1 U10194 ( .A1(n8623), .A2(n8620), .B1(n12839), .B2(n8625), .ZN(n8619) );
  NOR2_X1 U10195 ( .A1(n12839), .A2(n13466), .ZN(n8620) );
  NAND2_X1 U10196 ( .A1(n13584), .A2(n8622), .ZN(n8621) );
  NOR2_X1 U10197 ( .A1(n8623), .A2(n12839), .ZN(n8622) );
  INV_X1 U10198 ( .A(n12839), .ZN(n8624) );
  NAND2_X1 U10199 ( .A1(n16051), .A2(n10459), .ZN(n8632) );
  NAND2_X1 U10200 ( .A1(n8628), .A2(n8631), .ZN(n10626) );
  MUX2_X1 U10201 ( .A(P3_REG1_REG_1__SCAN_IN), .B(P3_REG2_REG_1__SCAN_IN), .S(
        n8633), .Z(n10074) );
  MUX2_X1 U10202 ( .A(n8387), .B(n8388), .S(n8633), .Z(n9953) );
  MUX2_X1 U10203 ( .A(P3_REG1_REG_2__SCAN_IN), .B(P3_REG2_REG_2__SCAN_IN), .S(
        n8633), .Z(n10259) );
  MUX2_X1 U10204 ( .A(P3_REG1_REG_3__SCAN_IN), .B(P3_REG2_REG_3__SCAN_IN), .S(
        n8633), .Z(n10287) );
  MUX2_X1 U10205 ( .A(P3_REG1_REG_4__SCAN_IN), .B(P3_REG2_REG_4__SCAN_IN), .S(
        n8633), .Z(n10292) );
  MUX2_X1 U10206 ( .A(P3_REG1_REG_5__SCAN_IN), .B(P3_REG2_REG_5__SCAN_IN), .S(
        n8633), .Z(n10489) );
  MUX2_X1 U10207 ( .A(P3_REG1_REG_7__SCAN_IN), .B(P3_REG2_REG_7__SCAN_IN), .S(
        n8633), .Z(n10563) );
  MUX2_X1 U10208 ( .A(n8909), .B(n8913), .S(n8633), .Z(n10698) );
  MUX2_X1 U10209 ( .A(n16278), .B(n10948), .S(n8633), .Z(n10949) );
  MUX2_X1 U10210 ( .A(n16317), .B(n11995), .S(n8633), .Z(n13635) );
  NOR2_X1 U10211 ( .A1(n11035), .A2(n8638), .ZN(n8637) );
  INV_X1 U10212 ( .A(n13473), .ZN(n8650) );
  INV_X1 U10213 ( .A(n8659), .ZN(n13057) );
  NAND2_X1 U10214 ( .A1(n8676), .A2(n12566), .ZN(n10983) );
  NAND2_X1 U10215 ( .A1(n13456), .A2(n13455), .ZN(n8686) );
  NAND3_X1 U10216 ( .A1(n8686), .A2(n8685), .A3(n8684), .ZN(P2_U3328) );
  AOI21_X1 U10217 ( .B1(n8711), .B2(n8710), .A(n8709), .ZN(n8708) );
  INV_X1 U10218 ( .A(n13240), .ZN(n8709) );
  INV_X1 U10219 ( .A(n13239), .ZN(n8712) );
  INV_X1 U10220 ( .A(n10104), .ZN(n10108) );
  AND2_X1 U10221 ( .A1(n10157), .A2(n9702), .ZN(n10168) );
  NOR2_X1 U10222 ( .A1(n10157), .A2(n9696), .ZN(P1_U4016) );
  NAND2_X1 U10223 ( .A1(n8956), .A2(n8394), .ZN(n12029) );
  OR2_X1 U10224 ( .A1(n9698), .A2(n15253), .ZN(n10132) );
  AND2_X1 U10225 ( .A1(n15253), .A2(n9693), .ZN(n9695) );
  INV_X1 U10226 ( .A(n10526), .ZN(n10248) );
  INV_X1 U10227 ( .A(n7427), .ZN(n12431) );
  INV_X1 U10228 ( .A(n8056), .ZN(n9619) );
  INV_X1 U10229 ( .A(n9742), .ZN(n13346) );
  OR2_X1 U10230 ( .A1(n16415), .A2(n16311), .ZN(n14102) );
  INV_X1 U10231 ( .A(n14102), .ZN(n9325) );
  NAND2_X2 U10232 ( .A1(n11094), .A2(n16113), .ZN(n16121) );
  INV_X1 U10233 ( .A(n14030), .ZN(n9313) );
  AND2_X2 U10234 ( .A1(n11090), .A2(n9308), .ZN(n16407) );
  INV_X1 U10235 ( .A(n8812), .ZN(n9097) );
  NOR2_X1 U10236 ( .A1(n9057), .A2(n9040), .ZN(n8715) );
  INV_X1 U10237 ( .A(n13901), .ZN(n9246) );
  AND2_X2 U10238 ( .A1(n13116), .A2(n9661), .ZN(n8716) );
  NAND2_X1 U10239 ( .A1(n10203), .A2(n14510), .ZN(n14549) );
  AND2_X1 U10240 ( .A1(n14101), .A2(n13475), .ZN(n8717) );
  AND2_X1 U10241 ( .A1(n14947), .A2(n13071), .ZN(n8718) );
  OR2_X1 U10242 ( .A1(n15132), .A2(n13054), .ZN(n8719) );
  OR2_X1 U10243 ( .A1(n15132), .A2(n14836), .ZN(n8720) );
  AND2_X2 U10244 ( .A1(n10932), .A2(n16161), .ZN(n16347) );
  INV_X1 U10245 ( .A(n16347), .ZN(n16159) );
  AND3_X1 U10246 ( .A1(n9845), .A2(n15649), .A3(n15650), .ZN(n8721) );
  INV_X1 U10247 ( .A(n13073), .ZN(n13056) );
  AND2_X1 U10248 ( .A1(n9770), .A2(n9717), .ZN(n8722) );
  OR2_X1 U10249 ( .A1(n14068), .A2(n13611), .ZN(n8723) );
  NAND2_X1 U10250 ( .A1(n13119), .A2(n9890), .ZN(n13117) );
  OAI21_X1 U10251 ( .B1(n13130), .B2(n13131), .A(n13129), .ZN(n13133) );
  INV_X1 U10252 ( .A(n13205), .ZN(n13206) );
  OR4_X1 U10253 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n10139) );
  INV_X1 U10254 ( .A(n13922), .ZN(n9244) );
  INV_X1 U10255 ( .A(n13769), .ZN(n13770) );
  INV_X1 U10256 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8783) );
  AND4_X1 U10257 ( .A1(n9618), .A2(n9535), .A3(n9534), .A4(n9533), .ZN(n9536)
         );
  INV_X1 U10258 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n15648) );
  INV_X1 U10259 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n13518) );
  OR2_X1 U10260 ( .A1(n9071), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9084) );
  OAI22_X1 U10261 ( .A1(n13776), .A2(n16103), .B1(n13734), .B2(n13025), .ZN(
        n9269) );
  AND2_X1 U10262 ( .A1(n14068), .A2(n13848), .ZN(n12962) );
  INV_X1 U10263 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10029) );
  NAND2_X1 U10264 ( .A1(n10793), .A2(n9660), .ZN(n13351) );
  OR2_X1 U10265 ( .A1(n9620), .A2(n9333), .ZN(n9334) );
  NAND2_X1 U10266 ( .A1(n10156), .A2(n14862), .ZN(n10159) );
  INV_X1 U10267 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n11365) );
  INV_X1 U10268 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9349) );
  INV_X1 U10269 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9347) );
  OR2_X1 U10270 ( .A1(n12808), .A2(n13913), .ZN(n12809) );
  INV_X1 U10271 ( .A(n10314), .ZN(n10453) );
  INV_X1 U10272 ( .A(n13752), .ZN(n13757) );
  OR2_X1 U10273 ( .A1(n9009), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9025) );
  INV_X1 U10274 ( .A(n10454), .ZN(n12863) );
  INV_X1 U10275 ( .A(n13000), .ZN(n9235) );
  NOR2_X1 U10276 ( .A1(n12279), .A2(n12278), .ZN(n13100) );
  INV_X1 U10277 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n9539) );
  NOR2_X1 U10278 ( .A1(n13298), .A2(n13297), .ZN(n13307) );
  OR2_X1 U10279 ( .A1(n11929), .A2(n11928), .ZN(n12279) );
  OR2_X1 U10280 ( .A1(n9885), .A2(n13350), .ZN(n9802) );
  INV_X1 U10281 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n11789) );
  OR2_X1 U10282 ( .A1(n12384), .A2(n12383), .ZN(n12385) );
  INV_X1 U10283 ( .A(n10974), .ZN(n10973) );
  NAND2_X1 U10284 ( .A1(n12402), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n12404) );
  INV_X1 U10285 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n12184) );
  AND2_X1 U10286 ( .A1(n12754), .A2(n12784), .ZN(n10936) );
  INV_X1 U10287 ( .A(n14787), .ZN(n14807) );
  NAND2_X1 U10288 ( .A1(n16332), .A2(n10944), .ZN(n10172) );
  INV_X1 U10289 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10525) );
  OR2_X1 U10290 ( .A1(n15730), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n15680) );
  OR2_X1 U10291 ( .A1(n9128), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9139) );
  AND2_X1 U10292 ( .A1(n8910), .A2(n10705), .ZN(n8927) );
  INV_X1 U10293 ( .A(n13801), .ZN(n13775) );
  NAND2_X1 U10294 ( .A1(n10463), .A2(n10462), .ZN(n13600) );
  INV_X1 U10295 ( .A(n13733), .ZN(n13021) );
  INV_X1 U10296 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n15349) );
  INV_X1 U10297 ( .A(n15983), .ZN(n13662) );
  INV_X1 U10298 ( .A(n15961), .ZN(n15982) );
  OR2_X1 U10299 ( .A1(n9120), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9128) );
  INV_X1 U10300 ( .A(n9223), .ZN(n12997) );
  NAND2_X1 U10301 ( .A1(n8860), .A2(n8859), .ZN(n11418) );
  AND2_X1 U10302 ( .A1(n11088), .A2(n11087), .ZN(n11089) );
  OR2_X1 U10303 ( .A1(n9500), .A2(n9300), .ZN(n9319) );
  AND2_X1 U10304 ( .A1(n9316), .A2(n13033), .ZN(n16107) );
  INV_X1 U10305 ( .A(n13943), .ZN(n16101) );
  AOI21_X1 U10306 ( .B1(n9175), .B2(n9173), .A(n8771), .ZN(n9191) );
  INV_X1 U10307 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n11819) );
  NAND2_X1 U10308 ( .A1(n11253), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n11338) );
  INV_X1 U10309 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10925) );
  INV_X1 U10310 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11705) );
  INV_X1 U10311 ( .A(n14195), .ZN(n14244) );
  AND2_X1 U10312 ( .A1(n13381), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n14333) );
  OR2_X1 U10313 ( .A1(n14413), .A2(n13309), .ZN(n13314) );
  NOR2_X1 U10314 ( .A1(n11765), .A2(n11959), .ZN(n11838) );
  INV_X1 U10315 ( .A(n9571), .ZN(n9558) );
  INV_X1 U10316 ( .A(n14523), .ZN(n14439) );
  AND2_X1 U10317 ( .A1(n9807), .A2(n9806), .ZN(n14486) );
  NAND2_X1 U10318 ( .A1(n9617), .A2(n9622), .ZN(n9625) );
  OR2_X1 U10319 ( .A1(n12404), .A2(n14779), .ZN(n12340) );
  INV_X1 U10320 ( .A(n12716), .ZN(n10151) );
  AND2_X1 U10321 ( .A1(n12328), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n12427) );
  INV_X1 U10322 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n15674) );
  INV_X1 U10323 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n15686) );
  INV_X1 U10324 ( .A(n12734), .ZN(n11600) );
  INV_X1 U10325 ( .A(n12729), .ZN(n11052) );
  NAND2_X1 U10326 ( .A1(n10112), .A2(n10944), .ZN(n16142) );
  AND2_X1 U10327 ( .A1(n16029), .A2(n10153), .ZN(n16366) );
  OR2_X1 U10328 ( .A1(n11098), .A2(n16038), .ZN(n16158) );
  INV_X1 U10329 ( .A(n10177), .ZN(n10145) );
  NAND2_X1 U10330 ( .A1(n12293), .A2(n12292), .ZN(n12457) );
  INV_X1 U10331 ( .A(n10821), .ZN(n10822) );
  OR2_X1 U10332 ( .A1(n8944), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8958) );
  NAND2_X1 U10333 ( .A1(n10339), .A2(n10338), .ZN(n13568) );
  INV_X1 U10334 ( .A(n13595), .ZN(n13606) );
  AND2_X1 U10335 ( .A1(n12995), .A2(n8808), .ZN(n12840) );
  INV_X1 U10336 ( .A(n15991), .ZN(n15970) );
  INV_X1 U10337 ( .A(n15984), .ZN(n13713) );
  INV_X1 U10338 ( .A(n13036), .ZN(n11093) );
  INV_X1 U10339 ( .A(n16407), .ZN(n9309) );
  NOR2_X1 U10340 ( .A1(n9309), .A2(n16274), .ZN(n16259) );
  AND3_X1 U10341 ( .A1(n10349), .A2(n9301), .A3(n9319), .ZN(n11090) );
  INV_X1 U10342 ( .A(n16178), .ZN(n16229) );
  XNOR2_X1 U10343 ( .A(n9206), .B(P3_IR_REG_22__SCAN_IN), .ZN(n13040) );
  INV_X1 U10344 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9202) );
  AND2_X1 U10345 ( .A1(n9550), .A2(n9549), .ZN(n9571) );
  NAND2_X1 U10346 ( .A1(n9741), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14218) );
  INV_X1 U10347 ( .A(n14657), .ZN(n14427) );
  NAND2_X1 U10348 ( .A1(n9630), .A2(n14510), .ZN(n14246) );
  AND4_X1 U10349 ( .A1(n13340), .A2(n13339), .A3(n13338), .A4(n13337), .ZN(
        n14180) );
  AND2_X1 U10350 ( .A1(n13258), .A2(n13257), .ZN(n14487) );
  INV_X1 U10351 ( .A(n15817), .ZN(n15830) );
  OR2_X1 U10352 ( .A1(n9566), .A2(n13458), .ZN(n15813) );
  AND2_X1 U10353 ( .A1(n15785), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15838) );
  INV_X1 U10354 ( .A(n7431), .ZN(n14507) );
  AND2_X1 U10355 ( .A1(n9805), .A2(n9660), .ZN(n14520) );
  NOR2_X1 U10356 ( .A1(n16405), .A2(n10204), .ZN(n16401) );
  OR2_X1 U10357 ( .A1(n14520), .A2(n13099), .ZN(n16348) );
  AND2_X1 U10358 ( .A1(n9600), .A2(n11530), .ZN(n9645) );
  OAI21_X1 U10359 ( .B1(n9542), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9341) );
  AND2_X1 U10360 ( .A1(n9496), .A2(n9674), .ZN(n10797) );
  AND2_X1 U10361 ( .A1(n10095), .A2(P2_U3088), .ZN(n11529) );
  INV_X1 U10362 ( .A(n14829), .ZN(n14796) );
  NAND2_X1 U10363 ( .A1(n10169), .A2(n16161), .ZN(n14826) );
  AND4_X1 U10364 ( .A1(n12530), .A2(n12529), .A3(n12528), .A4(n12527), .ZN(
        n12541) );
  INV_X1 U10365 ( .A(n12526), .ZN(n12334) );
  INV_X1 U10366 ( .A(n16022), .ZN(n14900) );
  INV_X1 U10367 ( .A(n16347), .ZN(n16086) );
  AND2_X1 U10368 ( .A1(n16159), .A2(n16194), .ZN(n15090) );
  INV_X1 U10369 ( .A(n16366), .ZN(n16378) );
  INV_X1 U10370 ( .A(n16332), .ZN(n16369) );
  INV_X1 U10371 ( .A(n16190), .ZN(n16383) );
  NAND2_X1 U10372 ( .A1(n10111), .A2(n10110), .ZN(n16194) );
  NOR2_X1 U10373 ( .A1(n12715), .A2(n12752), .ZN(n16332) );
  XNOR2_X1 U10374 ( .A(n9358), .B(P1_IR_REG_23__SCAN_IN), .ZN(n10175) );
  OR2_X1 U10375 ( .A1(n10757), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n10818) );
  AND2_X1 U10376 ( .A1(n9507), .A2(n9490), .ZN(n11363) );
  AND2_X1 U10377 ( .A1(n9960), .A2(n9959), .ZN(n15961) );
  INV_X1 U10378 ( .A(n13568), .ZN(n13604) );
  AND2_X1 U10379 ( .A1(n12995), .A2(n9268), .ZN(n13025) );
  OAI211_X1 U10380 ( .C1(n12992), .C2(n13842), .A(n9123), .B(n9122), .ZN(
        n13611) );
  INV_X1 U10381 ( .A(n11860), .ZN(n13616) );
  INV_X1 U10382 ( .A(n11306), .ZN(n13619) );
  INV_X1 U10383 ( .A(P3_U3897), .ZN(n13623) );
  INV_X1 U10384 ( .A(n15931), .ZN(n15993) );
  NAND2_X1 U10385 ( .A1(n16121), .A2(n16120), .ZN(n13871) );
  INV_X1 U10386 ( .A(n13967), .ZN(n13937) );
  AOI21_X1 U10387 ( .B1(n9310), .B2(n9313), .A(n9312), .ZN(n9314) );
  NAND2_X1 U10388 ( .A1(n16407), .A2(n16200), .ZN(n14030) );
  OR2_X1 U10389 ( .A1(n16415), .A2(n16274), .ZN(n14106) );
  AND2_X2 U10390 ( .A1(n9322), .A2(n9321), .ZN(n16415) );
  NAND2_X1 U10391 ( .A1(n14109), .A2(n9500), .ZN(n9501) );
  AND2_X1 U10392 ( .A1(n10331), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14109) );
  INV_X1 U10393 ( .A(SI_25_), .ZN(n15461) );
  INV_X1 U10394 ( .A(SI_16_), .ZN(n10774) );
  INV_X1 U10395 ( .A(SI_11_), .ZN(n9519) );
  AND2_X1 U10396 ( .A1(n9571), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15800) );
  INV_X1 U10397 ( .A(n14246), .ZN(n12244) );
  NAND2_X1 U10398 ( .A1(n10202), .A2(n9650), .ZN(n14248) );
  INV_X1 U10399 ( .A(n14180), .ZN(n14356) );
  INV_X1 U10400 ( .A(n14345), .ZN(n14344) );
  INV_X1 U10401 ( .A(n13226), .ZN(n14251) );
  AND3_X1 U10402 ( .A1(n15841), .A2(n15840), .A3(n15839), .ZN(n15843) );
  INV_X1 U10403 ( .A(n15838), .ZN(n14306) );
  OR2_X1 U10404 ( .A1(n16405), .A2(n14301), .ZN(n14539) );
  AND3_X1 U10405 ( .A1(n14533), .A2(n14532), .A3(n14531), .ZN(n14623) );
  NAND2_X1 U10406 ( .A1(n16358), .A2(n16170), .ZN(n14631) );
  INV_X1 U10407 ( .A(n16358), .ZN(n16357) );
  OR2_X1 U10410 ( .A1(n15781), .A2(n15779), .ZN(n15780) );
  INV_X1 U10411 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11829) );
  OR2_X1 U10412 ( .A1(n13081), .A2(n10853), .ZN(n14809) );
  INV_X1 U10413 ( .A(n14826), .ZN(n14804) );
  NAND2_X1 U10414 ( .A1(n10166), .A2(n10152), .ZN(n14829) );
  OR2_X1 U10415 ( .A1(n12020), .A2(n12019), .ZN(n14846) );
  OR2_X1 U10416 ( .A1(n9923), .A2(n12781), .ZN(n15852) );
  OR2_X1 U10417 ( .A1(n9923), .A2(n10361), .ZN(n16022) );
  XNOR2_X1 U10418 ( .A(n13057), .B(n13056), .ZN(n15112) );
  INV_X1 U10419 ( .A(n15090), .ZN(n15070) );
  NAND2_X1 U10420 ( .A1(n16086), .A2(n11099), .ZN(n15054) );
  INV_X1 U10421 ( .A(n16387), .ZN(n16385) );
  INV_X1 U10422 ( .A(n16391), .ZN(n16388) );
  AND2_X2 U10423 ( .A1(n10856), .A2(n10855), .ZN(n16391) );
  INV_X1 U10424 ( .A(n9696), .ZN(n9702) );
  INV_X1 U10425 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10825) );
  INV_X1 U10426 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9775) );
  AND2_X1 U10427 ( .A1(n14109), .A2(n9359), .ZN(P3_U3897) );
  INV_X1 U10428 ( .A(n14267), .ZN(P2_U3947) );
  INV_X1 U10429 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n15247) );
  INV_X1 U10430 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9402) );
  NAND2_X1 U10431 ( .A1(n9402), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8725) );
  INV_X1 U10432 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9721) );
  NAND2_X1 U10433 ( .A1(n9721), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8726) );
  INV_X1 U10434 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8727) );
  NAND2_X1 U10435 ( .A1(n8727), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8728) );
  NAND2_X1 U10436 ( .A1(n9399), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8730) );
  NAND2_X1 U10437 ( .A1(n9437), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8732) );
  NAND2_X1 U10438 ( .A1(n9449), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8734) );
  NAND2_X1 U10439 ( .A1(n8940), .A2(n8938), .ZN(n8738) );
  NAND2_X1 U10440 ( .A1(n8736), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8737) );
  XNOR2_X1 U10441 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n8951) );
  NAND2_X1 U10442 ( .A1(n8952), .A2(n8951), .ZN(n8740) );
  NAND2_X1 U10443 ( .A1(n9509), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8739) );
  XNOR2_X1 U10444 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8964) );
  NAND2_X1 U10445 ( .A1(n9518), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8741) );
  XNOR2_X1 U10446 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n8977) );
  NAND2_X1 U10447 ( .A1(n9714), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8742) );
  NAND2_X1 U10448 ( .A1(n8743), .A2(n9775), .ZN(n8744) );
  XNOR2_X1 U10449 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8989) );
  NAND2_X1 U10450 ( .A1(n9877), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8746) );
  XNOR2_X1 U10451 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n9017) );
  NAND2_X1 U10452 ( .A1(n10250), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8747) );
  XNOR2_X1 U10453 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .ZN(n9032) );
  NAND2_X1 U10454 ( .A1(n10525), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8749) );
  NAND2_X1 U10455 ( .A1(n10761), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8751) );
  INV_X1 U10456 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10759) );
  NAND2_X1 U10457 ( .A1(n10759), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8750) );
  NAND2_X1 U10458 ( .A1(n8751), .A2(n8750), .ZN(n9048) );
  NAND2_X1 U10459 ( .A1(n10825), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8752) );
  NAND2_X1 U10460 ( .A1(n10830), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8753) );
  XNOR2_X1 U10461 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .ZN(n9076) );
  INV_X1 U10462 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11009) );
  NAND2_X1 U10463 ( .A1(n11009), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U10464 ( .A1(n8757), .A2(n13096), .ZN(n8758) );
  INV_X1 U10465 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12325) );
  NAND2_X1 U10466 ( .A1(n12325), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8760) );
  INV_X1 U10467 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n13249) );
  NAND2_X1 U10468 ( .A1(n13249), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8759) );
  NAND2_X1 U10469 ( .A1(n8760), .A2(n8759), .ZN(n9102) );
  XNOR2_X1 U10470 ( .A(n13263), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n9116) );
  NAND2_X1 U10471 ( .A1(n13263), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8761) );
  XNOR2_X1 U10472 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n9124) );
  INV_X1 U10473 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n13279) );
  NAND2_X1 U10474 ( .A1(n13279), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8762) );
  NAND2_X1 U10475 ( .A1(n8763), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8764) );
  INV_X1 U10476 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13294) );
  INV_X1 U10477 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n15261) );
  NAND2_X1 U10478 ( .A1(n15261), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8766) );
  INV_X1 U10479 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n14692) );
  NAND2_X1 U10480 ( .A1(n14692), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8765) );
  AND2_X1 U10481 ( .A1(n8766), .A2(n8765), .ZN(n9147) );
  INV_X1 U10482 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15254) );
  NAND2_X1 U10483 ( .A1(n15254), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8768) );
  INV_X1 U10484 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14687) );
  NAND2_X1 U10485 ( .A1(n14687), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8767) );
  AND2_X1 U10486 ( .A1(n8768), .A2(n8767), .ZN(n9161) );
  INV_X1 U10487 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15252) );
  NAND2_X1 U10488 ( .A1(n15252), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8770) );
  INV_X1 U10489 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13333) );
  NAND2_X1 U10490 ( .A1(n13333), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8769) );
  AND2_X1 U10491 ( .A1(n8770), .A2(n8769), .ZN(n9173) );
  INV_X1 U10492 ( .A(n8770), .ZN(n8771) );
  INV_X1 U10493 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13377) );
  AOI22_X1 U10494 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(
        P1_DATAO_REG_28__SCAN_IN), .B1(n13377), .B2(n15247), .ZN(n9189) );
  NOR2_X1 U10495 ( .A1(n9191), .A2(n9189), .ZN(n8772) );
  INV_X1 U10496 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13364) );
  INV_X1 U10497 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n12537) );
  AOI22_X1 U10498 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(
        P1_DATAO_REG_29__SCAN_IN), .B1(n13364), .B2(n12537), .ZN(n12976) );
  INV_X1 U10499 ( .A(n12976), .ZN(n8773) );
  XNOR2_X1 U10500 ( .A(n12977), .B(n8773), .ZN(n14117) );
  NOR2_X1 U10501 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), 
        .ZN(n8785) );
  NAND2_X1 U10502 ( .A1(n14117), .A2(n8822), .ZN(n8798) );
  NAND2_X1 U10503 ( .A1(n9092), .A2(SI_29_), .ZN(n8797) );
  NAND2_X1 U10504 ( .A1(n8798), .A2(n8797), .ZN(n9310) );
  NAND2_X1 U10505 ( .A1(n8862), .A2(n15338), .ZN(n8879) );
  NAND2_X1 U10506 ( .A1(n9008), .A2(n15349), .ZN(n9009) );
  INV_X1 U10507 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n15346) );
  INV_X1 U10508 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n9108) );
  INV_X1 U10509 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9153) );
  NAND2_X1 U10510 ( .A1(n9154), .A2(n9153), .ZN(n9166) );
  INV_X1 U10511 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n9194) );
  NAND2_X1 U10512 ( .A1(n13744), .A2(n9201), .ZN(n12995) );
  INV_X1 U10513 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9311) );
  AND2_X2 U10514 ( .A1(n13465), .A2(n14120), .ZN(n8812) );
  NAND2_X1 U10515 ( .A1(n8812), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8806) );
  NAND2_X1 U10516 ( .A1(n9130), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8805) );
  OAI211_X1 U10517 ( .C1(n9311), .C2(n12988), .A(n8806), .B(n8805), .ZN(n8807)
         );
  INV_X1 U10518 ( .A(n8807), .ZN(n8808) );
  OR2_X1 U10519 ( .A1(n9310), .A2(n12840), .ZN(n13023) );
  NAND2_X1 U10520 ( .A1(n9310), .A2(n12840), .ZN(n13028) );
  NAND2_X1 U10521 ( .A1(n13023), .A2(n13028), .ZN(n12849) );
  NAND2_X1 U10522 ( .A1(n8812), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8810) );
  INV_X1 U10523 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10354) );
  OR2_X1 U10524 ( .A1(n9041), .A2(n10354), .ZN(n8809) );
  XNOR2_X1 U10525 ( .A(n9631), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n8811) );
  MUX2_X1 U10526 ( .A(n8811), .B(SI_0_), .S(n8006), .Z(n14121) );
  MUX2_X1 U10527 ( .A(P3_IR_REG_0__SCAN_IN), .B(n14121), .S(n9949), .Z(n16055)
         );
  NAND2_X1 U10528 ( .A1(n8812), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8818) );
  INV_X1 U10529 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n8813) );
  INV_X1 U10530 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n8814) );
  OR2_X1 U10531 ( .A1(n12992), .A2(n8814), .ZN(n8816) );
  INV_X1 U10532 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n16070) );
  INV_X1 U10533 ( .A(SI_1_), .ZN(n9457) );
  OAI21_X1 U10534 ( .B1(n8821), .B2(n8820), .A(n8819), .ZN(n9455) );
  INV_X1 U10535 ( .A(n9949), .ZN(n8985) );
  NAND2_X1 U10536 ( .A1(n16104), .A2(n8825), .ZN(n12868) );
  NAND2_X1 U10537 ( .A1(n8812), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8831) );
  INV_X1 U10538 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n8826) );
  OR2_X1 U10539 ( .A1(n12988), .A2(n8826), .ZN(n8830) );
  INV_X1 U10540 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n8827) );
  OR2_X1 U10541 ( .A1(n12992), .A2(n8827), .ZN(n8829) );
  INV_X1 U10542 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n16114) );
  OR2_X1 U10543 ( .A1(n9041), .A2(n16114), .ZN(n8828) );
  XNOR2_X1 U10544 ( .A(n8833), .B(n8832), .ZN(n9420) );
  OAI22_X1 U10545 ( .A1(n8873), .A2(n9420), .B1(n10076), .B2(n9949), .ZN(n8836) );
  NOR2_X1 U10546 ( .A1(n8874), .A2(SI_2_), .ZN(n8835) );
  NOR2_X1 U10547 ( .A1(n8836), .A2(n8835), .ZN(n10625) );
  NAND2_X1 U10548 ( .A1(n16052), .A2(n10625), .ZN(n12875) );
  INV_X1 U10549 ( .A(n16052), .ZN(n13622) );
  INV_X1 U10550 ( .A(n10625), .ZN(n16116) );
  NAND2_X1 U10551 ( .A1(n8812), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8841) );
  INV_X1 U10552 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n8837) );
  OR2_X1 U10553 ( .A1(n12988), .A2(n8837), .ZN(n8840) );
  INV_X1 U10554 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11327) );
  OR2_X1 U10555 ( .A1(n12992), .A2(n11327), .ZN(n8839) );
  XNOR2_X1 U10556 ( .A(n8843), .B(n8842), .ZN(n9440) );
  NAND2_X1 U10557 ( .A1(n8844), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8845) );
  XNOR2_X1 U10558 ( .A(n8845), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10289) );
  OAI22_X1 U10559 ( .A1(n8873), .A2(n9440), .B1(n10289), .B2(n9949), .ZN(n8847) );
  NOR2_X1 U10560 ( .A1(n8874), .A2(SI_3_), .ZN(n8846) );
  NAND2_X1 U10561 ( .A1(n16102), .A2(n11329), .ZN(n12877) );
  INV_X1 U10562 ( .A(n16102), .ZN(n13621) );
  INV_X1 U10563 ( .A(n11329), .ZN(n8848) );
  NAND2_X1 U10564 ( .A1(n8812), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8853) );
  AND2_X1 U10565 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8849) );
  NOR2_X1 U10566 ( .A1(n8862), .A2(n8849), .ZN(n11039) );
  OR2_X1 U10567 ( .A1(n9041), .A2(n11039), .ZN(n8852) );
  NAND2_X1 U10568 ( .A1(n9263), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8851) );
  NAND2_X1 U10569 ( .A1(n9130), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8850) );
  XNOR2_X1 U10570 ( .A(n8855), .B(n8854), .ZN(n9474) );
  INV_X1 U10571 ( .A(SI_4_), .ZN(n15495) );
  NAND2_X1 U10572 ( .A1(n9092), .A2(n15495), .ZN(n8858) );
  INV_X1 U10573 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8856) );
  NAND2_X1 U10574 ( .A1(n8985), .A2(n10485), .ZN(n8857) );
  XNOR2_X1 U10575 ( .A(n13620), .B(n12881), .ZN(n13004) );
  INV_X1 U10576 ( .A(n13004), .ZN(n11218) );
  NAND2_X1 U10577 ( .A1(n11215), .A2(n11218), .ZN(n8860) );
  INV_X1 U10578 ( .A(n12881), .ZN(n16182) );
  NAND2_X1 U10579 ( .A1(n11209), .A2(n16182), .ZN(n8859) );
  NAND2_X1 U10580 ( .A1(n8812), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8868) );
  INV_X1 U10581 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n8861) );
  OR2_X1 U10582 ( .A1(n12988), .A2(n8861), .ZN(n8867) );
  OR2_X1 U10583 ( .A1(n8862), .A2(n15338), .ZN(n8863) );
  AND2_X1 U10584 ( .A1(n8879), .A2(n8863), .ZN(n11419) );
  OR2_X1 U10585 ( .A1(n9041), .A2(n11419), .ZN(n8866) );
  INV_X1 U10586 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n8864) );
  OR2_X1 U10587 ( .A1(n12992), .A2(n8864), .ZN(n8865) );
  XNOR2_X1 U10588 ( .A(n8870), .B(n8869), .ZN(n9442) );
  OR2_X1 U10589 ( .A1(n8871), .A2(n14112), .ZN(n8872) );
  OAI22_X1 U10590 ( .A1(n8873), .A2(n9442), .B1(n10497), .B2(n9949), .ZN(n8876) );
  NOR2_X1 U10591 ( .A1(n8874), .A2(SI_5_), .ZN(n8875) );
  INV_X1 U10592 ( .A(n16199), .ZN(n11420) );
  NAND2_X1 U10593 ( .A1(n13619), .A2(n11420), .ZN(n12887) );
  NAND2_X1 U10594 ( .A1(n11306), .A2(n16199), .ZN(n12886) );
  NAND2_X1 U10595 ( .A1(n11418), .A2(n12997), .ZN(n8877) );
  INV_X1 U10596 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n8878) );
  OR2_X1 U10597 ( .A1(n12988), .A2(n8878), .ZN(n8885) );
  NAND2_X1 U10598 ( .A1(n8879), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8880) );
  AND2_X1 U10599 ( .A1(n8894), .A2(n8880), .ZN(n11534) );
  OR2_X1 U10600 ( .A1(n9041), .A2(n11534), .ZN(n8884) );
  INV_X1 U10601 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n8881) );
  OR2_X1 U10602 ( .A1(n12992), .A2(n8881), .ZN(n8883) );
  NAND2_X1 U10603 ( .A1(n8812), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8882) );
  NAND2_X1 U10604 ( .A1(n9092), .A2(SI_6_), .ZN(n8893) );
  XNOR2_X1 U10605 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n8886) );
  XNOR2_X1 U10606 ( .A(n8887), .B(n8886), .ZN(n9458) );
  NAND2_X1 U10607 ( .A1(n8822), .A2(n9458), .ZN(n8892) );
  NAND2_X1 U10608 ( .A1(n8871), .A2(n8888), .ZN(n8903) );
  NAND2_X1 U10609 ( .A1(n8903), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8890) );
  XNOR2_X1 U10610 ( .A(n8890), .B(n8889), .ZN(n10573) );
  INV_X1 U10611 ( .A(n10573), .ZN(n10514) );
  NAND2_X1 U10612 ( .A1(n8985), .A2(n10514), .ZN(n8891) );
  INV_X1 U10613 ( .A(n13618), .ZN(n11626) );
  INV_X1 U10614 ( .A(n16215), .ZN(n11309) );
  NAND2_X1 U10615 ( .A1(n11626), .A2(n11309), .ZN(n12891) );
  AND2_X1 U10616 ( .A1(n8894), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8895) );
  NOR2_X1 U10617 ( .A1(n8910), .A2(n8895), .ZN(n11631) );
  OR2_X1 U10618 ( .A1(n9086), .A2(n11631), .ZN(n8900) );
  INV_X1 U10619 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n8896) );
  OR2_X1 U10620 ( .A1(n12992), .A2(n8896), .ZN(n8899) );
  NAND2_X1 U10621 ( .A1(n8812), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8898) );
  NAND2_X1 U10622 ( .A1(n9263), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8897) );
  NAND4_X1 U10623 ( .A1(n8900), .A2(n8899), .A3(n8898), .A4(n8897), .ZN(n13617) );
  XNOR2_X1 U10624 ( .A(n8902), .B(n8901), .ZN(n9461) );
  NAND2_X1 U10625 ( .A1(n8822), .A2(n9461), .ZN(n8906) );
  NAND2_X1 U10626 ( .A1(n8920), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8904) );
  XNOR2_X1 U10627 ( .A(n8904), .B(P3_IR_REG_7__SCAN_IN), .ZN(n10708) );
  INV_X1 U10628 ( .A(n10708), .ZN(n10562) );
  NAND2_X1 U10629 ( .A1(n8985), .A2(n10562), .ZN(n8905) );
  OAI211_X1 U10630 ( .C1(SI_7_), .C2(n9080), .A(n8906), .B(n8905), .ZN(n16231)
         );
  XNOR2_X1 U10631 ( .A(n13617), .B(n16231), .ZN(n13005) );
  INV_X1 U10632 ( .A(n13005), .ZN(n12894) );
  INV_X1 U10633 ( .A(n13617), .ZN(n11670) );
  INV_X1 U10634 ( .A(n16231), .ZN(n12895) );
  NAND2_X1 U10635 ( .A1(n11670), .A2(n12895), .ZN(n8907) );
  NAND2_X1 U10636 ( .A1(n8908), .A2(n8907), .ZN(n11669) );
  NAND2_X1 U10637 ( .A1(n8812), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8917) );
  INV_X1 U10638 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n8909) );
  OR2_X1 U10639 ( .A1(n12988), .A2(n8909), .ZN(n8916) );
  NOR2_X1 U10640 ( .A1(n8910), .A2(n10705), .ZN(n8911) );
  OR2_X1 U10641 ( .A1(n8927), .A2(n8911), .ZN(n11677) );
  INV_X1 U10642 ( .A(n11677), .ZN(n8912) );
  OR2_X1 U10643 ( .A1(n9086), .A2(n8912), .ZN(n8915) );
  INV_X1 U10644 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n8913) );
  OR2_X1 U10645 ( .A1(n12992), .A2(n8913), .ZN(n8914) );
  XNOR2_X1 U10646 ( .A(n8919), .B(n8918), .ZN(n9473) );
  NAND2_X1 U10647 ( .A1(n9092), .A2(SI_8_), .ZN(n8926) );
  NOR2_X1 U10648 ( .A1(n8920), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8923) );
  OR2_X1 U10649 ( .A1(n8923), .A2(n14112), .ZN(n8921) );
  MUX2_X1 U10650 ( .A(n8921), .B(P3_IR_REG_31__SCAN_IN), .S(n8922), .Z(n8924)
         );
  NAND2_X1 U10651 ( .A1(n8923), .A2(n8922), .ZN(n8933) );
  INV_X1 U10652 ( .A(n10958), .ZN(n10717) );
  NAND2_X1 U10653 ( .A1(n8985), .A2(n10717), .ZN(n8925) );
  OAI211_X1 U10654 ( .C1(n8873), .C2(n9473), .A(n8926), .B(n8925), .ZN(n11678)
         );
  NAND2_X1 U10655 ( .A1(n11860), .A2(n11678), .ZN(n12901) );
  INV_X1 U10656 ( .A(n11678), .ZN(n16257) );
  NAND2_X1 U10657 ( .A1(n13616), .A2(n16257), .ZN(n12902) );
  NAND2_X1 U10658 ( .A1(n8812), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8932) );
  OR2_X1 U10659 ( .A1(n8927), .A2(n15536), .ZN(n8928) );
  AND2_X1 U10660 ( .A1(n8944), .A2(n8928), .ZN(n11864) );
  OR2_X1 U10661 ( .A1(n9086), .A2(n11864), .ZN(n8931) );
  NAND2_X1 U10662 ( .A1(n9263), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8930) );
  NAND2_X1 U10663 ( .A1(n9130), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8929) );
  NAND4_X1 U10664 ( .A1(n8932), .A2(n8931), .A3(n8930), .A4(n8929), .ZN(n13615) );
  NAND2_X1 U10665 ( .A1(n8933), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8934) );
  MUX2_X1 U10666 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8934), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n8937) );
  INV_X1 U10667 ( .A(n8935), .ZN(n8936) );
  NAND2_X1 U10668 ( .A1(n8937), .A2(n8936), .ZN(n10959) );
  OAI22_X1 U10669 ( .A1(n9080), .A2(SI_9_), .B1(n11121), .B2(n9949), .ZN(n8942) );
  INV_X1 U10670 ( .A(n8938), .ZN(n8939) );
  XNOR2_X1 U10671 ( .A(n8940), .B(n8939), .ZN(n9438) );
  NOR2_X1 U10672 ( .A1(n8873), .A2(n9438), .ZN(n8941) );
  NOR2_X1 U10673 ( .A1(n8942), .A2(n8941), .ZN(n11863) );
  INV_X1 U10674 ( .A(n11863), .ZN(n16273) );
  NOR2_X1 U10675 ( .A1(n13615), .A2(n16273), .ZN(n12905) );
  NAND2_X1 U10676 ( .A1(n13615), .A2(n16273), .ZN(n12907) );
  INV_X1 U10677 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n8943) );
  OR2_X1 U10678 ( .A1(n12988), .A2(n8943), .ZN(n8950) );
  NAND2_X1 U10679 ( .A1(n8944), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8945) );
  AND2_X1 U10680 ( .A1(n8958), .A2(n8945), .ZN(n12035) );
  OR2_X1 U10681 ( .A1(n9041), .A2(n12035), .ZN(n8949) );
  INV_X1 U10682 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n8946) );
  OR2_X1 U10683 ( .A1(n12992), .A2(n8946), .ZN(n8948) );
  NAND2_X1 U10684 ( .A1(n8812), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8947) );
  NAND4_X1 U10685 ( .A1(n8950), .A2(n8949), .A3(n8948), .A4(n8947), .ZN(n13614) );
  XNOR2_X1 U10686 ( .A(n8952), .B(n8951), .ZN(n16289) );
  NAND2_X1 U10687 ( .A1(n8822), .A2(n16289), .ZN(n8955) );
  OR2_X1 U10688 ( .A1(n8935), .A2(n14112), .ZN(n8953) );
  XNOR2_X1 U10689 ( .A(n8953), .B(n8966), .ZN(n16294) );
  NAND2_X1 U10690 ( .A1(n8985), .A2(n16294), .ZN(n8954) );
  OAI211_X1 U10691 ( .C1(SI_10_), .C2(n9080), .A(n8955), .B(n8954), .ZN(n16295) );
  XNOR2_X1 U10692 ( .A(n13614), .B(n16295), .ZN(n13011) );
  INV_X1 U10693 ( .A(n13614), .ZN(n12910) );
  INV_X1 U10694 ( .A(n16295), .ZN(n9238) );
  NAND2_X1 U10695 ( .A1(n12910), .A2(n9238), .ZN(n8957) );
  NAND2_X1 U10696 ( .A1(n8812), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8963) );
  NAND2_X1 U10697 ( .A1(n8958), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8959) );
  AND2_X1 U10698 ( .A1(n8971), .A2(n8959), .ZN(n12103) );
  OR2_X1 U10699 ( .A1(n9086), .A2(n12103), .ZN(n8962) );
  NAND2_X1 U10700 ( .A1(n9263), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8961) );
  NAND2_X1 U10701 ( .A1(n9130), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8960) );
  NAND4_X1 U10702 ( .A1(n8963), .A2(n8962), .A3(n8961), .A4(n8960), .ZN(n13613) );
  XNOR2_X1 U10703 ( .A(n8965), .B(n8964), .ZN(n9470) );
  NAND2_X1 U10704 ( .A1(n8822), .A2(n9470), .ZN(n8969) );
  NAND2_X1 U10705 ( .A1(n8935), .A2(n8966), .ZN(n8979) );
  NAND2_X1 U10706 ( .A1(n8979), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8967) );
  XNOR2_X1 U10707 ( .A(n8967), .B(P3_IR_REG_11__SCAN_IN), .ZN(n13655) );
  INV_X1 U10708 ( .A(n13655), .ZN(n11466) );
  NAND2_X1 U10709 ( .A1(n8985), .A2(n11466), .ZN(n8968) );
  OAI211_X1 U10710 ( .C1(SI_11_), .C2(n9080), .A(n8969), .B(n8968), .ZN(n16312) );
  INV_X1 U10711 ( .A(n16312), .ZN(n8970) );
  NAND2_X1 U10712 ( .A1(n8384), .A2(n8970), .ZN(n12917) );
  NAND2_X1 U10713 ( .A1(n13613), .A2(n16312), .ZN(n12916) );
  NAND2_X1 U10714 ( .A1(n11994), .A2(n13008), .ZN(n11993) );
  NAND2_X1 U10715 ( .A1(n11993), .A2(n12917), .ZN(n12108) );
  NAND2_X1 U10716 ( .A1(n9263), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8976) );
  AND2_X1 U10717 ( .A1(n8971), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8972) );
  NOR2_X1 U10718 ( .A1(n9008), .A2(n8972), .ZN(n12165) );
  OR2_X1 U10719 ( .A1(n9041), .A2(n12165), .ZN(n8975) );
  NAND2_X1 U10720 ( .A1(n9130), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8974) );
  NAND2_X1 U10721 ( .A1(n8812), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8973) );
  NAND4_X1 U10722 ( .A1(n8976), .A2(n8975), .A3(n8974), .A4(n8973), .ZN(n13612) );
  XNOR2_X1 U10723 ( .A(n8978), .B(n8977), .ZN(n9471) );
  NAND2_X1 U10724 ( .A1(n8822), .A2(n9471), .ZN(n8988) );
  NAND2_X1 U10725 ( .A1(n9092), .A2(n15485), .ZN(n8987) );
  INV_X1 U10726 ( .A(n9002), .ZN(n8984) );
  NAND2_X1 U10727 ( .A1(n8980), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8982) );
  MUX2_X1 U10728 ( .A(n8982), .B(P3_IR_REG_31__SCAN_IN), .S(n8981), .Z(n8983)
         );
  NAND2_X1 U10729 ( .A1(n8984), .A2(n8983), .ZN(n15926) );
  NAND2_X1 U10730 ( .A1(n8985), .A2(n15926), .ZN(n8986) );
  NAND2_X1 U10731 ( .A1(n13959), .A2(n12156), .ZN(n12920) );
  NAND2_X1 U10732 ( .A1(n13612), .A2(n14031), .ZN(n12921) );
  XNOR2_X1 U10733 ( .A(n8990), .B(n8989), .ZN(n9499) );
  NAND2_X1 U10734 ( .A1(n9499), .A2(n8822), .ZN(n8995) );
  INV_X1 U10735 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9003) );
  NAND2_X1 U10736 ( .A1(n9002), .A2(n9003), .ZN(n9019) );
  NAND2_X1 U10737 ( .A1(n9019), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8992) );
  INV_X1 U10738 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8991) );
  XNOR2_X1 U10739 ( .A(n8992), .B(n8991), .ZN(n15958) );
  INV_X1 U10740 ( .A(n15958), .ZN(n13634) );
  OAI22_X1 U10741 ( .A1(n9080), .A2(SI_14_), .B1(n13634), .B2(n9949), .ZN(
        n8993) );
  INV_X1 U10742 ( .A(n8993), .ZN(n8994) );
  NAND2_X1 U10743 ( .A1(n9009), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8996) );
  AND2_X1 U10744 ( .A1(n9025), .A2(n8996), .ZN(n13950) );
  OR2_X1 U10745 ( .A1(n9086), .A2(n13950), .ZN(n9000) );
  INV_X1 U10746 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13951) );
  OR2_X1 U10747 ( .A1(n12992), .A2(n13951), .ZN(n8999) );
  NAND2_X1 U10748 ( .A1(n8812), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8998) );
  NAND2_X1 U10749 ( .A1(n9263), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8997) );
  NAND4_X1 U10750 ( .A1(n9000), .A2(n8999), .A3(n8998), .A4(n8997), .ZN(n13927) );
  OR2_X1 U10751 ( .A1(n14097), .A2(n13927), .ZN(n12925) );
  NAND2_X1 U10752 ( .A1(n14097), .A2(n13927), .ZN(n9015) );
  INV_X1 U10753 ( .A(n13948), .ZN(n13939) );
  XNOR2_X1 U10754 ( .A(n9001), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n9481) );
  NAND2_X1 U10755 ( .A1(n9481), .A2(n8822), .ZN(n9007) );
  OR2_X1 U10756 ( .A1(n9002), .A2(n14112), .ZN(n9004) );
  XNOR2_X1 U10757 ( .A(n9004), .B(n9003), .ZN(n15944) );
  INV_X1 U10758 ( .A(n15944), .ZN(n13659) );
  OAI22_X1 U10759 ( .A1(n9080), .A2(SI_13_), .B1(n13659), .B2(n9949), .ZN(
        n9005) );
  INV_X1 U10760 ( .A(n9005), .ZN(n9006) );
  NAND2_X1 U10761 ( .A1(n8812), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9014) );
  OR2_X1 U10762 ( .A1(n9008), .A2(n15349), .ZN(n9010) );
  AND2_X1 U10763 ( .A1(n9010), .A2(n9009), .ZN(n13964) );
  OR2_X1 U10764 ( .A1(n9041), .A2(n13964), .ZN(n9013) );
  NAND2_X1 U10765 ( .A1(n9263), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n9012) );
  NAND2_X1 U10766 ( .A1(n9130), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n9011) );
  NAND4_X1 U10767 ( .A1(n9014), .A2(n9013), .A3(n9012), .A4(n9011), .ZN(n13942) );
  AND2_X1 U10768 ( .A1(n14101), .A2(n13942), .ZN(n13947) );
  NOR2_X1 U10769 ( .A1(n13939), .A2(n13947), .ZN(n12927) );
  NOR2_X1 U10770 ( .A1(n14101), .A2(n13942), .ZN(n12793) );
  NAND2_X1 U10771 ( .A1(n9015), .A2(n12793), .ZN(n9016) );
  XNOR2_X1 U10772 ( .A(n9018), .B(n9017), .ZN(n9502) );
  NAND2_X1 U10773 ( .A1(n9502), .A2(n8822), .ZN(n9024) );
  OAI21_X1 U10774 ( .B1(n9019), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9021) );
  INV_X1 U10775 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n9020) );
  XNOR2_X1 U10776 ( .A(n9021), .B(n9020), .ZN(n15983) );
  OAI22_X1 U10777 ( .A1(n9080), .A2(SI_15_), .B1(n13662), .B2(n9949), .ZN(
        n9022) );
  INV_X1 U10778 ( .A(n9022), .ZN(n9023) );
  NAND2_X1 U10779 ( .A1(n9024), .A2(n9023), .ZN(n14017) );
  INV_X1 U10780 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n15987) );
  OR2_X1 U10781 ( .A1(n12988), .A2(n15987), .ZN(n9030) );
  AND2_X1 U10782 ( .A1(n9025), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9026) );
  NOR2_X1 U10783 ( .A1(n9039), .A2(n9026), .ZN(n13931) );
  OR2_X1 U10784 ( .A1(n9086), .A2(n13931), .ZN(n9029) );
  INV_X1 U10785 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n15980) );
  OR2_X1 U10786 ( .A1(n12992), .A2(n15980), .ZN(n9028) );
  NAND2_X1 U10787 ( .A1(n8812), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9027) );
  NAND4_X1 U10788 ( .A1(n9030), .A2(n9029), .A3(n9028), .A4(n9027), .ZN(n13944) );
  OR2_X1 U10789 ( .A1(n14017), .A2(n13944), .ZN(n12932) );
  NAND2_X1 U10790 ( .A1(n14017), .A2(n13944), .ZN(n12933) );
  NAND2_X1 U10791 ( .A1(n13921), .A2(n13922), .ZN(n9031) );
  XNOR2_X1 U10792 ( .A(n9033), .B(n7697), .ZN(n9703) );
  NAND2_X1 U10793 ( .A1(n9703), .A2(n8822), .ZN(n9038) );
  NAND2_X1 U10794 ( .A1(n9034), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9035) );
  OAI22_X1 U10795 ( .A1(n9080), .A2(n10774), .B1(n9949), .B2(n13676), .ZN(
        n9036) );
  INV_X1 U10796 ( .A(n9036), .ZN(n9037) );
  NAND2_X1 U10797 ( .A1(n8812), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9045) );
  INV_X1 U10798 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13646) );
  OR2_X1 U10799 ( .A1(n12988), .A2(n13646), .ZN(n9044) );
  NOR2_X1 U10800 ( .A1(n9039), .A2(n13518), .ZN(n9040) );
  OR2_X1 U10801 ( .A1(n9086), .A2(n8715), .ZN(n9043) );
  INV_X1 U10802 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13916) );
  OR2_X1 U10803 ( .A1(n12992), .A2(n13916), .ZN(n9042) );
  XNOR2_X1 U10804 ( .A(n13918), .B(n13899), .ZN(n13910) );
  NAND2_X1 U10805 ( .A1(n13909), .A2(n7729), .ZN(n9047) );
  NAND2_X1 U10806 ( .A1(n13918), .A2(n13899), .ZN(n9046) );
  INV_X1 U10807 ( .A(n9048), .ZN(n9049) );
  XNOR2_X1 U10808 ( .A(n9050), .B(n9049), .ZN(n9692) );
  NAND2_X1 U10809 ( .A1(n9692), .A2(n8822), .ZN(n9056) );
  INV_X1 U10810 ( .A(n9051), .ZN(n9052) );
  NAND2_X1 U10811 ( .A1(n9052), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9053) );
  XNOR2_X1 U10812 ( .A(n9053), .B(P3_IR_REG_17__SCAN_IN), .ZN(n13706) );
  OAI22_X1 U10813 ( .A1(n9080), .A2(SI_17_), .B1(n13706), .B2(n9949), .ZN(
        n9054) );
  INV_X1 U10814 ( .A(n9054), .ZN(n9055) );
  NAND2_X1 U10815 ( .A1(n8812), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n9062) );
  INV_X1 U10816 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n14011) );
  OR2_X1 U10817 ( .A1(n12988), .A2(n14011), .ZN(n9061) );
  OR2_X1 U10818 ( .A1(n9057), .A2(n15531), .ZN(n9058) );
  AND2_X1 U10819 ( .A1(n9071), .A2(n9058), .ZN(n13903) );
  OR2_X1 U10820 ( .A1(n9086), .A2(n13903), .ZN(n9060) );
  INV_X1 U10821 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13904) );
  OR2_X1 U10822 ( .A1(n12992), .A2(n13904), .ZN(n9059) );
  XNOR2_X1 U10823 ( .A(n14089), .B(n12807), .ZN(n13901) );
  NAND2_X1 U10824 ( .A1(n13902), .A2(n13901), .ZN(n9063) );
  OR2_X1 U10825 ( .A1(n14089), .A2(n13913), .ZN(n12940) );
  NAND2_X1 U10826 ( .A1(n9063), .A2(n12940), .ZN(n13894) );
  AOI22_X1 U10827 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n10830), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n10825), .ZN(n9064) );
  XNOR2_X1 U10828 ( .A(n9065), .B(n9064), .ZN(n9814) );
  NAND2_X1 U10829 ( .A1(n9814), .A2(n8822), .ZN(n9070) );
  NAND2_X1 U10830 ( .A1(n9066), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9067) );
  XNOR2_X1 U10831 ( .A(n9067), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13721) );
  OAI22_X1 U10832 ( .A1(n9080), .A2(n11001), .B1(n9949), .B2(n13719), .ZN(
        n9068) );
  INV_X1 U10833 ( .A(n9068), .ZN(n9069) );
  NAND2_X1 U10834 ( .A1(n8812), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n9075) );
  INV_X1 U10835 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13709) );
  OR2_X1 U10836 ( .A1(n12988), .A2(n13709), .ZN(n9074) );
  INV_X1 U10837 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n15549) );
  XNOR2_X1 U10838 ( .A(n9071), .B(n15549), .ZN(n13889) );
  OR2_X1 U10839 ( .A1(n9086), .A2(n13889), .ZN(n9073) );
  INV_X1 U10840 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13890) );
  OR2_X1 U10841 ( .A1(n12992), .A2(n13890), .ZN(n9072) );
  OR2_X1 U10842 ( .A1(n14005), .A2(n13900), .ZN(n12939) );
  NAND2_X1 U10843 ( .A1(n14005), .A2(n13900), .ZN(n12942) );
  NAND2_X1 U10844 ( .A1(n12939), .A2(n12942), .ZN(n13885) );
  INV_X1 U10845 ( .A(n13885), .ZN(n13893) );
  XNOR2_X1 U10846 ( .A(n9077), .B(n9076), .ZN(n9883) );
  NAND2_X1 U10847 ( .A1(n9883), .A2(n8822), .ZN(n9083) );
  INV_X1 U10848 ( .A(n9203), .ZN(n9078) );
  NAND2_X1 U10849 ( .A1(n9078), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9079) );
  OAI22_X1 U10850 ( .A1(n9080), .A2(n15473), .B1(n13733), .B2(n9949), .ZN(
        n9081) );
  INV_X1 U10851 ( .A(n9081), .ZN(n9082) );
  AND2_X1 U10852 ( .A1(n9084), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9085) );
  NOR2_X1 U10853 ( .A1(n9095), .A2(n9085), .ZN(n13879) );
  OR2_X1 U10854 ( .A1(n9086), .A2(n13879), .ZN(n9090) );
  INV_X1 U10855 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13880) );
  OR2_X1 U10856 ( .A1(n12992), .A2(n13880), .ZN(n9089) );
  NAND2_X1 U10857 ( .A1(n9263), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n9088) );
  NAND2_X1 U10858 ( .A1(n8812), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9087) );
  NAND4_X1 U10859 ( .A1(n9090), .A2(n9089), .A3(n9088), .A4(n9087), .ZN(n13887) );
  OR2_X1 U10860 ( .A1(n14001), .A2(n13574), .ZN(n12946) );
  NAND2_X1 U10861 ( .A1(n14001), .A2(n13574), .ZN(n12947) );
  XNOR2_X1 U10862 ( .A(n9091), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n10312) );
  NAND2_X1 U10863 ( .A1(n10312), .A2(n8822), .ZN(n9094) );
  NAND2_X1 U10864 ( .A1(n9092), .A2(SI_20_), .ZN(n9093) );
  NOR2_X1 U10865 ( .A1(n9095), .A2(n15346), .ZN(n9096) );
  OR2_X1 U10866 ( .A1(n9109), .A2(n9096), .ZN(n13867) );
  NAND2_X1 U10867 ( .A1(n13867), .A2(n9201), .ZN(n9101) );
  NAND2_X1 U10868 ( .A1(n9263), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n9100) );
  INV_X1 U10869 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n13866) );
  OR2_X1 U10870 ( .A1(n12992), .A2(n13866), .ZN(n9099) );
  INV_X1 U10871 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n14079) );
  OR2_X1 U10872 ( .A1(n9097), .A2(n14079), .ZN(n9098) );
  OR2_X1 U10873 ( .A1(n14080), .A2(n13847), .ZN(n12951) );
  NAND2_X1 U10874 ( .A1(n14080), .A2(n13847), .ZN(n12952) );
  NAND2_X1 U10875 ( .A1(n12951), .A2(n12952), .ZN(n13858) );
  INV_X1 U10876 ( .A(n13858), .ZN(n13860) );
  NAND2_X1 U10877 ( .A1(n9103), .A2(n9102), .ZN(n9104) );
  NAND2_X1 U10878 ( .A1(n9105), .A2(n9104), .ZN(n10356) );
  OR2_X1 U10879 ( .A1(n10356), .A2(n8873), .ZN(n9107) );
  NAND2_X1 U10880 ( .A1(n9092), .A2(SI_21_), .ZN(n9106) );
  OR2_X1 U10881 ( .A1(n9109), .A2(n9108), .ZN(n9110) );
  NAND2_X1 U10882 ( .A1(n9120), .A2(n9110), .ZN(n13855) );
  NAND2_X1 U10883 ( .A1(n13855), .A2(n9201), .ZN(n9114) );
  NAND2_X1 U10884 ( .A1(n9263), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n9113) );
  NAND2_X1 U10885 ( .A1(n9130), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n9112) );
  NAND2_X1 U10886 ( .A1(n8812), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n9111) );
  NAND4_X1 U10887 ( .A1(n9114), .A2(n9113), .A3(n9112), .A4(n9111), .ZN(n13862) );
  OR2_X1 U10888 ( .A1(n14074), .A2(n13837), .ZN(n12955) );
  NAND2_X1 U10889 ( .A1(n14074), .A2(n13837), .ZN(n12956) );
  NAND2_X1 U10890 ( .A1(n13846), .A2(n13850), .ZN(n9115) );
  XNOR2_X1 U10891 ( .A(n9117), .B(n9116), .ZN(n10532) );
  NAND2_X1 U10892 ( .A1(n10532), .A2(n8822), .ZN(n9119) );
  NAND2_X1 U10893 ( .A1(n9092), .A2(SI_22_), .ZN(n9118) );
  INV_X1 U10894 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n13842) );
  NAND2_X1 U10895 ( .A1(n9120), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9121) );
  NAND2_X1 U10896 ( .A1(n9128), .A2(n9121), .ZN(n13843) );
  NAND2_X1 U10897 ( .A1(n13843), .A2(n9201), .ZN(n9123) );
  AOI22_X1 U10898 ( .A1(n8812), .A2(P3_REG0_REG_22__SCAN_IN), .B1(n9263), .B2(
        P3_REG1_REG_22__SCAN_IN), .ZN(n9122) );
  XNOR2_X1 U10899 ( .A(n9125), .B(n9124), .ZN(n10850) );
  NAND2_X1 U10900 ( .A1(n10850), .A2(n8822), .ZN(n9127) );
  NAND2_X1 U10901 ( .A1(n9092), .A2(SI_23_), .ZN(n9126) );
  NAND2_X1 U10902 ( .A1(n9128), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9129) );
  NAND2_X1 U10903 ( .A1(n9139), .A2(n9129), .ZN(n13827) );
  NAND2_X1 U10904 ( .A1(n13827), .A2(n9201), .ZN(n9133) );
  AOI22_X1 U10905 ( .A1(n9130), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n9263), .B2(
        P3_REG1_REG_23__SCAN_IN), .ZN(n9132) );
  NAND2_X1 U10906 ( .A1(n8812), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n9131) );
  NAND2_X1 U10907 ( .A1(n13482), .A2(n13838), .ZN(n12862) );
  INV_X1 U10908 ( .A(n13825), .ZN(n9134) );
  XNOR2_X1 U10909 ( .A(n9136), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n11291) );
  NAND2_X1 U10910 ( .A1(n11291), .A2(n8822), .ZN(n9138) );
  NAND2_X1 U10911 ( .A1(n9092), .A2(SI_24_), .ZN(n9137) );
  INV_X1 U10912 ( .A(n9154), .ZN(n9141) );
  NAND2_X1 U10913 ( .A1(n9139), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9140) );
  NAND2_X1 U10914 ( .A1(n9141), .A2(n9140), .ZN(n13820) );
  NAND2_X1 U10915 ( .A1(n13820), .A2(n9201), .ZN(n9146) );
  INV_X1 U10916 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n13819) );
  NAND2_X1 U10917 ( .A1(n8812), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n9143) );
  NAND2_X1 U10918 ( .A1(n9263), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9142) );
  OAI211_X1 U10919 ( .C1(n13819), .C2(n12992), .A(n9143), .B(n9142), .ZN(n9144) );
  INV_X1 U10920 ( .A(n9144), .ZN(n9145) );
  NAND2_X1 U10921 ( .A1(n14058), .A2(n8379), .ZN(n12859) );
  NAND2_X1 U10922 ( .A1(n9150), .A2(n9149), .ZN(n11392) );
  NAND2_X1 U10923 ( .A1(n9092), .A2(SI_25_), .ZN(n9151) );
  OR2_X1 U10924 ( .A1(n9154), .A2(n9153), .ZN(n9155) );
  NAND2_X1 U10925 ( .A1(n9166), .A2(n9155), .ZN(n13808) );
  INV_X1 U10926 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n9158) );
  NAND2_X1 U10927 ( .A1(n8812), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n9157) );
  NAND2_X1 U10928 ( .A1(n9263), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9156) );
  OAI211_X1 U10929 ( .C1(n9158), .C2(n12992), .A(n9157), .B(n9156), .ZN(n9159)
         );
  INV_X1 U10930 ( .A(n9258), .ZN(n9160) );
  OR2_X1 U10931 ( .A1(n9162), .A2(n9161), .ZN(n9163) );
  NAND2_X1 U10932 ( .A1(n9092), .A2(SI_26_), .ZN(n9165) );
  NAND2_X1 U10933 ( .A1(n9166), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9167) );
  NAND2_X1 U10934 ( .A1(n9178), .A2(n9167), .ZN(n13792) );
  NAND2_X1 U10935 ( .A1(n13792), .A2(n9201), .ZN(n9172) );
  INV_X1 U10936 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n13791) );
  NAND2_X1 U10937 ( .A1(n9263), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9169) );
  NAND2_X1 U10938 ( .A1(n8812), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n9168) );
  OAI211_X1 U10939 ( .C1(n12992), .C2(n13791), .A(n9169), .B(n9168), .ZN(n9170) );
  INV_X1 U10940 ( .A(n9170), .ZN(n9171) );
  INV_X1 U10941 ( .A(n9173), .ZN(n9174) );
  NAND2_X1 U10942 ( .A1(n11869), .A2(n8822), .ZN(n9177) );
  NAND2_X1 U10943 ( .A1(n9092), .A2(SI_27_), .ZN(n9176) );
  INV_X1 U10944 ( .A(n9195), .ZN(n9180) );
  NAND2_X1 U10945 ( .A1(n9178), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9179) );
  NAND2_X1 U10946 ( .A1(n9180), .A2(n9179), .ZN(n13781) );
  NAND2_X1 U10947 ( .A1(n13781), .A2(n9201), .ZN(n9185) );
  INV_X1 U10948 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n13780) );
  NAND2_X1 U10949 ( .A1(n9263), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9182) );
  NAND2_X1 U10950 ( .A1(n8812), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n9181) );
  OAI211_X1 U10951 ( .C1(n13780), .C2(n12992), .A(n9182), .B(n9181), .ZN(n9183) );
  INV_X1 U10952 ( .A(n9183), .ZN(n9184) );
  NAND2_X2 U10953 ( .A1(n9185), .A2(n9184), .ZN(n13787) );
  INV_X1 U10954 ( .A(n13787), .ZN(n12842) );
  NAND2_X1 U10955 ( .A1(n8258), .A2(n9257), .ZN(n9186) );
  OAI211_X1 U10956 ( .C1(n14042), .C2(n12842), .A(n9186), .B(n12850), .ZN(
        n9188) );
  NAND2_X1 U10957 ( .A1(n14042), .A2(n12842), .ZN(n9187) );
  NAND2_X1 U10958 ( .A1(n13768), .A2(n12855), .ZN(n13758) );
  INV_X1 U10959 ( .A(n9189), .ZN(n9190) );
  XNOR2_X1 U10960 ( .A(n9191), .B(n9190), .ZN(n11871) );
  NAND2_X1 U10961 ( .A1(n11871), .A2(n8822), .ZN(n9193) );
  NAND2_X1 U10962 ( .A1(n9092), .A2(SI_28_), .ZN(n9192) );
  NOR2_X1 U10963 ( .A1(n9195), .A2(n9194), .ZN(n9196) );
  INV_X1 U10964 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n9199) );
  NAND2_X1 U10965 ( .A1(n9263), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9198) );
  NAND2_X1 U10966 ( .A1(n8812), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n9197) );
  OAI211_X1 U10967 ( .C1(n9199), .C2(n12992), .A(n9198), .B(n9197), .ZN(n9200)
         );
  OR2_X1 U10968 ( .A1(n9222), .A2(n13776), .ZN(n12969) );
  NAND2_X1 U10969 ( .A1(n9222), .A2(n13776), .ZN(n12970) );
  NAND2_X1 U10970 ( .A1(n13758), .A2(n13757), .ZN(n13760) );
  NAND2_X1 U10971 ( .A1(n9272), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9206) );
  NAND2_X1 U10972 ( .A1(n9213), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9208) );
  MUX2_X1 U10973 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9208), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n9209) );
  INV_X1 U10974 ( .A(n9210), .ZN(n9211) );
  NAND2_X1 U10975 ( .A1(n9211), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9212) );
  NAND2_X1 U10976 ( .A1(n10454), .A2(n10314), .ZN(n9215) );
  XNOR2_X1 U10977 ( .A(n13040), .B(n9215), .ZN(n9217) );
  NAND2_X1 U10978 ( .A1(n10454), .A2(n13733), .ZN(n9216) );
  NAND2_X1 U10979 ( .A1(n9217), .A2(n9216), .ZN(n10340) );
  INV_X1 U10980 ( .A(n13040), .ZN(n9221) );
  INV_X1 U10981 ( .A(n16200), .ZN(n16311) );
  NAND2_X1 U10982 ( .A1(n10314), .A2(n13733), .ZN(n12996) );
  INV_X1 U10983 ( .A(n12996), .ZN(n9315) );
  AND2_X1 U10984 ( .A1(n16311), .A2(n9315), .ZN(n9218) );
  NAND2_X1 U10985 ( .A1(n10340), .A2(n9218), .ZN(n9220) );
  AND2_X1 U10986 ( .A1(n12996), .A2(n13733), .ZN(n9219) );
  NAND2_X1 U10987 ( .A1(n13040), .A2(n9219), .ZN(n9302) );
  NAND2_X1 U10988 ( .A1(n9221), .A2(n13036), .ZN(n16274) );
  NAND2_X1 U10989 ( .A1(n11306), .A2(n11420), .ZN(n11535) );
  AND2_X1 U10990 ( .A1(n12888), .A2(n11535), .ZN(n9224) );
  NAND2_X1 U10991 ( .A1(n13620), .A2(n16182), .ZN(n11412) );
  AND2_X1 U10992 ( .A1(n9224), .A2(n11414), .ZN(n9232) );
  NAND2_X1 U10993 ( .A1(n13624), .A2(n16055), .ZN(n9225) );
  NAND2_X1 U10994 ( .A1(n16104), .A2(n7738), .ZN(n9226) );
  NAND2_X1 U10995 ( .A1(n16052), .A2(n16116), .ZN(n9227) );
  NAND2_X1 U10996 ( .A1(n13621), .A2(n11329), .ZN(n11216) );
  AND2_X1 U10997 ( .A1(n11216), .A2(n9230), .ZN(n9231) );
  NAND2_X1 U10998 ( .A1(n11217), .A2(n9231), .ZN(n11415) );
  NAND2_X1 U10999 ( .A1(n9232), .A2(n11415), .ZN(n11537) );
  NAND2_X1 U11000 ( .A1(n13618), .A2(n11309), .ZN(n9233) );
  NAND2_X1 U11001 ( .A1(n11537), .A2(n9233), .ZN(n11314) );
  NAND2_X1 U11002 ( .A1(n13617), .A2(n12895), .ZN(n9234) );
  NAND2_X1 U11003 ( .A1(n11313), .A2(n9234), .ZN(n11671) );
  NAND2_X1 U11004 ( .A1(n11860), .A2(n16257), .ZN(n9237) );
  NAND2_X1 U11005 ( .A1(n13614), .A2(n9238), .ZN(n9239) );
  NAND2_X1 U11006 ( .A1(n13959), .A2(n14031), .ZN(n9240) );
  NAND2_X1 U11007 ( .A1(n9241), .A2(n9240), .ZN(n13956) );
  NAND2_X1 U11008 ( .A1(n9242), .A2(n13942), .ZN(n12797) );
  INV_X1 U11009 ( .A(n13942), .ZN(n13475) );
  INV_X1 U11010 ( .A(n13927), .ZN(n13958) );
  OR2_X1 U11011 ( .A1(n14097), .A2(n13958), .ZN(n9243) );
  NAND2_X1 U11012 ( .A1(n13938), .A2(n9243), .ZN(n13923) );
  NAND2_X1 U11013 ( .A1(n14017), .A2(n13519), .ZN(n9245) );
  OR2_X1 U11014 ( .A1(n14005), .A2(n13873), .ZN(n9248) );
  NOR2_X1 U11015 ( .A1(n14001), .A2(n13887), .ZN(n9249) );
  INV_X1 U11016 ( .A(n14001), .ZN(n13878) );
  NAND2_X1 U11017 ( .A1(n13861), .A2(n13858), .ZN(n9251) );
  NAND2_X1 U11018 ( .A1(n14080), .A2(n13874), .ZN(n9250) );
  OR2_X1 U11019 ( .A1(n14074), .A2(n13862), .ZN(n12817) );
  NAND2_X1 U11020 ( .A1(n14068), .A2(n13611), .ZN(n9252) );
  NAND2_X1 U11021 ( .A1(n13823), .A2(n13825), .ZN(n9255) );
  INV_X1 U11022 ( .A(n13838), .ZN(n13815) );
  NAND2_X1 U11023 ( .A1(n13482), .A2(n13815), .ZN(n9254) );
  AND2_X1 U11024 ( .A1(n14058), .A2(n13610), .ZN(n9256) );
  NAND2_X1 U11025 ( .A1(n14048), .A2(n13801), .ZN(n9259) );
  NAND2_X1 U11026 ( .A1(n9260), .A2(n9259), .ZN(n13772) );
  NAND2_X1 U11027 ( .A1(n13040), .A2(n13021), .ZN(n9316) );
  NAND2_X1 U11028 ( .A1(n12863), .A2(n10453), .ZN(n13033) );
  INV_X1 U11029 ( .A(n13037), .ZN(n9951) );
  NAND2_X1 U11030 ( .A1(n9951), .A2(n13038), .ZN(n9954) );
  NAND2_X1 U11031 ( .A1(n9954), .A2(n9949), .ZN(n9261) );
  INV_X1 U11032 ( .A(n9261), .ZN(n10462) );
  NAND2_X1 U11033 ( .A1(n9951), .A2(P3_B_REG_SCAN_IN), .ZN(n9262) );
  NAND2_X1 U11034 ( .A1(n13943), .A2(n9262), .ZN(n13734) );
  INV_X1 U11035 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n9266) );
  NAND2_X1 U11036 ( .A1(n8812), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9265) );
  NAND2_X1 U11037 ( .A1(n9263), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9264) );
  OAI211_X1 U11038 ( .C1(n9266), .C2(n12992), .A(n9265), .B(n9264), .ZN(n9267)
         );
  INV_X1 U11039 ( .A(n9267), .ZN(n9268) );
  INV_X1 U11040 ( .A(n9269), .ZN(n9270) );
  NAND2_X1 U11041 ( .A1(n7469), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9275) );
  MUX2_X1 U11042 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9276), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n9277) );
  NAND2_X1 U11043 ( .A1(n9278), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9279) );
  MUX2_X1 U11044 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9279), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n9280) );
  AND2_X1 U11045 ( .A1(n9280), .A2(n7469), .ZN(n9282) );
  NAND3_X1 U11046 ( .A1(n9285), .A2(n9281), .A3(n9282), .ZN(n10332) );
  XNOR2_X1 U11047 ( .A(n11294), .B(P3_B_REG_SCAN_IN), .ZN(n9283) );
  NAND2_X1 U11048 ( .A1(n9283), .A2(n11393), .ZN(n9284) );
  INV_X1 U11049 ( .A(n9285), .ZN(n11597) );
  NAND2_X1 U11050 ( .A1(n11597), .A2(n11393), .ZN(n9286) );
  NAND2_X1 U11051 ( .A1(n11597), .A2(n11294), .ZN(n9288) );
  XNOR2_X1 U11052 ( .A(n14108), .B(n10457), .ZN(n9301) );
  NOR2_X1 U11053 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .ZN(
        n9293) );
  NOR4_X1 U11054 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n9292) );
  NOR4_X1 U11055 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n9291) );
  NOR4_X1 U11056 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n9290) );
  NAND4_X1 U11057 ( .A1(n9293), .A2(n9292), .A3(n9291), .A4(n9290), .ZN(n9299)
         );
  NOR4_X1 U11058 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n9297) );
  NOR4_X1 U11059 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n9296) );
  NOR4_X1 U11060 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n9295) );
  NOR4_X1 U11061 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n9294) );
  NAND4_X1 U11062 ( .A1(n9297), .A2(n9296), .A3(n9295), .A4(n9294), .ZN(n9298)
         );
  NOR2_X1 U11063 ( .A1(n9299), .A2(n9298), .ZN(n9300) );
  NAND2_X1 U11064 ( .A1(n12974), .A2(n12996), .ZN(n10333) );
  NAND2_X1 U11065 ( .A1(n12960), .A2(n9302), .ZN(n11086) );
  NAND2_X1 U11066 ( .A1(n10333), .A2(n11086), .ZN(n11085) );
  NAND2_X1 U11067 ( .A1(n11085), .A2(n14108), .ZN(n9307) );
  INV_X1 U11068 ( .A(n11086), .ZN(n9304) );
  NAND3_X1 U11069 ( .A1(n16200), .A2(n10314), .A3(n12996), .ZN(n9303) );
  NAND2_X1 U11070 ( .A1(n9304), .A2(n9303), .ZN(n9305) );
  INV_X1 U11071 ( .A(n14108), .ZN(n11084) );
  NAND2_X1 U11072 ( .A1(n9305), .A2(n11084), .ZN(n9306) );
  AND2_X1 U11073 ( .A1(n9307), .A2(n9306), .ZN(n9308) );
  INV_X1 U11074 ( .A(n9310), .ZN(n13746) );
  NOR2_X1 U11075 ( .A1(n16407), .A2(n9311), .ZN(n9312) );
  INV_X1 U11076 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9324) );
  AND2_X1 U11077 ( .A1(n12974), .A2(n9315), .ZN(n10633) );
  NAND2_X1 U11078 ( .A1(n10349), .A2(n10633), .ZN(n13039) );
  NAND2_X1 U11079 ( .A1(n10454), .A2(n10453), .ZN(n13034) );
  NOR2_X1 U11080 ( .A1(n9316), .A2(n13034), .ZN(n10341) );
  NAND2_X1 U11081 ( .A1(n10349), .A2(n10341), .ZN(n9317) );
  NAND2_X1 U11082 ( .A1(n13039), .A2(n9317), .ZN(n9318) );
  INV_X1 U11083 ( .A(n10457), .ZN(n14110) );
  AND3_X1 U11084 ( .A1(n14110), .A2(n14108), .A3(n9319), .ZN(n10348) );
  NAND2_X1 U11085 ( .A1(n9318), .A2(n10348), .ZN(n9322) );
  NAND2_X1 U11086 ( .A1(n10457), .A2(n9319), .ZN(n9320) );
  NOR2_X1 U11087 ( .A1(n9320), .A2(n14108), .ZN(n10345) );
  NAND3_X1 U11088 ( .A1(n10345), .A2(n10349), .A3(n10340), .ZN(n9321) );
  NOR2_X1 U11089 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), 
        .ZN(n9329) );
  NOR2_X2 U11090 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n9531) );
  NAND2_X1 U11091 ( .A1(n9531), .A2(n9618), .ZN(n9333) );
  NAND2_X1 U11092 ( .A1(n9543), .A2(n9335), .ZN(n9541) );
  NAND2_X1 U11093 ( .A1(n9341), .A2(n9529), .ZN(n9336) );
  XNOR2_X1 U11094 ( .A(n9341), .B(n9529), .ZN(n11721) );
  INV_X1 U11095 ( .A(n9600), .ZN(n9343) );
  NAND2_X1 U11096 ( .A1(n9542), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9342) );
  NAND2_X1 U11097 ( .A1(n9343), .A2(n11530), .ZN(n9550) );
  OR2_X2 U11098 ( .A1(n9550), .A2(P2_U3088), .ZN(n14267) );
  NAND2_X1 U11099 ( .A1(n9352), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9351) );
  MUX2_X1 U11100 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9351), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n9353) );
  AND2_X2 U11101 ( .A1(n9353), .A2(n9354), .ZN(n9698) );
  NAND2_X1 U11102 ( .A1(n9357), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9358) );
  INV_X1 U11103 ( .A(n10332), .ZN(n9359) );
  INV_X2 U11104 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NAND2_X2 U11105 ( .A1(n10095), .A2(P1_U3086), .ZN(n15262) );
  INV_X1 U11106 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10088) );
  NOR2_X1 U11107 ( .A1(n10095), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15248) );
  INV_X2 U11108 ( .A(n15248), .ZN(n15260) );
  XNOR2_X1 U11109 ( .A(n9366), .B(SI_1_), .ZN(n9378) );
  XNOR2_X1 U11110 ( .A(n9378), .B(n9377), .ZN(n10087) );
  INV_X1 U11111 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n15622) );
  NAND2_X1 U11112 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9361) );
  XNOR2_X1 U11113 ( .A(n15622), .B(n9361), .ZN(n14867) );
  OAI222_X1 U11114 ( .A1(n15262), .A2(n10088), .B1(n15260), .B2(n10087), .C1(
        n14867), .C2(P1_U3086), .ZN(P1_U3354) );
  INV_X1 U11115 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10102) );
  INV_X1 U11116 ( .A(SI_2_), .ZN(n15502) );
  OAI21_X1 U11117 ( .B1(SI_1_), .B2(n15502), .A(n9362), .ZN(n9364) );
  OAI21_X1 U11118 ( .B1(SI_2_), .B2(n9457), .A(n9366), .ZN(n9363) );
  NAND2_X1 U11119 ( .A1(n9364), .A2(n9363), .ZN(n9369) );
  INV_X1 U11120 ( .A(n9377), .ZN(n9365) );
  OAI211_X1 U11121 ( .C1(SI_1_), .C2(n9366), .A(n9365), .B(n15502), .ZN(n9368)
         );
  NAND2_X1 U11122 ( .A1(n9366), .A2(SI_1_), .ZN(n9376) );
  NAND3_X1 U11123 ( .A1(n9376), .A2(SI_2_), .A3(n9377), .ZN(n9367) );
  MUX2_X1 U11124 ( .A(n10102), .B(n9721), .S(n12709), .Z(n9373) );
  XNOR2_X1 U11125 ( .A(n9375), .B(n9373), .ZN(n10101) );
  INV_X1 U11126 ( .A(n10101), .ZN(n9406) );
  INV_X1 U11127 ( .A(n9370), .ZN(n9371) );
  NAND2_X1 U11128 ( .A1(n9371), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9372) );
  XNOR2_X1 U11129 ( .A(n9372), .B(n15627), .ZN(n10103) );
  OAI222_X1 U11130 ( .A1(n15262), .A2(n10102), .B1(n15260), .B2(n9406), .C1(
        P1_U3086), .C2(n10103), .ZN(P1_U3353) );
  INV_X1 U11131 ( .A(n9373), .ZN(n9374) );
  NAND2_X1 U11132 ( .A1(n9375), .A2(n9374), .ZN(n9381) );
  OAI21_X1 U11133 ( .B1(n9378), .B2(n9377), .A(n9376), .ZN(n9379) );
  NAND2_X1 U11134 ( .A1(n9379), .A2(SI_2_), .ZN(n9380) );
  XNOR2_X1 U11135 ( .A(n9387), .B(SI_3_), .ZN(n9384) );
  XNOR2_X1 U11136 ( .A(n9386), .B(n9384), .ZN(n10721) );
  INV_X1 U11137 ( .A(n10721), .ZN(n9394) );
  NAND2_X1 U11138 ( .A1(n9382), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9383) );
  XNOR2_X1 U11139 ( .A(n9383), .B(n9344), .ZN(n10722) );
  OAI222_X1 U11140 ( .A1(n15262), .A2(n8047), .B1(n15260), .B2(n9394), .C1(
        P1_U3086), .C2(n10722), .ZN(P1_U3352) );
  INV_X1 U11141 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9391) );
  INV_X1 U11142 ( .A(n9384), .ZN(n9385) );
  NAND2_X1 U11143 ( .A1(n9387), .A2(SI_3_), .ZN(n9388) );
  MUX2_X1 U11144 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n12709), .Z(n9409) );
  XNOR2_X1 U11145 ( .A(n9409), .B(SI_4_), .ZN(n9407) );
  INV_X1 U11146 ( .A(n10865), .ZN(n9398) );
  NAND2_X1 U11147 ( .A1(n9389), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9390) );
  XNOR2_X1 U11148 ( .A(n9390), .B(P1_IR_REG_4__SCAN_IN), .ZN(n16003) );
  INV_X1 U11149 ( .A(n16003), .ZN(n16021) );
  OAI222_X1 U11150 ( .A1(n15262), .A2(n9391), .B1(n15260), .B2(n9398), .C1(
        P1_U3086), .C2(n16021), .ZN(P1_U3351) );
  INV_X2 U11151 ( .A(n11529), .ZN(n14691) );
  OR2_X1 U11152 ( .A1(n9396), .A2(n14676), .ZN(n9392) );
  XNOR2_X1 U11153 ( .A(n9392), .B(P2_IR_REG_3__SCAN_IN), .ZN(n9729) );
  AOI22_X1 U11154 ( .A1(n9729), .A2(P2_STATE_REG_SCAN_IN), .B1(n14685), .B2(
        P1_DATAO_REG_3__SCAN_IN), .ZN(n9393) );
  OAI21_X1 U11155 ( .B1(n9394), .B2(n14691), .A(n9393), .ZN(P2_U3324) );
  INV_X2 U11156 ( .A(n14685), .ZN(n14693) );
  NAND2_X1 U11157 ( .A1(n9396), .A2(n9395), .ZN(n9415) );
  NAND2_X1 U11158 ( .A1(n9415), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9397) );
  XNOR2_X1 U11159 ( .A(n9397), .B(P2_IR_REG_4__SCAN_IN), .ZN(n9784) );
  INV_X1 U11160 ( .A(n9784), .ZN(n9583) );
  OAI222_X1 U11161 ( .A1(n14693), .A2(n9399), .B1(n14691), .B2(n9398), .C1(
        P2_U3088), .C2(n9583), .ZN(P2_U3323) );
  INV_X1 U11162 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n9401) );
  NAND2_X1 U11163 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9400) );
  OAI222_X1 U11164 ( .A1(n14693), .A2(n9402), .B1(n14691), .B2(n10087), .C1(
        n15786), .C2(P2_U3088), .ZN(P2_U3326) );
  OAI222_X1 U11165 ( .A1(n14693), .A2(n9721), .B1(n14691), .B2(n9406), .C1(
        P2_U3088), .C2(n9723), .ZN(P2_U3325) );
  INV_X1 U11166 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9414) );
  INV_X1 U11167 ( .A(n9407), .ZN(n9408) );
  MUX2_X1 U11168 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n12298), .Z(n9425) );
  XNOR2_X1 U11169 ( .A(n9425), .B(SI_5_), .ZN(n9422) );
  XNOR2_X1 U11170 ( .A(n9424), .B(n9422), .ZN(n10869) );
  INV_X1 U11171 ( .A(n10869), .ZN(n9417) );
  INV_X1 U11172 ( .A(n9410), .ZN(n9412) );
  NAND2_X1 U11173 ( .A1(n9412), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9411) );
  MUX2_X1 U11174 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9411), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n9413) );
  AND2_X1 U11175 ( .A1(n9413), .A2(n9432), .ZN(n10870) );
  INV_X1 U11176 ( .A(n10870), .ZN(n9964) );
  OAI222_X1 U11177 ( .A1(n15262), .A2(n9414), .B1(n15260), .B2(n9417), .C1(
        P1_U3086), .C2(n9964), .ZN(P1_U3350) );
  OR2_X1 U11178 ( .A1(n9495), .A2(n14676), .ZN(n9416) );
  XNOR2_X1 U11179 ( .A(n9416), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9817) );
  INV_X1 U11180 ( .A(n9817), .ZN(n9574) );
  OAI222_X1 U11181 ( .A1(n14693), .A2(n9418), .B1(n14691), .B2(n9417), .C1(
        P2_U3088), .C2(n9574), .ZN(P2_U3322) );
  INV_X1 U11182 ( .A(n10076), .ZN(n10268) );
  INV_X1 U11183 ( .A(n9420), .ZN(n9421) );
  OAI222_X1 U11184 ( .A1(n10268), .A2(P3_U3151), .B1(n14119), .B2(n9421), .C1(
        n15502), .C2(n13462), .ZN(P3_U3293) );
  INV_X1 U11185 ( .A(n9422), .ZN(n9423) );
  NAND2_X1 U11186 ( .A1(n9425), .A2(SI_5_), .ZN(n9426) );
  MUX2_X1 U11187 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n12298), .Z(n9447) );
  XNOR2_X1 U11188 ( .A(n9447), .B(SI_6_), .ZN(n9444) );
  XNOR2_X1 U11189 ( .A(n9446), .B(n9444), .ZN(n10879) );
  INV_X1 U11190 ( .A(n10879), .ZN(n9436) );
  NAND2_X1 U11191 ( .A1(n9495), .A2(n9427), .ZN(n9450) );
  NAND2_X1 U11192 ( .A1(n9450), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9428) );
  XNOR2_X1 U11193 ( .A(n9428), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10022) );
  INV_X1 U11194 ( .A(n10022), .ZN(n9429) );
  OAI222_X1 U11195 ( .A1(n14693), .A2(n9430), .B1(n14691), .B2(n9436), .C1(
        P2_U3088), .C2(n9429), .ZN(P2_U3321) );
  NAND2_X1 U11196 ( .A1(n9432), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9431) );
  MUX2_X1 U11197 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9431), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n9435) );
  INV_X1 U11198 ( .A(n9432), .ZN(n9434) );
  INV_X1 U11199 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9433) );
  NAND2_X1 U11200 ( .A1(n9434), .A2(n9433), .ZN(n9468) );
  NAND2_X1 U11201 ( .A1(n9435), .A2(n9468), .ZN(n10011) );
  OAI222_X1 U11202 ( .A1(n15262), .A2(n9437), .B1(n15260), .B2(n9436), .C1(
        P1_U3086), .C2(n10011), .ZN(P1_U3349) );
  INV_X1 U11203 ( .A(n14119), .ZN(n16291) );
  INV_X1 U11204 ( .A(n13462), .ZN(n16290) );
  AOI222_X1 U11205 ( .A1(n9438), .A2(n16291), .B1(SI_9_), .B2(n16290), .C1(
        n11121), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9439) );
  INV_X1 U11206 ( .A(n9439), .ZN(P3_U3286) );
  AOI222_X1 U11207 ( .A1(n9440), .A2(n16291), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10289), .C1(SI_3_), .C2(n16290), .ZN(n9441) );
  INV_X1 U11208 ( .A(n9441), .ZN(P3_U3292) );
  AOI222_X1 U11209 ( .A1(n9442), .A2(n16291), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10497), .C1(SI_5_), .C2(n16290), .ZN(n9443) );
  INV_X1 U11210 ( .A(n9443), .ZN(P3_U3290) );
  INV_X1 U11211 ( .A(n9444), .ZN(n9445) );
  MUX2_X1 U11212 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n12298), .Z(n9466) );
  XNOR2_X1 U11213 ( .A(n9466), .B(SI_7_), .ZN(n9463) );
  XNOR2_X1 U11214 ( .A(n9465), .B(n9463), .ZN(n11045) );
  INV_X1 U11215 ( .A(n11045), .ZN(n9453) );
  NAND2_X1 U11216 ( .A1(n9468), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9448) );
  XNOR2_X1 U11217 ( .A(n9448), .B(P1_IR_REG_7__SCAN_IN), .ZN(n14883) );
  INV_X1 U11218 ( .A(n14883), .ZN(n9975) );
  OAI222_X1 U11219 ( .A1(n15262), .A2(n9449), .B1(n15260), .B2(n9453), .C1(
        P1_U3086), .C2(n9975), .ZN(P1_U3348) );
  INV_X1 U11220 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9454) );
  NAND2_X1 U11221 ( .A1(n9476), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9451) );
  XNOR2_X1 U11222 ( .A(n9451), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10397) );
  INV_X1 U11223 ( .A(n10397), .ZN(n9452) );
  OAI222_X1 U11224 ( .A1(n14693), .A2(n9454), .B1(n14691), .B2(n9453), .C1(
        P2_U3088), .C2(n9452), .ZN(P2_U3320) );
  AOI22_X1 U11225 ( .A1(n16291), .A2(n9455), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n8065), .ZN(n9456) );
  OAI21_X1 U11226 ( .B1(n9457), .B2(n13462), .A(n9456), .ZN(P3_U3294) );
  INV_X1 U11227 ( .A(n9458), .ZN(n9460) );
  INV_X1 U11228 ( .A(SI_6_), .ZN(n9459) );
  OAI222_X1 U11229 ( .A1(P3_U3151), .A2(n10573), .B1(n14119), .B2(n9460), .C1(
        n9459), .C2(n13462), .ZN(P3_U3289) );
  INV_X1 U11230 ( .A(SI_7_), .ZN(n9462) );
  OAI222_X1 U11231 ( .A1(P3_U3151), .A2(n10562), .B1(n13462), .B2(n9462), .C1(
        n14119), .C2(n9461), .ZN(P3_U3288) );
  INV_X1 U11232 ( .A(n9463), .ZN(n9464) );
  NAND2_X1 U11233 ( .A1(n9466), .A2(SI_7_), .ZN(n9467) );
  MUX2_X1 U11234 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n12298), .Z(n9486) );
  XNOR2_X1 U11235 ( .A(n9486), .B(SI_8_), .ZN(n9483) );
  XNOR2_X1 U11236 ( .A(n9485), .B(n9483), .ZN(n11356) );
  INV_X1 U11237 ( .A(n11356), .ZN(n9479) );
  NAND2_X1 U11238 ( .A1(n9526), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9487) );
  XNOR2_X1 U11239 ( .A(n9487), .B(P1_IR_REG_8__SCAN_IN), .ZN(n11357) );
  INV_X1 U11240 ( .A(n15262), .ZN(n10530) );
  AOI22_X1 U11241 ( .A1(n11357), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10530), .ZN(n9469) );
  OAI21_X1 U11242 ( .B1(n9479), .B2(n15260), .A(n9469), .ZN(P1_U3347) );
  OAI222_X1 U11243 ( .A1(P3_U3151), .A2(n11466), .B1(n13462), .B2(n9519), .C1(
        n14119), .C2(n9470), .ZN(P3_U3284) );
  OAI222_X1 U11244 ( .A1(P3_U3151), .A2(n15926), .B1(n13462), .B2(n15485), 
        .C1(n14119), .C2(n9471), .ZN(P3_U3283) );
  INV_X1 U11245 ( .A(SI_8_), .ZN(n9472) );
  OAI222_X1 U11246 ( .A1(n14119), .A2(n9473), .B1(n13462), .B2(n9472), .C1(
        P3_U3151), .C2(n10958), .ZN(P3_U3287) );
  INV_X1 U11247 ( .A(n9474), .ZN(n9475) );
  OAI222_X1 U11248 ( .A1(n10485), .A2(P3_U3151), .B1(n14119), .B2(n9475), .C1(
        n15495), .C2(n13462), .ZN(P3_U3291) );
  INV_X1 U11249 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9480) );
  NAND2_X1 U11250 ( .A1(n9492), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9477) );
  XNOR2_X1 U11251 ( .A(n9477), .B(P2_IR_REG_8__SCAN_IN), .ZN(n15822) );
  INV_X1 U11252 ( .A(n15822), .ZN(n9478) );
  OAI222_X1 U11253 ( .A1(n14693), .A2(n9480), .B1(n14691), .B2(n9479), .C1(
        P2_U3088), .C2(n9478), .ZN(P2_U3319) );
  INV_X1 U11254 ( .A(SI_13_), .ZN(n9482) );
  OAI222_X1 U11255 ( .A1(P3_U3151), .A2(n15944), .B1(n13462), .B2(n9482), .C1(
        n14119), .C2(n9481), .ZN(P3_U3282) );
  INV_X1 U11256 ( .A(n9483), .ZN(n9484) );
  MUX2_X1 U11257 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n12298), .Z(n9504) );
  INV_X1 U11258 ( .A(n11362), .ZN(n9497) );
  NAND2_X1 U11259 ( .A1(n9487), .A2(n15635), .ZN(n9488) );
  NAND2_X1 U11260 ( .A1(n9488), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9489) );
  NAND2_X1 U11261 ( .A1(n9489), .A2(n9523), .ZN(n9507) );
  OR2_X1 U11262 ( .A1(n9489), .A2(n9523), .ZN(n9490) );
  AOI22_X1 U11263 ( .A1(n11363), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n10530), .ZN(n9491) );
  OAI21_X1 U11264 ( .B1(n9497), .B2(n15260), .A(n9491), .ZN(P1_U3346) );
  INV_X1 U11265 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9498) );
  OAI21_X1 U11266 ( .B1(n9492), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9493) );
  MUX2_X1 U11267 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9493), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n9496) );
  NAND2_X1 U11268 ( .A1(n9495), .A2(n9494), .ZN(n9674) );
  INV_X1 U11269 ( .A(n10797), .ZN(n10189) );
  OAI222_X1 U11270 ( .A1(n14693), .A2(n9498), .B1(n14691), .B2(n9497), .C1(
        P2_U3088), .C2(n10189), .ZN(P2_U3318) );
  OAI222_X1 U11271 ( .A1(P3_U3151), .A2(n15958), .B1(n13462), .B2(n9871), .C1(
        n14119), .C2(n9499), .ZN(P3_U3281) );
  AND2_X1 U11272 ( .A1(n9501), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U11273 ( .A1(n9501), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U11274 ( .A1(n9501), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U11275 ( .A1(n9501), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U11276 ( .A1(n9501), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U11277 ( .A1(n9501), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U11278 ( .A1(n9501), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U11279 ( .A1(n9501), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U11280 ( .A1(n9501), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U11281 ( .A1(n9501), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U11282 ( .A1(n9501), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U11283 ( .A1(n9501), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U11284 ( .A1(n9501), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U11285 ( .A1(n9501), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U11286 ( .A1(n9501), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U11287 ( .A1(n9501), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U11288 ( .A1(n9501), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U11289 ( .A1(n9501), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U11290 ( .A1(n9501), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U11291 ( .A1(n9501), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U11292 ( .A1(n9501), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U11293 ( .A1(n9501), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U11294 ( .A1(n9501), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U11295 ( .A1(n9501), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U11296 ( .A1(n9501), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U11297 ( .A1(n9501), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U11298 ( .A1(n9501), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U11299 ( .A1(n9501), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U11300 ( .A1(n9501), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U11301 ( .A1(n9501), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  OAI222_X1 U11302 ( .A1(P3_U3151), .A2(n15983), .B1(n13462), .B2(n10244), 
        .C1(n14119), .C2(n9502), .ZN(P3_U3280) );
  NAND2_X1 U11303 ( .A1(n9505), .A2(SI_9_), .ZN(n9506) );
  MUX2_X1 U11304 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n12298), .Z(n9516) );
  XNOR2_X1 U11305 ( .A(n9516), .B(SI_10_), .ZN(n9513) );
  XNOR2_X1 U11306 ( .A(n9515), .B(n9513), .ZN(n11545) );
  INV_X1 U11307 ( .A(n11545), .ZN(n9511) );
  NAND2_X1 U11308 ( .A1(n9507), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9508) );
  XNOR2_X1 U11309 ( .A(n9508), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11546) );
  INV_X1 U11310 ( .A(n11546), .ZN(n10452) );
  OAI222_X1 U11311 ( .A1(n15262), .A2(n9509), .B1(n15260), .B2(n9511), .C1(
        P1_U3086), .C2(n10452), .ZN(P1_U3345) );
  INV_X1 U11312 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9512) );
  NAND2_X1 U11313 ( .A1(n9674), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9510) );
  XNOR2_X1 U11314 ( .A(n9510), .B(P2_IR_REG_10__SCAN_IN), .ZN(n11134) );
  INV_X1 U11315 ( .A(n11134), .ZN(n10652) );
  OAI222_X1 U11316 ( .A1(n14693), .A2(n9512), .B1(n14691), .B2(n9511), .C1(
        P2_U3088), .C2(n10652), .ZN(P2_U3317) );
  INV_X1 U11317 ( .A(n9513), .ZN(n9514) );
  NAND2_X1 U11318 ( .A1(n9516), .A2(SI_10_), .ZN(n9517) );
  MUX2_X1 U11319 ( .A(n9518), .B(n9678), .S(n12298), .Z(n9520) );
  NAND2_X1 U11320 ( .A1(n9520), .A2(n9519), .ZN(n9713) );
  INV_X1 U11321 ( .A(n9520), .ZN(n9521) );
  NAND2_X1 U11322 ( .A1(n9521), .A2(SI_11_), .ZN(n9522) );
  NAND2_X1 U11323 ( .A1(n9713), .A2(n9522), .ZN(n9711) );
  XNOR2_X1 U11324 ( .A(n9712), .B(n9711), .ZN(n11550) );
  INV_X1 U11325 ( .A(n11550), .ZN(n9677) );
  NAND3_X1 U11326 ( .A1(n15635), .A2(n9524), .A3(n9523), .ZN(n9525) );
  NAND2_X1 U11327 ( .A1(n9718), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9527) );
  XNOR2_X1 U11328 ( .A(n9527), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U11329 ( .A1(n11551), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10530), .ZN(n9528) );
  OAI21_X1 U11330 ( .B1(n9677), .B2(n15260), .A(n9528), .ZN(P1_U3344) );
  NOR2_X1 U11331 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n9530) );
  NOR2_X1 U11332 ( .A1(n9543), .A2(n14676), .ZN(n9617) );
  INV_X1 U11333 ( .A(n9617), .ZN(n9544) );
  NAND2_X1 U11334 ( .A1(n9670), .A2(n11530), .ZN(n9548) );
  NAND2_X1 U11335 ( .A1(n9548), .A2(n11830), .ZN(n9549) );
  AND2_X1 U11336 ( .A1(n9547), .A2(n9558), .ZN(n15785) );
  INV_X1 U11337 ( .A(n9723), .ZN(n15809) );
  INV_X1 U11338 ( .A(n15786), .ZN(n9562) );
  INV_X1 U11339 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9551) );
  NAND2_X1 U11340 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n15795) );
  NOR2_X1 U11341 ( .A1(n15794), .A2(n15795), .ZN(n15793) );
  INV_X1 U11342 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9552) );
  MUX2_X1 U11343 ( .A(n9552), .B(P2_REG2_REG_2__SCAN_IN), .S(n9723), .Z(n9553)
         );
  INV_X1 U11344 ( .A(n9553), .ZN(n15805) );
  NOR2_X1 U11345 ( .A1(n15806), .A2(n15805), .ZN(n15804) );
  AOI21_X1 U11346 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n15809), .A(n15804), .ZN(
        n9687) );
  INV_X1 U11347 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9554) );
  MUX2_X1 U11348 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n9554), .S(n9729), .Z(n9555)
         );
  INV_X1 U11349 ( .A(n9555), .ZN(n9686) );
  NOR2_X1 U11350 ( .A1(n9687), .A2(n9686), .ZN(n9685) );
  INV_X1 U11351 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9556) );
  MUX2_X1 U11352 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n9556), .S(n9784), .Z(n9557)
         );
  INV_X1 U11353 ( .A(n9557), .ZN(n9576) );
  NOR2_X1 U11354 ( .A1(n9577), .A2(n9576), .ZN(n9575) );
  AOI21_X1 U11355 ( .B1(n9784), .B2(P2_REG2_REG_4__SCAN_IN), .A(n9575), .ZN(
        n9560) );
  XNOR2_X1 U11356 ( .A(n9817), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n9559) );
  NOR2_X1 U11357 ( .A1(n9547), .A2(P2_U3088), .ZN(n14684) );
  NAND2_X1 U11358 ( .A1(n9558), .A2(n14684), .ZN(n9566) );
  NOR2_X1 U11359 ( .A1(n9560), .A2(n9559), .ZN(n9587) );
  AOI211_X1 U11360 ( .C1(n9560), .C2(n9559), .A(n15817), .B(n9587), .ZN(n9570)
         );
  INV_X1 U11361 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9561) );
  MUX2_X1 U11362 ( .A(n9561), .B(P2_REG1_REG_1__SCAN_IN), .S(n15786), .Z(
        n15789) );
  INV_X1 U11363 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9563) );
  MUX2_X1 U11364 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n9563), .S(n9723), .Z(n15802) );
  NOR2_X1 U11365 ( .A1(n15803), .A2(n15802), .ZN(n15801) );
  INV_X1 U11366 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9564) );
  MUX2_X1 U11367 ( .A(n9564), .B(P2_REG1_REG_3__SCAN_IN), .S(n9729), .Z(n9683)
         );
  NOR2_X1 U11368 ( .A1(n9684), .A2(n9683), .ZN(n9682) );
  INV_X1 U11369 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9565) );
  MUX2_X1 U11370 ( .A(n9565), .B(P2_REG1_REG_4__SCAN_IN), .S(n9784), .Z(n9579)
         );
  XNOR2_X1 U11371 ( .A(n9817), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n9567) );
  INV_X1 U11372 ( .A(n14314), .ZN(n13458) );
  AOI211_X1 U11373 ( .C1(n9568), .C2(n9567), .A(n15813), .B(n9590), .ZN(n9569)
         );
  NOR2_X1 U11374 ( .A1(n9570), .A2(n9569), .ZN(n9573) );
  AND2_X1 U11375 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n9836) );
  AOI21_X1 U11376 ( .B1(n15800), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n9836), .ZN(
        n9572) );
  OAI211_X1 U11377 ( .C1(n9574), .C2(n14306), .A(n9573), .B(n9572), .ZN(
        P2_U3219) );
  AOI211_X1 U11378 ( .C1(n9577), .C2(n9576), .A(n9575), .B(n15817), .ZN(n9586)
         );
  AOI211_X1 U11379 ( .C1(n9580), .C2(n9579), .A(n9578), .B(n15813), .ZN(n9585)
         );
  NAND2_X1 U11380 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n9582) );
  NAND2_X1 U11381 ( .A1(n15800), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n9581) );
  OAI211_X1 U11382 ( .C1(n14306), .C2(n9583), .A(n9582), .B(n9581), .ZN(n9584)
         );
  OR3_X1 U11383 ( .A1(n9586), .A2(n9585), .A3(n9584), .ZN(P2_U3218) );
  XNOR2_X1 U11384 ( .A(n10022), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n9588) );
  NOR2_X1 U11385 ( .A1(n9589), .A2(n9588), .ZN(n9758) );
  AOI211_X1 U11386 ( .C1(n9589), .C2(n9588), .A(n15817), .B(n9758), .ZN(n9599)
         );
  INV_X1 U11387 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9591) );
  MUX2_X1 U11388 ( .A(n9591), .B(P2_REG1_REG_6__SCAN_IN), .S(n10022), .Z(n9592) );
  NOR2_X1 U11389 ( .A1(n9593), .A2(n9592), .ZN(n9761) );
  AOI211_X1 U11390 ( .C1(n9593), .C2(n9592), .A(n15813), .B(n9761), .ZN(n9598)
         );
  INV_X1 U11391 ( .A(n15800), .ZN(n15844) );
  INV_X1 U11392 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n9596) );
  NAND2_X1 U11393 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n9595) );
  NAND2_X1 U11394 ( .A1(n15838), .A2(n10022), .ZN(n9594) );
  OAI211_X1 U11395 ( .C1(n15844), .C2(n9596), .A(n9595), .B(n9594), .ZN(n9597)
         );
  OR3_X1 U11396 ( .A1(n9599), .A2(n9598), .A3(n9597), .ZN(P2_U3220) );
  INV_X1 U11397 ( .A(P2_B_REG_SCAN_IN), .ZN(n14313) );
  XOR2_X1 U11398 ( .A(n14313), .B(n11721), .Z(n9601) );
  AND2_X1 U11399 ( .A1(n14690), .A2(n9601), .ZN(n9602) );
  OR2_X1 U11400 ( .A1(n14688), .A2(n9602), .ZN(n9614) );
  INV_X1 U11401 ( .A(n9614), .ZN(n15779) );
  INV_X1 U11402 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15778) );
  AOI22_X1 U11403 ( .A1(n15779), .A2(n15778), .B1(n14688), .B2(n14690), .ZN(
        n9801) );
  NOR4_X1 U11404 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n9606) );
  NOR4_X1 U11405 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n9605) );
  NOR4_X1 U11406 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n9604) );
  NOR4_X1 U11407 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9603) );
  NAND4_X1 U11408 ( .A1(n9606), .A2(n9605), .A3(n9604), .A4(n9603), .ZN(n9612)
         );
  NOR2_X1 U11409 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n9610) );
  NOR4_X1 U11410 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9609) );
  NOR4_X1 U11411 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n9608) );
  NOR4_X1 U11412 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n9607) );
  NAND4_X1 U11413 ( .A1(n9610), .A2(n9609), .A3(n9608), .A4(n9607), .ZN(n9611)
         );
  OAI21_X1 U11414 ( .B1(n9612), .B2(n9611), .A(n15779), .ZN(n9803) );
  NAND2_X1 U11415 ( .A1(n9801), .A2(n9803), .ZN(n9644) );
  INV_X1 U11416 ( .A(n9644), .ZN(n9613) );
  AND2_X1 U11417 ( .A1(n15784), .A2(n9613), .ZN(n10202) );
  NOR2_X1 U11418 ( .A1(n9614), .A2(P2_D_REG_0__SCAN_IN), .ZN(n9616) );
  AND2_X1 U11419 ( .A1(n14688), .A2(n11721), .ZN(n9615) );
  INV_X1 U11420 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9622) );
  NAND2_X1 U11421 ( .A1(n9628), .A2(n9627), .ZN(n9621) );
  NAND2_X1 U11422 ( .A1(n9621), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9623) );
  NAND2_X1 U11423 ( .A1(n9623), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n9624) );
  NAND2_X1 U11424 ( .A1(n9809), .A2(n13421), .ZN(n10418) );
  NOR2_X1 U11425 ( .A1(n15783), .A2(n10418), .ZN(n9626) );
  NAND2_X1 U11426 ( .A1(n10202), .A2(n9626), .ZN(n9630) );
  XNOR2_X1 U11427 ( .A(n9628), .B(n9627), .ZN(n9660) );
  INV_X1 U11428 ( .A(n9802), .ZN(n9629) );
  INV_X1 U11429 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9633) );
  NAND2_X1 U11430 ( .A1(n10095), .A2(SI_0_), .ZN(n9632) );
  XNOR2_X1 U11431 ( .A(n9632), .B(n9631), .ZN(n14694) );
  MUX2_X1 U11432 ( .A(n9633), .B(n14694), .S(n11830), .Z(n13121) );
  NOR2_X1 U11433 ( .A1(n15783), .A2(n13351), .ZN(n9634) );
  NAND2_X1 U11434 ( .A1(n9670), .A2(n9547), .ZN(n14523) );
  NAND2_X1 U11435 ( .A1(n14195), .A2(n14439), .ZN(n14217) );
  INV_X1 U11436 ( .A(n14217), .ZN(n14225) );
  AND2_X2 U11437 ( .A1(n9638), .A2(n9639), .ZN(n9789) );
  NAND2_X1 U11438 ( .A1(n9789), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9643) );
  INV_X1 U11439 ( .A(n9639), .ZN(n14680) );
  AND2_X4 U11440 ( .A1(n14680), .A2(n9638), .ZN(n9742) );
  NAND2_X1 U11441 ( .A1(n9742), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9642) );
  NAND2_X1 U11442 ( .A1(n9732), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n9641) );
  NAND2_X1 U11443 ( .A1(n9744), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9640) );
  OAI21_X1 U11444 ( .B1(n15783), .B2(n9644), .A(n9802), .ZN(n9647) );
  NAND2_X1 U11445 ( .A1(n9670), .A2(n13351), .ZN(n10200) );
  AND2_X1 U11446 ( .A1(n9645), .A2(n10200), .ZN(n9646) );
  NAND2_X1 U11447 ( .A1(n9647), .A2(n9646), .ZN(n9741) );
  OR2_X1 U11448 ( .A1(n9741), .A2(P2_U3088), .ZN(n14226) );
  AOI22_X1 U11449 ( .A1(n14225), .A2(n14266), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n14226), .ZN(n9658) );
  NAND2_X1 U11450 ( .A1(n9809), .A2(n13351), .ZN(n16353) );
  INV_X1 U11451 ( .A(n9670), .ZN(n9648) );
  NAND2_X1 U11452 ( .A1(n16353), .A2(n9648), .ZN(n9649) );
  NOR2_X1 U11453 ( .A1(n15783), .A2(n9649), .ZN(n9650) );
  INV_X1 U11454 ( .A(n14248), .ZN(n14232) );
  NAND2_X1 U11455 ( .A1(n9742), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9654) );
  NAND2_X1 U11456 ( .A1(n9732), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n9653) );
  NAND2_X1 U11457 ( .A1(n9789), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n9652) );
  NAND2_X1 U11458 ( .A1(n9744), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9651) );
  INV_X1 U11459 ( .A(n13121), .ZN(n9890) );
  AND2_X1 U11460 ( .A1(n14268), .A2(n9890), .ZN(n9889) );
  NAND2_X1 U11461 ( .A1(n9889), .A2(n7431), .ZN(n9662) );
  INV_X1 U11462 ( .A(n14268), .ZN(n9655) );
  OAI21_X1 U11463 ( .B1(n9655), .B2(n14507), .A(n13121), .ZN(n9656) );
  NAND3_X1 U11464 ( .A1(n14232), .A2(n9662), .A3(n9656), .ZN(n9657) );
  OAI211_X1 U11465 ( .C1(n12244), .C2(n13121), .A(n9658), .B(n9657), .ZN(
        P2_U3204) );
  NAND2_X1 U11466 ( .A1(n10793), .A2(n13350), .ZN(n13116) );
  NAND2_X1 U11467 ( .A1(n13090), .A2(n9660), .ZN(n9661) );
  INV_X1 U11468 ( .A(n8716), .ZN(n9823) );
  XNOR2_X1 U11469 ( .A(n14547), .B(n9823), .ZN(n9724) );
  NOR2_X1 U11470 ( .A1(n9664), .A2(n9663), .ZN(n14231) );
  AOI21_X1 U11471 ( .B1(n9664), .B2(n9663), .A(n14231), .ZN(n9673) );
  NAND2_X1 U11472 ( .A1(n9742), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9668) );
  NAND2_X1 U11473 ( .A1(n9732), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n9667) );
  NAND2_X1 U11474 ( .A1(n9789), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n9666) );
  NAND2_X1 U11475 ( .A1(n9744), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9665) );
  AOI22_X1 U11476 ( .A1(n14225), .A2(n14265), .B1(n14547), .B2(n14246), .ZN(
        n9672) );
  INV_X1 U11477 ( .A(n9547), .ZN(n9669) );
  NAND2_X1 U11478 ( .A1(n14195), .A2(n14438), .ZN(n14219) );
  INV_X1 U11479 ( .A(n14219), .ZN(n14227) );
  AOI22_X1 U11480 ( .A1(n14227), .A2(n14268), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n14226), .ZN(n9671) );
  OAI211_X1 U11481 ( .C1(n9673), .C2(n14248), .A(n9672), .B(n9671), .ZN(
        P2_U3194) );
  NAND2_X1 U11482 ( .A1(n9754), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9675) );
  XNOR2_X1 U11483 ( .A(n9675), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11243) );
  INV_X1 U11484 ( .A(n11243), .ZN(n9676) );
  OAI222_X1 U11485 ( .A1(n14693), .A2(n9678), .B1(n14691), .B2(n9677), .C1(
        P2_U3088), .C2(n9676), .ZN(P2_U3316) );
  INV_X1 U11486 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15864) );
  INV_X1 U11487 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9679) );
  NOR2_X1 U11488 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9679), .ZN(n9749) );
  INV_X1 U11489 ( .A(n9749), .ZN(n9681) );
  NAND2_X1 U11490 ( .A1(n15838), .A2(n9729), .ZN(n9680) );
  OAI211_X1 U11491 ( .C1(n15844), .C2(n15864), .A(n9681), .B(n9680), .ZN(n9690) );
  AOI211_X1 U11492 ( .C1(n9684), .C2(n9683), .A(n9682), .B(n15813), .ZN(n9689)
         );
  AOI211_X1 U11493 ( .C1(n9687), .C2(n9686), .A(n9685), .B(n15817), .ZN(n9688)
         );
  OR3_X1 U11494 ( .A1(n9690), .A2(n9689), .A3(n9688), .ZN(P2_U3217) );
  AOI22_X1 U11495 ( .A1(n13706), .A2(P3_STATE_REG_SCAN_IN), .B1(SI_17_), .B2(
        n16290), .ZN(n9691) );
  OAI21_X1 U11496 ( .B1(n9692), .B2(n14119), .A(n9691), .ZN(P3_U3278) );
  INV_X1 U11497 ( .A(P1_B_REG_SCAN_IN), .ZN(n13077) );
  NAND2_X1 U11498 ( .A1(n9698), .A2(n13077), .ZN(n9693) );
  INV_X1 U11499 ( .A(n9700), .ZN(n15258) );
  INV_X1 U11500 ( .A(n9698), .ZN(n11720) );
  NAND3_X1 U11501 ( .A1(n15258), .A2(P1_B_REG_SCAN_IN), .A3(n11720), .ZN(n9694) );
  INV_X1 U11502 ( .A(n10144), .ZN(n9697) );
  NAND2_X1 U11503 ( .A1(n9697), .A2(n10168), .ZN(n15775) );
  INV_X1 U11504 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10131) );
  INV_X1 U11505 ( .A(n10132), .ZN(n9699) );
  AOI22_X1 U11506 ( .A1(n15775), .A2(n10131), .B1(n9702), .B2(n9699), .ZN(
        P1_U3445) );
  INV_X1 U11507 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10128) );
  OR2_X1 U11508 ( .A1(n15253), .A2(n9700), .ZN(n10129) );
  INV_X1 U11509 ( .A(n10129), .ZN(n9701) );
  AOI22_X1 U11510 ( .A1(n15775), .A2(n10128), .B1(n9702), .B2(n9701), .ZN(
        P1_U3446) );
  INV_X1 U11511 ( .A(n9703), .ZN(n9704) );
  OAI222_X1 U11512 ( .A1(P3_U3151), .A2(n13676), .B1(n13462), .B2(n10774), 
        .C1(n14119), .C2(n9704), .ZN(P3_U3279) );
  INV_X1 U11513 ( .A(n15813), .ZN(n15835) );
  AOI22_X1 U11514 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n15830), .B1(n15835), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n9708) );
  INV_X1 U11515 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9706) );
  OAI21_X1 U11516 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n15813), .A(n14306), .ZN(
        n9705) );
  AOI21_X1 U11517 ( .B1(n15830), .B2(n9706), .A(n9705), .ZN(n9707) );
  MUX2_X1 U11518 ( .A(n9708), .B(n9707), .S(P2_IR_REG_0__SCAN_IN), .Z(n9710)
         );
  AOI22_X1 U11519 ( .A1(n15800), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n9709) );
  NAND2_X1 U11520 ( .A1(n9710), .A2(n9709), .ZN(P2_U3214) );
  MUX2_X1 U11521 ( .A(n9714), .B(n9757), .S(n12298), .Z(n9715) );
  NAND2_X1 U11522 ( .A1(n9715), .A2(n15485), .ZN(n9770) );
  INV_X1 U11523 ( .A(n9715), .ZN(n9716) );
  NAND2_X1 U11524 ( .A1(n9716), .A2(SI_12_), .ZN(n9717) );
  INV_X1 U11525 ( .A(n11562), .ZN(n9756) );
  OAI21_X1 U11526 ( .B1(n9718), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9771) );
  XNOR2_X1 U11527 ( .A(n9771), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U11528 ( .A1(n11563), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n10530), .ZN(n9719) );
  OAI21_X1 U11529 ( .B1(n9756), .B2(n15260), .A(n9719), .ZN(P1_U3343) );
  NAND2_X1 U11530 ( .A1(n14265), .A2(n7431), .ZN(n9726) );
  INV_X1 U11531 ( .A(n9726), .ZN(n9728) );
  XNOR2_X1 U11532 ( .A(n14224), .B(n9823), .ZN(n9727) );
  NOR2_X1 U11533 ( .A1(n9725), .A2(n9724), .ZN(n14230) );
  XNOR2_X1 U11534 ( .A(n9727), .B(n9726), .ZN(n14229) );
  OAI21_X1 U11535 ( .B1(n14231), .B2(n14230), .A(n14229), .ZN(n14228) );
  OAI21_X1 U11536 ( .B1(n9728), .B2(n9727), .A(n14228), .ZN(n9740) );
  NAND2_X1 U11537 ( .A1(n10721), .A2(n7434), .ZN(n9731) );
  AOI22_X1 U11538 ( .A1(n7430), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n13109), 
        .B2(n9729), .ZN(n9730) );
  INV_X2 U11539 ( .A(n8716), .ZN(n11516) );
  XNOR2_X1 U11540 ( .A(n16169), .B(n11516), .ZN(n9738) );
  NAND2_X1 U11541 ( .A1(n9789), .A2(n9679), .ZN(n9736) );
  NAND2_X1 U11542 ( .A1(n9742), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9735) );
  NAND2_X1 U11543 ( .A1(n9732), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n9734) );
  NAND2_X1 U11544 ( .A1(n13368), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9733) );
  NAND4_X1 U11545 ( .A1(n9736), .A2(n9735), .A3(n9734), .A4(n9733), .ZN(n14264) );
  INV_X2 U11546 ( .A(n14147), .ZN(n14445) );
  AND2_X1 U11547 ( .A1(n14264), .A2(n14445), .ZN(n9737) );
  NAND2_X1 U11548 ( .A1(n9738), .A2(n9737), .ZN(n9781) );
  OAI21_X1 U11549 ( .B1(n9738), .B2(n9737), .A(n9781), .ZN(n9739) );
  AOI211_X1 U11550 ( .C1(n9740), .C2(n9739), .A(n14248), .B(n9783), .ZN(n9753)
         );
  NAND2_X1 U11551 ( .A1(n9742), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9748) );
  NOR2_X1 U11552 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9743) );
  NOR2_X1 U11553 ( .A1(n9790), .A2(n9743), .ZN(n9788) );
  NAND2_X1 U11554 ( .A1(n11931), .A2(n9788), .ZN(n9747) );
  NAND2_X1 U11555 ( .A1(n9732), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9746) );
  NAND2_X1 U11556 ( .A1(n9744), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9745) );
  AOI22_X1 U11557 ( .A1(n14227), .A2(n14265), .B1(n14225), .B2(n14263), .ZN(
        n9751) );
  AOI21_X1 U11558 ( .B1(n14246), .B2(n16169), .A(n9749), .ZN(n9750) );
  OAI211_X1 U11559 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n14218), .A(n9751), .B(
        n9750), .ZN(n9752) );
  OR2_X1 U11560 ( .A1(n9753), .A2(n9752), .ZN(P2_U3190) );
  OR2_X1 U11561 ( .A1(n9754), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n9776) );
  NAND2_X1 U11562 ( .A1(n9776), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9755) );
  XNOR2_X1 U11563 ( .A(n9755), .B(P2_IR_REG_12__SCAN_IN), .ZN(n11431) );
  INV_X1 U11564 ( .A(n11431), .ZN(n11075) );
  OAI222_X1 U11565 ( .A1(n14693), .A2(n9757), .B1(n14691), .B2(n9756), .C1(
        n11075), .C2(P2_U3088), .ZN(P2_U3315) );
  AOI21_X1 U11566 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n10022), .A(n9758), .ZN(
        n9760) );
  XNOR2_X1 U11567 ( .A(n10397), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n9759) );
  NOR2_X1 U11568 ( .A1(n9760), .A2(n9759), .ZN(n10183) );
  AOI211_X1 U11569 ( .C1(n9760), .C2(n9759), .A(n15817), .B(n10183), .ZN(n9768) );
  INV_X1 U11570 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9762) );
  MUX2_X1 U11571 ( .A(n9762), .B(P2_REG1_REG_7__SCAN_IN), .S(n10397), .Z(n9763) );
  NOR2_X1 U11572 ( .A1(n9764), .A2(n9763), .ZN(n10192) );
  AOI211_X1 U11573 ( .C1(n9764), .C2(n9763), .A(n15813), .B(n10192), .ZN(n9767) );
  INV_X1 U11574 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n15737) );
  NAND2_X1 U11575 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n10411) );
  NAND2_X1 U11576 ( .A1(n15838), .A2(n10397), .ZN(n9765) );
  OAI211_X1 U11577 ( .C1(n15844), .C2(n15737), .A(n10411), .B(n9765), .ZN(
        n9766) );
  OR3_X1 U11578 ( .A1(n9768), .A2(n9767), .A3(n9766), .ZN(P2_U3221) );
  MUX2_X1 U11579 ( .A(n9775), .B(n9780), .S(n12298), .Z(n9868) );
  XNOR2_X1 U11580 ( .A(n9868), .B(SI_13_), .ZN(n9865) );
  INV_X1 U11581 ( .A(n11780), .ZN(n9779) );
  NAND2_X1 U11582 ( .A1(n9771), .A2(n15639), .ZN(n9772) );
  NAND2_X1 U11583 ( .A1(n9772), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9773) );
  INV_X1 U11584 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n15646) );
  NAND2_X1 U11585 ( .A1(n9773), .A2(n15646), .ZN(n9875) );
  OR2_X1 U11586 ( .A1(n9773), .A2(n15646), .ZN(n9774) );
  INV_X1 U11587 ( .A(n11781), .ZN(n11185) );
  OAI222_X1 U11588 ( .A1(n15262), .A2(n9775), .B1(n15260), .B2(n9779), .C1(
        n11185), .C2(P1_U3086), .ZN(P1_U3342) );
  NOR2_X1 U11589 ( .A1(n9776), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n9879) );
  OR2_X1 U11590 ( .A1(n9879), .A2(n14676), .ZN(n9777) );
  XNOR2_X1 U11591 ( .A(n9777), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11691) );
  INV_X1 U11592 ( .A(n11691), .ZN(n9778) );
  OAI222_X1 U11593 ( .A1(n14693), .A2(n9780), .B1(n14691), .B2(n9779), .C1(
        n9778), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U11594 ( .A(n9781), .ZN(n9782) );
  NAND2_X1 U11595 ( .A1(n10865), .A2(n9720), .ZN(n9786) );
  AOI22_X1 U11596 ( .A1(n9659), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n13109), 
        .B2(n9784), .ZN(n9785) );
  XNOR2_X1 U11597 ( .A(n13146), .B(n11516), .ZN(n9820) );
  NAND2_X1 U11598 ( .A1(n14263), .A2(n7431), .ZN(n9821) );
  XNOR2_X1 U11599 ( .A(n9820), .B(n9821), .ZN(n9787) );
  OAI21_X1 U11600 ( .B1(n7605), .B2(n9787), .A(n9826), .ZN(n9799) );
  INV_X1 U11601 ( .A(n9788), .ZN(n10419) );
  NAND2_X1 U11602 ( .A1(n9742), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9795) );
  NOR2_X1 U11603 ( .A1(n9790), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9791) );
  NOR2_X1 U11604 ( .A1(n9828), .A2(n9791), .ZN(n10600) );
  NAND2_X1 U11605 ( .A1(n11931), .A2(n10600), .ZN(n9794) );
  NAND2_X1 U11606 ( .A1(n13386), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9793) );
  NAND2_X1 U11607 ( .A1(n13368), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9792) );
  NAND4_X1 U11608 ( .A1(n9795), .A2(n9794), .A3(n9793), .A4(n9792), .ZN(n14262) );
  INV_X1 U11609 ( .A(n14262), .ZN(n13157) );
  OAI22_X1 U11610 ( .A1(n8013), .A2(n14521), .B1(n13157), .B2(n14523), .ZN(
        n9910) );
  AOI22_X1 U11611 ( .A1(n14195), .A2(n9910), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3088), .ZN(n9797) );
  NAND2_X1 U11612 ( .A1(n14246), .A2(n13146), .ZN(n9796) );
  OAI211_X1 U11613 ( .C1(n14218), .C2(n10419), .A(n9797), .B(n9796), .ZN(n9798) );
  AOI21_X1 U11614 ( .B1(n9799), .B2(n14232), .A(n9798), .ZN(n9800) );
  INV_X1 U11615 ( .A(n9800), .ZN(P2_U3202) );
  INV_X1 U11616 ( .A(n15784), .ZN(n15781) );
  OR2_X1 U11617 ( .A1(n9801), .A2(n15781), .ZN(n15776) );
  NAND3_X1 U11618 ( .A1(n9803), .A2(n9802), .A3(n10200), .ZN(n9804) );
  NOR2_X1 U11619 ( .A1(n15776), .A2(n9804), .ZN(n9897) );
  INV_X1 U11620 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9813) );
  XNOR2_X1 U11621 ( .A(n14268), .B(n9890), .ZN(n13422) );
  XNOR2_X1 U11622 ( .A(n13116), .B(n13090), .ZN(n9805) );
  NAND2_X1 U11623 ( .A1(n13090), .A2(n14301), .ZN(n9807) );
  NAND2_X1 U11624 ( .A1(n13421), .A2(n13350), .ZN(n9806) );
  NOR2_X1 U11625 ( .A1(n14520), .A2(n14529), .ZN(n9808) );
  INV_X1 U11626 ( .A(n14266), .ZN(n10664) );
  OAI22_X1 U11627 ( .A1(n13422), .A2(n9808), .B1(n10664), .B2(n14523), .ZN(
        n10207) );
  INV_X1 U11628 ( .A(n9809), .ZN(n9810) );
  NOR2_X1 U11629 ( .A1(n9810), .A2(n13121), .ZN(n9811) );
  NOR2_X1 U11630 ( .A1(n10207), .A2(n9811), .ZN(n10205) );
  OAI21_X1 U11631 ( .B1(n13422), .B2(n9885), .A(n10205), .ZN(n14637) );
  NAND2_X1 U11632 ( .A1(n14668), .A2(n14637), .ZN(n9812) );
  OAI21_X1 U11633 ( .B1(n14668), .B2(n9813), .A(n9812), .ZN(P2_U3430) );
  INV_X1 U11634 ( .A(n9814), .ZN(n9815) );
  OAI222_X1 U11635 ( .A1(P3_U3151), .A2(n13719), .B1(n13462), .B2(n11001), 
        .C1(n14119), .C2(n9815), .ZN(P3_U3277) );
  INV_X1 U11636 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n15389) );
  NAND2_X1 U11637 ( .A1(n13944), .A2(P3_U3897), .ZN(n9816) );
  OAI21_X1 U11638 ( .B1(P3_U3897), .B2(n15389), .A(n9816), .ZN(P3_U3506) );
  NAND2_X1 U11639 ( .A1(n10869), .A2(n9720), .ZN(n9819) );
  AOI22_X1 U11640 ( .A1(n9659), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n13109), 
        .B2(n9817), .ZN(n9818) );
  NAND2_X1 U11641 ( .A1(n9819), .A2(n9818), .ZN(n13155) );
  INV_X1 U11642 ( .A(n13155), .ZN(n10603) );
  INV_X1 U11643 ( .A(n9820), .ZN(n9822) );
  NAND2_X1 U11644 ( .A1(n9822), .A2(n9821), .ZN(n9824) );
  NAND2_X1 U11645 ( .A1(n14262), .A2(n7431), .ZN(n10020) );
  XNOR2_X1 U11646 ( .A(n13155), .B(n9823), .ZN(n10019) );
  XOR2_X1 U11647 ( .A(n10020), .B(n10019), .Z(n9825) );
  AND3_X1 U11648 ( .A1(n9826), .A2(n9825), .A3(n9824), .ZN(n9827) );
  NAND2_X1 U11649 ( .A1(n9828), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10030) );
  OAI21_X1 U11650 ( .B1(n9828), .B2(P2_REG3_REG_6__SCAN_IN), .A(n10030), .ZN(
        n10039) );
  INV_X1 U11651 ( .A(n10039), .ZN(n16222) );
  NAND2_X1 U11652 ( .A1(n11931), .A2(n16222), .ZN(n9833) );
  NAND2_X1 U11653 ( .A1(n9742), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9832) );
  NAND2_X1 U11654 ( .A1(n13386), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n9831) );
  INV_X2 U11655 ( .A(n9829), .ZN(n13368) );
  NAND2_X1 U11656 ( .A1(n13368), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9830) );
  NAND4_X1 U11657 ( .A1(n9833), .A2(n9832), .A3(n9831), .A4(n9830), .ZN(n14261) );
  INV_X1 U11658 ( .A(n14263), .ZN(n10218) );
  INV_X1 U11659 ( .A(n10600), .ZN(n9834) );
  OAI22_X1 U11660 ( .A1(n14219), .A2(n10218), .B1(n9834), .B2(n14218), .ZN(
        n9835) );
  AOI211_X1 U11661 ( .C1(n14225), .C2(n14261), .A(n9836), .B(n9835), .ZN(n9837) );
  OAI211_X1 U11662 ( .C1(n10603), .C2(n12244), .A(n9838), .B(n9837), .ZN(
        P2_U3199) );
  INV_X1 U11663 ( .A(n10168), .ZN(n9839) );
  NAND2_X1 U11664 ( .A1(n10175), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12774) );
  NAND2_X1 U11665 ( .A1(n9839), .A2(n12774), .ZN(n9856) );
  NAND2_X1 U11666 ( .A1(n9348), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9840) );
  INV_X1 U11667 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9841) );
  NAND3_X1 U11668 ( .A1(n9347), .A2(n15658), .A3(n9841), .ZN(n9842) );
  OAI21_X1 U11669 ( .B1(n10821), .B2(n9842), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9843) );
  NAND2_X1 U11670 ( .A1(n12540), .A2(n15263), .ZN(n12716) );
  OR2_X1 U11671 ( .A1(n12716), .A2(n10175), .ZN(n9853) );
  NAND3_X1 U11672 ( .A1(n9845), .A2(n9844), .A3(n15649), .ZN(n9850) );
  NOR2_X1 U11673 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), 
        .ZN(n9849) );
  NOR2_X1 U11674 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .ZN(n9848) );
  NOR2_X1 U11675 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n9847) );
  NOR2_X1 U11676 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n9846) );
  NAND2_X1 U11677 ( .A1(n9853), .A2(n12316), .ZN(n9854) );
  NAND2_X1 U11678 ( .A1(n9856), .A2(n9854), .ZN(n16028) );
  INV_X1 U11679 ( .A(n16028), .ZN(n14866) );
  INV_X1 U11680 ( .A(n9854), .ZN(n9855) );
  NAND2_X1 U11681 ( .A1(n9856), .A2(n9855), .ZN(n9923) );
  NOR2_X1 U11682 ( .A1(n13078), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9857) );
  OR2_X1 U11683 ( .A1(n9857), .A2(n15245), .ZN(n10358) );
  INV_X1 U11684 ( .A(n10358), .ZN(n9859) );
  INV_X1 U11685 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n16035) );
  NAND2_X1 U11686 ( .A1(n13078), .A2(n16035), .ZN(n9858) );
  NAND2_X1 U11687 ( .A1(n9859), .A2(n9858), .ZN(n9860) );
  MUX2_X1 U11688 ( .A(n9860), .B(n9859), .S(P1_IR_REG_0__SCAN_IN), .Z(n9861)
         );
  INV_X1 U11689 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n16043) );
  OAI22_X1 U11690 ( .A1(n9923), .A2(n9861), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n16043), .ZN(n9862) );
  AOI21_X1 U11691 ( .B1(n14866), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n9862), .ZN(
        n9864) );
  INV_X1 U11692 ( .A(n13078), .ZN(n12781) );
  INV_X1 U11693 ( .A(n15852), .ZN(n16018) );
  NAND3_X1 U11694 ( .A1(n16018), .A2(P1_IR_REG_0__SCAN_IN), .A3(n16035), .ZN(
        n9863) );
  NAND2_X1 U11695 ( .A1(n9864), .A2(n9863), .ZN(P1_U3243) );
  INV_X1 U11696 ( .A(n9865), .ZN(n9866) );
  INV_X1 U11697 ( .A(n9868), .ZN(n9869) );
  NAND2_X1 U11698 ( .A1(n9869), .A2(SI_13_), .ZN(n9870) );
  MUX2_X1 U11699 ( .A(n9877), .B(n9882), .S(n12298), .Z(n9872) );
  INV_X1 U11700 ( .A(n9872), .ZN(n9873) );
  NAND2_X1 U11701 ( .A1(n9873), .A2(SI_14_), .ZN(n9874) );
  NAND2_X1 U11702 ( .A1(n10243), .A2(n9874), .ZN(n10241) );
  XNOR2_X1 U11703 ( .A(n10242), .B(n10241), .ZN(n12002) );
  INV_X1 U11704 ( .A(n12002), .ZN(n9881) );
  NAND2_X1 U11705 ( .A1(n9875), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9876) );
  INV_X1 U11706 ( .A(n14901), .ZN(n11188) );
  OAI222_X1 U11707 ( .A1(n15262), .A2(n9877), .B1(n15260), .B2(n9881), .C1(
        P1_U3086), .C2(n11188), .ZN(P1_U3341) );
  INV_X1 U11708 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n9878) );
  NAND2_X1 U11709 ( .A1(n9879), .A2(n9878), .ZN(n10251) );
  NAND2_X1 U11710 ( .A1(n10251), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9880) );
  XNOR2_X1 U11711 ( .A(n9880), .B(P2_IR_REG_14__SCAN_IN), .ZN(n12221) );
  INV_X1 U11712 ( .A(n12221), .ZN(n11639) );
  OAI222_X1 U11713 ( .A1(n14693), .A2(n9882), .B1(n14691), .B2(n9881), .C1(
        P2_U3088), .C2(n11639), .ZN(P2_U3313) );
  INV_X1 U11714 ( .A(n9883), .ZN(n9884) );
  OAI222_X1 U11715 ( .A1(P3_U3151), .A2(n13733), .B1(n14119), .B2(n9884), .C1(
        n15473), .C2(n13462), .ZN(P3_U3276) );
  INV_X1 U11716 ( .A(n7424), .ZN(n9887) );
  INV_X1 U11717 ( .A(n9889), .ZN(n9886) );
  NAND2_X1 U11718 ( .A1(n9887), .A2(n9886), .ZN(n9900) );
  INV_X1 U11719 ( .A(n9900), .ZN(n9888) );
  AOI21_X1 U11720 ( .B1(n9889), .B2(n7424), .A(n9888), .ZN(n9895) );
  INV_X1 U11721 ( .A(n9895), .ZN(n14545) );
  AOI211_X1 U11722 ( .C1(n9890), .C2(n14547), .A(n7431), .B(n10666), .ZN(
        n14546) );
  INV_X1 U11723 ( .A(n14520), .ZN(n12045) );
  AOI22_X1 U11724 ( .A1(n14438), .A2(n14268), .B1(n14265), .B2(n14439), .ZN(
        n9894) );
  NOR2_X1 U11725 ( .A1(n14268), .A2(n13121), .ZN(n9891) );
  OAI21_X1 U11726 ( .B1(n9891), .B2(n7424), .A(n10659), .ZN(n9892) );
  NAND2_X1 U11727 ( .A1(n9892), .A2(n14529), .ZN(n9893) );
  OAI211_X1 U11728 ( .C1(n9895), .C2(n12045), .A(n9894), .B(n9893), .ZN(n14548) );
  AOI211_X1 U11729 ( .C1(n13099), .C2(n14545), .A(n14546), .B(n14548), .ZN(
        n10286) );
  INV_X1 U11730 ( .A(n15783), .ZN(n9896) );
  INV_X1 U11731 ( .A(n14631), .ZN(n11917) );
  AOI22_X1 U11732 ( .A1(n11917), .A2(n14547), .B1(n16357), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n9898) );
  OAI21_X1 U11733 ( .B1(n10286), .B2(n16357), .A(n9898), .ZN(P2_U3500) );
  NAND2_X1 U11734 ( .A1(n10664), .A2(n10283), .ZN(n9899) );
  NAND2_X1 U11735 ( .A1(n9900), .A2(n9899), .ZN(n10657) );
  INV_X1 U11736 ( .A(n14265), .ZN(n9902) );
  NAND2_X1 U11737 ( .A1(n9902), .A2(n14224), .ZN(n9906) );
  NAND2_X1 U11738 ( .A1(n14265), .A2(n16127), .ZN(n9901) );
  NAND2_X1 U11739 ( .A1(n9902), .A2(n16127), .ZN(n9903) );
  NAND2_X1 U11740 ( .A1(n8013), .A2(n10436), .ZN(n9904) );
  NAND2_X1 U11741 ( .A1(n9905), .A2(n13425), .ZN(n10211) );
  OAI21_X1 U11742 ( .B1(n9905), .B2(n13425), .A(n10211), .ZN(n10416) );
  NAND2_X1 U11743 ( .A1(n10666), .A2(n16127), .ZN(n10665) );
  OR2_X1 U11744 ( .A1(n10665), .A2(n16169), .ZN(n10434) );
  AOI211_X1 U11745 ( .C1(n13146), .C2(n10434), .A(n14445), .B(n10214), .ZN(
        n10422) );
  NAND2_X1 U11746 ( .A1(n10664), .A2(n14547), .ZN(n10658) );
  NAND2_X1 U11747 ( .A1(n8013), .A2(n16169), .ZN(n9907) );
  NAND2_X1 U11748 ( .A1(n10430), .A2(n9907), .ZN(n9909) );
  INV_X1 U11749 ( .A(n13425), .ZN(n9908) );
  OAI21_X1 U11750 ( .B1(n9909), .B2(n9908), .A(n10217), .ZN(n9911) );
  AOI21_X1 U11751 ( .B1(n9911), .B2(n14529), .A(n9910), .ZN(n10423) );
  INV_X1 U11752 ( .A(n10423), .ZN(n9912) );
  AOI211_X1 U11753 ( .C1(n16348), .C2(n10416), .A(n10422), .B(n9912), .ZN(
        n10240) );
  AOI22_X1 U11754 ( .A1(n11917), .A2(n13146), .B1(n16357), .B2(
        P2_REG1_REG_4__SCAN_IN), .ZN(n9913) );
  OAI21_X1 U11755 ( .B1(n10240), .B2(n16357), .A(n9913), .ZN(P2_U3503) );
  CLKBUF_X2 U11756 ( .A(P1_U4016), .Z(n14861) );
  NOR2_X1 U11757 ( .A1(n14866), .A2(n14861), .ZN(P1_U3085) );
  INV_X1 U11758 ( .A(n15245), .ZN(n10361) );
  INV_X1 U11759 ( .A(n10722), .ZN(n9932) );
  INV_X1 U11760 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10739) );
  OAI22_X1 U11761 ( .A1(n16028), .A2(n15674), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10739), .ZN(n9922) );
  INV_X1 U11762 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9914) );
  MUX2_X1 U11763 ( .A(n9914), .B(P1_REG1_REG_1__SCAN_IN), .S(n14867), .Z(n9916) );
  AND2_X1 U11764 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9915) );
  NAND2_X1 U11765 ( .A1(n9916), .A2(n9915), .ZN(n14870) );
  OR2_X1 U11766 ( .A1(n14867), .A2(n9914), .ZN(n9917) );
  NAND2_X1 U11767 ( .A1(n14870), .A2(n9917), .ZN(n10364) );
  XNOR2_X1 U11768 ( .A(n10103), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n10363) );
  INV_X1 U11769 ( .A(n10103), .ZN(n10371) );
  AOI22_X1 U11770 ( .A1(n10364), .A2(n10363), .B1(n10371), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n9920) );
  INV_X1 U11771 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n16150) );
  MUX2_X1 U11772 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n16150), .S(n10722), .Z(
        n9919) );
  OR2_X1 U11773 ( .A1(n9920), .A2(n9919), .ZN(n16015) );
  INV_X1 U11774 ( .A(n16015), .ZN(n9918) );
  AOI211_X1 U11775 ( .C1(n9920), .C2(n9919), .A(n9918), .B(n15852), .ZN(n9921)
         );
  AOI211_X1 U11776 ( .C1(n14900), .C2(n9932), .A(n9922), .B(n9921), .ZN(n9931)
         );
  NOR2_X1 U11777 ( .A1(n9923), .A2(n13078), .ZN(n12064) );
  INV_X1 U11778 ( .A(n12064), .ZN(n9924) );
  XNOR2_X1 U11779 ( .A(n14867), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n14865) );
  AND2_X1 U11780 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14864) );
  NAND2_X1 U11781 ( .A1(n14865), .A2(n14864), .ZN(n14863) );
  INV_X1 U11782 ( .A(n14867), .ZN(n14871) );
  NAND2_X1 U11783 ( .A1(n14871), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9925) );
  NAND2_X1 U11784 ( .A1(n14863), .A2(n9925), .ZN(n10366) );
  INV_X1 U11785 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n15094) );
  MUX2_X1 U11786 ( .A(n15094), .B(P1_REG2_REG_2__SCAN_IN), .S(n10103), .Z(
        n10367) );
  NAND2_X1 U11787 ( .A1(n10366), .A2(n10367), .ZN(n10365) );
  NAND2_X1 U11788 ( .A1(n10371), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9926) );
  INV_X1 U11789 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9939) );
  MUX2_X1 U11790 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9939), .S(n10722), .Z(n9927) );
  AOI21_X1 U11791 ( .B1(n10365), .B2(n9926), .A(n9927), .ZN(n16011) );
  INV_X1 U11792 ( .A(n16011), .ZN(n9929) );
  NAND3_X1 U11793 ( .A1(n10365), .A2(n9927), .A3(n9926), .ZN(n9928) );
  NAND3_X1 U11794 ( .A1(n7422), .A2(n9929), .A3(n9928), .ZN(n9930) );
  NAND2_X1 U11795 ( .A1(n9931), .A2(n9930), .ZN(P1_U3246) );
  INV_X1 U11796 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n16212) );
  MUX2_X1 U11797 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n16212), .S(n10870), .Z(
        n9934) );
  NAND2_X1 U11798 ( .A1(n9932), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n16014) );
  INV_X1 U11799 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n16196) );
  MUX2_X1 U11800 ( .A(n16196), .B(P1_REG1_REG_4__SCAN_IN), .S(n16003), .Z(
        n16013) );
  AOI21_X1 U11801 ( .B1(n16015), .B2(n16014), .A(n16013), .ZN(n16012) );
  AOI21_X1 U11802 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n16003), .A(n16012), .ZN(
        n9933) );
  NAND2_X1 U11803 ( .A1(n9933), .A2(n9934), .ZN(n9973) );
  OAI21_X1 U11804 ( .B1(n9934), .B2(n9933), .A(n9973), .ZN(n9938) );
  INV_X1 U11805 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9936) );
  NAND2_X1 U11806 ( .A1(n14900), .A2(n10870), .ZN(n9935) );
  NAND2_X1 U11807 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n11021) );
  OAI211_X1 U11808 ( .C1(n9936), .C2(n16028), .A(n9935), .B(n11021), .ZN(n9937) );
  AOI21_X1 U11809 ( .B1(n16018), .B2(n9938), .A(n9937), .ZN(n9946) );
  NOR2_X1 U11810 ( .A1(n10722), .A2(n9939), .ZN(n16005) );
  INV_X1 U11811 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n16004) );
  MUX2_X1 U11812 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n16004), .S(n16003), .Z(
        n9940) );
  OAI21_X1 U11813 ( .B1(n16011), .B2(n16005), .A(n9940), .ZN(n16008) );
  NAND2_X1 U11814 ( .A1(n16003), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9942) );
  INV_X1 U11815 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9963) );
  MUX2_X1 U11816 ( .A(n9963), .B(P1_REG2_REG_5__SCAN_IN), .S(n10870), .Z(n9941) );
  AOI21_X1 U11817 ( .B1(n16008), .B2(n9942), .A(n9941), .ZN(n10003) );
  INV_X1 U11818 ( .A(n10003), .ZN(n9944) );
  NAND3_X1 U11819 ( .A1(n16008), .A2(n9942), .A3(n9941), .ZN(n9943) );
  NAND3_X1 U11820 ( .A1(n7422), .A2(n9944), .A3(n9943), .ZN(n9945) );
  NAND2_X1 U11821 ( .A1(n9946), .A2(n9945), .ZN(P1_U3248) );
  OR2_X1 U11822 ( .A1(n10331), .A2(P3_U3151), .ZN(n13043) );
  INV_X1 U11823 ( .A(n13043), .ZN(n9947) );
  OR2_X1 U11824 ( .A1(n10349), .A2(n9947), .ZN(n9960) );
  NAND2_X1 U11825 ( .A1(n12974), .A2(n10331), .ZN(n9948) );
  NAND2_X1 U11826 ( .A1(n9949), .A2(n9948), .ZN(n9959) );
  INV_X1 U11827 ( .A(n9959), .ZN(n9950) );
  AND2_X1 U11828 ( .A1(n9960), .A2(n9950), .ZN(n9956) );
  INV_X1 U11829 ( .A(n9956), .ZN(n9952) );
  MUX2_X1 U11830 ( .A(n9952), .B(n13623), .S(n9951), .Z(n15984) );
  AND2_X1 U11831 ( .A1(n9953), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10316) );
  NOR2_X1 U11832 ( .A1(n9953), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9958) );
  INV_X1 U11833 ( .A(n9954), .ZN(n9955) );
  INV_X1 U11834 ( .A(n15966), .ZN(n15999) );
  NAND2_X1 U11835 ( .A1(P3_U3897), .A2(n13037), .ZN(n15991) );
  NAND3_X1 U11836 ( .A1(n15999), .A2(n15993), .A3(n15991), .ZN(n9957) );
  OAI21_X1 U11837 ( .B1(n10316), .B2(n9958), .A(n9957), .ZN(n9962) );
  AOI22_X1 U11838 ( .A1(n15961), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n9961) );
  OAI211_X1 U11839 ( .C1(n15984), .C2(n8391), .A(n9962), .B(n9961), .ZN(
        P3_U3182) );
  NOR2_X1 U11840 ( .A1(n9964), .A2(n9963), .ZN(n9999) );
  MUX2_X1 U11841 ( .A(n9998), .B(P1_REG2_REG_6__SCAN_IN), .S(n10011), .Z(n9965) );
  OAI21_X1 U11842 ( .B1(n10003), .B2(n9999), .A(n9965), .ZN(n14878) );
  INV_X1 U11843 ( .A(n10011), .ZN(n10880) );
  NAND2_X1 U11844 ( .A1(n10880), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n14877) );
  INV_X1 U11845 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9966) );
  MUX2_X1 U11846 ( .A(n9966), .B(P1_REG2_REG_7__SCAN_IN), .S(n14883), .Z(
        n14876) );
  AOI21_X1 U11847 ( .B1(n14878), .B2(n14877), .A(n14876), .ZN(n9989) );
  NOR2_X1 U11848 ( .A1(n9975), .A2(n9966), .ZN(n9990) );
  INV_X1 U11849 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9967) );
  MUX2_X1 U11850 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n9967), .S(n11357), .Z(n9968) );
  OAI21_X1 U11851 ( .B1(n9989), .B2(n9990), .A(n9968), .ZN(n9994) );
  NAND2_X1 U11852 ( .A1(n11357), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9971) );
  INV_X1 U11853 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9969) );
  MUX2_X1 U11854 ( .A(n9969), .B(P1_REG2_REG_9__SCAN_IN), .S(n11363), .Z(n9970) );
  AOI21_X1 U11855 ( .B1(n9994), .B2(n9971), .A(n9970), .ZN(n10044) );
  NAND3_X1 U11856 ( .A1(n9994), .A2(n9971), .A3(n9970), .ZN(n9972) );
  NAND2_X1 U11857 ( .A1(n7422), .A2(n9972), .ZN(n9984) );
  INV_X1 U11858 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n14884) );
  OAI21_X1 U11859 ( .B1(n10870), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9973), .ZN(
        n10004) );
  INV_X1 U11860 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10910) );
  MUX2_X1 U11861 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10910), .S(n10011), .Z(
        n10005) );
  NOR2_X1 U11862 ( .A1(n10004), .A2(n10005), .ZN(n14890) );
  AND2_X1 U11863 ( .A1(n10880), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n14885) );
  MUX2_X1 U11864 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n14884), .S(n14883), .Z(
        n9974) );
  OAI21_X1 U11865 ( .B1(n14890), .B2(n14885), .A(n9974), .ZN(n14888) );
  OAI21_X1 U11866 ( .B1(n14884), .B2(n9975), .A(n14888), .ZN(n9986) );
  INV_X1 U11867 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9976) );
  MUX2_X1 U11868 ( .A(n9976), .B(P1_REG1_REG_8__SCAN_IN), .S(n11357), .Z(n9987) );
  NOR2_X1 U11869 ( .A1(n9986), .A2(n9987), .ZN(n9985) );
  NOR2_X1 U11870 ( .A1(n11357), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9977) );
  INV_X1 U11871 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n16286) );
  MUX2_X1 U11872 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n16286), .S(n11363), .Z(
        n9978) );
  OAI21_X1 U11873 ( .B1(n9985), .B2(n9977), .A(n9978), .ZN(n10050) );
  INV_X1 U11874 ( .A(n10050), .ZN(n9980) );
  NOR3_X1 U11875 ( .A1(n9985), .A2(n9978), .A3(n9977), .ZN(n9979) );
  OAI21_X1 U11876 ( .B1(n9980), .B2(n9979), .A(n16018), .ZN(n9983) );
  INV_X1 U11877 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n15706) );
  NAND2_X1 U11878 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n11874) );
  OAI21_X1 U11879 ( .B1(n16028), .B2(n15706), .A(n11874), .ZN(n9981) );
  AOI21_X1 U11880 ( .B1(n11363), .B2(n14900), .A(n9981), .ZN(n9982) );
  OAI211_X1 U11881 ( .C1(n10044), .C2(n9984), .A(n9983), .B(n9982), .ZN(
        P1_U3252) );
  AOI21_X1 U11882 ( .B1(n9987), .B2(n9986), .A(n9985), .ZN(n9997) );
  NAND2_X1 U11883 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11493) );
  OAI21_X1 U11884 ( .B1(n16028), .B2(n15686), .A(n11493), .ZN(n9988) );
  AOI21_X1 U11885 ( .B1(n11357), .B2(n14900), .A(n9988), .ZN(n9996) );
  INV_X1 U11886 ( .A(n9989), .ZN(n14880) );
  INV_X1 U11887 ( .A(n9990), .ZN(n9992) );
  MUX2_X1 U11888 ( .A(n9967), .B(P1_REG2_REG_8__SCAN_IN), .S(n11357), .Z(n9991) );
  NAND3_X1 U11889 ( .A1(n14880), .A2(n9992), .A3(n9991), .ZN(n9993) );
  NAND3_X1 U11890 ( .A1(n7422), .A2(n9994), .A3(n9993), .ZN(n9995) );
  OAI211_X1 U11891 ( .C1(n9997), .C2(n15852), .A(n9996), .B(n9995), .ZN(
        P1_U3251) );
  INV_X1 U11892 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9998) );
  MUX2_X1 U11893 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9998), .S(n10011), .Z(
        n10001) );
  INV_X1 U11894 ( .A(n9999), .ZN(n10000) );
  NAND2_X1 U11895 ( .A1(n10001), .A2(n10000), .ZN(n10002) );
  OAI211_X1 U11896 ( .C1(n10003), .C2(n10002), .A(n7422), .B(n14878), .ZN(
        n10010) );
  NAND2_X1 U11897 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n11178) );
  AOI211_X1 U11898 ( .C1(n10005), .C2(n10004), .A(n14890), .B(n15852), .ZN(
        n10006) );
  INV_X1 U11899 ( .A(n10006), .ZN(n10007) );
  NAND2_X1 U11900 ( .A1(n11178), .A2(n10007), .ZN(n10008) );
  AOI21_X1 U11901 ( .B1(n14866), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10008), .ZN(
        n10009) );
  OAI211_X1 U11902 ( .C1(n16022), .C2(n10011), .A(n10010), .B(n10009), .ZN(
        P1_U3249) );
  INV_X1 U11903 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n12982) );
  NOR2_X2 U11904 ( .A1(n10015), .A2(n15238), .ZN(n10081) );
  INV_X1 U11905 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n14912) );
  INV_X2 U11906 ( .A(n12018), .ZN(n12524) );
  NAND2_X1 U11907 ( .A1(n12524), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n10017) );
  NAND2_X1 U11908 ( .A1(n12686), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n10016) );
  OAI211_X1 U11909 ( .C1(n12431), .C2(n14912), .A(n10017), .B(n10016), .ZN(
        n14914) );
  NAND2_X1 U11910 ( .A1(n14861), .A2(n14914), .ZN(n10018) );
  OAI21_X1 U11911 ( .B1(n14861), .B2(n12982), .A(n10018), .ZN(P1_U3591) );
  INV_X1 U11912 ( .A(n10019), .ZN(n10021) );
  NAND2_X1 U11913 ( .A1(n10879), .A2(n9720), .ZN(n10024) );
  AOI22_X1 U11914 ( .A1(n9659), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n13109), 
        .B2(n10022), .ZN(n10023) );
  XNOR2_X1 U11915 ( .A(n16223), .B(n8716), .ZN(n10026) );
  NAND2_X1 U11916 ( .A1(n14261), .A2(n7431), .ZN(n10025) );
  NOR2_X1 U11917 ( .A1(n10026), .A2(n10025), .ZN(n10400) );
  AOI21_X1 U11918 ( .B1(n10026), .B2(n10025), .A(n10400), .ZN(n10027) );
  OAI211_X1 U11919 ( .C1(n10028), .C2(n10027), .A(n10402), .B(n14232), .ZN(
        n10042) );
  NAND2_X1 U11920 ( .A1(n9742), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10035) );
  AND2_X1 U11921 ( .A1(n10030), .A2(n10029), .ZN(n10031) );
  NOR2_X1 U11922 ( .A1(n10405), .A2(n10031), .ZN(n16248) );
  NAND2_X1 U11923 ( .A1(n11931), .A2(n16248), .ZN(n10034) );
  NAND2_X1 U11924 ( .A1(n13386), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n10033) );
  NAND2_X1 U11925 ( .A1(n13368), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10032) );
  NAND4_X1 U11926 ( .A1(n10035), .A2(n10034), .A3(n10033), .A4(n10032), .ZN(
        n14260) );
  NAND2_X1 U11927 ( .A1(n14260), .A2(n14439), .ZN(n10037) );
  NAND2_X1 U11928 ( .A1(n14262), .A2(n14438), .ZN(n10036) );
  NAND2_X1 U11929 ( .A1(n10037), .A2(n10036), .ZN(n10590) );
  AOI22_X1 U11930 ( .A1(n14195), .A2(n10590), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10038) );
  OAI21_X1 U11931 ( .B1(n10039), .B2(n14218), .A(n10038), .ZN(n10040) );
  AOI21_X1 U11932 ( .B1(n16223), .B2(n14246), .A(n10040), .ZN(n10041) );
  NAND2_X1 U11933 ( .A1(n10042), .A2(n10041), .ZN(P2_U3211) );
  INV_X1 U11934 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10043) );
  MUX2_X1 U11935 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n10043), .S(n11563), .Z(
        n10048) );
  AOI21_X1 U11936 ( .B1(n11363), .B2(P1_REG2_REG_9__SCAN_IN), .A(n10044), .ZN(
        n10445) );
  INV_X1 U11937 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10045) );
  MUX2_X1 U11938 ( .A(n10045), .B(P1_REG2_REG_10__SCAN_IN), .S(n11546), .Z(
        n10444) );
  OR2_X1 U11939 ( .A1(n10445), .A2(n10444), .ZN(n10446) );
  NAND2_X1 U11940 ( .A1(n11546), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10380) );
  INV_X1 U11941 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10046) );
  MUX2_X1 U11942 ( .A(n10046), .B(P1_REG2_REG_11__SCAN_IN), .S(n11551), .Z(
        n10379) );
  AOI21_X1 U11943 ( .B1(n10446), .B2(n10380), .A(n10379), .ZN(n10382) );
  AOI21_X1 U11944 ( .B1(n11551), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10382), 
        .ZN(n10047) );
  NAND2_X1 U11945 ( .A1(n10047), .A2(n10048), .ZN(n10390) );
  OAI21_X1 U11946 ( .B1(n10048), .B2(n10047), .A(n10390), .ZN(n10057) );
  INV_X1 U11947 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n15695) );
  NAND2_X1 U11948 ( .A1(n14900), .A2(n11563), .ZN(n10049) );
  NAND2_X1 U11949 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n12127)
         );
  OAI211_X1 U11950 ( .C1(n15695), .C2(n16028), .A(n10049), .B(n12127), .ZN(
        n10056) );
  INV_X1 U11951 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n11610) );
  OAI21_X1 U11952 ( .B1(n11363), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10050), .ZN(
        n10441) );
  MUX2_X1 U11953 ( .A(n11610), .B(P1_REG1_REG_10__SCAN_IN), .S(n11546), .Z(
        n10440) );
  OR2_X1 U11954 ( .A1(n10441), .A2(n10440), .ZN(n10442) );
  OAI21_X1 U11955 ( .B1(n11610), .B2(n10452), .A(n10442), .ZN(n10377) );
  INV_X1 U11956 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10051) );
  MUX2_X1 U11957 ( .A(n10051), .B(P1_REG1_REG_11__SCAN_IN), .S(n11551), .Z(
        n10378) );
  NOR2_X1 U11958 ( .A1(n10377), .A2(n10378), .ZN(n10376) );
  NOR2_X1 U11959 ( .A1(n11551), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10052) );
  INV_X1 U11960 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n16373) );
  MUX2_X1 U11961 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n16373), .S(n11563), .Z(
        n10053) );
  OAI21_X1 U11962 ( .B1(n10376), .B2(n10052), .A(n10053), .ZN(n10387) );
  OR3_X1 U11963 ( .A1(n10376), .A2(n10053), .A3(n10052), .ZN(n10054) );
  AOI21_X1 U11964 ( .B1(n10387), .B2(n10054), .A(n15852), .ZN(n10055) );
  AOI211_X1 U11965 ( .C1(n7422), .C2(n10057), .A(n10056), .B(n10055), .ZN(
        n10058) );
  INV_X1 U11966 ( .A(n10058), .ZN(P1_U3255) );
  XNOR2_X1 U11967 ( .A(n10076), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n10063) );
  NAND2_X1 U11968 ( .A1(n8391), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10059) );
  NAND2_X1 U11969 ( .A1(n10327), .A2(n10059), .ZN(n10060) );
  NAND2_X1 U11970 ( .A1(n10060), .A2(n10061), .ZN(n10322) );
  NAND2_X1 U11971 ( .A1(n10324), .A2(n10061), .ZN(n10062) );
  NAND2_X1 U11972 ( .A1(n10063), .A2(n10062), .ZN(n10263) );
  OAI21_X1 U11973 ( .B1(n10063), .B2(n10062), .A(n10263), .ZN(n10073) );
  XNOR2_X1 U11974 ( .A(n10076), .B(P3_REG1_REG_2__SCAN_IN), .ZN(n10068) );
  NAND2_X1 U11975 ( .A1(n8391), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10064) );
  NAND2_X1 U11976 ( .A1(n10065), .A2(n10066), .ZN(n10319) );
  NAND2_X1 U11977 ( .A1(n10317), .A2(n10066), .ZN(n10067) );
  NAND2_X1 U11978 ( .A1(n10068), .A2(n10067), .ZN(n10270) );
  OAI21_X1 U11979 ( .B1(n10068), .B2(n10067), .A(n10270), .ZN(n10069) );
  AND2_X1 U11980 ( .A1(n15931), .A2(n10069), .ZN(n10072) );
  INV_X1 U11981 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10070) );
  OAI22_X1 U11982 ( .A1(n15982), .A2(n10070), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n16114), .ZN(n10071) );
  AOI211_X1 U11983 ( .C1(n15966), .C2(n10073), .A(n10072), .B(n10071), .ZN(
        n10079) );
  XNOR2_X1 U11984 ( .A(n10074), .B(n8065), .ZN(n10315) );
  INV_X1 U11985 ( .A(n10074), .ZN(n10075) );
  AOI22_X1 U11986 ( .A1(n10315), .A2(n10316), .B1(n8065), .B2(n10075), .ZN(
        n10261) );
  XOR2_X1 U11987 ( .A(n10076), .B(n10259), .Z(n10260) );
  XNOR2_X1 U11988 ( .A(n10261), .B(n10260), .ZN(n10077) );
  NAND2_X1 U11989 ( .A1(n10077), .A2(n15970), .ZN(n10078) );
  OAI211_X1 U11990 ( .C1(n15984), .C2(n10268), .A(n10079), .B(n10078), .ZN(
        P3_U3184) );
  NAND2_X1 U11991 ( .A1(n12526), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n10086) );
  NAND2_X1 U11992 ( .A1(n7425), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10085) );
  NAND2_X1 U11993 ( .A1(n10114), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n10083) );
  NAND2_X1 U11994 ( .A1(n10089), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10082) );
  NAND2_X1 U11995 ( .A1(n7426), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10093) );
  NAND2_X1 U11996 ( .A1(n10089), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10092) );
  NAND2_X1 U11997 ( .A1(n10114), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n10090) );
  INV_X1 U11998 ( .A(SI_0_), .ZN(n10094) );
  NOR2_X1 U11999 ( .A1(n10095), .A2(n10094), .ZN(n10096) );
  XNOR2_X1 U12000 ( .A(n10096), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n15265) );
  MUX2_X1 U12001 ( .A(n8323), .B(n15265), .S(n12316), .Z(n16031) );
  NAND2_X1 U12002 ( .A1(n16073), .A2(n12546), .ZN(n10097) );
  NAND2_X1 U12003 ( .A1(n12526), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n10100) );
  NAND2_X1 U12004 ( .A1(n10114), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n10099) );
  NAND2_X1 U12005 ( .A1(n7427), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n10098) );
  XNOR2_X1 U12006 ( .A(n10891), .B(n12725), .ZN(n15089) );
  NAND2_X1 U12007 ( .A1(n10108), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10105) );
  MUX2_X1 U12008 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10105), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n10106) );
  INV_X1 U12009 ( .A(n16039), .ZN(n10165) );
  NAND2_X1 U12010 ( .A1(n12540), .A2(n10165), .ZN(n10111) );
  NAND2_X1 U12011 ( .A1(n10821), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10107) );
  MUX2_X1 U12012 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10107), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n10109) );
  NAND2_X1 U12013 ( .A1(n16038), .A2(n15263), .ZN(n10110) );
  NOR2_X1 U12014 ( .A1(n12540), .A2(n15263), .ZN(n16029) );
  NAND2_X1 U12015 ( .A1(n16039), .A2(n12752), .ZN(n10153) );
  NAND2_X1 U12016 ( .A1(n16039), .A2(n12784), .ZN(n12715) );
  INV_X1 U12017 ( .A(n12715), .ZN(n10112) );
  INV_X1 U12018 ( .A(n16144), .ZN(n10113) );
  AOI211_X1 U12019 ( .C1(n15095), .C2(n16077), .A(n16142), .B(n10113), .ZN(
        n15096) );
  INV_X1 U12020 ( .A(n15096), .ZN(n10121) );
  NAND2_X1 U12021 ( .A1(n7427), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n10118) );
  NAND2_X1 U12022 ( .A1(n10089), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10117) );
  NAND2_X1 U12023 ( .A1(n12526), .A2(n10739), .ZN(n10116) );
  NAND2_X1 U12024 ( .A1(n10114), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n10115) );
  NOR2_X1 U12025 ( .A1(n12716), .A2(n10361), .ZN(n14799) );
  NAND2_X1 U12026 ( .A1(n14858), .A2(n14799), .ZN(n10120) );
  NAND2_X1 U12027 ( .A1(n10151), .A2(n10361), .ZN(n14785) );
  NAND2_X1 U12028 ( .A1(n14860), .A2(n14806), .ZN(n10119) );
  AND2_X1 U12029 ( .A1(n10120), .A2(n10119), .ZN(n15093) );
  OAI211_X1 U12030 ( .C1(n10859), .C2(n16378), .A(n10121), .B(n15093), .ZN(
        n10127) );
  NAND2_X1 U12031 ( .A1(n15263), .A2(n12752), .ZN(n10122) );
  NAND2_X4 U12032 ( .A1(n12547), .A2(n10122), .ZN(n12518) );
  OAI21_X1 U12033 ( .B1(n12547), .B2(n12784), .A(n12518), .ZN(n11098) );
  INV_X1 U12034 ( .A(n16031), .ZN(n16078) );
  AND2_X1 U12035 ( .A1(n14862), .A2(n16078), .ZN(n16071) );
  NAND2_X1 U12036 ( .A1(n10123), .A2(n16090), .ZN(n10124) );
  XNOR2_X1 U12037 ( .A(n10858), .B(n10857), .ZN(n15091) );
  INV_X1 U12038 ( .A(n15091), .ZN(n10125) );
  AOI21_X1 U12039 ( .B1(n16369), .B2(n16158), .A(n10125), .ZN(n10126) );
  AOI211_X1 U12040 ( .C1(n15089), .C2(n16194), .A(n10127), .B(n10126), .ZN(
        n16125) );
  NAND2_X1 U12041 ( .A1(n10144), .A2(n10128), .ZN(n10130) );
  NAND2_X1 U12042 ( .A1(n10130), .A2(n10129), .ZN(n10149) );
  NAND2_X1 U12043 ( .A1(n10149), .A2(n10172), .ZN(n10854) );
  NAND2_X1 U12044 ( .A1(n10144), .A2(n10131), .ZN(n10133) );
  NAND2_X1 U12045 ( .A1(n10133), .A2(n10132), .ZN(n10853) );
  NOR2_X1 U12046 ( .A1(n10854), .A2(n10853), .ZN(n10146) );
  NOR4_X1 U12047 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n10142) );
  NOR4_X1 U12048 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n10141) );
  NOR4_X1 U12049 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n10137) );
  NOR4_X1 U12050 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n10136) );
  NOR4_X1 U12051 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n10135) );
  NOR4_X1 U12052 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n10134) );
  NAND4_X1 U12053 ( .A1(n10137), .A2(n10136), .A3(n10135), .A4(n10134), .ZN(
        n10138) );
  NOR4_X1 U12054 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        n10139), .A4(n10138), .ZN(n10140) );
  NAND3_X1 U12055 ( .A1(n10142), .A2(n10141), .A3(n10140), .ZN(n10143) );
  NAND2_X1 U12056 ( .A1(n10144), .A2(n10143), .ZN(n10171) );
  NAND2_X1 U12057 ( .A1(n10171), .A2(n10168), .ZN(n10150) );
  NAND2_X1 U12058 ( .A1(n10151), .A2(n10153), .ZN(n10177) );
  AND2_X2 U12059 ( .A1(n10146), .A2(n10855), .ZN(n16387) );
  NAND2_X1 U12060 ( .A1(n16385), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n10147) );
  OAI21_X1 U12061 ( .B1(n16125), .B2(n16385), .A(n10147), .ZN(P1_U3530) );
  INV_X1 U12062 ( .A(n10149), .ZN(n10148) );
  NAND2_X1 U12063 ( .A1(n10855), .A2(n10148), .ZN(n13081) );
  NAND2_X1 U12064 ( .A1(n14860), .A2(n14799), .ZN(n16032) );
  OR2_X1 U12065 ( .A1(n10853), .A2(n10149), .ZN(n10174) );
  NOR2_X1 U12066 ( .A1(n10174), .A2(n10150), .ZN(n10166) );
  NOR2_X1 U12067 ( .A1(n16366), .A2(n10151), .ZN(n10152) );
  INV_X1 U12068 ( .A(n11965), .ZN(n10155) );
  INV_X1 U12069 ( .A(n10153), .ZN(n10154) );
  NAND2_X1 U12070 ( .A1(n16029), .A2(n10154), .ZN(n12183) );
  INV_X1 U12071 ( .A(n12483), .ZN(n10156) );
  INV_X1 U12072 ( .A(n12547), .ZN(n10933) );
  INV_X1 U12073 ( .A(n10157), .ZN(n10160) );
  AOI22_X1 U12074 ( .A1(n11234), .A2(n16078), .B1(n10160), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n10158) );
  NAND2_X1 U12075 ( .A1(n10159), .A2(n10158), .ZN(n10163) );
  NAND2_X1 U12076 ( .A1(n10160), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10161) );
  OAI211_X1 U12077 ( .C1(n11965), .C2(n16031), .A(n10162), .B(n10161), .ZN(
        n10225) );
  NAND2_X1 U12078 ( .A1(n10163), .A2(n10225), .ZN(n10227) );
  OR2_X1 U12079 ( .A1(n10163), .A2(n10225), .ZN(n10164) );
  NAND2_X1 U12080 ( .A1(n10227), .A2(n10164), .ZN(n10357) );
  INV_X1 U12081 ( .A(n10357), .ZN(n10170) );
  AND2_X1 U12082 ( .A1(n10165), .A2(n10944), .ZN(n12754) );
  NAND2_X1 U12083 ( .A1(n10166), .A2(n10936), .ZN(n10169) );
  INV_X1 U12084 ( .A(n10172), .ZN(n10167) );
  AOI22_X1 U12085 ( .A1(n14796), .A2(n10170), .B1(n14826), .B2(n16078), .ZN(
        n10182) );
  INV_X1 U12086 ( .A(n10171), .ZN(n10173) );
  OAI21_X1 U12087 ( .B1(n10174), .B2(n10173), .A(n10172), .ZN(n10180) );
  INV_X1 U12088 ( .A(n10175), .ZN(n10176) );
  AND2_X1 U12089 ( .A1(n10177), .A2(n10176), .ZN(n10178) );
  NAND2_X1 U12090 ( .A1(n10157), .A2(n10178), .ZN(n12782) );
  INV_X1 U12091 ( .A(n12782), .ZN(n10179) );
  NAND2_X1 U12092 ( .A1(n10180), .A2(n10179), .ZN(n10738) );
  OR2_X1 U12093 ( .A1(n10738), .A2(P1_U3086), .ZN(n10309) );
  NAND2_X1 U12094 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n10309), .ZN(n10181) );
  OAI211_X1 U12095 ( .C1(n14809), .C2(n16032), .A(n10182), .B(n10181), .ZN(
        P1_U3232) );
  XOR2_X1 U12096 ( .A(n10797), .B(P2_REG2_REG_9__SCAN_IN), .Z(n10186) );
  INV_X1 U12097 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10184) );
  MUX2_X1 U12098 ( .A(n10184), .B(P2_REG2_REG_8__SCAN_IN), .S(n15822), .Z(
        n15818) );
  NOR2_X1 U12099 ( .A1(n15819), .A2(n15818), .ZN(n15816) );
  AOI21_X1 U12100 ( .B1(n15822), .B2(P2_REG2_REG_8__SCAN_IN), .A(n15816), .ZN(
        n10185) );
  NAND2_X1 U12101 ( .A1(n10185), .A2(n10186), .ZN(n10643) );
  OAI21_X1 U12102 ( .B1(n10186), .B2(n10185), .A(n10643), .ZN(n10191) );
  NAND2_X1 U12103 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n10188) );
  NAND2_X1 U12104 ( .A1(n15800), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n10187) );
  OAI211_X1 U12105 ( .C1(n14306), .C2(n10189), .A(n10188), .B(n10187), .ZN(
        n10190) );
  AOI21_X1 U12106 ( .B1(n10191), .B2(n15830), .A(n10190), .ZN(n10199) );
  INV_X1 U12107 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10193) );
  MUX2_X1 U12108 ( .A(n10193), .B(P2_REG1_REG_8__SCAN_IN), .S(n15822), .Z(
        n15814) );
  INV_X1 U12109 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10194) );
  MUX2_X1 U12110 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10194), .S(n10797), .Z(
        n10195) );
  OAI21_X1 U12111 ( .B1(n10196), .B2(n10195), .A(n10647), .ZN(n10197) );
  NAND2_X1 U12112 ( .A1(n10197), .A2(n15835), .ZN(n10198) );
  NAND2_X1 U12113 ( .A1(n10199), .A2(n10198), .ZN(P2_U3223) );
  AND2_X1 U12114 ( .A1(n15783), .A2(n10200), .ZN(n10201) );
  NAND2_X1 U12115 ( .A1(n10202), .A2(n10201), .ZN(n10203) );
  AND2_X1 U12116 ( .A1(n13091), .A2(n13350), .ZN(n10417) );
  INV_X1 U12117 ( .A(n10417), .ZN(n10204) );
  INV_X1 U12118 ( .A(n16401), .ZN(n14452) );
  AOI22_X1 U12119 ( .A1(n16405), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(n16394), .ZN(n10209) );
  INV_X1 U12120 ( .A(n10205), .ZN(n10206) );
  OAI211_X1 U12121 ( .C1(n7849), .C2(n10207), .A(n14549), .B(n10206), .ZN(
        n10208) );
  OAI211_X1 U12122 ( .C1(n14452), .C2(n13422), .A(n10209), .B(n10208), .ZN(
        P2_U3265) );
  OR2_X1 U12123 ( .A1(n14263), .A2(n13146), .ZN(n10210) );
  NAND2_X1 U12124 ( .A1(n10211), .A2(n10210), .ZN(n10212) );
  XNOR2_X1 U12125 ( .A(n13155), .B(n13157), .ZN(n13427) );
  NAND2_X1 U12126 ( .A1(n10212), .A2(n13427), .ZN(n10553) );
  OR2_X1 U12127 ( .A1(n10212), .A2(n13427), .ZN(n10213) );
  NAND2_X1 U12128 ( .A1(n10553), .A2(n10213), .ZN(n10605) );
  OAI21_X1 U12129 ( .B1(n10214), .B2(n10603), .A(n14507), .ZN(n10215) );
  AND2_X1 U12130 ( .A1(n10214), .A2(n10603), .ZN(n10583) );
  NOR2_X1 U12131 ( .A1(n10215), .A2(n10583), .ZN(n10599) );
  NAND2_X1 U12132 ( .A1(n13146), .A2(n10218), .ZN(n10216) );
  XNOR2_X1 U12133 ( .A(n10536), .B(n13427), .ZN(n10221) );
  INV_X1 U12134 ( .A(n14261), .ZN(n10674) );
  OAI22_X1 U12135 ( .A1(n10218), .A2(n14521), .B1(n10674), .B2(n14523), .ZN(
        n10219) );
  AOI21_X1 U12136 ( .B1(n10605), .B2(n14520), .A(n10219), .ZN(n10220) );
  OAI21_X1 U12137 ( .B1(n14486), .B2(n10221), .A(n10220), .ZN(n10598) );
  AOI211_X1 U12138 ( .C1(n13099), .C2(n10605), .A(n10599), .B(n10598), .ZN(
        n10258) );
  INV_X1 U12139 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10222) );
  OAI22_X1 U12140 ( .A1(n14631), .A2(n10603), .B1(n16358), .B2(n10222), .ZN(
        n10223) );
  INV_X1 U12141 ( .A(n10223), .ZN(n10224) );
  OAI21_X1 U12142 ( .B1(n10258), .B2(n16357), .A(n10224), .ZN(P2_U3504) );
  INV_X1 U12143 ( .A(n10225), .ZN(n10226) );
  OAI22_X1 U12144 ( .A1(n12483), .A2(n10123), .B1(n16090), .B2(n10228), .ZN(
        n10229) );
  INV_X1 U12145 ( .A(n10229), .ZN(n10230) );
  NAND2_X1 U12146 ( .A1(n10231), .A2(n10230), .ZN(n10232) );
  XNOR2_X1 U12147 ( .A(n10233), .B(n12203), .ZN(n10731) );
  OAI22_X1 U12148 ( .A1(n12483), .A2(n10860), .B1(n10859), .B2(n10228), .ZN(
        n10729) );
  XNOR2_X1 U12149 ( .A(n10731), .B(n10729), .ZN(n10727) );
  XOR2_X1 U12150 ( .A(n10727), .B(n10728), .Z(n10236) );
  OAI22_X1 U12151 ( .A1(n14804), .A2(n10859), .B1(n15093), .B2(n14809), .ZN(
        n10234) );
  AOI21_X1 U12152 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n10309), .A(n10234), .ZN(
        n10235) );
  OAI21_X1 U12153 ( .B1(n10236), .B2(n14829), .A(n10235), .ZN(P1_U3237) );
  NAND2_X1 U12154 ( .A1(n14668), .A2(n16170), .ZN(n14673) );
  INV_X1 U12155 ( .A(n14673), .ZN(n11915) );
  INV_X1 U12156 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10237) );
  NOR2_X1 U12157 ( .A1(n14668), .A2(n10237), .ZN(n10238) );
  AOI21_X1 U12158 ( .B1(n11915), .B2(n13146), .A(n10238), .ZN(n10239) );
  OAI21_X1 U12159 ( .B1(n10240), .B2(n16359), .A(n10239), .ZN(P2_U3442) );
  MUX2_X1 U12160 ( .A(n10250), .B(n11829), .S(n12298), .Z(n10245) );
  INV_X1 U12161 ( .A(n10245), .ZN(n10246) );
  NAND2_X1 U12162 ( .A1(n10246), .A2(SI_15_), .ZN(n10247) );
  XNOR2_X1 U12163 ( .A(n10522), .B(n10521), .ZN(n12075) );
  INV_X1 U12164 ( .A(n12075), .ZN(n10254) );
  NAND2_X1 U12165 ( .A1(n10248), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10249) );
  XNOR2_X1 U12166 ( .A(n10249), .B(P1_IR_REG_15__SCAN_IN), .ZN(n12076) );
  INV_X1 U12167 ( .A(n12076), .ZN(n15853) );
  OAI222_X1 U12168 ( .A1(n15262), .A2(n10250), .B1(n15260), .B2(n10254), .C1(
        n15853), .C2(P1_U3086), .ZN(P1_U3340) );
  OAI21_X1 U12169 ( .B1(n10251), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n10253) );
  INV_X1 U12170 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n10252) );
  XNOR2_X1 U12171 ( .A(n10253), .B(n10252), .ZN(n15836) );
  OAI222_X1 U12172 ( .A1(n14693), .A2(n11829), .B1(n14691), .B2(n10254), .C1(
        n15836), .C2(P2_U3088), .ZN(P2_U3312) );
  INV_X1 U12173 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10255) );
  OAI22_X1 U12174 ( .A1(n14673), .A2(n10603), .B1(n14668), .B2(n10255), .ZN(
        n10256) );
  INV_X1 U12175 ( .A(n10256), .ZN(n10257) );
  OAI21_X1 U12176 ( .B1(n10258), .B2(n16359), .A(n10257), .ZN(P2_U3445) );
  XNOR2_X1 U12177 ( .A(n10287), .B(n10289), .ZN(n10290) );
  OAI22_X1 U12178 ( .A1(n10261), .A2(n10260), .B1(n10259), .B2(n10268), .ZN(
        n10291) );
  XOR2_X1 U12179 ( .A(n10290), .B(n10291), .Z(n10281) );
  NAND2_X1 U12180 ( .A1(n10268), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10262) );
  NAND2_X1 U12181 ( .A1(n10263), .A2(n10262), .ZN(n10264) );
  INV_X1 U12182 ( .A(n10289), .ZN(n10271) );
  NAND2_X1 U12183 ( .A1(n10264), .A2(n10271), .ZN(n10478) );
  OAI21_X1 U12184 ( .B1(n10266), .B2(P3_REG2_REG_3__SCAN_IN), .A(n10480), .ZN(
        n10267) );
  NAND2_X1 U12185 ( .A1(n15966), .A2(n10267), .ZN(n10278) );
  NAND2_X1 U12186 ( .A1(n10268), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10269) );
  NAND2_X1 U12187 ( .A1(n10270), .A2(n10269), .ZN(n10272) );
  NAND2_X1 U12188 ( .A1(n10272), .A2(n10271), .ZN(n10472) );
  AND2_X1 U12189 ( .A1(n10273), .A2(n10472), .ZN(n10274) );
  OAI21_X1 U12190 ( .B1(n10274), .B2(P3_REG1_REG_3__SCAN_IN), .A(n10474), .ZN(
        n10275) );
  NAND2_X1 U12191 ( .A1(n15931), .A2(n10275), .ZN(n10277) );
  INV_X1 U12192 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n11328) );
  NOR2_X1 U12193 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11328), .ZN(n10770) );
  AOI21_X1 U12194 ( .B1(n15961), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10770), .ZN(
        n10276) );
  NAND3_X1 U12195 ( .A1(n10278), .A2(n10277), .A3(n10276), .ZN(n10279) );
  AOI21_X1 U12196 ( .B1(n10289), .B2(n13713), .A(n10279), .ZN(n10280) );
  OAI21_X1 U12197 ( .B1(n10281), .B2(n15991), .A(n10280), .ZN(P3_U3185) );
  INV_X1 U12198 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10282) );
  OAI22_X1 U12199 ( .A1(n14673), .A2(n10283), .B1(n14668), .B2(n10282), .ZN(
        n10284) );
  INV_X1 U12200 ( .A(n10284), .ZN(n10285) );
  OAI21_X1 U12201 ( .B1(n10286), .B2(n16359), .A(n10285), .ZN(P2_U3433) );
  XNOR2_X1 U12202 ( .A(n10489), .B(n10497), .ZN(n10491) );
  INV_X1 U12203 ( .A(n10287), .ZN(n10288) );
  AOI22_X1 U12204 ( .A1(n10291), .A2(n10290), .B1(n10289), .B2(n10288), .ZN(
        n10469) );
  XNOR2_X1 U12205 ( .A(n10292), .B(n10485), .ZN(n10468) );
  XOR2_X1 U12206 ( .A(n10491), .B(n10492), .Z(n10304) );
  XNOR2_X1 U12207 ( .A(n10485), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n10479) );
  AOI21_X1 U12208 ( .B1(n10480), .B2(n10478), .A(n10479), .ZN(n10482) );
  XNOR2_X1 U12209 ( .A(n10505), .B(n10497), .ZN(n10293) );
  AOI21_X1 U12210 ( .B1(n8864), .B2(n10293), .A(n10506), .ZN(n10301) );
  AND2_X1 U12211 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n11211) );
  AOI21_X1 U12212 ( .B1(n15961), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11211), .ZN(
        n10300) );
  NAND2_X1 U12213 ( .A1(n10474), .A2(n10472), .ZN(n10295) );
  INV_X1 U12214 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10294) );
  XNOR2_X1 U12215 ( .A(n10485), .B(n10294), .ZN(n10471) );
  NAND2_X1 U12216 ( .A1(n10295), .A2(n10471), .ZN(n10476) );
  NAND2_X1 U12217 ( .A1(n10485), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n10296) );
  NAND2_X1 U12218 ( .A1(n10476), .A2(n10296), .ZN(n10498) );
  NAND2_X1 U12219 ( .A1(n10297), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n10500) );
  OAI21_X1 U12220 ( .B1(n10297), .B2(P3_REG1_REG_5__SCAN_IN), .A(n10500), .ZN(
        n10298) );
  NAND2_X1 U12221 ( .A1(n15931), .A2(n10298), .ZN(n10299) );
  OAI211_X1 U12222 ( .C1(n15999), .C2(n10301), .A(n10300), .B(n10299), .ZN(
        n10302) );
  AOI21_X1 U12223 ( .B1(n10497), .B2(n13713), .A(n10302), .ZN(n10303) );
  OAI21_X1 U12224 ( .B1(n10304), .B2(n15991), .A(n10303), .ZN(P3_U3187) );
  XOR2_X1 U12225 ( .A(n10305), .B(n10306), .Z(n10311) );
  INV_X1 U12226 ( .A(n14799), .ZN(n14787) );
  NOR2_X1 U12227 ( .A1(n10860), .A2(n14787), .ZN(n16085) );
  AND2_X1 U12228 ( .A1(n14862), .A2(n14806), .ZN(n16076) );
  INV_X1 U12229 ( .A(n14809), .ZN(n14821) );
  OAI21_X1 U12230 ( .B1(n16085), .B2(n16076), .A(n14821), .ZN(n10307) );
  OAI21_X1 U12231 ( .B1(n14804), .B2(n16090), .A(n10307), .ZN(n10308) );
  AOI21_X1 U12232 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n10309), .A(n10308), .ZN(
        n10310) );
  OAI21_X1 U12233 ( .B1(n10311), .B2(n14829), .A(n10310), .ZN(P1_U3222) );
  INV_X1 U12234 ( .A(n10312), .ZN(n10313) );
  OAI222_X1 U12235 ( .A1(P3_U3151), .A2(n10314), .B1(n14119), .B2(n10313), 
        .C1(n15280), .C2(n13462), .ZN(P3_U3275) );
  XOR2_X1 U12236 ( .A(n10316), .B(n10315), .Z(n10329) );
  INV_X1 U12237 ( .A(n10317), .ZN(n10318) );
  AOI21_X1 U12238 ( .B1(n8813), .B2(n10319), .A(n10318), .ZN(n10321) );
  AOI22_X1 U12239 ( .A1(n15961), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10320) );
  OAI21_X1 U12240 ( .B1(n15993), .B2(n10321), .A(n10320), .ZN(n10326) );
  NAND2_X1 U12241 ( .A1(n10322), .A2(n8814), .ZN(n10323) );
  AOI21_X1 U12242 ( .B1(n10324), .B2(n10323), .A(n15999), .ZN(n10325) );
  AOI211_X1 U12243 ( .C1(n13713), .C2(n8065), .A(n10326), .B(n10325), .ZN(
        n10328) );
  OAI21_X1 U12244 ( .B1(n15991), .B2(n10329), .A(n10328), .ZN(P3_U3183) );
  INV_X1 U12245 ( .A(n10340), .ZN(n10336) );
  INV_X1 U12246 ( .A(n10341), .ZN(n10330) );
  OR2_X1 U12247 ( .A1(n10345), .A2(n10330), .ZN(n10335) );
  AND3_X1 U12248 ( .A1(n10333), .A2(n10332), .A3(n10331), .ZN(n10334) );
  OAI211_X1 U12249 ( .C1(n10348), .C2(n10336), .A(n10335), .B(n10334), .ZN(
        n10337) );
  NAND2_X1 U12250 ( .A1(n10337), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10339) );
  OR2_X1 U12251 ( .A1(n13039), .A2(n10345), .ZN(n10338) );
  NOR2_X1 U12252 ( .A1(n13568), .A2(P3_U3151), .ZN(n10632) );
  INV_X1 U12253 ( .A(n16055), .ZN(n10638) );
  NAND2_X1 U12254 ( .A1(n13624), .A2(n10638), .ZN(n12865) );
  AND2_X1 U12255 ( .A1(n16051), .A2(n12865), .ZN(n12999) );
  INV_X1 U12256 ( .A(n12999), .ZN(n10352) );
  NAND3_X1 U12257 ( .A1(n10348), .A2(n10340), .A3(n16311), .ZN(n10343) );
  NAND2_X1 U12258 ( .A1(n10345), .A2(n10341), .ZN(n10342) );
  NAND2_X1 U12259 ( .A1(n10343), .A2(n10342), .ZN(n10344) );
  INV_X1 U12260 ( .A(n10345), .ZN(n10346) );
  NOR2_X1 U12261 ( .A1(n10346), .A2(n13039), .ZN(n10463) );
  INV_X1 U12262 ( .A(n10463), .ZN(n10347) );
  INV_X1 U12263 ( .A(n13602), .ZN(n13575) );
  NOR2_X1 U12264 ( .A1(n10348), .A2(n13036), .ZN(n10350) );
  NAND2_X1 U12265 ( .A1(n10349), .A2(n16200), .ZN(n11091) );
  OAI22_X1 U12266 ( .A1(n13575), .A2(n16104), .B1(n10638), .B2(n13595), .ZN(
        n10351) );
  AOI21_X1 U12267 ( .B1(n10352), .B2(n13587), .A(n10351), .ZN(n10353) );
  OAI21_X1 U12268 ( .B1(n10632), .B2(n10354), .A(n10353), .ZN(P3_U3172) );
  INV_X1 U12269 ( .A(SI_21_), .ZN(n10355) );
  OAI222_X1 U12270 ( .A1(n14119), .A2(n10356), .B1(n13462), .B2(n10355), .C1(
        P3_U3151), .C2(n10454), .ZN(P3_U3274) );
  MUX2_X1 U12271 ( .A(n10357), .B(n14864), .S(n12781), .Z(n10362) );
  NAND2_X1 U12272 ( .A1(n10358), .A2(n8323), .ZN(n10359) );
  NAND2_X1 U12273 ( .A1(n14861), .A2(n10359), .ZN(n10360) );
  AOI21_X1 U12274 ( .B1(n10362), .B2(n10361), .A(n10360), .ZN(n16024) );
  XNOR2_X1 U12275 ( .A(n10364), .B(n10363), .ZN(n10374) );
  OAI211_X1 U12276 ( .C1(n10367), .C2(n10366), .A(n7422), .B(n10365), .ZN(
        n10373) );
  INV_X1 U12277 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10369) );
  INV_X1 U12278 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10368) );
  OAI22_X1 U12279 ( .A1(n16028), .A2(n10369), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10368), .ZN(n10370) );
  AOI21_X1 U12280 ( .B1(n10371), .B2(n14900), .A(n10370), .ZN(n10372) );
  OAI211_X1 U12281 ( .C1(n10374), .C2(n15852), .A(n10373), .B(n10372), .ZN(
        n10375) );
  OR2_X1 U12282 ( .A1(n16024), .A2(n10375), .ZN(P1_U3245) );
  AOI21_X1 U12283 ( .B1(n10378), .B2(n10377), .A(n10376), .ZN(n10386) );
  NAND2_X1 U12284 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n11986)
         );
  OAI21_X1 U12285 ( .B1(n16028), .B2(n15694), .A(n11986), .ZN(n10384) );
  AND3_X1 U12286 ( .A1(n10446), .A2(n10380), .A3(n10379), .ZN(n10381) );
  NOR3_X1 U12288 ( .A1(n10382), .A2(n10381), .A3(n16423), .ZN(n10383) );
  AOI211_X1 U12289 ( .C1(n14900), .C2(n11551), .A(n10384), .B(n10383), .ZN(
        n10385) );
  OAI21_X1 U12290 ( .B1(n10386), .B2(n15852), .A(n10385), .ZN(P1_U3254) );
  OAI21_X1 U12291 ( .B1(n11563), .B2(P1_REG1_REG_12__SCAN_IN), .A(n10387), 
        .ZN(n10389) );
  INV_X1 U12292 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n16386) );
  MUX2_X1 U12293 ( .A(n16386), .B(P1_REG1_REG_13__SCAN_IN), .S(n11781), .Z(
        n10388) );
  NOR2_X1 U12294 ( .A1(n10389), .A2(n10388), .ZN(n11195) );
  AOI211_X1 U12295 ( .C1(n10389), .C2(n10388), .A(n15852), .B(n11195), .ZN(
        n10396) );
  OAI21_X1 U12296 ( .B1(n11563), .B2(P1_REG2_REG_12__SCAN_IN), .A(n10390), 
        .ZN(n10392) );
  INV_X1 U12297 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11184) );
  MUX2_X1 U12298 ( .A(n11184), .B(P1_REG2_REG_13__SCAN_IN), .S(n11781), .Z(
        n10391) );
  NOR2_X1 U12299 ( .A1(n10392), .A2(n10391), .ZN(n14907) );
  AOI211_X1 U12300 ( .C1(n10392), .C2(n10391), .A(n16423), .B(n14907), .ZN(
        n10395) );
  INV_X1 U12301 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n15758) );
  NAND2_X1 U12302 ( .A1(n14900), .A2(n11781), .ZN(n10393) );
  NAND2_X1 U12303 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n12210)
         );
  OAI211_X1 U12304 ( .C1(n15758), .C2(n16028), .A(n10393), .B(n12210), .ZN(
        n10394) );
  OR3_X1 U12305 ( .A1(n10396), .A2(n10395), .A3(n10394), .ZN(P1_U3256) );
  NAND2_X1 U12306 ( .A1(n14260), .A2(n7431), .ZN(n10612) );
  NAND2_X1 U12307 ( .A1(n11045), .A2(n9720), .ZN(n10399) );
  AOI22_X1 U12308 ( .A1(n9659), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n13109), 
        .B2(n10397), .ZN(n10398) );
  XNOR2_X1 U12309 ( .A(n16246), .B(n11516), .ZN(n10614) );
  XOR2_X1 U12310 ( .A(n10612), .B(n10614), .Z(n10404) );
  INV_X1 U12311 ( .A(n10400), .ZN(n10401) );
  AOI21_X1 U12312 ( .B1(n10404), .B2(n10403), .A(n7604), .ZN(n10415) );
  NAND2_X1 U12313 ( .A1(n9742), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10410) );
  NAND2_X1 U12314 ( .A1(n10405), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n10542) );
  OR2_X1 U12315 ( .A1(n10405), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n10406) );
  AND2_X1 U12316 ( .A1(n10542), .A2(n10406), .ZN(n10622) );
  NAND2_X1 U12317 ( .A1(n11931), .A2(n10622), .ZN(n10409) );
  NAND2_X1 U12318 ( .A1(n13386), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n10408) );
  NAND2_X1 U12319 ( .A1(n13368), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10407) );
  NAND4_X1 U12320 ( .A1(n10410), .A2(n10409), .A3(n10408), .A4(n10407), .ZN(
        n14259) );
  INV_X1 U12321 ( .A(n14259), .ZN(n10794) );
  INV_X1 U12322 ( .A(n14218), .ZN(n14242) );
  AOI22_X1 U12323 ( .A1(n14227), .A2(n14261), .B1(n16248), .B2(n14242), .ZN(
        n10412) );
  OAI211_X1 U12324 ( .C1(n10794), .C2(n14217), .A(n10412), .B(n10411), .ZN(
        n10413) );
  AOI21_X1 U12325 ( .B1(n16246), .B2(n14246), .A(n10413), .ZN(n10414) );
  OAI21_X1 U12326 ( .B1(n10415), .B2(n14248), .A(n10414), .ZN(P2_U3185) );
  INV_X1 U12327 ( .A(n10416), .ZN(n10426) );
  INV_X2 U12328 ( .A(n14539), .ZN(n16306) );
  OR2_X2 U12329 ( .A1(n16405), .A2(n10418), .ZN(n16398) );
  INV_X1 U12330 ( .A(n13146), .ZN(n10420) );
  OAI22_X1 U12331 ( .A1(n16398), .A2(n10420), .B1(n10419), .B2(n14510), .ZN(
        n10421) );
  AOI21_X1 U12332 ( .B1(n16306), .B2(n10422), .A(n10421), .ZN(n10425) );
  MUX2_X1 U12333 ( .A(n9556), .B(n10423), .S(n14549), .Z(n10424) );
  OAI211_X1 U12334 ( .C1(n10426), .C2(n14497), .A(n10425), .B(n10424), .ZN(
        P2_U3261) );
  OAI21_X1 U12335 ( .B1(n10428), .B2(n13424), .A(n10427), .ZN(n10429) );
  INV_X1 U12336 ( .A(n10429), .ZN(n16173) );
  OAI21_X1 U12337 ( .B1(n10432), .B2(n10431), .A(n10430), .ZN(n10433) );
  AOI222_X1 U12338 ( .A1(n14529), .A2(n10433), .B1(n14263), .B2(n14439), .C1(
        n14265), .C2(n14438), .ZN(n16172) );
  MUX2_X1 U12339 ( .A(n9554), .B(n16172), .S(n14549), .Z(n10439) );
  AOI21_X1 U12340 ( .B1(n10665), .B2(n16169), .A(n7431), .ZN(n10435) );
  AND2_X1 U12341 ( .A1(n10435), .A2(n10434), .ZN(n16168) );
  OAI22_X1 U12342 ( .A1(n16398), .A2(n10436), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n14510), .ZN(n10437) );
  AOI21_X1 U12343 ( .B1(n16306), .B2(n16168), .A(n10437), .ZN(n10438) );
  OAI211_X1 U12344 ( .C1(n16173), .C2(n14497), .A(n10439), .B(n10438), .ZN(
        P2_U3262) );
  AOI21_X1 U12345 ( .B1(n10441), .B2(n10440), .A(n15852), .ZN(n10443) );
  NAND2_X1 U12346 ( .A1(n10443), .A2(n10442), .ZN(n10451) );
  NAND2_X1 U12347 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n11743)
         );
  AOI21_X1 U12348 ( .B1(n10445), .B2(n10444), .A(n16423), .ZN(n10447) );
  NAND2_X1 U12349 ( .A1(n10447), .A2(n10446), .ZN(n10448) );
  NAND2_X1 U12350 ( .A1(n11743), .A2(n10448), .ZN(n10449) );
  AOI21_X1 U12351 ( .B1(n14866), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n10449), 
        .ZN(n10450) );
  OAI211_X1 U12352 ( .C1(n16022), .C2(n10452), .A(n10451), .B(n10450), .ZN(
        P1_U3253) );
  OAI21_X1 U12353 ( .B1(n10454), .B2(n10453), .A(n12996), .ZN(n10455) );
  INV_X1 U12354 ( .A(n10455), .ZN(n10456) );
  MUX2_X1 U12355 ( .A(n8025), .B(n13624), .S(n16055), .Z(n10460) );
  NAND2_X1 U12356 ( .A1(n10638), .A2(n12836), .ZN(n10459) );
  AOI21_X1 U12357 ( .B1(n10461), .B2(n10460), .A(n7607), .ZN(n10467) );
  INV_X1 U12358 ( .A(n13600), .ZN(n13589) );
  OAI22_X1 U12359 ( .A1(n13575), .A2(n16052), .B1(n7738), .B2(n13595), .ZN(
        n10465) );
  NOR2_X1 U12360 ( .A1(n10632), .A2(n16070), .ZN(n10464) );
  AOI211_X1 U12361 ( .C1(n13589), .C2(n13624), .A(n10465), .B(n10464), .ZN(
        n10466) );
  OAI21_X1 U12362 ( .B1(n10467), .B2(n13608), .A(n10466), .ZN(P3_U3162) );
  XNOR2_X1 U12363 ( .A(n10469), .B(n10468), .ZN(n10487) );
  INV_X1 U12364 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10470) );
  NOR2_X1 U12365 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10470), .ZN(n11038) );
  INV_X1 U12366 ( .A(n10471), .ZN(n10473) );
  NAND3_X1 U12367 ( .A1(n10474), .A2(n10473), .A3(n10472), .ZN(n10475) );
  AOI21_X1 U12368 ( .B1(n10476), .B2(n10475), .A(n15993), .ZN(n10477) );
  AOI211_X1 U12369 ( .C1(n15961), .C2(P3_ADDR_REG_4__SCAN_IN), .A(n11038), .B(
        n10477), .ZN(n10484) );
  AND3_X1 U12370 ( .A1(n10480), .A2(n10479), .A3(n10478), .ZN(n10481) );
  OAI21_X1 U12371 ( .B1(n10482), .B2(n10481), .A(n15966), .ZN(n10483) );
  OAI211_X1 U12372 ( .C1(n15984), .C2(n10485), .A(n10484), .B(n10483), .ZN(
        n10486) );
  AOI21_X1 U12373 ( .B1(n15970), .B2(n10487), .A(n10486), .ZN(n10488) );
  INV_X1 U12374 ( .A(n10488), .ZN(P3_U3186) );
  INV_X1 U12375 ( .A(n10489), .ZN(n10490) );
  MUX2_X1 U12376 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n8634), .Z(n10493) );
  AND2_X1 U12377 ( .A1(n10493), .A2(n10573), .ZN(n10564) );
  INV_X1 U12378 ( .A(n10564), .ZN(n10495) );
  INV_X1 U12379 ( .A(n10493), .ZN(n10494) );
  NAND2_X1 U12380 ( .A1(n10494), .A2(n10514), .ZN(n10565) );
  NAND2_X1 U12381 ( .A1(n10495), .A2(n10565), .ZN(n10496) );
  XNOR2_X1 U12382 ( .A(n10566), .B(n10496), .ZN(n10519) );
  INV_X1 U12383 ( .A(n10497), .ZN(n10508) );
  NAND2_X1 U12384 ( .A1(n10498), .A2(n10508), .ZN(n10499) );
  AND2_X1 U12385 ( .A1(n10500), .A2(n10499), .ZN(n10503) );
  NAND2_X1 U12386 ( .A1(P3_REG1_REG_6__SCAN_IN), .A2(n10573), .ZN(n10501) );
  OAI21_X1 U12387 ( .B1(P3_REG1_REG_6__SCAN_IN), .B2(n10573), .A(n10501), .ZN(
        n10502) );
  AOI21_X1 U12388 ( .B1(n10503), .B2(n10502), .A(n10560), .ZN(n10517) );
  INV_X1 U12389 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n10504) );
  NOR2_X1 U12390 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10504), .ZN(n11308) );
  INV_X1 U12391 ( .A(n10505), .ZN(n10507) );
  NAND2_X1 U12392 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n10573), .ZN(n10509) );
  OAI21_X1 U12393 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n10573), .A(n10509), .ZN(
        n10510) );
  AOI21_X1 U12394 ( .B1(n10511), .B2(n10510), .A(n10572), .ZN(n10512) );
  NOR2_X1 U12395 ( .A1(n15999), .A2(n10512), .ZN(n10513) );
  AOI211_X1 U12396 ( .C1(n15961), .C2(P3_ADDR_REG_6__SCAN_IN), .A(n11308), .B(
        n10513), .ZN(n10516) );
  NAND2_X1 U12397 ( .A1(n13713), .A2(n10514), .ZN(n10515) );
  OAI211_X1 U12398 ( .C1(n10517), .C2(n15993), .A(n10516), .B(n10515), .ZN(
        n10518) );
  AOI21_X1 U12399 ( .B1(n10519), .B2(n15970), .A(n10518), .ZN(n10520) );
  INV_X1 U12400 ( .A(n10520), .ZN(P3_U3188) );
  XNOR2_X1 U12401 ( .A(n10777), .B(SI_16_), .ZN(n10751) );
  INV_X1 U12402 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10611) );
  MUX2_X1 U12403 ( .A(n10525), .B(n10611), .S(n12298), .Z(n10773) );
  XNOR2_X1 U12404 ( .A(n10751), .B(n10773), .ZN(n12175) );
  INV_X1 U12405 ( .A(n12175), .ZN(n10610) );
  INV_X1 U12406 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n15447) );
  NAND2_X1 U12407 ( .A1(n10526), .A2(n15447), .ZN(n10528) );
  NAND2_X1 U12408 ( .A1(n10528), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10527) );
  MUX2_X1 U12409 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10527), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n10529) );
  AND2_X1 U12410 ( .A1(n10529), .A2(n10757), .ZN(n12176) );
  AOI22_X1 U12411 ( .A1(n12176), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10530), .ZN(n10531) );
  OAI21_X1 U12412 ( .B1(n10610), .B2(n15260), .A(n10531), .ZN(P1_U3339) );
  INV_X1 U12413 ( .A(n10532), .ZN(n10534) );
  OAI22_X1 U12414 ( .A1(n13040), .A2(P3_U3151), .B1(SI_22_), .B2(n13462), .ZN(
        n10533) );
  AOI21_X1 U12415 ( .B1(n10534), .B2(n16291), .A(n10533), .ZN(P3_U3273) );
  OR2_X1 U12416 ( .A1(n13155), .A2(n13157), .ZN(n10535) );
  NAND2_X1 U12417 ( .A1(n13155), .A2(n13157), .ZN(n10537) );
  XNOR2_X1 U12418 ( .A(n16223), .B(n14261), .ZN(n13429) );
  INV_X1 U12419 ( .A(n14260), .ZN(n13167) );
  OR2_X1 U12420 ( .A1(n16246), .A2(n13167), .ZN(n10675) );
  INV_X1 U12421 ( .A(n10540), .ZN(n10541) );
  NAND2_X1 U12422 ( .A1(n11356), .A2(n9720), .ZN(n10539) );
  AOI22_X1 U12423 ( .A1(n9659), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n15822), 
        .B2(n13109), .ZN(n10538) );
  NAND2_X1 U12424 ( .A1(n10539), .A2(n10538), .ZN(n13178) );
  XNOR2_X1 U12425 ( .A(n13178), .B(n14259), .ZN(n13431) );
  INV_X1 U12426 ( .A(n13431), .ZN(n10554) );
  OAI21_X1 U12427 ( .B1(n10541), .B2(n13431), .A(n10796), .ZN(n10549) );
  NAND2_X1 U12428 ( .A1(n9742), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n10547) );
  NAND2_X1 U12429 ( .A1(n10542), .A2(n10925), .ZN(n10543) );
  AND2_X1 U12430 ( .A1(n10800), .A2(n10543), .ZN(n10928) );
  NAND2_X1 U12431 ( .A1(n11931), .A2(n10928), .ZN(n10546) );
  NAND2_X1 U12432 ( .A1(n13386), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n10545) );
  NAND2_X1 U12433 ( .A1(n13368), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10544) );
  NAND4_X1 U12434 ( .A1(n10547), .A2(n10546), .A3(n10545), .A4(n10544), .ZN(
        n14258) );
  AOI22_X1 U12435 ( .A1(n14439), .A2(n14258), .B1(n14260), .B2(n14438), .ZN(
        n10620) );
  INV_X1 U12436 ( .A(n10620), .ZN(n10548) );
  AOI21_X1 U12437 ( .B1(n10549), .B2(n14529), .A(n10548), .ZN(n16266) );
  INV_X1 U12438 ( .A(n16223), .ZN(n10594) );
  NAND2_X1 U12439 ( .A1(n10583), .A2(n10594), .ZN(n10684) );
  AOI21_X1 U12440 ( .B1(n10683), .B2(n13178), .A(n7431), .ZN(n10550) );
  AND2_X1 U12441 ( .A1(n10813), .A2(n10550), .ZN(n16264) );
  AOI22_X1 U12442 ( .A1(n16405), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n10622), 
        .B2(n16394), .ZN(n10551) );
  OAI21_X1 U12443 ( .B1(n16398), .B2(n8270), .A(n10551), .ZN(n10558) );
  OR2_X1 U12444 ( .A1(n13155), .A2(n14262), .ZN(n10552) );
  INV_X1 U12445 ( .A(n13429), .ZN(n10586) );
  OR2_X1 U12446 ( .A1(n16246), .A2(n14260), .ZN(n10672) );
  NAND2_X1 U12447 ( .A1(n16246), .A2(n14260), .ZN(n10671) );
  NOR2_X1 U12448 ( .A1(n10555), .A2(n10554), .ZN(n16263) );
  INV_X1 U12449 ( .A(n16269), .ZN(n10556) );
  NOR3_X1 U12450 ( .A1(n16263), .A2(n10556), .A3(n14497), .ZN(n10557) );
  AOI211_X1 U12451 ( .C1(n16264), .C2(n16306), .A(n10558), .B(n10557), .ZN(
        n10559) );
  OAI21_X1 U12452 ( .B1(n16405), .B2(n16266), .A(n10559), .ZN(P2_U3257) );
  INV_X1 U12453 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n16236) );
  XNOR2_X1 U12454 ( .A(n10691), .B(n10708), .ZN(n10561) );
  AOI21_X1 U12455 ( .B1(n16236), .B2(n10561), .A(n10692), .ZN(n10580) );
  NOR2_X1 U12456 ( .A1(n10563), .A2(n10562), .ZN(n10697) );
  AOI21_X1 U12457 ( .B1(n10563), .B2(n10562), .A(n10697), .ZN(n10568) );
  AOI21_X1 U12458 ( .B1(n10566), .B2(n10565), .A(n10564), .ZN(n10567) );
  NAND2_X1 U12459 ( .A1(n10567), .A2(n10568), .ZN(n10703) );
  OAI21_X1 U12460 ( .B1(n10568), .B2(n10567), .A(n10703), .ZN(n10569) );
  NAND2_X1 U12461 ( .A1(n10569), .A2(n15970), .ZN(n10579) );
  INV_X1 U12462 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n15682) );
  INV_X1 U12463 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n10570) );
  NOR2_X1 U12464 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10570), .ZN(n11628) );
  INV_X1 U12465 ( .A(n11628), .ZN(n10571) );
  OAI21_X1 U12466 ( .B1(n15982), .B2(n15682), .A(n10571), .ZN(n10577) );
  AOI21_X1 U12467 ( .B1(n8896), .B2(n10574), .A(n10709), .ZN(n10575) );
  NOR2_X1 U12468 ( .A1(n10575), .A2(n15999), .ZN(n10576) );
  AOI211_X1 U12469 ( .C1(n13713), .C2(n10708), .A(n10577), .B(n10576), .ZN(
        n10578) );
  OAI211_X1 U12470 ( .C1(n10580), .C2(n15993), .A(n10579), .B(n10578), .ZN(
        P3_U3189) );
  OAI21_X1 U12471 ( .B1(n10582), .B2(n10586), .A(n10581), .ZN(n16225) );
  INV_X1 U12472 ( .A(n10583), .ZN(n10585) );
  INV_X1 U12473 ( .A(n10684), .ZN(n10584) );
  AOI211_X1 U12474 ( .C1(n16223), .C2(n10585), .A(n7431), .B(n10584), .ZN(
        n16224) );
  XNOR2_X1 U12475 ( .A(n10587), .B(n10586), .ZN(n10588) );
  NOR2_X1 U12476 ( .A1(n10588), .A2(n14486), .ZN(n10589) );
  AOI211_X1 U12477 ( .C1(n14520), .C2(n16225), .A(n10590), .B(n10589), .ZN(
        n16228) );
  INV_X1 U12478 ( .A(n16228), .ZN(n10591) );
  AOI211_X1 U12479 ( .C1(n13099), .C2(n16225), .A(n16224), .B(n10591), .ZN(
        n10597) );
  AOI22_X1 U12480 ( .A1(n11917), .A2(n16223), .B1(n16357), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n10592) );
  OAI21_X1 U12481 ( .B1(n10597), .B2(n16357), .A(n10592), .ZN(P2_U3505) );
  INV_X1 U12482 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10593) );
  OAI22_X1 U12483 ( .A1(n14673), .A2(n10594), .B1(n14668), .B2(n10593), .ZN(
        n10595) );
  INV_X1 U12484 ( .A(n10595), .ZN(n10596) );
  OAI21_X1 U12485 ( .B1(n10597), .B2(n16359), .A(n10596), .ZN(P2_U3448) );
  INV_X1 U12486 ( .A(n10598), .ZN(n10607) );
  NAND2_X1 U12487 ( .A1(n16306), .A2(n10599), .ZN(n10602) );
  AOI22_X1 U12488 ( .A1(n16405), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n10600), 
        .B2(n16394), .ZN(n10601) );
  OAI211_X1 U12489 ( .C1(n10603), .C2(n16398), .A(n10602), .B(n10601), .ZN(
        n10604) );
  AOI21_X1 U12490 ( .B1(n16401), .B2(n10605), .A(n10604), .ZN(n10606) );
  OAI21_X1 U12491 ( .B1(n10607), .B2(n16405), .A(n10606), .ZN(P2_U3260) );
  XNOR2_X1 U12492 ( .A(n10608), .B(P2_IR_REG_16__SCAN_IN), .ZN(n14273) );
  INV_X1 U12493 ( .A(n14273), .ZN(n10609) );
  OAI222_X1 U12494 ( .A1(n14693), .A2(n10611), .B1(n14691), .B2(n10610), .C1(
        n10609), .C2(P2_U3088), .ZN(P2_U3311) );
  INV_X1 U12495 ( .A(n10612), .ZN(n10613) );
  NOR2_X1 U12496 ( .A1(n10614), .A2(n10613), .ZN(n10616) );
  XNOR2_X1 U12497 ( .A(n13178), .B(n11516), .ZN(n10919) );
  NAND2_X1 U12498 ( .A1(n14259), .A2(n14445), .ZN(n10917) );
  XNOR2_X1 U12499 ( .A(n10919), .B(n10917), .ZN(n10615) );
  INV_X1 U12500 ( .A(n10918), .ZN(n10618) );
  NOR3_X1 U12501 ( .A1(n7604), .A2(n10616), .A3(n10615), .ZN(n10617) );
  OAI21_X1 U12502 ( .B1(n10618), .B2(n10617), .A(n14232), .ZN(n10624) );
  INV_X1 U12503 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10619) );
  OAI22_X1 U12504 ( .A1(n14244), .A2(n10620), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10619), .ZN(n10621) );
  AOI21_X1 U12505 ( .B1(n10622), .B2(n14242), .A(n10621), .ZN(n10623) );
  OAI211_X1 U12506 ( .C1(n8270), .C2(n12244), .A(n10624), .B(n10623), .ZN(
        P2_U3193) );
  XNOR2_X1 U12507 ( .A(n10625), .B(n10763), .ZN(n10762) );
  XNOR2_X1 U12508 ( .A(n10762), .B(n13622), .ZN(n10627) );
  OAI21_X1 U12509 ( .B1(n10627), .B2(n10626), .A(n10766), .ZN(n10628) );
  NAND2_X1 U12510 ( .A1(n10628), .A2(n13587), .ZN(n10631) );
  OAI22_X1 U12511 ( .A1(n13575), .A2(n16102), .B1(n13595), .B2(n16116), .ZN(
        n10629) );
  AOI21_X1 U12512 ( .B1(n13589), .B2(n7428), .A(n10629), .ZN(n10630) );
  OAI211_X1 U12513 ( .C1(n10632), .C2(n16114), .A(n10631), .B(n10630), .ZN(
        P3_U3177) );
  OR3_X1 U12514 ( .A1(n12999), .A2(n16200), .A3(n10633), .ZN(n10634) );
  OAI21_X1 U12515 ( .B1(n16104), .B2(n16101), .A(n10634), .ZN(n11092) );
  OAI22_X1 U12516 ( .A1(n14030), .A2(n10638), .B1(n16407), .B2(n8387), .ZN(
        n10635) );
  AOI21_X1 U12517 ( .B1(n11092), .B2(n16407), .A(n10635), .ZN(n10636) );
  INV_X1 U12518 ( .A(n10636), .ZN(P3_U3459) );
  INV_X1 U12519 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10637) );
  OAI22_X1 U12520 ( .A1(n10638), .A2(n14102), .B1(n16410), .B2(n10637), .ZN(
        n10639) );
  AOI21_X1 U12521 ( .B1(n11092), .B2(n16410), .A(n10639), .ZN(n10640) );
  INV_X1 U12522 ( .A(n10640), .ZN(P3_U3390) );
  INV_X1 U12523 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10641) );
  MUX2_X1 U12524 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n10641), .S(n11134), .Z(
        n10642) );
  INV_X1 U12525 ( .A(n10642), .ZN(n10645) );
  NOR2_X1 U12526 ( .A1(n10644), .A2(n10645), .ZN(n10834) );
  AOI211_X1 U12527 ( .C1(n10645), .C2(n10644), .A(n15817), .B(n10834), .ZN(
        n10655) );
  INV_X1 U12528 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10646) );
  MUX2_X1 U12529 ( .A(n10646), .B(P2_REG1_REG_10__SCAN_IN), .S(n11134), .Z(
        n10649) );
  OAI21_X1 U12530 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n10797), .A(n10647), .ZN(
        n10648) );
  NOR2_X1 U12531 ( .A1(n10648), .A2(n10649), .ZN(n10842) );
  AOI211_X1 U12532 ( .C1(n10649), .C2(n10648), .A(n15813), .B(n10842), .ZN(
        n10654) );
  NAND2_X1 U12533 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n10651)
         );
  NAND2_X1 U12534 ( .A1(n15800), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n10650) );
  OAI211_X1 U12535 ( .C1(n14306), .C2(n10652), .A(n10651), .B(n10650), .ZN(
        n10653) );
  OR3_X1 U12536 ( .A1(n10655), .A2(n10654), .A3(n10653), .ZN(P2_U3224) );
  INV_X1 U12537 ( .A(n14497), .ZN(n14515) );
  OAI21_X1 U12538 ( .B1(n10657), .B2(n10660), .A(n10656), .ZN(n16130) );
  NAND3_X1 U12539 ( .A1(n10660), .A2(n10659), .A3(n10658), .ZN(n10661) );
  AND2_X1 U12540 ( .A1(n10662), .A2(n10661), .ZN(n10663) );
  OAI222_X1 U12541 ( .A1(n14523), .A2(n8013), .B1(n14521), .B2(n10664), .C1(
        n14486), .C2(n10663), .ZN(n16128) );
  MUX2_X1 U12542 ( .A(n16128), .B(P2_REG2_REG_2__SCAN_IN), .S(n16405), .Z(
        n10669) );
  OAI211_X1 U12543 ( .C1(n10666), .C2(n16127), .A(n14507), .B(n10665), .ZN(
        n16126) );
  INV_X1 U12544 ( .A(n16398), .ZN(n16303) );
  AOI22_X1 U12545 ( .A1(n16303), .A2(n14224), .B1(n16394), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n10667) );
  OAI21_X1 U12546 ( .B1(n14539), .B2(n16126), .A(n10667), .ZN(n10668) );
  AOI211_X1 U12547 ( .C1(n14515), .C2(n16130), .A(n10669), .B(n10668), .ZN(
        n10670) );
  INV_X1 U12548 ( .A(n10670), .ZN(P2_U3263) );
  NAND2_X1 U12549 ( .A1(n10672), .A2(n10671), .ZN(n13428) );
  XOR2_X1 U12550 ( .A(n13428), .B(n10673), .Z(n16253) );
  INV_X1 U12551 ( .A(n16253), .ZN(n10686) );
  OAI22_X1 U12552 ( .A1(n10794), .A2(n14523), .B1(n10674), .B2(n14521), .ZN(
        n10682) );
  INV_X1 U12553 ( .A(n13428), .ZN(n10680) );
  INV_X1 U12554 ( .A(n10675), .ZN(n10676) );
  NOR2_X1 U12555 ( .A1(n10677), .A2(n10676), .ZN(n10678) );
  AOI211_X1 U12556 ( .C1(n10680), .C2(n10679), .A(n14486), .B(n10678), .ZN(
        n10681) );
  AOI211_X1 U12557 ( .C1(n16253), .C2(n14520), .A(n10682), .B(n10681), .ZN(
        n16255) );
  AOI211_X1 U12558 ( .C1(n16246), .C2(n10684), .A(n7431), .B(n8271), .ZN(
        n16247) );
  AOI21_X1 U12559 ( .B1(n16170), .B2(n16246), .A(n16247), .ZN(n10685) );
  OAI211_X1 U12560 ( .C1(n9885), .C2(n10686), .A(n16255), .B(n10685), .ZN(
        n10688) );
  NAND2_X1 U12561 ( .A1(n10688), .A2(n16358), .ZN(n10687) );
  OAI21_X1 U12562 ( .B1(n16358), .B2(n9762), .A(n10687), .ZN(P2_U3506) );
  INV_X1 U12563 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10690) );
  NAND2_X1 U12564 ( .A1(n10688), .A2(n14668), .ZN(n10689) );
  OAI21_X1 U12565 ( .B1(n14668), .B2(n10690), .A(n10689), .ZN(P2_U3451) );
  NOR2_X1 U12566 ( .A1(n10708), .A2(n10691), .ZN(n10693) );
  NAND2_X1 U12567 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n10958), .ZN(n10694) );
  OAI21_X1 U12568 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n10958), .A(n10694), .ZN(
        n10695) );
  AOI21_X1 U12569 ( .B1(n10696), .B2(n10695), .A(n10945), .ZN(n10720) );
  INV_X1 U12570 ( .A(n10697), .ZN(n10702) );
  NAND2_X1 U12571 ( .A1(n10698), .A2(n10717), .ZN(n10947) );
  INV_X1 U12572 ( .A(n10698), .ZN(n10699) );
  NAND2_X1 U12573 ( .A1(n10699), .A2(n10958), .ZN(n10700) );
  NAND2_X1 U12574 ( .A1(n10947), .A2(n10700), .ZN(n10701) );
  AND3_X1 U12575 ( .A1(n10703), .A2(n10702), .A3(n10701), .ZN(n10704) );
  OAI21_X1 U12576 ( .B1(n10954), .B2(n10704), .A(n15970), .ZN(n10719) );
  INV_X1 U12577 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15667) );
  NOR2_X1 U12578 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10705), .ZN(n11619) );
  INV_X1 U12579 ( .A(n11619), .ZN(n10706) );
  OAI21_X1 U12580 ( .B1(n15982), .B2(n15667), .A(n10706), .ZN(n10716) );
  NOR2_X1 U12581 ( .A1(n10708), .A2(n10707), .ZN(n10710) );
  NAND2_X1 U12582 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n10958), .ZN(n10711) );
  OAI21_X1 U12583 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n10958), .A(n10711), .ZN(
        n10712) );
  AOI21_X1 U12584 ( .B1(n10713), .B2(n10712), .A(n10957), .ZN(n10714) );
  NOR2_X1 U12585 ( .A1(n10714), .A2(n15999), .ZN(n10715) );
  AOI211_X1 U12586 ( .C1(n13713), .C2(n10717), .A(n10716), .B(n10715), .ZN(
        n10718) );
  OAI211_X1 U12587 ( .C1(n10720), .C2(n15993), .A(n10719), .B(n10718), .ZN(
        P3_U3190) );
  NAND2_X1 U12588 ( .A1(n10721), .A2(n7644), .ZN(n10725) );
  OR2_X1 U12589 ( .A1(n12316), .A2(n10722), .ZN(n10724) );
  OR2_X1 U12590 ( .A1(n7433), .A2(n8047), .ZN(n10723) );
  OAI22_X1 U12591 ( .A1(n12561), .A2(n10228), .B1(n11965), .B2(n16162), .ZN(
        n10726) );
  XNOR2_X1 U12592 ( .A(n10726), .B(n12518), .ZN(n10970) );
  OAI22_X1 U12593 ( .A1(n12483), .A2(n12561), .B1(n16162), .B2(n10228), .ZN(
        n10969) );
  XNOR2_X1 U12594 ( .A(n10970), .B(n10969), .ZN(n10737) );
  INV_X1 U12595 ( .A(n10729), .ZN(n10730) );
  NAND2_X1 U12596 ( .A1(n10731), .A2(n10730), .ZN(n10732) );
  INV_X1 U12597 ( .A(n10972), .ZN(n10735) );
  AOI211_X1 U12598 ( .C1(n10737), .C2(n10736), .A(n14829), .B(n10735), .ZN(
        n10749) );
  INV_X1 U12599 ( .A(n14811), .ZN(n14824) );
  AOI22_X1 U12600 ( .A1(n14824), .A2(n10739), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_STATE_REG_SCAN_IN), .ZN(n10748) );
  NAND2_X1 U12601 ( .A1(n7427), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10744) );
  NAND2_X1 U12602 ( .A1(n12524), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10743) );
  NOR2_X1 U12603 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n10740) );
  NOR2_X1 U12604 ( .A1(n10873), .A2(n10740), .ZN(n11102) );
  NAND2_X1 U12605 ( .A1(n12526), .A2(n11102), .ZN(n10742) );
  NAND2_X1 U12606 ( .A1(n12686), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n10741) );
  NAND2_X1 U12607 ( .A1(n14857), .A2(n14807), .ZN(n10745) );
  OAI21_X1 U12608 ( .B1(n10860), .B2(n14785), .A(n10745), .ZN(n16139) );
  INV_X1 U12609 ( .A(n16139), .ZN(n10746) );
  OAI22_X1 U12610 ( .A1(n14804), .A2(n16162), .B1(n10746), .B2(n14809), .ZN(
        n10747) );
  OR3_X1 U12611 ( .A1(n10749), .A2(n10748), .A3(n10747), .ZN(P1_U3218) );
  INV_X1 U12612 ( .A(n10773), .ZN(n10778) );
  NOR2_X1 U12613 ( .A1(n10777), .A2(n10774), .ZN(n10750) );
  AOI21_X1 U12614 ( .B1(n10751), .B2(n10778), .A(n10750), .ZN(n10755) );
  MUX2_X1 U12615 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n12298), .Z(n10752) );
  NAND2_X1 U12616 ( .A1(n10752), .A2(SI_17_), .ZN(n10781) );
  INV_X1 U12617 ( .A(n10752), .ZN(n10753) );
  NAND2_X1 U12618 ( .A1(n10753), .A2(n15477), .ZN(n10779) );
  AND2_X1 U12619 ( .A1(n10781), .A2(n10779), .ZN(n10754) );
  XNOR2_X1 U12620 ( .A(n10755), .B(n10754), .ZN(n12248) );
  INV_X1 U12621 ( .A(n12248), .ZN(n10760) );
  NAND2_X1 U12622 ( .A1(n10757), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10756) );
  MUX2_X1 U12623 ( .A(n10756), .B(P1_IR_REG_31__SCAN_IN), .S(n15649), .Z(
        n10758) );
  NAND2_X1 U12624 ( .A1(n10758), .A2(n10818), .ZN(n11751) );
  OAI222_X1 U12625 ( .A1(n15262), .A2(n10759), .B1(n15260), .B2(n10760), .C1(
        P1_U3086), .C2(n11751), .ZN(P1_U3338) );
  XNOR2_X1 U12626 ( .A(n10827), .B(P2_IR_REG_17__SCAN_IN), .ZN(n14288) );
  INV_X1 U12627 ( .A(n14288), .ZN(n14281) );
  OAI222_X1 U12628 ( .A1(n14693), .A2(n10761), .B1(n14691), .B2(n10760), .C1(
        P2_U3088), .C2(n14281), .ZN(P2_U3310) );
  NAND2_X1 U12629 ( .A1(n10762), .A2(n16052), .ZN(n10764) );
  AND2_X1 U12630 ( .A1(n10766), .A2(n10764), .ZN(n10768) );
  XNOR2_X1 U12631 ( .A(n11027), .B(n13621), .ZN(n10767) );
  AND2_X1 U12632 ( .A1(n10767), .A2(n10764), .ZN(n10765) );
  OAI211_X1 U12633 ( .C1(n10768), .C2(n10767), .A(n13587), .B(n11030), .ZN(
        n10772) );
  OAI22_X1 U12634 ( .A1(n13575), .A2(n11209), .B1(n16052), .B2(n13600), .ZN(
        n10769) );
  AOI211_X1 U12635 ( .C1(n13606), .C2(n11329), .A(n10770), .B(n10769), .ZN(
        n10771) );
  OAI211_X1 U12636 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n13604), .A(n10772), .B(
        n10771), .ZN(P3_U3158) );
  OAI21_X1 U12637 ( .B1(n10774), .B2(n10773), .A(n10781), .ZN(n10775) );
  INV_X1 U12638 ( .A(n10775), .ZN(n10776) );
  NOR2_X1 U12639 ( .A1(n10778), .A2(SI_16_), .ZN(n10782) );
  INV_X1 U12640 ( .A(n10779), .ZN(n10780) );
  AOI21_X1 U12641 ( .B1(n10782), .B2(n10781), .A(n10780), .ZN(n10783) );
  MUX2_X1 U12642 ( .A(n10825), .B(n10830), .S(n8006), .Z(n10824) );
  MUX2_X1 U12643 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n8006), .Z(n10786) );
  NAND2_X1 U12644 ( .A1(n10786), .A2(SI_19_), .ZN(n11006) );
  OAI21_X1 U12645 ( .B1(n11001), .B2(n10824), .A(n11006), .ZN(n10784) );
  INV_X1 U12646 ( .A(n10784), .ZN(n10785) );
  INV_X1 U12647 ( .A(n10824), .ZN(n10999) );
  NOR2_X1 U12648 ( .A1(n10999), .A2(SI_18_), .ZN(n10789) );
  INV_X1 U12649 ( .A(n10786), .ZN(n10787) );
  NAND2_X1 U12650 ( .A1(n10787), .A2(n15473), .ZN(n11005) );
  INV_X1 U12651 ( .A(n11005), .ZN(n10788) );
  AOI21_X1 U12652 ( .B1(n10789), .B2(n11006), .A(n10788), .ZN(n10790) );
  MUX2_X1 U12653 ( .A(n12336), .B(n13096), .S(n8006), .Z(n10911) );
  XNOR2_X1 U12654 ( .A(n10911), .B(SI_20_), .ZN(n10792) );
  XNOR2_X1 U12655 ( .A(n10912), .B(n10792), .ZN(n13095) );
  INV_X1 U12656 ( .A(n13095), .ZN(n10833) );
  OAI222_X1 U12657 ( .A1(n14693), .A2(n13096), .B1(P2_U3088), .B2(n10793), 
        .C1(n10833), .C2(n14691), .ZN(P2_U3307) );
  NAND2_X1 U12658 ( .A1(n13178), .A2(n10794), .ZN(n10795) );
  NAND2_X1 U12659 ( .A1(n11362), .A2(n9720), .ZN(n10799) );
  AOI22_X1 U12660 ( .A1(n10797), .A2(n13109), .B1(n9659), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n10798) );
  INV_X1 U12661 ( .A(n14258), .ZN(n13185) );
  XNOR2_X1 U12662 ( .A(n13183), .B(n13185), .ZN(n13433) );
  INV_X1 U12663 ( .A(n13433), .ZN(n11246) );
  XNOR2_X1 U12664 ( .A(n11247), .B(n11246), .ZN(n10812) );
  NAND2_X1 U12665 ( .A1(n9742), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10805) );
  AND2_X1 U12666 ( .A1(n10800), .A2(n11151), .ZN(n10801) );
  NOR2_X1 U12667 ( .A1(n11144), .A2(n10801), .ZN(n16302) );
  NAND2_X1 U12668 ( .A1(n11931), .A2(n16302), .ZN(n10804) );
  NAND2_X1 U12669 ( .A1(n13386), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n10803) );
  NAND2_X1 U12670 ( .A1(n13368), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10802) );
  NAND4_X1 U12671 ( .A1(n10805), .A2(n10804), .A3(n10803), .A4(n10802), .ZN(
        n14257) );
  NAND2_X1 U12672 ( .A1(n14257), .A2(n14439), .ZN(n10807) );
  NAND2_X1 U12673 ( .A1(n14259), .A2(n14438), .ZN(n10806) );
  NAND2_X1 U12674 ( .A1(n10807), .A2(n10806), .ZN(n10924) );
  NAND2_X1 U12675 ( .A1(n13178), .A2(n14259), .ZN(n10808) );
  OR2_X1 U12676 ( .A1(n10809), .A2(n13433), .ZN(n10810) );
  NAND2_X1 U12677 ( .A1(n11266), .A2(n10810), .ZN(n11159) );
  NOR2_X1 U12678 ( .A1(n11159), .A2(n12045), .ZN(n10811) );
  AOI211_X1 U12679 ( .C1(n14529), .C2(n10812), .A(n10924), .B(n10811), .ZN(
        n11158) );
  AOI211_X1 U12680 ( .C1(n13183), .C2(n10813), .A(n14445), .B(n11282), .ZN(
        n11156) );
  INV_X1 U12681 ( .A(n13183), .ZN(n10931) );
  AOI22_X1 U12682 ( .A1(n16405), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n10928), 
        .B2(n16394), .ZN(n10814) );
  OAI21_X1 U12683 ( .B1(n10931), .B2(n16398), .A(n10814), .ZN(n10816) );
  NOR2_X1 U12684 ( .A1(n11159), .A2(n14452), .ZN(n10815) );
  AOI211_X1 U12685 ( .C1(n11156), .C2(n16306), .A(n10816), .B(n10815), .ZN(
        n10817) );
  OAI21_X1 U12686 ( .B1(n11158), .B2(n16405), .A(n10817), .ZN(P2_U3256) );
  NAND2_X1 U12687 ( .A1(n10818), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10819) );
  MUX2_X1 U12688 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10819), .S(
        P1_IR_REG_18__SCAN_IN), .Z(n10820) );
  INV_X1 U12689 ( .A(n10820), .ZN(n10823) );
  NOR2_X1 U12690 ( .A1(n10823), .A2(n10822), .ZN(n12351) );
  INV_X1 U12691 ( .A(n12351), .ZN(n11759) );
  XNOR2_X1 U12692 ( .A(n11002), .B(SI_18_), .ZN(n11000) );
  XNOR2_X1 U12693 ( .A(n11000), .B(n10824), .ZN(n12350) );
  INV_X1 U12694 ( .A(n12350), .ZN(n10831) );
  OAI222_X1 U12695 ( .A1(P1_U3086), .A2(n11759), .B1(n15260), .B2(n10831), 
        .C1(n10825), .C2(n15262), .ZN(P1_U3337) );
  INV_X1 U12696 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n10826) );
  NAND2_X1 U12697 ( .A1(n10827), .A2(n10826), .ZN(n10828) );
  NAND2_X1 U12698 ( .A1(n10828), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10829) );
  XNOR2_X1 U12699 ( .A(n10829), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14286) );
  INV_X1 U12700 ( .A(n14286), .ZN(n14294) );
  OAI222_X1 U12701 ( .A1(P2_U3088), .A2(n14294), .B1(n14691), .B2(n10831), 
        .C1(n10830), .C2(n14693), .ZN(P2_U3309) );
  NAND2_X1 U12702 ( .A1(n13623), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n10832) );
  OAI21_X1 U12703 ( .B1(n13025), .B2(n13623), .A(n10832), .ZN(P3_U3521) );
  OAI222_X1 U12704 ( .A1(n15262), .A2(n12336), .B1(P1_U3086), .B2(n16039), 
        .C1(n15260), .C2(n10833), .ZN(P1_U3335) );
  INV_X1 U12705 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10835) );
  MUX2_X1 U12706 ( .A(n10835), .B(P2_REG2_REG_11__SCAN_IN), .S(n11243), .Z(
        n10836) );
  INV_X1 U12707 ( .A(n10836), .ZN(n10837) );
  NAND2_X1 U12708 ( .A1(n10838), .A2(n10837), .ZN(n11078) );
  OAI21_X1 U12709 ( .B1(n10838), .B2(n10837), .A(n11078), .ZN(n10848) );
  NAND2_X1 U12710 ( .A1(n15838), .A2(n11243), .ZN(n10841) );
  NAND2_X1 U12711 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n10840)
         );
  NAND2_X1 U12712 ( .A1(n15800), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n10839) );
  NAND3_X1 U12713 ( .A1(n10841), .A2(n10840), .A3(n10839), .ZN(n10847) );
  INV_X1 U12714 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10843) );
  MUX2_X1 U12715 ( .A(n10843), .B(P2_REG1_REG_11__SCAN_IN), .S(n11243), .Z(
        n10844) );
  AOI211_X1 U12716 ( .C1(n10845), .C2(n10844), .A(n15813), .B(n11070), .ZN(
        n10846) );
  AOI211_X1 U12717 ( .C1(n15830), .C2(n10848), .A(n10847), .B(n10846), .ZN(
        n10849) );
  INV_X1 U12718 ( .A(n10849), .ZN(P2_U3225) );
  INV_X1 U12719 ( .A(SI_23_), .ZN(n10852) );
  NAND2_X1 U12720 ( .A1(n10850), .A2(n16291), .ZN(n10851) );
  OAI211_X1 U12721 ( .C1(n10852), .C2(n13462), .A(n10851), .B(n13043), .ZN(
        P3_U3272) );
  INV_X1 U12722 ( .A(n10853), .ZN(n13080) );
  NOR2_X1 U12723 ( .A1(n13080), .A2(n10854), .ZN(n10856) );
  INV_X1 U12724 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10907) );
  NAND2_X1 U12725 ( .A1(n10860), .A2(n10859), .ZN(n10861) );
  XNOR2_X1 U12726 ( .A(n14858), .B(n16143), .ZN(n16137) );
  INV_X1 U12727 ( .A(n16137), .ZN(n10862) );
  NAND2_X1 U12728 ( .A1(n16136), .A2(n10862), .ZN(n10864) );
  NAND2_X1 U12729 ( .A1(n12561), .A2(n16162), .ZN(n10863) );
  INV_X1 U12730 ( .A(n14857), .ZN(n12542) );
  NAND2_X1 U12731 ( .A1(n10865), .A2(n12491), .ZN(n10867) );
  AOI22_X1 U12733 ( .A1(n12399), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n12398), 
        .B2(n16003), .ZN(n10866) );
  NAND2_X1 U12734 ( .A1(n10867), .A2(n10866), .ZN(n12544) );
  NAND2_X1 U12735 ( .A1(n10869), .A2(n12491), .ZN(n10872) );
  AOI22_X1 U12736 ( .A1(n12399), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n12398), 
        .B2(n10870), .ZN(n10871) );
  NAND2_X1 U12737 ( .A1(n10872), .A2(n10871), .ZN(n12570) );
  NAND2_X1 U12738 ( .A1(n7426), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10877) );
  NAND2_X1 U12739 ( .A1(n12524), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n10876) );
  NAND2_X1 U12740 ( .A1(n10873), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10884) );
  OAI21_X1 U12741 ( .B1(n10873), .B2(P1_REG3_REG_5__SCAN_IN), .A(n10884), .ZN(
        n11022) );
  INV_X1 U12742 ( .A(n11022), .ZN(n10993) );
  NAND2_X1 U12743 ( .A1(n12526), .A2(n10993), .ZN(n10875) );
  NAND2_X1 U12744 ( .A1(n12686), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n10874) );
  INV_X1 U12745 ( .A(n12570), .ZN(n16208) );
  INV_X1 U12746 ( .A(n14856), .ZN(n11016) );
  NAND2_X1 U12747 ( .A1(n16208), .A2(n11016), .ZN(n10878) );
  NAND2_X1 U12748 ( .A1(n10879), .A2(n12491), .ZN(n10882) );
  AOI22_X1 U12749 ( .A1(n12399), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n12398), 
        .B2(n10880), .ZN(n10881) );
  NAND2_X1 U12750 ( .A1(n10882), .A2(n10881), .ZN(n12575) );
  NAND2_X1 U12751 ( .A1(n7427), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10889) );
  NAND2_X1 U12752 ( .A1(n12524), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10888) );
  NOR2_X1 U12753 ( .A1(n10884), .A2(n10883), .ZN(n10896) );
  AND2_X1 U12754 ( .A1(n10884), .A2(n10883), .ZN(n10885) );
  NOR2_X1 U12755 ( .A1(n10896), .A2(n10885), .ZN(n11177) );
  NAND2_X1 U12756 ( .A1(n12526), .A2(n11177), .ZN(n10887) );
  NAND2_X1 U12757 ( .A1(n12686), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n10886) );
  NAND4_X1 U12758 ( .A1(n10889), .A2(n10888), .A3(n10887), .A4(n10886), .ZN(
        n14855) );
  XNOR2_X1 U12759 ( .A(n12575), .B(n14855), .ZN(n12728) );
  OAI21_X1 U12760 ( .B1(n10890), .B2(n8337), .A(n11044), .ZN(n10904) );
  INV_X1 U12761 ( .A(n10904), .ZN(n10943) );
  NAND2_X1 U12762 ( .A1(n14858), .A2(n16162), .ZN(n10892) );
  INV_X2 U12763 ( .A(n12544), .ZN(n16189) );
  AND2_X1 U12764 ( .A1(n14857), .A2(n16189), .ZN(n10893) );
  OAI22_X1 U12765 ( .A1(n11106), .A2(n10893), .B1(n16189), .B2(n14857), .ZN(
        n10982) );
  NAND2_X1 U12766 ( .A1(n10982), .A2(n12566), .ZN(n10895) );
  NAND2_X1 U12767 ( .A1(n11016), .A2(n12570), .ZN(n10894) );
  NAND2_X1 U12768 ( .A1(n10895), .A2(n10894), .ZN(n11049) );
  XNOR2_X1 U12769 ( .A(n11049), .B(n8337), .ZN(n10902) );
  NAND2_X1 U12770 ( .A1(n7426), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10901) );
  NAND2_X1 U12771 ( .A1(n12524), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10900) );
  NAND2_X1 U12772 ( .A1(n10896), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n11054) );
  OR2_X1 U12773 ( .A1(n10896), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10897) );
  AND2_X1 U12774 ( .A1(n11054), .A2(n10897), .ZN(n16239) );
  NAND2_X1 U12775 ( .A1(n12526), .A2(n16239), .ZN(n10899) );
  NAND2_X1 U12776 ( .A1(n12686), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n10898) );
  NAND4_X1 U12777 ( .A1(n10901), .A2(n10900), .A3(n10899), .A4(n10898), .ZN(
        n14854) );
  AOI22_X1 U12778 ( .A1(n14807), .A2(n14854), .B1(n14856), .B2(n14806), .ZN(
        n11180) );
  OAI21_X1 U12779 ( .B1(n10902), .B2(n16379), .A(n11180), .ZN(n10903) );
  AOI21_X1 U12780 ( .B1(n16372), .B2(n10904), .A(n10903), .ZN(n10935) );
  AOI211_X1 U12781 ( .C1(n12575), .C2(n10991), .A(n16142), .B(n11062), .ZN(
        n10940) );
  AOI21_X1 U12782 ( .B1(n16366), .B2(n12575), .A(n10940), .ZN(n10905) );
  OAI211_X1 U12783 ( .C1(n10943), .C2(n16369), .A(n10935), .B(n10905), .ZN(
        n10908) );
  NAND2_X1 U12784 ( .A1(n10908), .A2(n16391), .ZN(n10906) );
  OAI21_X1 U12785 ( .B1(n16391), .B2(n10907), .A(n10906), .ZN(P1_U3477) );
  NAND2_X1 U12786 ( .A1(n10908), .A2(n16387), .ZN(n10909) );
  OAI21_X1 U12787 ( .B1(n16387), .B2(n10910), .A(n10909), .ZN(P1_U3534) );
  MUX2_X1 U12788 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n8006), .Z(n10913) );
  NAND2_X1 U12789 ( .A1(n10913), .A2(SI_21_), .ZN(n11320) );
  OAI21_X1 U12790 ( .B1(SI_21_), .B2(n10913), .A(n11320), .ZN(n10914) );
  NAND2_X1 U12791 ( .A1(n10915), .A2(n10914), .ZN(n10916) );
  NAND2_X1 U12792 ( .A1(n11321), .A2(n10916), .ZN(n13248) );
  INV_X1 U12793 ( .A(n13350), .ZN(n13451) );
  OAI222_X1 U12794 ( .A1(n14693), .A2(n13249), .B1(n14691), .B2(n13248), .C1(
        n13451), .C2(P2_U3088), .ZN(P2_U3306) );
  XNOR2_X1 U12795 ( .A(n13183), .B(n11516), .ZN(n11139) );
  NAND2_X1 U12796 ( .A1(n14258), .A2(n14445), .ZN(n11137) );
  XNOR2_X1 U12797 ( .A(n11139), .B(n11137), .ZN(n10922) );
  INV_X1 U12798 ( .A(n10917), .ZN(n10920) );
  OAI21_X1 U12799 ( .B1(n10920), .B2(n10919), .A(n10918), .ZN(n10921) );
  NAND2_X1 U12800 ( .A1(n10921), .A2(n10922), .ZN(n11138) );
  OAI21_X1 U12801 ( .B1(n10922), .B2(n10921), .A(n11138), .ZN(n10923) );
  NAND2_X1 U12802 ( .A1(n10923), .A2(n14232), .ZN(n10930) );
  INV_X1 U12803 ( .A(n10924), .ZN(n10926) );
  OAI22_X1 U12804 ( .A1(n14244), .A2(n10926), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10925), .ZN(n10927) );
  AOI21_X1 U12805 ( .B1(n10928), .B2(n14242), .A(n10927), .ZN(n10929) );
  OAI211_X1 U12806 ( .C1(n10931), .C2(n12244), .A(n10930), .B(n10929), .ZN(
        P2_U3203) );
  OR2_X1 U12807 ( .A1(n13081), .A2(n13080), .ZN(n10932) );
  NAND2_X1 U12808 ( .A1(n10933), .A2(n16038), .ZN(n12718) );
  INV_X1 U12809 ( .A(n12718), .ZN(n10934) );
  NAND2_X1 U12810 ( .A1(n16086), .A2(n10934), .ZN(n16045) );
  MUX2_X1 U12811 ( .A(n9998), .B(n10935), .S(n16159), .Z(n10942) );
  INV_X1 U12812 ( .A(n12575), .ZN(n10938) );
  INV_X1 U12813 ( .A(n11177), .ZN(n10937) );
  OAI22_X1 U12814 ( .A1(n16163), .A2(n10938), .B1(n10937), .B2(n16161), .ZN(
        n10939) );
  AOI21_X1 U12815 ( .B1(n16341), .B2(n10940), .A(n10939), .ZN(n10941) );
  OAI211_X1 U12816 ( .C1(n10943), .C2(n16045), .A(n10942), .B(n10941), .ZN(
        P1_U3287) );
  OAI222_X1 U12817 ( .A1(n15262), .A2(n12325), .B1(P1_U3086), .B2(n10944), 
        .C1(n15260), .C2(n13248), .ZN(P1_U3334) );
  INV_X1 U12818 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n16278) );
  AOI21_X1 U12819 ( .B1(n16278), .B2(n10946), .A(n11110), .ZN(n10967) );
  INV_X1 U12820 ( .A(n10947), .ZN(n10953) );
  INV_X1 U12821 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n10948) );
  NAND2_X1 U12822 ( .A1(n10949), .A2(n11121), .ZN(n11114) );
  INV_X1 U12823 ( .A(n10949), .ZN(n10950) );
  NAND2_X1 U12824 ( .A1(n10950), .A2(n10959), .ZN(n10951) );
  AND2_X1 U12825 ( .A1(n11114), .A2(n10951), .ZN(n10952) );
  INV_X1 U12826 ( .A(n11115), .ZN(n10956) );
  NOR3_X1 U12827 ( .A1(n10954), .A2(n10953), .A3(n10952), .ZN(n10955) );
  OAI21_X1 U12828 ( .B1(n10956), .B2(n10955), .A(n15970), .ZN(n10966) );
  AOI21_X1 U12829 ( .B1(n10948), .B2(n10960), .A(n11122), .ZN(n10963) );
  NOR2_X1 U12830 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15536), .ZN(n11862) );
  AOI21_X1 U12831 ( .B1(n15961), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n11862), .ZN(
        n10962) );
  NAND2_X1 U12832 ( .A1(n13713), .A2(n11121), .ZN(n10961) );
  OAI211_X1 U12833 ( .C1(n10963), .C2(n15999), .A(n10962), .B(n10961), .ZN(
        n10964) );
  INV_X1 U12834 ( .A(n10964), .ZN(n10965) );
  OAI211_X1 U12835 ( .C1(n10967), .C2(n15993), .A(n10966), .B(n10965), .ZN(
        P3_U3191) );
  OAI22_X1 U12836 ( .A1(n12542), .A2(n10228), .B1(n8012), .B2(n16189), .ZN(
        n10968) );
  XNOR2_X1 U12837 ( .A(n10968), .B(n12518), .ZN(n11012) );
  NAND2_X1 U12838 ( .A1(n10970), .A2(n10969), .ZN(n10971) );
  OAI22_X1 U12839 ( .A1(n12483), .A2(n12542), .B1(n16189), .B2(n10228), .ZN(
        n10974) );
  NAND2_X1 U12840 ( .A1(n11013), .A2(n11014), .ZN(n10976) );
  XOR2_X1 U12841 ( .A(n11012), .B(n10976), .Z(n10981) );
  NAND2_X1 U12842 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n16025) );
  NAND2_X1 U12843 ( .A1(n14856), .A2(n14807), .ZN(n10977) );
  OAI21_X1 U12844 ( .B1(n12561), .B2(n14785), .A(n10977), .ZN(n16186) );
  NAND2_X1 U12845 ( .A1(n14821), .A2(n16186), .ZN(n10978) );
  OAI211_X1 U12846 ( .C1(n14804), .C2(n16189), .A(n16025), .B(n10978), .ZN(
        n10979) );
  AOI21_X1 U12847 ( .B1(n11102), .B2(n14811), .A(n10979), .ZN(n10980) );
  OAI21_X1 U12848 ( .B1(n10981), .B2(n14829), .A(n10980), .ZN(P1_U3230) );
  XNOR2_X1 U12849 ( .A(n10982), .B(n8675), .ZN(n10989) );
  NAND2_X1 U12850 ( .A1(n10984), .A2(n10983), .ZN(n16211) );
  NAND2_X1 U12851 ( .A1(n16211), .A2(n16372), .ZN(n10988) );
  NAND2_X1 U12852 ( .A1(n14855), .A2(n14807), .ZN(n10986) );
  NAND2_X1 U12853 ( .A1(n14857), .A2(n14806), .ZN(n10985) );
  NAND2_X1 U12854 ( .A1(n10986), .A2(n10985), .ZN(n11019) );
  INV_X1 U12855 ( .A(n11019), .ZN(n10987) );
  OAI211_X1 U12856 ( .C1(n10989), .C2(n16379), .A(n10988), .B(n10987), .ZN(
        n16209) );
  MUX2_X1 U12857 ( .A(n16209), .B(P1_REG2_REG_5__SCAN_IN), .S(n16347), .Z(
        n10990) );
  INV_X1 U12858 ( .A(n10990), .ZN(n10998) );
  INV_X1 U12859 ( .A(n16045), .ZN(n16342) );
  AOI21_X1 U12860 ( .B1(n11101), .B2(n12570), .A(n16142), .ZN(n10992) );
  AND2_X1 U12861 ( .A1(n10992), .A2(n10991), .ZN(n16206) );
  NAND2_X1 U12862 ( .A1(n16341), .A2(n16206), .ZN(n10995) );
  INV_X1 U12863 ( .A(n16161), .ZN(n16336) );
  NAND2_X1 U12864 ( .A1(n16336), .A2(n10993), .ZN(n10994) );
  OAI211_X1 U12865 ( .C1(n16208), .C2(n16163), .A(n10995), .B(n10994), .ZN(
        n10996) );
  AOI21_X1 U12866 ( .B1(n16211), .B2(n16342), .A(n10996), .ZN(n10997) );
  NAND2_X1 U12867 ( .A1(n10998), .A2(n10997), .ZN(P1_U3288) );
  NAND2_X1 U12868 ( .A1(n11000), .A2(n10999), .ZN(n11004) );
  OR2_X1 U12869 ( .A1(n11002), .A2(n11001), .ZN(n11003) );
  NAND2_X1 U12870 ( .A1(n11004), .A2(n11003), .ZN(n11008) );
  NAND2_X1 U12871 ( .A1(n11006), .A2(n11005), .ZN(n11007) );
  INV_X1 U12872 ( .A(n13108), .ZN(n11010) );
  OAI222_X1 U12873 ( .A1(n14693), .A2(n11009), .B1(n14691), .B2(n11010), .C1(
        P2_U3088), .C2(n9660), .ZN(P2_U3308) );
  INV_X1 U12874 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11011) );
  OAI222_X1 U12875 ( .A1(n15262), .A2(n11011), .B1(n15260), .B2(n11010), .C1(
        n12752), .C2(P1_U3086), .ZN(P1_U3336) );
  NAND2_X1 U12876 ( .A1(n11013), .A2(n11012), .ZN(n11015) );
  OAI22_X1 U12877 ( .A1(n12483), .A2(n11016), .B1(n16208), .B2(n10228), .ZN(
        n11172) );
  OAI22_X1 U12878 ( .A1(n16208), .A2(n8012), .B1(n10228), .B2(n11016), .ZN(
        n11017) );
  XNOR2_X1 U12879 ( .A(n11017), .B(n12518), .ZN(n11173) );
  XOR2_X1 U12880 ( .A(n11172), .B(n11173), .Z(n11018) );
  NAND2_X1 U12881 ( .A1(n14821), .A2(n11019), .ZN(n11020) );
  OAI211_X1 U12882 ( .C1(n14824), .C2(n11022), .A(n11021), .B(n11020), .ZN(
        n11023) );
  AOI21_X1 U12883 ( .B1(n12570), .B2(n14826), .A(n11023), .ZN(n11024) );
  OAI21_X1 U12884 ( .B1(n11025), .B2(n14829), .A(n11024), .ZN(P1_U3227) );
  NAND2_X1 U12885 ( .A1(n13623), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n11026) );
  OAI21_X1 U12886 ( .B1(n13776), .B2(n13623), .A(n11026), .ZN(P3_U3519) );
  INV_X1 U12887 ( .A(n11027), .ZN(n11028) );
  NAND2_X1 U12888 ( .A1(n11028), .A2(n13621), .ZN(n11029) );
  XNOR2_X1 U12889 ( .A(n12881), .B(n12836), .ZN(n11031) );
  NAND2_X1 U12890 ( .A1(n11031), .A2(n11209), .ZN(n11204) );
  INV_X1 U12891 ( .A(n11031), .ZN(n11032) );
  NAND2_X1 U12892 ( .A1(n11032), .A2(n13620), .ZN(n11033) );
  NAND2_X1 U12893 ( .A1(n11204), .A2(n11033), .ZN(n11035) );
  INV_X1 U12894 ( .A(n11205), .ZN(n11034) );
  AOI21_X1 U12895 ( .B1(n11036), .B2(n11035), .A(n11034), .ZN(n11042) );
  OAI22_X1 U12896 ( .A1(n13575), .A2(n11306), .B1(n16102), .B2(n13600), .ZN(
        n11037) );
  AOI211_X1 U12897 ( .C1(n13606), .C2(n16182), .A(n11038), .B(n11037), .ZN(
        n11041) );
  INV_X1 U12898 ( .A(n11039), .ZN(n11224) );
  NAND2_X1 U12899 ( .A1(n13568), .A2(n11224), .ZN(n11040) );
  OAI211_X1 U12900 ( .C1(n11042), .C2(n13608), .A(n11041), .B(n11040), .ZN(
        P3_U3170) );
  INV_X1 U12901 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n11067) );
  OR2_X1 U12902 ( .A1(n12575), .A2(n14855), .ZN(n11043) );
  NAND2_X1 U12903 ( .A1(n11044), .A2(n11043), .ZN(n11048) );
  NAND2_X1 U12904 ( .A1(n11045), .A2(n12491), .ZN(n11047) );
  AOI22_X1 U12905 ( .A1(n12399), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n12398), 
        .B2(n14883), .ZN(n11046) );
  NAND2_X1 U12906 ( .A1(n11047), .A2(n11046), .ZN(n16240) );
  XNOR2_X1 U12907 ( .A(n16240), .B(n14854), .ZN(n12729) );
  NAND2_X1 U12908 ( .A1(n11048), .A2(n11052), .ZN(n11373) );
  OAI21_X1 U12909 ( .B1(n11048), .B2(n11052), .A(n11373), .ZN(n16242) );
  INV_X1 U12910 ( .A(n16242), .ZN(n11065) );
  INV_X1 U12911 ( .A(n14855), .ZN(n11050) );
  NAND2_X1 U12912 ( .A1(n12575), .A2(n11050), .ZN(n11051) );
  XNOR2_X1 U12913 ( .A(n11355), .B(n11052), .ZN(n11060) );
  NAND2_X1 U12914 ( .A1(n7426), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n11059) );
  NAND2_X1 U12915 ( .A1(n12524), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n11058) );
  INV_X1 U12916 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n11053) );
  NAND2_X1 U12917 ( .A1(n11054), .A2(n11053), .ZN(n11055) );
  AND2_X1 U12918 ( .A1(n11366), .A2(n11055), .ZN(n11492) );
  NAND2_X1 U12919 ( .A1(n12526), .A2(n11492), .ZN(n11057) );
  NAND2_X1 U12920 ( .A1(n12686), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n11056) );
  NAND4_X1 U12921 ( .A1(n11059), .A2(n11058), .A3(n11057), .A4(n11056), .ZN(
        n14853) );
  AOI22_X1 U12922 ( .A1(n14807), .A2(n14853), .B1(n14855), .B2(n14806), .ZN(
        n11239) );
  OAI21_X1 U12923 ( .B1(n11060), .B2(n16379), .A(n11239), .ZN(n11061) );
  AOI21_X1 U12924 ( .B1(n16372), .B2(n16242), .A(n11061), .ZN(n16245) );
  INV_X1 U12925 ( .A(n11062), .ZN(n11063) );
  AOI211_X1 U12926 ( .C1(n16240), .C2(n11063), .A(n16142), .B(n11398), .ZN(
        n16241) );
  AOI21_X1 U12927 ( .B1(n16366), .B2(n16240), .A(n16241), .ZN(n11064) );
  OAI211_X1 U12928 ( .C1(n11065), .C2(n16369), .A(n16245), .B(n11064), .ZN(
        n11068) );
  NAND2_X1 U12929 ( .A1(n11068), .A2(n16391), .ZN(n11066) );
  OAI21_X1 U12930 ( .B1(n16391), .B2(n11067), .A(n11066), .ZN(P1_U3480) );
  NAND2_X1 U12931 ( .A1(n11068), .A2(n16387), .ZN(n11069) );
  OAI21_X1 U12932 ( .B1(n16387), .B2(n14884), .A(n11069), .ZN(P1_U3535) );
  INV_X1 U12933 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11071) );
  MUX2_X1 U12934 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n11071), .S(n11431), .Z(
        n11072) );
  OAI21_X1 U12935 ( .B1(n11073), .B2(n11072), .A(n11425), .ZN(n11077) );
  NAND2_X1 U12936 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n11520)
         );
  NAND2_X1 U12937 ( .A1(n15800), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n11074) );
  OAI211_X1 U12938 ( .C1(n14306), .C2(n11075), .A(n11520), .B(n11074), .ZN(
        n11076) );
  AOI21_X1 U12939 ( .B1(n11077), .B2(n15835), .A(n11076), .ZN(n11083) );
  XOR2_X1 U12940 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n11431), .Z(n11080) );
  OAI21_X1 U12941 ( .B1(n11243), .B2(P2_REG2_REG_11__SCAN_IN), .A(n11078), 
        .ZN(n11079) );
  NAND2_X1 U12942 ( .A1(n11079), .A2(n11080), .ZN(n11430) );
  OAI21_X1 U12943 ( .B1(n11080), .B2(n11079), .A(n11430), .ZN(n11081) );
  NAND2_X1 U12944 ( .A1(n11081), .A2(n15830), .ZN(n11082) );
  NAND2_X1 U12945 ( .A1(n11083), .A2(n11082), .ZN(P2_U3226) );
  NAND2_X1 U12946 ( .A1(n11085), .A2(n11084), .ZN(n11088) );
  NAND2_X1 U12947 ( .A1(n14108), .A2(n11086), .ZN(n11087) );
  NAND2_X1 U12948 ( .A1(n11090), .A2(n11089), .ZN(n11094) );
  NAND2_X1 U12949 ( .A1(n11092), .A2(n16121), .ZN(n11096) );
  NAND2_X1 U12950 ( .A1(n16200), .A2(n11093), .ZN(n16115) );
  INV_X1 U12951 ( .A(n13963), .ZN(n13933) );
  AOI22_X1 U12952 ( .A1(n13933), .A2(n16055), .B1(n13868), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n11095) );
  OAI211_X1 U12953 ( .C1(n8388), .C2(n16121), .A(n11096), .B(n11095), .ZN(
        P3_U3233) );
  XNOR2_X1 U12954 ( .A(n14857), .B(n12544), .ZN(n12565) );
  XNOR2_X1 U12955 ( .A(n11097), .B(n12565), .ZN(n16191) );
  INV_X1 U12956 ( .A(n11098), .ZN(n11099) );
  OR2_X1 U12957 ( .A1(n16141), .A2(n16189), .ZN(n11100) );
  AND3_X1 U12958 ( .A1(n11101), .A2(n11100), .A3(n16322), .ZN(n16185) );
  MUX2_X1 U12959 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n16186), .S(n16159), .Z(
        n11105) );
  INV_X1 U12960 ( .A(n11102), .ZN(n11103) );
  OAI22_X1 U12961 ( .A1(n16163), .A2(n16189), .B1(n16161), .B2(n11103), .ZN(
        n11104) );
  AOI211_X1 U12962 ( .C1(n16185), .C2(n16341), .A(n11105), .B(n11104), .ZN(
        n11108) );
  INV_X1 U12963 ( .A(n12565), .ZN(n12726) );
  XNOR2_X1 U12964 ( .A(n11106), .B(n12726), .ZN(n16195) );
  NAND2_X1 U12965 ( .A1(n16195), .A2(n15090), .ZN(n11107) );
  OAI211_X1 U12966 ( .C1(n16191), .C2(n15054), .A(n11108), .B(n11107), .ZN(
        P1_U3289) );
  NOR2_X1 U12967 ( .A1(n11121), .A2(n11109), .ZN(n11111) );
  NOR2_X1 U12968 ( .A1(n11111), .A2(n11110), .ZN(n11113) );
  INV_X1 U12969 ( .A(n16294), .ZN(n11126) );
  AOI22_X1 U12970 ( .A1(n11126), .A2(P3_REG1_REG_10__SCAN_IN), .B1(n8943), 
        .B2(n16294), .ZN(n11112) );
  AOI21_X1 U12971 ( .B1(n11113), .B2(n11112), .A(n11454), .ZN(n11133) );
  NAND2_X1 U12972 ( .A1(n11115), .A2(n11114), .ZN(n11118) );
  MUX2_X1 U12973 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n8634), .Z(n11116) );
  NOR2_X1 U12974 ( .A1(n11116), .A2(n16294), .ZN(n11460) );
  AOI21_X1 U12975 ( .B1(n11116), .B2(n16294), .A(n11460), .ZN(n11117) );
  AND2_X1 U12976 ( .A1(n11118), .A2(n11117), .ZN(n11459) );
  NOR2_X1 U12977 ( .A1(n11118), .A2(n11117), .ZN(n11119) );
  OAI21_X1 U12978 ( .B1(n11459), .B2(n11119), .A(n15970), .ZN(n11132) );
  AOI22_X1 U12979 ( .A1(n11126), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n8946), 
        .B2(n16294), .ZN(n11123) );
  AOI21_X1 U12980 ( .B1(n11124), .B2(n11123), .A(n11456), .ZN(n11129) );
  INV_X1 U12981 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n11125) );
  NOR2_X1 U12982 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11125), .ZN(n11899) );
  AOI21_X1 U12983 ( .B1(n15961), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11899), 
        .ZN(n11128) );
  NAND2_X1 U12984 ( .A1(n13713), .A2(n11126), .ZN(n11127) );
  OAI211_X1 U12985 ( .C1(n11129), .C2(n15999), .A(n11128), .B(n11127), .ZN(
        n11130) );
  INV_X1 U12986 ( .A(n11130), .ZN(n11131) );
  OAI211_X1 U12987 ( .C1(n11133), .C2(n15993), .A(n11132), .B(n11131), .ZN(
        P3_U3192) );
  NAND2_X1 U12988 ( .A1(n11545), .A2(n9720), .ZN(n11136) );
  AOI22_X1 U12989 ( .A1(n9659), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n13109), 
        .B2(n11134), .ZN(n11135) );
  INV_X1 U12990 ( .A(n16304), .ZN(n11262) );
  XNOR2_X1 U12991 ( .A(n16304), .B(n11516), .ZN(n11507) );
  NAND2_X1 U12992 ( .A1(n14257), .A2(n7431), .ZN(n11505) );
  XNOR2_X1 U12993 ( .A(n11507), .B(n11505), .ZN(n11142) );
  INV_X1 U12994 ( .A(n11137), .ZN(n11140) );
  OAI21_X1 U12995 ( .B1(n11140), .B2(n11139), .A(n11138), .ZN(n11141) );
  OAI21_X1 U12996 ( .B1(n11142), .B2(n11141), .A(n11506), .ZN(n11143) );
  NAND2_X1 U12997 ( .A1(n11143), .A2(n14232), .ZN(n11155) );
  NAND2_X1 U12998 ( .A1(n9742), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n11150) );
  NOR2_X1 U12999 ( .A1(n11144), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n11145) );
  OR2_X1 U13000 ( .A1(n11253), .A2(n11145), .ZN(n11502) );
  INV_X1 U13001 ( .A(n11502), .ZN(n11146) );
  NAND2_X1 U13002 ( .A1(n11931), .A2(n11146), .ZN(n11149) );
  NAND2_X1 U13003 ( .A1(n13386), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n11148) );
  NAND2_X1 U13004 ( .A1(n13368), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n11147) );
  NAND4_X1 U13005 ( .A1(n11150), .A2(n11149), .A3(n11148), .A4(n11147), .ZN(
        n14256) );
  INV_X1 U13006 ( .A(n14256), .ZN(n11335) );
  OAI22_X1 U13007 ( .A1(n13185), .A2(n14521), .B1(n11335), .B2(n14523), .ZN(
        n11281) );
  INV_X1 U13008 ( .A(n11281), .ZN(n11152) );
  OAI22_X1 U13009 ( .A1(n14244), .A2(n11152), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11151), .ZN(n11153) );
  AOI21_X1 U13010 ( .B1(n16302), .B2(n14242), .A(n11153), .ZN(n11154) );
  OAI211_X1 U13011 ( .C1(n11262), .C2(n12244), .A(n11155), .B(n11154), .ZN(
        P2_U3189) );
  AOI21_X1 U13012 ( .B1(n16170), .B2(n13183), .A(n11156), .ZN(n11157) );
  OAI211_X1 U13013 ( .C1(n9885), .C2(n11159), .A(n11158), .B(n11157), .ZN(
        n11161) );
  NAND2_X1 U13014 ( .A1(n11161), .A2(n16358), .ZN(n11160) );
  OAI21_X1 U13015 ( .B1(n16358), .B2(n10194), .A(n11160), .ZN(P2_U3508) );
  INV_X1 U13016 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11163) );
  NAND2_X1 U13017 ( .A1(n11161), .A2(n14668), .ZN(n11162) );
  OAI21_X1 U13018 ( .B1(n14668), .B2(n11163), .A(n11162), .ZN(P2_U3457) );
  AOI22_X1 U13019 ( .A1(n12520), .A2(n14855), .B1(n8541), .B2(n12575), .ZN(
        n11168) );
  NAND2_X1 U13020 ( .A1(n12575), .A2(n12494), .ZN(n11165) );
  NAND2_X1 U13021 ( .A1(n11165), .A2(n11164), .ZN(n11166) );
  XNOR2_X1 U13022 ( .A(n11166), .B(n12203), .ZN(n11167) );
  NAND2_X1 U13023 ( .A1(n11168), .A2(n11167), .ZN(n11227) );
  INV_X1 U13024 ( .A(n11167), .ZN(n11170) );
  INV_X1 U13025 ( .A(n11168), .ZN(n11169) );
  NAND2_X1 U13026 ( .A1(n11170), .A2(n11169), .ZN(n11229) );
  NAND2_X1 U13027 ( .A1(n11227), .A2(n11229), .ZN(n11176) );
  OR2_X1 U13028 ( .A1(n11173), .A2(n11172), .ZN(n11171) );
  NAND2_X1 U13029 ( .A1(n11173), .A2(n11172), .ZN(n11174) );
  XOR2_X1 U13030 ( .A(n11228), .B(n11176), .Z(n11183) );
  NAND2_X1 U13031 ( .A1(n14811), .A2(n11177), .ZN(n11179) );
  OAI211_X1 U13032 ( .C1(n11180), .C2(n14809), .A(n11179), .B(n11178), .ZN(
        n11181) );
  AOI21_X1 U13033 ( .B1(n12575), .B2(n14826), .A(n11181), .ZN(n11182) );
  OAI21_X1 U13034 ( .B1(n11183), .B2(n14829), .A(n11182), .ZN(P1_U3239) );
  INV_X1 U13035 ( .A(n12176), .ZN(n11203) );
  NOR2_X1 U13036 ( .A1(n11185), .A2(n11184), .ZN(n14902) );
  INV_X1 U13037 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11186) );
  MUX2_X1 U13038 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n11186), .S(n14901), .Z(
        n11187) );
  OAI21_X1 U13039 ( .B1(n14907), .B2(n14902), .A(n11187), .ZN(n14905) );
  OAI21_X1 U13040 ( .B1(n11186), .B2(n11188), .A(n14905), .ZN(n11189) );
  INV_X1 U13041 ( .A(n11189), .ZN(n11190) );
  XNOR2_X1 U13042 ( .A(n11189), .B(n12076), .ZN(n15848) );
  NOR2_X1 U13043 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n15848), .ZN(n15847) );
  AOI21_X1 U13044 ( .B1(n11190), .B2(n15853), .A(n15847), .ZN(n11194) );
  INV_X1 U13045 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11192) );
  NAND2_X1 U13046 ( .A1(n12176), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11441) );
  INV_X1 U13047 ( .A(n11441), .ZN(n11191) );
  AOI21_X1 U13048 ( .B1(n11192), .B2(n11203), .A(n11191), .ZN(n11193) );
  NAND2_X1 U13049 ( .A1(n11193), .A2(n11194), .ZN(n11440) );
  OAI211_X1 U13050 ( .C1(n11194), .C2(n11193), .A(n7422), .B(n11440), .ZN(
        n11202) );
  NAND2_X1 U13051 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14751)
         );
  AOI21_X1 U13052 ( .B1(n11781), .B2(P1_REG1_REG_13__SCAN_IN), .A(n11195), 
        .ZN(n14895) );
  XOR2_X1 U13053 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n14901), .Z(n14896) );
  NAND2_X1 U13054 ( .A1(n14895), .A2(n14896), .ZN(n14894) );
  OAI21_X1 U13055 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n14901), .A(n14894), 
        .ZN(n11196) );
  XOR2_X1 U13056 ( .A(n12076), .B(n11196), .Z(n15846) );
  NOR2_X1 U13057 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n15846), .ZN(n15845) );
  AOI21_X1 U13058 ( .B1(n15853), .B2(n11196), .A(n15845), .ZN(n11198) );
  XOR2_X1 U13059 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n12176), .Z(n11197) );
  NAND2_X1 U13060 ( .A1(n11197), .A2(n11198), .ZN(n11447) );
  OAI211_X1 U13061 ( .C1(n11198), .C2(n11197), .A(n16018), .B(n11447), .ZN(
        n11199) );
  NAND2_X1 U13062 ( .A1(n14751), .A2(n11199), .ZN(n11200) );
  AOI21_X1 U13063 ( .B1(n14866), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11200), 
        .ZN(n11201) );
  OAI211_X1 U13064 ( .C1(n16022), .C2(n11203), .A(n11202), .B(n11201), .ZN(
        P1_U3259) );
  XNOR2_X1 U13065 ( .A(n16199), .B(n10763), .ZN(n11301) );
  XNOR2_X1 U13066 ( .A(n11301), .B(n13619), .ZN(n11207) );
  OAI21_X1 U13067 ( .B1(n11207), .B2(n11206), .A(n11303), .ZN(n11208) );
  NAND2_X1 U13068 ( .A1(n11208), .A2(n13587), .ZN(n11213) );
  OAI22_X1 U13069 ( .A1(n13575), .A2(n11626), .B1(n11209), .B2(n13600), .ZN(
        n11210) );
  AOI211_X1 U13070 ( .C1(n13606), .C2(n16199), .A(n11211), .B(n11210), .ZN(
        n11212) );
  OAI211_X1 U13071 ( .C1(n11419), .C2(n13604), .A(n11213), .B(n11212), .ZN(
        P3_U3167) );
  NAND2_X1 U13072 ( .A1(n12863), .A2(n13036), .ZN(n11676) );
  NAND2_X1 U13073 ( .A1(n16178), .A2(n11676), .ZN(n11214) );
  XNOR2_X1 U13074 ( .A(n11215), .B(n13004), .ZN(n16177) );
  INV_X1 U13075 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11223) );
  NAND2_X1 U13076 ( .A1(n11217), .A2(n11216), .ZN(n11220) );
  INV_X1 U13077 ( .A(n11220), .ZN(n11219) );
  AOI21_X1 U13078 ( .B1(n11219), .B2(n11218), .A(n16107), .ZN(n11222) );
  NAND2_X1 U13079 ( .A1(n11220), .A2(n13004), .ZN(n11413) );
  OAI22_X1 U13080 ( .A1(n16102), .A2(n16103), .B1(n11306), .B2(n16101), .ZN(
        n11221) );
  AOI21_X1 U13081 ( .B1(n11222), .B2(n11413), .A(n11221), .ZN(n16179) );
  MUX2_X1 U13082 ( .A(n11223), .B(n16179), .S(n16121), .Z(n11226) );
  AOI22_X1 U13083 ( .A1(n13933), .A2(n16182), .B1(n13868), .B2(n11224), .ZN(
        n11225) );
  OAI211_X1 U13084 ( .C1(n13937), .C2(n16177), .A(n11226), .B(n11225), .ZN(
        P3_U3229) );
  NAND2_X1 U13085 ( .A1(n11228), .A2(n11227), .ZN(n11230) );
  NAND2_X1 U13086 ( .A1(n16240), .A2(n12494), .ZN(n11232) );
  NAND2_X1 U13087 ( .A1(n11232), .A2(n11231), .ZN(n11233) );
  XNOR2_X1 U13088 ( .A(n11233), .B(n12203), .ZN(n11484) );
  NAND2_X1 U13089 ( .A1(n16240), .A2(n8541), .ZN(n11236) );
  NAND2_X1 U13090 ( .A1(n12520), .A2(n14854), .ZN(n11235) );
  NAND2_X1 U13091 ( .A1(n11236), .A2(n11235), .ZN(n11485) );
  XNOR2_X1 U13092 ( .A(n11484), .B(n11485), .ZN(n11237) );
  OAI211_X1 U13093 ( .C1(n11238), .C2(n11237), .A(n11488), .B(n14796), .ZN(
        n11242) );
  NAND2_X1 U13094 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n14881) );
  OAI21_X1 U13095 ( .B1(n14809), .B2(n11239), .A(n14881), .ZN(n11240) );
  AOI21_X1 U13096 ( .B1(n16239), .B2(n14811), .A(n11240), .ZN(n11241) );
  OAI211_X1 U13097 ( .C1(n8342), .C2(n14804), .A(n11242), .B(n11241), .ZN(
        P1_U3213) );
  NAND2_X1 U13098 ( .A1(n11550), .A2(n9720), .ZN(n11245) );
  AOI22_X1 U13099 ( .A1(n9659), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n13109), 
        .B2(n11243), .ZN(n11244) );
  XNOR2_X1 U13100 ( .A(n13197), .B(n11335), .ZN(n13435) );
  NAND2_X1 U13101 ( .A1(n13183), .A2(n13185), .ZN(n11248) );
  INV_X1 U13102 ( .A(n14257), .ZN(n11249) );
  XNOR2_X1 U13103 ( .A(n16304), .B(n11249), .ZN(n13434) );
  OR2_X1 U13104 ( .A1(n16304), .A2(n11249), .ZN(n11250) );
  INV_X1 U13105 ( .A(n11337), .ZN(n11251) );
  AOI21_X1 U13106 ( .B1(n13435), .B2(n11252), .A(n11251), .ZN(n11261) );
  OR2_X1 U13107 ( .A1(n11253), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n11254) );
  AND2_X1 U13108 ( .A1(n11338), .A2(n11254), .ZN(n11523) );
  NAND2_X1 U13109 ( .A1(n11931), .A2(n11523), .ZN(n11258) );
  NAND2_X1 U13110 ( .A1(n9742), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n11257) );
  NAND2_X1 U13111 ( .A1(n13386), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n11256) );
  NAND2_X1 U13112 ( .A1(n13368), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n11255) );
  NAND4_X1 U13113 ( .A1(n11258), .A2(n11257), .A3(n11256), .A4(n11255), .ZN(
        n14255) );
  NAND2_X1 U13114 ( .A1(n14255), .A2(n14439), .ZN(n11260) );
  NAND2_X1 U13115 ( .A1(n14257), .A2(n14438), .ZN(n11259) );
  AND2_X1 U13116 ( .A1(n11260), .A2(n11259), .ZN(n11499) );
  OAI21_X1 U13117 ( .B1(n11261), .B2(n14486), .A(n11499), .ZN(n16356) );
  INV_X1 U13118 ( .A(n16356), .ZN(n11273) );
  OAI22_X1 U13119 ( .A1(n14549), .A2(n10835), .B1(n11502), .B2(n14510), .ZN(
        n11265) );
  INV_X1 U13120 ( .A(n11263), .ZN(n11283) );
  INV_X1 U13121 ( .A(n13197), .ZN(n16354) );
  OAI211_X1 U13122 ( .C1(n11283), .C2(n16354), .A(n14507), .B(n11347), .ZN(
        n16351) );
  NOR2_X1 U13123 ( .A1(n16351), .A2(n14539), .ZN(n11264) );
  AOI211_X1 U13124 ( .C1(n16303), .C2(n13197), .A(n11265), .B(n11264), .ZN(
        n11272) );
  INV_X1 U13125 ( .A(n13434), .ZN(n11267) );
  OR2_X1 U13126 ( .A1(n16304), .A2(n14257), .ZN(n11268) );
  INV_X1 U13127 ( .A(n13435), .ZN(n11269) );
  NAND2_X1 U13128 ( .A1(n11270), .A2(n11269), .ZN(n16349) );
  NAND3_X1 U13129 ( .A1(n16350), .A2(n16349), .A3(n14515), .ZN(n11271) );
  OAI211_X1 U13130 ( .C1(n11273), .C2(n16405), .A(n11272), .B(n11271), .ZN(
        P2_U3254) );
  INV_X1 U13131 ( .A(n11274), .ZN(n11276) );
  OAI21_X1 U13132 ( .B1(n11276), .B2(n13434), .A(n11275), .ZN(n16307) );
  INV_X1 U13133 ( .A(n16307), .ZN(n11286) );
  INV_X1 U13134 ( .A(n11277), .ZN(n11278) );
  AOI211_X1 U13135 ( .C1(n13434), .C2(n11279), .A(n14486), .B(n11278), .ZN(
        n11280) );
  AOI211_X1 U13136 ( .C1(n14520), .C2(n16307), .A(n11281), .B(n11280), .ZN(
        n16310) );
  INV_X1 U13137 ( .A(n11282), .ZN(n11284) );
  AOI211_X1 U13138 ( .C1(n16304), .C2(n11284), .A(n7431), .B(n11283), .ZN(
        n16305) );
  AOI21_X1 U13139 ( .B1(n16170), .B2(n16304), .A(n16305), .ZN(n11285) );
  OAI211_X1 U13140 ( .C1(n11286), .C2(n9885), .A(n16310), .B(n11285), .ZN(
        n11288) );
  NAND2_X1 U13141 ( .A1(n11288), .A2(n16358), .ZN(n11287) );
  OAI21_X1 U13142 ( .B1(n16358), .B2(n10646), .A(n11287), .ZN(P2_U3509) );
  INV_X1 U13143 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11290) );
  NAND2_X1 U13144 ( .A1(n11288), .A2(n14668), .ZN(n11289) );
  OAI21_X1 U13145 ( .B1(n14668), .B2(n11290), .A(n11289), .ZN(P2_U3460) );
  INV_X1 U13146 ( .A(SI_24_), .ZN(n11293) );
  INV_X1 U13147 ( .A(n11291), .ZN(n11292) );
  OAI222_X1 U13148 ( .A1(P3_U3151), .A2(n11294), .B1(n13462), .B2(n11293), 
        .C1(n14119), .C2(n11292), .ZN(P3_U3271) );
  XOR2_X1 U13149 ( .A(n13001), .B(n11295), .Z(n11296) );
  AOI222_X1 U13150 ( .A1(n16054), .A2(n11296), .B1(n13620), .B2(n13943), .C1(
        n13622), .C2(n13941), .ZN(n11326) );
  XNOR2_X1 U13151 ( .A(n13001), .B(n11297), .ZN(n16133) );
  AOI22_X1 U13152 ( .A1(n16133), .A2(n16229), .B1(n16200), .B2(n11329), .ZN(
        n11298) );
  NAND2_X1 U13153 ( .A1(n11326), .A2(n11298), .ZN(n16134) );
  INV_X1 U13154 ( .A(n16134), .ZN(n11300) );
  INV_X1 U13155 ( .A(n14106), .ZN(n11685) );
  AOI22_X1 U13156 ( .A1(n16133), .A2(n11685), .B1(P3_REG0_REG_3__SCAN_IN), 
        .B2(n16415), .ZN(n11299) );
  OAI21_X1 U13157 ( .B1(n11300), .B2(n16415), .A(n11299), .ZN(P3_U3399) );
  NAND2_X1 U13158 ( .A1(n11301), .A2(n11306), .ZN(n11302) );
  XNOR2_X1 U13159 ( .A(n16215), .B(n8025), .ZN(n11611) );
  XNOR2_X1 U13160 ( .A(n11611), .B(n11626), .ZN(n11304) );
  OAI211_X1 U13161 ( .C1(n11305), .C2(n11304), .A(n11613), .B(n13587), .ZN(
        n11311) );
  OAI22_X1 U13162 ( .A1(n13575), .A2(n11670), .B1(n11306), .B2(n13600), .ZN(
        n11307) );
  AOI211_X1 U13163 ( .C1(n13606), .C2(n11309), .A(n11308), .B(n11307), .ZN(
        n11310) );
  OAI211_X1 U13164 ( .C1(n11534), .C2(n13604), .A(n11311), .B(n11310), .ZN(
        P3_U3179) );
  XNOR2_X1 U13165 ( .A(n11312), .B(n13005), .ZN(n16232) );
  OAI211_X1 U13166 ( .C1(n11314), .C2(n13005), .A(n11313), .B(n16054), .ZN(
        n11316) );
  AOI22_X1 U13167 ( .A1(n13616), .A2(n13943), .B1(n13941), .B2(n13618), .ZN(
        n11315) );
  NAND2_X1 U13168 ( .A1(n11316), .A2(n11315), .ZN(n16235) );
  NAND2_X1 U13169 ( .A1(n16235), .A2(n16121), .ZN(n11319) );
  OAI22_X1 U13170 ( .A1(n13963), .A2(n16231), .B1(n11631), .B2(n16113), .ZN(
        n11317) );
  AOI21_X1 U13171 ( .B1(P3_REG2_REG_7__SCAN_IN), .B2(n16123), .A(n11317), .ZN(
        n11318) );
  OAI211_X1 U13172 ( .C1(n13937), .C2(n16232), .A(n11319), .B(n11318), .ZN(
        P3_U3226) );
  INV_X1 U13173 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n11323) );
  MUX2_X1 U13174 ( .A(n11323), .B(n13263), .S(n8006), .Z(n11324) );
  NAND2_X1 U13175 ( .A1(n12314), .A2(n11324), .ZN(n11325) );
  NAND2_X1 U13176 ( .A1(n11527), .A2(n11325), .ZN(n13262) );
  OAI222_X1 U13177 ( .A1(n14693), .A2(n13263), .B1(P2_U3088), .B2(n13093), 
        .C1(n14691), .C2(n13262), .ZN(P2_U3305) );
  INV_X1 U13178 ( .A(n16133), .ZN(n11332) );
  MUX2_X1 U13179 ( .A(n11327), .B(n11326), .S(n16121), .Z(n11331) );
  AOI22_X1 U13180 ( .A1(n13933), .A2(n11329), .B1(n13868), .B2(n11328), .ZN(
        n11330) );
  OAI211_X1 U13181 ( .C1(n13937), .C2(n11332), .A(n11331), .B(n11330), .ZN(
        P3_U3230) );
  NAND2_X1 U13182 ( .A1(n11562), .A2(n9720), .ZN(n11334) );
  AOI22_X1 U13183 ( .A1(n9659), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n11431), 
        .B2(n13109), .ZN(n11333) );
  XNOR2_X1 U13184 ( .A(n13202), .B(n14255), .ZN(n13436) );
  NAND2_X1 U13185 ( .A1(n13197), .A2(n11335), .ZN(n11336) );
  XOR2_X1 U13186 ( .A(n11762), .B(n13436), .Z(n11344) );
  NAND2_X1 U13187 ( .A1(n11338), .A2(n11705), .ZN(n11339) );
  AND2_X1 U13188 ( .A1(n11698), .A2(n11339), .ZN(n16395) );
  NAND2_X1 U13189 ( .A1(n16395), .A2(n11931), .ZN(n11343) );
  NAND2_X1 U13190 ( .A1(n9742), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11342) );
  NAND2_X1 U13191 ( .A1(n13386), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n11341) );
  NAND2_X1 U13192 ( .A1(n13368), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11340) );
  NAND4_X1 U13193 ( .A1(n11343), .A2(n11342), .A3(n11341), .A4(n11340), .ZN(
        n14254) );
  AOI22_X1 U13194 ( .A1(n14439), .A2(n14254), .B1(n14256), .B2(n14438), .ZN(
        n11521) );
  OAI21_X1 U13195 ( .B1(n11344), .B2(n14486), .A(n11521), .ZN(n11661) );
  INV_X1 U13196 ( .A(n11661), .ZN(n11352) );
  NAND2_X1 U13197 ( .A1(n13197), .A2(n14256), .ZN(n11345) );
  XNOR2_X1 U13198 ( .A(n11772), .B(n13436), .ZN(n11663) );
  INV_X1 U13199 ( .A(n13202), .ZN(n11526) );
  INV_X1 U13200 ( .A(n11907), .ZN(n11346) );
  AOI211_X1 U13201 ( .C1(n13202), .C2(n11347), .A(n14445), .B(n11346), .ZN(
        n11662) );
  NAND2_X1 U13202 ( .A1(n11662), .A2(n16306), .ZN(n11349) );
  AOI22_X1 U13203 ( .A1(n16405), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n11523), 
        .B2(n16394), .ZN(n11348) );
  OAI211_X1 U13204 ( .C1(n11526), .C2(n16398), .A(n11349), .B(n11348), .ZN(
        n11350) );
  AOI21_X1 U13205 ( .B1(n11663), .B2(n14515), .A(n11350), .ZN(n11351) );
  OAI21_X1 U13206 ( .B1(n11352), .B2(n16405), .A(n11351), .ZN(P2_U3253) );
  INV_X1 U13207 ( .A(n14854), .ZN(n11353) );
  AND2_X1 U13208 ( .A1(n16240), .A2(n11353), .ZN(n11354) );
  NAND2_X1 U13209 ( .A1(n11356), .A2(n12491), .ZN(n11359) );
  AOI22_X1 U13210 ( .A1(n12399), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n12398), 
        .B2(n11357), .ZN(n11358) );
  NAND2_X1 U13211 ( .A1(n11359), .A2(n11358), .ZN(n12583) );
  XNOR2_X1 U13212 ( .A(n12583), .B(n14853), .ZN(n12731) );
  INV_X1 U13213 ( .A(n14853), .ZN(n11482) );
  OR2_X1 U13214 ( .A1(n12583), .A2(n11482), .ZN(n11360) );
  NAND2_X1 U13215 ( .A1(n11361), .A2(n11360), .ZN(n11574) );
  AOI22_X1 U13216 ( .A1(n12399), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n11363), 
        .B2(n12398), .ZN(n11364) );
  NAND2_X1 U13217 ( .A1(n10089), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n11371) );
  NAND2_X1 U13218 ( .A1(n7427), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n11370) );
  AND2_X1 U13219 ( .A1(n11366), .A2(n11365), .ZN(n11367) );
  NOR2_X1 U13220 ( .A1(n11376), .A2(n11367), .ZN(n11873) );
  NAND2_X1 U13221 ( .A1(n12526), .A2(n11873), .ZN(n11369) );
  NAND2_X1 U13222 ( .A1(n12686), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n11368) );
  NAND4_X1 U13223 ( .A1(n11371), .A2(n11370), .A3(n11369), .A4(n11368), .ZN(
        n14852) );
  INV_X1 U13224 ( .A(n14852), .ZN(n11575) );
  XNOR2_X1 U13225 ( .A(n11574), .B(n8658), .ZN(n11385) );
  OR2_X1 U13226 ( .A1(n16240), .A2(n14854), .ZN(n11372) );
  OR2_X1 U13227 ( .A1(n12583), .A2(n14853), .ZN(n11374) );
  OAI21_X1 U13228 ( .B1(n11375), .B2(n12733), .A(n11544), .ZN(n16285) );
  NAND2_X1 U13229 ( .A1(n16285), .A2(n16372), .ZN(n11384) );
  NAND2_X1 U13230 ( .A1(n7427), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n11381) );
  NAND2_X1 U13231 ( .A1(n10089), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n11380) );
  NOR2_X1 U13232 ( .A1(n11376), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11377) );
  OR2_X1 U13233 ( .A1(n11554), .A2(n11377), .ZN(n11744) );
  INV_X1 U13234 ( .A(n11744), .ZN(n11651) );
  NAND2_X1 U13235 ( .A1(n12526), .A2(n11651), .ZN(n11379) );
  NAND2_X1 U13236 ( .A1(n12686), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n11378) );
  NAND4_X1 U13237 ( .A1(n11381), .A2(n11380), .A3(n11379), .A4(n11378), .ZN(
        n14851) );
  NAND2_X1 U13238 ( .A1(n14851), .A2(n14799), .ZN(n11383) );
  NAND2_X1 U13239 ( .A1(n14853), .A2(n14806), .ZN(n11382) );
  AND2_X1 U13240 ( .A1(n11383), .A2(n11382), .ZN(n11876) );
  OAI211_X1 U13241 ( .C1(n16379), .C2(n11385), .A(n11384), .B(n11876), .ZN(
        n16283) );
  INV_X1 U13242 ( .A(n16283), .ZN(n11391) );
  INV_X1 U13243 ( .A(n12592), .ZN(n16282) );
  INV_X1 U13244 ( .A(n12583), .ZN(n11399) );
  INV_X1 U13245 ( .A(n11397), .ZN(n11386) );
  OAI211_X1 U13246 ( .C1(n16282), .C2(n11386), .A(n16322), .B(n11603), .ZN(
        n16281) );
  AOI22_X1 U13247 ( .A1(n16347), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n11873), 
        .B2(n16336), .ZN(n11388) );
  NAND2_X1 U13248 ( .A1(n16337), .A2(n12592), .ZN(n11387) );
  OAI211_X1 U13249 ( .C1(n16281), .C2(n15051), .A(n11388), .B(n11387), .ZN(
        n11389) );
  AOI21_X1 U13250 ( .B1(n16285), .B2(n16342), .A(n11389), .ZN(n11390) );
  OAI21_X1 U13251 ( .B1(n11391), .B2(n16347), .A(n11390), .ZN(P1_U3284) );
  OAI222_X1 U13252 ( .A1(P3_U3151), .A2(n11393), .B1(n14119), .B2(n11392), 
        .C1(n15461), .C2(n13462), .ZN(P3_U3270) );
  INV_X1 U13253 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n11409) );
  OR2_X1 U13254 ( .A1(n11394), .A2(n7429), .ZN(n11395) );
  NAND2_X1 U13255 ( .A1(n11396), .A2(n11395), .ZN(n11477) );
  OAI211_X1 U13256 ( .C1(n11398), .C2(n11399), .A(n16322), .B(n11397), .ZN(
        n11473) );
  OAI21_X1 U13257 ( .B1(n11399), .B2(n16378), .A(n11473), .ZN(n11407) );
  XNOR2_X1 U13258 ( .A(n11400), .B(n7429), .ZN(n11404) );
  NAND2_X1 U13259 ( .A1(n14852), .A2(n14807), .ZN(n11402) );
  NAND2_X1 U13260 ( .A1(n14854), .A2(n14806), .ZN(n11401) );
  AND2_X1 U13261 ( .A1(n11402), .A2(n11401), .ZN(n11495) );
  INV_X1 U13262 ( .A(n11495), .ZN(n11403) );
  AOI21_X1 U13263 ( .B1(n11404), .B2(n16194), .A(n11403), .ZN(n11406) );
  NAND2_X1 U13264 ( .A1(n11477), .A2(n16372), .ZN(n11405) );
  NAND2_X1 U13265 ( .A1(n11406), .A2(n11405), .ZN(n11474) );
  AOI211_X1 U13266 ( .C1(n16332), .C2(n11477), .A(n11407), .B(n11474), .ZN(
        n11410) );
  OR2_X1 U13267 ( .A1(n11410), .A2(n16388), .ZN(n11408) );
  OAI21_X1 U13268 ( .B1(n16391), .B2(n11409), .A(n11408), .ZN(P1_U3483) );
  OR2_X1 U13269 ( .A1(n11410), .A2(n16385), .ZN(n11411) );
  OAI21_X1 U13270 ( .B1(n16387), .B2(n9976), .A(n11411), .ZN(P1_U3536) );
  AND2_X1 U13271 ( .A1(n11413), .A2(n11412), .ZN(n11416) );
  AND2_X1 U13272 ( .A1(n11415), .A2(n11414), .ZN(n11536) );
  OAI21_X1 U13273 ( .B1(n11416), .B2(n9223), .A(n11536), .ZN(n11417) );
  AOI222_X1 U13274 ( .A1(n16054), .A2(n11417), .B1(n13620), .B2(n13941), .C1(
        n13618), .C2(n13943), .ZN(n16203) );
  XNOR2_X1 U13275 ( .A(n11418), .B(n12997), .ZN(n16201) );
  NOR2_X1 U13276 ( .A1(n16121), .A2(n8864), .ZN(n11422) );
  OAI22_X1 U13277 ( .A1(n11420), .A2(n13963), .B1(n11419), .B2(n16113), .ZN(
        n11421) );
  AOI211_X1 U13278 ( .C1(n16201), .C2(n13967), .A(n11422), .B(n11421), .ZN(
        n11423) );
  OAI21_X1 U13279 ( .B1(n16203), .B2(n16123), .A(n11423), .ZN(P3_U3228) );
  INV_X1 U13280 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11424) );
  MUX2_X1 U13281 ( .A(n11424), .B(P2_REG1_REG_13__SCAN_IN), .S(n11691), .Z(
        n11427) );
  NOR2_X1 U13282 ( .A1(n11426), .A2(n11427), .ZN(n11640) );
  AOI211_X1 U13283 ( .C1(n11427), .C2(n11426), .A(n15813), .B(n11640), .ZN(
        n11439) );
  INV_X1 U13284 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11428) );
  MUX2_X1 U13285 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n11428), .S(n11691), .Z(
        n11429) );
  INV_X1 U13286 ( .A(n11429), .ZN(n11433) );
  OAI21_X1 U13287 ( .B1(n11431), .B2(P2_REG2_REG_12__SCAN_IN), .A(n11430), 
        .ZN(n11432) );
  NOR2_X1 U13288 ( .A1(n11432), .A2(n11433), .ZN(n11632) );
  AOI211_X1 U13289 ( .C1(n11433), .C2(n11432), .A(n15817), .B(n11632), .ZN(
        n11438) );
  NAND2_X1 U13290 ( .A1(n15838), .A2(n11691), .ZN(n11436) );
  NAND2_X1 U13291 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n11435)
         );
  NAND2_X1 U13292 ( .A1(n15800), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n11434) );
  NAND3_X1 U13293 ( .A1(n11436), .A2(n11435), .A3(n11434), .ZN(n11437) );
  OR3_X1 U13294 ( .A1(n11439), .A2(n11438), .A3(n11437), .ZN(P2_U3227) );
  NAND2_X1 U13295 ( .A1(n11441), .A2(n11440), .ZN(n11446) );
  NAND2_X1 U13296 ( .A1(n11751), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11442) );
  OAI21_X1 U13297 ( .B1(n11751), .B2(P1_REG2_REG_17__SCAN_IN), .A(n11442), 
        .ZN(n11445) );
  INV_X1 U13298 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n11444) );
  NAND2_X1 U13299 ( .A1(n11751), .A2(n11444), .ZN(n11443) );
  OAI211_X1 U13300 ( .C1(n11444), .C2(n11751), .A(n11446), .B(n11443), .ZN(
        n11748) );
  OAI211_X1 U13301 ( .C1(n11446), .C2(n11445), .A(n11748), .B(n7422), .ZN(
        n11453) );
  NAND2_X1 U13302 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14763)
         );
  INV_X1 U13303 ( .A(n11447), .ZN(n11448) );
  AOI21_X1 U13304 ( .B1(n12176), .B2(P1_REG1_REG_16__SCAN_IN), .A(n11448), 
        .ZN(n11752) );
  INV_X1 U13305 ( .A(n11751), .ZN(n12249) );
  XNOR2_X1 U13306 ( .A(n12249), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n11753) );
  XOR2_X1 U13307 ( .A(n11752), .B(n11753), .Z(n11449) );
  NAND2_X1 U13308 ( .A1(n16018), .A2(n11449), .ZN(n11450) );
  NAND2_X1 U13309 ( .A1(n14763), .A2(n11450), .ZN(n11451) );
  AOI21_X1 U13310 ( .B1(n14866), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n11451), 
        .ZN(n11452) );
  OAI211_X1 U13311 ( .C1(n16022), .C2(n11751), .A(n11453), .B(n11452), .ZN(
        P1_U3260) );
  INV_X1 U13312 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n16317) );
  AOI21_X1 U13313 ( .B1(n16317), .B2(n11455), .A(n13656), .ZN(n11471) );
  INV_X1 U13314 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11995) );
  AOI21_X1 U13315 ( .B1(n11995), .B2(n11457), .A(n13625), .ZN(n11458) );
  NOR2_X1 U13316 ( .A1(n11458), .A2(n15999), .ZN(n11469) );
  XNOR2_X1 U13317 ( .A(n13635), .B(n13655), .ZN(n11461) );
  NAND2_X1 U13318 ( .A1(n11461), .A2(n11462), .ZN(n11463) );
  AOI21_X1 U13319 ( .B1(n11463), .B2(n13636), .A(n15991), .ZN(n11468) );
  INV_X1 U13320 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11464) );
  NOR2_X1 U13321 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11464), .ZN(n12100) );
  AOI21_X1 U13322 ( .B1(n15961), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n12100), 
        .ZN(n11465) );
  OAI21_X1 U13323 ( .B1(n15984), .B2(n11466), .A(n11465), .ZN(n11467) );
  NOR3_X1 U13324 ( .A1(n11469), .A2(n11468), .A3(n11467), .ZN(n11470) );
  OAI21_X1 U13325 ( .B1(n11471), .B2(n15993), .A(n11470), .ZN(P3_U3193) );
  AOI22_X1 U13326 ( .A1(n16337), .A2(n12583), .B1(n11492), .B2(n16336), .ZN(
        n11472) );
  OAI21_X1 U13327 ( .B1(n15051), .B2(n11473), .A(n11472), .ZN(n11476) );
  MUX2_X1 U13328 ( .A(n11474), .B(P1_REG2_REG_8__SCAN_IN), .S(n16347), .Z(
        n11475) );
  AOI211_X1 U13329 ( .C1(n16342), .C2(n11477), .A(n11476), .B(n11475), .ZN(
        n11478) );
  INV_X1 U13330 ( .A(n11478), .ZN(P1_U3285) );
  NAND2_X1 U13331 ( .A1(n12583), .A2(n12494), .ZN(n11480) );
  NAND2_X1 U13332 ( .A1(n11480), .A2(n11479), .ZN(n11481) );
  XNOR2_X1 U13333 ( .A(n11481), .B(n12203), .ZN(n11723) );
  NOR2_X1 U13334 ( .A1(n12483), .A2(n11482), .ZN(n11483) );
  AOI21_X1 U13335 ( .B1(n12583), .B2(n8541), .A(n11483), .ZN(n11722) );
  XNOR2_X1 U13336 ( .A(n11723), .B(n11722), .ZN(n11491) );
  INV_X1 U13337 ( .A(n11484), .ZN(n11486) );
  NAND2_X1 U13338 ( .A1(n11486), .A2(n11485), .ZN(n11487) );
  INV_X1 U13339 ( .A(n11725), .ZN(n11489) );
  AOI21_X1 U13340 ( .B1(n11491), .B2(n11490), .A(n11489), .ZN(n11498) );
  NAND2_X1 U13341 ( .A1(n14811), .A2(n11492), .ZN(n11494) );
  OAI211_X1 U13342 ( .C1(n11495), .C2(n14809), .A(n11494), .B(n11493), .ZN(
        n11496) );
  AOI21_X1 U13343 ( .B1(n12583), .B2(n14826), .A(n11496), .ZN(n11497) );
  OAI21_X1 U13344 ( .B1(n11498), .B2(n14829), .A(n11497), .ZN(P1_U3221) );
  INV_X1 U13345 ( .A(n11499), .ZN(n11500) );
  AOI22_X1 U13346 ( .A1(n14195), .A2(n11500), .B1(P2_REG3_REG_11__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11501) );
  OAI21_X1 U13347 ( .B1(n11502), .B2(n14218), .A(n11501), .ZN(n11512) );
  XNOR2_X1 U13348 ( .A(n13197), .B(n11516), .ZN(n11504) );
  AND2_X1 U13349 ( .A1(n14256), .A2(n14445), .ZN(n11503) );
  NAND2_X1 U13350 ( .A1(n11504), .A2(n11503), .ZN(n11514) );
  OAI21_X1 U13351 ( .B1(n11504), .B2(n11503), .A(n11514), .ZN(n11510) );
  INV_X1 U13352 ( .A(n11505), .ZN(n11508) );
  AOI211_X1 U13353 ( .C1(n11510), .C2(n11509), .A(n14248), .B(n11515), .ZN(
        n11511) );
  AOI211_X1 U13354 ( .C1(n13197), .C2(n14246), .A(n11512), .B(n11511), .ZN(
        n11513) );
  INV_X1 U13355 ( .A(n11513), .ZN(P2_U3208) );
  XNOR2_X1 U13356 ( .A(n13202), .B(n11516), .ZN(n11689) );
  NAND2_X1 U13357 ( .A1(n14255), .A2(n14445), .ZN(n11687) );
  XNOR2_X1 U13358 ( .A(n11689), .B(n11687), .ZN(n11517) );
  OAI21_X1 U13359 ( .B1(n11518), .B2(n11517), .A(n11688), .ZN(n11519) );
  NAND2_X1 U13360 ( .A1(n11519), .A2(n14232), .ZN(n11525) );
  OAI21_X1 U13361 ( .B1(n14244), .B2(n11521), .A(n11520), .ZN(n11522) );
  AOI21_X1 U13362 ( .B1(n11523), .B2(n14242), .A(n11522), .ZN(n11524) );
  OAI211_X1 U13363 ( .C1(n11526), .C2(n12244), .A(n11525), .B(n11524), .ZN(
        P2_U3196) );
  MUX2_X1 U13364 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n8006), .Z(n11528) );
  NAND2_X1 U13365 ( .A1(n11528), .A2(SI_23_), .ZN(n11713) );
  OAI21_X1 U13366 ( .B1(SI_23_), .B2(n11528), .A(n11713), .ZN(n11710) );
  XNOR2_X1 U13367 ( .A(n11712), .B(n11710), .ZN(n13278) );
  NAND2_X1 U13368 ( .A1(n13278), .A2(n11529), .ZN(n11531) );
  OR2_X1 U13369 ( .A1(n11530), .A2(P2_U3088), .ZN(n13460) );
  OAI211_X1 U13370 ( .C1(n13279), .C2(n14693), .A(n11531), .B(n13460), .ZN(
        P2_U3304) );
  INV_X1 U13371 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n12424) );
  NAND2_X1 U13372 ( .A1(n13278), .A2(n15248), .ZN(n11532) );
  OAI211_X1 U13373 ( .C1(n12424), .C2(n15262), .A(n11532), .B(n12774), .ZN(
        P1_U3332) );
  XNOR2_X1 U13374 ( .A(n11533), .B(n13006), .ZN(n16219) );
  OAI22_X1 U13375 ( .A1(n13963), .A2(n16215), .B1(n11534), .B2(n16113), .ZN(
        n11542) );
  AND2_X1 U13376 ( .A1(n11536), .A2(n11535), .ZN(n11538) );
  OAI211_X1 U13377 ( .C1(n11538), .C2(n12888), .A(n11537), .B(n16054), .ZN(
        n11540) );
  AOI22_X1 U13378 ( .A1(n13619), .A2(n13941), .B1(n13943), .B2(n13617), .ZN(
        n11539) );
  NAND2_X1 U13379 ( .A1(n11540), .A2(n11539), .ZN(n16217) );
  MUX2_X1 U13380 ( .A(n16217), .B(P3_REG2_REG_6__SCAN_IN), .S(n16123), .Z(
        n11541) );
  AOI211_X1 U13381 ( .C1(n13967), .C2(n16219), .A(n11542), .B(n11541), .ZN(
        n11543) );
  INV_X1 U13382 ( .A(n11543), .ZN(P3_U3227) );
  INV_X2 U13383 ( .A(n8724), .ZN(n12491) );
  NAND2_X1 U13384 ( .A1(n11545), .A2(n12491), .ZN(n11548) );
  AOI22_X1 U13385 ( .A1(n11546), .A2(n12398), .B1(n12399), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n11547) );
  XNOR2_X1 U13386 ( .A(n12601), .B(n14851), .ZN(n12734) );
  OR2_X1 U13387 ( .A1(n12601), .A2(n14851), .ZN(n11549) );
  NAND2_X1 U13388 ( .A1(n11550), .A2(n12491), .ZN(n11553) );
  AOI22_X1 U13389 ( .A1(n12399), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n12398), 
        .B2(n11551), .ZN(n11552) );
  NAND2_X1 U13390 ( .A1(n12524), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n11559) );
  NAND2_X1 U13391 ( .A1(n7427), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11558) );
  OR2_X1 U13392 ( .A1(n11554), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n11555) );
  AND2_X1 U13393 ( .A1(n11567), .A2(n11555), .ZN(n16335) );
  NAND2_X1 U13394 ( .A1(n12526), .A2(n16335), .ZN(n11557) );
  NAND2_X1 U13395 ( .A1(n12686), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n11556) );
  OAI21_X1 U13396 ( .B1(n16320), .B2(n16324), .A(n12606), .ZN(n11561) );
  NAND2_X1 U13397 ( .A1(n16320), .A2(n16324), .ZN(n11560) );
  NAND2_X1 U13398 ( .A1(n11561), .A2(n11560), .ZN(n11786) );
  NAND2_X1 U13399 ( .A1(n11562), .A2(n12491), .ZN(n11565) );
  AOI22_X1 U13400 ( .A1(n12398), .A2(n11563), .B1(n12399), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n11564) );
  NAND2_X1 U13401 ( .A1(n12524), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11572) );
  NAND2_X1 U13402 ( .A1(n12686), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n11571) );
  INV_X1 U13403 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n11566) );
  NAND2_X1 U13404 ( .A1(n11567), .A2(n11566), .ZN(n11568) );
  AND2_X1 U13405 ( .A1(n11583), .A2(n11568), .ZN(n12130) );
  NAND2_X1 U13406 ( .A1(n12526), .A2(n12130), .ZN(n11570) );
  NAND2_X1 U13407 ( .A1(n7426), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11569) );
  NAND4_X1 U13408 ( .A1(n11572), .A2(n11571), .A3(n11570), .A4(n11569), .ZN(
        n14849) );
  XNOR2_X1 U13409 ( .A(n11786), .B(n12736), .ZN(n16368) );
  NAND2_X1 U13410 ( .A1(n16086), .A2(n16372), .ZN(n11573) );
  AND2_X1 U13411 ( .A1(n16045), .A2(n11573), .ZN(n15088) );
  NAND2_X1 U13412 ( .A1(n11574), .A2(n8658), .ZN(n11577) );
  OR2_X1 U13413 ( .A1(n12592), .A2(n11575), .ZN(n11576) );
  NAND2_X1 U13414 ( .A1(n11577), .A2(n11576), .ZN(n11601) );
  NAND2_X1 U13415 ( .A1(n11601), .A2(n12734), .ZN(n11579) );
  INV_X1 U13416 ( .A(n14851), .ZN(n11739) );
  OR2_X1 U13417 ( .A1(n12601), .A2(n11739), .ZN(n11578) );
  AND2_X1 U13418 ( .A1(n16324), .A2(n14850), .ZN(n11580) );
  OR2_X1 U13419 ( .A1(n16324), .A2(n14850), .ZN(n11581) );
  INV_X1 U13420 ( .A(n12736), .ZN(n11785) );
  OAI211_X1 U13421 ( .C1(n7591), .C2(n12736), .A(n16194), .B(n11779), .ZN(
        n11590) );
  NAND2_X1 U13422 ( .A1(n10089), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11588) );
  NAND2_X1 U13423 ( .A1(n12686), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n11587) );
  INV_X1 U13424 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n11582) );
  NAND2_X1 U13425 ( .A1(n11583), .A2(n11582), .ZN(n11584) );
  AND2_X1 U13426 ( .A1(n11790), .A2(n11584), .ZN(n12212) );
  NAND2_X1 U13427 ( .A1(n12526), .A2(n12212), .ZN(n11586) );
  NAND2_X1 U13428 ( .A1(n7426), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11585) );
  NAND4_X1 U13429 ( .A1(n11588), .A2(n11587), .A3(n11586), .A4(n11585), .ZN(
        n14848) );
  AND2_X1 U13430 ( .A1(n14848), .A2(n14807), .ZN(n11589) );
  AOI21_X1 U13431 ( .B1(n14850), .B2(n14806), .A(n11589), .ZN(n12128) );
  NAND2_X1 U13432 ( .A1(n11590), .A2(n12128), .ZN(n16363) );
  INV_X1 U13433 ( .A(n16365), .ZN(n12133) );
  NAND2_X1 U13434 ( .A1(n16324), .A2(n16323), .ZN(n16321) );
  AOI211_X1 U13435 ( .C1(n16365), .C2(n16321), .A(n16142), .B(n7672), .ZN(
        n16364) );
  NAND2_X1 U13436 ( .A1(n16364), .A2(n16341), .ZN(n11592) );
  AOI22_X1 U13437 ( .A1(n16347), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n12130), 
        .B2(n16336), .ZN(n11591) );
  OAI211_X1 U13438 ( .C1(n12133), .C2(n16163), .A(n11592), .B(n11591), .ZN(
        n11593) );
  AOI21_X1 U13439 ( .B1(n16363), .B2(n16159), .A(n11593), .ZN(n11594) );
  OAI21_X1 U13440 ( .B1(n16368), .B2(n15088), .A(n11594), .ZN(P1_U3281) );
  INV_X1 U13441 ( .A(SI_26_), .ZN(n11596) );
  OAI222_X1 U13442 ( .A1(P3_U3151), .A2(n11597), .B1(n13462), .B2(n11596), 
        .C1(n14119), .C2(n11595), .ZN(P3_U3269) );
  INV_X1 U13443 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n11607) );
  OAI21_X1 U13444 ( .B1(n11599), .B2(n11600), .A(n11598), .ZN(n11659) );
  INV_X1 U13445 ( .A(n11659), .ZN(n11605) );
  XNOR2_X1 U13446 ( .A(n11601), .B(n11600), .ZN(n11602) );
  AOI22_X1 U13447 ( .A1(n11659), .A2(n16372), .B1(n11602), .B2(n16194), .ZN(
        n11656) );
  NAND2_X1 U13448 ( .A1(n14850), .A2(n14807), .ZN(n11648) );
  NAND2_X1 U13449 ( .A1(n14852), .A2(n14806), .ZN(n11655) );
  NAND2_X1 U13450 ( .A1(n11648), .A2(n11655), .ZN(n11741) );
  AOI211_X1 U13451 ( .C1(n12601), .C2(n11603), .A(n16142), .B(n16323), .ZN(
        n11650) );
  AOI211_X1 U13452 ( .C1(n16366), .C2(n12601), .A(n11741), .B(n11650), .ZN(
        n11604) );
  OAI211_X1 U13453 ( .C1(n11605), .C2(n16369), .A(n11656), .B(n11604), .ZN(
        n11608) );
  NAND2_X1 U13454 ( .A1(n11608), .A2(n16391), .ZN(n11606) );
  OAI21_X1 U13455 ( .B1(n16391), .B2(n11607), .A(n11606), .ZN(P1_U3489) );
  NAND2_X1 U13456 ( .A1(n11608), .A2(n16387), .ZN(n11609) );
  OAI21_X1 U13457 ( .B1(n16387), .B2(n11610), .A(n11609), .ZN(P1_U3538) );
  NAND2_X1 U13458 ( .A1(n11611), .A2(n13618), .ZN(n11612) );
  XNOR2_X1 U13459 ( .A(n16231), .B(n12836), .ZN(n11614) );
  XNOR2_X1 U13460 ( .A(n11614), .B(n13617), .ZN(n11623) );
  NAND2_X1 U13461 ( .A1(n11624), .A2(n11623), .ZN(n11617) );
  INV_X1 U13462 ( .A(n11614), .ZN(n11615) );
  NAND2_X1 U13463 ( .A1(n11615), .A2(n13617), .ZN(n11616) );
  XNOR2_X1 U13464 ( .A(n11678), .B(n12836), .ZN(n11855) );
  XNOR2_X1 U13465 ( .A(n11855), .B(n11860), .ZN(n11853) );
  XNOR2_X1 U13466 ( .A(n11854), .B(n11853), .ZN(n11622) );
  OAI22_X1 U13467 ( .A1(n13575), .A2(n12031), .B1(n11670), .B2(n13600), .ZN(
        n11618) );
  AOI211_X1 U13468 ( .C1(n13606), .C2(n11678), .A(n11619), .B(n11618), .ZN(
        n11621) );
  NAND2_X1 U13469 ( .A1(n13568), .A2(n11677), .ZN(n11620) );
  OAI211_X1 U13470 ( .C1(n11622), .C2(n13608), .A(n11621), .B(n11620), .ZN(
        P3_U3161) );
  XOR2_X1 U13471 ( .A(n11624), .B(n11623), .Z(n11625) );
  NAND2_X1 U13472 ( .A1(n11625), .A2(n13587), .ZN(n11630) );
  OAI22_X1 U13473 ( .A1(n13575), .A2(n11860), .B1(n11626), .B2(n13600), .ZN(
        n11627) );
  AOI211_X1 U13474 ( .C1(n13606), .C2(n12895), .A(n11628), .B(n11627), .ZN(
        n11629) );
  OAI211_X1 U13475 ( .C1(n11631), .C2(n13604), .A(n11630), .B(n11629), .ZN(
        P3_U3153) );
  INV_X1 U13476 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11633) );
  MUX2_X1 U13477 ( .A(n11633), .B(P2_REG2_REG_14__SCAN_IN), .S(n12221), .Z(
        n11634) );
  INV_X1 U13478 ( .A(n11634), .ZN(n11635) );
  NAND2_X1 U13479 ( .A1(n11635), .A2(n11636), .ZN(n12220) );
  OAI21_X1 U13480 ( .B1(n11636), .B2(n11635), .A(n12220), .ZN(n11646) );
  NAND2_X1 U13481 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n11638)
         );
  NAND2_X1 U13482 ( .A1(n15800), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n11637) );
  OAI211_X1 U13483 ( .C1(n14306), .C2(n11639), .A(n11638), .B(n11637), .ZN(
        n11645) );
  INV_X1 U13484 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11641) );
  MUX2_X1 U13485 ( .A(n11641), .B(P2_REG1_REG_14__SCAN_IN), .S(n12221), .Z(
        n11642) );
  AOI211_X1 U13486 ( .C1(n11643), .C2(n11642), .A(n12215), .B(n15813), .ZN(
        n11644) );
  AOI211_X1 U13487 ( .C1(n15830), .C2(n11646), .A(n11645), .B(n11644), .ZN(
        n11647) );
  INV_X1 U13488 ( .A(n11647), .ZN(P2_U3228) );
  INV_X1 U13489 ( .A(n12601), .ZN(n11654) );
  INV_X1 U13490 ( .A(n11648), .ZN(n11649) );
  OAI21_X1 U13491 ( .B1(n11650), .B2(n11649), .A(n16341), .ZN(n11653) );
  AOI22_X1 U13492 ( .A1(n16347), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n11651), 
        .B2(n16336), .ZN(n11652) );
  OAI211_X1 U13493 ( .C1(n11654), .C2(n16163), .A(n11653), .B(n11652), .ZN(
        n11658) );
  AOI21_X1 U13494 ( .B1(n11656), .B2(n11655), .A(n16347), .ZN(n11657) );
  AOI211_X1 U13495 ( .C1(n16342), .C2(n11659), .A(n11658), .B(n11657), .ZN(
        n11660) );
  INV_X1 U13496 ( .A(n11660), .ZN(P1_U3283) );
  AOI211_X1 U13497 ( .C1(n16348), .C2(n11663), .A(n11662), .B(n11661), .ZN(
        n11668) );
  INV_X1 U13498 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11664) );
  NOR2_X1 U13499 ( .A1(n14668), .A2(n11664), .ZN(n11665) );
  AOI21_X1 U13500 ( .B1(n13202), .B2(n11915), .A(n11665), .ZN(n11666) );
  OAI21_X1 U13501 ( .B1(n11668), .B2(n16359), .A(n11666), .ZN(P2_U3466) );
  AOI22_X1 U13502 ( .A1(n13202), .A2(n11917), .B1(n16357), .B2(
        P2_REG1_REG_12__SCAN_IN), .ZN(n11667) );
  OAI21_X1 U13503 ( .B1(n11668), .B2(n16357), .A(n11667), .ZN(P2_U3511) );
  XNOR2_X1 U13504 ( .A(n11669), .B(n13000), .ZN(n16258) );
  OAI22_X1 U13505 ( .A1(n11670), .A2(n16103), .B1(n12031), .B2(n16101), .ZN(
        n11675) );
  NAND2_X1 U13506 ( .A1(n11671), .A2(n13000), .ZN(n11672) );
  AOI21_X1 U13507 ( .B1(n11673), .B2(n11672), .A(n16107), .ZN(n11674) );
  AOI211_X1 U13508 ( .C1(n16258), .C2(n16229), .A(n11675), .B(n11674), .ZN(
        n16256) );
  INV_X2 U13509 ( .A(n16121), .ZN(n16123) );
  INV_X1 U13510 ( .A(n11676), .ZN(n16120) );
  INV_X1 U13511 ( .A(n13871), .ZN(n11681) );
  AOI22_X1 U13512 ( .A1(n13933), .A2(n11678), .B1(n13868), .B2(n11677), .ZN(
        n11679) );
  OAI21_X1 U13513 ( .B1(n8913), .B2(n16121), .A(n11679), .ZN(n11680) );
  AOI21_X1 U13514 ( .B1(n16258), .B2(n11681), .A(n11680), .ZN(n11682) );
  OAI21_X1 U13515 ( .B1(n16256), .B2(n16123), .A(n11682), .ZN(P3_U3225) );
  INV_X1 U13516 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n11683) );
  OAI22_X1 U13517 ( .A1(n16257), .A2(n14102), .B1(n16410), .B2(n11683), .ZN(
        n11684) );
  AOI21_X1 U13518 ( .B1(n16258), .B2(n11685), .A(n11684), .ZN(n11686) );
  OAI21_X1 U13519 ( .B1(n16256), .B2(n16415), .A(n11686), .ZN(P3_U3414) );
  INV_X1 U13520 ( .A(n11687), .ZN(n11690) );
  NAND2_X1 U13521 ( .A1(n11780), .A2(n9720), .ZN(n11693) );
  AOI22_X1 U13522 ( .A1(n11691), .A2(n13109), .B1(n9659), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n11692) );
  NAND2_X2 U13523 ( .A1(n11693), .A2(n11692), .ZN(n16392) );
  XNOR2_X1 U13524 ( .A(n16392), .B(n11516), .ZN(n11695) );
  AND2_X1 U13525 ( .A1(n14254), .A2(n14445), .ZN(n11694) );
  NOR2_X1 U13526 ( .A1(n11695), .A2(n11694), .ZN(n11815) );
  INV_X1 U13527 ( .A(n11815), .ZN(n11696) );
  NAND2_X1 U13528 ( .A1(n11695), .A2(n11694), .ZN(n11814) );
  NAND2_X1 U13529 ( .A1(n11696), .A2(n11814), .ZN(n11697) );
  XNOR2_X1 U13530 ( .A(n11816), .B(n11697), .ZN(n11709) );
  NAND2_X1 U13531 ( .A1(n11698), .A2(n11819), .ZN(n11699) );
  AND2_X1 U13532 ( .A1(n11765), .A2(n11699), .ZN(n11823) );
  NAND2_X1 U13533 ( .A1(n11823), .A2(n11931), .ZN(n11704) );
  NAND2_X1 U13534 ( .A1(n9742), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n11701) );
  NAND2_X1 U13535 ( .A1(n13386), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n11700) );
  AND2_X1 U13536 ( .A1(n11701), .A2(n11700), .ZN(n11703) );
  NAND2_X1 U13537 ( .A1(n13368), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n11702) );
  AOI22_X1 U13538 ( .A1(n14253), .A2(n14439), .B1(n14438), .B2(n14255), .ZN(
        n11909) );
  OAI22_X1 U13539 ( .A1(n14244), .A2(n11909), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11705), .ZN(n11706) );
  AOI21_X1 U13540 ( .B1(n16395), .B2(n14242), .A(n11706), .ZN(n11708) );
  NAND2_X1 U13541 ( .A1(n16392), .A2(n14246), .ZN(n11707) );
  OAI211_X1 U13542 ( .C1(n11709), .C2(n14248), .A(n11708), .B(n11707), .ZN(
        P2_U3206) );
  INV_X1 U13543 ( .A(n11710), .ZN(n11711) );
  NAND2_X1 U13544 ( .A1(n11712), .A2(n11711), .ZN(n11714) );
  NAND2_X1 U13545 ( .A1(n11714), .A2(n11713), .ZN(n11718) );
  MUX2_X1 U13546 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n8006), .Z(n11715) );
  NAND2_X1 U13547 ( .A1(n11715), .A2(SI_24_), .ZN(n12292) );
  OAI21_X1 U13548 ( .B1(SI_24_), .B2(n11715), .A(n12292), .ZN(n11716) );
  INV_X1 U13549 ( .A(n11716), .ZN(n11717) );
  OR2_X1 U13550 ( .A1(n11718), .A2(n11717), .ZN(n11719) );
  NAND2_X1 U13551 ( .A1(n12293), .A2(n11719), .ZN(n13293) );
  OAI222_X1 U13552 ( .A1(n11720), .A2(P1_U3086), .B1(n15260), .B2(n13293), 
        .C1(n7719), .C2(n15262), .ZN(P1_U3331) );
  OAI222_X1 U13553 ( .A1(n11721), .A2(P2_U3088), .B1(n14691), .B2(n13293), 
        .C1(n13294), .C2(n14693), .ZN(P2_U3303) );
  NAND2_X1 U13554 ( .A1(n11723), .A2(n11722), .ZN(n11724) );
  NAND2_X1 U13555 ( .A1(n12592), .A2(n12494), .ZN(n11727) );
  NAND2_X1 U13556 ( .A1(n11727), .A2(n11726), .ZN(n11728) );
  XNOR2_X1 U13557 ( .A(n11728), .B(n12518), .ZN(n11731) );
  NAND2_X1 U13558 ( .A1(n12592), .A2(n8541), .ZN(n11730) );
  NAND2_X1 U13559 ( .A1(n12520), .A2(n14852), .ZN(n11729) );
  NAND2_X1 U13560 ( .A1(n11730), .A2(n11729), .ZN(n11732) );
  NAND2_X1 U13561 ( .A1(n11731), .A2(n11732), .ZN(n11877) );
  NAND2_X1 U13562 ( .A1(n11880), .A2(n11877), .ZN(n11735) );
  INV_X1 U13563 ( .A(n11731), .ZN(n11734) );
  INV_X1 U13564 ( .A(n11732), .ZN(n11733) );
  NAND2_X1 U13565 ( .A1(n11734), .A2(n11733), .ZN(n11878) );
  NAND2_X1 U13566 ( .A1(n12601), .A2(n12494), .ZN(n11737) );
  NAND2_X1 U13567 ( .A1(n8541), .A2(n14851), .ZN(n11736) );
  NAND2_X1 U13568 ( .A1(n11737), .A2(n11736), .ZN(n11738) );
  XNOR2_X1 U13569 ( .A(n11738), .B(n12203), .ZN(n11976) );
  NOR2_X1 U13570 ( .A1(n12483), .A2(n11739), .ZN(n11740) );
  AOI21_X1 U13571 ( .B1(n12601), .B2(n8541), .A(n11740), .ZN(n11977) );
  XNOR2_X1 U13572 ( .A(n11976), .B(n11977), .ZN(n11975) );
  XNOR2_X1 U13573 ( .A(n11974), .B(n11975), .ZN(n11747) );
  NAND2_X1 U13574 ( .A1(n14821), .A2(n11741), .ZN(n11742) );
  OAI211_X1 U13575 ( .C1(n14824), .C2(n11744), .A(n11743), .B(n11742), .ZN(
        n11745) );
  AOI21_X1 U13576 ( .B1(n12601), .B2(n14826), .A(n11745), .ZN(n11746) );
  OAI21_X1 U13577 ( .B1(n11747), .B2(n14829), .A(n11746), .ZN(P1_U3217) );
  OAI21_X1 U13578 ( .B1(n11444), .B2(n11751), .A(n11748), .ZN(n12060) );
  XOR2_X1 U13579 ( .A(n12351), .B(n12060), .Z(n11749) );
  NAND2_X1 U13580 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n11749), .ZN(n12062) );
  OAI211_X1 U13581 ( .C1(n11749), .C2(P1_REG2_REG_18__SCAN_IN), .A(n7422), .B(
        n12062), .ZN(n11758) );
  NAND2_X1 U13582 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14800)
         );
  INV_X1 U13583 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n11750) );
  OAI22_X1 U13584 ( .A1(n11753), .A2(n11752), .B1(n11751), .B2(n11750), .ZN(
        n12056) );
  XNOR2_X1 U13585 ( .A(n11759), .B(n12056), .ZN(n11754) );
  NAND2_X1 U13586 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n11754), .ZN(n12057) );
  OAI211_X1 U13587 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n11754), .A(n16018), 
        .B(n12057), .ZN(n11755) );
  NAND2_X1 U13588 ( .A1(n14800), .A2(n11755), .ZN(n11756) );
  AOI21_X1 U13589 ( .B1(n14866), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n11756), 
        .ZN(n11757) );
  OAI211_X1 U13590 ( .C1(n16022), .C2(n11759), .A(n11758), .B(n11757), .ZN(
        P1_U3261) );
  NAND2_X1 U13591 ( .A1(n12002), .A2(n9720), .ZN(n11761) );
  AOI22_X1 U13592 ( .A1(n12221), .A2(n13109), .B1(n9659), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n11760) );
  AND2_X2 U13593 ( .A1(n11761), .A2(n11760), .ZN(n13216) );
  XNOR2_X1 U13594 ( .A(n13217), .B(n14253), .ZN(n13439) );
  INV_X1 U13595 ( .A(n14255), .ZN(n13204) );
  NAND2_X1 U13596 ( .A1(n13202), .A2(n13204), .ZN(n11763) );
  XNOR2_X1 U13597 ( .A(n16392), .B(n14254), .ZN(n13437) );
  INV_X1 U13598 ( .A(n14254), .ZN(n11764) );
  XOR2_X1 U13599 ( .A(n11836), .B(n13439), .Z(n11768) );
  INV_X1 U13600 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n11959) );
  OR2_X1 U13601 ( .A1(n7554), .A2(n11838), .ZN(n11960) );
  INV_X1 U13602 ( .A(n11931), .ZN(n13309) );
  AOI22_X1 U13603 ( .A1(n9742), .A2(P2_REG1_REG_15__SCAN_IN), .B1(n13386), 
        .B2(P2_REG0_REG_15__SCAN_IN), .ZN(n11767) );
  NAND2_X1 U13604 ( .A1(n13368), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n11766) );
  OAI211_X1 U13605 ( .C1(n11960), .C2(n13309), .A(n11767), .B(n11766), .ZN(
        n14252) );
  AOI22_X1 U13606 ( .A1(n14252), .A2(n14439), .B1(n14438), .B2(n14254), .ZN(
        n11820) );
  OAI21_X1 U13607 ( .B1(n11768), .B2(n14486), .A(n11820), .ZN(n11885) );
  AOI21_X1 U13608 ( .B1(n11823), .B2(n16394), .A(n11885), .ZN(n11777) );
  INV_X1 U13609 ( .A(n11906), .ZN(n11770) );
  NAND2_X1 U13610 ( .A1(n13216), .A2(n11906), .ZN(n11846) );
  INV_X1 U13611 ( .A(n11846), .ZN(n11769) );
  AOI211_X1 U13612 ( .C1(n13217), .C2(n11770), .A(n14445), .B(n11769), .ZN(
        n11886) );
  OAI22_X1 U13613 ( .A1(n13216), .A2(n16398), .B1(n14549), .B2(n11633), .ZN(
        n11771) );
  AOI21_X1 U13614 ( .B1(n11886), .B2(n16306), .A(n11771), .ZN(n11776) );
  NAND2_X1 U13615 ( .A1(n13202), .A2(n14255), .ZN(n11773) );
  NAND2_X1 U13616 ( .A1(n16392), .A2(n14254), .ZN(n11774) );
  XNOR2_X1 U13617 ( .A(n11826), .B(n13439), .ZN(n11887) );
  NAND2_X1 U13618 ( .A1(n11887), .A2(n14515), .ZN(n11775) );
  OAI211_X1 U13619 ( .C1(n11777), .C2(n16405), .A(n11776), .B(n11775), .ZN(
        P2_U3251) );
  INV_X1 U13620 ( .A(n14849), .ZN(n12120) );
  OR2_X1 U13621 ( .A1(n16365), .A2(n12120), .ZN(n11778) );
  NAND2_X1 U13622 ( .A1(n11779), .A2(n11778), .ZN(n11784) );
  AOI22_X1 U13623 ( .A1(n11781), .A2(n12398), .B1(n12399), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n11782) );
  INV_X1 U13624 ( .A(n14848), .ZN(n12205) );
  XNOR2_X1 U13625 ( .A(n12616), .B(n12205), .ZN(n12738) );
  OAI21_X1 U13626 ( .B1(n11784), .B2(n11783), .A(n12001), .ZN(n16380) );
  NAND2_X1 U13627 ( .A1(n11786), .A2(n11785), .ZN(n11788) );
  OR2_X1 U13628 ( .A1(n16365), .A2(n14849), .ZN(n11787) );
  XNOR2_X1 U13629 ( .A(n12005), .B(n12738), .ZN(n16384) );
  NAND2_X1 U13630 ( .A1(n16384), .A2(n15058), .ZN(n11801) );
  NAND2_X1 U13631 ( .A1(n7426), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11795) );
  AND2_X1 U13632 ( .A1(n11790), .A2(n11789), .ZN(n11791) );
  NOR2_X1 U13633 ( .A1(n12013), .A2(n11791), .ZN(n14710) );
  NAND2_X1 U13634 ( .A1(n14710), .A2(n12526), .ZN(n11794) );
  NAND2_X1 U13635 ( .A1(n10089), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11793) );
  NAND2_X1 U13636 ( .A1(n12686), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n11792) );
  NAND4_X1 U13637 ( .A1(n11795), .A2(n11794), .A3(n11793), .A4(n11792), .ZN(
        n14847) );
  AOI22_X1 U13638 ( .A1(n14807), .A2(n14847), .B1(n14849), .B2(n14806), .ZN(
        n16376) );
  INV_X1 U13639 ( .A(n16376), .ZN(n11796) );
  AOI22_X1 U13640 ( .A1(n16086), .A2(n11796), .B1(n12212), .B2(n16336), .ZN(
        n11797) );
  OAI21_X1 U13641 ( .B1(n11184), .B2(n16159), .A(n11797), .ZN(n11799) );
  OAI211_X1 U13642 ( .C1(n7671), .C2(n7672), .A(n16322), .B(n12010), .ZN(
        n16377) );
  NOR2_X1 U13643 ( .A1(n16377), .A2(n15051), .ZN(n11798) );
  AOI211_X1 U13644 ( .C1(n16337), .C2(n12616), .A(n11799), .B(n11798), .ZN(
        n11800) );
  OAI211_X1 U13645 ( .C1(n16380), .C2(n15070), .A(n11801), .B(n11800), .ZN(
        P1_U3280) );
  INV_X1 U13646 ( .A(n12907), .ZN(n11802) );
  NOR2_X1 U13647 ( .A1(n11802), .A2(n12905), .ZN(n12998) );
  XNOR2_X1 U13648 ( .A(n11803), .B(n12998), .ZN(n11806) );
  INV_X1 U13649 ( .A(n11806), .ZN(n16275) );
  XNOR2_X1 U13650 ( .A(n11804), .B(n12998), .ZN(n11808) );
  OAI22_X1 U13651 ( .A1(n12910), .A2(n16101), .B1(n11860), .B2(n16103), .ZN(
        n11805) );
  AOI21_X1 U13652 ( .B1(n11806), .B2(n16229), .A(n11805), .ZN(n11807) );
  OAI21_X1 U13653 ( .B1(n11808), .B2(n16107), .A(n11807), .ZN(n16277) );
  NAND2_X1 U13654 ( .A1(n16277), .A2(n16121), .ZN(n11811) );
  OAI22_X1 U13655 ( .A1(n16273), .A2(n13963), .B1(n11864), .B2(n16113), .ZN(
        n11809) );
  AOI21_X1 U13656 ( .B1(n16123), .B2(P3_REG2_REG_9__SCAN_IN), .A(n11809), .ZN(
        n11810) );
  OAI211_X1 U13657 ( .C1(n16275), .C2(n13871), .A(n11811), .B(n11810), .ZN(
        P3_U3224) );
  XNOR2_X1 U13658 ( .A(n13216), .B(n11516), .ZN(n11813) );
  NAND2_X1 U13659 ( .A1(n14253), .A2(n14445), .ZN(n11812) );
  NAND2_X1 U13660 ( .A1(n11813), .A2(n11812), .ZN(n11956) );
  OAI21_X1 U13661 ( .B1(n11813), .B2(n11812), .A(n11956), .ZN(n11818) );
  AOI21_X1 U13662 ( .B1(n11818), .B2(n11817), .A(n11958), .ZN(n11825) );
  OAI22_X1 U13663 ( .A1(n14244), .A2(n11820), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11819), .ZN(n11822) );
  NOR2_X1 U13664 ( .A1(n13216), .A2(n12244), .ZN(n11821) );
  AOI211_X1 U13665 ( .C1(n14242), .C2(n11823), .A(n11822), .B(n11821), .ZN(
        n11824) );
  OAI21_X1 U13666 ( .B1(n11825), .B2(n14248), .A(n11824), .ZN(P2_U3187) );
  NAND2_X1 U13667 ( .A1(n13216), .A2(n13215), .ZN(n11827) );
  NAND2_X1 U13668 ( .A1(n12075), .A2(n9720), .ZN(n11833) );
  OAI22_X1 U13669 ( .A1(n15836), .A2(n11830), .B1(n8004), .B2(n11829), .ZN(
        n11831) );
  INV_X1 U13670 ( .A(n11831), .ZN(n11832) );
  INV_X1 U13671 ( .A(n14252), .ZN(n13222) );
  XNOR2_X1 U13672 ( .A(n13221), .B(n13222), .ZN(n13441) );
  OAI21_X1 U13673 ( .B1(n11834), .B2(n13441), .A(n11947), .ZN(n12136) );
  INV_X1 U13674 ( .A(n12136), .ZN(n11852) );
  NOR2_X1 U13675 ( .A1(n13216), .A2(n14253), .ZN(n11835) );
  NAND2_X1 U13676 ( .A1(n13216), .A2(n14253), .ZN(n11837) );
  XNOR2_X1 U13677 ( .A(n11920), .B(n7816), .ZN(n11845) );
  OR2_X1 U13678 ( .A1(n11838), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n11839) );
  NAND2_X1 U13679 ( .A1(n11838), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n11929) );
  AND2_X1 U13680 ( .A1(n11839), .A2(n11929), .ZN(n12150) );
  NAND2_X1 U13681 ( .A1(n12150), .A2(n9789), .ZN(n11842) );
  AOI22_X1 U13682 ( .A1(n9742), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n13386), 
        .B2(P2_REG0_REG_16__SCAN_IN), .ZN(n11841) );
  NAND2_X1 U13683 ( .A1(n13368), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n11840) );
  OAI22_X1 U13684 ( .A1(n13226), .A2(n14523), .B1(n13215), .B2(n14521), .ZN(
        n11843) );
  AOI21_X1 U13685 ( .B1(n12136), .B2(n14520), .A(n11843), .ZN(n11844) );
  OAI21_X1 U13686 ( .B1(n14486), .B2(n11845), .A(n11844), .ZN(n12134) );
  NAND2_X1 U13687 ( .A1(n12134), .A2(n14549), .ZN(n11851) );
  AOI211_X1 U13688 ( .C1(n13221), .C2(n11846), .A(n14445), .B(n12048), .ZN(
        n12135) );
  INV_X1 U13689 ( .A(n13221), .ZN(n13223) );
  INV_X1 U13690 ( .A(n11960), .ZN(n11847) );
  AOI22_X1 U13691 ( .A1(n16405), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n11847), 
        .B2(n16394), .ZN(n11848) );
  OAI21_X1 U13692 ( .B1(n13223), .B2(n16398), .A(n11848), .ZN(n11849) );
  AOI21_X1 U13693 ( .B1(n12135), .B2(n16306), .A(n11849), .ZN(n11850) );
  OAI211_X1 U13694 ( .C1(n11852), .C2(n14452), .A(n11851), .B(n11850), .ZN(
        P2_U3250) );
  XNOR2_X1 U13695 ( .A(n11863), .B(n8025), .ZN(n11893) );
  XNOR2_X1 U13696 ( .A(n11893), .B(n12031), .ZN(n11859) );
  NAND2_X1 U13697 ( .A1(n13616), .A2(n11855), .ZN(n11856) );
  INV_X1 U13698 ( .A(n11896), .ZN(n11857) );
  AOI21_X1 U13699 ( .B1(n11859), .B2(n11858), .A(n11857), .ZN(n11868) );
  OAI22_X1 U13700 ( .A1(n13575), .A2(n12910), .B1(n11860), .B2(n13600), .ZN(
        n11861) );
  AOI211_X1 U13701 ( .C1(n13606), .C2(n11863), .A(n11862), .B(n11861), .ZN(
        n11867) );
  INV_X1 U13702 ( .A(n11864), .ZN(n11865) );
  NAND2_X1 U13703 ( .A1(n13568), .A2(n11865), .ZN(n11866) );
  OAI211_X1 U13704 ( .C1(n11868), .C2(n13608), .A(n11867), .B(n11866), .ZN(
        P3_U3171) );
  INV_X1 U13705 ( .A(n11869), .ZN(n11870) );
  INV_X1 U13706 ( .A(SI_27_), .ZN(n15460) );
  OAI222_X1 U13707 ( .A1(P3_U3151), .A2(n8634), .B1(n14119), .B2(n11870), .C1(
        n15460), .C2(n13462), .ZN(P3_U3268) );
  INV_X1 U13708 ( .A(SI_28_), .ZN(n12305) );
  INV_X1 U13709 ( .A(n11871), .ZN(n11872) );
  OAI222_X1 U13710 ( .A1(n13462), .A2(n12305), .B1(P3_U3151), .B2(n13037), 
        .C1(n14119), .C2(n11872), .ZN(P3_U3267) );
  NAND2_X1 U13711 ( .A1(n14811), .A2(n11873), .ZN(n11875) );
  OAI211_X1 U13712 ( .C1(n11876), .C2(n14809), .A(n11875), .B(n11874), .ZN(
        n11883) );
  NAND2_X1 U13713 ( .A1(n11878), .A2(n11877), .ZN(n11879) );
  XNOR2_X1 U13714 ( .A(n11880), .B(n11879), .ZN(n11881) );
  NOR2_X1 U13715 ( .A1(n11881), .A2(n14829), .ZN(n11882) );
  AOI211_X1 U13716 ( .C1(n12592), .C2(n14826), .A(n11883), .B(n11882), .ZN(
        n11884) );
  INV_X1 U13717 ( .A(n11884), .ZN(P1_U3231) );
  AOI211_X1 U13718 ( .C1(n16348), .C2(n11887), .A(n11886), .B(n11885), .ZN(
        n11892) );
  INV_X1 U13719 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n11888) );
  OAI22_X1 U13720 ( .A1(n13216), .A2(n14673), .B1(n14668), .B2(n11888), .ZN(
        n11889) );
  INV_X1 U13721 ( .A(n11889), .ZN(n11890) );
  OAI21_X1 U13722 ( .B1(n11892), .B2(n16359), .A(n11890), .ZN(P2_U3472) );
  AOI22_X1 U13723 ( .A1(n13217), .A2(n11917), .B1(n16357), .B2(
        P2_REG1_REG_14__SCAN_IN), .ZN(n11891) );
  OAI21_X1 U13724 ( .B1(n11892), .B2(n16357), .A(n11891), .ZN(P2_U3513) );
  NAND2_X1 U13725 ( .A1(n11893), .A2(n12031), .ZN(n11894) );
  AND2_X1 U13726 ( .A1(n11896), .A2(n11894), .ZN(n11898) );
  XNOR2_X1 U13727 ( .A(n16295), .B(n12836), .ZN(n12096) );
  XNOR2_X1 U13728 ( .A(n12096), .B(n13614), .ZN(n11897) );
  AND2_X1 U13729 ( .A1(n11897), .A2(n11894), .ZN(n11895) );
  OAI211_X1 U13730 ( .C1(n11898), .C2(n11897), .A(n13587), .B(n12099), .ZN(
        n11904) );
  AOI21_X1 U13731 ( .B1(n13602), .B2(n13613), .A(n11899), .ZN(n11901) );
  NAND2_X1 U13732 ( .A1(n13589), .A2(n13615), .ZN(n11900) );
  OAI211_X1 U13733 ( .C1(n13595), .C2(n16295), .A(n11901), .B(n11900), .ZN(
        n11902) );
  INV_X1 U13734 ( .A(n11902), .ZN(n11903) );
  OAI211_X1 U13735 ( .C1(n12035), .C2(n13604), .A(n11904), .B(n11903), .ZN(
        P3_U3157) );
  XNOR2_X1 U13736 ( .A(n11905), .B(n13437), .ZN(n16402) );
  AOI211_X1 U13737 ( .C1(n16392), .C2(n11907), .A(n7431), .B(n11906), .ZN(
        n16393) );
  XNOR2_X1 U13738 ( .A(n11908), .B(n7782), .ZN(n11910) );
  OAI21_X1 U13739 ( .B1(n11910), .B2(n14486), .A(n11909), .ZN(n11911) );
  AOI21_X1 U13740 ( .B1(n16402), .B2(n14520), .A(n11911), .ZN(n16404) );
  INV_X1 U13741 ( .A(n16404), .ZN(n11912) );
  AOI211_X1 U13742 ( .C1(n13099), .C2(n16402), .A(n16393), .B(n11912), .ZN(
        n11919) );
  INV_X1 U13743 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11913) );
  NOR2_X1 U13744 ( .A1(n14668), .A2(n11913), .ZN(n11914) );
  AOI21_X1 U13745 ( .B1(n16392), .B2(n11915), .A(n11914), .ZN(n11916) );
  OAI21_X1 U13746 ( .B1(n11919), .B2(n16359), .A(n11916), .ZN(P2_U3469) );
  AOI22_X1 U13747 ( .A1(n16392), .A2(n11917), .B1(n16357), .B2(
        P2_REG1_REG_13__SCAN_IN), .ZN(n11918) );
  OAI21_X1 U13748 ( .B1(n11919), .B2(n16357), .A(n11918), .ZN(P2_U3512) );
  OR2_X1 U13749 ( .A1(n13221), .A2(n13222), .ZN(n11921) );
  NAND2_X1 U13750 ( .A1(n11922), .A2(n11921), .ZN(n12040) );
  NAND2_X1 U13751 ( .A1(n12175), .A2(n9720), .ZN(n11924) );
  AOI22_X1 U13752 ( .A1(n9659), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n13109), 
        .B2(n14273), .ZN(n11923) );
  NAND2_X1 U13753 ( .A1(n13227), .A2(n14251), .ZN(n11925) );
  NAND2_X1 U13754 ( .A1(n12248), .A2(n9720), .ZN(n11927) );
  AOI22_X1 U13755 ( .A1(n9659), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n13109), 
        .B2(n14288), .ZN(n11926) );
  INV_X1 U13756 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n11928) );
  NAND2_X1 U13757 ( .A1(n11929), .A2(n11928), .ZN(n11930) );
  AND2_X1 U13758 ( .A1(n12279), .A2(n11930), .ZN(n11950) );
  NAND2_X1 U13759 ( .A1(n11950), .A2(n11931), .ZN(n11936) );
  INV_X1 U13760 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n14629) );
  NAND2_X1 U13761 ( .A1(n13386), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n11933) );
  NAND2_X1 U13762 ( .A1(n13368), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11932) );
  OAI211_X1 U13763 ( .C1(n14629), .C2(n13346), .A(n11933), .B(n11932), .ZN(
        n11934) );
  INV_X1 U13764 ( .A(n11934), .ZN(n11935) );
  NAND2_X1 U13765 ( .A1(n11936), .A2(n11935), .ZN(n14324) );
  XNOR2_X1 U13766 ( .A(n14336), .B(n14324), .ZN(n14338) );
  INV_X1 U13767 ( .A(n14338), .ZN(n11937) );
  XNOR2_X1 U13768 ( .A(n14339), .B(n11937), .ZN(n11945) );
  XNOR2_X1 U13769 ( .A(n12279), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n14540) );
  NAND2_X1 U13770 ( .A1(n14540), .A2(n9789), .ZN(n11943) );
  INV_X1 U13771 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n11940) );
  NAND2_X1 U13772 ( .A1(n9742), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n11939) );
  NAND2_X1 U13773 ( .A1(n13386), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n11938) );
  OAI211_X1 U13774 ( .C1(n11940), .C2(n9829), .A(n11939), .B(n11938), .ZN(
        n11941) );
  INV_X1 U13775 ( .A(n11941), .ZN(n11942) );
  OAI22_X1 U13776 ( .A1(n14326), .A2(n14523), .B1(n13226), .B2(n14521), .ZN(
        n11944) );
  AOI21_X1 U13777 ( .B1(n11945), .B2(n14529), .A(n11944), .ZN(n14626) );
  OR2_X1 U13778 ( .A1(n13221), .A2(n14252), .ZN(n11946) );
  OR2_X1 U13779 ( .A1(n13227), .A2(n13226), .ZN(n11948) );
  XNOR2_X1 U13780 ( .A(n14323), .B(n14338), .ZN(n14624) );
  NAND2_X1 U13781 ( .A1(n14336), .A2(n12049), .ZN(n11949) );
  NAND3_X1 U13782 ( .A1(n14535), .A2(n14507), .A3(n11949), .ZN(n14625) );
  INV_X1 U13783 ( .A(n11950), .ZN(n12240) );
  NAND2_X1 U13784 ( .A1(n16405), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11951) );
  OAI21_X1 U13785 ( .B1(n14510), .B2(n12240), .A(n11951), .ZN(n11952) );
  AOI21_X1 U13786 ( .B1(n14336), .B2(n16303), .A(n11952), .ZN(n11953) );
  OAI21_X1 U13787 ( .B1(n14625), .B2(n14539), .A(n11953), .ZN(n11954) );
  AOI21_X1 U13788 ( .B1(n14624), .B2(n14515), .A(n11954), .ZN(n11955) );
  OAI21_X1 U13789 ( .B1(n16405), .B2(n14626), .A(n11955), .ZN(P2_U3248) );
  INV_X1 U13790 ( .A(n11956), .ZN(n11957) );
  XNOR2_X1 U13791 ( .A(n13221), .B(n11516), .ZN(n12144) );
  NAND2_X1 U13792 ( .A1(n14252), .A2(n7431), .ZN(n12143) );
  XNOR2_X1 U13793 ( .A(n12144), .B(n12143), .ZN(n12146) );
  XNOR2_X1 U13794 ( .A(n7580), .B(n12146), .ZN(n11964) );
  OAI22_X1 U13795 ( .A1(n14217), .A2(n13226), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11959), .ZN(n11962) );
  OAI22_X1 U13796 ( .A1(n14219), .A2(n13215), .B1(n11960), .B2(n14218), .ZN(
        n11961) );
  AOI211_X1 U13797 ( .C1(n13221), .C2(n14246), .A(n11962), .B(n11961), .ZN(
        n11963) );
  OAI21_X1 U13798 ( .B1(n11964), .B2(n14248), .A(n11963), .ZN(P2_U3213) );
  OAI22_X1 U13799 ( .A1(n16324), .A2(n8012), .B1(n12606), .B2(n10228), .ZN(
        n11966) );
  XNOR2_X1 U13800 ( .A(n11966), .B(n12203), .ZN(n11969) );
  OR2_X1 U13801 ( .A1(n16324), .A2(n10228), .ZN(n11968) );
  NAND2_X1 U13802 ( .A1(n12520), .A2(n14850), .ZN(n11967) );
  AND2_X1 U13803 ( .A1(n11968), .A2(n11967), .ZN(n11970) );
  NAND2_X1 U13804 ( .A1(n11969), .A2(n11970), .ZN(n12122) );
  INV_X1 U13805 ( .A(n11969), .ZN(n11972) );
  INV_X1 U13806 ( .A(n11970), .ZN(n11971) );
  NAND2_X1 U13807 ( .A1(n11972), .A2(n11971), .ZN(n11973) );
  NAND2_X1 U13808 ( .A1(n12122), .A2(n11973), .ZN(n11985) );
  INV_X1 U13809 ( .A(n11976), .ZN(n11979) );
  INV_X1 U13810 ( .A(n11977), .ZN(n11978) );
  NAND2_X1 U13811 ( .A1(n11979), .A2(n11978), .ZN(n11980) );
  INV_X1 U13812 ( .A(n11985), .ZN(n11982) );
  INV_X1 U13813 ( .A(n12123), .ZN(n11983) );
  AOI21_X1 U13814 ( .B1(n11985), .B2(n11984), .A(n11983), .ZN(n11990) );
  AOI22_X1 U13815 ( .A1(n14806), .A2(n14851), .B1(n14849), .B2(n14799), .ZN(
        n16327) );
  NAND2_X1 U13816 ( .A1(n14811), .A2(n16335), .ZN(n11987) );
  OAI211_X1 U13817 ( .C1(n16327), .C2(n14809), .A(n11987), .B(n11986), .ZN(
        n11988) );
  AOI21_X1 U13818 ( .B1(n16338), .B2(n14826), .A(n11988), .ZN(n11989) );
  OAI21_X1 U13819 ( .B1(n11990), .B2(n14829), .A(n11989), .ZN(P1_U3236) );
  INV_X1 U13820 ( .A(n13008), .ZN(n12913) );
  XNOR2_X1 U13821 ( .A(n11991), .B(n12913), .ZN(n11992) );
  OAI222_X1 U13822 ( .A1(n16101), .A2(n13959), .B1(n16103), .B2(n12910), .C1(
        n11992), .C2(n16107), .ZN(n16313) );
  INV_X1 U13823 ( .A(n16313), .ZN(n11999) );
  OAI21_X1 U13824 ( .B1(n11994), .B2(n13008), .A(n11993), .ZN(n16315) );
  NOR2_X1 U13825 ( .A1(n13963), .A2(n16312), .ZN(n11997) );
  OAI22_X1 U13826 ( .A1(n16121), .A2(n11995), .B1(n12103), .B2(n16113), .ZN(
        n11996) );
  AOI211_X1 U13827 ( .C1(n16315), .C2(n13967), .A(n11997), .B(n11996), .ZN(
        n11998) );
  OAI21_X1 U13828 ( .B1(n11999), .B2(n16123), .A(n11998), .ZN(P3_U3222) );
  OR2_X1 U13829 ( .A1(n12616), .A2(n12205), .ZN(n12000) );
  NAND2_X1 U13830 ( .A1(n12002), .A2(n12491), .ZN(n12004) );
  AOI22_X1 U13831 ( .A1(n14901), .A2(n12398), .B1(n12399), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n12003) );
  XNOR2_X1 U13832 ( .A(n14705), .B(n14847), .ZN(n12739) );
  XNOR2_X1 U13833 ( .A(n12074), .B(n12739), .ZN(n15217) );
  OR2_X1 U13834 ( .A1(n12616), .A2(n14848), .ZN(n12006) );
  INV_X1 U13835 ( .A(n12080), .ZN(n12008) );
  AOI21_X1 U13836 ( .B1(n12739), .B2(n12009), .A(n12008), .ZN(n15215) );
  NAND2_X1 U13837 ( .A1(n15215), .A2(n15058), .ZN(n12026) );
  NAND2_X1 U13838 ( .A1(n14705), .A2(n12010), .ZN(n12011) );
  NAND2_X1 U13839 ( .A1(n12011), .A2(n16322), .ZN(n12012) );
  NOR2_X1 U13840 ( .A1(n12081), .A2(n12012), .ZN(n15214) );
  NAND2_X1 U13841 ( .A1(n14705), .A2(n16337), .ZN(n12023) );
  NAND2_X1 U13842 ( .A1(n12013), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n12083) );
  OR2_X1 U13843 ( .A1(n12013), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n12014) );
  NAND2_X1 U13844 ( .A1(n12083), .A2(n12014), .ZN(n14823) );
  INV_X1 U13845 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n12092) );
  OAI22_X1 U13846 ( .A1(n14823), .A2(n12334), .B1(n12431), .B2(n12092), .ZN(
        n12020) );
  INV_X1 U13847 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n12017) );
  INV_X1 U13848 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n12015) );
  OAI22_X1 U13849 ( .A1(n12018), .A2(n12017), .B1(n12016), .B2(n12015), .ZN(
        n12019) );
  AOI22_X1 U13850 ( .A1(n14799), .A2(n14846), .B1(n14848), .B2(n14806), .ZN(
        n15211) );
  INV_X1 U13851 ( .A(n15211), .ZN(n12021) );
  AOI22_X1 U13852 ( .A1(n16086), .A2(n12021), .B1(n14710), .B2(n16336), .ZN(
        n12022) );
  OAI211_X1 U13853 ( .C1(n11186), .C2(n16159), .A(n12023), .B(n12022), .ZN(
        n12024) );
  AOI21_X1 U13854 ( .B1(n15214), .B2(n16341), .A(n12024), .ZN(n12025) );
  OAI211_X1 U13855 ( .C1(n15217), .C2(n15070), .A(n12026), .B(n12025), .ZN(
        P1_U3279) );
  NAND2_X1 U13856 ( .A1(n12027), .A2(n13011), .ZN(n12028) );
  NAND2_X1 U13857 ( .A1(n12029), .A2(n12028), .ZN(n16298) );
  INV_X1 U13858 ( .A(n16298), .ZN(n12039) );
  XNOR2_X1 U13859 ( .A(n12030), .B(n13011), .ZN(n12034) );
  OAI22_X1 U13860 ( .A1(n12031), .A2(n16103), .B1(n8384), .B2(n16101), .ZN(
        n12032) );
  AOI21_X1 U13861 ( .B1(n16298), .B2(n16229), .A(n12032), .ZN(n12033) );
  OAI21_X1 U13862 ( .B1(n12034), .B2(n16107), .A(n12033), .ZN(n16296) );
  NAND2_X1 U13863 ( .A1(n16296), .A2(n16121), .ZN(n12038) );
  OAI22_X1 U13864 ( .A1(n13963), .A2(n16295), .B1(n12035), .B2(n16113), .ZN(
        n12036) );
  AOI21_X1 U13865 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n16123), .A(n12036), 
        .ZN(n12037) );
  OAI211_X1 U13866 ( .C1(n12039), .C2(n13871), .A(n12038), .B(n12037), .ZN(
        P3_U3223) );
  XOR2_X1 U13867 ( .A(n12040), .B(n13442), .Z(n12047) );
  NAND2_X1 U13868 ( .A1(n12041), .A2(n13442), .ZN(n12042) );
  NAND2_X1 U13869 ( .A1(n12043), .A2(n12042), .ZN(n14636) );
  AOI22_X1 U13870 ( .A1(n14324), .A2(n14439), .B1(n14438), .B2(n14252), .ZN(
        n12044) );
  OAI21_X1 U13871 ( .B1(n14636), .B2(n12045), .A(n12044), .ZN(n12046) );
  AOI21_X1 U13872 ( .B1(n12047), .B2(n14529), .A(n12046), .ZN(n14635) );
  INV_X1 U13873 ( .A(n12048), .ZN(n12051) );
  INV_X1 U13874 ( .A(n12049), .ZN(n12050) );
  AOI211_X1 U13875 ( .C1(n14633), .C2(n12051), .A(n14445), .B(n12050), .ZN(
        n14632) );
  AOI22_X1 U13876 ( .A1(n16405), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n12150), 
        .B2(n16394), .ZN(n12052) );
  OAI21_X1 U13877 ( .B1(n13227), .B2(n16398), .A(n12052), .ZN(n12054) );
  NOR2_X1 U13878 ( .A1(n14636), .A2(n14452), .ZN(n12053) );
  AOI211_X1 U13879 ( .C1(n14632), .C2(n16306), .A(n12054), .B(n12053), .ZN(
        n12055) );
  OAI21_X1 U13880 ( .B1(n16405), .B2(n14635), .A(n12055), .ZN(P2_U3249) );
  NAND2_X1 U13881 ( .A1(n12351), .A2(n12056), .ZN(n12058) );
  NAND2_X1 U13882 ( .A1(n12058), .A2(n12057), .ZN(n12059) );
  XOR2_X1 U13883 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n12059), .Z(n12069) );
  NAND2_X1 U13884 ( .A1(n12351), .A2(n12060), .ZN(n12061) );
  NAND2_X1 U13885 ( .A1(n12062), .A2(n12061), .ZN(n12063) );
  XOR2_X1 U13886 ( .A(n12063), .B(P1_REG2_REG_19__SCAN_IN), .Z(n12068) );
  INV_X1 U13887 ( .A(n12068), .ZN(n12065) );
  NAND2_X1 U13888 ( .A1(n12065), .A2(n12064), .ZN(n12066) );
  OAI211_X1 U13889 ( .C1(n12069), .C2(n15852), .A(n12066), .B(n16022), .ZN(
        n12067) );
  INV_X1 U13890 ( .A(n12067), .ZN(n12071) );
  AOI22_X1 U13891 ( .A1(n12069), .A2(n16018), .B1(n7422), .B2(n12068), .ZN(
        n12070) );
  MUX2_X1 U13892 ( .A(n12071), .B(n12070), .S(n12752), .Z(n12072) );
  NAND2_X1 U13893 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14724)
         );
  OAI211_X1 U13894 ( .C1(n8795), .C2(n16028), .A(n12072), .B(n14724), .ZN(
        P1_U3262) );
  INV_X1 U13895 ( .A(n14847), .ZN(n12366) );
  NAND2_X1 U13896 ( .A1(n14705), .A2(n12366), .ZN(n12073) );
  NAND2_X1 U13897 ( .A1(n12075), .A2(n12491), .ZN(n12078) );
  AOI22_X1 U13898 ( .A1(n12399), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n12398), 
        .B2(n12076), .ZN(n12077) );
  XNOR2_X1 U13899 ( .A(n14827), .B(n14846), .ZN(n12740) );
  XNOR2_X1 U13900 ( .A(n12179), .B(n12740), .ZN(n15210) );
  NAND2_X1 U13901 ( .A1(n14705), .A2(n14847), .ZN(n12079) );
  OAI21_X1 U13902 ( .B1(n7586), .B2(n8673), .A(n12174), .ZN(n15208) );
  INV_X1 U13903 ( .A(n14827), .ZN(n15206) );
  OAI211_X1 U13904 ( .C1(n15206), .C2(n12081), .A(n16322), .B(n12182), .ZN(
        n15205) );
  NOR2_X1 U13905 ( .A1(n15205), .A2(n15051), .ZN(n12094) );
  NAND2_X1 U13906 ( .A1(n14827), .A2(n16337), .ZN(n12091) );
  INV_X1 U13907 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n12082) );
  NAND2_X1 U13908 ( .A1(n12083), .A2(n12082), .ZN(n12084) );
  NAND2_X1 U13909 ( .A1(n12185), .A2(n12084), .ZN(n14750) );
  AOI22_X1 U13910 ( .A1(n12524), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n7426), 
        .B2(P1_REG2_REG_16__SCAN_IN), .ZN(n12086) );
  NAND2_X1 U13911 ( .A1(n12686), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n12085) );
  OAI211_X1 U13912 ( .C1(n14750), .C2(n12334), .A(n12086), .B(n12085), .ZN(
        n14845) );
  NAND2_X1 U13913 ( .A1(n14845), .A2(n14799), .ZN(n12088) );
  NAND2_X1 U13914 ( .A1(n14847), .A2(n14806), .ZN(n12087) );
  NAND2_X1 U13915 ( .A1(n12088), .A2(n12087), .ZN(n15203) );
  NOR2_X1 U13916 ( .A1(n16161), .A2(n14823), .ZN(n12089) );
  AOI21_X1 U13917 ( .B1(n16159), .B2(n15203), .A(n12089), .ZN(n12090) );
  OAI211_X1 U13918 ( .C1(n16159), .C2(n12092), .A(n12091), .B(n12090), .ZN(
        n12093) );
  AOI211_X1 U13919 ( .C1(n15208), .C2(n15058), .A(n12094), .B(n12093), .ZN(
        n12095) );
  OAI21_X1 U13920 ( .B1(n15070), .B2(n15210), .A(n12095), .ZN(P1_U3278) );
  INV_X1 U13921 ( .A(n12096), .ZN(n12097) );
  NAND2_X1 U13922 ( .A1(n12097), .A2(n13614), .ZN(n12098) );
  NAND2_X1 U13923 ( .A1(n12099), .A2(n12098), .ZN(n12158) );
  XNOR2_X1 U13924 ( .A(n16312), .B(n12836), .ZN(n12159) );
  XNOR2_X1 U13925 ( .A(n12159), .B(n13613), .ZN(n12157) );
  XOR2_X1 U13926 ( .A(n12158), .B(n12157), .Z(n12106) );
  NOR2_X1 U13927 ( .A1(n13595), .A2(n16312), .ZN(n12105) );
  AOI21_X1 U13928 ( .B1(n13602), .B2(n13612), .A(n12100), .ZN(n12102) );
  NAND2_X1 U13929 ( .A1(n13589), .A2(n13614), .ZN(n12101) );
  OAI211_X1 U13930 ( .C1(n12103), .C2(n13604), .A(n12102), .B(n12101), .ZN(
        n12104) );
  AOI211_X1 U13931 ( .C1(n12106), .C2(n13587), .A(n12105), .B(n12104), .ZN(
        n12107) );
  INV_X1 U13932 ( .A(n12107), .ZN(P3_U3176) );
  OR2_X1 U13933 ( .A1(n12108), .A2(n13010), .ZN(n12109) );
  NAND2_X1 U13934 ( .A1(n12110), .A2(n12109), .ZN(n14034) );
  INV_X1 U13935 ( .A(n14034), .ZN(n14107) );
  XNOR2_X1 U13936 ( .A(n12111), .B(n13010), .ZN(n12112) );
  OAI222_X1 U13937 ( .A1(n16103), .A2(n8384), .B1(n16101), .B2(n13475), .C1(
        n16107), .C2(n12112), .ZN(n14032) );
  NAND2_X1 U13938 ( .A1(n14032), .A2(n16121), .ZN(n12116) );
  INV_X1 U13939 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12113) );
  OAI22_X1 U13940 ( .A1(n16121), .A2(n12113), .B1(n12165), .B2(n16113), .ZN(
        n12114) );
  AOI21_X1 U13941 ( .B1(n12156), .B2(n13933), .A(n12114), .ZN(n12115) );
  OAI211_X1 U13942 ( .C1(n14107), .C2(n13937), .A(n12116), .B(n12115), .ZN(
        P3_U3221) );
  NAND2_X1 U13943 ( .A1(n16365), .A2(n12494), .ZN(n12118) );
  NAND2_X1 U13944 ( .A1(n12118), .A2(n12117), .ZN(n12119) );
  XNOR2_X1 U13945 ( .A(n12119), .B(n12518), .ZN(n12196) );
  NOR2_X1 U13946 ( .A1(n12483), .A2(n12120), .ZN(n12121) );
  AOI21_X1 U13947 ( .B1(n16365), .B2(n8541), .A(n12121), .ZN(n12197) );
  XNOR2_X1 U13948 ( .A(n12196), .B(n12197), .ZN(n12125) );
  OAI21_X1 U13949 ( .B1(n12125), .B2(n12124), .A(n12200), .ZN(n12126) );
  NAND2_X1 U13950 ( .A1(n12126), .A2(n14796), .ZN(n12132) );
  OAI21_X1 U13951 ( .B1(n14809), .B2(n12128), .A(n12127), .ZN(n12129) );
  AOI21_X1 U13952 ( .B1(n12130), .B2(n14811), .A(n12129), .ZN(n12131) );
  OAI211_X1 U13953 ( .C1(n12133), .C2(n14804), .A(n12132), .B(n12131), .ZN(
        P1_U3224) );
  INV_X1 U13954 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n15832) );
  AOI211_X1 U13955 ( .C1(n13099), .C2(n12136), .A(n12135), .B(n12134), .ZN(
        n12138) );
  MUX2_X1 U13956 ( .A(n15832), .B(n12138), .S(n16358), .Z(n12137) );
  OAI21_X1 U13957 ( .B1(n13223), .B2(n14631), .A(n12137), .ZN(P2_U3514) );
  INV_X1 U13958 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n12139) );
  MUX2_X1 U13959 ( .A(n12139), .B(n12138), .S(n14668), .Z(n12140) );
  OAI21_X1 U13960 ( .B1(n13223), .B2(n14673), .A(n12140), .ZN(P2_U3475) );
  NOR2_X1 U13961 ( .A1(n13226), .A2(n14507), .ZN(n12142) );
  XNOR2_X1 U13962 ( .A(n13227), .B(n8716), .ZN(n12141) );
  NOR2_X1 U13963 ( .A1(n12141), .A2(n12142), .ZN(n12234) );
  AOI21_X1 U13964 ( .B1(n12142), .B2(n12141), .A(n12234), .ZN(n12148) );
  INV_X1 U13965 ( .A(n12143), .ZN(n12145) );
  OAI21_X1 U13966 ( .B1(n12148), .B2(n12147), .A(n12236), .ZN(n12149) );
  NAND2_X1 U13967 ( .A1(n12149), .A2(n14232), .ZN(n12155) );
  NAND2_X1 U13968 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n12228)
         );
  INV_X1 U13969 ( .A(n12228), .ZN(n12153) );
  INV_X1 U13970 ( .A(n12150), .ZN(n12151) );
  OAI22_X1 U13971 ( .A1(n14219), .A2(n13222), .B1(n12151), .B2(n14218), .ZN(
        n12152) );
  AOI211_X1 U13972 ( .C1(n14225), .C2(n14324), .A(n12153), .B(n12152), .ZN(
        n12154) );
  OAI211_X1 U13973 ( .C1(n13227), .C2(n12244), .A(n12155), .B(n12154), .ZN(
        P2_U3198) );
  XNOR2_X1 U13974 ( .A(n12156), .B(n8025), .ZN(n12794) );
  XNOR2_X1 U13975 ( .A(n12794), .B(n13959), .ZN(n12164) );
  INV_X1 U13976 ( .A(n12159), .ZN(n12160) );
  NAND2_X1 U13977 ( .A1(n12160), .A2(n13613), .ZN(n12161) );
  INV_X1 U13978 ( .A(n13557), .ZN(n12162) );
  AOI21_X1 U13979 ( .B1(n12164), .B2(n12163), .A(n12162), .ZN(n12172) );
  INV_X1 U13980 ( .A(n12165), .ZN(n12170) );
  NOR2_X1 U13981 ( .A1(n14031), .A2(n13595), .ZN(n12169) );
  NAND2_X1 U13982 ( .A1(n13602), .A2(n13942), .ZN(n12167) );
  INV_X1 U13983 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n12166) );
  OR2_X1 U13984 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12166), .ZN(n15927) );
  OAI211_X1 U13985 ( .C1(n8384), .C2(n13600), .A(n12167), .B(n15927), .ZN(
        n12168) );
  AOI211_X1 U13986 ( .C1(n12170), .C2(n13568), .A(n12169), .B(n12168), .ZN(
        n12171) );
  OAI21_X1 U13987 ( .B1(n12172), .B2(n13608), .A(n12171), .ZN(P3_U3164) );
  OR2_X1 U13988 ( .A1(n14827), .A2(n14846), .ZN(n12173) );
  NAND2_X1 U13989 ( .A1(n12175), .A2(n12491), .ZN(n12178) );
  AOI22_X1 U13990 ( .A1(n12399), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n12398), 
        .B2(n12176), .ZN(n12177) );
  INV_X1 U13991 ( .A(n14845), .ZN(n12265) );
  XNOR2_X1 U13992 ( .A(n14745), .B(n12265), .ZN(n12743) );
  XOR2_X1 U13993 ( .A(n12245), .B(n12743), .Z(n15202) );
  NAND2_X1 U13994 ( .A1(n12179), .A2(n12740), .ZN(n12181) );
  INV_X1 U13995 ( .A(n14846), .ZN(n12375) );
  OR2_X1 U13996 ( .A1(n14827), .A2(n12375), .ZN(n12180) );
  XNOR2_X1 U13997 ( .A(n12252), .B(n12743), .ZN(n15199) );
  AOI21_X1 U13998 ( .B1(n14745), .B2(n12182), .A(n8189), .ZN(n15198) );
  INV_X1 U13999 ( .A(n12183), .ZN(n12191) );
  AND2_X1 U14000 ( .A1(n12185), .A2(n12184), .ZN(n12186) );
  OR2_X1 U14001 ( .A1(n12186), .A2(n12258), .ZN(n14764) );
  AOI22_X1 U14002 ( .A1(n12524), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n7427), 
        .B2(P1_REG2_REG_17__SCAN_IN), .ZN(n12188) );
  NAND2_X1 U14003 ( .A1(n12686), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n12187) );
  OAI211_X1 U14004 ( .C1(n14764), .C2(n12334), .A(n12188), .B(n12187), .ZN(
        n14844) );
  AND2_X1 U14005 ( .A1(n14846), .A2(n14806), .ZN(n12189) );
  AOI21_X1 U14006 ( .B1(n14844), .B2(n14807), .A(n12189), .ZN(n15195) );
  OAI21_X1 U14007 ( .B1(n14750), .B2(n16161), .A(n15195), .ZN(n12190) );
  AOI21_X1 U14008 ( .B1(n15198), .B2(n12191), .A(n12190), .ZN(n12193) );
  AOI22_X1 U14009 ( .A1(n14745), .A2(n16337), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(n16347), .ZN(n12192) );
  OAI21_X1 U14010 ( .B1(n12193), .B2(n16347), .A(n12192), .ZN(n12194) );
  AOI21_X1 U14011 ( .B1(n15199), .B2(n15090), .A(n12194), .ZN(n12195) );
  OAI21_X1 U14012 ( .B1(n15202), .B2(n15054), .A(n12195), .ZN(P1_U3277) );
  INV_X1 U14013 ( .A(n12196), .ZN(n12198) );
  NAND2_X1 U14014 ( .A1(n12198), .A2(n12197), .ZN(n12199) );
  NAND2_X1 U14015 ( .A1(n12616), .A2(n12494), .ZN(n12202) );
  NAND2_X1 U14016 ( .A1(n12202), .A2(n12201), .ZN(n12204) );
  XNOR2_X1 U14017 ( .A(n12204), .B(n12203), .ZN(n12357) );
  NOR2_X1 U14018 ( .A1(n12483), .A2(n12205), .ZN(n12206) );
  AOI21_X1 U14019 ( .B1(n12616), .B2(n8541), .A(n12206), .ZN(n12358) );
  XNOR2_X1 U14020 ( .A(n12357), .B(n12358), .ZN(n12208) );
  AOI21_X1 U14021 ( .B1(n12207), .B2(n12208), .A(n14829), .ZN(n12209) );
  NAND2_X1 U14022 ( .A1(n12209), .A2(n12362), .ZN(n12214) );
  OAI21_X1 U14023 ( .B1(n14809), .B2(n16376), .A(n12210), .ZN(n12211) );
  AOI21_X1 U14024 ( .B1(n12212), .B2(n14811), .A(n12211), .ZN(n12213) );
  OAI211_X1 U14025 ( .C1(n7671), .C2(n14804), .A(n12214), .B(n12213), .ZN(
        P1_U3234) );
  NOR2_X1 U14026 ( .A1(n12216), .A2(n15836), .ZN(n12217) );
  XNOR2_X1 U14027 ( .A(n14273), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n12218) );
  NOR2_X1 U14028 ( .A1(n12219), .A2(n12218), .ZN(n14269) );
  AOI211_X1 U14029 ( .C1(n12219), .C2(n12218), .A(n14269), .B(n15813), .ZN(
        n12231) );
  OAI21_X1 U14030 ( .B1(n12221), .B2(P2_REG2_REG_14__SCAN_IN), .A(n12220), 
        .ZN(n12222) );
  NOR2_X1 U14031 ( .A1(n15836), .A2(n12222), .ZN(n12223) );
  INV_X1 U14032 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n15827) );
  XNOR2_X1 U14033 ( .A(n15836), .B(n12222), .ZN(n15828) );
  NOR2_X1 U14034 ( .A1(n15827), .A2(n15828), .ZN(n15826) );
  NAND2_X1 U14035 ( .A1(n14273), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n12224) );
  OAI21_X1 U14036 ( .B1(n14273), .B2(P2_REG2_REG_16__SCAN_IN), .A(n12224), 
        .ZN(n12225) );
  NOR2_X1 U14037 ( .A1(n12226), .A2(n12225), .ZN(n14272) );
  AOI211_X1 U14038 ( .C1(n12226), .C2(n12225), .A(n14272), .B(n15817), .ZN(
        n12230) );
  INV_X1 U14039 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15772) );
  NAND2_X1 U14040 ( .A1(n15838), .A2(n14273), .ZN(n12227) );
  OAI211_X1 U14041 ( .C1(n15844), .C2(n15772), .A(n12228), .B(n12227), .ZN(
        n12229) );
  OR3_X1 U14042 ( .A1(n12231), .A2(n12230), .A3(n12229), .ZN(P2_U3230) );
  AND2_X1 U14043 ( .A1(n14324), .A2(n7431), .ZN(n12233) );
  XNOR2_X1 U14044 ( .A(n14336), .B(n11516), .ZN(n12232) );
  NOR2_X1 U14045 ( .A1(n12232), .A2(n12233), .ZN(n12272) );
  AOI21_X1 U14046 ( .B1(n12233), .B2(n12232), .A(n12272), .ZN(n12238) );
  INV_X1 U14047 ( .A(n12234), .ZN(n12235) );
  OAI21_X1 U14048 ( .B1(n12238), .B2(n12237), .A(n12274), .ZN(n12239) );
  NAND2_X1 U14049 ( .A1(n12239), .A2(n14232), .ZN(n12243) );
  INV_X1 U14050 ( .A(n14326), .ZN(n14340) );
  AND2_X1 U14051 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3088), .ZN(n14278) );
  OAI22_X1 U14052 ( .A1(n14219), .A2(n13226), .B1(n12240), .B2(n14218), .ZN(
        n12241) );
  AOI211_X1 U14053 ( .C1(n14225), .C2(n14340), .A(n14278), .B(n12241), .ZN(
        n12242) );
  OAI211_X1 U14054 ( .C1(n14674), .C2(n12244), .A(n12243), .B(n12242), .ZN(
        P2_U3200) );
  OR2_X1 U14055 ( .A1(n14745), .A2(n14845), .ZN(n12246) );
  NAND2_X1 U14056 ( .A1(n12248), .A2(n12491), .ZN(n12251) );
  AOI22_X1 U14057 ( .A1(n12399), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n12398), 
        .B2(n12249), .ZN(n12250) );
  INV_X1 U14058 ( .A(n14844), .ZN(n13058) );
  XNOR2_X1 U14059 ( .A(n15190), .B(n13058), .ZN(n12744) );
  INV_X1 U14060 ( .A(n12744), .ZN(n12254) );
  OAI21_X1 U14061 ( .B1(n7589), .B2(n12744), .A(n13045), .ZN(n15194) );
  NAND2_X1 U14062 ( .A1(n14745), .A2(n12265), .ZN(n12253) );
  OAI21_X1 U14063 ( .B1(n12255), .B2(n12254), .A(n13060), .ZN(n15191) );
  INV_X1 U14064 ( .A(n15081), .ZN(n12256) );
  AOI211_X1 U14065 ( .C1(n15190), .C2(n12257), .A(n16142), .B(n12256), .ZN(
        n15188) );
  NAND2_X1 U14066 ( .A1(n15188), .A2(n16341), .ZN(n12269) );
  NOR2_X1 U14067 ( .A1(n12258), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n12259) );
  OR2_X1 U14068 ( .A1(n12402), .A2(n12259), .ZN(n14798) );
  INV_X1 U14069 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n12262) );
  NAND2_X1 U14070 ( .A1(n12524), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n12261) );
  NAND2_X1 U14071 ( .A1(n12686), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n12260) );
  OAI211_X1 U14072 ( .C1(n12431), .C2(n12262), .A(n12261), .B(n12260), .ZN(
        n12263) );
  INV_X1 U14073 ( .A(n12263), .ZN(n12264) );
  OAI21_X1 U14074 ( .B1(n14798), .B2(n12334), .A(n12264), .ZN(n14843) );
  INV_X1 U14075 ( .A(n14843), .ZN(n13061) );
  OAI22_X1 U14076 ( .A1(n13061), .A2(n14787), .B1(n12265), .B2(n14785), .ZN(
        n15189) );
  INV_X1 U14077 ( .A(n15189), .ZN(n12266) );
  OAI22_X1 U14078 ( .A1(n16347), .A2(n12266), .B1(n14764), .B2(n16161), .ZN(
        n12267) );
  AOI21_X1 U14079 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n16347), .A(n12267), 
        .ZN(n12268) );
  OAI211_X1 U14080 ( .C1(n8188), .C2(n16163), .A(n12269), .B(n12268), .ZN(
        n12270) );
  AOI21_X1 U14081 ( .B1(n15090), .B2(n15191), .A(n12270), .ZN(n12271) );
  OAI21_X1 U14082 ( .B1(n15194), .B2(n15054), .A(n12271), .ZN(P1_U3276) );
  INV_X1 U14083 ( .A(n12272), .ZN(n12273) );
  NAND2_X1 U14084 ( .A1(n12350), .A2(n9720), .ZN(n12276) );
  AOI22_X1 U14085 ( .A1(n9659), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n13109), 
        .B2(n14286), .ZN(n12275) );
  XNOR2_X1 U14086 ( .A(n14619), .B(n8716), .ZN(n14122) );
  NOR2_X1 U14087 ( .A1(n14326), .A2(n14507), .ZN(n14123) );
  XNOR2_X1 U14088 ( .A(n14122), .B(n14123), .ZN(n14124) );
  XNOR2_X1 U14089 ( .A(n14125), .B(n14124), .ZN(n12291) );
  INV_X1 U14090 ( .A(n12279), .ZN(n12277) );
  AOI21_X1 U14091 ( .B1(n12277), .B2(P2_REG3_REG_18__SCAN_IN), .A(
        P2_REG3_REG_19__SCAN_IN), .ZN(n12280) );
  NAND2_X1 U14092 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n12278) );
  OR2_X1 U14093 ( .A1(n12280), .A2(n13100), .ZN(n14509) );
  INV_X1 U14094 ( .A(n14509), .ZN(n12281) );
  NAND2_X1 U14095 ( .A1(n12281), .A2(n11931), .ZN(n12287) );
  INV_X1 U14096 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n12284) );
  NAND2_X1 U14097 ( .A1(n9742), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n12283) );
  NAND2_X1 U14098 ( .A1(n13386), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n12282) );
  OAI211_X1 U14099 ( .C1(n12284), .C2(n9829), .A(n12283), .B(n12282), .ZN(
        n12285) );
  INV_X1 U14100 ( .A(n12285), .ZN(n12286) );
  AOI22_X1 U14101 ( .A1(n14227), .A2(n14324), .B1(n14540), .B2(n14242), .ZN(
        n12288) );
  NAND2_X1 U14102 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3088), .ZN(n14283)
         );
  OAI211_X1 U14103 ( .C1(n14524), .C2(n14217), .A(n12288), .B(n14283), .ZN(
        n12289) );
  AOI21_X1 U14104 ( .B1(n14536), .B2(n14246), .A(n12289), .ZN(n12290) );
  OAI21_X1 U14105 ( .B1(n12291), .B2(n14248), .A(n12290), .ZN(P2_U3210) );
  MUX2_X1 U14106 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n8006), .Z(n12294) );
  XNOR2_X1 U14107 ( .A(n12294), .B(SI_25_), .ZN(n12456) );
  INV_X1 U14108 ( .A(n12294), .ZN(n12295) );
  NAND2_X1 U14109 ( .A1(n12295), .A2(n15461), .ZN(n12296) );
  MUX2_X1 U14110 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n12298), .Z(n12299) );
  NAND2_X1 U14111 ( .A1(n12299), .A2(SI_26_), .ZN(n12300) );
  OAI21_X1 U14112 ( .B1(SI_26_), .B2(n12299), .A(n12300), .ZN(n12471) );
  MUX2_X1 U14113 ( .A(n15252), .B(n13333), .S(n8006), .Z(n12309) );
  NOR2_X1 U14114 ( .A1(n12309), .A2(n15460), .ZN(n12301) );
  NAND2_X1 U14115 ( .A1(n12309), .A2(n15460), .ZN(n12302) );
  MUX2_X1 U14116 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n8006), .Z(n12304) );
  XNOR2_X1 U14117 ( .A(n12304), .B(n12305), .ZN(n12506) );
  INV_X1 U14118 ( .A(n12304), .ZN(n12306) );
  NAND2_X1 U14119 ( .A1(n12306), .A2(n12305), .ZN(n12307) );
  MUX2_X1 U14120 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n8006), .Z(n12693) );
  INV_X1 U14121 ( .A(SI_29_), .ZN(n15456) );
  XNOR2_X1 U14122 ( .A(n12693), .B(n15456), .ZN(n12691) );
  INV_X1 U14123 ( .A(n13363), .ZN(n12847) );
  OAI222_X1 U14124 ( .A1(n15262), .A2(n12537), .B1(P1_U3086), .B2(n12308), 
        .C1(n15260), .C2(n12847), .ZN(P1_U3326) );
  INV_X1 U14125 ( .A(n12309), .ZN(n12310) );
  XNOR2_X1 U14126 ( .A(n12310), .B(SI_27_), .ZN(n12311) );
  INV_X1 U14127 ( .A(n15249), .ZN(n12313) );
  OAI222_X1 U14128 ( .A1(n14693), .A2(n13333), .B1(n14691), .B2(n12313), .C1(
        P2_U3088), .C2(n14314), .ZN(P2_U3300) );
  OR2_X1 U14129 ( .A1(n12314), .A2(n8006), .ZN(n12315) );
  XNOR2_X1 U14130 ( .A(n12315), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15264) );
  INV_X1 U14131 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14779) );
  INV_X1 U14132 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14733) );
  NOR2_X1 U14133 ( .A1(n12328), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n12317) );
  OR2_X1 U14134 ( .A1(n12427), .A2(n12317), .ZN(n15017) );
  INV_X1 U14135 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n15018) );
  NAND2_X1 U14136 ( .A1(n10089), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n12319) );
  NAND2_X1 U14137 ( .A1(n12686), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n12318) );
  OAI211_X1 U14138 ( .C1(n12431), .C2(n15018), .A(n12319), .B(n12318), .ZN(
        n12320) );
  INV_X1 U14139 ( .A(n12320), .ZN(n12321) );
  OAI21_X1 U14140 ( .B1(n15017), .B2(n12334), .A(n12321), .ZN(n14839) );
  INV_X1 U14141 ( .A(n14839), .ZN(n14715) );
  OAI22_X1 U14142 ( .A1(n15021), .A2(n10228), .B1(n14715), .B2(n12483), .ZN(
        n12420) );
  INV_X1 U14143 ( .A(n12420), .ZN(n12423) );
  NAND2_X1 U14144 ( .A1(n15155), .A2(n12494), .ZN(n12323) );
  NAND2_X1 U14145 ( .A1(n14839), .A2(n8541), .ZN(n12322) );
  NAND2_X1 U14146 ( .A1(n12323), .A2(n12322), .ZN(n12324) );
  XNOR2_X1 U14147 ( .A(n12324), .B(n12518), .ZN(n12421) );
  INV_X1 U14148 ( .A(n12421), .ZN(n12422) );
  OR2_X1 U14149 ( .A1(n13248), .A2(n8724), .ZN(n12327) );
  OR2_X1 U14150 ( .A1(n7433), .A2(n12325), .ZN(n12326) );
  AND2_X1 U14151 ( .A1(n12340), .A2(n14733), .ZN(n12329) );
  OR2_X1 U14152 ( .A1(n12329), .A2(n12328), .ZN(n15031) );
  INV_X1 U14153 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n15035) );
  NAND2_X1 U14154 ( .A1(n10089), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n12331) );
  NAND2_X1 U14155 ( .A1(n12686), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n12330) );
  OAI211_X1 U14156 ( .C1(n12431), .C2(n15035), .A(n12331), .B(n12330), .ZN(
        n12332) );
  INV_X1 U14157 ( .A(n12332), .ZN(n12333) );
  OAI21_X1 U14158 ( .B1(n15031), .B2(n12334), .A(n12333), .ZN(n14840) );
  AOI22_X1 U14159 ( .A1(n15159), .A2(n8541), .B1(n12520), .B2(n14840), .ZN(
        n12419) );
  AOI22_X1 U14160 ( .A1(n15159), .A2(n12494), .B1(n8541), .B2(n14840), .ZN(
        n12335) );
  XNOR2_X1 U14161 ( .A(n12335), .B(n12518), .ZN(n12418) );
  NAND2_X1 U14162 ( .A1(n13095), .A2(n12491), .ZN(n12338) );
  OR2_X1 U14163 ( .A1(n7432), .A2(n12336), .ZN(n12337) );
  NAND2_X1 U14164 ( .A1(n12404), .A2(n14779), .ZN(n12339) );
  AND2_X1 U14165 ( .A1(n12340), .A2(n12339), .ZN(n15044) );
  NAND2_X1 U14166 ( .A1(n15044), .A2(n12526), .ZN(n12345) );
  INV_X1 U14167 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n15047) );
  NAND2_X1 U14168 ( .A1(n10089), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n12342) );
  NAND2_X1 U14169 ( .A1(n12686), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n12341) );
  OAI211_X1 U14170 ( .C1(n15047), .C2(n12431), .A(n12342), .B(n12341), .ZN(
        n12343) );
  INV_X1 U14171 ( .A(n12343), .ZN(n12344) );
  NAND2_X1 U14172 ( .A1(n12345), .A2(n12344), .ZN(n14841) );
  AND2_X1 U14173 ( .A1(n14841), .A2(n12520), .ZN(n12346) );
  AOI21_X1 U14174 ( .B1(n15049), .B2(n8541), .A(n12346), .ZN(n12417) );
  NAND2_X1 U14175 ( .A1(n15049), .A2(n12494), .ZN(n12348) );
  NAND2_X1 U14176 ( .A1(n14841), .A2(n8541), .ZN(n12347) );
  NAND2_X1 U14177 ( .A1(n12348), .A2(n12347), .ZN(n12349) );
  XNOR2_X1 U14178 ( .A(n12349), .B(n12518), .ZN(n12416) );
  NAND2_X1 U14179 ( .A1(n12350), .A2(n12491), .ZN(n12353) );
  AOI22_X1 U14180 ( .A1(n12351), .A2(n12398), .B1(n12399), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n12352) );
  AOI22_X1 U14181 ( .A1(n15184), .A2(n8541), .B1(n12520), .B2(n14843), .ZN(
        n12395) );
  INV_X1 U14182 ( .A(n12395), .ZN(n12397) );
  NAND2_X1 U14183 ( .A1(n15184), .A2(n12494), .ZN(n12355) );
  NAND2_X1 U14184 ( .A1(n14843), .A2(n8541), .ZN(n12354) );
  NAND2_X1 U14185 ( .A1(n12355), .A2(n12354), .ZN(n12356) );
  XNOR2_X1 U14186 ( .A(n12356), .B(n12518), .ZN(n12396) );
  INV_X1 U14187 ( .A(n12357), .ZN(n12360) );
  INV_X1 U14188 ( .A(n12358), .ZN(n12359) );
  NAND2_X1 U14189 ( .A1(n12360), .A2(n12359), .ZN(n12361) );
  NAND2_X1 U14190 ( .A1(n14705), .A2(n12494), .ZN(n12364) );
  NAND2_X1 U14191 ( .A1(n12364), .A2(n12363), .ZN(n12365) );
  XNOR2_X1 U14192 ( .A(n12365), .B(n12518), .ZN(n12368) );
  NOR2_X1 U14193 ( .A1(n12483), .A2(n12366), .ZN(n12367) );
  AOI21_X1 U14194 ( .B1(n14705), .B2(n8541), .A(n12367), .ZN(n12369) );
  XNOR2_X1 U14195 ( .A(n12368), .B(n12369), .ZN(n14707) );
  INV_X1 U14196 ( .A(n12368), .ZN(n12370) );
  NAND2_X1 U14197 ( .A1(n12370), .A2(n12369), .ZN(n12371) );
  NAND2_X1 U14198 ( .A1(n14827), .A2(n12494), .ZN(n12373) );
  NAND2_X1 U14199 ( .A1(n12373), .A2(n12372), .ZN(n12374) );
  XNOR2_X1 U14200 ( .A(n12374), .B(n12518), .ZN(n12377) );
  NOR2_X1 U14201 ( .A1(n12483), .A2(n12375), .ZN(n12376) );
  AOI21_X1 U14202 ( .B1(n14827), .B2(n8541), .A(n12376), .ZN(n14816) );
  INV_X1 U14203 ( .A(n12377), .ZN(n12378) );
  NAND2_X1 U14204 ( .A1(n14745), .A2(n12494), .ZN(n12380) );
  NAND2_X1 U14205 ( .A1(n12380), .A2(n12379), .ZN(n12381) );
  XNOR2_X1 U14206 ( .A(n12381), .B(n12518), .ZN(n12384) );
  AOI22_X1 U14207 ( .A1(n14745), .A2(n8541), .B1(n12520), .B2(n14845), .ZN(
        n12382) );
  XNOR2_X1 U14208 ( .A(n12384), .B(n12382), .ZN(n14748) );
  INV_X1 U14209 ( .A(n12382), .ZN(n12383) );
  NAND2_X1 U14210 ( .A1(n15190), .A2(n12494), .ZN(n12387) );
  NAND2_X1 U14211 ( .A1(n14844), .A2(n8541), .ZN(n12386) );
  NAND2_X1 U14212 ( .A1(n12387), .A2(n12386), .ZN(n12388) );
  XNOR2_X1 U14213 ( .A(n12388), .B(n12518), .ZN(n12391) );
  NAND2_X1 U14214 ( .A1(n15190), .A2(n8541), .ZN(n12390) );
  NAND2_X1 U14215 ( .A1(n12520), .A2(n14844), .ZN(n12389) );
  NAND2_X1 U14216 ( .A1(n12390), .A2(n12389), .ZN(n12392) );
  NAND2_X1 U14217 ( .A1(n12391), .A2(n12392), .ZN(n14758) );
  INV_X1 U14218 ( .A(n12391), .ZN(n12394) );
  INV_X1 U14219 ( .A(n12392), .ZN(n12393) );
  NAND2_X1 U14220 ( .A1(n12394), .A2(n12393), .ZN(n14760) );
  XNOR2_X1 U14221 ( .A(n12396), .B(n12395), .ZN(n14795) );
  NAND2_X1 U14222 ( .A1(n13108), .A2(n12491), .ZN(n12401) );
  AOI22_X1 U14223 ( .A1(n12399), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n12398), 
        .B2(n16038), .ZN(n12400) );
  NAND2_X1 U14224 ( .A1(n15174), .A2(n12494), .ZN(n12411) );
  OR2_X1 U14225 ( .A1(n12402), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n12403) );
  AND2_X1 U14226 ( .A1(n12404), .A2(n12403), .ZN(n15062) );
  NAND2_X1 U14227 ( .A1(n15062), .A2(n12526), .ZN(n12409) );
  INV_X1 U14228 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n15066) );
  NAND2_X1 U14229 ( .A1(n12524), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n12406) );
  NAND2_X1 U14230 ( .A1(n12686), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n12405) );
  OAI211_X1 U14231 ( .C1(n12431), .C2(n15066), .A(n12406), .B(n12405), .ZN(
        n12407) );
  INV_X1 U14232 ( .A(n12407), .ZN(n12408) );
  NAND2_X1 U14233 ( .A1(n12409), .A2(n12408), .ZN(n14842) );
  NAND2_X1 U14234 ( .A1(n14842), .A2(n8541), .ZN(n12410) );
  NAND2_X1 U14235 ( .A1(n12411), .A2(n12410), .ZN(n12412) );
  XNOR2_X1 U14236 ( .A(n12412), .B(n12518), .ZN(n12413) );
  AOI22_X1 U14237 ( .A1(n15174), .A2(n8541), .B1(n12520), .B2(n14842), .ZN(
        n12414) );
  XNOR2_X1 U14238 ( .A(n12413), .B(n12414), .ZN(n14722) );
  INV_X1 U14239 ( .A(n12413), .ZN(n12415) );
  XNOR2_X1 U14240 ( .A(n12416), .B(n12417), .ZN(n14777) );
  XNOR2_X1 U14241 ( .A(n12418), .B(n12419), .ZN(n14731) );
  XNOR2_X1 U14242 ( .A(n12421), .B(n12420), .ZN(n14784) );
  NAND2_X1 U14243 ( .A1(n13278), .A2(n12491), .ZN(n12426) );
  OR2_X1 U14244 ( .A1(n7432), .A2(n12424), .ZN(n12425) );
  OR2_X1 U14245 ( .A1(n12427), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n12428) );
  NAND2_X1 U14246 ( .A1(n12427), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n12444) );
  AND2_X1 U14247 ( .A1(n12428), .A2(n12444), .ZN(n15001) );
  NAND2_X1 U14248 ( .A1(n15001), .A2(n12526), .ZN(n12434) );
  INV_X1 U14249 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n15004) );
  NAND2_X1 U14250 ( .A1(n12524), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n12430) );
  NAND2_X1 U14251 ( .A1(n12686), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n12429) );
  OAI211_X1 U14252 ( .C1(n12431), .C2(n15004), .A(n12430), .B(n12429), .ZN(
        n12432) );
  INV_X1 U14253 ( .A(n12432), .ZN(n12433) );
  NAND2_X1 U14254 ( .A1(n12434), .A2(n12433), .ZN(n14838) );
  AOI22_X1 U14255 ( .A1(n15147), .A2(n8541), .B1(n12520), .B2(n14838), .ZN(
        n12438) );
  NAND2_X1 U14256 ( .A1(n15147), .A2(n12494), .ZN(n12436) );
  NAND2_X1 U14257 ( .A1(n14838), .A2(n8541), .ZN(n12435) );
  NAND2_X1 U14258 ( .A1(n12436), .A2(n12435), .ZN(n12437) );
  XNOR2_X1 U14259 ( .A(n12437), .B(n12518), .ZN(n12440) );
  XOR2_X1 U14260 ( .A(n12438), .B(n12440), .Z(n14713) );
  INV_X1 U14261 ( .A(n12438), .ZN(n12439) );
  OR2_X1 U14262 ( .A1(n13293), .A2(n8724), .ZN(n12442) );
  OR2_X1 U14263 ( .A1(n7433), .A2(n7719), .ZN(n12441) );
  NAND2_X1 U14264 ( .A1(n7426), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n12448) );
  NAND2_X1 U14265 ( .A1(n12524), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n12447) );
  INV_X1 U14266 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14771) );
  INV_X1 U14267 ( .A(n12444), .ZN(n12443) );
  NAND2_X1 U14268 ( .A1(n12443), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n12461) );
  AOI21_X1 U14269 ( .B1(n14771), .B2(n12444), .A(n12460), .ZN(n14993) );
  NAND2_X1 U14270 ( .A1(n12526), .A2(n14993), .ZN(n12446) );
  NAND2_X1 U14271 ( .A1(n12686), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n12445) );
  NAND4_X1 U14272 ( .A1(n12448), .A2(n12447), .A3(n12446), .A4(n12445), .ZN(
        n14837) );
  INV_X1 U14273 ( .A(n14837), .ZN(n14714) );
  OAI22_X1 U14274 ( .A1(n14992), .A2(n10228), .B1(n14714), .B2(n12483), .ZN(
        n12453) );
  NAND2_X1 U14275 ( .A1(n15138), .A2(n12494), .ZN(n12450) );
  NAND2_X1 U14276 ( .A1(n12450), .A2(n12449), .ZN(n12451) );
  XNOR2_X1 U14277 ( .A(n12451), .B(n12518), .ZN(n12452) );
  XOR2_X1 U14278 ( .A(n12453), .B(n12452), .Z(n14769) );
  INV_X1 U14279 ( .A(n12452), .ZN(n12455) );
  INV_X1 U14280 ( .A(n12453), .ZN(n12454) );
  XNOR2_X1 U14281 ( .A(n12457), .B(n12456), .ZN(n14689) );
  NAND2_X1 U14282 ( .A1(n14689), .A2(n12491), .ZN(n12459) );
  OR2_X1 U14283 ( .A1(n7432), .A2(n15261), .ZN(n12458) );
  NAND2_X1 U14284 ( .A1(n14972), .A2(n12494), .ZN(n12467) );
  NAND2_X1 U14285 ( .A1(n7427), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n12465) );
  NAND2_X1 U14286 ( .A1(n12524), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n12464) );
  INV_X1 U14287 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14740) );
  NAND2_X1 U14288 ( .A1(n12460), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n12478) );
  INV_X1 U14289 ( .A(n12478), .ZN(n12477) );
  AOI21_X1 U14290 ( .B1(n14740), .B2(n12461), .A(n12477), .ZN(n14973) );
  NAND2_X1 U14291 ( .A1(n12526), .A2(n14973), .ZN(n12463) );
  NAND2_X1 U14292 ( .A1(n12686), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n12462) );
  NAND4_X1 U14293 ( .A1(n12465), .A2(n12464), .A3(n12463), .A4(n12462), .ZN(
        n14836) );
  NAND2_X1 U14294 ( .A1(n12467), .A2(n12466), .ZN(n12468) );
  XNOR2_X1 U14295 ( .A(n12468), .B(n12518), .ZN(n12470) );
  INV_X1 U14296 ( .A(n14836), .ZN(n13054) );
  OAI22_X1 U14297 ( .A1(n15132), .A2(n10228), .B1(n13054), .B2(n12483), .ZN(
        n12469) );
  XNOR2_X1 U14298 ( .A(n12470), .B(n12469), .ZN(n14739) );
  NAND2_X1 U14299 ( .A1(n12472), .A2(n12471), .ZN(n12473) );
  NAND2_X1 U14300 ( .A1(n12474), .A2(n12473), .ZN(n15255) );
  OR2_X1 U14301 ( .A1(n7433), .A2(n15254), .ZN(n12475) );
  NAND2_X1 U14302 ( .A1(n7427), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n12482) );
  NAND2_X1 U14303 ( .A1(n12524), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n12481) );
  INV_X1 U14304 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14808) );
  NAND2_X1 U14305 ( .A1(n12477), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n12495) );
  INV_X1 U14306 ( .A(n12495), .ZN(n12510) );
  AOI21_X1 U14307 ( .B1(n14808), .B2(n12478), .A(n12510), .ZN(n14959) );
  NAND2_X1 U14308 ( .A1(n12526), .A2(n14959), .ZN(n12480) );
  NAND2_X1 U14309 ( .A1(n12686), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n12479) );
  NAND4_X1 U14310 ( .A1(n12482), .A2(n12481), .A3(n12480), .A4(n12479), .ZN(
        n14835) );
  OAI22_X1 U14311 ( .A1(n15126), .A2(n10228), .B1(n14698), .B2(n12483), .ZN(
        n12488) );
  NAND2_X1 U14312 ( .A1(n14812), .A2(n12494), .ZN(n12485) );
  NAND2_X1 U14313 ( .A1(n12485), .A2(n12484), .ZN(n12486) );
  XNOR2_X1 U14314 ( .A(n12486), .B(n12518), .ZN(n12487) );
  INV_X1 U14315 ( .A(n12487), .ZN(n12490) );
  INV_X1 U14316 ( .A(n12488), .ZN(n12489) );
  NAND2_X1 U14317 ( .A1(n15249), .A2(n12491), .ZN(n12493) );
  OR2_X1 U14318 ( .A1(n7433), .A2(n15252), .ZN(n12492) );
  NAND2_X1 U14319 ( .A1(n15119), .A2(n12494), .ZN(n12501) );
  NAND2_X1 U14320 ( .A1(n10089), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n12499) );
  NAND2_X1 U14321 ( .A1(n12686), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n12498) );
  XNOR2_X1 U14322 ( .A(P1_REG3_REG_27__SCAN_IN), .B(n12495), .ZN(n14944) );
  NAND2_X1 U14323 ( .A1(n12526), .A2(n14944), .ZN(n12497) );
  NAND2_X1 U14324 ( .A1(n7426), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n12496) );
  NAND4_X1 U14325 ( .A1(n12499), .A2(n12498), .A3(n12497), .A4(n12496), .ZN(
        n14834) );
  NAND2_X1 U14326 ( .A1(n8541), .A2(n14834), .ZN(n12500) );
  NAND2_X1 U14327 ( .A1(n12501), .A2(n12500), .ZN(n12502) );
  XNOR2_X1 U14328 ( .A(n12502), .B(n12518), .ZN(n12504) );
  INV_X1 U14329 ( .A(n15119), .ZN(n14947) );
  INV_X1 U14330 ( .A(n14834), .ZN(n13071) );
  OAI22_X1 U14331 ( .A1(n14947), .A2(n10228), .B1(n13071), .B2(n12483), .ZN(
        n12503) );
  XNOR2_X1 U14332 ( .A(n12504), .B(n12503), .ZN(n14697) );
  NAND2_X1 U14333 ( .A1(n14683), .A2(n12491), .ZN(n12509) );
  OR2_X1 U14334 ( .A1(n7432), .A2(n15247), .ZN(n12508) );
  NAND2_X1 U14335 ( .A1(n7426), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n12517) );
  NAND2_X1 U14336 ( .A1(n12524), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n12516) );
  NAND2_X1 U14337 ( .A1(n12511), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n12525) );
  INV_X1 U14338 ( .A(n12511), .ZN(n12512) );
  INV_X1 U14339 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n12532) );
  NAND2_X1 U14340 ( .A1(n12512), .A2(n12532), .ZN(n12513) );
  NAND2_X1 U14341 ( .A1(n12526), .A2(n14927), .ZN(n12515) );
  NAND2_X1 U14342 ( .A1(n12686), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n12514) );
  NAND4_X1 U14343 ( .A1(n12517), .A2(n12516), .A3(n12515), .A4(n12514), .ZN(
        n14833) );
  AOI22_X1 U14344 ( .A1(n15115), .A2(n12494), .B1(n8541), .B2(n14833), .ZN(
        n12519) );
  XNOR2_X1 U14345 ( .A(n12519), .B(n12518), .ZN(n12522) );
  AOI22_X1 U14346 ( .A1(n15115), .A2(n8541), .B1(n12520), .B2(n14833), .ZN(
        n12521) );
  XNOR2_X1 U14347 ( .A(n12522), .B(n12521), .ZN(n12523) );
  NAND2_X1 U14348 ( .A1(n12524), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n12530) );
  NAND2_X1 U14349 ( .A1(n12686), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n12529) );
  INV_X1 U14350 ( .A(n12525), .ZN(n13083) );
  NAND2_X1 U14351 ( .A1(n12526), .A2(n13083), .ZN(n12528) );
  NAND2_X1 U14352 ( .A1(n7427), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n12527) );
  INV_X1 U14353 ( .A(n12541), .ZN(n14832) );
  AND2_X1 U14354 ( .A1(n14834), .A2(n14806), .ZN(n12531) );
  AOI21_X1 U14355 ( .B1(n14832), .B2(n14799), .A(n12531), .ZN(n14935) );
  OAI22_X1 U14356 ( .A1(n14809), .A2(n14935), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12532), .ZN(n12533) );
  AOI21_X1 U14357 ( .B1(n14927), .B2(n14811), .A(n12533), .ZN(n12535) );
  NAND2_X1 U14358 ( .A1(n15115), .A2(n14826), .ZN(n12534) );
  NAND2_X1 U14359 ( .A1(n13363), .A2(n12491), .ZN(n12539) );
  OR2_X1 U14360 ( .A1(n7432), .A2(n12537), .ZN(n12538) );
  XNOR2_X1 U14361 ( .A(n15263), .B(n12752), .ZN(n12703) );
  MUX2_X1 U14362 ( .A(n16039), .B(n12540), .S(n12703), .Z(n12543) );
  MUX2_X1 U14363 ( .A(n15108), .B(n12541), .S(n12551), .Z(n12684) );
  MUX2_X1 U14364 ( .A(n14851), .B(n12601), .S(n12551), .Z(n12605) );
  AOI21_X1 U14365 ( .B1(n12542), .B2(n12682), .A(n16189), .ZN(n12568) );
  AOI21_X1 U14366 ( .B1(n14857), .B2(n12551), .A(n12544), .ZN(n12567) );
  NAND3_X1 U14367 ( .A1(n12546), .A2(n12556), .A3(n12555), .ZN(n12545) );
  INV_X1 U14368 ( .A(n12546), .ZN(n16072) );
  NAND2_X1 U14369 ( .A1(n16072), .A2(n12547), .ZN(n12548) );
  NAND2_X1 U14370 ( .A1(n14862), .A2(n16031), .ZN(n12724) );
  NAND3_X1 U14371 ( .A1(n12548), .A2(n12682), .A3(n12724), .ZN(n12549) );
  NAND3_X1 U14372 ( .A1(n12553), .A2(n12552), .A3(n12551), .ZN(n12559) );
  INV_X1 U14373 ( .A(n12556), .ZN(n12554) );
  NAND2_X1 U14374 ( .A1(n12554), .A2(n12551), .ZN(n12558) );
  NAND3_X1 U14375 ( .A1(n12556), .A2(n12555), .A3(n12682), .ZN(n12557) );
  MUX2_X1 U14376 ( .A(n12561), .B(n16162), .S(n12682), .Z(n12563) );
  MUX2_X1 U14377 ( .A(n14858), .B(n16143), .S(n12551), .Z(n12562) );
  NAND2_X1 U14378 ( .A1(n14856), .A2(n12682), .ZN(n12569) );
  NAND2_X1 U14379 ( .A1(n16208), .A2(n12569), .ZN(n12572) );
  OAI21_X1 U14380 ( .B1(n14856), .B2(n12682), .A(n12570), .ZN(n12571) );
  NAND2_X1 U14381 ( .A1(n12572), .A2(n12571), .ZN(n12573) );
  MUX2_X1 U14382 ( .A(n14855), .B(n12575), .S(n12551), .Z(n12578) );
  NAND2_X1 U14383 ( .A1(n12579), .A2(n12578), .ZN(n12577) );
  MUX2_X1 U14384 ( .A(n14855), .B(n12575), .S(n12705), .Z(n12576) );
  NAND2_X1 U14385 ( .A1(n12577), .A2(n12576), .ZN(n12580) );
  MUX2_X1 U14386 ( .A(n14854), .B(n16240), .S(n12705), .Z(n12582) );
  MUX2_X1 U14387 ( .A(n14854), .B(n16240), .S(n12551), .Z(n12581) );
  MUX2_X1 U14388 ( .A(n14853), .B(n12583), .S(n12551), .Z(n12587) );
  NAND2_X1 U14389 ( .A1(n12586), .A2(n12587), .ZN(n12585) );
  MUX2_X1 U14390 ( .A(n14853), .B(n12583), .S(n12705), .Z(n12584) );
  NAND2_X1 U14391 ( .A1(n12585), .A2(n12584), .ZN(n12591) );
  INV_X1 U14392 ( .A(n12586), .ZN(n12589) );
  INV_X1 U14393 ( .A(n12587), .ZN(n12588) );
  NAND2_X1 U14394 ( .A1(n12589), .A2(n12588), .ZN(n12590) );
  NAND2_X1 U14395 ( .A1(n12591), .A2(n12590), .ZN(n12595) );
  INV_X1 U14396 ( .A(n12551), .ZN(n12705) );
  MUX2_X1 U14397 ( .A(n14852), .B(n12592), .S(n12705), .Z(n12596) );
  NAND2_X1 U14398 ( .A1(n12595), .A2(n12596), .ZN(n12594) );
  MUX2_X1 U14399 ( .A(n14852), .B(n12592), .S(n12551), .Z(n12593) );
  NAND2_X1 U14400 ( .A1(n12594), .A2(n12593), .ZN(n12600) );
  INV_X1 U14401 ( .A(n12595), .ZN(n12598) );
  INV_X1 U14402 ( .A(n12596), .ZN(n12597) );
  NAND2_X1 U14403 ( .A1(n12598), .A2(n12597), .ZN(n12599) );
  NAND2_X1 U14404 ( .A1(n12604), .A2(n12605), .ZN(n12603) );
  MUX2_X1 U14405 ( .A(n14851), .B(n12601), .S(n12705), .Z(n12602) );
  MUX2_X1 U14406 ( .A(n12606), .B(n16324), .S(n12705), .Z(n12609) );
  NAND2_X1 U14407 ( .A1(n12609), .A2(n12608), .ZN(n12607) );
  INV_X1 U14408 ( .A(n12608), .ZN(n12611) );
  INV_X1 U14409 ( .A(n12609), .ZN(n12610) );
  NAND3_X1 U14410 ( .A1(n12736), .A2(n12611), .A3(n12610), .ZN(n12615) );
  AND2_X1 U14411 ( .A1(n14849), .A2(n12551), .ZN(n12613) );
  OAI21_X1 U14412 ( .B1(n12551), .B2(n14849), .A(n16365), .ZN(n12612) );
  OAI21_X1 U14413 ( .B1(n12613), .B2(n16365), .A(n12612), .ZN(n12614) );
  MUX2_X1 U14414 ( .A(n14848), .B(n12616), .S(n12705), .Z(n12619) );
  NAND2_X1 U14415 ( .A1(n12620), .A2(n12619), .ZN(n12618) );
  MUX2_X1 U14416 ( .A(n14848), .B(n12616), .S(n12551), .Z(n12617) );
  NAND2_X1 U14417 ( .A1(n12618), .A2(n12617), .ZN(n12621) );
  MUX2_X1 U14418 ( .A(n14847), .B(n14705), .S(n12551), .Z(n12623) );
  MUX2_X1 U14419 ( .A(n14847), .B(n14705), .S(n12705), .Z(n12622) );
  MUX2_X1 U14420 ( .A(n14846), .B(n14827), .S(n12705), .Z(n12626) );
  MUX2_X1 U14421 ( .A(n14846), .B(n14827), .S(n12551), .Z(n12624) );
  INV_X1 U14422 ( .A(n12626), .ZN(n12627) );
  MUX2_X1 U14423 ( .A(n14845), .B(n14745), .S(n12551), .Z(n12631) );
  MUX2_X1 U14424 ( .A(n14845), .B(n14745), .S(n12705), .Z(n12628) );
  MUX2_X1 U14425 ( .A(n14844), .B(n15190), .S(n12705), .Z(n12633) );
  MUX2_X1 U14426 ( .A(n14844), .B(n15190), .S(n12551), .Z(n12632) );
  MUX2_X1 U14427 ( .A(n14843), .B(n15184), .S(n12551), .Z(n12636) );
  MUX2_X1 U14428 ( .A(n14843), .B(n15184), .S(n12705), .Z(n12634) );
  MUX2_X1 U14429 ( .A(n14842), .B(n15174), .S(n12705), .Z(n12638) );
  MUX2_X1 U14430 ( .A(n14842), .B(n15174), .S(n12551), .Z(n12637) );
  INV_X1 U14431 ( .A(n12638), .ZN(n12639) );
  MUX2_X1 U14432 ( .A(n14841), .B(n15049), .S(n12551), .Z(n12643) );
  MUX2_X1 U14433 ( .A(n14841), .B(n15049), .S(n12705), .Z(n12640) );
  NAND2_X1 U14434 ( .A1(n12641), .A2(n12640), .ZN(n12647) );
  INV_X1 U14435 ( .A(n12642), .ZN(n12645) );
  INV_X1 U14436 ( .A(n12643), .ZN(n12644) );
  NAND2_X1 U14437 ( .A1(n12645), .A2(n12644), .ZN(n12646) );
  MUX2_X1 U14438 ( .A(n14840), .B(n15159), .S(n12705), .Z(n12650) );
  NAND2_X1 U14439 ( .A1(n12651), .A2(n12650), .ZN(n12649) );
  MUX2_X1 U14440 ( .A(n14840), .B(n15159), .S(n12551), .Z(n12648) );
  NAND2_X1 U14441 ( .A1(n12649), .A2(n12648), .ZN(n12652) );
  MUX2_X1 U14442 ( .A(n14839), .B(n15155), .S(n12551), .Z(n12654) );
  MUX2_X1 U14443 ( .A(n14839), .B(n15155), .S(n12705), .Z(n12653) );
  MUX2_X1 U14444 ( .A(n14838), .B(n15147), .S(n12682), .Z(n12656) );
  MUX2_X1 U14445 ( .A(n14838), .B(n15147), .S(n12551), .Z(n12655) );
  INV_X1 U14446 ( .A(n12656), .ZN(n12657) );
  MUX2_X1 U14447 ( .A(n15138), .B(n14837), .S(n12682), .Z(n12660) );
  MUX2_X1 U14448 ( .A(n14837), .B(n15138), .S(n12682), .Z(n12658) );
  MUX2_X1 U14449 ( .A(n14836), .B(n14972), .S(n12682), .Z(n12662) );
  MUX2_X1 U14450 ( .A(n14836), .B(n14972), .S(n12551), .Z(n12661) );
  MUX2_X1 U14451 ( .A(n14812), .B(n14835), .S(n12551), .Z(n12668) );
  INV_X1 U14452 ( .A(n12668), .ZN(n12663) );
  MUX2_X1 U14453 ( .A(n14812), .B(n14835), .S(n12682), .Z(n12664) );
  INV_X1 U14454 ( .A(n12664), .ZN(n12665) );
  NAND2_X1 U14455 ( .A1(n12666), .A2(n12665), .ZN(n12671) );
  INV_X1 U14456 ( .A(n12667), .ZN(n12669) );
  NAND2_X1 U14457 ( .A1(n12669), .A2(n12668), .ZN(n12670) );
  MUX2_X1 U14458 ( .A(n14834), .B(n15119), .S(n12682), .Z(n12673) );
  MUX2_X1 U14459 ( .A(n14834), .B(n15119), .S(n12551), .Z(n12672) );
  MUX2_X1 U14460 ( .A(n14833), .B(n15115), .S(n12551), .Z(n12677) );
  NAND2_X1 U14461 ( .A1(n12676), .A2(n12677), .ZN(n12675) );
  MUX2_X1 U14462 ( .A(n14833), .B(n15115), .S(n12682), .Z(n12674) );
  NAND2_X1 U14463 ( .A1(n12675), .A2(n12674), .ZN(n12681) );
  INV_X1 U14464 ( .A(n12676), .ZN(n12679) );
  INV_X1 U14465 ( .A(n12677), .ZN(n12678) );
  NAND2_X1 U14466 ( .A1(n12679), .A2(n12678), .ZN(n12680) );
  MUX2_X1 U14467 ( .A(n13076), .B(n14832), .S(n12682), .Z(n12683) );
  NAND2_X1 U14468 ( .A1(n10089), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n12689) );
  NAND2_X1 U14469 ( .A1(n7426), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n12688) );
  NAND2_X1 U14470 ( .A1(n12686), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n12687) );
  AND3_X1 U14471 ( .A1(n12689), .A2(n12688), .A3(n12687), .ZN(n12722) );
  INV_X1 U14472 ( .A(n12722), .ZN(n14831) );
  OAI21_X1 U14473 ( .B1(n14914), .B2(n16039), .A(n14831), .ZN(n12690) );
  INV_X1 U14474 ( .A(n12690), .ZN(n12702) );
  INV_X1 U14475 ( .A(n12693), .ZN(n12694) );
  NAND2_X1 U14476 ( .A1(n12694), .A2(n15456), .ZN(n12695) );
  MUX2_X1 U14477 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n8006), .Z(n12696) );
  NAND2_X1 U14478 ( .A1(n12696), .A2(SI_30_), .ZN(n12707) );
  OAI21_X1 U14479 ( .B1(n12696), .B2(SI_30_), .A(n12707), .ZN(n12697) );
  NAND2_X1 U14480 ( .A1(n12698), .A2(n12697), .ZN(n12699) );
  NAND2_X1 U14481 ( .A1(n14681), .A2(n12491), .ZN(n12701) );
  INV_X1 U14482 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n15244) );
  OR2_X1 U14483 ( .A1(n7432), .A2(n15244), .ZN(n12700) );
  MUX2_X1 U14484 ( .A(n12702), .B(n14911), .S(n12551), .Z(n12775) );
  INV_X1 U14485 ( .A(n12775), .ZN(n12720) );
  OAI21_X1 U14486 ( .B1(n14914), .B2(n12703), .A(n14831), .ZN(n12704) );
  INV_X1 U14487 ( .A(n12704), .ZN(n12706) );
  MUX2_X1 U14488 ( .A(n12706), .B(n14911), .S(n12705), .Z(n12779) );
  MUX2_X1 U14489 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8006), .Z(n12710) );
  XNOR2_X1 U14490 ( .A(n12710), .B(SI_31_), .ZN(n12711) );
  NAND2_X1 U14491 ( .A1(n15236), .A2(n12491), .ZN(n12714) );
  INV_X1 U14492 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n15241) );
  OR2_X1 U14493 ( .A1(n7433), .A2(n15241), .ZN(n12713) );
  XNOR2_X1 U14494 ( .A(n15101), .B(n14914), .ZN(n12772) );
  NAND2_X1 U14495 ( .A1(n12716), .A2(n12715), .ZN(n12717) );
  AND2_X1 U14496 ( .A1(n12718), .A2(n12717), .ZN(n12756) );
  NAND2_X1 U14497 ( .A1(n12772), .A2(n12756), .ZN(n12777) );
  INV_X1 U14498 ( .A(n12777), .ZN(n12719) );
  INV_X1 U14499 ( .A(n12774), .ZN(n12785) );
  OAI211_X1 U14500 ( .C1(n12720), .C2(n12779), .A(n12719), .B(n12785), .ZN(
        n12791) );
  NAND2_X1 U14501 ( .A1(n15101), .A2(n12551), .ZN(n12758) );
  OR2_X1 U14502 ( .A1(n15101), .A2(n12551), .ZN(n12762) );
  INV_X1 U14503 ( .A(n14914), .ZN(n12759) );
  NOR2_X1 U14504 ( .A1(n12762), .A2(n12759), .ZN(n12757) );
  INV_X1 U14505 ( .A(n12757), .ZN(n12721) );
  INV_X1 U14506 ( .A(n12756), .ZN(n12761) );
  INV_X1 U14507 ( .A(n12754), .ZN(n12765) );
  AND2_X1 U14508 ( .A1(n12761), .A2(n12765), .ZN(n12773) );
  OAI211_X1 U14509 ( .C1(n14914), .C2(n12758), .A(n12721), .B(n12773), .ZN(
        n12780) );
  NAND2_X1 U14510 ( .A1(n12775), .A2(n12785), .ZN(n12778) );
  NOR2_X1 U14511 ( .A1(n12780), .A2(n12778), .ZN(n12770) );
  XNOR2_X1 U14512 ( .A(n14911), .B(n12722), .ZN(n12750) );
  NAND2_X1 U14513 ( .A1(n15115), .A2(n14833), .ZN(n13055) );
  OR2_X1 U14514 ( .A1(n15115), .A2(n14833), .ZN(n12723) );
  NAND2_X1 U14515 ( .A1(n13055), .A2(n12723), .ZN(n14933) );
  XNOR2_X1 U14516 ( .A(n14812), .B(n14698), .ZN(n14955) );
  XNOR2_X1 U14517 ( .A(n15138), .B(n14837), .ZN(n14980) );
  XNOR2_X1 U14518 ( .A(n15021), .B(n14715), .ZN(n15011) );
  INV_X1 U14519 ( .A(n14840), .ZN(n14786) );
  XNOR2_X1 U14520 ( .A(n15159), .B(n14786), .ZN(n15028) );
  XNOR2_X1 U14521 ( .A(n15049), .B(n14841), .ZN(n13064) );
  AND2_X1 U14522 ( .A1(n16072), .A2(n12724), .ZN(n16044) );
  NAND4_X1 U14523 ( .A1(n16073), .A2(n16044), .A3(n12725), .A4(n16137), .ZN(
        n12727) );
  NOR3_X1 U14524 ( .A1(n12727), .A2(n8675), .A3(n12726), .ZN(n12730) );
  NAND4_X1 U14525 ( .A1(n12731), .A2(n12730), .A3(n12729), .A4(n12728), .ZN(
        n12732) );
  NOR2_X1 U14526 ( .A1(n12733), .A2(n12732), .ZN(n12735) );
  XNOR2_X1 U14527 ( .A(n16338), .B(n14850), .ZN(n16325) );
  NAND4_X1 U14528 ( .A1(n12736), .A2(n12735), .A3(n16325), .A4(n12734), .ZN(
        n12737) );
  NOR2_X1 U14529 ( .A1(n12738), .A2(n12737), .ZN(n12741) );
  NAND4_X1 U14530 ( .A1(n13064), .A2(n12741), .A3(n12740), .A4(n12739), .ZN(
        n12742) );
  OR4_X1 U14531 ( .A1(n15028), .A2(n12744), .A3(n12743), .A4(n12742), .ZN(
        n12745) );
  INV_X1 U14532 ( .A(n14842), .ZN(n13063) );
  XNOR2_X1 U14533 ( .A(n15174), .B(n13063), .ZN(n15056) );
  XNOR2_X1 U14534 ( .A(n15184), .B(n13061), .ZN(n15076) );
  NOR3_X1 U14535 ( .A1(n12745), .A2(n15056), .A3(n15076), .ZN(n12746) );
  XNOR2_X1 U14536 ( .A(n15147), .B(n14838), .ZN(n15007) );
  NAND4_X1 U14537 ( .A1(n14980), .A2(n15011), .A3(n12746), .A4(n15007), .ZN(
        n12747) );
  NOR2_X1 U14538 ( .A1(n14955), .A2(n12747), .ZN(n12748) );
  XNOR2_X1 U14539 ( .A(n15119), .B(n14834), .ZN(n14949) );
  XNOR2_X1 U14540 ( .A(n14972), .B(n14836), .ZN(n14970) );
  NAND4_X1 U14541 ( .A1(n14933), .A2(n12748), .A3(n14949), .A4(n14970), .ZN(
        n12749) );
  NOR2_X1 U14542 ( .A1(n12750), .A2(n12749), .ZN(n12751) );
  XNOR2_X1 U14543 ( .A(n13076), .B(n14832), .ZN(n13073) );
  NAND3_X1 U14544 ( .A1(n12772), .A2(n12751), .A3(n13073), .ZN(n12753) );
  XNOR2_X1 U14545 ( .A(n12753), .B(n12752), .ZN(n12755) );
  NAND2_X1 U14546 ( .A1(n12755), .A2(n12754), .ZN(n12768) );
  NAND2_X1 U14547 ( .A1(n12757), .A2(n12756), .ZN(n12766) );
  XNOR2_X1 U14548 ( .A(n12758), .B(n12761), .ZN(n12760) );
  NAND2_X1 U14549 ( .A1(n12760), .A2(n12759), .ZN(n12764) );
  NAND3_X1 U14550 ( .A1(n12762), .A2(n14914), .A3(n12761), .ZN(n12763) );
  NAND4_X1 U14551 ( .A1(n12766), .A2(n12765), .A3(n12764), .A4(n12763), .ZN(
        n12767) );
  NAND2_X1 U14552 ( .A1(n12768), .A2(n12767), .ZN(n12771) );
  NOR3_X1 U14553 ( .A1(n12771), .A2(n12779), .A3(n12774), .ZN(n12769) );
  AOI211_X1 U14554 ( .C1(n12773), .C2(n12772), .A(n12774), .B(n12771), .ZN(
        n12789) );
  INV_X1 U14555 ( .A(n12779), .ZN(n12776) );
  NOR4_X1 U14556 ( .A1(n12777), .A2(n12776), .A3(n12775), .A4(n12774), .ZN(
        n12788) );
  NOR3_X1 U14557 ( .A1(n12780), .A2(n12779), .A3(n12778), .ZN(n12787) );
  NAND2_X1 U14558 ( .A1(n12781), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15250) );
  NOR3_X1 U14559 ( .A1(n12782), .A2(n15250), .A3(n14785), .ZN(n12783) );
  AOI211_X1 U14560 ( .C1(n12785), .C2(n12784), .A(n13077), .B(n12783), .ZN(
        n12786) );
  NOR4_X1 U14561 ( .A1(n12789), .A2(n12788), .A3(n12787), .A4(n12786), .ZN(
        n12790) );
  XNOR2_X1 U14562 ( .A(n14001), .B(n8025), .ZN(n12812) );
  INV_X1 U14563 ( .A(n12812), .ZN(n12813) );
  XNOR2_X1 U14564 ( .A(n14005), .B(n8025), .ZN(n12810) );
  INV_X1 U14565 ( .A(n12810), .ZN(n12811) );
  XNOR2_X1 U14566 ( .A(n14017), .B(n12836), .ZN(n13597) );
  XNOR2_X1 U14567 ( .A(n13961), .B(n12836), .ZN(n13559) );
  NAND2_X1 U14568 ( .A1(n12794), .A2(n13959), .ZN(n13556) );
  AND2_X1 U14569 ( .A1(n13559), .A2(n13556), .ZN(n12795) );
  INV_X1 U14570 ( .A(n13947), .ZN(n12796) );
  MUX2_X1 U14571 ( .A(n12797), .B(n12796), .S(n8025), .Z(n12798) );
  XNOR2_X1 U14572 ( .A(n14097), .B(n12836), .ZN(n12799) );
  NAND2_X1 U14573 ( .A1(n12799), .A2(n13958), .ZN(n12802) );
  INV_X1 U14574 ( .A(n12799), .ZN(n12800) );
  NAND2_X1 U14575 ( .A1(n12800), .A2(n13927), .ZN(n12801) );
  NAND2_X1 U14576 ( .A1(n12802), .A2(n12801), .ZN(n13473) );
  XNOR2_X1 U14577 ( .A(n13918), .B(n12836), .ZN(n12803) );
  NAND2_X1 U14578 ( .A1(n12803), .A2(n13928), .ZN(n13514) );
  INV_X1 U14579 ( .A(n12803), .ZN(n12804) );
  NAND2_X1 U14580 ( .A1(n12804), .A2(n13899), .ZN(n13525) );
  NAND3_X1 U14581 ( .A1(n13514), .A2(n13519), .A3(n13597), .ZN(n12805) );
  XNOR2_X1 U14582 ( .A(n14089), .B(n8025), .ZN(n12808) );
  XNOR2_X1 U14583 ( .A(n12808), .B(n12807), .ZN(n13526) );
  XNOR2_X1 U14584 ( .A(n12810), .B(n13900), .ZN(n13580) );
  XNOR2_X1 U14585 ( .A(n12812), .B(n13887), .ZN(n13490) );
  XNOR2_X1 U14586 ( .A(n14080), .B(n12836), .ZN(n13548) );
  NAND2_X1 U14587 ( .A1(n13548), .A2(n13874), .ZN(n12815) );
  INV_X1 U14588 ( .A(n13548), .ZN(n12814) );
  XNOR2_X1 U14589 ( .A(n14074), .B(n8025), .ZN(n12816) );
  NOR2_X1 U14590 ( .A1(n12816), .A2(n13837), .ZN(n13498) );
  MUX2_X1 U14591 ( .A(n12817), .B(n12956), .S(n8025), .Z(n13497) );
  XNOR2_X1 U14592 ( .A(n14068), .B(n8025), .ZN(n12818) );
  INV_X1 U14593 ( .A(n12820), .ZN(n12821) );
  XOR2_X1 U14594 ( .A(n8025), .B(n13482), .Z(n12822) );
  NOR2_X1 U14595 ( .A1(n12823), .A2(n12822), .ZN(n12825) );
  INV_X1 U14596 ( .A(n12825), .ZN(n13538) );
  XNOR2_X1 U14597 ( .A(n14058), .B(n8025), .ZN(n12826) );
  NAND2_X1 U14598 ( .A1(n12826), .A2(n8379), .ZN(n12829) );
  INV_X1 U14599 ( .A(n12826), .ZN(n12827) );
  NAND2_X1 U14600 ( .A1(n12827), .A2(n13610), .ZN(n12828) );
  NAND2_X1 U14601 ( .A1(n12829), .A2(n12828), .ZN(n13537) );
  INV_X1 U14602 ( .A(n12829), .ZN(n13508) );
  XNOR2_X1 U14603 ( .A(n13809), .B(n8025), .ZN(n12830) );
  NAND2_X1 U14604 ( .A1(n12830), .A2(n13543), .ZN(n12833) );
  INV_X1 U14605 ( .A(n12830), .ZN(n12831) );
  NAND2_X1 U14606 ( .A1(n12831), .A2(n8037), .ZN(n12832) );
  XNOR2_X1 U14607 ( .A(n14048), .B(n12836), .ZN(n12834) );
  NOR2_X1 U14608 ( .A1(n12834), .A2(n13801), .ZN(n12835) );
  AOI21_X1 U14609 ( .B1(n12834), .B2(n13801), .A(n12835), .ZN(n13586) );
  XNOR2_X1 U14610 ( .A(n14042), .B(n12836), .ZN(n12837) );
  NOR2_X1 U14611 ( .A1(n12837), .A2(n13787), .ZN(n12838) );
  XNOR2_X1 U14612 ( .A(n13752), .B(n8025), .ZN(n12839) );
  INV_X1 U14613 ( .A(n12840), .ZN(n13754) );
  AOI22_X1 U14614 ( .A1(n13761), .A2(n13568), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12841) );
  OAI21_X1 U14615 ( .B1(n12842), .B2(n13600), .A(n12841), .ZN(n12844) );
  NOR2_X1 U14616 ( .A1(n14039), .A2(n13595), .ZN(n12843) );
  AOI211_X1 U14617 ( .C1(n13602), .C2(n13754), .A(n12844), .B(n12843), .ZN(
        n12845) );
  OAI21_X1 U14618 ( .B1(n12846), .B2(n13608), .A(n12845), .ZN(P3_U3160) );
  OAI222_X1 U14619 ( .A1(n12848), .A2(P2_U3088), .B1(n14691), .B2(n12847), 
        .C1(n13364), .C2(n14693), .ZN(P2_U3298) );
  INV_X1 U14620 ( .A(n12849), .ZN(n13018) );
  INV_X1 U14621 ( .A(n12850), .ZN(n12852) );
  NAND3_X1 U14622 ( .A1(n12854), .A2(n13771), .A3(n12853), .ZN(n12860) );
  NAND2_X1 U14623 ( .A1(n12860), .A2(n12855), .ZN(n12858) );
  INV_X1 U14624 ( .A(n12855), .ZN(n12856) );
  NOR2_X1 U14625 ( .A1(n7447), .A2(n12856), .ZN(n12857) );
  OR2_X1 U14626 ( .A1(n12860), .A2(n8257), .ZN(n13019) );
  INV_X1 U14627 ( .A(n13019), .ZN(n12967) );
  MUX2_X1 U14628 ( .A(n12862), .B(n12861), .S(n12974), .Z(n12966) );
  INV_X1 U14629 ( .A(n12870), .ZN(n12880) );
  NAND3_X1 U14630 ( .A1(n12866), .A2(n12865), .A3(n12863), .ZN(n12864) );
  AOI21_X1 U14631 ( .B1(n16100), .B2(n12864), .A(n16099), .ZN(n12874) );
  INV_X1 U14632 ( .A(n12865), .ZN(n12869) );
  INV_X1 U14633 ( .A(n12866), .ZN(n12867) );
  AOI21_X1 U14634 ( .B1(n12869), .B2(n12868), .A(n12867), .ZN(n12872) );
  OAI211_X1 U14635 ( .C1(n12872), .C2(n16099), .A(n12871), .B(n12870), .ZN(
        n12873) );
  MUX2_X1 U14636 ( .A(n12874), .B(n12873), .S(n12974), .Z(n12878) );
  AOI21_X1 U14637 ( .B1(n12877), .B2(n12875), .A(n12974), .ZN(n12876) );
  AOI21_X1 U14638 ( .B1(n12878), .B2(n12877), .A(n12876), .ZN(n12879) );
  AOI21_X1 U14639 ( .B1(n12880), .B2(n12960), .A(n12879), .ZN(n12885) );
  NAND2_X1 U14640 ( .A1(n16182), .A2(n12974), .ZN(n12883) );
  NAND2_X1 U14641 ( .A1(n12881), .A2(n12960), .ZN(n12882) );
  MUX2_X1 U14642 ( .A(n12883), .B(n12882), .S(n13620), .Z(n12884) );
  OAI211_X1 U14643 ( .C1(n12885), .C2(n13004), .A(n12997), .B(n12884), .ZN(
        n12890) );
  MUX2_X1 U14644 ( .A(n12887), .B(n12886), .S(n12960), .Z(n12889) );
  AOI21_X1 U14645 ( .B1(n12890), .B2(n12889), .A(n12888), .ZN(n12900) );
  NAND2_X1 U14646 ( .A1(n13618), .A2(n16215), .ZN(n12892) );
  MUX2_X1 U14647 ( .A(n12892), .B(n12891), .S(n12960), .Z(n12893) );
  NAND2_X1 U14648 ( .A1(n12894), .A2(n12893), .ZN(n12899) );
  NAND2_X1 U14649 ( .A1(n12895), .A2(n12974), .ZN(n12897) );
  NAND2_X1 U14650 ( .A1(n16231), .A2(n12960), .ZN(n12896) );
  MUX2_X1 U14651 ( .A(n12897), .B(n12896), .S(n13617), .Z(n12898) );
  OAI211_X1 U14652 ( .C1(n12900), .C2(n12899), .A(n13000), .B(n12898), .ZN(
        n12904) );
  MUX2_X1 U14653 ( .A(n12902), .B(n12901), .S(n12960), .Z(n12903) );
  NAND3_X1 U14654 ( .A1(n12904), .A2(n12998), .A3(n12903), .ZN(n12909) );
  INV_X1 U14655 ( .A(n12905), .ZN(n12906) );
  MUX2_X1 U14656 ( .A(n12907), .B(n12906), .S(n12974), .Z(n12908) );
  AOI21_X1 U14657 ( .B1(n12909), .B2(n12908), .A(n13011), .ZN(n12915) );
  NOR2_X1 U14658 ( .A1(n13614), .A2(n12960), .ZN(n12912) );
  NOR2_X1 U14659 ( .A1(n12910), .A2(n12974), .ZN(n12911) );
  MUX2_X1 U14660 ( .A(n12912), .B(n12911), .S(n16295), .Z(n12914) );
  NOR3_X1 U14661 ( .A1(n12915), .A2(n12914), .A3(n12913), .ZN(n12924) );
  NAND2_X1 U14662 ( .A1(n12921), .A2(n12916), .ZN(n12919) );
  NAND2_X1 U14663 ( .A1(n12920), .A2(n12917), .ZN(n12918) );
  MUX2_X1 U14664 ( .A(n12919), .B(n12918), .S(n12960), .Z(n12923) );
  MUX2_X1 U14665 ( .A(n12921), .B(n12920), .S(n12974), .Z(n12922) );
  OAI21_X1 U14666 ( .B1(n12924), .B2(n12923), .A(n12922), .ZN(n12931) );
  NOR2_X1 U14667 ( .A1(n13939), .A2(n13961), .ZN(n12930) );
  INV_X1 U14668 ( .A(n12925), .ZN(n12926) );
  NOR2_X1 U14669 ( .A1(n12927), .A2(n12926), .ZN(n12928) );
  MUX2_X1 U14670 ( .A(n7597), .B(n12928), .S(n12960), .Z(n12929) );
  AOI21_X1 U14671 ( .B1(n12931), .B2(n12930), .A(n12929), .ZN(n12935) );
  MUX2_X1 U14672 ( .A(n12933), .B(n12932), .S(n12974), .Z(n12934) );
  OAI211_X1 U14673 ( .C1(n12935), .C2(n9244), .A(n7729), .B(n12934), .ZN(
        n12938) );
  INV_X1 U14674 ( .A(n13918), .ZN(n14013) );
  MUX2_X1 U14675 ( .A(n12960), .B(n14013), .S(n13928), .Z(n12936) );
  OAI21_X1 U14676 ( .B1(n12974), .B2(n13918), .A(n12936), .ZN(n12937) );
  AOI211_X1 U14677 ( .C1(n12938), .C2(n12937), .A(n13885), .B(n9246), .ZN(
        n12950) );
  INV_X1 U14678 ( .A(n12939), .ZN(n12941) );
  OAI211_X1 U14679 ( .C1(n12941), .C2(n12940), .A(n12947), .B(n12942), .ZN(
        n12945) );
  AOI21_X1 U14680 ( .B1(n13913), .B2(n14089), .A(n12941), .ZN(n12943) );
  OAI21_X1 U14681 ( .B1(n12943), .B2(n8195), .A(n12946), .ZN(n12944) );
  MUX2_X1 U14682 ( .A(n12945), .B(n12944), .S(n12974), .Z(n12949) );
  MUX2_X1 U14683 ( .A(n12947), .B(n12946), .S(n12960), .Z(n12948) );
  OAI211_X1 U14684 ( .C1(n12950), .C2(n12949), .A(n13860), .B(n12948), .ZN(
        n12954) );
  MUX2_X1 U14685 ( .A(n12952), .B(n12951), .S(n12974), .Z(n12953) );
  NAND3_X1 U14686 ( .A1(n12954), .A2(n13850), .A3(n12953), .ZN(n12959) );
  MUX2_X1 U14687 ( .A(n12956), .B(n12955), .S(n12960), .Z(n12958) );
  INV_X1 U14688 ( .A(n12957), .ZN(n12961) );
  AOI21_X1 U14689 ( .B1(n12959), .B2(n12958), .A(n13834), .ZN(n12964) );
  MUX2_X1 U14690 ( .A(n12962), .B(n12961), .S(n12960), .Z(n12963) );
  OR3_X1 U14691 ( .A1(n12964), .A2(n12963), .A3(n13825), .ZN(n12965) );
  MUX2_X1 U14692 ( .A(n12970), .B(n12969), .S(n12974), .Z(n12971) );
  NAND3_X1 U14693 ( .A1(n13018), .A2(n12972), .A3(n12971), .ZN(n12973) );
  AND2_X1 U14694 ( .A1(n12973), .A2(n13028), .ZN(n12975) );
  INV_X1 U14695 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n14682) );
  OAI22_X1 U14696 ( .A1(n15244), .A2(n14682), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12980) );
  XNOR2_X1 U14697 ( .A(n12979), .B(n12980), .ZN(n13464) );
  NAND2_X1 U14698 ( .A1(n9092), .A2(SI_30_), .ZN(n12978) );
  NAND2_X1 U14699 ( .A1(n16409), .A2(n13025), .ZN(n13017) );
  OAI21_X1 U14700 ( .B1(n14682), .B2(P2_DATAO_REG_30__SCAN_IN), .A(n12981), 
        .ZN(n12984) );
  AOI22_X1 U14701 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(
        P1_DATAO_REG_31__SCAN_IN), .B1(n12982), .B2(n15241), .ZN(n12983) );
  XNOR2_X1 U14702 ( .A(n12984), .B(n12983), .ZN(n14111) );
  NAND2_X1 U14703 ( .A1(n14111), .A2(n8822), .ZN(n12986) );
  NAND2_X1 U14704 ( .A1(n9092), .A2(SI_31_), .ZN(n12985) );
  INV_X1 U14705 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12991) );
  NAND2_X1 U14706 ( .A1(n8812), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12990) );
  INV_X1 U14707 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12987) );
  OR2_X1 U14708 ( .A1(n12988), .A2(n12987), .ZN(n12989) );
  OAI211_X1 U14709 ( .C1(n12992), .C2(n12991), .A(n12990), .B(n12989), .ZN(
        n12993) );
  INV_X1 U14710 ( .A(n12993), .ZN(n12994) );
  NAND2_X1 U14711 ( .A1(n12995), .A2(n12994), .ZN(n13736) );
  OR2_X1 U14712 ( .A1(n16409), .A2(n13025), .ZN(n13029) );
  OAI21_X1 U14713 ( .B1(n13739), .B2(n13736), .A(n13029), .ZN(n13020) );
  NAND2_X1 U14714 ( .A1(n13739), .A2(n13736), .ZN(n13027) );
  INV_X1 U14715 ( .A(n16099), .ZN(n16097) );
  NAND3_X1 U14716 ( .A1(n12998), .A2(n16097), .A3(n12997), .ZN(n13003) );
  INV_X1 U14717 ( .A(n16050), .ZN(n16056) );
  NAND4_X1 U14718 ( .A1(n16056), .A2(n13001), .A3(n13000), .A4(n12999), .ZN(
        n13002) );
  NOR2_X1 U14719 ( .A1(n13003), .A2(n13002), .ZN(n13009) );
  NOR2_X1 U14720 ( .A1(n13005), .A2(n13004), .ZN(n13007) );
  NAND4_X1 U14721 ( .A1(n13009), .A2(n13008), .A3(n13007), .A4(n13006), .ZN(
        n13012) );
  NOR4_X1 U14722 ( .A1(n13012), .A2(n13011), .A3(n8200), .A4(n13961), .ZN(
        n13013) );
  NAND4_X1 U14723 ( .A1(n13013), .A2(n13922), .A3(n13948), .A4(n7729), .ZN(
        n13014) );
  NOR2_X1 U14724 ( .A1(n13885), .A2(n13014), .ZN(n13015) );
  NAND4_X1 U14725 ( .A1(n13850), .A2(n13901), .A3(n13876), .A4(n13015), .ZN(
        n13016) );
  XNOR2_X1 U14726 ( .A(n13022), .B(n13021), .ZN(n13035) );
  INV_X1 U14727 ( .A(n13736), .ZN(n13030) );
  OAI21_X1 U14728 ( .B1(n13025), .B2(n13030), .A(n16409), .ZN(n13026) );
  INV_X1 U14729 ( .A(n13029), .ZN(n13031) );
  OAI21_X1 U14730 ( .B1(n13031), .B2(n13030), .A(n16416), .ZN(n13032) );
  NOR3_X1 U14731 ( .A1(n13039), .A2(n13038), .A3(n13037), .ZN(n13042) );
  OAI21_X1 U14732 ( .B1(n13043), .B2(n13040), .A(P3_B_REG_SCAN_IN), .ZN(n13041) );
  NAND2_X1 U14733 ( .A1(n15190), .A2(n14844), .ZN(n13044) );
  OR2_X1 U14734 ( .A1(n15184), .A2(n14843), .ZN(n13046) );
  OR2_X1 U14735 ( .A1(n15174), .A2(n14842), .ZN(n13047) );
  NAND2_X1 U14736 ( .A1(n15049), .A2(n14841), .ZN(n13049) );
  OR2_X1 U14737 ( .A1(n15159), .A2(n14840), .ZN(n13050) );
  INV_X1 U14738 ( .A(n15011), .ZN(n15013) );
  OR2_X1 U14739 ( .A1(n15155), .A2(n14839), .ZN(n13051) );
  NAND2_X1 U14740 ( .A1(n15147), .A2(n14838), .ZN(n13053) );
  INV_X1 U14741 ( .A(n14970), .ZN(n14967) );
  NAND2_X1 U14742 ( .A1(n14966), .A2(n8719), .ZN(n14956) );
  INV_X1 U14743 ( .A(n14933), .ZN(n14923) );
  NAND2_X1 U14744 ( .A1(n15190), .A2(n13058), .ZN(n13059) );
  OR2_X1 U14745 ( .A1(n15184), .A2(n13061), .ZN(n13062) );
  INV_X1 U14746 ( .A(n13064), .ZN(n15042) );
  OR2_X2 U14747 ( .A1(n15041), .A2(n15042), .ZN(n15040) );
  INV_X1 U14748 ( .A(n14841), .ZN(n13065) );
  OR2_X1 U14749 ( .A1(n15049), .A2(n13065), .ZN(n13066) );
  NAND2_X1 U14750 ( .A1(n15155), .A2(n14715), .ZN(n13067) );
  INV_X1 U14751 ( .A(n14838), .ZN(n14788) );
  NAND2_X1 U14752 ( .A1(n15147), .A2(n14788), .ZN(n13069) );
  INV_X1 U14753 ( .A(n14980), .ZN(n14984) );
  OAI21_X1 U14754 ( .B1(n14698), .B2(n14812), .A(n14953), .ZN(n13070) );
  NAND2_X1 U14755 ( .A1(n14934), .A2(n14933), .ZN(n14932) );
  INV_X1 U14756 ( .A(n14833), .ZN(n14699) );
  INV_X1 U14757 ( .A(n15115), .ZN(n13075) );
  AOI211_X1 U14758 ( .C1(n13076), .C2(n14926), .A(n16142), .B(n14918), .ZN(
        n15110) );
  NAND2_X1 U14759 ( .A1(n15110), .A2(n16341), .ZN(n13087) );
  NAND2_X1 U14760 ( .A1(n14833), .A2(n14806), .ZN(n15106) );
  OR2_X1 U14761 ( .A1(n13078), .A2(n13077), .ZN(n13079) );
  AND2_X1 U14762 ( .A1(n14807), .A2(n13079), .ZN(n14913) );
  NAND2_X1 U14763 ( .A1(n14831), .A2(n14913), .ZN(n15107) );
  NOR3_X1 U14764 ( .A1(n13081), .A2(n13080), .A3(n15107), .ZN(n13082) );
  AOI21_X1 U14765 ( .B1(n16336), .B2(n13083), .A(n13082), .ZN(n13084) );
  OAI21_X1 U14766 ( .B1(n16347), .B2(n15106), .A(n13084), .ZN(n13085) );
  AOI21_X1 U14767 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n16347), .A(n13085), 
        .ZN(n13086) );
  OAI211_X1 U14768 ( .C1(n15108), .C2(n16163), .A(n13087), .B(n13086), .ZN(
        n13088) );
  AOI21_X1 U14769 ( .B1(n15111), .B2(n15090), .A(n13088), .ZN(n13089) );
  OAI21_X1 U14770 ( .B1(n15112), .B2(n15054), .A(n13089), .ZN(P1_U3356) );
  NAND2_X1 U14771 ( .A1(n13091), .A2(n13090), .ZN(n13352) );
  NAND3_X1 U14772 ( .A1(n13421), .A2(n13350), .A3(n14301), .ZN(n13092) );
  NAND2_X1 U14773 ( .A1(n13352), .A2(n13092), .ZN(n13418) );
  INV_X1 U14774 ( .A(n13116), .ZN(n13119) );
  NAND2_X1 U14775 ( .A1(n13119), .A2(n13093), .ZN(n13094) );
  AOI22_X1 U14776 ( .A1(n13094), .A2(n14301), .B1(n13451), .B2(n13421), .ZN(
        n13417) );
  NAND2_X1 U14777 ( .A1(n13095), .A2(n9720), .ZN(n13098) );
  OR2_X1 U14778 ( .A1(n8004), .A2(n13096), .ZN(n13097) );
  INV_X4 U14779 ( .A(n13349), .ZN(n13360) );
  NOR2_X1 U14780 ( .A1(n13100), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n13101) );
  OR2_X1 U14781 ( .A1(n13268), .A2(n13101), .ZN(n14209) );
  INV_X1 U14782 ( .A(n14209), .ZN(n14491) );
  NAND2_X1 U14783 ( .A1(n14491), .A2(n9789), .ZN(n13107) );
  INV_X1 U14784 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n13104) );
  NAND2_X1 U14785 ( .A1(n13368), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n13103) );
  NAND2_X1 U14786 ( .A1(n13386), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n13102) );
  OAI211_X1 U14787 ( .C1(n13346), .C2(n13104), .A(n13103), .B(n13102), .ZN(
        n13105) );
  INV_X1 U14788 ( .A(n13105), .ZN(n13106) );
  INV_X1 U14789 ( .A(n13242), .ZN(n13247) );
  NAND2_X1 U14790 ( .A1(n13108), .A2(n9720), .ZN(n13111) );
  AOI22_X1 U14791 ( .A1(n9659), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n13109), 
        .B2(n14301), .ZN(n13110) );
  OAI22_X1 U14792 ( .A1(n14667), .A2(n13411), .B1(n14524), .B2(n13341), .ZN(
        n13240) );
  NAND2_X1 U14793 ( .A1(n13349), .A2(n14224), .ZN(n13113) );
  NAND2_X1 U14794 ( .A1(n14265), .A2(n13360), .ZN(n13112) );
  NAND2_X1 U14795 ( .A1(n13360), .A2(n14224), .ZN(n13115) );
  NAND2_X1 U14796 ( .A1(n13349), .A2(n14265), .ZN(n13114) );
  NAND2_X1 U14797 ( .A1(n13115), .A2(n13114), .ZN(n13135) );
  NAND2_X1 U14798 ( .A1(n13136), .A2(n13135), .ZN(n13134) );
  NAND2_X1 U14799 ( .A1(n13118), .A2(n13117), .ZN(n13120) );
  NAND2_X1 U14800 ( .A1(n9885), .A2(n13119), .ZN(n13122) );
  NAND2_X1 U14801 ( .A1(n13120), .A2(n13122), .ZN(n13124) );
  NAND2_X1 U14802 ( .A1(n13124), .A2(n13123), .ZN(n13130) );
  NAND2_X1 U14803 ( .A1(n13349), .A2(n14547), .ZN(n13126) );
  NAND2_X1 U14804 ( .A1(n14266), .A2(n13360), .ZN(n13125) );
  NAND2_X1 U14805 ( .A1(n13349), .A2(n14266), .ZN(n13128) );
  NAND2_X1 U14806 ( .A1(n13360), .A2(n14547), .ZN(n13127) );
  NAND2_X1 U14807 ( .A1(n13128), .A2(n13127), .ZN(n13129) );
  NAND2_X1 U14808 ( .A1(n13131), .A2(n13130), .ZN(n13132) );
  NAND3_X1 U14809 ( .A1(n13134), .A2(n13133), .A3(n13132), .ZN(n13140) );
  INV_X1 U14810 ( .A(n13135), .ZN(n13138) );
  INV_X1 U14811 ( .A(n13136), .ZN(n13137) );
  NAND2_X1 U14812 ( .A1(n13138), .A2(n13137), .ZN(n13139) );
  NAND2_X1 U14813 ( .A1(n13349), .A2(n16169), .ZN(n13142) );
  NAND2_X1 U14814 ( .A1(n14264), .A2(n13360), .ZN(n13141) );
  NAND2_X1 U14815 ( .A1(n13142), .A2(n13141), .ZN(n13147) );
  INV_X1 U14816 ( .A(n13360), .ZN(n13392) );
  AOI22_X1 U14817 ( .A1(n14264), .A2(n13392), .B1(n13360), .B2(n16169), .ZN(
        n13143) );
  NAND2_X1 U14818 ( .A1(n13146), .A2(n13360), .ZN(n13145) );
  NAND2_X1 U14819 ( .A1(n13349), .A2(n14263), .ZN(n13144) );
  NAND2_X1 U14820 ( .A1(n13145), .A2(n13144), .ZN(n13148) );
  AOI22_X1 U14821 ( .A1(n13146), .A2(n13392), .B1(n13360), .B2(n14263), .ZN(
        n13149) );
  INV_X1 U14822 ( .A(n13148), .ZN(n13151) );
  INV_X1 U14823 ( .A(n13149), .ZN(n13150) );
  NAND2_X1 U14824 ( .A1(n13151), .A2(n13150), .ZN(n13152) );
  NAND2_X1 U14825 ( .A1(n13155), .A2(n13392), .ZN(n13154) );
  NAND2_X1 U14826 ( .A1(n14262), .A2(n13360), .ZN(n13153) );
  NAND2_X1 U14827 ( .A1(n13155), .A2(n13360), .ZN(n13156) );
  OAI21_X1 U14828 ( .B1(n13157), .B2(n13360), .A(n13156), .ZN(n13158) );
  NAND2_X1 U14829 ( .A1(n16223), .A2(n13360), .ZN(n13161) );
  NAND2_X1 U14830 ( .A1(n13392), .A2(n14261), .ZN(n13160) );
  NAND2_X1 U14831 ( .A1(n13161), .A2(n13160), .ZN(n13163) );
  AOI22_X1 U14832 ( .A1(n16223), .A2(n13392), .B1(n13360), .B2(n14261), .ZN(
        n13162) );
  NAND2_X1 U14833 ( .A1(n16246), .A2(n13341), .ZN(n13165) );
  NAND2_X1 U14834 ( .A1(n14260), .A2(n13360), .ZN(n13164) );
  NAND2_X1 U14835 ( .A1(n13165), .A2(n13164), .ZN(n13171) );
  NAND2_X1 U14836 ( .A1(n13170), .A2(n13171), .ZN(n13169) );
  NAND2_X1 U14837 ( .A1(n16246), .A2(n13360), .ZN(n13166) );
  OAI21_X1 U14838 ( .B1(n13167), .B2(n13360), .A(n13166), .ZN(n13168) );
  NAND2_X1 U14839 ( .A1(n13169), .A2(n13168), .ZN(n13175) );
  INV_X1 U14840 ( .A(n13170), .ZN(n13173) );
  INV_X1 U14841 ( .A(n13171), .ZN(n13172) );
  NAND2_X1 U14842 ( .A1(n13173), .A2(n13172), .ZN(n13174) );
  NAND2_X1 U14843 ( .A1(n13178), .A2(n13360), .ZN(n13177) );
  NAND2_X1 U14844 ( .A1(n13349), .A2(n14259), .ZN(n13176) );
  NAND2_X1 U14845 ( .A1(n13177), .A2(n13176), .ZN(n13180) );
  AOI22_X1 U14846 ( .A1(n13178), .A2(n13392), .B1(n13360), .B2(n14259), .ZN(
        n13179) );
  NAND2_X1 U14847 ( .A1(n13183), .A2(n13341), .ZN(n13182) );
  NAND2_X1 U14848 ( .A1(n14258), .A2(n13360), .ZN(n13181) );
  NAND2_X1 U14849 ( .A1(n13182), .A2(n13181), .ZN(n13187) );
  NAND2_X1 U14850 ( .A1(n13183), .A2(n13360), .ZN(n13184) );
  OAI21_X1 U14851 ( .B1(n13185), .B2(n13360), .A(n13184), .ZN(n13186) );
  NAND2_X1 U14852 ( .A1(n16304), .A2(n13360), .ZN(n13189) );
  NAND2_X1 U14853 ( .A1(n13349), .A2(n14257), .ZN(n13188) );
  NAND2_X1 U14854 ( .A1(n13189), .A2(n13188), .ZN(n13191) );
  AOI22_X1 U14855 ( .A1(n16304), .A2(n13392), .B1(n13360), .B2(n14257), .ZN(
        n13190) );
  NOR2_X1 U14856 ( .A1(n13192), .A2(n13191), .ZN(n13193) );
  NAND2_X1 U14857 ( .A1(n13197), .A2(n13341), .ZN(n13196) );
  NAND2_X1 U14858 ( .A1(n14256), .A2(n13411), .ZN(n13195) );
  AOI22_X1 U14859 ( .A1(n13197), .A2(n13411), .B1(n14256), .B2(n13341), .ZN(
        n13198) );
  NAND2_X1 U14860 ( .A1(n13202), .A2(n13360), .ZN(n13201) );
  NAND2_X1 U14861 ( .A1(n13349), .A2(n14255), .ZN(n13200) );
  NAND2_X1 U14862 ( .A1(n13201), .A2(n13200), .ZN(n13207) );
  NAND2_X1 U14863 ( .A1(n13202), .A2(n13341), .ZN(n13203) );
  OAI21_X1 U14864 ( .B1(n13204), .B2(n13341), .A(n13203), .ZN(n13205) );
  NAND2_X1 U14865 ( .A1(n16392), .A2(n13341), .ZN(n13209) );
  NAND2_X1 U14866 ( .A1(n14254), .A2(n13360), .ZN(n13208) );
  NAND2_X1 U14867 ( .A1(n13209), .A2(n13208), .ZN(n13213) );
  AOI22_X1 U14868 ( .A1(n16392), .A2(n13411), .B1(n14254), .B2(n13341), .ZN(
        n13210) );
  INV_X1 U14869 ( .A(n13210), .ZN(n13211) );
  INV_X1 U14870 ( .A(n13213), .ZN(n13214) );
  OAI22_X1 U14871 ( .A1(n13216), .A2(n13341), .B1(n13215), .B2(n13411), .ZN(
        n13219) );
  AOI22_X1 U14872 ( .A1(n13217), .A2(n13392), .B1(n13411), .B2(n14253), .ZN(
        n13218) );
  AOI22_X1 U14873 ( .A1(n13221), .A2(n13392), .B1(n13360), .B2(n14252), .ZN(
        n13225) );
  OAI22_X1 U14874 ( .A1(n13223), .A2(n13341), .B1(n13222), .B2(n13411), .ZN(
        n13224) );
  INV_X1 U14875 ( .A(n13230), .ZN(n13233) );
  OAI22_X1 U14876 ( .A1(n13227), .A2(n13341), .B1(n13226), .B2(n13411), .ZN(
        n13229) );
  INV_X1 U14877 ( .A(n13229), .ZN(n13232) );
  AOI22_X1 U14878 ( .A1(n14633), .A2(n13341), .B1(n13360), .B2(n14251), .ZN(
        n13228) );
  AOI21_X1 U14879 ( .B1(n13230), .B2(n13229), .A(n13228), .ZN(n13231) );
  AOI22_X1 U14880 ( .A1(n14336), .A2(n13341), .B1(n13360), .B2(n14324), .ZN(
        n13235) );
  INV_X1 U14881 ( .A(n14324), .ZN(n14522) );
  OAI22_X1 U14882 ( .A1(n14674), .A2(n13341), .B1(n14522), .B2(n13411), .ZN(
        n13234) );
  OAI22_X1 U14883 ( .A1(n14619), .A2(n13341), .B1(n14326), .B2(n13411), .ZN(
        n13237) );
  OAI22_X1 U14884 ( .A1(n14619), .A2(n13411), .B1(n14326), .B2(n13341), .ZN(
        n13239) );
  INV_X1 U14885 ( .A(n13237), .ZN(n13238) );
  OAI22_X1 U14886 ( .A1(n14667), .A2(n13341), .B1(n14524), .B2(n13411), .ZN(
        n13241) );
  NAND2_X1 U14887 ( .A1(n13243), .A2(n13242), .ZN(n13245) );
  OAI22_X1 U14888 ( .A1(n14493), .A2(n13411), .B1(n14345), .B2(n13341), .ZN(
        n13244) );
  AOI22_X1 U14889 ( .A1(n13247), .A2(n13246), .B1(n13245), .B2(n13244), .ZN(
        n13260) );
  OR2_X1 U14890 ( .A1(n13248), .A2(n13321), .ZN(n13251) );
  OR2_X1 U14891 ( .A1(n8004), .A2(n13249), .ZN(n13250) );
  INV_X1 U14892 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13252) );
  XNOR2_X1 U14893 ( .A(n13268), .B(n13252), .ZN(n14474) );
  NAND2_X1 U14894 ( .A1(n14474), .A2(n9789), .ZN(n13258) );
  INV_X1 U14895 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n13255) );
  NAND2_X1 U14896 ( .A1(n13386), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n13254) );
  NAND2_X1 U14897 ( .A1(n13368), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n13253) );
  OAI211_X1 U14898 ( .C1(n13255), .C2(n13346), .A(n13254), .B(n13253), .ZN(
        n13256) );
  INV_X1 U14899 ( .A(n13256), .ZN(n13257) );
  OAI22_X1 U14900 ( .A1(n14476), .A2(n13411), .B1(n14487), .B2(n13341), .ZN(
        n13259) );
  OAI22_X1 U14901 ( .A1(n14476), .A2(n13341), .B1(n14487), .B2(n13411), .ZN(
        n13261) );
  OR2_X1 U14902 ( .A1(n8004), .A2(n13263), .ZN(n13264) );
  NAND2_X1 U14903 ( .A1(n13268), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n13266) );
  INV_X1 U14904 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n14216) );
  NAND2_X1 U14905 ( .A1(n13266), .A2(n14216), .ZN(n13269) );
  AND2_X1 U14906 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .ZN(n13267) );
  NAND2_X1 U14907 ( .A1(n13268), .A2(n13267), .ZN(n13281) );
  NAND2_X1 U14908 ( .A1(n13269), .A2(n13281), .ZN(n14459) );
  OR2_X1 U14909 ( .A1(n14459), .A2(n13309), .ZN(n13275) );
  INV_X1 U14910 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n13272) );
  NAND2_X1 U14911 ( .A1(n13368), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n13271) );
  NAND2_X1 U14912 ( .A1(n13386), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n13270) );
  OAI211_X1 U14913 ( .C1(n13346), .C2(n13272), .A(n13271), .B(n13270), .ZN(
        n13273) );
  INV_X1 U14914 ( .A(n13273), .ZN(n13274) );
  NAND2_X1 U14915 ( .A1(n13275), .A2(n13274), .ZN(n14437) );
  AOI22_X1 U14916 ( .A1(n14599), .A2(n13411), .B1(n14437), .B2(n13341), .ZN(
        n13276) );
  INV_X1 U14917 ( .A(n14599), .ZN(n14463) );
  OAI22_X1 U14918 ( .A1(n14463), .A2(n13411), .B1(n14350), .B2(n13341), .ZN(
        n13277) );
  OR2_X1 U14919 ( .A1(n8004), .A2(n13279), .ZN(n13280) );
  INV_X1 U14920 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n14159) );
  NAND2_X1 U14921 ( .A1(n13281), .A2(n14159), .ZN(n13282) );
  AND2_X1 U14922 ( .A1(n13298), .A2(n13282), .ZN(n14447) );
  NAND2_X1 U14923 ( .A1(n14447), .A2(n9789), .ZN(n13287) );
  INV_X1 U14924 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n14595) );
  NAND2_X1 U14925 ( .A1(n13386), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n13284) );
  NAND2_X1 U14926 ( .A1(n13368), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n13283) );
  OAI211_X1 U14927 ( .C1(n14595), .C2(n13346), .A(n13284), .B(n13283), .ZN(
        n13285) );
  INV_X1 U14928 ( .A(n13285), .ZN(n13286) );
  NAND2_X1 U14929 ( .A1(n13287), .A2(n13286), .ZN(n14352) );
  AOI22_X1 U14930 ( .A1(n14446), .A2(n13341), .B1(n13360), .B2(n14352), .ZN(
        n13290) );
  AOI22_X1 U14931 ( .A1(n14446), .A2(n13411), .B1(n14352), .B2(n13341), .ZN(
        n13288) );
  INV_X1 U14932 ( .A(n13288), .ZN(n13289) );
  NAND2_X1 U14933 ( .A1(n13291), .A2(n13290), .ZN(n13292) );
  OR2_X1 U14934 ( .A1(n13293), .A2(n13321), .ZN(n13296) );
  OR2_X1 U14935 ( .A1(n8004), .A2(n13294), .ZN(n13295) );
  INV_X1 U14936 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13297) );
  AND2_X1 U14937 ( .A1(n13298), .A2(n13297), .ZN(n13299) );
  NOR2_X1 U14938 ( .A1(n13299), .A2(n13307), .ZN(n14428) );
  INV_X1 U14939 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n14590) );
  NAND2_X1 U14940 ( .A1(n13368), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n13301) );
  NAND2_X1 U14941 ( .A1(n13386), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n13300) );
  OAI211_X1 U14942 ( .C1(n13346), .C2(n14590), .A(n13301), .B(n13300), .ZN(
        n13302) );
  AOI21_X1 U14943 ( .B1(n14428), .B2(n9789), .A(n13302), .ZN(n14353) );
  OAI22_X1 U14944 ( .A1(n14657), .A2(n13360), .B1(n14353), .B2(n13341), .ZN(
        n13303) );
  NAND2_X1 U14945 ( .A1(n14689), .A2(n9720), .ZN(n13306) );
  OR2_X1 U14946 ( .A1(n8004), .A2(n14692), .ZN(n13305) );
  OR2_X1 U14947 ( .A1(n13307), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n13308) );
  NAND2_X1 U14948 ( .A1(n13307), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n13325) );
  NAND2_X1 U14949 ( .A1(n13308), .A2(n13325), .ZN(n14413) );
  INV_X1 U14950 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n14585) );
  NAND2_X1 U14951 ( .A1(n13368), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n13311) );
  NAND2_X1 U14952 ( .A1(n13386), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n13310) );
  OAI211_X1 U14953 ( .C1(n13346), .C2(n14585), .A(n13311), .B(n13310), .ZN(
        n13312) );
  INV_X1 U14954 ( .A(n13312), .ZN(n13313) );
  OAI22_X1 U14955 ( .A1(n14653), .A2(n13360), .B1(n13315), .B2(n13341), .ZN(
        n13318) );
  AOI22_X1 U14956 ( .A1(n14412), .A2(n13411), .B1(n14354), .B2(n13341), .ZN(
        n13316) );
  AOI21_X1 U14957 ( .B1(n13319), .B2(n13318), .A(n13316), .ZN(n13317) );
  NOR2_X1 U14958 ( .A1(n13319), .A2(n13318), .ZN(n13320) );
  OR2_X1 U14959 ( .A1(n15255), .A2(n13321), .ZN(n13323) );
  OR2_X1 U14960 ( .A1(n8004), .A2(n14687), .ZN(n13322) );
  NAND2_X1 U14961 ( .A1(n9742), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n13330) );
  INV_X1 U14962 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13326) );
  INV_X1 U14963 ( .A(n13325), .ZN(n13324) );
  NAND2_X1 U14964 ( .A1(n13324), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n13336) );
  INV_X1 U14965 ( .A(n13336), .ZN(n13367) );
  AOI21_X1 U14966 ( .B1(n13326), .B2(n13325), .A(n13367), .ZN(n14398) );
  NAND2_X1 U14967 ( .A1(n9789), .A2(n14398), .ZN(n13329) );
  NAND2_X1 U14968 ( .A1(n13386), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n13328) );
  NAND2_X1 U14969 ( .A1(n13368), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n13327) );
  OAI22_X1 U14970 ( .A1(n14401), .A2(n13341), .B1(n14355), .B2(n13360), .ZN(
        n13331) );
  AOI22_X1 U14971 ( .A1(n14580), .A2(n13392), .B1(n13360), .B2(n14330), .ZN(
        n13332) );
  NAND2_X1 U14972 ( .A1(n15249), .A2(n9720), .ZN(n13335) );
  OR2_X1 U14973 ( .A1(n8004), .A2(n13333), .ZN(n13334) );
  NAND2_X1 U14974 ( .A1(n9742), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n13340) );
  XNOR2_X1 U14975 ( .A(P2_REG3_REG_27__SCAN_IN), .B(n13336), .ZN(n14151) );
  NAND2_X1 U14976 ( .A1(n11931), .A2(n14151), .ZN(n13339) );
  NAND2_X1 U14977 ( .A1(n13386), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n13338) );
  NAND2_X1 U14978 ( .A1(n13368), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n13337) );
  AOI22_X1 U14979 ( .A1(n14574), .A2(n13341), .B1(n13360), .B2(n14356), .ZN(
        n13406) );
  OAI22_X1 U14980 ( .A1(n14383), .A2(n13341), .B1(n14180), .B2(n13360), .ZN(
        n13405) );
  NAND2_X1 U14981 ( .A1(n15236), .A2(n9720), .ZN(n13343) );
  OR2_X1 U14982 ( .A1(n8004), .A2(n12982), .ZN(n13342) );
  INV_X1 U14983 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n14556) );
  NAND2_X1 U14984 ( .A1(n13368), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n13345) );
  NAND2_X1 U14985 ( .A1(n13386), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n13344) );
  OAI211_X1 U14986 ( .C1(n13346), .C2(n14556), .A(n13345), .B(n13344), .ZN(
        n14316) );
  XNOR2_X1 U14987 ( .A(n14311), .B(n14316), .ZN(n13449) );
  NAND2_X1 U14988 ( .A1(n14681), .A2(n9720), .ZN(n13348) );
  OR2_X1 U14989 ( .A1(n8004), .A2(n14682), .ZN(n13347) );
  NAND2_X1 U14990 ( .A1(n13349), .A2(n14316), .ZN(n13410) );
  AND2_X1 U14991 ( .A1(n13351), .A2(n13350), .ZN(n13353) );
  AND2_X1 U14992 ( .A1(n13353), .A2(n13352), .ZN(n13357) );
  NAND2_X1 U14993 ( .A1(n9742), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n13356) );
  NAND2_X1 U14994 ( .A1(n13368), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n13355) );
  NAND2_X1 U14995 ( .A1(n13386), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n13354) );
  AND3_X1 U14996 ( .A1(n13356), .A2(n13355), .A3(n13354), .ZN(n13359) );
  AOI21_X1 U14997 ( .B1(n13410), .B2(n13357), .A(n13359), .ZN(n13358) );
  AOI21_X1 U14998 ( .B1(n14310), .B2(n13411), .A(n13358), .ZN(n13409) );
  NAND2_X1 U14999 ( .A1(n14310), .A2(n13341), .ZN(n13362) );
  INV_X1 U15000 ( .A(n13359), .ZN(n14362) );
  NAND2_X1 U15001 ( .A1(n13360), .A2(n14362), .ZN(n13361) );
  NAND2_X1 U15002 ( .A1(n13362), .A2(n13361), .ZN(n13408) );
  NAND2_X1 U15003 ( .A1(n13363), .A2(n9720), .ZN(n13366) );
  OR2_X1 U15004 ( .A1(n8004), .A2(n13364), .ZN(n13365) );
  NAND2_X1 U15005 ( .A1(n9742), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n13372) );
  NAND2_X1 U15006 ( .A1(n9789), .A2(n14333), .ZN(n13371) );
  NAND2_X1 U15007 ( .A1(n13386), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n13370) );
  NAND2_X1 U15008 ( .A1(n13368), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n13369) );
  NAND4_X1 U15009 ( .A1(n13372), .A2(n13371), .A3(n13370), .A4(n13369), .ZN(
        n14250) );
  AND2_X1 U15010 ( .A1(n13392), .A2(n14250), .ZN(n13373) );
  AOI21_X1 U15011 ( .B1(n14563), .B2(n13411), .A(n13373), .ZN(n13402) );
  NAND2_X1 U15012 ( .A1(n14563), .A2(n13341), .ZN(n13375) );
  NAND2_X1 U15013 ( .A1(n14250), .A2(n13360), .ZN(n13374) );
  NAND2_X1 U15014 ( .A1(n13375), .A2(n13374), .ZN(n13401) );
  OAI22_X1 U15015 ( .A1(n13409), .A2(n13408), .B1(n13402), .B2(n13401), .ZN(
        n13376) );
  NAND2_X1 U15016 ( .A1(n13449), .A2(n13376), .ZN(n13403) );
  NAND2_X1 U15017 ( .A1(n14683), .A2(n9720), .ZN(n13380) );
  OR2_X1 U15018 ( .A1(n8004), .A2(n13377), .ZN(n13379) );
  INV_X1 U15019 ( .A(n14333), .ZN(n13385) );
  INV_X1 U15020 ( .A(n13381), .ZN(n13383) );
  INV_X1 U15021 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n13382) );
  NAND2_X1 U15022 ( .A1(n13383), .A2(n13382), .ZN(n13384) );
  NAND2_X1 U15023 ( .A1(n9789), .A2(n14371), .ZN(n13390) );
  NAND2_X1 U15024 ( .A1(n9742), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n13389) );
  NAND2_X1 U15025 ( .A1(n13386), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n13388) );
  NAND2_X1 U15026 ( .A1(n13368), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n13387) );
  NAND4_X1 U15027 ( .A1(n13390), .A2(n13389), .A3(n13388), .A4(n13387), .ZN(
        n14363) );
  AND2_X1 U15028 ( .A1(n14363), .A2(n13411), .ZN(n13391) );
  AOI21_X1 U15029 ( .B1(n14569), .B2(n13392), .A(n13391), .ZN(n13398) );
  NAND2_X1 U15030 ( .A1(n14569), .A2(n13360), .ZN(n13394) );
  NAND2_X1 U15031 ( .A1(n13392), .A2(n14363), .ZN(n13393) );
  NAND2_X1 U15032 ( .A1(n13394), .A2(n13393), .ZN(n13397) );
  NAND2_X1 U15033 ( .A1(n13398), .A2(n13397), .ZN(n13395) );
  AOI21_X1 U15034 ( .B1(n13406), .B2(n13405), .A(n13407), .ZN(n13396) );
  INV_X1 U15035 ( .A(n13397), .ZN(n13400) );
  INV_X1 U15036 ( .A(n13398), .ZN(n13399) );
  AOI22_X1 U15037 ( .A1(n13402), .A2(n13401), .B1(n13400), .B2(n13399), .ZN(
        n13404) );
  INV_X1 U15038 ( .A(n13410), .ZN(n13412) );
  NOR2_X1 U15039 ( .A1(n13412), .A2(n13411), .ZN(n13415) );
  INV_X1 U15040 ( .A(n14316), .ZN(n13413) );
  NOR2_X1 U15041 ( .A1(n13413), .A2(n13341), .ZN(n13414) );
  MUX2_X1 U15042 ( .A(n13415), .B(n13414), .S(n14641), .Z(n13416) );
  INV_X1 U15043 ( .A(n14363), .ZN(n14152) );
  NAND2_X1 U15044 ( .A1(n14569), .A2(n14152), .ZN(n13419) );
  NAND2_X1 U15045 ( .A1(n14357), .A2(n13419), .ZN(n14368) );
  XNOR2_X1 U15046 ( .A(n14574), .B(n14180), .ZN(n14384) );
  XOR2_X1 U15047 ( .A(n14354), .B(n14412), .Z(n14407) );
  XNOR2_X1 U15048 ( .A(n14580), .B(n14330), .ZN(n14393) );
  XNOR2_X1 U15049 ( .A(n14599), .B(n14350), .ZN(n14464) );
  OR2_X1 U15050 ( .A1(n14603), .A2(n14487), .ZN(n14347) );
  NAND2_X1 U15051 ( .A1(n14603), .A2(n14487), .ZN(n14348) );
  NAND2_X1 U15052 ( .A1(n14347), .A2(n14348), .ZN(n14477) );
  NAND4_X1 U15053 ( .A1(n13423), .A2(n13422), .A3(n13421), .A4(n7424), .ZN(
        n13426) );
  NOR4_X1 U15054 ( .A1(n13427), .A2(n13426), .A3(n13425), .A4(n13424), .ZN(
        n13430) );
  NAND4_X1 U15055 ( .A1(n13431), .A2(n13430), .A3(n13429), .A4(n13428), .ZN(
        n13432) );
  NOR4_X1 U15056 ( .A1(n13435), .A2(n13434), .A3(n13433), .A4(n13432), .ZN(
        n13438) );
  NAND4_X1 U15057 ( .A1(n13439), .A2(n13438), .A3(n13437), .A4(n13436), .ZN(
        n13440) );
  NOR3_X1 U15058 ( .A1(n14477), .A2(n13441), .A3(n13440), .ZN(n13443) );
  XNOR2_X1 U15059 ( .A(n14609), .B(n14344), .ZN(n14484) );
  NAND4_X1 U15060 ( .A1(n13443), .A2(n14338), .A3(n13442), .A4(n14484), .ZN(
        n13444) );
  XNOR2_X1 U15061 ( .A(n14505), .B(n14524), .ZN(n14501) );
  XNOR2_X1 U15062 ( .A(n14536), .B(n14326), .ZN(n14526) );
  NOR4_X1 U15063 ( .A1(n14464), .A2(n13444), .A3(n14501), .A4(n14526), .ZN(
        n13445) );
  INV_X1 U15064 ( .A(n14353), .ZN(n14440) );
  XNOR2_X1 U15065 ( .A(n14427), .B(n14440), .ZN(n14420) );
  NAND4_X1 U15066 ( .A1(n14393), .A2(n13445), .A3(n14436), .A4(n14420), .ZN(
        n13446) );
  NOR4_X1 U15067 ( .A1(n14368), .A2(n14384), .A3(n14407), .A4(n13446), .ZN(
        n13448) );
  XNOR2_X1 U15068 ( .A(n14563), .B(n14250), .ZN(n14359) );
  XNOR2_X1 U15069 ( .A(n14310), .B(n14362), .ZN(n13447) );
  NAND4_X1 U15070 ( .A1(n13449), .A2(n13448), .A3(n14359), .A4(n13447), .ZN(
        n13450) );
  XNOR2_X1 U15071 ( .A(n13450), .B(n14301), .ZN(n13452) );
  NAND2_X1 U15072 ( .A1(n13452), .A2(n13451), .ZN(n13453) );
  AOI21_X1 U15073 ( .B1(n13454), .B2(n13091), .A(n13453), .ZN(n13456) );
  INV_X1 U15074 ( .A(n13460), .ZN(n13455) );
  INV_X1 U15075 ( .A(n13351), .ZN(n13457) );
  NAND4_X1 U15076 ( .A1(n15784), .A2(n13458), .A3(n13457), .A4(n14438), .ZN(
        n13459) );
  OAI211_X1 U15077 ( .C1(n13090), .C2(n13460), .A(n13459), .B(P2_B_REG_SCAN_IN), .ZN(n13461) );
  INV_X1 U15078 ( .A(SI_30_), .ZN(n13463) );
  OAI222_X1 U15079 ( .A1(P3_U3151), .A2(n13465), .B1(n14119), .B2(n13464), 
        .C1(n13463), .C2(n13462), .ZN(P3_U3265) );
  INV_X1 U15080 ( .A(n14042), .ZN(n13471) );
  INV_X1 U15081 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n13467) );
  OAI22_X1 U15082 ( .A1(n13775), .A2(n13600), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13467), .ZN(n13469) );
  NOR2_X1 U15083 ( .A1(n13776), .A2(n13575), .ZN(n13468) );
  AOI211_X1 U15084 ( .C1(n13781), .C2(n13568), .A(n13469), .B(n13468), .ZN(
        n13470) );
  AOI21_X1 U15085 ( .B1(n13473), .B2(n13472), .A(n7606), .ZN(n13481) );
  INV_X1 U15086 ( .A(n14097), .ZN(n13479) );
  INV_X1 U15087 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n13474) );
  NOR2_X1 U15088 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13474), .ZN(n15960) );
  NOR2_X1 U15089 ( .A1(n13475), .A2(n13600), .ZN(n13476) );
  AOI211_X1 U15090 ( .C1(n13602), .C2(n13944), .A(n15960), .B(n13476), .ZN(
        n13477) );
  OAI21_X1 U15091 ( .B1(n13950), .B2(n13604), .A(n13477), .ZN(n13478) );
  AOI21_X1 U15092 ( .B1(n13479), .B2(n13606), .A(n13478), .ZN(n13480) );
  OAI21_X1 U15093 ( .B1(n13481), .B2(n13608), .A(n13480), .ZN(P3_U3155) );
  INV_X1 U15094 ( .A(n13482), .ZN(n14065) );
  OAI21_X1 U15095 ( .B1(n13838), .B2(n13483), .A(n13539), .ZN(n13484) );
  NAND2_X1 U15096 ( .A1(n13484), .A2(n13587), .ZN(n13488) );
  AOI22_X1 U15097 ( .A1(n13611), .A2(n13589), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13485) );
  OAI21_X1 U15098 ( .B1(n8379), .B2(n13575), .A(n13485), .ZN(n13486) );
  AOI21_X1 U15099 ( .B1(n13827), .B2(n13568), .A(n13486), .ZN(n13487) );
  OAI211_X1 U15100 ( .C1(n14065), .C2(n13595), .A(n13488), .B(n13487), .ZN(
        P3_U3156) );
  OAI21_X1 U15101 ( .B1(n13491), .B2(n13490), .A(n13489), .ZN(n13492) );
  NAND2_X1 U15102 ( .A1(n13492), .A2(n13587), .ZN(n13496) );
  NOR2_X1 U15103 ( .A1(n13604), .A2(n13879), .ZN(n13494) );
  NAND2_X1 U15104 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13729)
         );
  OAI21_X1 U15105 ( .B1(n13575), .B2(n13847), .A(n13729), .ZN(n13493) );
  AOI211_X1 U15106 ( .C1(n13589), .C2(n13873), .A(n13494), .B(n13493), .ZN(
        n13495) );
  OAI211_X1 U15107 ( .C1(n13878), .C2(n13595), .A(n13496), .B(n13495), .ZN(
        P3_U3159) );
  INV_X1 U15108 ( .A(n13497), .ZN(n13499) );
  NOR2_X1 U15109 ( .A1(n13499), .A2(n13498), .ZN(n13500) );
  XNOR2_X1 U15110 ( .A(n13501), .B(n13500), .ZN(n13506) );
  AOI22_X1 U15111 ( .A1(n13874), .A2(n13589), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13503) );
  NAND2_X1 U15112 ( .A1(n13568), .A2(n13855), .ZN(n13502) );
  OAI211_X1 U15113 ( .C1(n13848), .C2(n13575), .A(n13503), .B(n13502), .ZN(
        n13504) );
  AOI21_X1 U15114 ( .B1(n14074), .B2(n13606), .A(n13504), .ZN(n13505) );
  OAI21_X1 U15115 ( .B1(n13506), .B2(n13608), .A(n13505), .ZN(P3_U3163) );
  NOR3_X1 U15116 ( .A1(n13541), .A2(n13508), .A3(n13507), .ZN(n13509) );
  OAI21_X1 U15117 ( .B1(n7493), .B2(n13509), .A(n13587), .ZN(n13513) );
  AOI22_X1 U15118 ( .A1(n13610), .A2(n13589), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13510) );
  OAI21_X1 U15119 ( .B1(n13775), .B2(n13575), .A(n13510), .ZN(n13511) );
  AOI21_X1 U15120 ( .B1(n13808), .B2(n13568), .A(n13511), .ZN(n13512) );
  OAI211_X1 U15121 ( .C1(n8038), .C2(n13595), .A(n13513), .B(n13512), .ZN(
        P3_U3165) );
  NAND2_X1 U15122 ( .A1(n13514), .A2(n13525), .ZN(n13517) );
  XNOR2_X1 U15123 ( .A(n13515), .B(n13519), .ZN(n13598) );
  OAI22_X1 U15124 ( .A1(n13598), .A2(n13597), .B1(n13519), .B2(n13515), .ZN(
        n13516) );
  NOR2_X1 U15125 ( .A1(n13516), .A2(n13517), .ZN(n13528) );
  AOI21_X1 U15126 ( .B1(n13517), .B2(n13516), .A(n13528), .ZN(n13524) );
  NOR2_X1 U15127 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13518), .ZN(n13652) );
  NOR2_X1 U15128 ( .A1(n13519), .A2(n13600), .ZN(n13520) );
  AOI211_X1 U15129 ( .C1(n13602), .C2(n13913), .A(n13652), .B(n13520), .ZN(
        n13521) );
  OAI21_X1 U15130 ( .B1(n8715), .B2(n13604), .A(n13521), .ZN(n13522) );
  AOI21_X1 U15131 ( .B1(n13606), .B2(n13918), .A(n13522), .ZN(n13523) );
  OAI21_X1 U15132 ( .B1(n13524), .B2(n13608), .A(n13523), .ZN(P3_U3166) );
  INV_X1 U15133 ( .A(n13525), .ZN(n13527) );
  NOR3_X1 U15134 ( .A1(n13528), .A2(n13527), .A3(n13526), .ZN(n13531) );
  INV_X1 U15135 ( .A(n13529), .ZN(n13530) );
  OAI21_X1 U15136 ( .B1(n13531), .B2(n13530), .A(n13587), .ZN(n13536) );
  NOR2_X1 U15137 ( .A1(n13604), .A2(n13903), .ZN(n13534) );
  NAND2_X1 U15138 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13679)
         );
  OAI21_X1 U15139 ( .B1(n13575), .B2(n13900), .A(n13679), .ZN(n13533) );
  AOI211_X1 U15140 ( .C1(n13589), .C2(n13928), .A(n13534), .B(n13533), .ZN(
        n13535) );
  OAI211_X1 U15141 ( .C1(n13595), .C2(n14089), .A(n13536), .B(n13535), .ZN(
        P3_U3168) );
  AND3_X1 U15142 ( .A1(n13539), .A2(n13538), .A3(n13537), .ZN(n13540) );
  OAI21_X1 U15143 ( .B1(n13541), .B2(n13540), .A(n13587), .ZN(n13547) );
  INV_X1 U15144 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n13542) );
  OAI22_X1 U15145 ( .A1(n13838), .A2(n13600), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13542), .ZN(n13545) );
  NOR2_X1 U15146 ( .A1(n13543), .A2(n13575), .ZN(n13544) );
  AOI211_X1 U15147 ( .C1(n13820), .C2(n13568), .A(n13545), .B(n13544), .ZN(
        n13546) );
  OAI211_X1 U15148 ( .C1(n8380), .C2(n13595), .A(n13547), .B(n13546), .ZN(
        P3_U3169) );
  XNOR2_X1 U15149 ( .A(n13548), .B(n13874), .ZN(n13549) );
  XNOR2_X1 U15150 ( .A(n13550), .B(n13549), .ZN(n13555) );
  AOI22_X1 U15151 ( .A1(n13602), .A2(n13862), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13552) );
  NAND2_X1 U15152 ( .A1(n13568), .A2(n13867), .ZN(n13551) );
  OAI211_X1 U15153 ( .C1(n13574), .C2(n13600), .A(n13552), .B(n13551), .ZN(
        n13553) );
  AOI21_X1 U15154 ( .B1(n14080), .B2(n13606), .A(n13553), .ZN(n13554) );
  OAI21_X1 U15155 ( .B1(n13555), .B2(n13608), .A(n13554), .ZN(P3_U3173) );
  AND2_X1 U15156 ( .A1(n13557), .A2(n13556), .ZN(n13560) );
  OAI211_X1 U15157 ( .C1(n13560), .C2(n13559), .A(n13587), .B(n13558), .ZN(
        n13565) );
  NOR2_X1 U15158 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15349), .ZN(n15955) );
  AOI21_X1 U15159 ( .B1(n13602), .B2(n13927), .A(n15955), .ZN(n13562) );
  NAND2_X1 U15160 ( .A1(n13589), .A2(n13612), .ZN(n13561) );
  OAI211_X1 U15161 ( .C1(n13964), .C2(n13604), .A(n13562), .B(n13561), .ZN(
        n13563) );
  INV_X1 U15162 ( .A(n13563), .ZN(n13564) );
  OAI211_X1 U15163 ( .C1(n13595), .C2(n14101), .A(n13565), .B(n13564), .ZN(
        P3_U3174) );
  AOI21_X1 U15164 ( .B1(n13611), .B2(n13567), .A(n13566), .ZN(n13573) );
  AOI22_X1 U15165 ( .A1(n13589), .A2(n13862), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13570) );
  NAND2_X1 U15166 ( .A1(n13568), .A2(n13843), .ZN(n13569) );
  OAI211_X1 U15167 ( .C1(n13838), .C2(n13575), .A(n13570), .B(n13569), .ZN(
        n13571) );
  AOI21_X1 U15168 ( .B1(n14068), .B2(n13606), .A(n13571), .ZN(n13572) );
  OAI21_X1 U15169 ( .B1(n13573), .B2(n13608), .A(n13572), .ZN(P3_U3175) );
  NAND2_X1 U15170 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13702)
         );
  OAI21_X1 U15171 ( .B1(n13575), .B2(n13574), .A(n13702), .ZN(n13576) );
  AOI21_X1 U15172 ( .B1(n13589), .B2(n13913), .A(n13576), .ZN(n13577) );
  OAI21_X1 U15173 ( .B1(n13604), .B2(n13889), .A(n13577), .ZN(n13582) );
  AOI211_X1 U15174 ( .C1(n13580), .C2(n13579), .A(n13608), .B(n13578), .ZN(
        n13581) );
  AOI211_X1 U15175 ( .C1(n13606), .C2(n14005), .A(n13582), .B(n13581), .ZN(
        n13583) );
  INV_X1 U15176 ( .A(n13583), .ZN(P3_U3178) );
  INV_X1 U15177 ( .A(n14048), .ZN(n13596) );
  OAI21_X1 U15178 ( .B1(n13586), .B2(n13585), .A(n13584), .ZN(n13588) );
  NAND2_X1 U15179 ( .A1(n13588), .A2(n13587), .ZN(n13594) );
  INV_X1 U15180 ( .A(n13792), .ZN(n13591) );
  AOI22_X1 U15181 ( .A1(n8037), .A2(n13589), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13590) );
  OAI21_X1 U15182 ( .B1(n13591), .B2(n13604), .A(n13590), .ZN(n13592) );
  AOI21_X1 U15183 ( .B1(n13602), .B2(n13787), .A(n13592), .ZN(n13593) );
  OAI211_X1 U15184 ( .C1(n13596), .C2(n13595), .A(n13594), .B(n13593), .ZN(
        P3_U3180) );
  XNOR2_X1 U15185 ( .A(n13598), .B(n13597), .ZN(n13609) );
  INV_X1 U15186 ( .A(n14017), .ZN(n13934) );
  INV_X1 U15187 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n13599) );
  NOR2_X1 U15188 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13599), .ZN(n15997) );
  NOR2_X1 U15189 ( .A1(n13958), .A2(n13600), .ZN(n13601) );
  AOI211_X1 U15190 ( .C1(n13602), .C2(n13928), .A(n15997), .B(n13601), .ZN(
        n13603) );
  OAI21_X1 U15191 ( .B1(n13931), .B2(n13604), .A(n13603), .ZN(n13605) );
  AOI21_X1 U15192 ( .B1(n13934), .B2(n13606), .A(n13605), .ZN(n13607) );
  OAI21_X1 U15193 ( .B1(n13609), .B2(n13608), .A(n13607), .ZN(P3_U3181) );
  MUX2_X1 U15194 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n13736), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U15195 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n13754), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U15196 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n13787), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15197 ( .A(n13801), .B(P3_DATAO_REG_26__SCAN_IN), .S(n13623), .Z(
        P3_U3517) );
  MUX2_X1 U15198 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n8037), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U15199 ( .A(n13610), .B(P3_DATAO_REG_24__SCAN_IN), .S(n13623), .Z(
        P3_U3515) );
  MUX2_X1 U15200 ( .A(n13815), .B(P3_DATAO_REG_23__SCAN_IN), .S(n13623), .Z(
        P3_U3514) );
  MUX2_X1 U15201 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n13611), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15202 ( .A(n13862), .B(P3_DATAO_REG_21__SCAN_IN), .S(n13623), .Z(
        P3_U3512) );
  MUX2_X1 U15203 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13874), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15204 ( .A(n13887), .B(P3_DATAO_REG_19__SCAN_IN), .S(n13623), .Z(
        P3_U3510) );
  MUX2_X1 U15205 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13873), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15206 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13913), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U15207 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13928), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U15208 ( .A(n13927), .B(P3_DATAO_REG_14__SCAN_IN), .S(n13623), .Z(
        P3_U3505) );
  MUX2_X1 U15209 ( .A(n13942), .B(P3_DATAO_REG_13__SCAN_IN), .S(n13623), .Z(
        P3_U3504) );
  MUX2_X1 U15210 ( .A(n13612), .B(P3_DATAO_REG_12__SCAN_IN), .S(n13623), .Z(
        P3_U3503) );
  MUX2_X1 U15211 ( .A(n13613), .B(P3_DATAO_REG_11__SCAN_IN), .S(n13623), .Z(
        P3_U3502) );
  MUX2_X1 U15212 ( .A(n13614), .B(P3_DATAO_REG_10__SCAN_IN), .S(n13623), .Z(
        P3_U3501) );
  MUX2_X1 U15213 ( .A(n13615), .B(P3_DATAO_REG_9__SCAN_IN), .S(n13623), .Z(
        P3_U3500) );
  MUX2_X1 U15214 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n13616), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U15215 ( .A(n13617), .B(P3_DATAO_REG_7__SCAN_IN), .S(n13623), .Z(
        P3_U3498) );
  MUX2_X1 U15216 ( .A(n13618), .B(P3_DATAO_REG_6__SCAN_IN), .S(n13623), .Z(
        P3_U3497) );
  MUX2_X1 U15217 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n13619), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U15218 ( .A(n13620), .B(P3_DATAO_REG_4__SCAN_IN), .S(n13623), .Z(
        P3_U3495) );
  MUX2_X1 U15219 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n13621), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15220 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n13622), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15221 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n7428), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15222 ( .A(n13624), .B(P3_DATAO_REG_0__SCAN_IN), .S(n13623), .Z(
        P3_U3491) );
  NAND2_X1 U15223 ( .A1(n15926), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n13638) );
  OAI21_X1 U15224 ( .B1(n15926), .B2(P3_REG2_REG_12__SCAN_IN), .A(n13638), 
        .ZN(n15922) );
  INV_X1 U15225 ( .A(n15921), .ZN(n13626) );
  AND2_X1 U15226 ( .A1(n15944), .A2(n13627), .ZN(n13628) );
  INV_X1 U15227 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n15942) );
  NOR2_X1 U15228 ( .A1(n15942), .A2(n15941), .ZN(n15940) );
  NAND2_X1 U15229 ( .A1(P3_REG2_REG_14__SCAN_IN), .A2(n15958), .ZN(n13629) );
  OAI21_X1 U15230 ( .B1(P3_REG2_REG_14__SCAN_IN), .B2(n15958), .A(n13629), 
        .ZN(n15967) );
  NOR2_X1 U15231 ( .A1(n15968), .A2(n15967), .ZN(n15969) );
  NOR2_X1 U15232 ( .A1(n13662), .A2(n13630), .ZN(n13631) );
  NAND2_X1 U15233 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n13676), .ZN(n13632) );
  OAI21_X1 U15234 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n13676), .A(n13632), 
        .ZN(n13633) );
  AOI21_X1 U15235 ( .B1(n7504), .B2(n13633), .A(n13675), .ZN(n13672) );
  INV_X1 U15236 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n14025) );
  MUX2_X1 U15237 ( .A(n13951), .B(n14025), .S(n8634), .Z(n13642) );
  OR2_X1 U15238 ( .A1(n13634), .A2(n13642), .ZN(n13643) );
  MUX2_X1 U15239 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n8634), .Z(n13640) );
  INV_X1 U15240 ( .A(n13640), .ZN(n13641) );
  NAND2_X1 U15241 ( .A1(n13635), .A2(n13655), .ZN(n13637) );
  NAND2_X1 U15242 ( .A1(n13637), .A2(n13636), .ZN(n15933) );
  NAND2_X1 U15243 ( .A1(n15926), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n13657) );
  OAI21_X1 U15244 ( .B1(n15926), .B2(P3_REG1_REG_12__SCAN_IN), .A(n13657), 
        .ZN(n15924) );
  MUX2_X1 U15245 ( .A(n15922), .B(n15924), .S(n8634), .Z(n15934) );
  OR2_X2 U15246 ( .A1(n15933), .A2(n15934), .ZN(n15935) );
  MUX2_X1 U15247 ( .A(n13638), .B(n13657), .S(n8634), .Z(n13639) );
  NAND2_X1 U15248 ( .A1(n15935), .A2(n13639), .ZN(n15949) );
  XNOR2_X1 U15249 ( .A(n13640), .B(n15944), .ZN(n15950) );
  NOR2_X1 U15250 ( .A1(n15949), .A2(n15950), .ZN(n15948) );
  AOI21_X1 U15251 ( .B1(n13659), .B2(n13641), .A(n15948), .ZN(n15973) );
  XNOR2_X1 U15252 ( .A(n13642), .B(n15958), .ZN(n15972) );
  NOR2_X1 U15253 ( .A1(n15983), .A2(n13644), .ZN(n13645) );
  MUX2_X1 U15254 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n8634), .Z(n15989) );
  XNOR2_X1 U15255 ( .A(n15983), .B(n13644), .ZN(n15990) );
  NOR2_X1 U15256 ( .A1(n13645), .A2(n15988), .ZN(n13681) );
  MUX2_X1 U15257 ( .A(n13916), .B(n13646), .S(n8634), .Z(n13648) );
  INV_X1 U15258 ( .A(n13676), .ZN(n13647) );
  NAND2_X1 U15259 ( .A1(n13648), .A2(n13647), .ZN(n13680) );
  MUX2_X1 U15260 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n8634), .Z(n13649) );
  AND2_X1 U15261 ( .A1(n13649), .A2(n13676), .ZN(n13682) );
  INV_X1 U15262 ( .A(n13682), .ZN(n13650) );
  NAND2_X1 U15263 ( .A1(n13680), .A2(n13650), .ZN(n13651) );
  XNOR2_X1 U15264 ( .A(n13681), .B(n13651), .ZN(n13670) );
  AOI21_X1 U15265 ( .B1(n15961), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n13652), 
        .ZN(n13653) );
  OAI21_X1 U15266 ( .B1(n15984), .B2(n13676), .A(n13653), .ZN(n13669) );
  AND2_X1 U15267 ( .A1(n15944), .A2(n13658), .ZN(n13660) );
  INV_X1 U15268 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n15947) );
  NOR2_X1 U15269 ( .A1(n13660), .A2(n15945), .ZN(n15964) );
  NAND2_X1 U15270 ( .A1(P3_REG1_REG_14__SCAN_IN), .A2(n15958), .ZN(n13661) );
  OAI21_X1 U15271 ( .B1(n15958), .B2(P3_REG1_REG_14__SCAN_IN), .A(n13661), 
        .ZN(n15963) );
  NOR2_X1 U15272 ( .A1(n15964), .A2(n15963), .ZN(n15962) );
  NAND2_X1 U15273 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n13676), .ZN(n13664) );
  OAI21_X1 U15274 ( .B1(P3_REG1_REG_16__SCAN_IN), .B2(n13676), .A(n13664), 
        .ZN(n13665) );
  AOI21_X1 U15275 ( .B1(n13666), .B2(n13665), .A(n13673), .ZN(n13667) );
  NOR2_X1 U15276 ( .A1(n13667), .A2(n15993), .ZN(n13668) );
  AOI211_X1 U15277 ( .C1(n15970), .C2(n13670), .A(n13669), .B(n13668), .ZN(
        n13671) );
  OAI21_X1 U15278 ( .B1(n13672), .B2(n15999), .A(n13671), .ZN(P3_U3198) );
  XNOR2_X1 U15279 ( .A(n13705), .B(n13706), .ZN(n13674) );
  AOI21_X1 U15280 ( .B1(n14011), .B2(n13674), .A(n13707), .ZN(n13691) );
  NOR2_X1 U15281 ( .A1(n8016), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n13678) );
  OAI21_X1 U15282 ( .B1(n13678), .B2(n13692), .A(n15966), .ZN(n13690) );
  INV_X1 U15283 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n15903) );
  OAI21_X1 U15284 ( .B1(n15982), .B2(n15903), .A(n13679), .ZN(n13688) );
  OAI21_X1 U15285 ( .B1(n13682), .B2(n13681), .A(n13680), .ZN(n13686) );
  MUX2_X1 U15286 ( .A(n13904), .B(n14011), .S(n8634), .Z(n13683) );
  NOR2_X1 U15287 ( .A1(n13683), .A2(n13706), .ZN(n13697) );
  AOI21_X1 U15288 ( .B1(n13706), .B2(n13683), .A(n13697), .ZN(n13684) );
  INV_X1 U15289 ( .A(n13684), .ZN(n13685) );
  NOR2_X1 U15290 ( .A1(n13686), .A2(n13685), .ZN(n13696) );
  AOI211_X1 U15291 ( .C1(n13686), .C2(n13685), .A(n13696), .B(n15991), .ZN(
        n13687) );
  AOI211_X1 U15292 ( .C1(n13713), .C2(n13706), .A(n13688), .B(n13687), .ZN(
        n13689) );
  OAI211_X1 U15293 ( .C1(n13691), .C2(n15993), .A(n13690), .B(n13689), .ZN(
        P3_U3199) );
  NAND2_X1 U15294 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n13719), .ZN(n13693) );
  OAI21_X1 U15295 ( .B1(P3_REG2_REG_18__SCAN_IN), .B2(n13719), .A(n13693), 
        .ZN(n13694) );
  AOI21_X1 U15296 ( .B1(n13695), .B2(n13694), .A(n13718), .ZN(n13714) );
  NAND2_X1 U15297 ( .A1(n15961), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n13704) );
  INV_X1 U15298 ( .A(n13720), .ZN(n13698) );
  MUX2_X1 U15299 ( .A(n13890), .B(n13709), .S(n8634), .Z(n13699) );
  NAND2_X1 U15300 ( .A1(n13699), .A2(n13700), .ZN(n13723) );
  OAI21_X1 U15301 ( .B1(n13700), .B2(n13699), .A(n13723), .ZN(n13701) );
  NAND2_X1 U15302 ( .A1(n15970), .A2(n13701), .ZN(n13703) );
  NAND3_X1 U15303 ( .A1(n13704), .A2(n13703), .A3(n13702), .ZN(n13712) );
  NOR2_X1 U15304 ( .A1(n13706), .A2(n13705), .ZN(n13708) );
  AOI22_X1 U15305 ( .A1(n13721), .A2(P3_REG1_REG_18__SCAN_IN), .B1(n13709), 
        .B2(n13719), .ZN(n13710) );
  XNOR2_X1 U15306 ( .A(n13733), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13724) );
  XNOR2_X1 U15307 ( .A(n13716), .B(n13724), .ZN(n13717) );
  NAND2_X1 U15308 ( .A1(n13717), .A2(n15931), .ZN(n13732) );
  MUX2_X1 U15309 ( .A(n13880), .B(P3_REG2_REG_19__SCAN_IN), .S(n13733), .Z(
        n13725) );
  NAND2_X1 U15310 ( .A1(n13721), .A2(n13720), .ZN(n13722) );
  NAND2_X1 U15311 ( .A1(n13723), .A2(n13722), .ZN(n13727) );
  MUX2_X1 U15312 ( .A(n13725), .B(n13724), .S(n8634), .Z(n13726) );
  XNOR2_X1 U15313 ( .A(n13727), .B(n13726), .ZN(n13728) );
  OAI21_X1 U15314 ( .B1(n15982), .B2(n8402), .A(n13729), .ZN(n13730) );
  AOI21_X1 U15315 ( .B1(n13868), .B2(n13744), .A(n16123), .ZN(n13737) );
  INV_X1 U15316 ( .A(n13734), .ZN(n13735) );
  NAND2_X1 U15317 ( .A1(n13736), .A2(n13735), .ZN(n16406) );
  NAND2_X1 U15318 ( .A1(n13737), .A2(n16406), .ZN(n13740) );
  OAI21_X1 U15319 ( .B1(P3_REG2_REG_31__SCAN_IN), .B2(n16121), .A(n13740), 
        .ZN(n13738) );
  OAI21_X1 U15320 ( .B1(n13739), .B2(n13963), .A(n13738), .ZN(P3_U3202) );
  INV_X1 U15321 ( .A(n16409), .ZN(n13742) );
  OAI21_X1 U15322 ( .B1(P3_REG2_REG_30__SCAN_IN), .B2(n16121), .A(n13740), 
        .ZN(n13741) );
  OAI21_X1 U15323 ( .B1(n13742), .B2(n13963), .A(n13741), .ZN(P3_U3203) );
  INV_X1 U15324 ( .A(n13743), .ZN(n13750) );
  AOI22_X1 U15325 ( .A1(n13744), .A2(n13868), .B1(P3_REG2_REG_29__SCAN_IN), 
        .B2(n16123), .ZN(n13745) );
  OAI21_X1 U15326 ( .B1(n13746), .B2(n13963), .A(n13745), .ZN(n13747) );
  AOI21_X1 U15327 ( .B1(n13748), .B2(n13967), .A(n13747), .ZN(n13749) );
  OAI21_X1 U15328 ( .B1(n13750), .B2(n16123), .A(n13749), .ZN(P3_U3204) );
  AOI22_X1 U15329 ( .A1(n13754), .A2(n13943), .B1(n13941), .B2(n13787), .ZN(
        n13755) );
  OR2_X1 U15330 ( .A1(n13758), .A2(n13757), .ZN(n13759) );
  NAND2_X1 U15331 ( .A1(n13760), .A2(n13759), .ZN(n13970) );
  AOI22_X1 U15332 ( .A1(n13761), .A2(n13868), .B1(n16123), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n13762) );
  OAI21_X1 U15333 ( .B1(n14039), .B2(n13963), .A(n13762), .ZN(n13763) );
  AOI21_X1 U15334 ( .B1(n13970), .B2(n13967), .A(n13763), .ZN(n13764) );
  OAI21_X1 U15335 ( .B1(n13972), .B2(n16123), .A(n13764), .ZN(P3_U3205) );
  NAND2_X1 U15336 ( .A1(n13766), .A2(n13765), .ZN(n13767) );
  NAND2_X1 U15337 ( .A1(n13768), .A2(n13767), .ZN(n13975) );
  INV_X1 U15338 ( .A(n13975), .ZN(n14045) );
  NAND2_X1 U15339 ( .A1(n13772), .A2(n13771), .ZN(n13773) );
  NAND2_X1 U15340 ( .A1(n13770), .A2(n13773), .ZN(n13774) );
  NAND2_X1 U15341 ( .A1(n13774), .A2(n16054), .ZN(n13779) );
  OAI22_X1 U15342 ( .A1(n13776), .A2(n16101), .B1(n13775), .B2(n16103), .ZN(
        n13777) );
  AOI21_X1 U15343 ( .B1(n13975), .B2(n16229), .A(n13777), .ZN(n13778) );
  MUX2_X1 U15344 ( .A(n14041), .B(n13780), .S(n16123), .Z(n13783) );
  AOI22_X1 U15345 ( .A1(n14042), .A2(n13933), .B1(n13868), .B2(n13781), .ZN(
        n13782) );
  OAI211_X1 U15346 ( .C1(n14045), .C2(n13871), .A(n13783), .B(n13782), .ZN(
        P3_U3206) );
  XOR2_X1 U15347 ( .A(n13786), .B(n13785), .Z(n13790) );
  AOI22_X1 U15348 ( .A1(n13787), .A2(n13943), .B1(n13941), .B2(n8037), .ZN(
        n13788) );
  OAI21_X1 U15349 ( .B1(n14051), .B2(n16178), .A(n13788), .ZN(n13789) );
  AOI21_X1 U15350 ( .B1(n13790), .B2(n16054), .A(n13789), .ZN(n14047) );
  MUX2_X1 U15351 ( .A(n14047), .B(n13791), .S(n16123), .Z(n13794) );
  AOI22_X1 U15352 ( .A1(n14048), .A2(n13933), .B1(n13868), .B2(n13792), .ZN(
        n13793) );
  OAI211_X1 U15353 ( .C1(n14051), .C2(n13871), .A(n13794), .B(n13793), .ZN(
        P3_U3207) );
  XNOR2_X1 U15354 ( .A(n13796), .B(n13795), .ZN(n13804) );
  INV_X1 U15355 ( .A(n13804), .ZN(n14053) );
  NAND2_X1 U15356 ( .A1(n13798), .A2(n13797), .ZN(n13799) );
  NAND3_X1 U15357 ( .A1(n13800), .A2(n16054), .A3(n13799), .ZN(n13806) );
  NAND2_X1 U15358 ( .A1(n13801), .A2(n13943), .ZN(n13802) );
  OAI21_X1 U15359 ( .B1(n8379), .B2(n16103), .A(n13802), .ZN(n13803) );
  AOI21_X1 U15360 ( .B1(n13804), .B2(n16229), .A(n13803), .ZN(n13805) );
  NAND2_X1 U15361 ( .A1(n13806), .A2(n13805), .ZN(n14052) );
  MUX2_X1 U15362 ( .A(n14052), .B(P3_REG2_REG_25__SCAN_IN), .S(n16123), .Z(
        n13807) );
  INV_X1 U15363 ( .A(n13807), .ZN(n13811) );
  AOI22_X1 U15364 ( .A1(n13809), .A2(n13933), .B1(n13868), .B2(n13808), .ZN(
        n13810) );
  OAI211_X1 U15365 ( .C1(n14053), .C2(n13871), .A(n13811), .B(n13810), .ZN(
        P3_U3208) );
  XNOR2_X1 U15366 ( .A(n13812), .B(n13813), .ZN(n14061) );
  XNOR2_X1 U15367 ( .A(n13814), .B(n13813), .ZN(n13818) );
  AOI22_X1 U15368 ( .A1(n8037), .A2(n13943), .B1(n13941), .B2(n13815), .ZN(
        n13816) );
  OAI21_X1 U15369 ( .B1(n14061), .B2(n16178), .A(n13816), .ZN(n13817) );
  AOI21_X1 U15370 ( .B1(n13818), .B2(n16054), .A(n13817), .ZN(n14057) );
  MUX2_X1 U15371 ( .A(n14057), .B(n13819), .S(n16123), .Z(n13822) );
  AOI22_X1 U15372 ( .A1(n14058), .A2(n13933), .B1(n13868), .B2(n13820), .ZN(
        n13821) );
  OAI211_X1 U15373 ( .C1(n14061), .C2(n13871), .A(n13822), .B(n13821), .ZN(
        P3_U3209) );
  XNOR2_X1 U15374 ( .A(n13823), .B(n13825), .ZN(n13824) );
  OAI222_X1 U15375 ( .A1(n16101), .A2(n8379), .B1(n16103), .B2(n13848), .C1(
        n13824), .C2(n16107), .ZN(n13986) );
  INV_X1 U15376 ( .A(n13986), .ZN(n13831) );
  XNOR2_X1 U15377 ( .A(n13826), .B(n13825), .ZN(n13987) );
  AOI22_X1 U15378 ( .A1(n16123), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n13827), 
        .B2(n13868), .ZN(n13828) );
  OAI21_X1 U15379 ( .B1(n14065), .B2(n13963), .A(n13828), .ZN(n13829) );
  AOI21_X1 U15380 ( .B1(n13987), .B2(n13967), .A(n13829), .ZN(n13830) );
  OAI21_X1 U15381 ( .B1(n13831), .B2(n16123), .A(n13830), .ZN(P3_U3210) );
  INV_X1 U15382 ( .A(n13834), .ZN(n13832) );
  XNOR2_X1 U15383 ( .A(n13833), .B(n13832), .ZN(n13991) );
  INV_X1 U15384 ( .A(n13991), .ZN(n14071) );
  XNOR2_X1 U15385 ( .A(n13835), .B(n13834), .ZN(n13836) );
  NAND2_X1 U15386 ( .A1(n13836), .A2(n16054), .ZN(n13841) );
  OAI22_X1 U15387 ( .A1(n13838), .A2(n16101), .B1(n13837), .B2(n16103), .ZN(
        n13839) );
  AOI21_X1 U15388 ( .B1(n13991), .B2(n16229), .A(n13839), .ZN(n13840) );
  MUX2_X1 U15389 ( .A(n14066), .B(n13842), .S(n16123), .Z(n13845) );
  AOI22_X1 U15390 ( .A1(n14068), .A2(n13933), .B1(n13868), .B2(n13843), .ZN(
        n13844) );
  OAI211_X1 U15391 ( .C1(n14071), .C2(n13871), .A(n13845), .B(n13844), .ZN(
        P3_U3211) );
  XNOR2_X1 U15392 ( .A(n13846), .B(n13850), .ZN(n13995) );
  INV_X1 U15393 ( .A(n13995), .ZN(n14077) );
  INV_X1 U15394 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n13854) );
  OAI22_X1 U15395 ( .A1(n13848), .A2(n16101), .B1(n13847), .B2(n16103), .ZN(
        n13853) );
  XOR2_X1 U15396 ( .A(n13850), .B(n13849), .Z(n13851) );
  NOR2_X1 U15397 ( .A1(n13851), .A2(n16107), .ZN(n13852) );
  AOI211_X1 U15398 ( .C1(n13995), .C2(n16229), .A(n13853), .B(n13852), .ZN(
        n14072) );
  MUX2_X1 U15399 ( .A(n13854), .B(n14072), .S(n16121), .Z(n13857) );
  AOI22_X1 U15400 ( .A1(n14074), .A2(n13933), .B1(n13868), .B2(n13855), .ZN(
        n13856) );
  OAI211_X1 U15401 ( .C1(n14077), .C2(n13871), .A(n13857), .B(n13856), .ZN(
        P3_U3212) );
  XNOR2_X1 U15402 ( .A(n13859), .B(n13858), .ZN(n14083) );
  XNOR2_X1 U15403 ( .A(n13861), .B(n13860), .ZN(n13865) );
  AOI22_X1 U15404 ( .A1(n13862), .A2(n13943), .B1(n13887), .B2(n13941), .ZN(
        n13863) );
  OAI21_X1 U15405 ( .B1(n14083), .B2(n16178), .A(n13863), .ZN(n13864) );
  AOI21_X1 U15406 ( .B1(n13865), .B2(n16054), .A(n13864), .ZN(n14078) );
  MUX2_X1 U15407 ( .A(n13866), .B(n14078), .S(n16121), .Z(n13870) );
  AOI22_X1 U15408 ( .A1(n14080), .A2(n13933), .B1(n13868), .B2(n13867), .ZN(
        n13869) );
  OAI211_X1 U15409 ( .C1(n14083), .C2(n13871), .A(n13870), .B(n13869), .ZN(
        P3_U3213) );
  XOR2_X1 U15410 ( .A(n13872), .B(n13876), .Z(n13875) );
  AOI222_X1 U15411 ( .A1(n16054), .A2(n13875), .B1(n13874), .B2(n13943), .C1(
        n13873), .C2(n13941), .ZN(n14004) );
  XNOR2_X1 U15412 ( .A(n13877), .B(n13876), .ZN(n14002) );
  NOR2_X1 U15413 ( .A1(n13878), .A2(n13963), .ZN(n13882) );
  OAI22_X1 U15414 ( .A1(n16121), .A2(n13880), .B1(n13879), .B2(n16113), .ZN(
        n13881) );
  AOI211_X1 U15415 ( .C1(n14002), .C2(n13967), .A(n13882), .B(n13881), .ZN(
        n13883) );
  OAI21_X1 U15416 ( .B1(n14004), .B2(n16123), .A(n13883), .ZN(P3_U3214) );
  OAI21_X1 U15417 ( .B1(n13886), .B2(n13885), .A(n13884), .ZN(n13888) );
  AOI222_X1 U15418 ( .A1(n16054), .A2(n13888), .B1(n13887), .B2(n13943), .C1(
        n13913), .C2(n13941), .ZN(n14008) );
  OAI22_X1 U15419 ( .A1(n16121), .A2(n13890), .B1(n13889), .B2(n16113), .ZN(
        n13891) );
  AOI21_X1 U15420 ( .B1(n14005), .B2(n13933), .A(n13891), .ZN(n13896) );
  OAI21_X1 U15421 ( .B1(n13894), .B2(n13893), .A(n13892), .ZN(n14006) );
  NAND2_X1 U15422 ( .A1(n14006), .A2(n13967), .ZN(n13895) );
  OAI211_X1 U15423 ( .C1(n14008), .C2(n16123), .A(n13896), .B(n13895), .ZN(
        P3_U3215) );
  XNOR2_X1 U15424 ( .A(n13897), .B(n13901), .ZN(n13898) );
  OAI222_X1 U15425 ( .A1(n16101), .A2(n13900), .B1(n16103), .B2(n13899), .C1(
        n16107), .C2(n13898), .ZN(n14009) );
  INV_X1 U15426 ( .A(n14009), .ZN(n13908) );
  XNOR2_X1 U15427 ( .A(n13902), .B(n13901), .ZN(n14010) );
  NOR2_X1 U15428 ( .A1(n14089), .A2(n13963), .ZN(n13906) );
  OAI22_X1 U15429 ( .A1(n16121), .A2(n13904), .B1(n13903), .B2(n16113), .ZN(
        n13905) );
  AOI211_X1 U15430 ( .C1(n14010), .C2(n13967), .A(n13906), .B(n13905), .ZN(
        n13907) );
  OAI21_X1 U15431 ( .B1(n13908), .B2(n16123), .A(n13907), .ZN(P3_U3216) );
  XNOR2_X1 U15432 ( .A(n13909), .B(n13910), .ZN(n14014) );
  XNOR2_X1 U15433 ( .A(n13911), .B(n13910), .ZN(n13912) );
  NAND2_X1 U15434 ( .A1(n13912), .A2(n16054), .ZN(n13915) );
  AOI22_X1 U15435 ( .A1(n13913), .A2(n13943), .B1(n13941), .B2(n13944), .ZN(
        n13914) );
  NAND2_X1 U15436 ( .A1(n13915), .A2(n13914), .ZN(n14016) );
  NAND2_X1 U15437 ( .A1(n14016), .A2(n16121), .ZN(n13920) );
  OAI22_X1 U15438 ( .A1(n16121), .A2(n13916), .B1(n8715), .B2(n16113), .ZN(
        n13917) );
  AOI21_X1 U15439 ( .B1(n13918), .B2(n13933), .A(n13917), .ZN(n13919) );
  OAI211_X1 U15440 ( .C1(n14014), .C2(n13937), .A(n13920), .B(n13919), .ZN(
        P3_U3217) );
  XNOR2_X1 U15441 ( .A(n13921), .B(n9244), .ZN(n14019) );
  NAND2_X1 U15442 ( .A1(n13923), .A2(n13922), .ZN(n13924) );
  NAND2_X1 U15443 ( .A1(n13925), .A2(n13924), .ZN(n13926) );
  NAND2_X1 U15444 ( .A1(n13926), .A2(n16054), .ZN(n13930) );
  AOI22_X1 U15445 ( .A1(n13928), .A2(n13943), .B1(n13941), .B2(n13927), .ZN(
        n13929) );
  NAND2_X1 U15446 ( .A1(n13930), .A2(n13929), .ZN(n14021) );
  NAND2_X1 U15447 ( .A1(n14021), .A2(n16121), .ZN(n13936) );
  OAI22_X1 U15448 ( .A1(n16121), .A2(n15980), .B1(n13931), .B2(n16113), .ZN(
        n13932) );
  AOI21_X1 U15449 ( .B1(n13934), .B2(n13933), .A(n13932), .ZN(n13935) );
  OAI211_X1 U15450 ( .C1(n14019), .C2(n13937), .A(n13936), .B(n13935), .ZN(
        P3_U3218) );
  OAI211_X1 U15451 ( .C1(n13940), .C2(n13939), .A(n16054), .B(n13938), .ZN(
        n13946) );
  AOI22_X1 U15452 ( .A1(n13944), .A2(n13943), .B1(n13942), .B2(n13941), .ZN(
        n13945) );
  NAND2_X1 U15453 ( .A1(n13946), .A2(n13945), .ZN(n14023) );
  INV_X1 U15454 ( .A(n14023), .ZN(n13955) );
  NOR2_X1 U15455 ( .A1(n13962), .A2(n13961), .ZN(n13960) );
  NOR2_X1 U15456 ( .A1(n13960), .A2(n13947), .ZN(n13949) );
  XNOR2_X1 U15457 ( .A(n13949), .B(n13948), .ZN(n14024) );
  NOR2_X1 U15458 ( .A1(n14097), .A2(n13963), .ZN(n13953) );
  OAI22_X1 U15459 ( .A1(n16121), .A2(n13951), .B1(n13950), .B2(n16113), .ZN(
        n13952) );
  AOI211_X1 U15460 ( .C1(n14024), .C2(n13967), .A(n13953), .B(n13952), .ZN(
        n13954) );
  OAI21_X1 U15461 ( .B1(n13955), .B2(n16123), .A(n13954), .ZN(P3_U3219) );
  XOR2_X1 U15462 ( .A(n13956), .B(n13961), .Z(n13957) );
  OAI222_X1 U15463 ( .A1(n16103), .A2(n13959), .B1(n16101), .B2(n13958), .C1(
        n16107), .C2(n13957), .ZN(n14027) );
  INV_X1 U15464 ( .A(n14027), .ZN(n13969) );
  AOI21_X1 U15465 ( .B1(n13962), .B2(n13961), .A(n13960), .ZN(n14028) );
  NOR2_X1 U15466 ( .A1(n14101), .A2(n13963), .ZN(n13966) );
  OAI22_X1 U15467 ( .A1(n16121), .A2(n15942), .B1(n13964), .B2(n16113), .ZN(
        n13965) );
  AOI211_X1 U15468 ( .C1(n14028), .C2(n13967), .A(n13966), .B(n13965), .ZN(
        n13968) );
  OAI21_X1 U15469 ( .B1(n13969), .B2(n16123), .A(n13968), .ZN(P3_U3220) );
  NAND2_X1 U15470 ( .A1(n13970), .A2(n16316), .ZN(n13971) );
  OAI21_X1 U15471 ( .B1(n14039), .B2(n14030), .A(n13973), .ZN(P3_U3487) );
  INV_X1 U15472 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13974) );
  MUX2_X1 U15473 ( .A(n13974), .B(n14041), .S(n16407), .Z(n13977) );
  AOI22_X1 U15474 ( .A1(n13975), .A2(n16259), .B1(n9313), .B2(n14042), .ZN(
        n13976) );
  NAND2_X1 U15475 ( .A1(n13977), .A2(n13976), .ZN(P3_U3486) );
  INV_X1 U15476 ( .A(n16259), .ZN(n14037) );
  INV_X1 U15477 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13978) );
  MUX2_X1 U15478 ( .A(n14047), .B(n13978), .S(n9309), .Z(n13980) );
  NAND2_X1 U15479 ( .A1(n14048), .A2(n9313), .ZN(n13979) );
  OAI211_X1 U15480 ( .C1(n14051), .C2(n14037), .A(n13980), .B(n13979), .ZN(
        P3_U3485) );
  MUX2_X1 U15481 ( .A(n14052), .B(P3_REG1_REG_25__SCAN_IN), .S(n9309), .Z(
        n13982) );
  OAI22_X1 U15482 ( .A1(n14053), .A2(n14037), .B1(n8038), .B2(n14030), .ZN(
        n13981) );
  OR2_X1 U15483 ( .A1(n13982), .A2(n13981), .ZN(P3_U3484) );
  INV_X1 U15484 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13983) );
  MUX2_X1 U15485 ( .A(n14057), .B(n13983), .S(n9309), .Z(n13985) );
  NAND2_X1 U15486 ( .A1(n14058), .A2(n9313), .ZN(n13984) );
  OAI211_X1 U15487 ( .C1(n14061), .C2(n14037), .A(n13985), .B(n13984), .ZN(
        P3_U3483) );
  INV_X1 U15488 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13988) );
  AOI21_X1 U15489 ( .B1(n16316), .B2(n13987), .A(n13986), .ZN(n14062) );
  MUX2_X1 U15490 ( .A(n13988), .B(n14062), .S(n16407), .Z(n13989) );
  OAI21_X1 U15491 ( .B1(n14065), .B2(n14030), .A(n13989), .ZN(P3_U3482) );
  INV_X1 U15492 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13990) );
  MUX2_X1 U15493 ( .A(n13990), .B(n14066), .S(n16407), .Z(n13993) );
  AOI22_X1 U15494 ( .A1(n13991), .A2(n16259), .B1(n9313), .B2(n14068), .ZN(
        n13992) );
  NAND2_X1 U15495 ( .A1(n13993), .A2(n13992), .ZN(P3_U3481) );
  INV_X1 U15496 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13994) );
  MUX2_X1 U15497 ( .A(n13994), .B(n14072), .S(n16407), .Z(n13997) );
  AOI22_X1 U15498 ( .A1(n13995), .A2(n16259), .B1(n9313), .B2(n14074), .ZN(
        n13996) );
  NAND2_X1 U15499 ( .A1(n13997), .A2(n13996), .ZN(P3_U3480) );
  INV_X1 U15500 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13998) );
  MUX2_X1 U15501 ( .A(n13998), .B(n14078), .S(n16407), .Z(n14000) );
  NAND2_X1 U15502 ( .A1(n14080), .A2(n9313), .ZN(n13999) );
  OAI211_X1 U15503 ( .C1(n14083), .C2(n14037), .A(n14000), .B(n13999), .ZN(
        P3_U3479) );
  AOI22_X1 U15504 ( .A1(n14002), .A2(n16316), .B1(n16200), .B2(n14001), .ZN(
        n14003) );
  NAND2_X1 U15505 ( .A1(n14004), .A2(n14003), .ZN(n14084) );
  MUX2_X1 U15506 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n14084), .S(n16407), .Z(
        P3_U3478) );
  AOI22_X1 U15507 ( .A1(n14006), .A2(n16316), .B1(n16200), .B2(n14005), .ZN(
        n14007) );
  NAND2_X1 U15508 ( .A1(n14008), .A2(n14007), .ZN(n14085) );
  MUX2_X1 U15509 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n14085), .S(n16407), .Z(
        P3_U3477) );
  AOI21_X1 U15510 ( .B1(n14010), .B2(n16316), .A(n14009), .ZN(n14086) );
  MUX2_X1 U15511 ( .A(n14011), .B(n14086), .S(n16407), .Z(n14012) );
  OAI21_X1 U15512 ( .B1(n14030), .B2(n14089), .A(n14012), .ZN(P3_U3476) );
  INV_X1 U15513 ( .A(n16316), .ZN(n14018) );
  OAI22_X1 U15514 ( .A1(n14014), .A2(n14018), .B1(n14013), .B2(n16311), .ZN(
        n14015) );
  MUX2_X1 U15515 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n14090), .S(n16407), .Z(
        P3_U3475) );
  OAI22_X1 U15516 ( .A1(n14019), .A2(n14018), .B1(n16311), .B2(n14017), .ZN(
        n14020) );
  NOR2_X1 U15517 ( .A1(n14021), .A2(n14020), .ZN(n14091) );
  MUX2_X1 U15518 ( .A(n15987), .B(n14091), .S(n16407), .Z(n14022) );
  INV_X1 U15519 ( .A(n14022), .ZN(P3_U3474) );
  AOI21_X1 U15520 ( .B1(n16316), .B2(n14024), .A(n14023), .ZN(n14094) );
  MUX2_X1 U15521 ( .A(n14025), .B(n14094), .S(n16407), .Z(n14026) );
  OAI21_X1 U15522 ( .B1(n14030), .B2(n14097), .A(n14026), .ZN(P3_U3473) );
  AOI21_X1 U15523 ( .B1(n14028), .B2(n16316), .A(n14027), .ZN(n14098) );
  MUX2_X1 U15524 ( .A(n15947), .B(n14098), .S(n16407), .Z(n14029) );
  OAI21_X1 U15525 ( .B1(n14030), .B2(n14101), .A(n14029), .ZN(P3_U3472) );
  INV_X1 U15526 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14035) );
  NOR2_X1 U15527 ( .A1(n14031), .A2(n16311), .ZN(n14033) );
  AOI211_X1 U15528 ( .C1(n16229), .C2(n14034), .A(n14033), .B(n14032), .ZN(
        n14103) );
  MUX2_X1 U15529 ( .A(n14035), .B(n14103), .S(n16407), .Z(n14036) );
  OAI21_X1 U15530 ( .B1(n14107), .B2(n14037), .A(n14036), .ZN(P3_U3471) );
  INV_X1 U15531 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n14040) );
  MUX2_X1 U15532 ( .A(n14041), .B(n14040), .S(n16415), .Z(n14044) );
  NAND2_X1 U15533 ( .A1(n14042), .A2(n9325), .ZN(n14043) );
  OAI211_X1 U15534 ( .C1(n14045), .C2(n14106), .A(n14044), .B(n14043), .ZN(
        P3_U3454) );
  INV_X1 U15535 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n14046) );
  MUX2_X1 U15536 ( .A(n14047), .B(n14046), .S(n16415), .Z(n14050) );
  NAND2_X1 U15537 ( .A1(n14048), .A2(n9325), .ZN(n14049) );
  OAI211_X1 U15538 ( .C1(n14051), .C2(n14106), .A(n14050), .B(n14049), .ZN(
        P3_U3453) );
  MUX2_X1 U15539 ( .A(n14052), .B(P3_REG0_REG_25__SCAN_IN), .S(n16415), .Z(
        n14055) );
  OAI22_X1 U15540 ( .A1(n14053), .A2(n14106), .B1(n8038), .B2(n14102), .ZN(
        n14054) );
  OR2_X1 U15541 ( .A1(n14055), .A2(n14054), .ZN(P3_U3452) );
  INV_X1 U15542 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n14056) );
  MUX2_X1 U15543 ( .A(n14057), .B(n14056), .S(n16415), .Z(n14060) );
  NAND2_X1 U15544 ( .A1(n14058), .A2(n9325), .ZN(n14059) );
  OAI211_X1 U15545 ( .C1(n14061), .C2(n14106), .A(n14060), .B(n14059), .ZN(
        P3_U3451) );
  INV_X1 U15546 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n14063) );
  MUX2_X1 U15547 ( .A(n14063), .B(n14062), .S(n16410), .Z(n14064) );
  OAI21_X1 U15548 ( .B1(n14065), .B2(n14102), .A(n14064), .ZN(P3_U3450) );
  INV_X1 U15549 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n14067) );
  MUX2_X1 U15550 ( .A(n14067), .B(n14066), .S(n16410), .Z(n14070) );
  NAND2_X1 U15551 ( .A1(n14068), .A2(n9325), .ZN(n14069) );
  OAI211_X1 U15552 ( .C1(n14071), .C2(n14106), .A(n14070), .B(n14069), .ZN(
        P3_U3449) );
  INV_X1 U15553 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n14073) );
  MUX2_X1 U15554 ( .A(n14073), .B(n14072), .S(n16410), .Z(n14076) );
  NAND2_X1 U15555 ( .A1(n14074), .A2(n9325), .ZN(n14075) );
  OAI211_X1 U15556 ( .C1(n14077), .C2(n14106), .A(n14076), .B(n14075), .ZN(
        P3_U3448) );
  MUX2_X1 U15557 ( .A(n14079), .B(n14078), .S(n16410), .Z(n14082) );
  NAND2_X1 U15558 ( .A1(n14080), .A2(n9325), .ZN(n14081) );
  OAI211_X1 U15559 ( .C1(n14083), .C2(n14106), .A(n14082), .B(n14081), .ZN(
        P3_U3447) );
  MUX2_X1 U15560 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n14084), .S(n16410), .Z(
        P3_U3446) );
  MUX2_X1 U15561 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n14085), .S(n16410), .Z(
        P3_U3444) );
  INV_X1 U15562 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n14087) );
  MUX2_X1 U15563 ( .A(n14087), .B(n14086), .S(n16410), .Z(n14088) );
  OAI21_X1 U15564 ( .B1(n14102), .B2(n14089), .A(n14088), .ZN(P3_U3441) );
  MUX2_X1 U15565 ( .A(n14090), .B(P3_REG0_REG_16__SCAN_IN), .S(n16415), .Z(
        P3_U3438) );
  INV_X1 U15566 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n14092) );
  MUX2_X1 U15567 ( .A(n14092), .B(n14091), .S(n16410), .Z(n14093) );
  INV_X1 U15568 ( .A(n14093), .ZN(P3_U3435) );
  INV_X1 U15569 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n14095) );
  MUX2_X1 U15570 ( .A(n14095), .B(n14094), .S(n16410), .Z(n14096) );
  OAI21_X1 U15571 ( .B1(n14102), .B2(n14097), .A(n14096), .ZN(P3_U3432) );
  INV_X1 U15572 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14099) );
  MUX2_X1 U15573 ( .A(n14099), .B(n14098), .S(n16410), .Z(n14100) );
  OAI21_X1 U15574 ( .B1(n14102), .B2(n14101), .A(n14100), .ZN(P3_U3429) );
  INV_X1 U15575 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14104) );
  MUX2_X1 U15576 ( .A(n14104), .B(n14103), .S(n16410), .Z(n14105) );
  OAI21_X1 U15577 ( .B1(n14107), .B2(n14106), .A(n14105), .ZN(P3_U3426) );
  MUX2_X1 U15578 ( .A(P3_D_REG_1__SCAN_IN), .B(n14108), .S(n14109), .Z(
        P3_U3377) );
  MUX2_X1 U15579 ( .A(P3_D_REG_0__SCAN_IN), .B(n14110), .S(n14109), .Z(
        P3_U3376) );
  INV_X1 U15580 ( .A(n14111), .ZN(n14116) );
  NOR4_X1 U15581 ( .A1(n14113), .A2(P3_IR_REG_30__SCAN_IN), .A3(n14112), .A4(
        P3_U3151), .ZN(n14114) );
  AOI21_X1 U15582 ( .B1(n16290), .B2(SI_31_), .A(n14114), .ZN(n14115) );
  OAI21_X1 U15583 ( .B1(n14116), .B2(n14119), .A(n14115), .ZN(P3_U3264) );
  INV_X1 U15584 ( .A(n14117), .ZN(n14118) );
  OAI222_X1 U15585 ( .A1(n13462), .A2(n15456), .B1(P3_U3151), .B2(n14120), 
        .C1(n14119), .C2(n14118), .ZN(P3_U3266) );
  MUX2_X1 U15586 ( .A(n14121), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  XNOR2_X1 U15587 ( .A(n14667), .B(n11516), .ZN(n14126) );
  NOR2_X1 U15588 ( .A1(n14524), .A2(n14507), .ZN(n14128) );
  XNOR2_X1 U15589 ( .A(n14126), .B(n14128), .ZN(n14165) );
  INV_X1 U15590 ( .A(n14126), .ZN(n14127) );
  XNOR2_X1 U15591 ( .A(n14493), .B(n8716), .ZN(n14129) );
  NOR2_X1 U15592 ( .A1(n14345), .A2(n14507), .ZN(n14130) );
  XNOR2_X1 U15593 ( .A(n14129), .B(n14130), .ZN(n14206) );
  XNOR2_X1 U15594 ( .A(n14476), .B(n11516), .ZN(n14131) );
  NOR2_X1 U15595 ( .A1(n14487), .A2(n14507), .ZN(n14133) );
  XNOR2_X1 U15596 ( .A(n14131), .B(n14133), .ZN(n14186) );
  INV_X1 U15597 ( .A(n14131), .ZN(n14132) );
  XNOR2_X1 U15598 ( .A(n14599), .B(n11516), .ZN(n14135) );
  XNOR2_X1 U15599 ( .A(n14134), .B(n14135), .ZN(n14215) );
  AND2_X1 U15600 ( .A1(n14437), .A2(n14445), .ZN(n14214) );
  XNOR2_X1 U15601 ( .A(n14446), .B(n11516), .ZN(n14136) );
  XNOR2_X1 U15602 ( .A(n14137), .B(n14136), .ZN(n14158) );
  INV_X1 U15603 ( .A(n14352), .ZN(n14456) );
  NOR2_X1 U15604 ( .A1(n14456), .A2(n14507), .ZN(n14157) );
  XNOR2_X1 U15605 ( .A(n14657), .B(n11516), .ZN(n14138) );
  NOR2_X1 U15606 ( .A1(n14353), .A2(n14507), .ZN(n14139) );
  XNOR2_X1 U15607 ( .A(n14138), .B(n14139), .ZN(n14200) );
  INV_X1 U15608 ( .A(n14138), .ZN(n14140) );
  NAND2_X1 U15609 ( .A1(n14140), .A2(n14139), .ZN(n14141) );
  XNOR2_X1 U15610 ( .A(n14412), .B(n11516), .ZN(n14144) );
  NAND2_X1 U15611 ( .A1(n14354), .A2(n14445), .ZN(n14142) );
  XNOR2_X1 U15612 ( .A(n14144), .B(n14142), .ZN(n14193) );
  INV_X1 U15613 ( .A(n14142), .ZN(n14143) );
  NAND2_X1 U15614 ( .A1(n14144), .A2(n14143), .ZN(n14145) );
  NAND2_X1 U15615 ( .A1(n14146), .A2(n14145), .ZN(n14240) );
  XNOR2_X1 U15616 ( .A(n14401), .B(n11516), .ZN(n14149) );
  OR2_X1 U15617 ( .A1(n14355), .A2(n14147), .ZN(n14148) );
  NAND2_X1 U15618 ( .A1(n14149), .A2(n14148), .ZN(n14150) );
  OAI21_X1 U15619 ( .B1(n14149), .B2(n14148), .A(n14150), .ZN(n14241) );
  XNOR2_X1 U15620 ( .A(n14383), .B(n11516), .ZN(n14174) );
  NAND2_X1 U15621 ( .A1(n14356), .A2(n14445), .ZN(n14173) );
  XNOR2_X1 U15622 ( .A(n14174), .B(n14173), .ZN(n14175) );
  XNOR2_X1 U15623 ( .A(n14176), .B(n14175), .ZN(n14156) );
  INV_X1 U15624 ( .A(n14151), .ZN(n14380) );
  OAI22_X1 U15625 ( .A1(n14152), .A2(n14523), .B1(n14355), .B2(n14521), .ZN(
        n14386) );
  AOI22_X1 U15626 ( .A1(n14195), .A2(n14386), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14153) );
  OAI21_X1 U15627 ( .B1(n14380), .B2(n14218), .A(n14153), .ZN(n14154) );
  AOI21_X1 U15628 ( .B1(n14574), .B2(n14246), .A(n14154), .ZN(n14155) );
  OAI21_X1 U15629 ( .B1(n14156), .B2(n14248), .A(n14155), .ZN(P2_U3186) );
  XNOR2_X1 U15630 ( .A(n14158), .B(n14157), .ZN(n14164) );
  OAI22_X1 U15631 ( .A1(n14353), .A2(n14217), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14159), .ZN(n14162) );
  INV_X1 U15632 ( .A(n14447), .ZN(n14160) );
  OAI22_X1 U15633 ( .A1(n14350), .A2(n14219), .B1(n14160), .B2(n14218), .ZN(
        n14161) );
  AOI211_X1 U15634 ( .C1(n14446), .C2(n14246), .A(n14162), .B(n14161), .ZN(
        n14163) );
  OAI21_X1 U15635 ( .B1(n14164), .B2(n14248), .A(n14163), .ZN(P2_U3188) );
  XNOR2_X1 U15636 ( .A(n14166), .B(n14165), .ZN(n14172) );
  OR2_X1 U15637 ( .A1(n14345), .A2(n14523), .ZN(n14168) );
  OR2_X1 U15638 ( .A1(n14326), .A2(n14521), .ZN(n14167) );
  NAND2_X1 U15639 ( .A1(n14168), .A2(n14167), .ZN(n14499) );
  AND2_X1 U15640 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n14304) );
  AOI21_X1 U15641 ( .B1(n14499), .B2(n14195), .A(n14304), .ZN(n14169) );
  OAI21_X1 U15642 ( .B1(n14509), .B2(n14218), .A(n14169), .ZN(n14170) );
  AOI21_X1 U15643 ( .B1(n14505), .B2(n14246), .A(n14170), .ZN(n14171) );
  OAI21_X1 U15644 ( .B1(n14172), .B2(n14248), .A(n14171), .ZN(P2_U3191) );
  NAND2_X1 U15645 ( .A1(n14363), .A2(n14445), .ZN(n14177) );
  XNOR2_X1 U15646 ( .A(n14177), .B(n11516), .ZN(n14178) );
  XNOR2_X1 U15647 ( .A(n14569), .B(n14178), .ZN(n14179) );
  INV_X1 U15648 ( .A(n14371), .ZN(n14183) );
  INV_X1 U15649 ( .A(n14250), .ZN(n14181) );
  OAI22_X1 U15650 ( .A1(n14181), .A2(n14523), .B1(n14180), .B2(n14521), .ZN(
        n14369) );
  AOI22_X1 U15651 ( .A1(n14195), .A2(n14369), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14182) );
  OAI21_X1 U15652 ( .B1(n14183), .B2(n14218), .A(n14182), .ZN(n14184) );
  AOI21_X1 U15653 ( .B1(n14569), .B2(n14246), .A(n14184), .ZN(n14185) );
  XNOR2_X1 U15654 ( .A(n14187), .B(n14186), .ZN(n14192) );
  INV_X1 U15655 ( .A(n14474), .ZN(n14189) );
  OAI22_X1 U15656 ( .A1(n14350), .A2(n14523), .B1(n14345), .B2(n14521), .ZN(
        n14470) );
  AOI22_X1 U15657 ( .A1(n14470), .A2(n14195), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14188) );
  OAI21_X1 U15658 ( .B1(n14189), .B2(n14218), .A(n14188), .ZN(n14190) );
  AOI21_X1 U15659 ( .B1(n14603), .B2(n14246), .A(n14190), .ZN(n14191) );
  OAI21_X1 U15660 ( .B1(n14192), .B2(n14248), .A(n14191), .ZN(P2_U3195) );
  XNOR2_X1 U15661 ( .A(n14194), .B(n14193), .ZN(n14199) );
  OAI22_X1 U15662 ( .A1(n14353), .A2(n14521), .B1(n14355), .B2(n14523), .ZN(
        n14408) );
  AOI22_X1 U15663 ( .A1(n14408), .A2(n14195), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14196) );
  OAI21_X1 U15664 ( .B1(n14413), .B2(n14218), .A(n14196), .ZN(n14197) );
  AOI21_X1 U15665 ( .B1(n14412), .B2(n14246), .A(n14197), .ZN(n14198) );
  OAI21_X1 U15666 ( .B1(n14199), .B2(n14248), .A(n14198), .ZN(P2_U3197) );
  XNOR2_X1 U15667 ( .A(n14201), .B(n14200), .ZN(n14205) );
  AOI22_X1 U15668 ( .A1(n14354), .A2(n14439), .B1(n14438), .B2(n14352), .ZN(
        n14424) );
  AOI22_X1 U15669 ( .A1(n14428), .A2(n14242), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14202) );
  OAI21_X1 U15670 ( .B1(n14424), .B2(n14244), .A(n14202), .ZN(n14203) );
  AOI21_X1 U15671 ( .B1(n14427), .B2(n14246), .A(n14203), .ZN(n14204) );
  OAI21_X1 U15672 ( .B1(n14205), .B2(n14248), .A(n14204), .ZN(P2_U3201) );
  XNOR2_X1 U15673 ( .A(n14207), .B(n14206), .ZN(n14213) );
  INV_X1 U15674 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n14208) );
  OAI22_X1 U15675 ( .A1(n14487), .A2(n14217), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14208), .ZN(n14211) );
  OAI22_X1 U15676 ( .A1(n14219), .A2(n14524), .B1(n14209), .B2(n14218), .ZN(
        n14210) );
  AOI211_X1 U15677 ( .C1(n14609), .C2(n14246), .A(n14211), .B(n14210), .ZN(
        n14212) );
  OAI21_X1 U15678 ( .B1(n14213), .B2(n14248), .A(n14212), .ZN(P2_U3205) );
  XNOR2_X1 U15679 ( .A(n14215), .B(n14214), .ZN(n14223) );
  OAI22_X1 U15680 ( .A1(n14456), .A2(n14217), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14216), .ZN(n14221) );
  OAI22_X1 U15681 ( .A1(n14487), .A2(n14219), .B1(n14218), .B2(n14459), .ZN(
        n14220) );
  AOI211_X1 U15682 ( .C1(n14599), .C2(n14246), .A(n14221), .B(n14220), .ZN(
        n14222) );
  OAI21_X1 U15683 ( .B1(n14223), .B2(n14248), .A(n14222), .ZN(P2_U3207) );
  AOI22_X1 U15684 ( .A1(n14225), .A2(n14264), .B1(n14224), .B2(n14246), .ZN(
        n14237) );
  AOI22_X1 U15685 ( .A1(n14227), .A2(n14266), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n14226), .ZN(n14236) );
  INV_X1 U15686 ( .A(n14228), .ZN(n14234) );
  NOR3_X1 U15687 ( .A1(n14231), .A2(n14230), .A3(n14229), .ZN(n14233) );
  OAI21_X1 U15688 ( .B1(n14234), .B2(n14233), .A(n14232), .ZN(n14235) );
  NAND3_X1 U15689 ( .A1(n14237), .A2(n14236), .A3(n14235), .ZN(P2_U3209) );
  INV_X1 U15690 ( .A(n14238), .ZN(n14239) );
  AOI21_X1 U15691 ( .B1(n14241), .B2(n14240), .A(n14239), .ZN(n14249) );
  AOI22_X1 U15692 ( .A1(n14354), .A2(n14438), .B1(n14439), .B2(n14356), .ZN(
        n14394) );
  AOI22_X1 U15693 ( .A1(n14242), .A2(n14398), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14243) );
  OAI21_X1 U15694 ( .B1(n14394), .B2(n14244), .A(n14243), .ZN(n14245) );
  AOI21_X1 U15695 ( .B1(n14580), .B2(n14246), .A(n14245), .ZN(n14247) );
  OAI21_X1 U15696 ( .B1(n14249), .B2(n14248), .A(n14247), .ZN(P2_U3212) );
  MUX2_X1 U15697 ( .A(n14316), .B(P2_DATAO_REG_31__SCAN_IN), .S(n14267), .Z(
        P2_U3562) );
  MUX2_X1 U15698 ( .A(n14362), .B(P2_DATAO_REG_30__SCAN_IN), .S(n14267), .Z(
        P2_U3561) );
  MUX2_X1 U15699 ( .A(n14250), .B(P2_DATAO_REG_29__SCAN_IN), .S(n14267), .Z(
        P2_U3560) );
  MUX2_X1 U15700 ( .A(n14363), .B(P2_DATAO_REG_28__SCAN_IN), .S(n14267), .Z(
        P2_U3559) );
  MUX2_X1 U15701 ( .A(n14356), .B(P2_DATAO_REG_27__SCAN_IN), .S(n14267), .Z(
        P2_U3558) );
  MUX2_X1 U15702 ( .A(n14330), .B(P2_DATAO_REG_26__SCAN_IN), .S(n14267), .Z(
        P2_U3557) );
  MUX2_X1 U15703 ( .A(n14354), .B(P2_DATAO_REG_25__SCAN_IN), .S(n14267), .Z(
        P2_U3556) );
  MUX2_X1 U15704 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n14440), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U15705 ( .A(n14352), .B(P2_DATAO_REG_23__SCAN_IN), .S(n14267), .Z(
        P2_U3554) );
  MUX2_X1 U15706 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n14437), .S(P2_U3947), .Z(
        P2_U3553) );
  INV_X1 U15707 ( .A(n14487), .ZN(n14329) );
  MUX2_X1 U15708 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n14329), .S(P2_U3947), .Z(
        P2_U3552) );
  MUX2_X1 U15709 ( .A(n14344), .B(P2_DATAO_REG_20__SCAN_IN), .S(n14267), .Z(
        P2_U3551) );
  INV_X1 U15710 ( .A(n14524), .ZN(n14343) );
  MUX2_X1 U15711 ( .A(n14343), .B(P2_DATAO_REG_19__SCAN_IN), .S(n14267), .Z(
        P2_U3550) );
  MUX2_X1 U15712 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n14340), .S(P2_U3947), .Z(
        P2_U3549) );
  MUX2_X1 U15713 ( .A(n14324), .B(P2_DATAO_REG_17__SCAN_IN), .S(n14267), .Z(
        P2_U3548) );
  MUX2_X1 U15714 ( .A(n14251), .B(P2_DATAO_REG_16__SCAN_IN), .S(n14267), .Z(
        P2_U3547) );
  MUX2_X1 U15715 ( .A(n14252), .B(P2_DATAO_REG_15__SCAN_IN), .S(n14267), .Z(
        P2_U3546) );
  MUX2_X1 U15716 ( .A(n14253), .B(P2_DATAO_REG_14__SCAN_IN), .S(n14267), .Z(
        P2_U3545) );
  MUX2_X1 U15717 ( .A(n14254), .B(P2_DATAO_REG_13__SCAN_IN), .S(n14267), .Z(
        P2_U3544) );
  MUX2_X1 U15718 ( .A(n14255), .B(P2_DATAO_REG_12__SCAN_IN), .S(n14267), .Z(
        P2_U3543) );
  MUX2_X1 U15719 ( .A(n14256), .B(P2_DATAO_REG_11__SCAN_IN), .S(n14267), .Z(
        P2_U3542) );
  MUX2_X1 U15720 ( .A(n14257), .B(P2_DATAO_REG_10__SCAN_IN), .S(n14267), .Z(
        P2_U3541) );
  MUX2_X1 U15721 ( .A(n14258), .B(P2_DATAO_REG_9__SCAN_IN), .S(n14267), .Z(
        P2_U3540) );
  MUX2_X1 U15722 ( .A(n14259), .B(P2_DATAO_REG_8__SCAN_IN), .S(n14267), .Z(
        P2_U3539) );
  MUX2_X1 U15723 ( .A(n14260), .B(P2_DATAO_REG_7__SCAN_IN), .S(n14267), .Z(
        P2_U3538) );
  MUX2_X1 U15724 ( .A(n14261), .B(P2_DATAO_REG_6__SCAN_IN), .S(n14267), .Z(
        P2_U3537) );
  MUX2_X1 U15725 ( .A(n14262), .B(P2_DATAO_REG_5__SCAN_IN), .S(n14267), .Z(
        P2_U3536) );
  MUX2_X1 U15726 ( .A(n14263), .B(P2_DATAO_REG_4__SCAN_IN), .S(n14267), .Z(
        P2_U3535) );
  MUX2_X1 U15727 ( .A(n14264), .B(P2_DATAO_REG_3__SCAN_IN), .S(n14267), .Z(
        P2_U3534) );
  MUX2_X1 U15728 ( .A(n14265), .B(P2_DATAO_REG_2__SCAN_IN), .S(n14267), .Z(
        P2_U3533) );
  MUX2_X1 U15729 ( .A(n14266), .B(P2_DATAO_REG_1__SCAN_IN), .S(n14267), .Z(
        P2_U3532) );
  MUX2_X1 U15730 ( .A(n14268), .B(P2_DATAO_REG_0__SCAN_IN), .S(n14267), .Z(
        P2_U3531) );
  AOI21_X1 U15731 ( .B1(n14273), .B2(P2_REG1_REG_16__SCAN_IN), .A(n14269), 
        .ZN(n14271) );
  XNOR2_X1 U15732 ( .A(n14288), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14270) );
  NOR2_X1 U15733 ( .A1(n14270), .A2(n14271), .ZN(n14287) );
  AOI211_X1 U15734 ( .C1(n14271), .C2(n14270), .A(n14287), .B(n15813), .ZN(
        n14277) );
  XNOR2_X1 U15735 ( .A(n14288), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n14274) );
  NOR2_X1 U15736 ( .A1(n14274), .A2(n14275), .ZN(n14282) );
  AOI211_X1 U15737 ( .C1(n14275), .C2(n14274), .A(n14282), .B(n15817), .ZN(
        n14276) );
  NOR2_X1 U15738 ( .A1(n14277), .A2(n14276), .ZN(n14280) );
  AOI21_X1 U15739 ( .B1(n15800), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n14278), 
        .ZN(n14279) );
  OAI211_X1 U15740 ( .C1(n14281), .C2(n14306), .A(n14280), .B(n14279), .ZN(
        P2_U3231) );
  XNOR2_X1 U15741 ( .A(n14295), .B(n14294), .ZN(n14293) );
  XNOR2_X1 U15742 ( .A(n14293), .B(n11940), .ZN(n14292) );
  INV_X1 U15743 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n14284) );
  OAI21_X1 U15744 ( .B1(n15844), .B2(n14284), .A(n14283), .ZN(n14285) );
  AOI21_X1 U15745 ( .B1(n14286), .B2(n15838), .A(n14285), .ZN(n14291) );
  OAI211_X1 U15746 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n14289), .A(n15835), 
        .B(n14300), .ZN(n14290) );
  OAI211_X1 U15747 ( .C1(n15817), .C2(n14292), .A(n14291), .B(n14290), .ZN(
        P2_U3232) );
  MUX2_X1 U15748 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n12284), .S(n9660), .Z(
        n14297) );
  INV_X1 U15749 ( .A(n14293), .ZN(n14296) );
  INV_X1 U15750 ( .A(n14298), .ZN(n14299) );
  NAND2_X1 U15751 ( .A1(n14300), .A2(n14299), .ZN(n14303) );
  XNOR2_X1 U15752 ( .A(n14301), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n14302) );
  AOI21_X1 U15753 ( .B1(n15800), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n14304), 
        .ZN(n14305) );
  OAI21_X1 U15754 ( .B1(n14306), .B2(n9660), .A(n14305), .ZN(n14307) );
  OAI21_X1 U15755 ( .B1(n14309), .B2(n15817), .A(n14308), .ZN(P2_U3233) );
  INV_X1 U15756 ( .A(n14563), .ZN(n14335) );
  NAND2_X1 U15757 ( .A1(n14490), .A2(n14476), .ZN(n14473) );
  XNOR2_X1 U15758 ( .A(n14319), .B(n14311), .ZN(n14312) );
  NOR2_X1 U15759 ( .A1(n14312), .A2(n14445), .ZN(n14555) );
  NAND2_X1 U15760 ( .A1(n14555), .A2(n16306), .ZN(n14318) );
  NOR2_X1 U15761 ( .A1(n14314), .A2(n14313), .ZN(n14315) );
  NOR2_X1 U15762 ( .A1(n14523), .A2(n14315), .ZN(n14361) );
  AND2_X1 U15763 ( .A1(n14361), .A2(n14316), .ZN(n14554) );
  INV_X1 U15764 ( .A(n14554), .ZN(n14558) );
  NOR2_X1 U15765 ( .A1(n16405), .A2(n14558), .ZN(n14321) );
  AOI21_X1 U15766 ( .B1(n16405), .B2(P2_REG2_REG_31__SCAN_IN), .A(n14321), 
        .ZN(n14317) );
  OAI211_X1 U15767 ( .C1(n14641), .C2(n16398), .A(n14318), .B(n14317), .ZN(
        P2_U3234) );
  OAI211_X1 U15768 ( .C1(n14645), .C2(n7458), .A(n14507), .B(n14319), .ZN(
        n14559) );
  NOR2_X1 U15769 ( .A1(n14645), .A2(n16398), .ZN(n14320) );
  AOI211_X1 U15770 ( .C1(n16405), .C2(P2_REG2_REG_30__SCAN_IN), .A(n14321), 
        .B(n14320), .ZN(n14322) );
  OAI21_X1 U15771 ( .B1(n14539), .B2(n14559), .A(n14322), .ZN(P2_U3235) );
  OR2_X1 U15772 ( .A1(n14336), .A2(n14324), .ZN(n14325) );
  NAND2_X1 U15773 ( .A1(n14517), .A2(n14526), .ZN(n14519) );
  NAND2_X1 U15774 ( .A1(n14619), .A2(n14326), .ZN(n14327) );
  NAND2_X1 U15775 ( .A1(n14519), .A2(n14327), .ZN(n14502) );
  NAND2_X1 U15776 ( .A1(n14502), .A2(n14501), .ZN(n14504) );
  NAND2_X1 U15777 ( .A1(n14609), .A2(n14344), .ZN(n14328) );
  INV_X1 U15778 ( .A(n14420), .ZN(n14422) );
  OAI21_X1 U15779 ( .B1(n14363), .B2(n14569), .A(n14365), .ZN(n14331) );
  INV_X1 U15780 ( .A(n14370), .ZN(n14332) );
  AOI22_X1 U15781 ( .A1(n16405), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n14333), 
        .B2(n16394), .ZN(n14334) );
  OAI21_X1 U15782 ( .B1(n14335), .B2(n16398), .A(n14334), .ZN(n14364) );
  NOR2_X1 U15783 ( .A1(n14336), .A2(n14522), .ZN(n14337) );
  NAND2_X1 U15784 ( .A1(n14619), .A2(n14340), .ZN(n14342) );
  NOR2_X1 U15785 ( .A1(n14619), .A2(n14340), .ZN(n14341) );
  NOR2_X1 U15786 ( .A1(n14493), .A2(n14344), .ZN(n14346) );
  INV_X1 U15787 ( .A(n14347), .ZN(n14349) );
  INV_X1 U15788 ( .A(n14357), .ZN(n14358) );
  INV_X1 U15789 ( .A(n14569), .ZN(n14374) );
  AOI211_X1 U15790 ( .C1(n14569), .C2(n14378), .A(n14445), .B(n14370), .ZN(
        n14568) );
  NAND2_X1 U15791 ( .A1(n14568), .A2(n16306), .ZN(n14373) );
  AOI22_X1 U15792 ( .A1(n16405), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n14371), 
        .B2(n16394), .ZN(n14372) );
  OAI211_X1 U15793 ( .C1(n14374), .C2(n16398), .A(n14373), .B(n14372), .ZN(
        n14375) );
  AOI21_X1 U15794 ( .B1(n14567), .B2(n16401), .A(n14375), .ZN(n14376) );
  OAI21_X1 U15795 ( .B1(n14571), .B2(n16405), .A(n14376), .ZN(P2_U3237) );
  XNOR2_X1 U15796 ( .A(n14377), .B(n14384), .ZN(n14577) );
  OAI211_X1 U15797 ( .C1(n14383), .C2(n14396), .A(n14507), .B(n14378), .ZN(
        n14379) );
  INV_X1 U15798 ( .A(n14379), .ZN(n14573) );
  NOR2_X1 U15799 ( .A1(n14510), .A2(n14380), .ZN(n14381) );
  AOI21_X1 U15800 ( .B1(n16405), .B2(P2_REG2_REG_27__SCAN_IN), .A(n14381), 
        .ZN(n14382) );
  OAI21_X1 U15801 ( .B1(n14383), .B2(n16398), .A(n14382), .ZN(n14389) );
  XNOR2_X1 U15802 ( .A(n14385), .B(n14384), .ZN(n14387) );
  AOI21_X1 U15803 ( .B1(n14387), .B2(n14529), .A(n14386), .ZN(n14576) );
  NOR2_X1 U15804 ( .A1(n14576), .A2(n16405), .ZN(n14388) );
  AOI211_X1 U15805 ( .C1(n14573), .C2(n16306), .A(n14389), .B(n14388), .ZN(
        n14390) );
  OAI21_X1 U15806 ( .B1(n14497), .B2(n14577), .A(n14390), .ZN(P2_U3238) );
  XNOR2_X1 U15807 ( .A(n14391), .B(n14393), .ZN(n14581) );
  XOR2_X1 U15808 ( .A(n14393), .B(n14392), .Z(n14395) );
  OAI21_X1 U15809 ( .B1(n14395), .B2(n14486), .A(n14394), .ZN(n14578) );
  OAI21_X1 U15810 ( .B1(n14401), .B2(n14411), .A(n14507), .ZN(n14397) );
  NOR2_X1 U15811 ( .A1(n14397), .A2(n14396), .ZN(n14579) );
  NAND2_X1 U15812 ( .A1(n14579), .A2(n16306), .ZN(n14400) );
  AOI22_X1 U15813 ( .A1(n16405), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n14398), 
        .B2(n16394), .ZN(n14399) );
  OAI211_X1 U15814 ( .C1(n14401), .C2(n16398), .A(n14400), .B(n14399), .ZN(
        n14402) );
  AOI21_X1 U15815 ( .B1(n14578), .B2(n14549), .A(n14402), .ZN(n14403) );
  OAI21_X1 U15816 ( .B1(n14497), .B2(n14581), .A(n14403), .ZN(P2_U3239) );
  OAI21_X1 U15817 ( .B1(n14405), .B2(n14407), .A(n14404), .ZN(n14584) );
  INV_X1 U15818 ( .A(n14584), .ZN(n14419) );
  XOR2_X1 U15819 ( .A(n14406), .B(n14407), .Z(n14410) );
  INV_X1 U15820 ( .A(n14408), .ZN(n14409) );
  OAI21_X1 U15821 ( .B1(n14410), .B2(n14486), .A(n14409), .ZN(n14582) );
  NAND2_X1 U15822 ( .A1(n14582), .A2(n14549), .ZN(n14418) );
  AOI211_X1 U15823 ( .C1(n14412), .C2(n8266), .A(n14445), .B(n14411), .ZN(
        n14583) );
  INV_X1 U15824 ( .A(n14413), .ZN(n14414) );
  AOI22_X1 U15825 ( .A1(n14414), .A2(n16394), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n16405), .ZN(n14415) );
  OAI21_X1 U15826 ( .B1(n14653), .B2(n16398), .A(n14415), .ZN(n14416) );
  AOI21_X1 U15827 ( .B1(n14583), .B2(n16306), .A(n14416), .ZN(n14417) );
  OAI211_X1 U15828 ( .C1(n14419), .C2(n14497), .A(n14418), .B(n14417), .ZN(
        P2_U3240) );
  XNOR2_X1 U15829 ( .A(n14421), .B(n14420), .ZN(n14589) );
  INV_X1 U15830 ( .A(n14589), .ZN(n14433) );
  XNOR2_X1 U15831 ( .A(n14423), .B(n14422), .ZN(n14425) );
  OAI21_X1 U15832 ( .B1(n14425), .B2(n14486), .A(n14424), .ZN(n14587) );
  NAND2_X1 U15833 ( .A1(n14587), .A2(n14549), .ZN(n14432) );
  AOI211_X1 U15834 ( .C1(n14427), .C2(n8267), .A(n14445), .B(n14426), .ZN(
        n14588) );
  AOI22_X1 U15835 ( .A1(n14428), .A2(n16394), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n16405), .ZN(n14429) );
  OAI21_X1 U15836 ( .B1(n14657), .B2(n16398), .A(n14429), .ZN(n14430) );
  AOI21_X1 U15837 ( .B1(n14588), .B2(n16306), .A(n14430), .ZN(n14431) );
  OAI211_X1 U15838 ( .C1(n14433), .C2(n14497), .A(n14432), .B(n14431), .ZN(
        P2_U3241) );
  XOR2_X1 U15839 ( .A(n14436), .B(n14434), .Z(n14594) );
  INV_X1 U15840 ( .A(n14594), .ZN(n14453) );
  XOR2_X1 U15841 ( .A(n14436), .B(n14435), .Z(n14443) );
  NAND2_X1 U15842 ( .A1(n14594), .A2(n14520), .ZN(n14442) );
  AOI22_X1 U15843 ( .A1(n14440), .A2(n14439), .B1(n14438), .B2(n14437), .ZN(
        n14441) );
  OAI211_X1 U15844 ( .C1(n14443), .C2(n14486), .A(n14442), .B(n14441), .ZN(
        n14592) );
  NAND2_X1 U15845 ( .A1(n14592), .A2(n14549), .ZN(n14451) );
  AOI211_X1 U15846 ( .C1(n14446), .C2(n14457), .A(n14445), .B(n14444), .ZN(
        n14593) );
  AOI22_X1 U15847 ( .A1(P2_REG2_REG_23__SCAN_IN), .A2(n16405), .B1(n14447), 
        .B2(n16394), .ZN(n14448) );
  OAI21_X1 U15848 ( .B1(n8265), .B2(n16398), .A(n14448), .ZN(n14449) );
  AOI21_X1 U15849 ( .B1(n14593), .B2(n16306), .A(n14449), .ZN(n14450) );
  OAI211_X1 U15850 ( .C1(n14453), .C2(n14452), .A(n14451), .B(n14450), .ZN(
        P2_U3242) );
  XNOR2_X1 U15851 ( .A(n14454), .B(n14464), .ZN(n14455) );
  OAI222_X1 U15852 ( .A1(n14521), .A2(n14487), .B1(n14523), .B2(n14456), .C1(
        n14486), .C2(n14455), .ZN(n14597) );
  AOI21_X1 U15853 ( .B1(n14473), .B2(n14599), .A(n7431), .ZN(n14458) );
  AND2_X1 U15854 ( .A1(n14458), .A2(n14457), .ZN(n14598) );
  NAND2_X1 U15855 ( .A1(n14598), .A2(n16306), .ZN(n14462) );
  INV_X1 U15856 ( .A(n14459), .ZN(n14460) );
  AOI22_X1 U15857 ( .A1(n16405), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n14460), 
        .B2(n16394), .ZN(n14461) );
  OAI211_X1 U15858 ( .C1(n14463), .C2(n16398), .A(n14462), .B(n14461), .ZN(
        n14467) );
  XNOR2_X1 U15859 ( .A(n14465), .B(n14464), .ZN(n14601) );
  NOR2_X1 U15860 ( .A1(n14601), .A2(n14497), .ZN(n14466) );
  AOI211_X1 U15861 ( .C1(n14549), .C2(n14597), .A(n14467), .B(n14466), .ZN(
        n14468) );
  INV_X1 U15862 ( .A(n14468), .ZN(P2_U3243) );
  XNOR2_X1 U15863 ( .A(n14469), .B(n14477), .ZN(n14471) );
  AOI21_X1 U15864 ( .B1(n14471), .B2(n14529), .A(n14470), .ZN(n14605) );
  OR2_X1 U15865 ( .A1(n14490), .A2(n14476), .ZN(n14472) );
  AND3_X1 U15866 ( .A1(n14473), .A2(n14507), .A3(n14472), .ZN(n14602) );
  AOI22_X1 U15867 ( .A1(n16405), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n14474), 
        .B2(n16394), .ZN(n14475) );
  OAI21_X1 U15868 ( .B1(n14476), .B2(n16398), .A(n14475), .ZN(n14480) );
  XNOR2_X1 U15869 ( .A(n14478), .B(n14477), .ZN(n14606) );
  NOR2_X1 U15870 ( .A1(n14606), .A2(n14497), .ZN(n14479) );
  AOI211_X1 U15871 ( .C1(n14602), .C2(n16306), .A(n14480), .B(n14479), .ZN(
        n14481) );
  OAI21_X1 U15872 ( .B1(n16405), .B2(n14605), .A(n14481), .ZN(P2_U3244) );
  XNOR2_X1 U15873 ( .A(n14482), .B(n14484), .ZN(n14611) );
  XOR2_X1 U15874 ( .A(n14484), .B(n14483), .Z(n14485) );
  OAI222_X1 U15875 ( .A1(n14523), .A2(n14487), .B1(n14521), .B2(n14524), .C1(
        n14486), .C2(n14485), .ZN(n14607) );
  NAND2_X1 U15876 ( .A1(n14607), .A2(n14549), .ZN(n14496) );
  NAND2_X1 U15877 ( .A1(n14508), .A2(n14609), .ZN(n14488) );
  NAND2_X1 U15878 ( .A1(n14488), .A2(n14507), .ZN(n14489) );
  NOR2_X1 U15879 ( .A1(n14490), .A2(n14489), .ZN(n14608) );
  AOI22_X1 U15880 ( .A1(n16405), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14491), 
        .B2(n16394), .ZN(n14492) );
  OAI21_X1 U15881 ( .B1(n14493), .B2(n16398), .A(n14492), .ZN(n14494) );
  AOI21_X1 U15882 ( .B1(n14608), .B2(n16306), .A(n14494), .ZN(n14495) );
  OAI211_X1 U15883 ( .C1(n14611), .C2(n14497), .A(n14496), .B(n14495), .ZN(
        P2_U3245) );
  XNOR2_X1 U15884 ( .A(n14498), .B(n14501), .ZN(n14500) );
  AOI21_X1 U15885 ( .B1(n14500), .B2(n14529), .A(n14499), .ZN(n14614) );
  OR2_X1 U15886 ( .A1(n14502), .A2(n14501), .ZN(n14503) );
  NAND2_X1 U15887 ( .A1(n14504), .A2(n14503), .ZN(n14612) );
  NAND2_X1 U15888 ( .A1(n14505), .A2(n14537), .ZN(n14506) );
  NAND3_X1 U15889 ( .A1(n14508), .A2(n14507), .A3(n14506), .ZN(n14613) );
  NOR2_X1 U15890 ( .A1(n14613), .A2(n14539), .ZN(n14514) );
  NOR2_X1 U15891 ( .A1(n14510), .A2(n14509), .ZN(n14511) );
  AOI21_X1 U15892 ( .B1(n16405), .B2(P2_REG2_REG_19__SCAN_IN), .A(n14511), 
        .ZN(n14512) );
  OAI21_X1 U15893 ( .B1(n14667), .B2(n16398), .A(n14512), .ZN(n14513) );
  AOI211_X1 U15894 ( .C1(n14612), .C2(n14515), .A(n14514), .B(n14513), .ZN(
        n14516) );
  OAI21_X1 U15895 ( .B1(n16405), .B2(n14614), .A(n14516), .ZN(P2_U3246) );
  OR2_X1 U15896 ( .A1(n14517), .A2(n14526), .ZN(n14518) );
  NAND2_X1 U15897 ( .A1(n14519), .A2(n14518), .ZN(n14621) );
  NAND2_X1 U15898 ( .A1(n14621), .A2(n14520), .ZN(n14533) );
  OAI22_X1 U15899 ( .A1(n14524), .A2(n14523), .B1(n14522), .B2(n14521), .ZN(
        n14525) );
  INV_X1 U15900 ( .A(n14525), .ZN(n14532) );
  INV_X1 U15901 ( .A(n14526), .ZN(n14527) );
  XNOR2_X1 U15902 ( .A(n14528), .B(n14527), .ZN(n14530) );
  NAND2_X1 U15903 ( .A1(n14530), .A2(n14529), .ZN(n14531) );
  AOI21_X1 U15904 ( .B1(n14536), .B2(n14535), .A(n7431), .ZN(n14538) );
  NAND2_X1 U15905 ( .A1(n14538), .A2(n14537), .ZN(n14618) );
  NOR2_X1 U15906 ( .A1(n14618), .A2(n14539), .ZN(n14543) );
  AOI22_X1 U15907 ( .A1(n16405), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14540), 
        .B2(n16394), .ZN(n14541) );
  OAI21_X1 U15908 ( .B1(n14619), .B2(n16398), .A(n14541), .ZN(n14542) );
  AOI211_X1 U15909 ( .C1(n14621), .C2(n16401), .A(n14543), .B(n14542), .ZN(
        n14544) );
  OAI21_X1 U15910 ( .B1(n14623), .B2(n16405), .A(n14544), .ZN(P2_U3247) );
  AOI22_X1 U15911 ( .A1(n16306), .A2(n14546), .B1(n16401), .B2(n14545), .ZN(
        n14553) );
  AOI22_X1 U15912 ( .A1(n16303), .A2(n14547), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n16394), .ZN(n14552) );
  INV_X1 U15913 ( .A(n14548), .ZN(n14550) );
  MUX2_X1 U15914 ( .A(n9551), .B(n14550), .S(n14549), .Z(n14551) );
  NAND3_X1 U15915 ( .A1(n14553), .A2(n14552), .A3(n14551), .ZN(P2_U3264) );
  NOR2_X1 U15916 ( .A1(n14555), .A2(n14554), .ZN(n14638) );
  MUX2_X1 U15917 ( .A(n14556), .B(n14638), .S(n16358), .Z(n14557) );
  OAI21_X1 U15918 ( .B1(n14641), .B2(n14631), .A(n14557), .ZN(P2_U3530) );
  NAND2_X1 U15919 ( .A1(n14559), .A2(n14558), .ZN(n14642) );
  MUX2_X1 U15920 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n14642), .S(n16358), .Z(
        n14560) );
  INV_X1 U15921 ( .A(n14560), .ZN(n14561) );
  OAI21_X1 U15922 ( .B1(n14645), .B2(n14631), .A(n14561), .ZN(P2_U3529) );
  AOI21_X1 U15923 ( .B1(n16170), .B2(n14563), .A(n14562), .ZN(n14564) );
  INV_X1 U15924 ( .A(n14567), .ZN(n14572) );
  AOI21_X1 U15925 ( .B1(n16170), .B2(n14569), .A(n14568), .ZN(n14570) );
  OAI211_X1 U15926 ( .C1(n14572), .C2(n9885), .A(n14571), .B(n14570), .ZN(
        n14647) );
  MUX2_X1 U15927 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n14647), .S(n16358), .Z(
        P2_U3527) );
  AOI21_X1 U15928 ( .B1(n16170), .B2(n14574), .A(n14573), .ZN(n14575) );
  OAI211_X1 U15929 ( .C1(n16262), .C2(n14577), .A(n14576), .B(n14575), .ZN(
        n14648) );
  MUX2_X1 U15930 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14648), .S(n16358), .Z(
        P2_U3526) );
  MUX2_X1 U15931 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14649), .S(n16358), .Z(
        P2_U3525) );
  AOI211_X1 U15932 ( .C1(n16348), .C2(n14584), .A(n14583), .B(n14582), .ZN(
        n14650) );
  MUX2_X1 U15933 ( .A(n14585), .B(n14650), .S(n16358), .Z(n14586) );
  OAI21_X1 U15934 ( .B1(n14653), .B2(n14631), .A(n14586), .ZN(P2_U3524) );
  AOI211_X1 U15935 ( .C1(n16348), .C2(n14589), .A(n14588), .B(n14587), .ZN(
        n14654) );
  MUX2_X1 U15936 ( .A(n14590), .B(n14654), .S(n16358), .Z(n14591) );
  OAI21_X1 U15937 ( .B1(n14657), .B2(n14631), .A(n14591), .ZN(P2_U3523) );
  AOI211_X1 U15938 ( .C1(n13099), .C2(n14594), .A(n14593), .B(n14592), .ZN(
        n14658) );
  MUX2_X1 U15939 ( .A(n14595), .B(n14658), .S(n16358), .Z(n14596) );
  OAI21_X1 U15940 ( .B1(n8265), .B2(n14631), .A(n14596), .ZN(P2_U3522) );
  AOI211_X1 U15941 ( .C1(n16170), .C2(n14599), .A(n14598), .B(n14597), .ZN(
        n14600) );
  OAI21_X1 U15942 ( .B1(n16262), .B2(n14601), .A(n14600), .ZN(n14661) );
  MUX2_X1 U15943 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14661), .S(n16358), .Z(
        P2_U3521) );
  AOI21_X1 U15944 ( .B1(n16170), .B2(n14603), .A(n14602), .ZN(n14604) );
  OAI211_X1 U15945 ( .C1(n14606), .C2(n16262), .A(n14605), .B(n14604), .ZN(
        n14662) );
  MUX2_X1 U15946 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14662), .S(n16358), .Z(
        P2_U3520) );
  AOI211_X1 U15947 ( .C1(n16170), .C2(n14609), .A(n14608), .B(n14607), .ZN(
        n14610) );
  OAI21_X1 U15948 ( .B1(n16262), .B2(n14611), .A(n14610), .ZN(n14663) );
  MUX2_X1 U15949 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14663), .S(n16358), .Z(
        P2_U3519) );
  NAND2_X1 U15950 ( .A1(n14612), .A2(n16348), .ZN(n14615) );
  NAND3_X1 U15951 ( .A1(n14615), .A2(n14614), .A3(n14613), .ZN(n14664) );
  MUX2_X1 U15952 ( .A(n14664), .B(P2_REG1_REG_19__SCAN_IN), .S(n16357), .Z(
        n14616) );
  INV_X1 U15953 ( .A(n14616), .ZN(n14617) );
  OAI21_X1 U15954 ( .B1(n14667), .B2(n14631), .A(n14617), .ZN(P2_U3518) );
  OAI21_X1 U15955 ( .B1(n14619), .B2(n16353), .A(n14618), .ZN(n14620) );
  AOI21_X1 U15956 ( .B1(n14621), .B2(n13099), .A(n14620), .ZN(n14622) );
  NAND2_X1 U15957 ( .A1(n14623), .A2(n14622), .ZN(n14669) );
  MUX2_X1 U15958 ( .A(n14669), .B(P2_REG1_REG_18__SCAN_IN), .S(n16357), .Z(
        P2_U3517) );
  NAND2_X1 U15959 ( .A1(n14624), .A2(n16348), .ZN(n14628) );
  AND2_X1 U15960 ( .A1(n14626), .A2(n14625), .ZN(n14627) );
  AND2_X1 U15961 ( .A1(n14628), .A2(n14627), .ZN(n14670) );
  MUX2_X1 U15962 ( .A(n14629), .B(n14670), .S(n16358), .Z(n14630) );
  OAI21_X1 U15963 ( .B1(n14674), .B2(n14631), .A(n14630), .ZN(P2_U3516) );
  AOI21_X1 U15964 ( .B1(n16170), .B2(n14633), .A(n14632), .ZN(n14634) );
  OAI211_X1 U15965 ( .C1(n9885), .C2(n14636), .A(n14635), .B(n14634), .ZN(
        n14675) );
  MUX2_X1 U15966 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14675), .S(n16358), .Z(
        P2_U3515) );
  MUX2_X1 U15967 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n14637), .S(n16358), .Z(
        P2_U3499) );
  INV_X1 U15968 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n14639) );
  MUX2_X1 U15969 ( .A(n14639), .B(n14638), .S(n14668), .Z(n14640) );
  OAI21_X1 U15970 ( .B1(n14641), .B2(n14673), .A(n14640), .ZN(P2_U3498) );
  MUX2_X1 U15971 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n14642), .S(n14668), .Z(
        n14643) );
  INV_X1 U15972 ( .A(n14643), .ZN(n14644) );
  OAI21_X1 U15973 ( .B1(n14645), .B2(n14673), .A(n14644), .ZN(P2_U3497) );
  MUX2_X1 U15974 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n14647), .S(n14668), .Z(
        P2_U3495) );
  MUX2_X1 U15975 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14648), .S(n14668), .Z(
        P2_U3494) );
  MUX2_X1 U15976 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14649), .S(n14668), .Z(
        P2_U3493) );
  INV_X1 U15977 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n14651) );
  MUX2_X1 U15978 ( .A(n14651), .B(n14650), .S(n14668), .Z(n14652) );
  OAI21_X1 U15979 ( .B1(n14653), .B2(n14673), .A(n14652), .ZN(P2_U3492) );
  INV_X1 U15980 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n14655) );
  MUX2_X1 U15981 ( .A(n14655), .B(n14654), .S(n14668), .Z(n14656) );
  OAI21_X1 U15982 ( .B1(n14657), .B2(n14673), .A(n14656), .ZN(P2_U3491) );
  INV_X1 U15983 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n14659) );
  MUX2_X1 U15984 ( .A(n14659), .B(n14658), .S(n14668), .Z(n14660) );
  OAI21_X1 U15985 ( .B1(n8265), .B2(n14673), .A(n14660), .ZN(P2_U3490) );
  MUX2_X1 U15986 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14661), .S(n14668), .Z(
        P2_U3489) );
  MUX2_X1 U15987 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14662), .S(n14668), .Z(
        P2_U3488) );
  MUX2_X1 U15988 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14663), .S(n14668), .Z(
        P2_U3487) );
  MUX2_X1 U15989 ( .A(n14664), .B(P2_REG0_REG_19__SCAN_IN), .S(n16359), .Z(
        n14665) );
  INV_X1 U15990 ( .A(n14665), .ZN(n14666) );
  OAI21_X1 U15991 ( .B1(n14667), .B2(n14673), .A(n14666), .ZN(P2_U3486) );
  MUX2_X1 U15992 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14669), .S(n14668), .Z(
        P2_U3484) );
  INV_X1 U15993 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n14671) );
  MUX2_X1 U15994 ( .A(n14671), .B(n14670), .S(n14668), .Z(n14672) );
  OAI21_X1 U15995 ( .B1(n14674), .B2(n14673), .A(n14672), .ZN(P2_U3481) );
  MUX2_X1 U15996 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14675), .S(n14668), .Z(
        P2_U3478) );
  INV_X1 U15997 ( .A(n15236), .ZN(n14679) );
  NOR4_X1 U15998 ( .A1(n9636), .A2(P2_IR_REG_30__SCAN_IN), .A3(n14676), .A4(
        P2_U3088), .ZN(n14677) );
  AOI21_X1 U15999 ( .B1(n14685), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14677), 
        .ZN(n14678) );
  OAI21_X1 U16000 ( .B1(n14679), .B2(n14691), .A(n14678), .ZN(P2_U3296) );
  INV_X1 U16001 ( .A(n14681), .ZN(n15242) );
  OAI222_X1 U16002 ( .A1(n14680), .A2(P2_U3088), .B1(n14691), .B2(n15242), 
        .C1(n14682), .C2(n14693), .ZN(P2_U3297) );
  INV_X1 U16003 ( .A(n14683), .ZN(n15246) );
  AOI21_X1 U16004 ( .B1(n14685), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n14684), 
        .ZN(n14686) );
  OAI21_X1 U16005 ( .B1(n15246), .B2(n14691), .A(n14686), .ZN(P2_U3299) );
  OAI222_X1 U16006 ( .A1(n14688), .A2(P2_U3088), .B1(n14691), .B2(n15255), 
        .C1(n14687), .C2(n14693), .ZN(P2_U3301) );
  INV_X1 U16007 ( .A(n14689), .ZN(n15259) );
  OAI222_X1 U16008 ( .A1(n14693), .A2(n14692), .B1(n14691), .B2(n15259), .C1(
        n14690), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U16009 ( .A(n14694), .ZN(n14695) );
  MUX2_X1 U16010 ( .A(n14695), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XOR2_X1 U16011 ( .A(n14697), .B(n14696), .Z(n14704) );
  INV_X1 U16012 ( .A(n14944), .ZN(n14701) );
  OAI22_X1 U16013 ( .A1(n14699), .A2(n14787), .B1(n14698), .B2(n14785), .ZN(
        n15118) );
  AOI22_X1 U16014 ( .A1(n14821), .A2(n15118), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14700) );
  OAI21_X1 U16015 ( .B1(n14701), .B2(n14824), .A(n14700), .ZN(n14702) );
  AOI21_X1 U16016 ( .B1(n15119), .B2(n14826), .A(n14702), .ZN(n14703) );
  OAI21_X1 U16017 ( .B1(n14704), .B2(n14829), .A(n14703), .ZN(P1_U3214) );
  INV_X1 U16018 ( .A(n14705), .ZN(n15212) );
  OAI21_X1 U16019 ( .B1(n14707), .B2(n7601), .A(n14706), .ZN(n14708) );
  NAND2_X1 U16020 ( .A1(n14708), .A2(n14796), .ZN(n14712) );
  NAND2_X1 U16021 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14898)
         );
  OAI21_X1 U16022 ( .B1(n14809), .B2(n15211), .A(n14898), .ZN(n14709) );
  AOI21_X1 U16023 ( .B1(n14710), .B2(n14811), .A(n14709), .ZN(n14711) );
  OAI211_X1 U16024 ( .C1(n15212), .C2(n14804), .A(n14712), .B(n14711), .ZN(
        P1_U3215) );
  XOR2_X1 U16025 ( .A(n14713), .B(n7445), .Z(n14720) );
  INV_X1 U16026 ( .A(n15001), .ZN(n14717) );
  OAI22_X1 U16027 ( .A1(n14715), .A2(n14785), .B1(n14714), .B2(n14787), .ZN(
        n15146) );
  AOI22_X1 U16028 ( .A1(n15146), .A2(n14821), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14716) );
  OAI21_X1 U16029 ( .B1(n14717), .B2(n14824), .A(n14716), .ZN(n14718) );
  AOI21_X1 U16030 ( .B1(n15147), .B2(n14826), .A(n14718), .ZN(n14719) );
  OAI21_X1 U16031 ( .B1(n14720), .B2(n14829), .A(n14719), .ZN(P1_U3216) );
  XOR2_X1 U16032 ( .A(n14721), .B(n14722), .Z(n14728) );
  AND2_X1 U16033 ( .A1(n14843), .A2(n14806), .ZN(n14723) );
  AOI21_X1 U16034 ( .B1(n14841), .B2(n14799), .A(n14723), .ZN(n15175) );
  NAND2_X1 U16035 ( .A1(n14811), .A2(n15062), .ZN(n14725) );
  OAI211_X1 U16036 ( .C1(n15175), .C2(n14809), .A(n14725), .B(n14724), .ZN(
        n14726) );
  AOI21_X1 U16037 ( .B1(n15174), .B2(n14826), .A(n14726), .ZN(n14727) );
  OAI21_X1 U16038 ( .B1(n14728), .B2(n14829), .A(n14727), .ZN(P1_U3219) );
  AOI21_X1 U16039 ( .B1(n14731), .B2(n14730), .A(n14729), .ZN(n14737) );
  NOR2_X1 U16040 ( .A1(n14824), .A2(n15031), .ZN(n14735) );
  AND2_X1 U16041 ( .A1(n14841), .A2(n14806), .ZN(n14732) );
  AOI21_X1 U16042 ( .B1(n14839), .B2(n14807), .A(n14732), .ZN(n15160) );
  OAI22_X1 U16043 ( .A1(n15160), .A2(n14809), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14733), .ZN(n14734) );
  AOI211_X1 U16044 ( .C1(n15159), .C2(n14826), .A(n14735), .B(n14734), .ZN(
        n14736) );
  OAI21_X1 U16045 ( .B1(n14737), .B2(n14829), .A(n14736), .ZN(P1_U3223) );
  XOR2_X1 U16046 ( .A(n14739), .B(n14738), .Z(n14744) );
  AOI22_X1 U16047 ( .A1(n14806), .A2(n14837), .B1(n14835), .B2(n14799), .ZN(
        n15131) );
  OAI22_X1 U16048 ( .A1(n14809), .A2(n15131), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14740), .ZN(n14741) );
  AOI21_X1 U16049 ( .B1(n14973), .B2(n14811), .A(n14741), .ZN(n14743) );
  NAND2_X1 U16050 ( .A1(n14972), .A2(n14826), .ZN(n14742) );
  OAI211_X1 U16051 ( .C1(n14744), .C2(n14829), .A(n14743), .B(n14742), .ZN(
        P1_U3225) );
  INV_X1 U16052 ( .A(n14745), .ZN(n15196) );
  OAI21_X1 U16053 ( .B1(n14748), .B2(n14747), .A(n14746), .ZN(n14749) );
  NAND2_X1 U16054 ( .A1(n14749), .A2(n14796), .ZN(n14755) );
  INV_X1 U16055 ( .A(n14750), .ZN(n14753) );
  OAI21_X1 U16056 ( .B1(n14809), .B2(n15195), .A(n14751), .ZN(n14752) );
  AOI21_X1 U16057 ( .B1(n14753), .B2(n14811), .A(n14752), .ZN(n14754) );
  OAI211_X1 U16058 ( .C1(n15196), .C2(n14804), .A(n14755), .B(n14754), .ZN(
        P1_U3226) );
  INV_X1 U16059 ( .A(n14756), .ZN(n14761) );
  AOI21_X1 U16060 ( .B1(n14758), .B2(n14760), .A(n14757), .ZN(n14759) );
  AOI21_X1 U16061 ( .B1(n14761), .B2(n14760), .A(n14759), .ZN(n14767) );
  NAND2_X1 U16062 ( .A1(n14821), .A2(n15189), .ZN(n14762) );
  OAI211_X1 U16063 ( .C1(n14824), .C2(n14764), .A(n14763), .B(n14762), .ZN(
        n14765) );
  AOI21_X1 U16064 ( .B1(n15190), .B2(n14826), .A(n14765), .ZN(n14766) );
  OAI21_X1 U16065 ( .B1(n14767), .B2(n14829), .A(n14766), .ZN(P1_U3228) );
  XOR2_X1 U16066 ( .A(n14769), .B(n14768), .Z(n14775) );
  AND2_X1 U16067 ( .A1(n14836), .A2(n14807), .ZN(n14770) );
  AOI21_X1 U16068 ( .B1(n14838), .B2(n14806), .A(n14770), .ZN(n14987) );
  OAI22_X1 U16069 ( .A1(n14987), .A2(n14809), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14771), .ZN(n14772) );
  AOI21_X1 U16070 ( .B1(n14993), .B2(n14811), .A(n14772), .ZN(n14774) );
  NAND2_X1 U16071 ( .A1(n15138), .A2(n14826), .ZN(n14773) );
  OAI211_X1 U16072 ( .C1(n14775), .C2(n14829), .A(n14774), .B(n14773), .ZN(
        P1_U3229) );
  OAI211_X1 U16073 ( .C1(n14778), .C2(n14777), .A(n14776), .B(n14796), .ZN(
        n14782) );
  AOI22_X1 U16074 ( .A1(n14840), .A2(n14807), .B1(n14806), .B2(n14842), .ZN(
        n15167) );
  OAI22_X1 U16075 ( .A1(n15167), .A2(n14809), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14779), .ZN(n14780) );
  AOI21_X1 U16076 ( .B1(n15044), .B2(n14811), .A(n14780), .ZN(n14781) );
  OAI211_X1 U16077 ( .C1(n15169), .C2(n14804), .A(n14782), .B(n14781), .ZN(
        P1_U3233) );
  AOI21_X1 U16078 ( .B1(n8051), .B2(n14784), .A(n14783), .ZN(n14792) );
  OAI22_X1 U16079 ( .A1(n14788), .A2(n14787), .B1(n14786), .B2(n14785), .ZN(
        n15154) );
  AOI22_X1 U16080 ( .A1(n15154), .A2(n14821), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14789) );
  OAI21_X1 U16081 ( .B1(n15017), .B2(n14824), .A(n14789), .ZN(n14790) );
  AOI21_X1 U16082 ( .B1(n15155), .B2(n14826), .A(n14790), .ZN(n14791) );
  OAI21_X1 U16083 ( .B1(n14792), .B2(n14829), .A(n14791), .ZN(P1_U3235) );
  INV_X1 U16084 ( .A(n15184), .ZN(n15085) );
  OAI21_X1 U16085 ( .B1(n14795), .B2(n14794), .A(n14793), .ZN(n14797) );
  NAND2_X1 U16086 ( .A1(n14797), .A2(n14796), .ZN(n14803) );
  INV_X1 U16087 ( .A(n14798), .ZN(n15082) );
  AOI22_X1 U16088 ( .A1(n14842), .A2(n14799), .B1(n14806), .B2(n14844), .ZN(
        n15072) );
  OAI21_X1 U16089 ( .B1(n14809), .B2(n15072), .A(n14800), .ZN(n14801) );
  AOI21_X1 U16090 ( .B1(n15082), .B2(n14811), .A(n14801), .ZN(n14802) );
  OAI211_X1 U16091 ( .C1(n15085), .C2(n14804), .A(n14803), .B(n14802), .ZN(
        P1_U3238) );
  AOI22_X1 U16092 ( .A1(n14807), .A2(n14834), .B1(n14836), .B2(n14806), .ZN(
        n15124) );
  OAI22_X1 U16093 ( .A1(n14809), .A2(n15124), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14808), .ZN(n14810) );
  AOI21_X1 U16094 ( .B1(n14959), .B2(n14811), .A(n14810), .ZN(n14814) );
  NAND2_X1 U16095 ( .A1(n14812), .A2(n14826), .ZN(n14813) );
  INV_X1 U16096 ( .A(n14815), .ZN(n14820) );
  AOI21_X1 U16097 ( .B1(n14817), .B2(n14819), .A(n14816), .ZN(n14818) );
  AOI21_X1 U16098 ( .B1(n14820), .B2(n14819), .A(n14818), .ZN(n14830) );
  NAND2_X1 U16099 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n15855)
         );
  NAND2_X1 U16100 ( .A1(n14821), .A2(n15203), .ZN(n14822) );
  OAI211_X1 U16101 ( .C1(n14824), .C2(n14823), .A(n15855), .B(n14822), .ZN(
        n14825) );
  AOI21_X1 U16102 ( .B1(n14827), .B2(n14826), .A(n14825), .ZN(n14828) );
  OAI21_X1 U16103 ( .B1(n14830), .B2(n14829), .A(n14828), .ZN(P1_U3241) );
  MUX2_X1 U16104 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14831), .S(n14861), .Z(
        P1_U3590) );
  MUX2_X1 U16105 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14832), .S(n14861), .Z(
        P1_U3589) );
  MUX2_X1 U16106 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14833), .S(n14861), .Z(
        P1_U3588) );
  MUX2_X1 U16107 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14834), .S(n14861), .Z(
        P1_U3587) );
  MUX2_X1 U16108 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14835), .S(n14861), .Z(
        P1_U3586) );
  MUX2_X1 U16109 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14836), .S(n14861), .Z(
        P1_U3585) );
  MUX2_X1 U16110 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14837), .S(n14861), .Z(
        P1_U3584) );
  MUX2_X1 U16111 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14838), .S(n14861), .Z(
        P1_U3583) );
  MUX2_X1 U16112 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14839), .S(n14861), .Z(
        P1_U3582) );
  MUX2_X1 U16113 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14840), .S(n14861), .Z(
        P1_U3581) );
  MUX2_X1 U16114 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14841), .S(n14861), .Z(
        P1_U3580) );
  MUX2_X1 U16115 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14842), .S(n14861), .Z(
        P1_U3579) );
  MUX2_X1 U16116 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14843), .S(n14861), .Z(
        P1_U3578) );
  MUX2_X1 U16117 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14844), .S(n14861), .Z(
        P1_U3577) );
  MUX2_X1 U16118 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14845), .S(n14861), .Z(
        P1_U3576) );
  MUX2_X1 U16119 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14846), .S(n14861), .Z(
        P1_U3575) );
  MUX2_X1 U16120 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14847), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16121 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14848), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16122 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14849), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16123 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14850), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16124 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14851), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16125 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14852), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16126 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14853), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16127 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14854), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16128 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14855), .S(n14861), .Z(
        P1_U3566) );
  MUX2_X1 U16129 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14856), .S(n14861), .Z(
        P1_U3565) );
  MUX2_X1 U16130 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14857), .S(n14861), .Z(
        P1_U3564) );
  MUX2_X1 U16131 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14858), .S(n14861), .Z(
        P1_U3563) );
  MUX2_X1 U16132 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14859), .S(n14861), .Z(
        P1_U3562) );
  MUX2_X1 U16133 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14860), .S(n14861), .Z(
        P1_U3561) );
  MUX2_X1 U16134 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14862), .S(n14861), .Z(
        P1_U3560) );
  OAI211_X1 U16135 ( .C1(n14865), .C2(n14864), .A(n7422), .B(n14863), .ZN(
        n14875) );
  AOI22_X1 U16136 ( .A1(n14866), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14874) );
  MUX2_X1 U16137 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9914), .S(n14867), .Z(
        n14868) );
  OAI21_X1 U16138 ( .B1(n16035), .B2(n8323), .A(n14868), .ZN(n14869) );
  NAND3_X1 U16139 ( .A1(n16018), .A2(n14870), .A3(n14869), .ZN(n14873) );
  NAND2_X1 U16140 ( .A1(n14900), .A2(n14871), .ZN(n14872) );
  NAND4_X1 U16141 ( .A1(n14875), .A2(n14874), .A3(n14873), .A4(n14872), .ZN(
        P1_U3244) );
  NAND3_X1 U16142 ( .A1(n14878), .A2(n14877), .A3(n14876), .ZN(n14879) );
  NAND3_X1 U16143 ( .A1(n7422), .A2(n14880), .A3(n14879), .ZN(n14893) );
  INV_X1 U16144 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n15739) );
  OAI21_X1 U16145 ( .B1(n16028), .B2(n15739), .A(n14881), .ZN(n14882) );
  AOI21_X1 U16146 ( .B1(n14883), .B2(n14900), .A(n14882), .ZN(n14892) );
  MUX2_X1 U16147 ( .A(n14884), .B(P1_REG1_REG_7__SCAN_IN), .S(n14883), .Z(
        n14887) );
  INV_X1 U16148 ( .A(n14885), .ZN(n14886) );
  NAND2_X1 U16149 ( .A1(n14887), .A2(n14886), .ZN(n14889) );
  OAI211_X1 U16150 ( .C1(n14890), .C2(n14889), .A(n16018), .B(n14888), .ZN(
        n14891) );
  NAND3_X1 U16151 ( .A1(n14893), .A2(n14892), .A3(n14891), .ZN(P1_U3250) );
  OAI21_X1 U16152 ( .B1(n14896), .B2(n14895), .A(n14894), .ZN(n14897) );
  NAND2_X1 U16153 ( .A1(n14897), .A2(n16018), .ZN(n14910) );
  INV_X1 U16154 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15699) );
  OAI21_X1 U16155 ( .B1(n16028), .B2(n15699), .A(n14898), .ZN(n14899) );
  AOI21_X1 U16156 ( .B1(n14901), .B2(n14900), .A(n14899), .ZN(n14909) );
  MUX2_X1 U16157 ( .A(n11186), .B(P1_REG2_REG_14__SCAN_IN), .S(n14901), .Z(
        n14904) );
  INV_X1 U16158 ( .A(n14902), .ZN(n14903) );
  NAND2_X1 U16159 ( .A1(n14904), .A2(n14903), .ZN(n14906) );
  OAI211_X1 U16160 ( .C1(n14907), .C2(n14906), .A(n14905), .B(n7422), .ZN(
        n14908) );
  NAND3_X1 U16161 ( .A1(n14910), .A2(n14909), .A3(n14908), .ZN(P1_U3257) );
  NOR2_X1 U16162 ( .A1(n16086), .A2(n14912), .ZN(n14915) );
  NAND2_X1 U16163 ( .A1(n14914), .A2(n14913), .ZN(n15103) );
  NOR2_X1 U16164 ( .A1(n16347), .A2(n15103), .ZN(n14920) );
  AOI211_X1 U16165 ( .C1(n15101), .C2(n16337), .A(n14915), .B(n14920), .ZN(
        n14916) );
  OAI21_X1 U16166 ( .B1(n15102), .B2(n15051), .A(n14916), .ZN(P1_U3263) );
  OAI211_X1 U16167 ( .C1(n15105), .C2(n14918), .A(n14917), .B(n16322), .ZN(
        n15104) );
  NOR2_X1 U16168 ( .A1(n15105), .A2(n16163), .ZN(n14919) );
  AOI211_X1 U16169 ( .C1(n16347), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14920), 
        .B(n14919), .ZN(n14921) );
  OAI21_X1 U16170 ( .B1(n15051), .B2(n15104), .A(n14921), .ZN(P1_U3264) );
  INV_X1 U16171 ( .A(n14943), .ZN(n14924) );
  AOI21_X1 U16172 ( .B1(n15115), .B2(n14924), .A(n16142), .ZN(n14925) );
  AND2_X1 U16173 ( .A1(n14926), .A2(n14925), .ZN(n15114) );
  INV_X1 U16174 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n14930) );
  NAND2_X1 U16175 ( .A1(n15115), .A2(n16337), .ZN(n14929) );
  NAND2_X1 U16176 ( .A1(n16336), .A2(n14927), .ZN(n14928) );
  OAI211_X1 U16177 ( .C1(n16159), .C2(n14930), .A(n14929), .B(n14928), .ZN(
        n14931) );
  AOI21_X1 U16178 ( .B1(n15114), .B2(n16341), .A(n14931), .ZN(n14938) );
  OAI211_X1 U16179 ( .C1(n14934), .C2(n14933), .A(n14932), .B(n16194), .ZN(
        n14936) );
  NAND2_X1 U16180 ( .A1(n15113), .A2(n16159), .ZN(n14937) );
  OAI211_X1 U16181 ( .C1(n15116), .C2(n15088), .A(n14938), .B(n14937), .ZN(
        P1_U3265) );
  AOI21_X1 U16182 ( .B1(n14949), .B2(n14940), .A(n14939), .ZN(n15123) );
  NAND2_X1 U16183 ( .A1(n15119), .A2(n14958), .ZN(n14941) );
  NAND2_X1 U16184 ( .A1(n14941), .A2(n16322), .ZN(n14942) );
  NOR2_X1 U16185 ( .A1(n14943), .A2(n14942), .ZN(n15117) );
  AOI22_X1 U16186 ( .A1(n16086), .A2(n15118), .B1(n16336), .B2(n14944), .ZN(
        n14946) );
  NAND2_X1 U16187 ( .A1(n16347), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n14945) );
  OAI211_X1 U16188 ( .C1(n14947), .C2(n16163), .A(n14946), .B(n14945), .ZN(
        n14948) );
  AOI21_X1 U16189 ( .B1(n15117), .B2(n16341), .A(n14948), .ZN(n14952) );
  XNOR2_X1 U16190 ( .A(n14950), .B(n14949), .ZN(n15120) );
  NAND2_X1 U16191 ( .A1(n15120), .A2(n15090), .ZN(n14951) );
  OAI211_X1 U16192 ( .C1(n15123), .C2(n15088), .A(n14952), .B(n14951), .ZN(
        P1_U3266) );
  XNOR2_X1 U16193 ( .A(n14953), .B(n14955), .ZN(n15130) );
  OAI21_X1 U16194 ( .B1(n14956), .B2(n14955), .A(n14954), .ZN(n14957) );
  INV_X1 U16195 ( .A(n14957), .ZN(n15128) );
  OAI211_X1 U16196 ( .C1(n15126), .C2(n7461), .A(n16322), .B(n14958), .ZN(
        n15125) );
  INV_X1 U16197 ( .A(n14959), .ZN(n14960) );
  OAI22_X1 U16198 ( .A1(n16347), .A2(n15124), .B1(n14960), .B2(n16161), .ZN(
        n14962) );
  NOR2_X1 U16199 ( .A1(n15126), .A2(n16163), .ZN(n14961) );
  AOI211_X1 U16200 ( .C1(n16347), .C2(P1_REG2_REG_26__SCAN_IN), .A(n14962), 
        .B(n14961), .ZN(n14963) );
  OAI21_X1 U16201 ( .B1(n15051), .B2(n15125), .A(n14963), .ZN(n14964) );
  AOI21_X1 U16202 ( .B1(n15128), .B2(n15058), .A(n14964), .ZN(n14965) );
  OAI21_X1 U16203 ( .B1(n15130), .B2(n15070), .A(n14965), .ZN(P1_U3267) );
  OAI21_X1 U16204 ( .B1(n14968), .B2(n14967), .A(n14966), .ZN(n15137) );
  OAI21_X1 U16205 ( .B1(n14971), .B2(n14970), .A(n14969), .ZN(n15135) );
  AOI211_X1 U16206 ( .C1(n14972), .C2(n14991), .A(n16142), .B(n7461), .ZN(
        n15134) );
  NAND2_X1 U16207 ( .A1(n15134), .A2(n16341), .ZN(n14977) );
  INV_X1 U16208 ( .A(n14973), .ZN(n14974) );
  OAI22_X1 U16209 ( .A1(n16347), .A2(n15131), .B1(n14974), .B2(n16161), .ZN(
        n14975) );
  AOI21_X1 U16210 ( .B1(P1_REG2_REG_25__SCAN_IN), .B2(n16347), .A(n14975), 
        .ZN(n14976) );
  OAI211_X1 U16211 ( .C1(n15132), .C2(n16163), .A(n14977), .B(n14976), .ZN(
        n14978) );
  AOI21_X1 U16212 ( .B1(n15135), .B2(n15090), .A(n14978), .ZN(n14979) );
  OAI21_X1 U16213 ( .B1(n15137), .B2(n15054), .A(n14979), .ZN(P1_U3268) );
  AND2_X1 U16214 ( .A1(n14981), .A2(n14980), .ZN(n14983) );
  NAND2_X1 U16215 ( .A1(n14985), .A2(n14984), .ZN(n14986) );
  NAND2_X1 U16216 ( .A1(n14986), .A2(n16194), .ZN(n14988) );
  OAI21_X1 U16217 ( .B1(n14989), .B2(n14988), .A(n14987), .ZN(n14990) );
  AOI21_X1 U16218 ( .B1(n15142), .B2(n16372), .A(n14990), .ZN(n15144) );
  OAI211_X1 U16219 ( .C1(n14992), .C2(n15000), .A(n16322), .B(n14991), .ZN(
        n15140) );
  AOI22_X1 U16220 ( .A1(n16347), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14993), 
        .B2(n16336), .ZN(n14995) );
  NAND2_X1 U16221 ( .A1(n15138), .A2(n16337), .ZN(n14994) );
  OAI211_X1 U16222 ( .C1(n15140), .C2(n15051), .A(n14995), .B(n14994), .ZN(
        n14996) );
  AOI21_X1 U16223 ( .B1(n15142), .B2(n16342), .A(n14996), .ZN(n14997) );
  OAI21_X1 U16224 ( .B1(n15144), .B2(n16347), .A(n14997), .ZN(P1_U3269) );
  INV_X1 U16225 ( .A(n15007), .ZN(n14999) );
  OAI21_X1 U16226 ( .B1(n7590), .B2(n14999), .A(n14998), .ZN(n15151) );
  AOI211_X1 U16227 ( .C1(n15147), .C2(n15015), .A(n16142), .B(n15000), .ZN(
        n15145) );
  NAND2_X1 U16228 ( .A1(n15147), .A2(n16337), .ZN(n15003) );
  AOI22_X1 U16229 ( .A1(n15146), .A2(n16159), .B1(n15001), .B2(n16336), .ZN(
        n15002) );
  OAI211_X1 U16230 ( .C1(n16159), .C2(n15004), .A(n15003), .B(n15002), .ZN(
        n15005) );
  AOI21_X1 U16231 ( .B1(n15145), .B2(n16341), .A(n15005), .ZN(n15010) );
  OAI21_X1 U16232 ( .B1(n15008), .B2(n15007), .A(n15006), .ZN(n15148) );
  NAND2_X1 U16233 ( .A1(n15148), .A2(n15090), .ZN(n15009) );
  OAI211_X1 U16234 ( .C1(n15151), .C2(n15054), .A(n15010), .B(n15009), .ZN(
        P1_U3270) );
  XNOR2_X1 U16235 ( .A(n15012), .B(n15011), .ZN(n15158) );
  XNOR2_X1 U16236 ( .A(n15014), .B(n15013), .ZN(n15152) );
  NAND2_X1 U16237 ( .A1(n15152), .A2(n15058), .ZN(n15024) );
  INV_X1 U16238 ( .A(n15015), .ZN(n15016) );
  AOI211_X1 U16239 ( .C1(n15155), .C2(n15029), .A(n16142), .B(n15016), .ZN(
        n15153) );
  OAI22_X1 U16240 ( .A1(n16086), .A2(n15018), .B1(n15017), .B2(n16161), .ZN(
        n15019) );
  AOI21_X1 U16241 ( .B1(n15154), .B2(n16159), .A(n15019), .ZN(n15020) );
  OAI21_X1 U16242 ( .B1(n15021), .B2(n16163), .A(n15020), .ZN(n15022) );
  AOI21_X1 U16243 ( .B1(n15153), .B2(n16341), .A(n15022), .ZN(n15023) );
  OAI211_X1 U16244 ( .C1(n15158), .C2(n15070), .A(n15024), .B(n15023), .ZN(
        P1_U3271) );
  XNOR2_X1 U16245 ( .A(n15026), .B(n15025), .ZN(n15166) );
  OAI21_X1 U16246 ( .B1(n7587), .B2(n15028), .A(n15027), .ZN(n15164) );
  AOI21_X1 U16247 ( .B1(n15043), .B2(n15159), .A(n16142), .ZN(n15030) );
  NAND2_X1 U16248 ( .A1(n15030), .A2(n15029), .ZN(n15161) );
  NOR2_X1 U16249 ( .A1(n15161), .A2(n15051), .ZN(n15037) );
  NAND2_X1 U16250 ( .A1(n15159), .A2(n16337), .ZN(n15034) );
  OAI22_X1 U16251 ( .A1(n15160), .A2(n16347), .B1(n15031), .B2(n16161), .ZN(
        n15032) );
  INV_X1 U16252 ( .A(n15032), .ZN(n15033) );
  OAI211_X1 U16253 ( .C1(n16159), .C2(n15035), .A(n15034), .B(n15033), .ZN(
        n15036) );
  AOI211_X1 U16254 ( .C1(n15164), .C2(n15058), .A(n15037), .B(n15036), .ZN(
        n15038) );
  OAI21_X1 U16255 ( .B1(n15070), .B2(n15166), .A(n15038), .ZN(P1_U3272) );
  OAI21_X1 U16256 ( .B1(n7584), .B2(n15042), .A(n15039), .ZN(n15173) );
  AOI21_X1 U16257 ( .B1(n15042), .B2(n15041), .A(n8326), .ZN(n15171) );
  OAI211_X1 U16258 ( .C1(n15061), .C2(n15169), .A(n15043), .B(n16322), .ZN(
        n15168) );
  INV_X1 U16259 ( .A(n15167), .ZN(n15045) );
  AOI22_X1 U16260 ( .A1(n15045), .A2(n16159), .B1(n15044), .B2(n16336), .ZN(
        n15046) );
  OAI21_X1 U16261 ( .B1(n15047), .B2(n16159), .A(n15046), .ZN(n15048) );
  AOI21_X1 U16262 ( .B1(n15049), .B2(n16337), .A(n15048), .ZN(n15050) );
  OAI21_X1 U16263 ( .B1(n15168), .B2(n15051), .A(n15050), .ZN(n15052) );
  AOI21_X1 U16264 ( .B1(n15171), .B2(n15090), .A(n15052), .ZN(n15053) );
  OAI21_X1 U16265 ( .B1(n15054), .B2(n15173), .A(n15053), .ZN(P1_U3273) );
  XOR2_X1 U16266 ( .A(n15056), .B(n15055), .Z(n15181) );
  XNOR2_X1 U16267 ( .A(n15057), .B(n15056), .ZN(n15179) );
  NAND2_X1 U16268 ( .A1(n15179), .A2(n15058), .ZN(n15069) );
  NAND2_X1 U16269 ( .A1(n15079), .A2(n15174), .ZN(n15059) );
  NAND2_X1 U16270 ( .A1(n15059), .A2(n16322), .ZN(n15060) );
  NOR2_X1 U16271 ( .A1(n15061), .A2(n15060), .ZN(n15178) );
  NAND2_X1 U16272 ( .A1(n15174), .A2(n16337), .ZN(n15065) );
  INV_X1 U16273 ( .A(n15175), .ZN(n15063) );
  AOI22_X1 U16274 ( .A1(n15063), .A2(n16159), .B1(n15062), .B2(n16336), .ZN(
        n15064) );
  OAI211_X1 U16275 ( .C1(n16159), .C2(n15066), .A(n15065), .B(n15064), .ZN(
        n15067) );
  AOI21_X1 U16276 ( .B1(n15178), .B2(n16341), .A(n15067), .ZN(n15068) );
  OAI211_X1 U16277 ( .C1(n15181), .C2(n15070), .A(n15069), .B(n15068), .ZN(
        P1_U3274) );
  OAI21_X1 U16278 ( .B1(n7585), .B2(n15076), .A(n15071), .ZN(n15182) );
  INV_X1 U16279 ( .A(n15072), .ZN(n15078) );
  INV_X1 U16280 ( .A(n15073), .ZN(n15074) );
  AOI211_X1 U16281 ( .C1(n15076), .C2(n15075), .A(n16379), .B(n15074), .ZN(
        n15077) );
  AOI211_X1 U16282 ( .C1(n16372), .C2(n15182), .A(n15078), .B(n15077), .ZN(
        n15186) );
  INV_X1 U16283 ( .A(n15079), .ZN(n15080) );
  AOI211_X1 U16284 ( .C1(n15184), .C2(n15081), .A(n16142), .B(n15080), .ZN(
        n15183) );
  NAND2_X1 U16285 ( .A1(n15183), .A2(n16341), .ZN(n15084) );
  AOI22_X1 U16286 ( .A1(n16347), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n15082), 
        .B2(n16336), .ZN(n15083) );
  OAI211_X1 U16287 ( .C1(n15085), .C2(n16163), .A(n15084), .B(n15083), .ZN(
        n15086) );
  AOI21_X1 U16288 ( .B1(n15182), .B2(n16342), .A(n15086), .ZN(n15087) );
  OAI21_X1 U16289 ( .B1(n15186), .B2(n16347), .A(n15087), .ZN(P1_U3275) );
  INV_X1 U16290 ( .A(n15088), .ZN(n15092) );
  AOI22_X1 U16291 ( .A1(n15092), .A2(n15091), .B1(n15090), .B2(n15089), .ZN(
        n15100) );
  MUX2_X1 U16292 ( .A(n15094), .B(n15093), .S(n16159), .Z(n15099) );
  AOI22_X1 U16293 ( .A1(n16337), .A2(n15095), .B1(n16336), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n15098) );
  NAND2_X1 U16294 ( .A1(n16341), .A2(n15096), .ZN(n15097) );
  NAND4_X1 U16295 ( .A1(n15100), .A2(n15099), .A3(n15098), .A4(n15097), .ZN(
        P1_U3291) );
  MUX2_X1 U16296 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15218), .S(n16387), .Z(
        P1_U3559) );
  OAI211_X1 U16297 ( .C1(n15105), .C2(n16378), .A(n15104), .B(n15103), .ZN(
        n15219) );
  MUX2_X1 U16298 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15219), .S(n16387), .Z(
        P1_U3558) );
  OAI211_X1 U16299 ( .C1(n15108), .C2(n16378), .A(n15107), .B(n15106), .ZN(
        n15109) );
  MUX2_X1 U16300 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n15220), .S(n16387), .Z(
        P1_U3557) );
  MUX2_X1 U16301 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15221), .S(n16387), .Z(
        P1_U3556) );
  AOI211_X1 U16302 ( .C1(n16366), .C2(n15119), .A(n15118), .B(n15117), .ZN(
        n15122) );
  NAND2_X1 U16303 ( .A1(n15120), .A2(n16194), .ZN(n15121) );
  OAI211_X1 U16304 ( .C1(n15123), .C2(n16190), .A(n15122), .B(n15121), .ZN(
        n15222) );
  MUX2_X1 U16305 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15222), .S(n16387), .Z(
        P1_U3555) );
  OAI211_X1 U16306 ( .C1(n15126), .C2(n16378), .A(n15125), .B(n15124), .ZN(
        n15127) );
  AOI21_X1 U16307 ( .B1(n15128), .B2(n16383), .A(n15127), .ZN(n15129) );
  OAI21_X1 U16308 ( .B1(n16379), .B2(n15130), .A(n15129), .ZN(n15223) );
  MUX2_X1 U16309 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15223), .S(n16387), .Z(
        P1_U3554) );
  OAI21_X1 U16310 ( .B1(n15132), .B2(n16378), .A(n15131), .ZN(n15133) );
  AOI211_X1 U16311 ( .C1(n15135), .C2(n16194), .A(n15134), .B(n15133), .ZN(
        n15136) );
  OAI21_X1 U16312 ( .B1(n15137), .B2(n16190), .A(n15136), .ZN(n15224) );
  MUX2_X1 U16313 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15224), .S(n16387), .Z(
        P1_U3553) );
  NAND2_X1 U16314 ( .A1(n15138), .A2(n16366), .ZN(n15139) );
  NAND2_X1 U16315 ( .A1(n15140), .A2(n15139), .ZN(n15141) );
  AOI21_X1 U16316 ( .B1(n15142), .B2(n16332), .A(n15141), .ZN(n15143) );
  NAND2_X1 U16317 ( .A1(n15144), .A2(n15143), .ZN(n15225) );
  MUX2_X1 U16318 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15225), .S(n16387), .Z(
        P1_U3552) );
  AOI211_X1 U16319 ( .C1(n16366), .C2(n15147), .A(n15146), .B(n15145), .ZN(
        n15150) );
  NAND2_X1 U16320 ( .A1(n15148), .A2(n16194), .ZN(n15149) );
  OAI211_X1 U16321 ( .C1(n15151), .C2(n16190), .A(n15150), .B(n15149), .ZN(
        n15226) );
  MUX2_X1 U16322 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15226), .S(n16387), .Z(
        P1_U3551) );
  NAND2_X1 U16323 ( .A1(n15152), .A2(n16383), .ZN(n15157) );
  AOI211_X1 U16324 ( .C1(n16366), .C2(n15155), .A(n15154), .B(n15153), .ZN(
        n15156) );
  OAI211_X1 U16325 ( .C1(n16379), .C2(n15158), .A(n15157), .B(n15156), .ZN(
        n15227) );
  MUX2_X1 U16326 ( .A(n15227), .B(P1_REG1_REG_22__SCAN_IN), .S(n16385), .Z(
        P1_U3550) );
  INV_X1 U16327 ( .A(n15159), .ZN(n15162) );
  OAI211_X1 U16328 ( .C1(n15162), .C2(n16378), .A(n15161), .B(n15160), .ZN(
        n15163) );
  AOI21_X1 U16329 ( .B1(n15164), .B2(n16383), .A(n15163), .ZN(n15165) );
  OAI21_X1 U16330 ( .B1(n16379), .B2(n15166), .A(n15165), .ZN(n15228) );
  MUX2_X1 U16331 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15228), .S(n16387), .Z(
        P1_U3549) );
  OAI211_X1 U16332 ( .C1(n15169), .C2(n16378), .A(n15168), .B(n15167), .ZN(
        n15170) );
  AOI21_X1 U16333 ( .B1(n15171), .B2(n16194), .A(n15170), .ZN(n15172) );
  OAI21_X1 U16334 ( .B1(n16190), .B2(n15173), .A(n15172), .ZN(n15229) );
  MUX2_X1 U16335 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15229), .S(n16387), .Z(
        P1_U3548) );
  NAND2_X1 U16336 ( .A1(n15174), .A2(n16366), .ZN(n15176) );
  NAND2_X1 U16337 ( .A1(n15176), .A2(n15175), .ZN(n15177) );
  AOI211_X1 U16338 ( .C1(n15179), .C2(n16383), .A(n15178), .B(n15177), .ZN(
        n15180) );
  OAI21_X1 U16339 ( .B1(n16379), .B2(n15181), .A(n15180), .ZN(n15230) );
  MUX2_X1 U16340 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15230), .S(n16387), .Z(
        P1_U3547) );
  INV_X1 U16341 ( .A(n15182), .ZN(n15187) );
  AOI21_X1 U16342 ( .B1(n16366), .B2(n15184), .A(n15183), .ZN(n15185) );
  OAI211_X1 U16343 ( .C1(n15187), .C2(n16369), .A(n15186), .B(n15185), .ZN(
        n15231) );
  MUX2_X1 U16344 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15231), .S(n16387), .Z(
        P1_U3546) );
  AOI211_X1 U16345 ( .C1(n16366), .C2(n15190), .A(n15189), .B(n15188), .ZN(
        n15193) );
  NAND2_X1 U16346 ( .A1(n15191), .A2(n16194), .ZN(n15192) );
  OAI211_X1 U16347 ( .C1(n15194), .C2(n16190), .A(n15193), .B(n15192), .ZN(
        n15232) );
  MUX2_X1 U16348 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15232), .S(n16387), .Z(
        P1_U3545) );
  OAI21_X1 U16349 ( .B1(n15196), .B2(n16378), .A(n15195), .ZN(n15197) );
  AOI21_X1 U16350 ( .B1(n15198), .B2(n16322), .A(n15197), .ZN(n15201) );
  NAND2_X1 U16351 ( .A1(n15199), .A2(n16194), .ZN(n15200) );
  OAI211_X1 U16352 ( .C1(n15202), .C2(n16190), .A(n15201), .B(n15200), .ZN(
        n15233) );
  MUX2_X1 U16353 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15233), .S(n16387), .Z(
        P1_U3544) );
  INV_X1 U16354 ( .A(n15203), .ZN(n15204) );
  OAI211_X1 U16355 ( .C1(n15206), .C2(n16378), .A(n15205), .B(n15204), .ZN(
        n15207) );
  AOI21_X1 U16356 ( .B1(n15208), .B2(n16383), .A(n15207), .ZN(n15209) );
  OAI21_X1 U16357 ( .B1(n16379), .B2(n15210), .A(n15209), .ZN(n15234) );
  MUX2_X1 U16358 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15234), .S(n16387), .Z(
        P1_U3543) );
  OAI21_X1 U16359 ( .B1(n15212), .B2(n16378), .A(n15211), .ZN(n15213) );
  AOI211_X1 U16360 ( .C1(n15215), .C2(n16383), .A(n15214), .B(n15213), .ZN(
        n15216) );
  OAI21_X1 U16361 ( .B1(n16379), .B2(n15217), .A(n15216), .ZN(n15235) );
  MUX2_X1 U16362 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15235), .S(n16387), .Z(
        P1_U3542) );
  MUX2_X1 U16363 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15218), .S(n16391), .Z(
        P1_U3527) );
  MUX2_X1 U16364 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15219), .S(n16391), .Z(
        P1_U3526) );
  MUX2_X1 U16365 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n15220), .S(n16391), .Z(
        P1_U3525) );
  MUX2_X1 U16366 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15222), .S(n16391), .Z(
        P1_U3523) );
  MUX2_X1 U16367 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15223), .S(n16391), .Z(
        P1_U3522) );
  MUX2_X1 U16368 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15224), .S(n16391), .Z(
        P1_U3521) );
  MUX2_X1 U16369 ( .A(n15225), .B(P1_REG0_REG_24__SCAN_IN), .S(n16388), .Z(
        P1_U3520) );
  MUX2_X1 U16370 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15226), .S(n16391), .Z(
        P1_U3519) );
  MUX2_X1 U16371 ( .A(n15227), .B(P1_REG0_REG_22__SCAN_IN), .S(n16388), .Z(
        P1_U3518) );
  MUX2_X1 U16372 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15228), .S(n16391), .Z(
        P1_U3517) );
  MUX2_X1 U16373 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15229), .S(n16391), .Z(
        P1_U3516) );
  MUX2_X1 U16374 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15230), .S(n16391), .Z(
        P1_U3515) );
  MUX2_X1 U16375 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15231), .S(n16391), .Z(
        P1_U3513) );
  MUX2_X1 U16376 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15232), .S(n16391), .Z(
        P1_U3510) );
  MUX2_X1 U16377 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15233), .S(n16391), .Z(
        P1_U3507) );
  MUX2_X1 U16378 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15234), .S(n16391), .Z(
        P1_U3504) );
  MUX2_X1 U16379 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15235), .S(n16391), .Z(
        P1_U3501) );
  NAND2_X1 U16380 ( .A1(n15236), .A2(n15248), .ZN(n15240) );
  NAND4_X1 U16381 ( .A1(n15238), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .A4(n15237), .ZN(n15239) );
  OAI211_X1 U16382 ( .C1(n15241), .C2(n15262), .A(n15240), .B(n15239), .ZN(
        P1_U3324) );
  OAI222_X1 U16383 ( .A1(n15262), .A2(n15244), .B1(P1_U3086), .B2(n15243), 
        .C1(n15260), .C2(n15242), .ZN(P1_U3325) );
  OAI222_X1 U16384 ( .A1(n15262), .A2(n15247), .B1(n15260), .B2(n15246), .C1(
        n15245), .C2(P1_U3086), .ZN(P1_U3327) );
  NAND2_X1 U16385 ( .A1(n15249), .A2(n15248), .ZN(n15251) );
  OAI211_X1 U16386 ( .C1(n15252), .C2(n15262), .A(n15251), .B(n15250), .ZN(
        P1_U3328) );
  INV_X1 U16387 ( .A(n15253), .ZN(n15256) );
  OAI222_X1 U16388 ( .A1(n15256), .A2(P1_U3086), .B1(n15260), .B2(n15255), 
        .C1(n15254), .C2(n15262), .ZN(P1_U3329) );
  OAI222_X1 U16389 ( .A1(n15262), .A2(n15261), .B1(n15260), .B2(n15259), .C1(
        n15258), .C2(P1_U3086), .ZN(P1_U3330) );
  MUX2_X1 U16390 ( .A(n15264), .B(n15263), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16391 ( .A(n15265), .ZN(n15266) );
  MUX2_X1 U16392 ( .A(n15266), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XOR2_X1 U16393 ( .A(SI_31_), .B(keyinput_129), .Z(n15269) );
  XOR2_X1 U16394 ( .A(P3_WR_REG_SCAN_IN), .B(keyinput_128), .Z(n15268) );
  XNOR2_X1 U16395 ( .A(SI_30_), .B(keyinput_130), .ZN(n15267) );
  NAND3_X1 U16396 ( .A1(n15269), .A2(n15268), .A3(n15267), .ZN(n15272) );
  XNOR2_X1 U16397 ( .A(n15456), .B(keyinput_131), .ZN(n15271) );
  XNOR2_X1 U16398 ( .A(SI_28_), .B(keyinput_132), .ZN(n15270) );
  AOI21_X1 U16399 ( .B1(n15272), .B2(n15271), .A(n15270), .ZN(n15279) );
  XNOR2_X1 U16400 ( .A(SI_27_), .B(keyinput_133), .ZN(n15278) );
  XOR2_X1 U16401 ( .A(SI_24_), .B(keyinput_136), .Z(n15276) );
  XNOR2_X1 U16402 ( .A(SI_23_), .B(keyinput_137), .ZN(n15275) );
  XNOR2_X1 U16403 ( .A(SI_26_), .B(keyinput_134), .ZN(n15274) );
  XNOR2_X1 U16404 ( .A(SI_25_), .B(keyinput_135), .ZN(n15273) );
  NOR4_X1 U16405 ( .A1(n15276), .A2(n15275), .A3(n15274), .A4(n15273), .ZN(
        n15277) );
  OAI21_X1 U16406 ( .B1(n15279), .B2(n15278), .A(n15277), .ZN(n15284) );
  XOR2_X1 U16407 ( .A(SI_21_), .B(keyinput_139), .Z(n15283) );
  XNOR2_X1 U16408 ( .A(n15280), .B(keyinput_140), .ZN(n15282) );
  XOR2_X1 U16409 ( .A(SI_22_), .B(keyinput_138), .Z(n15281) );
  NAND4_X1 U16410 ( .A1(n15284), .A2(n15283), .A3(n15282), .A4(n15281), .ZN(
        n15287) );
  XOR2_X1 U16411 ( .A(SI_18_), .B(keyinput_142), .Z(n15286) );
  XNOR2_X1 U16412 ( .A(SI_19_), .B(keyinput_141), .ZN(n15285) );
  NAND3_X1 U16413 ( .A1(n15287), .A2(n15286), .A3(n15285), .ZN(n15291) );
  XNOR2_X1 U16414 ( .A(n15477), .B(keyinput_143), .ZN(n15290) );
  XOR2_X1 U16415 ( .A(SI_16_), .B(keyinput_144), .Z(n15289) );
  XNOR2_X1 U16416 ( .A(SI_15_), .B(keyinput_145), .ZN(n15288) );
  NAND4_X1 U16417 ( .A1(n15291), .A2(n15290), .A3(n15289), .A4(n15288), .ZN(
        n15294) );
  XNOR2_X1 U16418 ( .A(SI_14_), .B(keyinput_146), .ZN(n15293) );
  XNOR2_X1 U16419 ( .A(SI_13_), .B(keyinput_147), .ZN(n15292) );
  AOI21_X1 U16420 ( .B1(n15294), .B2(n15293), .A(n15292), .ZN(n15300) );
  XNOR2_X1 U16421 ( .A(n15485), .B(keyinput_148), .ZN(n15299) );
  XOR2_X1 U16422 ( .A(SI_9_), .B(keyinput_151), .Z(n15297) );
  XNOR2_X1 U16423 ( .A(SI_10_), .B(keyinput_150), .ZN(n15296) );
  XNOR2_X1 U16424 ( .A(SI_11_), .B(keyinput_149), .ZN(n15295) );
  NOR3_X1 U16425 ( .A1(n15297), .A2(n15296), .A3(n15295), .ZN(n15298) );
  OAI21_X1 U16426 ( .B1(n15300), .B2(n15299), .A(n15298), .ZN(n15303) );
  XNOR2_X1 U16427 ( .A(SI_8_), .B(keyinput_152), .ZN(n15302) );
  XNOR2_X1 U16428 ( .A(SI_7_), .B(keyinput_153), .ZN(n15301) );
  AOI21_X1 U16429 ( .B1(n15303), .B2(n15302), .A(n15301), .ZN(n15309) );
  XOR2_X1 U16430 ( .A(SI_6_), .B(keyinput_154), .Z(n15308) );
  XOR2_X1 U16431 ( .A(SI_3_), .B(keyinput_157), .Z(n15306) );
  XNOR2_X1 U16432 ( .A(SI_5_), .B(keyinput_155), .ZN(n15305) );
  XNOR2_X1 U16433 ( .A(SI_4_), .B(keyinput_156), .ZN(n15304) );
  NOR3_X1 U16434 ( .A1(n15306), .A2(n15305), .A3(n15304), .ZN(n15307) );
  OAI21_X1 U16435 ( .B1(n15309), .B2(n15308), .A(n15307), .ZN(n15312) );
  XNOR2_X1 U16436 ( .A(n15502), .B(keyinput_158), .ZN(n15311) );
  XOR2_X1 U16437 ( .A(SI_1_), .B(keyinput_159), .Z(n15310) );
  AOI21_X1 U16438 ( .B1(n15312), .B2(n15311), .A(n15310), .ZN(n15318) );
  XNOR2_X1 U16439 ( .A(SI_0_), .B(keyinput_160), .ZN(n15317) );
  XNOR2_X1 U16440 ( .A(P3_U3151), .B(keyinput_162), .ZN(n15315) );
  INV_X1 U16441 ( .A(P3_RD_REG_SCAN_IN), .ZN(n16001) );
  XNOR2_X1 U16442 ( .A(n16001), .B(keyinput_161), .ZN(n15314) );
  XNOR2_X1 U16443 ( .A(P3_REG3_REG_7__SCAN_IN), .B(keyinput_163), .ZN(n15313)
         );
  NOR3_X1 U16444 ( .A1(n15315), .A2(n15314), .A3(n15313), .ZN(n15316) );
  OAI21_X1 U16445 ( .B1(n15318), .B2(n15317), .A(n15316), .ZN(n15325) );
  XOR2_X1 U16446 ( .A(P3_REG3_REG_10__SCAN_IN), .B(keyinput_167), .Z(n15322)
         );
  XOR2_X1 U16447 ( .A(P3_REG3_REG_23__SCAN_IN), .B(keyinput_166), .Z(n15321)
         );
  XNOR2_X1 U16448 ( .A(P3_REG3_REG_27__SCAN_IN), .B(keyinput_164), .ZN(n15320)
         );
  XNOR2_X1 U16449 ( .A(P3_REG3_REG_14__SCAN_IN), .B(keyinput_165), .ZN(n15319)
         );
  NOR4_X1 U16450 ( .A1(n15322), .A2(n15321), .A3(n15320), .A4(n15319), .ZN(
        n15324) );
  XNOR2_X1 U16451 ( .A(P3_REG3_REG_3__SCAN_IN), .B(keyinput_168), .ZN(n15323)
         );
  AOI21_X1 U16452 ( .B1(n15325), .B2(n15324), .A(n15323), .ZN(n15331) );
  XOR2_X1 U16453 ( .A(P3_REG3_REG_19__SCAN_IN), .B(keyinput_169), .Z(n15330)
         );
  XNOR2_X1 U16454 ( .A(P3_REG3_REG_8__SCAN_IN), .B(keyinput_171), .ZN(n15328)
         );
  XNOR2_X1 U16455 ( .A(P3_REG3_REG_1__SCAN_IN), .B(keyinput_172), .ZN(n15327)
         );
  XNOR2_X1 U16456 ( .A(P3_REG3_REG_28__SCAN_IN), .B(keyinput_170), .ZN(n15326)
         );
  NOR3_X1 U16457 ( .A1(n15328), .A2(n15327), .A3(n15326), .ZN(n15329) );
  OAI21_X1 U16458 ( .B1(n15331), .B2(n15330), .A(n15329), .ZN(n15334) );
  XNOR2_X1 U16459 ( .A(P3_REG3_REG_21__SCAN_IN), .B(keyinput_173), .ZN(n15333)
         );
  XOR2_X1 U16460 ( .A(P3_REG3_REG_12__SCAN_IN), .B(keyinput_174), .Z(n15332)
         );
  AOI21_X1 U16461 ( .B1(n15334), .B2(n15333), .A(n15332), .ZN(n15337) );
  XNOR2_X1 U16462 ( .A(P3_REG3_REG_16__SCAN_IN), .B(keyinput_176), .ZN(n15336)
         );
  XNOR2_X1 U16463 ( .A(P3_REG3_REG_25__SCAN_IN), .B(keyinput_175), .ZN(n15335)
         );
  NOR3_X1 U16464 ( .A1(n15337), .A2(n15336), .A3(n15335), .ZN(n15345) );
  XOR2_X1 U16465 ( .A(P3_REG3_REG_24__SCAN_IN), .B(keyinput_179), .Z(n15342)
         );
  XNOR2_X1 U16466 ( .A(n15338), .B(keyinput_177), .ZN(n15341) );
  XNOR2_X1 U16467 ( .A(P3_REG3_REG_4__SCAN_IN), .B(keyinput_180), .ZN(n15340)
         );
  XNOR2_X1 U16468 ( .A(P3_REG3_REG_17__SCAN_IN), .B(keyinput_178), .ZN(n15339)
         );
  NAND4_X1 U16469 ( .A1(n15342), .A2(n15341), .A3(n15340), .A4(n15339), .ZN(
        n15344) );
  XNOR2_X1 U16470 ( .A(P3_REG3_REG_9__SCAN_IN), .B(keyinput_181), .ZN(n15343)
         );
  OAI21_X1 U16471 ( .B1(n15345), .B2(n15344), .A(n15343), .ZN(n15355) );
  XOR2_X1 U16472 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_182), .Z(n15354) );
  INV_X1 U16473 ( .A(keyinput_185), .ZN(n15352) );
  XNOR2_X1 U16474 ( .A(n15346), .B(keyinput_183), .ZN(n15351) );
  INV_X1 U16475 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n15347) );
  OAI22_X1 U16476 ( .A1(n15347), .A2(keyinput_185), .B1(n15349), .B2(
        keyinput_184), .ZN(n15348) );
  AOI21_X1 U16477 ( .B1(n15349), .B2(keyinput_184), .A(n15348), .ZN(n15350) );
  OAI211_X1 U16478 ( .C1(P3_REG3_REG_22__SCAN_IN), .C2(n15352), .A(n15351), 
        .B(n15350), .ZN(n15353) );
  AOI21_X1 U16479 ( .B1(n15355), .B2(n15354), .A(n15353), .ZN(n15358) );
  XOR2_X1 U16480 ( .A(P3_REG3_REG_11__SCAN_IN), .B(keyinput_186), .Z(n15357)
         );
  XOR2_X1 U16481 ( .A(P3_REG3_REG_2__SCAN_IN), .B(keyinput_187), .Z(n15356) );
  NOR3_X1 U16482 ( .A1(n15358), .A2(n15357), .A3(n15356), .ZN(n15361) );
  XNOR2_X1 U16483 ( .A(n15549), .B(keyinput_188), .ZN(n15360) );
  XOR2_X1 U16484 ( .A(P3_REG3_REG_6__SCAN_IN), .B(keyinput_189), .Z(n15359) );
  OAI21_X1 U16485 ( .B1(n15361), .B2(n15360), .A(n15359), .ZN(n15364) );
  XOR2_X1 U16486 ( .A(P3_REG3_REG_26__SCAN_IN), .B(keyinput_190), .Z(n15363)
         );
  XNOR2_X1 U16487 ( .A(P3_REG3_REG_15__SCAN_IN), .B(keyinput_191), .ZN(n15362)
         );
  NAND3_X1 U16488 ( .A1(n15364), .A2(n15363), .A3(n15362), .ZN(n15367) );
  XOR2_X1 U16489 ( .A(P3_B_REG_SCAN_IN), .B(keyinput_192), .Z(n15366) );
  XOR2_X1 U16490 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(keyinput_193), .Z(n15365)
         );
  AOI21_X1 U16491 ( .B1(n15367), .B2(n15366), .A(n15365), .ZN(n15370) );
  XNOR2_X1 U16492 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(keyinput_194), .ZN(n15369) );
  XOR2_X1 U16493 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(keyinput_195), .Z(n15368)
         );
  OAI21_X1 U16494 ( .B1(n15370), .B2(n15369), .A(n15368), .ZN(n15373) );
  XOR2_X1 U16495 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(keyinput_196), .Z(n15372)
         );
  XNOR2_X1 U16496 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(keyinput_197), .ZN(n15371) );
  NAND3_X1 U16497 ( .A1(n15373), .A2(n15372), .A3(n15371), .ZN(n15376) );
  XNOR2_X1 U16498 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(keyinput_199), .ZN(n15375) );
  XNOR2_X1 U16499 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(keyinput_198), .ZN(n15374) );
  NAND3_X1 U16500 ( .A1(n15376), .A2(n15375), .A3(n15374), .ZN(n15379) );
  XOR2_X1 U16501 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(keyinput_200), .Z(n15378)
         );
  XNOR2_X1 U16502 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(keyinput_201), .ZN(n15377) );
  AOI21_X1 U16503 ( .B1(n15379), .B2(n15378), .A(n15377), .ZN(n15383) );
  XOR2_X1 U16504 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(keyinput_202), .Z(n15382)
         );
  XOR2_X1 U16505 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(keyinput_203), .Z(n15381)
         );
  XNOR2_X1 U16506 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(keyinput_204), .ZN(n15380) );
  NOR4_X1 U16507 ( .A1(n15383), .A2(n15382), .A3(n15381), .A4(n15380), .ZN(
        n15397) );
  XOR2_X1 U16508 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(keyinput_205), .Z(n15396)
         );
  AOI22_X1 U16509 ( .A1(P3_DATAO_REG_13__SCAN_IN), .A2(keyinput_211), .B1(
        P3_DATAO_REG_12__SCAN_IN), .B2(keyinput_212), .ZN(n15384) );
  OAI221_X1 U16510 ( .B1(P3_DATAO_REG_13__SCAN_IN), .B2(keyinput_211), .C1(
        P3_DATAO_REG_12__SCAN_IN), .C2(keyinput_212), .A(n15384), .ZN(n15387)
         );
  XNOR2_X1 U16511 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(keyinput_210), .ZN(n15386) );
  XNOR2_X1 U16512 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(keyinput_206), .ZN(n15385) );
  NOR3_X1 U16513 ( .A1(n15387), .A2(n15386), .A3(n15385), .ZN(n15395) );
  AOI22_X1 U16514 ( .A1(P3_DATAO_REG_16__SCAN_IN), .A2(keyinput_208), .B1(
        n15389), .B2(keyinput_209), .ZN(n15388) );
  OAI221_X1 U16515 ( .B1(P3_DATAO_REG_16__SCAN_IN), .B2(keyinput_208), .C1(
        n15389), .C2(keyinput_209), .A(n15388), .ZN(n15393) );
  XOR2_X1 U16516 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(keyinput_214), .Z(n15392)
         );
  XOR2_X1 U16517 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(keyinput_213), .Z(n15391)
         );
  XNOR2_X1 U16518 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(keyinput_207), .ZN(n15390) );
  NOR4_X1 U16519 ( .A1(n15393), .A2(n15392), .A3(n15391), .A4(n15390), .ZN(
        n15394) );
  OAI211_X1 U16520 ( .C1(n15397), .C2(n15396), .A(n15395), .B(n15394), .ZN(
        n15404) );
  XOR2_X1 U16521 ( .A(keyinput_217), .B(P3_DATAO_REG_7__SCAN_IN), .Z(n15400)
         );
  XOR2_X1 U16522 ( .A(keyinput_218), .B(P3_DATAO_REG_6__SCAN_IN), .Z(n15399)
         );
  XOR2_X1 U16523 ( .A(keyinput_219), .B(P3_DATAO_REG_5__SCAN_IN), .Z(n15398)
         );
  NOR3_X1 U16524 ( .A1(n15400), .A2(n15399), .A3(n15398), .ZN(n15403) );
  XNOR2_X1 U16525 ( .A(keyinput_216), .B(P3_DATAO_REG_8__SCAN_IN), .ZN(n15402)
         );
  XNOR2_X1 U16526 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(keyinput_215), .ZN(n15401)
         );
  NAND4_X1 U16527 ( .A1(n15404), .A2(n15403), .A3(n15402), .A4(n15401), .ZN(
        n15408) );
  XOR2_X1 U16528 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(keyinput_220), .Z(n15407)
         );
  XOR2_X1 U16529 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(keyinput_221), .Z(n15406)
         );
  XNOR2_X1 U16530 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(keyinput_222), .ZN(n15405)
         );
  AOI211_X1 U16531 ( .C1(n15408), .C2(n15407), .A(n15406), .B(n15405), .ZN(
        n15415) );
  XOR2_X1 U16532 ( .A(P3_ADDR_REG_0__SCAN_IN), .B(keyinput_225), .Z(n15411) );
  XOR2_X1 U16533 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(keyinput_223), .Z(n15410)
         );
  XNOR2_X1 U16534 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(keyinput_224), .ZN(n15409)
         );
  NAND3_X1 U16535 ( .A1(n15411), .A2(n15410), .A3(n15409), .ZN(n15414) );
  XOR2_X1 U16536 ( .A(P3_ADDR_REG_2__SCAN_IN), .B(keyinput_227), .Z(n15413) );
  XOR2_X1 U16537 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(keyinput_226), .Z(n15412) );
  OAI211_X1 U16538 ( .C1(n15415), .C2(n15414), .A(n15413), .B(n15412), .ZN(
        n15418) );
  XNOR2_X1 U16539 ( .A(P3_ADDR_REG_3__SCAN_IN), .B(keyinput_228), .ZN(n15417)
         );
  XOR2_X1 U16540 ( .A(P3_ADDR_REG_4__SCAN_IN), .B(keyinput_229), .Z(n15416) );
  AOI21_X1 U16541 ( .B1(n15418), .B2(n15417), .A(n15416), .ZN(n15421) );
  XOR2_X1 U16542 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(keyinput_231), .Z(n15420) );
  XNOR2_X1 U16543 ( .A(P3_ADDR_REG_5__SCAN_IN), .B(keyinput_230), .ZN(n15419)
         );
  NOR3_X1 U16544 ( .A1(n15421), .A2(n15420), .A3(n15419), .ZN(n15424) );
  XOR2_X1 U16545 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(keyinput_233), .Z(n15423) );
  XNOR2_X1 U16546 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(keyinput_232), .ZN(n15422)
         );
  NOR3_X1 U16547 ( .A1(n15424), .A2(n15423), .A3(n15422), .ZN(n15428) );
  XOR2_X1 U16548 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(keyinput_234), .Z(n15427) );
  XNOR2_X1 U16549 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_235), .ZN(n15426) );
  XNOR2_X1 U16550 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_236), .ZN(n15425) );
  OAI211_X1 U16551 ( .C1(n15428), .C2(n15427), .A(n15426), .B(n15425), .ZN(
        n15432) );
  XNOR2_X1 U16552 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_237), .ZN(n15431) );
  XNOR2_X1 U16553 ( .A(n9344), .B(keyinput_238), .ZN(n15430) );
  XNOR2_X1 U16554 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_239), .ZN(n15429) );
  AOI211_X1 U16555 ( .C1(n15432), .C2(n15431), .A(n15430), .B(n15429), .ZN(
        n15435) );
  XNOR2_X1 U16556 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_240), .ZN(n15434) );
  XNOR2_X1 U16557 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_241), .ZN(n15433) );
  NOR3_X1 U16558 ( .A1(n15435), .A2(n15434), .A3(n15433), .ZN(n15438) );
  XNOR2_X1 U16559 ( .A(n15635), .B(keyinput_243), .ZN(n15437) );
  XNOR2_X1 U16560 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_242), .ZN(n15436) );
  NOR3_X1 U16561 ( .A1(n15438), .A2(n15437), .A3(n15436), .ZN(n15445) );
  XOR2_X1 U16562 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_246), .Z(n15442) );
  XNOR2_X1 U16563 ( .A(n15639), .B(keyinput_247), .ZN(n15441) );
  XNOR2_X1 U16564 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_245), .ZN(n15440)
         );
  XNOR2_X1 U16565 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_244), .ZN(n15439) );
  NAND4_X1 U16566 ( .A1(n15442), .A2(n15441), .A3(n15440), .A4(n15439), .ZN(
        n15444) );
  XNOR2_X1 U16567 ( .A(n15646), .B(keyinput_248), .ZN(n15443) );
  OAI21_X1 U16568 ( .B1(n15445), .B2(n15444), .A(n15443), .ZN(n15452) );
  OAI22_X1 U16569 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput_252), .B1(
        P1_IR_REG_16__SCAN_IN), .B2(keyinput_251), .ZN(n15446) );
  AOI221_X1 U16570 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput_252), .C1(
        keyinput_251), .C2(P1_IR_REG_16__SCAN_IN), .A(n15446), .ZN(n15451) );
  XNOR2_X1 U16571 ( .A(n15447), .B(keyinput_250), .ZN(n15450) );
  OAI22_X1 U16572 ( .A1(n15650), .A2(keyinput_253), .B1(P1_IR_REG_14__SCAN_IN), 
        .B2(keyinput_249), .ZN(n15448) );
  AOI221_X1 U16573 ( .B1(n15650), .B2(keyinput_253), .C1(keyinput_249), .C2(
        P1_IR_REG_14__SCAN_IN), .A(n15448), .ZN(n15449) );
  NAND4_X1 U16574 ( .A1(n15452), .A2(n15451), .A3(n15450), .A4(n15449), .ZN(
        n15665) );
  XNOR2_X1 U16575 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_254), .ZN(n15664)
         );
  XNOR2_X1 U16576 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_255), .ZN(n15663)
         );
  XOR2_X1 U16577 ( .A(SI_30_), .B(keyinput_2), .Z(n15455) );
  XNOR2_X1 U16578 ( .A(SI_31_), .B(keyinput_1), .ZN(n15454) );
  XNOR2_X1 U16579 ( .A(P3_WR_REG_SCAN_IN), .B(keyinput_0), .ZN(n15453) );
  NOR3_X1 U16580 ( .A1(n15455), .A2(n15454), .A3(n15453), .ZN(n15459) );
  XNOR2_X1 U16581 ( .A(n15456), .B(keyinput_3), .ZN(n15458) );
  XNOR2_X1 U16582 ( .A(SI_28_), .B(keyinput_4), .ZN(n15457) );
  OAI21_X1 U16583 ( .B1(n15459), .B2(n15458), .A(n15457), .ZN(n15468) );
  XNOR2_X1 U16584 ( .A(n15460), .B(keyinput_5), .ZN(n15467) );
  XOR2_X1 U16585 ( .A(SI_23_), .B(keyinput_9), .Z(n15465) );
  XOR2_X1 U16586 ( .A(SI_26_), .B(keyinput_6), .Z(n15464) );
  XOR2_X1 U16587 ( .A(SI_24_), .B(keyinput_8), .Z(n15463) );
  XNOR2_X1 U16588 ( .A(n15461), .B(keyinput_7), .ZN(n15462) );
  NAND4_X1 U16589 ( .A1(n15465), .A2(n15464), .A3(n15463), .A4(n15462), .ZN(
        n15466) );
  AOI21_X1 U16590 ( .B1(n15468), .B2(n15467), .A(n15466), .ZN(n15472) );
  XOR2_X1 U16591 ( .A(SI_21_), .B(keyinput_11), .Z(n15471) );
  XOR2_X1 U16592 ( .A(SI_22_), .B(keyinput_10), .Z(n15470) );
  XNOR2_X1 U16593 ( .A(SI_20_), .B(keyinput_12), .ZN(n15469) );
  NOR4_X1 U16594 ( .A1(n15472), .A2(n15471), .A3(n15470), .A4(n15469), .ZN(
        n15476) );
  XNOR2_X1 U16595 ( .A(n15473), .B(keyinput_13), .ZN(n15475) );
  XNOR2_X1 U16596 ( .A(SI_18_), .B(keyinput_14), .ZN(n15474) );
  NOR3_X1 U16597 ( .A1(n15476), .A2(n15475), .A3(n15474), .ZN(n15481) );
  XOR2_X1 U16598 ( .A(SI_16_), .B(keyinput_16), .Z(n15480) );
  XNOR2_X1 U16599 ( .A(n15477), .B(keyinput_15), .ZN(n15479) );
  XNOR2_X1 U16600 ( .A(SI_15_), .B(keyinput_17), .ZN(n15478) );
  NOR4_X1 U16601 ( .A1(n15481), .A2(n15480), .A3(n15479), .A4(n15478), .ZN(
        n15484) );
  XNOR2_X1 U16602 ( .A(SI_14_), .B(keyinput_18), .ZN(n15483) );
  XNOR2_X1 U16603 ( .A(SI_13_), .B(keyinput_19), .ZN(n15482) );
  OAI21_X1 U16604 ( .B1(n15484), .B2(n15483), .A(n15482), .ZN(n15491) );
  XNOR2_X1 U16605 ( .A(n15485), .B(keyinput_20), .ZN(n15490) );
  XOR2_X1 U16606 ( .A(SI_9_), .B(keyinput_23), .Z(n15488) );
  XOR2_X1 U16607 ( .A(SI_10_), .B(keyinput_22), .Z(n15487) );
  XNOR2_X1 U16608 ( .A(SI_11_), .B(keyinput_21), .ZN(n15486) );
  NAND3_X1 U16609 ( .A1(n15488), .A2(n15487), .A3(n15486), .ZN(n15489) );
  AOI21_X1 U16610 ( .B1(n15491), .B2(n15490), .A(n15489), .ZN(n15494) );
  XNOR2_X1 U16611 ( .A(SI_8_), .B(keyinput_24), .ZN(n15493) );
  XNOR2_X1 U16612 ( .A(SI_7_), .B(keyinput_25), .ZN(n15492) );
  OAI21_X1 U16613 ( .B1(n15494), .B2(n15493), .A(n15492), .ZN(n15501) );
  XOR2_X1 U16614 ( .A(SI_6_), .B(keyinput_26), .Z(n15500) );
  XOR2_X1 U16615 ( .A(SI_5_), .B(keyinput_27), .Z(n15498) );
  XNOR2_X1 U16616 ( .A(n15495), .B(keyinput_28), .ZN(n15497) );
  XNOR2_X1 U16617 ( .A(SI_3_), .B(keyinput_29), .ZN(n15496) );
  NAND3_X1 U16618 ( .A1(n15498), .A2(n15497), .A3(n15496), .ZN(n15499) );
  AOI21_X1 U16619 ( .B1(n15501), .B2(n15500), .A(n15499), .ZN(n15505) );
  XNOR2_X1 U16620 ( .A(n15502), .B(keyinput_30), .ZN(n15504) );
  XOR2_X1 U16621 ( .A(SI_1_), .B(keyinput_31), .Z(n15503) );
  OAI21_X1 U16622 ( .B1(n15505), .B2(n15504), .A(n15503), .ZN(n15511) );
  XOR2_X1 U16623 ( .A(SI_0_), .B(keyinput_32), .Z(n15510) );
  XNOR2_X1 U16624 ( .A(P3_U3151), .B(keyinput_34), .ZN(n15508) );
  XNOR2_X1 U16625 ( .A(n16001), .B(keyinput_33), .ZN(n15507) );
  XNOR2_X1 U16626 ( .A(P3_REG3_REG_7__SCAN_IN), .B(keyinput_35), .ZN(n15506)
         );
  NAND3_X1 U16627 ( .A1(n15508), .A2(n15507), .A3(n15506), .ZN(n15509) );
  AOI21_X1 U16628 ( .B1(n15511), .B2(n15510), .A(n15509), .ZN(n15518) );
  XOR2_X1 U16629 ( .A(P3_REG3_REG_23__SCAN_IN), .B(keyinput_38), .Z(n15515) );
  XOR2_X1 U16630 ( .A(P3_REG3_REG_10__SCAN_IN), .B(keyinput_39), .Z(n15514) );
  XNOR2_X1 U16631 ( .A(P3_REG3_REG_14__SCAN_IN), .B(keyinput_37), .ZN(n15513)
         );
  XNOR2_X1 U16632 ( .A(P3_REG3_REG_27__SCAN_IN), .B(keyinput_36), .ZN(n15512)
         );
  NAND4_X1 U16633 ( .A1(n15515), .A2(n15514), .A3(n15513), .A4(n15512), .ZN(
        n15517) );
  XNOR2_X1 U16634 ( .A(P3_REG3_REG_3__SCAN_IN), .B(keyinput_40), .ZN(n15516)
         );
  OAI21_X1 U16635 ( .B1(n15518), .B2(n15517), .A(n15516), .ZN(n15524) );
  XOR2_X1 U16636 ( .A(P3_REG3_REG_19__SCAN_IN), .B(keyinput_41), .Z(n15523) );
  XNOR2_X1 U16637 ( .A(P3_REG3_REG_28__SCAN_IN), .B(keyinput_42), .ZN(n15521)
         );
  XNOR2_X1 U16638 ( .A(P3_REG3_REG_1__SCAN_IN), .B(keyinput_44), .ZN(n15520)
         );
  XNOR2_X1 U16639 ( .A(P3_REG3_REG_8__SCAN_IN), .B(keyinput_43), .ZN(n15519)
         );
  NAND3_X1 U16640 ( .A1(n15521), .A2(n15520), .A3(n15519), .ZN(n15522) );
  AOI21_X1 U16641 ( .B1(n15524), .B2(n15523), .A(n15522), .ZN(n15527) );
  XNOR2_X1 U16642 ( .A(P3_REG3_REG_21__SCAN_IN), .B(keyinput_45), .ZN(n15526)
         );
  XOR2_X1 U16643 ( .A(P3_REG3_REG_12__SCAN_IN), .B(keyinput_46), .Z(n15525) );
  OAI21_X1 U16644 ( .B1(n15527), .B2(n15526), .A(n15525), .ZN(n15530) );
  XNOR2_X1 U16645 ( .A(P3_REG3_REG_25__SCAN_IN), .B(keyinput_47), .ZN(n15529)
         );
  XNOR2_X1 U16646 ( .A(P3_REG3_REG_16__SCAN_IN), .B(keyinput_48), .ZN(n15528)
         );
  NAND3_X1 U16647 ( .A1(n15530), .A2(n15529), .A3(n15528), .ZN(n15539) );
  XOR2_X1 U16648 ( .A(P3_REG3_REG_4__SCAN_IN), .B(keyinput_52), .Z(n15535) );
  XNOR2_X1 U16649 ( .A(n15531), .B(keyinput_50), .ZN(n15534) );
  XNOR2_X1 U16650 ( .A(P3_REG3_REG_5__SCAN_IN), .B(keyinput_49), .ZN(n15533)
         );
  XNOR2_X1 U16651 ( .A(P3_REG3_REG_24__SCAN_IN), .B(keyinput_51), .ZN(n15532)
         );
  NOR4_X1 U16652 ( .A1(n15535), .A2(n15534), .A3(n15533), .A4(n15532), .ZN(
        n15538) );
  XNOR2_X1 U16653 ( .A(n15536), .B(keyinput_53), .ZN(n15537) );
  AOI21_X1 U16654 ( .B1(n15539), .B2(n15538), .A(n15537), .ZN(n15545) );
  XOR2_X1 U16655 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_54), .Z(n15544) );
  XNOR2_X1 U16656 ( .A(P3_REG3_REG_13__SCAN_IN), .B(keyinput_56), .ZN(n15542)
         );
  XNOR2_X1 U16657 ( .A(P3_REG3_REG_20__SCAN_IN), .B(keyinput_55), .ZN(n15541)
         );
  XNOR2_X1 U16658 ( .A(P3_REG3_REG_22__SCAN_IN), .B(keyinput_57), .ZN(n15540)
         );
  NOR3_X1 U16659 ( .A1(n15542), .A2(n15541), .A3(n15540), .ZN(n15543) );
  OAI21_X1 U16660 ( .B1(n15545), .B2(n15544), .A(n15543), .ZN(n15548) );
  XNOR2_X1 U16661 ( .A(P3_REG3_REG_11__SCAN_IN), .B(keyinput_58), .ZN(n15547)
         );
  XNOR2_X1 U16662 ( .A(P3_REG3_REG_2__SCAN_IN), .B(keyinput_59), .ZN(n15546)
         );
  NAND3_X1 U16663 ( .A1(n15548), .A2(n15547), .A3(n15546), .ZN(n15552) );
  XNOR2_X1 U16664 ( .A(n15549), .B(keyinput_60), .ZN(n15551) );
  XNOR2_X1 U16665 ( .A(P3_REG3_REG_6__SCAN_IN), .B(keyinput_61), .ZN(n15550)
         );
  AOI21_X1 U16666 ( .B1(n15552), .B2(n15551), .A(n15550), .ZN(n15555) );
  XOR2_X1 U16667 ( .A(P3_REG3_REG_15__SCAN_IN), .B(keyinput_63), .Z(n15554) );
  XNOR2_X1 U16668 ( .A(P3_REG3_REG_26__SCAN_IN), .B(keyinput_62), .ZN(n15553)
         );
  NOR3_X1 U16669 ( .A1(n15555), .A2(n15554), .A3(n15553), .ZN(n15558) );
  XOR2_X1 U16670 ( .A(P3_B_REG_SCAN_IN), .B(keyinput_64), .Z(n15557) );
  XOR2_X1 U16671 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(keyinput_65), .Z(n15556)
         );
  OAI21_X1 U16672 ( .B1(n15558), .B2(n15557), .A(n15556), .ZN(n15561) );
  XNOR2_X1 U16673 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(keyinput_66), .ZN(n15560)
         );
  XOR2_X1 U16674 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(keyinput_67), .Z(n15559)
         );
  AOI21_X1 U16675 ( .B1(n15561), .B2(n15560), .A(n15559), .ZN(n15564) );
  XOR2_X1 U16676 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(keyinput_68), .Z(n15563)
         );
  XNOR2_X1 U16677 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(keyinput_69), .ZN(n15562)
         );
  NOR3_X1 U16678 ( .A1(n15564), .A2(n15563), .A3(n15562), .ZN(n15567) );
  XOR2_X1 U16679 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(keyinput_70), .Z(n15566)
         );
  XNOR2_X1 U16680 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(keyinput_71), .ZN(n15565)
         );
  NOR3_X1 U16681 ( .A1(n15567), .A2(n15566), .A3(n15565), .ZN(n15570) );
  XNOR2_X1 U16682 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(keyinput_72), .ZN(n15569)
         );
  XNOR2_X1 U16683 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(keyinput_73), .ZN(n15568)
         );
  OAI21_X1 U16684 ( .B1(n15570), .B2(n15569), .A(n15568), .ZN(n15574) );
  XOR2_X1 U16685 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .Z(n15573)
         );
  XNOR2_X1 U16686 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(keyinput_74), .ZN(n15572)
         );
  XNOR2_X1 U16687 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(keyinput_76), .ZN(n15571)
         );
  NAND4_X1 U16688 ( .A1(n15574), .A2(n15573), .A3(n15572), .A4(n15571), .ZN(
        n15576) );
  XOR2_X1 U16689 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .Z(n15575)
         );
  NAND2_X1 U16690 ( .A1(n15576), .A2(n15575), .ZN(n15593) );
  OAI22_X1 U16691 ( .A1(keyinput_81), .A2(P3_DATAO_REG_15__SCAN_IN), .B1(
        P3_DATAO_REG_17__SCAN_IN), .B2(keyinput_79), .ZN(n15578) );
  OAI22_X1 U16692 ( .A1(keyinput_83), .A2(P3_DATAO_REG_13__SCAN_IN), .B1(
        P3_DATAO_REG_10__SCAN_IN), .B2(keyinput_86), .ZN(n15577) );
  OR2_X1 U16693 ( .A1(n15578), .A2(n15577), .ZN(n15587) );
  INV_X1 U16694 ( .A(keyinput_85), .ZN(n15579) );
  NAND2_X1 U16695 ( .A1(n15579), .A2(P3_DATAO_REG_11__SCAN_IN), .ZN(n15585) );
  INV_X1 U16696 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n15580) );
  AOI22_X1 U16697 ( .A1(keyinput_81), .A2(P3_DATAO_REG_15__SCAN_IN), .B1(
        n15580), .B2(keyinput_85), .ZN(n15583) );
  AOI22_X1 U16698 ( .A1(P3_DATAO_REG_17__SCAN_IN), .A2(keyinput_79), .B1(
        P3_DATAO_REG_18__SCAN_IN), .B2(keyinput_78), .ZN(n15582) );
  AOI22_X1 U16699 ( .A1(P3_DATAO_REG_10__SCAN_IN), .A2(keyinput_86), .B1(
        P3_DATAO_REG_13__SCAN_IN), .B2(keyinput_83), .ZN(n15581) );
  AND3_X1 U16700 ( .A1(n15583), .A2(n15582), .A3(n15581), .ZN(n15584) );
  OAI211_X1 U16701 ( .C1(P3_DATAO_REG_18__SCAN_IN), .C2(keyinput_78), .A(
        n15585), .B(n15584), .ZN(n15586) );
  NOR2_X1 U16702 ( .A1(n15587), .A2(n15586), .ZN(n15592) );
  XNOR2_X1 U16703 ( .A(keyinput_84), .B(P3_DATAO_REG_12__SCAN_IN), .ZN(n15589)
         );
  XNOR2_X1 U16704 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(keyinput_82), .ZN(n15588)
         );
  AND2_X1 U16705 ( .A1(n15589), .A2(n15588), .ZN(n15591) );
  XNOR2_X1 U16706 ( .A(keyinput_80), .B(P3_DATAO_REG_16__SCAN_IN), .ZN(n15590)
         );
  NAND4_X1 U16707 ( .A1(n15593), .A2(n15592), .A3(n15591), .A4(n15590), .ZN(
        n15601) );
  INV_X1 U16708 ( .A(P3_DATAO_REG_8__SCAN_IN), .ZN(n15595) );
  OAI22_X1 U16709 ( .A1(n15595), .A2(keyinput_88), .B1(P3_DATAO_REG_7__SCAN_IN), .B2(keyinput_89), .ZN(n15594) );
  AOI221_X1 U16710 ( .B1(n15595), .B2(keyinput_88), .C1(keyinput_89), .C2(
        P3_DATAO_REG_7__SCAN_IN), .A(n15594), .ZN(n15600) );
  XOR2_X1 U16711 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(keyinput_87), .Z(n15599) );
  INV_X1 U16712 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n15597) );
  OAI22_X1 U16713 ( .A1(n15597), .A2(keyinput_91), .B1(P3_DATAO_REG_6__SCAN_IN), .B2(keyinput_90), .ZN(n15596) );
  AOI221_X1 U16714 ( .B1(n15597), .B2(keyinput_91), .C1(keyinput_90), .C2(
        P3_DATAO_REG_6__SCAN_IN), .A(n15596), .ZN(n15598) );
  NAND4_X1 U16715 ( .A1(n15601), .A2(n15600), .A3(n15599), .A4(n15598), .ZN(
        n15605) );
  XNOR2_X1 U16716 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(keyinput_92), .ZN(n15604)
         );
  XOR2_X1 U16717 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(keyinput_93), .Z(n15603) );
  XOR2_X1 U16718 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(keyinput_94), .Z(n15602) );
  AOI211_X1 U16719 ( .C1(n15605), .C2(n15604), .A(n15603), .B(n15602), .ZN(
        n15612) );
  XOR2_X1 U16720 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(keyinput_95), .Z(n15608) );
  XNOR2_X1 U16721 ( .A(P3_ADDR_REG_0__SCAN_IN), .B(keyinput_97), .ZN(n15607)
         );
  XNOR2_X1 U16722 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(keyinput_96), .ZN(n15606)
         );
  NAND3_X1 U16723 ( .A1(n15608), .A2(n15607), .A3(n15606), .ZN(n15611) );
  XOR2_X1 U16724 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(keyinput_98), .Z(n15610) );
  XOR2_X1 U16725 ( .A(P3_ADDR_REG_2__SCAN_IN), .B(keyinput_99), .Z(n15609) );
  OAI211_X1 U16726 ( .C1(n15612), .C2(n15611), .A(n15610), .B(n15609), .ZN(
        n15615) );
  XNOR2_X1 U16727 ( .A(P3_ADDR_REG_3__SCAN_IN), .B(keyinput_100), .ZN(n15614)
         );
  XOR2_X1 U16728 ( .A(P3_ADDR_REG_4__SCAN_IN), .B(keyinput_101), .Z(n15613) );
  AOI21_X1 U16729 ( .B1(n15615), .B2(n15614), .A(n15613), .ZN(n15618) );
  XOR2_X1 U16730 ( .A(P3_ADDR_REG_5__SCAN_IN), .B(keyinput_102), .Z(n15617) );
  XOR2_X1 U16731 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(keyinput_103), .Z(n15616) );
  NOR3_X1 U16732 ( .A1(n15618), .A2(n15617), .A3(n15616), .ZN(n15621) );
  XOR2_X1 U16733 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(keyinput_104), .Z(n15620) );
  XOR2_X1 U16734 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(keyinput_105), .Z(n15619) );
  NOR3_X1 U16735 ( .A1(n15621), .A2(n15620), .A3(n15619), .ZN(n15626) );
  XNOR2_X1 U16736 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(keyinput_106), .ZN(n15625)
         );
  XNOR2_X1 U16737 ( .A(n15622), .B(keyinput_108), .ZN(n15624) );
  XNOR2_X1 U16738 ( .A(n8323), .B(keyinput_107), .ZN(n15623) );
  OAI211_X1 U16739 ( .C1(n15626), .C2(n15625), .A(n15624), .B(n15623), .ZN(
        n15631) );
  XNOR2_X1 U16740 ( .A(n15627), .B(keyinput_109), .ZN(n15630) );
  XOR2_X1 U16741 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_111), .Z(n15629) );
  XNOR2_X1 U16742 ( .A(n9344), .B(keyinput_110), .ZN(n15628) );
  AOI211_X1 U16743 ( .C1(n15631), .C2(n15630), .A(n15629), .B(n15628), .ZN(
        n15634) );
  XOR2_X1 U16744 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_112), .Z(n15633) );
  XNOR2_X1 U16745 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_113), .ZN(n15632) );
  NOR3_X1 U16746 ( .A1(n15634), .A2(n15633), .A3(n15632), .ZN(n15638) );
  XNOR2_X1 U16747 ( .A(n15635), .B(keyinput_115), .ZN(n15637) );
  XNOR2_X1 U16748 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_114), .ZN(n15636) );
  NOR3_X1 U16749 ( .A1(n15638), .A2(n15637), .A3(n15636), .ZN(n15645) );
  XNOR2_X1 U16750 ( .A(n15639), .B(keyinput_119), .ZN(n15644) );
  XNOR2_X1 U16751 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_117), .ZN(n15641)
         );
  XNOR2_X1 U16752 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_116), .ZN(n15640) );
  NAND2_X1 U16753 ( .A1(n15641), .A2(n15640), .ZN(n15643) );
  XNOR2_X1 U16754 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_118), .ZN(n15642)
         );
  NOR4_X1 U16755 ( .A1(n15645), .A2(n15644), .A3(n15643), .A4(n15642), .ZN(
        n15657) );
  XNOR2_X1 U16756 ( .A(n15646), .B(keyinput_120), .ZN(n15656) );
  OAI22_X1 U16757 ( .A1(n15648), .A2(keyinput_121), .B1(P1_IR_REG_15__SCAN_IN), 
        .B2(keyinput_122), .ZN(n15647) );
  AOI221_X1 U16758 ( .B1(n15648), .B2(keyinput_121), .C1(keyinput_122), .C2(
        P1_IR_REG_15__SCAN_IN), .A(n15647), .ZN(n15655) );
  XNOR2_X1 U16759 ( .A(n15649), .B(keyinput_124), .ZN(n15653) );
  XNOR2_X1 U16760 ( .A(n15650), .B(keyinput_125), .ZN(n15652) );
  XNOR2_X1 U16761 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_123), .ZN(n15651)
         );
  NOR3_X1 U16762 ( .A1(n15653), .A2(n15652), .A3(n15651), .ZN(n15654) );
  OAI211_X1 U16763 ( .C1(n15657), .C2(n15656), .A(n15655), .B(n15654), .ZN(
        n15661) );
  XNOR2_X1 U16764 ( .A(n15658), .B(keyinput_126), .ZN(n15660) );
  XNOR2_X1 U16765 ( .A(keyinput_255), .B(keyinput_127), .ZN(n15659) );
  AOI21_X1 U16766 ( .B1(n15661), .B2(n15660), .A(n15659), .ZN(n15662) );
  AOI211_X1 U16767 ( .C1(n15665), .C2(n15664), .A(n15663), .B(n15662), .ZN(
        n15704) );
  INV_X1 U16768 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n15703) );
  INV_X1 U16769 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15857) );
  INV_X1 U16770 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n15928) );
  INV_X1 U16771 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n15666) );
  XNOR2_X1 U16772 ( .A(n15666), .B(n15694), .ZN(n15749) );
  INV_X1 U16773 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n15692) );
  XNOR2_X1 U16774 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n15692), .ZN(n15746) );
  INV_X1 U16775 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n15687) );
  XNOR2_X1 U16776 ( .A(n15667), .B(P1_ADDR_REG_8__SCAN_IN), .ZN(n15740) );
  NOR2_X1 U16777 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n15708), .ZN(n15679) );
  NOR2_X1 U16778 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n15678), .ZN(n15668) );
  AOI21_X1 U16779 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(n15678), .A(n15668), .ZN(
        n15711) );
  NAND2_X1 U16780 ( .A1(n15717), .A2(n15716), .ZN(n15669) );
  NAND2_X1 U16781 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n15670), .ZN(n15671) );
  XNOR2_X1 U16782 ( .A(P3_ADDR_REG_2__SCAN_IN), .B(n15670), .ZN(n15714) );
  NAND2_X1 U16783 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n15672), .ZN(n15676) );
  INV_X1 U16784 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n15673) );
  NAND2_X1 U16785 ( .A1(n15723), .A2(n15674), .ZN(n15675) );
  NAND2_X1 U16786 ( .A1(n15676), .A2(n15675), .ZN(n15712) );
  NAND2_X1 U16787 ( .A1(n15711), .A2(n15712), .ZN(n15677) );
  NAND2_X1 U16788 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n15708), .ZN(n15707) );
  NAND2_X1 U16789 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n15681), .ZN(n15684) );
  XOR2_X1 U16790 ( .A(n15682), .B(n15681), .Z(n15738) );
  NAND2_X1 U16791 ( .A1(n15687), .A2(n15688), .ZN(n15690) );
  XNOR2_X1 U16792 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(n15688), .ZN(n15705) );
  NAND2_X1 U16793 ( .A1(n15705), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n15689) );
  NAND2_X1 U16794 ( .A1(n15749), .A2(n15750), .ZN(n15693) );
  NAND2_X1 U16795 ( .A1(P3_ADDR_REG_12__SCAN_IN), .A2(n15695), .ZN(n15696) );
  INV_X1 U16796 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15943) );
  NAND2_X1 U16797 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n15943), .ZN(n15697) );
  XNOR2_X1 U16798 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(n15699), .ZN(n15760) );
  NOR2_X1 U16799 ( .A1(n15761), .A2(n15760), .ZN(n15698) );
  AOI21_X1 U16800 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n15699), .A(n15698), 
        .ZN(n15763) );
  INV_X1 U16801 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n15981) );
  XNOR2_X1 U16802 ( .A(n15981), .B(P1_ADDR_REG_15__SCAN_IN), .ZN(n15762) );
  NOR2_X1 U16803 ( .A1(n15763), .A2(n15762), .ZN(n15700) );
  AOI21_X1 U16804 ( .B1(P3_ADDR_REG_15__SCAN_IN), .B2(n15857), .A(n15700), 
        .ZN(n15768) );
  INV_X1 U16805 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n15701) );
  XNOR2_X1 U16806 ( .A(n15701), .B(P1_ADDR_REG_16__SCAN_IN), .ZN(n15767) );
  NOR2_X1 U16807 ( .A1(n15768), .A2(n15767), .ZN(n15702) );
  AOI21_X1 U16808 ( .B1(P3_ADDR_REG_16__SCAN_IN), .B2(n15703), .A(n15702), 
        .ZN(n15905) );
  XOR2_X1 U16809 ( .A(n15905), .B(P1_ADDR_REG_17__SCAN_IN), .Z(n15904) );
  XNOR2_X1 U16810 ( .A(n15904), .B(P3_ADDR_REG_17__SCAN_IN), .ZN(n15901) );
  XOR2_X1 U16811 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n15901), .Z(n15902) );
  INV_X1 U16812 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15756) );
  INV_X1 U16813 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n15752) );
  INV_X1 U16814 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n15748) );
  XNOR2_X1 U16815 ( .A(n15706), .B(n15705), .ZN(n15744) );
  OAI21_X1 U16816 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(n15708), .A(n15707), .ZN(
        n15709) );
  XOR2_X1 U16817 ( .A(n15710), .B(n15709), .Z(n15728) );
  XNOR2_X1 U16818 ( .A(n15712), .B(n15711), .ZN(n15713) );
  NAND2_X1 U16819 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n15713), .ZN(n15726) );
  XOR2_X1 U16820 ( .A(n15713), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n15866) );
  XOR2_X1 U16821 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n15714), .Z(n15721) );
  INV_X1 U16822 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15858) );
  XNOR2_X1 U16823 ( .A(n15716), .B(n15717), .ZN(n15919) );
  OR2_X1 U16824 ( .A1(n7441), .A2(n15919), .ZN(n15719) );
  INV_X1 U16825 ( .A(n15918), .ZN(n15718) );
  AOI21_X1 U16826 ( .B1(n15719), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n15718), .ZN(
        n15720) );
  AND2_X1 U16827 ( .A1(n15721), .A2(n15720), .ZN(n15861) );
  NOR2_X1 U16828 ( .A1(n15721), .A2(n15720), .ZN(n15860) );
  NOR2_X1 U16829 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(n15860), .ZN(n15722) );
  NOR2_X1 U16830 ( .A1(n15861), .A2(n15722), .ZN(n15725) );
  NAND2_X1 U16831 ( .A1(n15728), .A2(n15727), .ZN(n15729) );
  XOR2_X1 U16832 ( .A(n15730), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n15732) );
  XOR2_X1 U16833 ( .A(n15732), .B(n15731), .Z(n15734) );
  NAND2_X1 U16834 ( .A1(n15733), .A2(n15734), .ZN(n15735) );
  XOR2_X1 U16835 ( .A(n15739), .B(n15738), .Z(n15868) );
  XOR2_X1 U16836 ( .A(n15741), .B(n15740), .Z(n15742) );
  NOR2_X1 U16837 ( .A1(n15743), .A2(n15742), .ZN(n15870) );
  XNOR2_X1 U16838 ( .A(n15746), .B(n15745), .ZN(n15877) );
  NAND2_X1 U16839 ( .A1(n15878), .A2(n15877), .ZN(n15747) );
  XOR2_X1 U16840 ( .A(n15750), .B(n15749), .Z(n15882) );
  NAND2_X1 U16841 ( .A1(n15881), .A2(n15882), .ZN(n15751) );
  NOR2_X1 U16842 ( .A1(n15881), .A2(n15882), .ZN(n15880) );
  XNOR2_X1 U16843 ( .A(n15928), .B(P1_ADDR_REG_12__SCAN_IN), .ZN(n15753) );
  XNOR2_X1 U16844 ( .A(n15754), .B(n15753), .ZN(n15885) );
  NAND2_X1 U16845 ( .A1(n15886), .A2(n15885), .ZN(n15755) );
  NOR2_X1 U16846 ( .A1(n15886), .A2(n15885), .ZN(n15884) );
  XOR2_X1 U16847 ( .A(n15757), .B(n15943), .Z(n15759) );
  XOR2_X1 U16848 ( .A(n15759), .B(n15758), .Z(n15889) );
  XNOR2_X1 U16849 ( .A(n15761), .B(n15760), .ZN(n15893) );
  NOR2_X1 U16850 ( .A1(n15894), .A2(n15893), .ZN(n15892) );
  XOR2_X1 U16851 ( .A(n15763), .B(n15762), .Z(n15765) );
  AND2_X1 U16852 ( .A1(n15764), .A2(n15765), .ZN(n15897) );
  XNOR2_X1 U16853 ( .A(n15768), .B(n15767), .ZN(n15769) );
  OR2_X1 U16854 ( .A1(n15770), .A2(n15769), .ZN(n15774) );
  XNOR2_X1 U16855 ( .A(n15770), .B(n15769), .ZN(n15900) );
  INV_X1 U16856 ( .A(n15900), .ZN(n15771) );
  AND2_X1 U16857 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15775), .ZN(P1_U3323) );
  AND2_X1 U16858 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15775), .ZN(P1_U3322) );
  AND2_X1 U16859 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15775), .ZN(P1_U3321) );
  AND2_X1 U16860 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15775), .ZN(P1_U3320) );
  AND2_X1 U16861 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15775), .ZN(P1_U3319) );
  AND2_X1 U16862 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15775), .ZN(P1_U3318) );
  AND2_X1 U16863 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15775), .ZN(P1_U3317) );
  AND2_X1 U16864 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15775), .ZN(P1_U3316) );
  AND2_X1 U16865 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15775), .ZN(P1_U3315) );
  AND2_X1 U16866 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15775), .ZN(P1_U3314) );
  AND2_X1 U16867 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15775), .ZN(P1_U3313) );
  AND2_X1 U16868 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15775), .ZN(P1_U3312) );
  AND2_X1 U16869 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15775), .ZN(P1_U3311) );
  AND2_X1 U16870 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15775), .ZN(P1_U3310) );
  AND2_X1 U16871 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15775), .ZN(P1_U3309) );
  AND2_X1 U16872 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15775), .ZN(P1_U3308) );
  AND2_X1 U16873 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15775), .ZN(P1_U3307) );
  AND2_X1 U16874 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15775), .ZN(P1_U3306) );
  AND2_X1 U16875 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15775), .ZN(P1_U3305) );
  AND2_X1 U16876 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15775), .ZN(P1_U3304) );
  AND2_X1 U16877 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15775), .ZN(P1_U3303) );
  AND2_X1 U16878 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15775), .ZN(P1_U3302) );
  AND2_X1 U16879 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15775), .ZN(P1_U3301) );
  AND2_X1 U16880 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15775), .ZN(P1_U3300) );
  AND2_X1 U16881 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15775), .ZN(P1_U3299) );
  AND2_X1 U16882 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15775), .ZN(P1_U3298) );
  AND2_X1 U16883 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15775), .ZN(P1_U3297) );
  AND2_X1 U16884 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15775), .ZN(P1_U3296) );
  AND2_X1 U16885 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15775), .ZN(P1_U3295) );
  AND2_X1 U16886 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15775), .ZN(P1_U3294) );
  INV_X1 U16887 ( .A(n15776), .ZN(n15777) );
  AOI21_X1 U16888 ( .B1(n15778), .B2(n15781), .A(n15777), .ZN(P2_U3417) );
  AND2_X1 U16889 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15780), .ZN(P2_U3295) );
  AND2_X1 U16890 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15780), .ZN(P2_U3294) );
  AND2_X1 U16891 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15780), .ZN(P2_U3293) );
  AND2_X1 U16892 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15780), .ZN(P2_U3292) );
  AND2_X1 U16893 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15780), .ZN(P2_U3291) );
  AND2_X1 U16894 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15780), .ZN(P2_U3290) );
  AND2_X1 U16895 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15780), .ZN(P2_U3289) );
  AND2_X1 U16896 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15780), .ZN(P2_U3288) );
  AND2_X1 U16897 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15780), .ZN(P2_U3287) );
  AND2_X1 U16898 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15780), .ZN(P2_U3286) );
  AND2_X1 U16899 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15780), .ZN(P2_U3285) );
  AND2_X1 U16900 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15780), .ZN(P2_U3284) );
  AND2_X1 U16901 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15780), .ZN(P2_U3283) );
  AND2_X1 U16902 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15780), .ZN(P2_U3282) );
  AND2_X1 U16903 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15780), .ZN(P2_U3281) );
  AND2_X1 U16904 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15780), .ZN(P2_U3280) );
  AND2_X1 U16905 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15780), .ZN(P2_U3279) );
  AND2_X1 U16906 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15780), .ZN(P2_U3278) );
  AND2_X1 U16907 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15780), .ZN(P2_U3277) );
  AND2_X1 U16908 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15780), .ZN(P2_U3276) );
  AND2_X1 U16909 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15780), .ZN(P2_U3275) );
  AND2_X1 U16910 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15780), .ZN(P2_U3274) );
  AND2_X1 U16911 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15780), .ZN(P2_U3273) );
  AND2_X1 U16912 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15780), .ZN(P2_U3272) );
  AND2_X1 U16913 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15780), .ZN(P2_U3271) );
  AND2_X1 U16914 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15780), .ZN(P2_U3270) );
  AND2_X1 U16915 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15780), .ZN(P2_U3269) );
  AND2_X1 U16916 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15780), .ZN(P2_U3268) );
  AND2_X1 U16917 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15780), .ZN(P2_U3267) );
  AND2_X1 U16918 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15780), .ZN(P2_U3266) );
  NOR2_X1 U16919 ( .A1(n15800), .A2(P2_U3947), .ZN(P2_U3087) );
  NOR2_X1 U16920 ( .A1(P3_U3897), .A2(n15961), .ZN(P3_U3150) );
  INV_X1 U16921 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15782) );
  AOI22_X1 U16922 ( .A1(n15784), .A2(n15783), .B1(n15782), .B2(n15781), .ZN(
        P2_U3416) );
  INV_X1 U16923 ( .A(n15785), .ZN(n15787) );
  OAI21_X1 U16924 ( .B1(n15787), .B2(n15786), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15788) );
  OAI21_X1 U16925 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15788), .ZN(n15799) );
  NAND2_X1 U16926 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n15792) );
  INV_X1 U16927 ( .A(n15789), .ZN(n15791) );
  AOI211_X1 U16928 ( .C1(n15792), .C2(n15791), .A(n15790), .B(n15813), .ZN(
        n15797) );
  AOI211_X1 U16929 ( .C1(n15795), .C2(n15794), .A(n15793), .B(n15817), .ZN(
        n15796) );
  AOI211_X1 U16930 ( .C1(n15800), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n15797), .B(
        n15796), .ZN(n15798) );
  NAND2_X1 U16931 ( .A1(n15799), .A2(n15798), .ZN(P2_U3215) );
  AOI22_X1 U16932 ( .A1(n15800), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n15811) );
  AOI211_X1 U16933 ( .C1(n15803), .C2(n15802), .A(n15801), .B(n15813), .ZN(
        n15808) );
  AOI211_X1 U16934 ( .C1(n15806), .C2(n15805), .A(n15804), .B(n15817), .ZN(
        n15807) );
  AOI211_X1 U16935 ( .C1(n15838), .C2(n15809), .A(n15808), .B(n15807), .ZN(
        n15810) );
  NAND2_X1 U16936 ( .A1(n15811), .A2(n15810), .ZN(P2_U3216) );
  INV_X1 U16937 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n15825) );
  AOI211_X1 U16938 ( .C1(n15815), .C2(n15814), .A(n15813), .B(n15812), .ZN(
        n15821) );
  AOI211_X1 U16939 ( .C1(n15819), .C2(n15818), .A(n15817), .B(n15816), .ZN(
        n15820) );
  AOI211_X1 U16940 ( .C1(n15838), .C2(n15822), .A(n15821), .B(n15820), .ZN(
        n15824) );
  NAND2_X1 U16941 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n15823) );
  OAI211_X1 U16942 ( .C1(n15825), .C2(n15844), .A(n15824), .B(n15823), .ZN(
        P2_U3222) );
  INV_X1 U16943 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15899) );
  AOI21_X1 U16944 ( .B1(n15828), .B2(n15827), .A(n15826), .ZN(n15829) );
  NAND2_X1 U16945 ( .A1(n15830), .A2(n15829), .ZN(n15841) );
  AOI21_X1 U16946 ( .B1(n15833), .B2(n15832), .A(n15831), .ZN(n15834) );
  NAND2_X1 U16947 ( .A1(n15835), .A2(n15834), .ZN(n15840) );
  INV_X1 U16948 ( .A(n15836), .ZN(n15837) );
  NAND2_X1 U16949 ( .A1(n15838), .A2(n15837), .ZN(n15839) );
  NAND2_X1 U16950 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n15842)
         );
  OAI211_X1 U16951 ( .C1(n15899), .C2(n15844), .A(n15843), .B(n15842), .ZN(
        P2_U3229) );
  AOI21_X1 U16952 ( .B1(n15846), .B2(P1_REG1_REG_15__SCAN_IN), .A(n15845), 
        .ZN(n15851) );
  AOI21_X1 U16953 ( .B1(n15848), .B2(P1_REG2_REG_15__SCAN_IN), .A(n15847), 
        .ZN(n15849) );
  OAI222_X1 U16954 ( .A1(n16022), .A2(n15853), .B1(n15852), .B2(n15851), .C1(
        n16423), .C2(n15849), .ZN(n15854) );
  INV_X1 U16955 ( .A(n15854), .ZN(n15856) );
  OAI211_X1 U16956 ( .C1(n15857), .C2(n16028), .A(n15856), .B(n15855), .ZN(
        P1_U3258) );
  AOI21_X1 U16957 ( .B1(n15859), .B2(n15858), .A(n7441), .ZN(SUB_1596_U53) );
  NOR2_X1 U16958 ( .A1(n15861), .A2(n15860), .ZN(n15862) );
  XOR2_X1 U16959 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n15862), .Z(SUB_1596_U61) );
  XOR2_X1 U16960 ( .A(n15864), .B(n15863), .Z(SUB_1596_U60) );
  XOR2_X1 U16961 ( .A(n15866), .B(n15865), .Z(SUB_1596_U59) );
  XOR2_X1 U16962 ( .A(n15867), .B(P2_ADDR_REG_5__SCAN_IN), .Z(SUB_1596_U58) );
  XNOR2_X1 U16963 ( .A(n15869), .B(n15868), .ZN(SUB_1596_U56) );
  NOR2_X1 U16964 ( .A1(n15871), .A2(n15870), .ZN(n15872) );
  XOR2_X1 U16965 ( .A(n15872), .B(P2_ADDR_REG_8__SCAN_IN), .Z(SUB_1596_U55) );
  NOR2_X1 U16966 ( .A1(n15874), .A2(n15873), .ZN(n15875) );
  XOR2_X1 U16967 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n15875), .Z(SUB_1596_U54) );
  AOI21_X1 U16968 ( .B1(n15878), .B2(n15877), .A(n15876), .ZN(n15879) );
  XOR2_X1 U16969 ( .A(n15879), .B(P2_ADDR_REG_10__SCAN_IN), .Z(SUB_1596_U70)
         );
  AOI21_X1 U16970 ( .B1(n15882), .B2(n15881), .A(n15880), .ZN(n15883) );
  XOR2_X1 U16971 ( .A(n15883), .B(P2_ADDR_REG_11__SCAN_IN), .Z(SUB_1596_U69)
         );
  AOI21_X1 U16972 ( .B1(n15886), .B2(n15885), .A(n15884), .ZN(n15887) );
  XOR2_X1 U16973 ( .A(n15887), .B(P2_ADDR_REG_12__SCAN_IN), .Z(SUB_1596_U68)
         );
  AOI21_X1 U16974 ( .B1(n15890), .B2(n15889), .A(n15888), .ZN(n15891) );
  XOR2_X1 U16975 ( .A(n15891), .B(P2_ADDR_REG_13__SCAN_IN), .Z(SUB_1596_U67)
         );
  AOI21_X1 U16976 ( .B1(n15894), .B2(n15893), .A(n15892), .ZN(n15895) );
  XOR2_X1 U16977 ( .A(n15895), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  NOR2_X1 U16978 ( .A1(n15897), .A2(n15896), .ZN(n15898) );
  XNOR2_X1 U16979 ( .A(n15899), .B(n15898), .ZN(SUB_1596_U65) );
  XNOR2_X1 U16980 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n15900), .ZN(SUB_1596_U64)
         );
  AOI22_X1 U16981 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n15905), .B1(n15904), 
        .B2(n15903), .ZN(n15913) );
  INV_X1 U16982 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15915) );
  NAND2_X1 U16983 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n15915), .ZN(n15906) );
  OAI21_X1 U16984 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n15915), .A(n15906), 
        .ZN(n15912) );
  XNOR2_X1 U16985 ( .A(n15913), .B(n15912), .ZN(n15908) );
  XOR2_X1 U16986 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n15907), .Z(SUB_1596_U62)
         );
  NAND2_X1 U16987 ( .A1(n15909), .A2(n15908), .ZN(n15910) );
  XNOR2_X1 U16988 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n15911) );
  NOR2_X1 U16989 ( .A1(n15913), .A2(n15912), .ZN(n15914) );
  AOI21_X1 U16990 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n15915), .A(n15914), 
        .ZN(n15916) );
  XOR2_X1 U16991 ( .A(n15917), .B(P2_ADDR_REG_6__SCAN_IN), .Z(SUB_1596_U57) );
  OAI21_X1 U16992 ( .B1(n15919), .B2(n7441), .A(n15918), .ZN(n15920) );
  XNOR2_X1 U16993 ( .A(n15920), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(SUB_1596_U5)
         );
  AOI21_X1 U16994 ( .B1(n15923), .B2(n15922), .A(n15921), .ZN(n15939) );
  XNOR2_X1 U16995 ( .A(n15925), .B(n15924), .ZN(n15932) );
  NOR2_X1 U16996 ( .A1(n15984), .A2(n15926), .ZN(n15930) );
  OAI21_X1 U16997 ( .B1(n15982), .B2(n15928), .A(n15927), .ZN(n15929) );
  AOI211_X1 U16998 ( .C1(n15932), .C2(n15931), .A(n15930), .B(n15929), .ZN(
        n15938) );
  AOI21_X1 U16999 ( .B1(n15934), .B2(n15933), .A(n15991), .ZN(n15936) );
  NAND2_X1 U17000 ( .A1(n15936), .A2(n15935), .ZN(n15937) );
  OAI211_X1 U17001 ( .C1(n15939), .C2(n15999), .A(n15938), .B(n15937), .ZN(
        P3_U3194) );
  AOI21_X1 U17002 ( .B1(n15942), .B2(n15941), .A(n15940), .ZN(n15957) );
  OAI22_X1 U17003 ( .A1(n15984), .A2(n15944), .B1(n15982), .B2(n15943), .ZN(
        n15954) );
  AOI21_X1 U17004 ( .B1(n15947), .B2(n15946), .A(n15945), .ZN(n15952) );
  AOI21_X1 U17005 ( .B1(n15950), .B2(n15949), .A(n15948), .ZN(n15951) );
  OAI22_X1 U17006 ( .A1(n15952), .A2(n15993), .B1(n15951), .B2(n15991), .ZN(
        n15953) );
  NOR3_X1 U17007 ( .A1(n15955), .A2(n15954), .A3(n15953), .ZN(n15956) );
  OAI21_X1 U17008 ( .B1(n15957), .B2(n15999), .A(n15956), .ZN(P3_U3195) );
  NOR2_X1 U17009 ( .A1(n15984), .A2(n15958), .ZN(n15959) );
  AOI211_X1 U17010 ( .C1(P3_ADDR_REG_14__SCAN_IN), .C2(n15961), .A(n15960), 
        .B(n15959), .ZN(n15977) );
  AOI21_X1 U17011 ( .B1(n15964), .B2(n15963), .A(n15962), .ZN(n15965) );
  OR2_X1 U17012 ( .A1(n15965), .A2(n15993), .ZN(n15976) );
  OAI221_X1 U17013 ( .B1(n15969), .B2(n15968), .C1(n15969), .C2(n15967), .A(
        n15966), .ZN(n15975) );
  OAI211_X1 U17014 ( .C1(n15973), .C2(n15972), .A(n15971), .B(n15970), .ZN(
        n15974) );
  NAND4_X1 U17015 ( .A1(n15977), .A2(n15976), .A3(n15975), .A4(n15974), .ZN(
        P3_U3196) );
  AOI21_X1 U17016 ( .B1(n15980), .B2(n15979), .A(n15978), .ZN(n16000) );
  OAI22_X1 U17017 ( .A1(n15984), .A2(n15983), .B1(n15982), .B2(n15981), .ZN(
        n15996) );
  AOI21_X1 U17018 ( .B1(n15987), .B2(n15986), .A(n15985), .ZN(n15994) );
  AOI21_X1 U17019 ( .B1(n15990), .B2(n15989), .A(n15988), .ZN(n15992) );
  OAI22_X1 U17020 ( .A1(n15994), .A2(n15993), .B1(n15992), .B2(n15991), .ZN(
        n15995) );
  NOR3_X1 U17021 ( .A1(n15997), .A2(n15996), .A3(n15995), .ZN(n15998) );
  OAI21_X1 U17022 ( .B1(n16000), .B2(n15999), .A(n15998), .ZN(P3_U3197) );
  INV_X1 U17023 ( .A(P1_RD_REG_SCAN_IN), .ZN(n16002) );
  OAI221_X1 U17024 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(n8796), .C2(n16002), .A(n16001), .ZN(U29) );
  INV_X1 U17025 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n16027) );
  MUX2_X1 U17026 ( .A(n16004), .B(P1_REG2_REG_4__SCAN_IN), .S(n16003), .Z(
        n16007) );
  INV_X1 U17027 ( .A(n16005), .ZN(n16006) );
  NAND2_X1 U17028 ( .A1(n16007), .A2(n16006), .ZN(n16010) );
  OAI211_X1 U17029 ( .C1(n16011), .C2(n16010), .A(n7422), .B(n16008), .ZN(
        n16020) );
  INV_X1 U17030 ( .A(n16012), .ZN(n16017) );
  NAND3_X1 U17031 ( .A1(n16015), .A2(n16014), .A3(n16013), .ZN(n16016) );
  NAND3_X1 U17032 ( .A1(n16018), .A2(n16017), .A3(n16016), .ZN(n16019) );
  OAI211_X1 U17033 ( .C1(n16022), .C2(n16021), .A(n16020), .B(n16019), .ZN(
        n16023) );
  NOR2_X1 U17034 ( .A1(n16024), .A2(n16023), .ZN(n16026) );
  OAI211_X1 U17035 ( .C1(n16028), .C2(n16027), .A(n16026), .B(n16025), .ZN(
        P1_U3247) );
  INV_X1 U17036 ( .A(n16044), .ZN(n16034) );
  INV_X1 U17037 ( .A(n16029), .ZN(n16030) );
  NOR2_X1 U17038 ( .A1(n16031), .A2(n16030), .ZN(n16042) );
  OAI21_X1 U17039 ( .B1(n16372), .B2(n16194), .A(n16034), .ZN(n16033) );
  NAND2_X1 U17040 ( .A1(n16033), .A2(n16032), .ZN(n16040) );
  AOI211_X1 U17041 ( .C1(n16332), .C2(n16034), .A(n16042), .B(n16040), .ZN(
        n16037) );
  AOI22_X1 U17042 ( .A1(n16387), .A2(n16037), .B1(n16035), .B2(n16385), .ZN(
        P1_U3528) );
  INV_X1 U17043 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n16036) );
  AOI22_X1 U17044 ( .A1(n16391), .A2(n16037), .B1(n16036), .B2(n16388), .ZN(
        P1_U3459) );
  NAND2_X1 U17045 ( .A1(n16039), .A2(n16038), .ZN(n16041) );
  AOI21_X1 U17046 ( .B1(n16042), .B2(n16041), .A(n16040), .ZN(n16049) );
  INV_X1 U17047 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n16048) );
  OAI22_X1 U17048 ( .A1(n16045), .A2(n16044), .B1(n16043), .B2(n16161), .ZN(
        n16046) );
  INV_X1 U17049 ( .A(n16046), .ZN(n16047) );
  OAI221_X1 U17050 ( .B1(n16347), .B2(n16049), .C1(n16159), .C2(n16048), .A(
        n16047), .ZN(P1_U3293) );
  XNOR2_X1 U17051 ( .A(n16051), .B(n16050), .ZN(n16065) );
  OAI22_X1 U17052 ( .A1(n16053), .A2(n16107), .B1(n16052), .B2(n16101), .ZN(
        n16060) );
  NAND3_X1 U17053 ( .A1(n16056), .A2(n16055), .A3(n16054), .ZN(n16058) );
  AOI21_X1 U17054 ( .B1(n16058), .B2(n16103), .A(n16057), .ZN(n16059) );
  AOI211_X1 U17055 ( .C1(n16229), .C2(n16065), .A(n16060), .B(n16059), .ZN(
        n16064) );
  INV_X1 U17056 ( .A(n16274), .ZN(n16299) );
  AOI22_X1 U17057 ( .A1(n16065), .A2(n16299), .B1(n16200), .B2(n8825), .ZN(
        n16061) );
  AND2_X1 U17058 ( .A1(n16064), .A2(n16061), .ZN(n16063) );
  AOI22_X1 U17059 ( .A1(n16407), .A2(n16063), .B1(n8813), .B2(n9309), .ZN(
        P3_U3460) );
  INV_X1 U17060 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n16062) );
  AOI22_X1 U17061 ( .A1(n16410), .A2(n16063), .B1(n16062), .B2(n16415), .ZN(
        P3_U3393) );
  INV_X1 U17062 ( .A(n16064), .ZN(n16068) );
  NAND2_X1 U17063 ( .A1(n16065), .A2(n16120), .ZN(n16066) );
  OAI211_X1 U17064 ( .C1(n7738), .C2(n16115), .A(n16066), .B(n16121), .ZN(
        n16067) );
  OAI22_X1 U17065 ( .A1(n16068), .A2(n16067), .B1(P3_REG2_REG_1__SCAN_IN), 
        .B2(n16121), .ZN(n16069) );
  OAI21_X1 U17066 ( .B1(n16070), .B2(n16113), .A(n16069), .ZN(P3_U3232) );
  XNOR2_X1 U17067 ( .A(n16073), .B(n16071), .ZN(n16093) );
  INV_X1 U17068 ( .A(n16093), .ZN(n16081) );
  XNOR2_X1 U17069 ( .A(n16072), .B(n16073), .ZN(n16074) );
  NOR2_X1 U17070 ( .A1(n16074), .A2(n16379), .ZN(n16075) );
  AOI211_X1 U17071 ( .C1(n16372), .C2(n16093), .A(n16076), .B(n16075), .ZN(
        n16096) );
  AOI211_X1 U17072 ( .C1(n16078), .C2(n16079), .A(n16142), .B(n8187), .ZN(
        n16092) );
  AOI211_X1 U17073 ( .C1(n16366), .C2(n16079), .A(n16085), .B(n16092), .ZN(
        n16080) );
  OAI211_X1 U17074 ( .C1(n16081), .C2(n16369), .A(n16096), .B(n16080), .ZN(
        n16082) );
  INV_X1 U17075 ( .A(n16082), .ZN(n16084) );
  AOI22_X1 U17076 ( .A1(n16387), .A2(n16084), .B1(n9914), .B2(n16385), .ZN(
        P1_U3529) );
  INV_X1 U17077 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n16083) );
  AOI22_X1 U17078 ( .A1(n16391), .A2(n16084), .B1(n16083), .B2(n16388), .ZN(
        P1_U3462) );
  AOI22_X1 U17079 ( .A1(n16086), .A2(n16085), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n16336), .ZN(n16089) );
  INV_X1 U17080 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n16087) );
  OR2_X1 U17081 ( .A1(n16159), .A2(n16087), .ZN(n16088) );
  OAI211_X1 U17082 ( .C1(n16163), .C2(n16090), .A(n16089), .B(n16088), .ZN(
        n16091) );
  INV_X1 U17083 ( .A(n16091), .ZN(n16095) );
  AOI22_X1 U17084 ( .A1(n16342), .A2(n16093), .B1(n16341), .B2(n16092), .ZN(
        n16094) );
  OAI211_X1 U17085 ( .C1(n16347), .C2(n16096), .A(n16095), .B(n16094), .ZN(
        P1_U3292) );
  XNOR2_X1 U17086 ( .A(n16098), .B(n16097), .ZN(n16108) );
  XNOR2_X1 U17087 ( .A(n16100), .B(n16099), .ZN(n16119) );
  OAI22_X1 U17088 ( .A1(n16104), .A2(n16103), .B1(n16102), .B2(n16101), .ZN(
        n16105) );
  AOI21_X1 U17089 ( .B1(n16119), .B2(n16229), .A(n16105), .ZN(n16106) );
  OAI21_X1 U17090 ( .B1(n16108), .B2(n16107), .A(n16106), .ZN(n16117) );
  INV_X1 U17091 ( .A(n16119), .ZN(n16109) );
  OAI22_X1 U17092 ( .A1(n16109), .A2(n16274), .B1(n16311), .B2(n16116), .ZN(
        n16110) );
  NOR2_X1 U17093 ( .A1(n16117), .A2(n16110), .ZN(n16112) );
  AOI22_X1 U17094 ( .A1(n16407), .A2(n16112), .B1(n8826), .B2(n9309), .ZN(
        P3_U3461) );
  INV_X1 U17095 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n16111) );
  AOI22_X1 U17096 ( .A1(n16410), .A2(n16112), .B1(n16111), .B2(n16415), .ZN(
        P3_U3396) );
  OAI22_X1 U17097 ( .A1(n16116), .A2(n16115), .B1(n16114), .B2(n16113), .ZN(
        n16118) );
  AOI211_X1 U17098 ( .C1(n16120), .C2(n16119), .A(n16118), .B(n16117), .ZN(
        n16122) );
  AOI22_X1 U17099 ( .A1(n16123), .A2(n8827), .B1(n16122), .B2(n16121), .ZN(
        P3_U3231) );
  INV_X1 U17100 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n16124) );
  AOI22_X1 U17101 ( .A1(n16391), .A2(n16125), .B1(n16124), .B2(n16388), .ZN(
        P1_U3465) );
  OAI21_X1 U17102 ( .B1(n16127), .B2(n16353), .A(n16126), .ZN(n16129) );
  AOI211_X1 U17103 ( .C1(n16348), .C2(n16130), .A(n16129), .B(n16128), .ZN(
        n16132) );
  AOI22_X1 U17104 ( .A1(n16358), .A2(n16132), .B1(n9563), .B2(n16357), .ZN(
        P2_U3501) );
  INV_X1 U17105 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n16131) );
  AOI22_X1 U17106 ( .A1(n14668), .A2(n16132), .B1(n16131), .B2(n16359), .ZN(
        P2_U3436) );
  AOI22_X1 U17107 ( .A1(n16134), .A2(n16407), .B1(n16259), .B2(n16133), .ZN(
        n16135) );
  OAI21_X1 U17108 ( .B1(n16407), .B2(n8837), .A(n16135), .ZN(P3_U3462) );
  XNOR2_X1 U17109 ( .A(n16136), .B(n16137), .ZN(n16157) );
  XNOR2_X1 U17110 ( .A(n16138), .B(n16137), .ZN(n16140) );
  AOI21_X1 U17111 ( .B1(n16140), .B2(n16194), .A(n16139), .ZN(n16156) );
  INV_X1 U17112 ( .A(n16141), .ZN(n16146) );
  AOI21_X1 U17113 ( .B1(n16144), .B2(n16143), .A(n16142), .ZN(n16145) );
  NAND2_X1 U17114 ( .A1(n16146), .A2(n16145), .ZN(n16153) );
  OR2_X1 U17115 ( .A1(n16162), .A2(n16378), .ZN(n16147) );
  AND2_X1 U17116 ( .A1(n16153), .A2(n16147), .ZN(n16148) );
  OAI211_X1 U17117 ( .C1(n16157), .C2(n16190), .A(n16156), .B(n16148), .ZN(
        n16149) );
  INV_X1 U17118 ( .A(n16149), .ZN(n16152) );
  AOI22_X1 U17119 ( .A1(n16387), .A2(n16152), .B1(n16150), .B2(n16385), .ZN(
        P1_U3531) );
  INV_X1 U17120 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n16151) );
  AOI22_X1 U17121 ( .A1(n16391), .A2(n16152), .B1(n16151), .B2(n16388), .ZN(
        P1_U3468) );
  INV_X1 U17122 ( .A(n16157), .ZN(n16155) );
  INV_X1 U17123 ( .A(n16153), .ZN(n16154) );
  AOI22_X1 U17124 ( .A1(n16342), .A2(n16155), .B1(n16341), .B2(n16154), .ZN(
        n16167) );
  OAI21_X1 U17125 ( .B1(n16158), .B2(n16157), .A(n16156), .ZN(n16160) );
  MUX2_X1 U17126 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n16160), .S(n16159), .Z(
        n16165) );
  OAI22_X1 U17127 ( .A1(n16163), .A2(n16162), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n16161), .ZN(n16164) );
  NOR2_X1 U17128 ( .A1(n16165), .A2(n16164), .ZN(n16166) );
  NAND2_X1 U17129 ( .A1(n16167), .A2(n16166), .ZN(P1_U3290) );
  AOI21_X1 U17130 ( .B1(n16170), .B2(n16169), .A(n16168), .ZN(n16171) );
  OAI211_X1 U17131 ( .C1(n16262), .C2(n16173), .A(n16172), .B(n16171), .ZN(
        n16174) );
  INV_X1 U17132 ( .A(n16174), .ZN(n16176) );
  AOI22_X1 U17133 ( .A1(n16358), .A2(n16176), .B1(n9564), .B2(n16357), .ZN(
        P2_U3502) );
  INV_X1 U17134 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n16175) );
  AOI22_X1 U17135 ( .A1(n14668), .A2(n16176), .B1(n16175), .B2(n16359), .ZN(
        P2_U3439) );
  AOI21_X1 U17136 ( .B1(n16178), .B2(n16274), .A(n16177), .ZN(n16181) );
  INV_X1 U17137 ( .A(n16179), .ZN(n16180) );
  AOI211_X1 U17138 ( .C1(n16200), .C2(n16182), .A(n16181), .B(n16180), .ZN(
        n16184) );
  AOI22_X1 U17139 ( .A1(n16407), .A2(n16184), .B1(n10294), .B2(n9309), .ZN(
        P3_U3463) );
  INV_X1 U17140 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n16183) );
  AOI22_X1 U17141 ( .A1(n16410), .A2(n16184), .B1(n16183), .B2(n16415), .ZN(
        P3_U3402) );
  INV_X1 U17142 ( .A(n16185), .ZN(n16188) );
  INV_X1 U17143 ( .A(n16186), .ZN(n16187) );
  OAI211_X1 U17144 ( .C1(n16189), .C2(n16378), .A(n16188), .B(n16187), .ZN(
        n16193) );
  NOR2_X1 U17145 ( .A1(n16191), .A2(n16190), .ZN(n16192) );
  AOI211_X1 U17146 ( .C1(n16195), .C2(n16194), .A(n16193), .B(n16192), .ZN(
        n16198) );
  AOI22_X1 U17147 ( .A1(n16387), .A2(n16198), .B1(n16196), .B2(n16385), .ZN(
        P1_U3532) );
  INV_X1 U17148 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n16197) );
  AOI22_X1 U17149 ( .A1(n16391), .A2(n16198), .B1(n16197), .B2(n16388), .ZN(
        P1_U3471) );
  AOI22_X1 U17150 ( .A1(n16201), .A2(n16316), .B1(n16200), .B2(n16199), .ZN(
        n16202) );
  AND2_X1 U17151 ( .A1(n16203), .A2(n16202), .ZN(n16205) );
  AOI22_X1 U17152 ( .A1(n16407), .A2(n16205), .B1(n8861), .B2(n9309), .ZN(
        P3_U3464) );
  INV_X1 U17153 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n16204) );
  AOI22_X1 U17154 ( .A1(n16410), .A2(n16205), .B1(n16204), .B2(n16415), .ZN(
        P3_U3405) );
  INV_X1 U17155 ( .A(n16206), .ZN(n16207) );
  OAI21_X1 U17156 ( .B1(n16208), .B2(n16378), .A(n16207), .ZN(n16210) );
  AOI211_X1 U17157 ( .C1(n16332), .C2(n16211), .A(n16210), .B(n16209), .ZN(
        n16214) );
  AOI22_X1 U17158 ( .A1(n16387), .A2(n16214), .B1(n16212), .B2(n16385), .ZN(
        P1_U3533) );
  INV_X1 U17159 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n16213) );
  AOI22_X1 U17160 ( .A1(n16391), .A2(n16214), .B1(n16213), .B2(n16388), .ZN(
        P1_U3474) );
  INV_X1 U17161 ( .A(n16219), .ZN(n16216) );
  OAI22_X1 U17162 ( .A1(n16216), .A2(n16274), .B1(n16215), .B2(n16311), .ZN(
        n16218) );
  AOI211_X1 U17163 ( .C1(n16229), .C2(n16219), .A(n16218), .B(n16217), .ZN(
        n16221) );
  AOI22_X1 U17164 ( .A1(n16407), .A2(n16221), .B1(n8878), .B2(n9309), .ZN(
        P3_U3465) );
  INV_X1 U17165 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n16220) );
  AOI22_X1 U17166 ( .A1(n16410), .A2(n16221), .B1(n16220), .B2(n16415), .ZN(
        P3_U3408) );
  AOI222_X1 U17167 ( .A1(n16223), .A2(n16303), .B1(P2_REG2_REG_6__SCAN_IN), 
        .B2(n16405), .C1(n16394), .C2(n16222), .ZN(n16227) );
  AOI22_X1 U17168 ( .A1(n16225), .A2(n16401), .B1(n16306), .B2(n16224), .ZN(
        n16226) );
  OAI211_X1 U17169 ( .C1(n16405), .C2(n16228), .A(n16227), .B(n16226), .ZN(
        P2_U3259) );
  INV_X1 U17170 ( .A(n16232), .ZN(n16230) );
  AND2_X1 U17171 ( .A1(n16230), .A2(n16229), .ZN(n16234) );
  OAI22_X1 U17172 ( .A1(n16232), .A2(n16274), .B1(n16311), .B2(n16231), .ZN(
        n16233) );
  NOR3_X1 U17173 ( .A1(n16235), .A2(n16234), .A3(n16233), .ZN(n16238) );
  AOI22_X1 U17174 ( .A1(n16407), .A2(n16238), .B1(n16236), .B2(n9309), .ZN(
        P3_U3466) );
  INV_X1 U17175 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n16237) );
  AOI22_X1 U17176 ( .A1(n16410), .A2(n16238), .B1(n16237), .B2(n16415), .ZN(
        P3_U3411) );
  AOI222_X1 U17177 ( .A1(n16240), .A2(n16337), .B1(P1_REG2_REG_7__SCAN_IN), 
        .B2(n16347), .C1(n16336), .C2(n16239), .ZN(n16244) );
  AOI22_X1 U17178 ( .A1(n16242), .A2(n16342), .B1(n16341), .B2(n16241), .ZN(
        n16243) );
  OAI211_X1 U17179 ( .C1(n16347), .C2(n16245), .A(n16244), .B(n16243), .ZN(
        P1_U3286) );
  INV_X1 U17180 ( .A(n16246), .ZN(n16251) );
  NAND2_X1 U17181 ( .A1(n16247), .A2(n16306), .ZN(n16250) );
  AOI22_X1 U17182 ( .A1(n16405), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n16248), 
        .B2(n16394), .ZN(n16249) );
  OAI211_X1 U17183 ( .C1(n16251), .C2(n16398), .A(n16250), .B(n16249), .ZN(
        n16252) );
  AOI21_X1 U17184 ( .B1(n16253), .B2(n16401), .A(n16252), .ZN(n16254) );
  OAI21_X1 U17185 ( .B1(n16405), .B2(n16255), .A(n16254), .ZN(P2_U3258) );
  OAI21_X1 U17186 ( .B1(n16257), .B2(n16311), .A(n16256), .ZN(n16260) );
  AOI22_X1 U17187 ( .A1(n16260), .A2(n16407), .B1(n16259), .B2(n16258), .ZN(
        n16261) );
  OAI21_X1 U17188 ( .B1(n16407), .B2(n8909), .A(n16261), .ZN(P3_U3467) );
  NOR2_X1 U17189 ( .A1(n16263), .A2(n16262), .ZN(n16270) );
  INV_X1 U17190 ( .A(n16264), .ZN(n16265) );
  OAI21_X1 U17191 ( .B1(n8270), .B2(n16353), .A(n16265), .ZN(n16268) );
  INV_X1 U17192 ( .A(n16266), .ZN(n16267) );
  AOI211_X1 U17193 ( .C1(n16270), .C2(n16269), .A(n16268), .B(n16267), .ZN(
        n16272) );
  AOI22_X1 U17194 ( .A1(n16358), .A2(n16272), .B1(n10193), .B2(n16357), .ZN(
        P2_U3507) );
  INV_X1 U17195 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n16271) );
  AOI22_X1 U17196 ( .A1(n14668), .A2(n16272), .B1(n16271), .B2(n16359), .ZN(
        P2_U3454) );
  OAI22_X1 U17197 ( .A1(n16275), .A2(n16274), .B1(n16311), .B2(n16273), .ZN(
        n16276) );
  NOR2_X1 U17198 ( .A1(n16277), .A2(n16276), .ZN(n16280) );
  AOI22_X1 U17199 ( .A1(n16407), .A2(n16280), .B1(n16278), .B2(n9309), .ZN(
        P3_U3468) );
  INV_X1 U17200 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n16279) );
  AOI22_X1 U17201 ( .A1(n16410), .A2(n16280), .B1(n16279), .B2(n16415), .ZN(
        P3_U3417) );
  OAI21_X1 U17202 ( .B1(n16282), .B2(n16378), .A(n16281), .ZN(n16284) );
  AOI211_X1 U17203 ( .C1(n16332), .C2(n16285), .A(n16284), .B(n16283), .ZN(
        n16288) );
  AOI22_X1 U17204 ( .A1(n16387), .A2(n16288), .B1(n16286), .B2(n16385), .ZN(
        P1_U3537) );
  INV_X1 U17205 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n16287) );
  AOI22_X1 U17206 ( .A1(n16391), .A2(n16288), .B1(n16287), .B2(n16388), .ZN(
        P1_U3486) );
  INV_X1 U17207 ( .A(n16289), .ZN(n16292) );
  AOI22_X1 U17208 ( .A1(n16292), .A2(n16291), .B1(SI_10_), .B2(n16290), .ZN(
        n16293) );
  OAI21_X1 U17209 ( .B1(P3_U3151), .B2(n16294), .A(n16293), .ZN(P3_U3285) );
  NOR2_X1 U17210 ( .A1(n16295), .A2(n16311), .ZN(n16297) );
  AOI211_X1 U17211 ( .C1(n16299), .C2(n16298), .A(n16297), .B(n16296), .ZN(
        n16301) );
  AOI22_X1 U17212 ( .A1(n16407), .A2(n16301), .B1(n8943), .B2(n9309), .ZN(
        P3_U3469) );
  INV_X1 U17213 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n16300) );
  AOI22_X1 U17214 ( .A1(n16410), .A2(n16301), .B1(n16300), .B2(n16415), .ZN(
        P3_U3420) );
  AOI222_X1 U17215 ( .A1(n16304), .A2(n16303), .B1(P2_REG2_REG_10__SCAN_IN), 
        .B2(n16405), .C1(n16394), .C2(n16302), .ZN(n16309) );
  AOI22_X1 U17216 ( .A1(n16307), .A2(n16401), .B1(n16306), .B2(n16305), .ZN(
        n16308) );
  OAI211_X1 U17217 ( .C1(n16405), .C2(n16310), .A(n16309), .B(n16308), .ZN(
        P2_U3255) );
  NOR2_X1 U17218 ( .A1(n16312), .A2(n16311), .ZN(n16314) );
  AOI211_X1 U17219 ( .C1(n16316), .C2(n16315), .A(n16314), .B(n16313), .ZN(
        n16319) );
  AOI22_X1 U17220 ( .A1(n16407), .A2(n16319), .B1(n16317), .B2(n9309), .ZN(
        P3_U3470) );
  INV_X1 U17221 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n16318) );
  AOI22_X1 U17222 ( .A1(n16410), .A2(n16319), .B1(n16318), .B2(n16415), .ZN(
        P3_U3423) );
  XOR2_X1 U17223 ( .A(n16320), .B(n16325), .Z(n16343) );
  OAI211_X1 U17224 ( .C1(n16324), .C2(n16323), .A(n16322), .B(n16321), .ZN(
        n16339) );
  OAI21_X1 U17225 ( .B1(n16324), .B2(n16378), .A(n16339), .ZN(n16331) );
  XNOR2_X1 U17226 ( .A(n16326), .B(n16325), .ZN(n16328) );
  OAI21_X1 U17227 ( .B1(n16328), .B2(n16379), .A(n16327), .ZN(n16329) );
  AOI21_X1 U17228 ( .B1(n16343), .B2(n16372), .A(n16329), .ZN(n16346) );
  INV_X1 U17229 ( .A(n16346), .ZN(n16330) );
  AOI211_X1 U17230 ( .C1(n16332), .C2(n16343), .A(n16331), .B(n16330), .ZN(
        n16334) );
  AOI22_X1 U17231 ( .A1(n16387), .A2(n16334), .B1(n10051), .B2(n16385), .ZN(
        P1_U3539) );
  INV_X1 U17232 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n16333) );
  AOI22_X1 U17233 ( .A1(n16391), .A2(n16334), .B1(n16333), .B2(n16388), .ZN(
        P1_U3492) );
  AOI222_X1 U17234 ( .A1(n16338), .A2(n16337), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n16347), .C1(n16336), .C2(n16335), .ZN(n16345) );
  INV_X1 U17235 ( .A(n16339), .ZN(n16340) );
  AOI22_X1 U17236 ( .A1(n16343), .A2(n16342), .B1(n16341), .B2(n16340), .ZN(
        n16344) );
  OAI211_X1 U17237 ( .C1(n16347), .C2(n16346), .A(n16345), .B(n16344), .ZN(
        P1_U3282) );
  NAND3_X1 U17238 ( .A1(n16350), .A2(n16349), .A3(n16348), .ZN(n16352) );
  OAI211_X1 U17239 ( .C1(n16354), .C2(n16353), .A(n16352), .B(n16351), .ZN(
        n16355) );
  NOR2_X1 U17240 ( .A1(n16356), .A2(n16355), .ZN(n16361) );
  AOI22_X1 U17241 ( .A1(n16358), .A2(n16361), .B1(n10843), .B2(n16357), .ZN(
        P2_U3510) );
  INV_X1 U17242 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n16360) );
  AOI22_X1 U17243 ( .A1(n14668), .A2(n16361), .B1(n16360), .B2(n16359), .ZN(
        P2_U3463) );
  INV_X1 U17244 ( .A(n16368), .ZN(n16371) );
  AOI211_X1 U17245 ( .C1(n16366), .C2(n16365), .A(n16364), .B(n16363), .ZN(
        n16367) );
  OAI21_X1 U17246 ( .B1(n16369), .B2(n16368), .A(n16367), .ZN(n16370) );
  AOI21_X1 U17247 ( .B1(n16372), .B2(n16371), .A(n16370), .ZN(n16375) );
  AOI22_X1 U17248 ( .A1(n16387), .A2(n16375), .B1(n16373), .B2(n16385), .ZN(
        P1_U3540) );
  INV_X1 U17249 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n16374) );
  AOI22_X1 U17250 ( .A1(n16391), .A2(n16375), .B1(n16374), .B2(n16388), .ZN(
        P1_U3495) );
  OAI211_X1 U17251 ( .C1(n7671), .C2(n16378), .A(n16377), .B(n16376), .ZN(
        n16382) );
  NOR2_X1 U17252 ( .A1(n16380), .A2(n16379), .ZN(n16381) );
  AOI211_X1 U17253 ( .C1(n16384), .C2(n16383), .A(n16382), .B(n16381), .ZN(
        n16390) );
  AOI22_X1 U17254 ( .A1(n16387), .A2(n16390), .B1(n16386), .B2(n16385), .ZN(
        P1_U3541) );
  INV_X1 U17255 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n16389) );
  AOI22_X1 U17256 ( .A1(n16391), .A2(n16390), .B1(n16389), .B2(n16388), .ZN(
        P1_U3498) );
  INV_X1 U17257 ( .A(n16392), .ZN(n16399) );
  NAND2_X1 U17258 ( .A1(n16393), .A2(n16306), .ZN(n16397) );
  AOI22_X1 U17259 ( .A1(n16405), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n16395), 
        .B2(n16394), .ZN(n16396) );
  OAI211_X1 U17260 ( .C1(n16399), .C2(n16398), .A(n16397), .B(n16396), .ZN(
        n16400) );
  AOI21_X1 U17261 ( .B1(n16402), .B2(n16401), .A(n16400), .ZN(n16403) );
  OAI21_X1 U17262 ( .B1(n16405), .B2(n16404), .A(n16403), .ZN(P2_U3252) );
  AOI22_X1 U17263 ( .A1(n16409), .A2(n9313), .B1(P3_REG1_REG_30__SCAN_IN), 
        .B2(n9309), .ZN(n16408) );
  INV_X1 U17264 ( .A(n16406), .ZN(n16411) );
  NAND2_X1 U17265 ( .A1(n16411), .A2(n16407), .ZN(n16413) );
  NAND2_X1 U17266 ( .A1(n16408), .A2(n16413), .ZN(P3_U3489) );
  AOI22_X1 U17267 ( .A1(n16409), .A2(n9325), .B1(P3_REG0_REG_30__SCAN_IN), 
        .B2(n16415), .ZN(n16412) );
  NAND2_X1 U17268 ( .A1(n16411), .A2(n16410), .ZN(n16417) );
  NAND2_X1 U17269 ( .A1(n16412), .A2(n16417), .ZN(P3_U3457) );
  AOI22_X1 U17270 ( .A1(n16416), .A2(n9313), .B1(P3_REG1_REG_31__SCAN_IN), 
        .B2(n9309), .ZN(n16414) );
  NAND2_X1 U17271 ( .A1(n16414), .A2(n16413), .ZN(P3_U3490) );
  AOI22_X1 U17272 ( .A1(n16416), .A2(n9325), .B1(n16415), .B2(
        P3_REG0_REG_31__SCAN_IN), .ZN(n16418) );
  NAND2_X1 U17273 ( .A1(n16418), .A2(n16417), .ZN(P3_U3458) );
  AOI21_X1 U17274 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n16419) );
  OAI21_X1 U17275 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n16419), 
        .ZN(U28) );
  CLKBUF_X1 U7534 ( .A(n8874), .Z(n9080) );
  OR2_X1 U7545 ( .A1(n14505), .A2(n14537), .ZN(n14508) );
  INV_X1 U7564 ( .A(n7433), .ZN(n12399) );
  CLKBUF_X1 U7577 ( .A(n10763), .Z(n8025) );
  AOI22_X1 U7752 ( .A1(n14215), .A2(n14214), .B1(n8061), .B2(n14135), .ZN(
        n14137) );
  CLKBUF_X2 U7869 ( .A(n12685), .Z(n7426) );
  OR2_X1 U8319 ( .A1(n9924), .A2(n15245), .ZN(n16423) );
  INV_X2 U10056 ( .A(n16359), .ZN(n14668) );
endmodule

