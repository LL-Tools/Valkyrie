

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput0, keyinput1, keyinput2, 
        keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, 
        keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, 
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, 
        keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, 
        keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, 
        keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, 
        keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, 
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, 
        keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, 
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, 
        keyinput63 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859;

  OR2_X1 U3393 ( .A1(n5194), .A2(n3066), .ZN(n5325) );
  NOR2_X1 U3394 ( .A1(n4248), .A2(n2961), .ZN(n3558) );
  BUF_X2 U3395 ( .A(n3292), .Z(n4079) );
  BUF_X2 U3396 ( .A(n3168), .Z(n4052) );
  CLKBUF_X2 U3397 ( .A(n3263), .Z(n4051) );
  CLKBUF_X2 U3398 ( .A(n3258), .Z(n4072) );
  CLKBUF_X2 U3399 ( .A(n3198), .Z(n2946) );
  CLKBUF_X2 U3400 ( .A(n3328), .Z(n3293) );
  CLKBUF_X2 U3401 ( .A(n3173), .Z(n4551) );
  CLKBUF_X2 U3402 ( .A(n3189), .Z(n4070) );
  CLKBUF_X2 U3403 ( .A(n3333), .Z(n3281) );
  CLKBUF_X2 U3404 ( .A(n3154), .Z(n4057) );
  CLKBUF_X1 U3405 ( .A(n3165), .Z(n4624) );
  NAND2_X1 U3406 ( .A1(n3167), .A2(n3221), .ZN(n3214) );
  AND2_X2 U3407 ( .A1(n4441), .A2(n4547), .ZN(n3258) );
  AND2_X2 U3408 ( .A1(n3107), .A2(n4441), .ZN(n3327) );
  CLKBUF_X2 U3409 ( .A(n3184), .Z(n4071) );
  CLKBUF_X2 U3410 ( .A(n4027), .Z(n4078) );
  INV_X1 U3411 ( .A(n3532), .ZN(n3540) );
  BUF_X1 U3412 ( .A(n3228), .Z(n2961) );
  OR2_X1 U3413 ( .A1(n3179), .A2(n3178), .ZN(n4638) );
  AND4_X1 U3414 ( .A1(n3141), .A2(n3140), .A3(n3139), .A4(n3138), .ZN(n3142)
         );
  XNOR2_X1 U3416 ( .A(n3456), .B(n3455), .ZN(n3604) );
  NAND2_X1 U3417 ( .A1(n3470), .A2(n3469), .ZN(n3471) );
  INV_X1 U3418 ( .A(n6398), .ZN(n6327) );
  CLKBUF_X3 U3419 ( .A(n4158), .Z(n4145) );
  AND2_X1 U3420 ( .A1(n4631), .A2(n4724), .ZN(n4726) );
  AND4_X1 U3421 ( .A1(n3193), .A2(n3192), .A3(n3191), .A4(n3190), .ZN(n3206)
         );
  NAND2_X1 U3422 ( .A1(n5697), .A2(n2988), .ZN(n5690) );
  OR2_X1 U3423 ( .A1(n5376), .A2(n5377), .ZN(n5374) );
  INV_X1 U3424 ( .A(n3492), .ZN(n4296) );
  XNOR2_X1 U3425 ( .A(n3471), .B(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3086)
         );
  AND2_X1 U3426 ( .A1(n5549), .A2(n5178), .ZN(n6398) );
  OR2_X1 U3427 ( .A1(n4236), .A2(n5439), .ZN(n4423) );
  NOR2_X1 U3428 ( .A1(n6449), .A2(n6421), .ZN(n6448) );
  INV_X1 U3429 ( .A(n5762), .ZN(n6501) );
  INV_X1 U3430 ( .A(n6399), .ZN(n6375) );
  INV_X1 U3431 ( .A(n6346), .ZN(n6371) );
  NAND2_X1 U3432 ( .A1(n5762), .A2(n4465), .ZN(n6510) );
  AND2_X2 U3433 ( .A1(n4441), .A2(n4548), .ZN(n3189) );
  BUF_X4 U3435 ( .A(n3221), .Z(n3235) );
  NAND2_X2 U3436 ( .A1(n3123), .A2(n3122), .ZN(n3237) );
  NAND2_X2 U3437 ( .A1(n3143), .A2(n3142), .ZN(n3210) );
  XNOR2_X2 U3438 ( .A(n3423), .B(n3422), .ZN(n4578) );
  INV_X1 U3439 ( .A(n3449), .ZN(n2963) );
  INV_X1 U3440 ( .A(n5330), .ZN(n6397) );
  INV_X4 U3441 ( .A(n4296), .ZN(n5808) );
  NAND2_X2 U3442 ( .A1(n5921), .A2(n5923), .ZN(n5958) );
  INV_X1 U3443 ( .A(n6510), .ZN(n5764) );
  NOR2_X2 U3444 ( .A1(n5623), .A2(n3054), .ZN(n5603) );
  NAND2_X2 U34450 ( .A1(n3351), .A2(n3350), .ZN(n3553) );
  INV_X2 U34460 ( .A(n3404), .ZN(n3411) );
  NAND2_X2 U34470 ( .A1(n3113), .A2(n3112), .ZN(n3221) );
  AND4_X1 U34480 ( .A1(n3158), .A2(n3157), .A3(n3156), .A4(n3155), .ZN(n3164)
         );
  BUF_X2 U3449 ( .A(n4077), .Z(n2971) );
  NAND2_X1 U3450 ( .A1(n4295), .A2(n5698), .ZN(n5697) );
  AND3_X1 U34510 ( .A1(REIP_REG_21__SCAN_IN), .A2(REIP_REG_20__SCAN_IN), .A3(
        n5430), .ZN(n5392) );
  OR2_X1 U34520 ( .A1(n3750), .A2(n3749), .ZN(n5728) );
  AOI21_X1 U34530 ( .B1(n5277), .B2(n6541), .A(n2999), .ZN(n2998) );
  NAND2_X1 U3454 ( .A1(n5861), .A2(n5924), .ZN(n5952) );
  NAND2_X1 U34550 ( .A1(n3595), .A2(n4454), .ZN(n4585) );
  XNOR2_X1 U34560 ( .A(n3476), .B(n3475), .ZN(n3614) );
  AND2_X1 U3457 ( .A1(n3576), .A2(n3862), .ZN(n3595) );
  BUF_X1 U3458 ( .A(n3402), .Z(n2953) );
  AND2_X1 U34590 ( .A1(n4132), .A2(n3080), .ZN(n4268) );
  NAND2_X1 U34600 ( .A1(n4895), .A2(n4894), .ZN(n4893) );
  INV_X2 U34610 ( .A(n4620), .ZN(n4121) );
  INV_X1 U34620 ( .A(n4638), .ZN(n2945) );
  CLKBUF_X2 U34630 ( .A(n3327), .Z(n2970) );
  CLKBUF_X2 U34640 ( .A(n3199), .Z(n3978) );
  INV_X2 U34650 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3225) );
  OR2_X1 U3466 ( .A1(n5682), .A2(n6520), .ZN(n4293) );
  OAI21_X1 U3467 ( .B1(n5252), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n3961), 
        .ZN(n3962) );
  XNOR2_X1 U34680 ( .A(n5690), .B(n5691), .ZN(n5826) );
  OR2_X1 U34690 ( .A1(n5745), .A2(n5744), .ZN(n5747) );
  AOI211_X1 U34700 ( .C1(n5764), .C2(n5336), .A(n4304), .B(n4303), .ZN(n4305)
         );
  OAI21_X1 U34710 ( .B1(n5743), .B2(n5744), .A(n5746), .ZN(n5731) );
  NOR2_X1 U34720 ( .A1(n3738), .A2(n3737), .ZN(n3739) );
  AOI21_X1 U34730 ( .B1(n5808), .B2(n5906), .A(n5769), .ZN(n5758) );
  NOR2_X1 U34740 ( .A1(n4295), .A2(n3960), .ZN(n4102) );
  AND2_X1 U3475 ( .A1(n5358), .A2(n4301), .ZN(n5197) );
  NAND2_X1 U3476 ( .A1(n3090), .A2(n3089), .ZN(n4295) );
  OR2_X1 U3477 ( .A1(n5594), .A2(n5593), .ZN(n6321) );
  NOR2_X1 U3478 ( .A1(n5194), .A2(n3067), .ZN(n5324) );
  OAI22_X1 U3479 ( .A1(n5602), .A2(n3712), .B1(n3711), .B2(n5608), .ZN(n3729)
         );
  AOI21_X1 U3480 ( .B1(n5800), .B2(n3015), .A(n3014), .ZN(n5767) );
  XNOR2_X1 U3481 ( .A(n5608), .B(n3711), .ZN(n5602) );
  NOR2_X1 U3482 ( .A1(n3002), .A2(n2997), .ZN(n2996) );
  OAI21_X1 U3483 ( .B1(n3001), .B2(n3000), .A(n2998), .ZN(n2997) );
  NAND2_X1 U3484 ( .A1(n4891), .A2(n5045), .ZN(n5133) );
  NAND2_X1 U3485 ( .A1(n5369), .A2(n5215), .ZN(n5333) );
  OR2_X1 U3486 ( .A1(n5846), .A2(n4275), .ZN(n5835) );
  OR2_X1 U3487 ( .A1(n2977), .A2(n2972), .ZN(n3091) );
  NAND2_X1 U3488 ( .A1(n2972), .A2(n2994), .ZN(n3089) );
  OR2_X1 U3489 ( .A1(n4311), .A2(n4289), .ZN(n5838) );
  OR2_X1 U3490 ( .A1(n5881), .A2(n6784), .ZN(n5873) );
  AND3_X1 U3491 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .A3(
        n5460), .ZN(n5430) );
  NAND2_X1 U3492 ( .A1(n3064), .A2(n3061), .ZN(n5045) );
  OR4_X1 U3493 ( .A1(n5126), .A2(n5125), .A3(n5124), .A4(n5123), .ZN(n6282) );
  NAND2_X1 U3494 ( .A1(n5264), .A2(n5263), .ZN(n5574) );
  OR2_X1 U3495 ( .A1(n6333), .A2(n5211), .ZN(n6319) );
  NAND2_X1 U3496 ( .A1(n3476), .A2(n3401), .ZN(n3492) );
  INV_X1 U3497 ( .A(n5228), .ZN(n5226) );
  OR2_X1 U3498 ( .A1(n3463), .A2(n2987), .ZN(n3476) );
  AND2_X1 U3499 ( .A1(n5958), .A2(n4517), .ZN(n6570) );
  NAND2_X2 U3500 ( .A1(n5155), .A2(n5154), .ZN(n6409) );
  INV_X1 U3501 ( .A(n3408), .ZN(n3402) );
  AND2_X1 U3502 ( .A1(n4268), .A2(n4267), .ZN(n5938) );
  NAND2_X1 U3503 ( .A1(n4268), .A2(n4262), .ZN(n5923) );
  NAND2_X1 U3504 ( .A1(n3416), .A2(n3417), .ZN(n4577) );
  NAND2_X1 U3505 ( .A1(n5150), .A2(n5149), .ZN(n6695) );
  NAND2_X1 U3506 ( .A1(n3315), .A2(n3314), .ZN(n3415) );
  OR3_X1 U3507 ( .A1(n4432), .A2(n4431), .A3(n4430), .ZN(n4561) );
  OR2_X1 U3508 ( .A1(n4714), .A2(n4457), .ZN(n5150) );
  NAND2_X1 U3509 ( .A1(n3081), .A2(n3080), .ZN(n4714) );
  CLKBUF_X1 U3510 ( .A(n4545), .Z(n6218) );
  AND2_X1 U3511 ( .A1(n3323), .A2(n2956), .ZN(n3324) );
  NAND2_X1 U3512 ( .A1(n3349), .A2(n3348), .ZN(n4610) );
  OR2_X1 U3513 ( .A1(n4587), .A2(n2983), .ZN(n4840) );
  OR2_X1 U3514 ( .A1(n3056), .A2(n2993), .ZN(n3055) );
  OR2_X1 U3515 ( .A1(n5047), .A2(n5135), .ZN(n3056) );
  CLKBUF_X1 U3516 ( .A(n3404), .Z(n5174) );
  OR2_X1 U3517 ( .A1(n3496), .A2(n3245), .ZN(n3532) );
  NAND2_X1 U3518 ( .A1(n4638), .A2(n4620), .ZN(n4158) );
  CLKBUF_X1 U3519 ( .A(n2950), .Z(n3245) );
  OR2_X1 U3520 ( .A1(n3287), .A2(n3286), .ZN(n3480) );
  INV_X1 U3521 ( .A(n4209), .ZN(n2947) );
  CLKBUF_X1 U3522 ( .A(n2948), .Z(n3215) );
  AND2_X1 U3523 ( .A1(n3136), .A2(n3135), .ZN(n3143) );
  AND4_X1 U3524 ( .A1(n3148), .A2(n3147), .A3(n3146), .A4(n3145), .ZN(n3153)
         );
  AND4_X1 U3525 ( .A1(n3117), .A2(n3116), .A3(n3115), .A4(n3114), .ZN(n3123)
         );
  AND4_X1 U3526 ( .A1(n3203), .A2(n3202), .A3(n3201), .A4(n3200), .ZN(n3204)
         );
  AND4_X1 U3527 ( .A1(n3121), .A2(n3120), .A3(n3119), .A4(n3118), .ZN(n3122)
         );
  AND4_X1 U3528 ( .A1(n3105), .A2(n3104), .A3(n3103), .A4(n3102), .ZN(n3113)
         );
  AND4_X1 U3529 ( .A1(n3197), .A2(n3196), .A3(n3195), .A4(n3194), .ZN(n3205)
         );
  AND4_X1 U3530 ( .A1(n3111), .A2(n3110), .A3(n3109), .A4(n3108), .ZN(n3112)
         );
  AND4_X1 U3531 ( .A1(n3162), .A2(n3161), .A3(n3160), .A4(n3159), .ZN(n3163)
         );
  BUF_X2 U3532 ( .A(n4069), .Z(n3983) );
  AND3_X1 U3533 ( .A1(n3134), .A2(n3133), .A3(n3132), .ZN(n3136) );
  AND2_X2 U3534 ( .A1(n4440), .A2(n4547), .ZN(n3154) );
  AND2_X2 U3535 ( .A1(n3106), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3107)
         );
  AND2_X2 U3536 ( .A1(n4537), .A2(n4547), .ZN(n3333) );
  AND2_X2 U3537 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4548) );
  AND2_X2 U3539 ( .A1(n5603), .A2(n5604), .ZN(n5165) );
  AND2_X2 U3540 ( .A1(n3249), .A2(n4620), .ZN(n4209) );
  AND2_X1 U3541 ( .A1(n4258), .A2(n3236), .ZN(n4256) );
  NAND2_X1 U3542 ( .A1(n4268), .A2(n5270), .ZN(n5921) );
  INV_X1 U3543 ( .A(n4158), .ZN(n5439) );
  NAND2_X1 U3544 ( .A1(n3325), .A2(n3324), .ZN(n2954) );
  AND2_X1 U3545 ( .A1(n3113), .A2(n3112), .ZN(n2948) );
  INV_X1 U3546 ( .A(n2950), .ZN(n3209) );
  INV_X1 U3547 ( .A(n3210), .ZN(n2949) );
  AND2_X2 U3548 ( .A1(n2967), .A2(n4121), .ZN(n3404) );
  NAND3_X2 U3549 ( .A1(n3257), .A2(n3256), .A3(n3255), .ZN(n3273) );
  NOR2_X2 U3550 ( .A1(n2951), .A2(n2952), .ZN(n2950) );
  NAND4_X1 U3551 ( .A1(n3127), .A2(n3124), .A3(n3125), .A4(n3126), .ZN(n2951)
         );
  NAND4_X1 U3552 ( .A1(n3128), .A2(n3130), .A3(n3129), .A4(n3131), .ZN(n2952)
         );
  NAND2_X1 U3553 ( .A1(n3325), .A2(n3324), .ZN(n4530) );
  NOR2_X2 U3554 ( .A1(n4893), .A2(n3055), .ZN(n5514) );
  NOR2_X2 U3555 ( .A1(n5425), .A2(n2985), .ZN(n4312) );
  CLKBUF_X1 U3556 ( .A(n6476), .Z(n2955) );
  INV_X1 U3558 ( .A(n2963), .ZN(n2957) );
  BUF_X1 U3559 ( .A(n4332), .Z(n2958) );
  BUF_X1 U3560 ( .A(n3232), .Z(n2959) );
  NAND2_X1 U3561 ( .A1(n2948), .A2(n3237), .ZN(n3211) );
  NAND2_X1 U3562 ( .A1(n4258), .A2(n2960), .ZN(n4134) );
  AND2_X1 U3563 ( .A1(n3236), .A2(n4726), .ZN(n2960) );
  NAND2_X1 U3564 ( .A1(n3234), .A2(n4121), .ZN(n4717) );
  NAND2_X1 U3565 ( .A1(n3246), .A2(n4638), .ZN(n3228) );
  NAND2_X1 U3566 ( .A1(n3210), .A2(n3167), .ZN(n3581) );
  AND2_X1 U3568 ( .A1(n3181), .A2(n3180), .ZN(n2962) );
  AND2_X1 U3569 ( .A1(n3181), .A2(n3180), .ZN(n3231) );
  INV_X1 U3570 ( .A(n3449), .ZN(n6502) );
  AND2_X1 U3571 ( .A1(n3318), .A2(n3243), .ZN(n2964) );
  AND2_X1 U3572 ( .A1(n2966), .A2(STATE2_REG_0__SCAN_IN), .ZN(n2965) );
  OAI211_X1 U3573 ( .C1(n4396), .C2(n3238), .A(n4136), .B(n4134), .ZN(n2966)
         );
  NAND2_X1 U3574 ( .A1(n3318), .A2(n3243), .ZN(n3316) );
  AND2_X4 U3575 ( .A1(n3225), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4441)
         );
  AND2_X4 U3577 ( .A1(n3107), .A2(n4565), .ZN(n3328) );
  AND2_X1 U3578 ( .A1(n3235), .A2(n4620), .ZN(n3399) );
  NAND4_X1 U3579 ( .A1(n3207), .A2(n3206), .A3(n3205), .A4(n3204), .ZN(n2967)
         );
  AND2_X1 U3581 ( .A1(n3107), .A2(n4537), .ZN(n2968) );
  AND2_X1 U3582 ( .A1(n3107), .A2(n4537), .ZN(n2969) );
  AND2_X2 U3583 ( .A1(n3100), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4440)
         );
  NAND2_X2 U3584 ( .A1(n3272), .A2(n3273), .ZN(n3317) );
  OAI21_X1 U3585 ( .B1(n4434), .B2(STATE2_REG_0__SCAN_IN), .A(n3270), .ZN(
        n3271) );
  AND2_X2 U3586 ( .A1(n4440), .A2(n4548), .ZN(n4077) );
  INV_X1 U3587 ( .A(n4353), .ZN(n3049) );
  INV_X1 U3588 ( .A(n3340), .ZN(n3418) );
  NOR2_X2 U3589 ( .A1(n4631), .A2(n6768), .ZN(n3726) );
  NAND2_X1 U3590 ( .A1(n3550), .A2(n3549), .ZN(n4111) );
  NAND2_X1 U3591 ( .A1(n4044), .A2(n3068), .ZN(n3067) );
  INV_X1 U3592 ( .A(n5326), .ZN(n3068) );
  INV_X1 U3593 ( .A(n4044), .ZN(n3066) );
  AND2_X1 U3594 ( .A1(n5443), .A2(n5438), .ZN(n4208) );
  OR2_X1 U3595 ( .A1(n4131), .A2(n4432), .ZN(n4132) );
  OR2_X1 U3596 ( .A1(n4133), .A2(n3559), .ZN(n5121) );
  INV_X1 U3597 ( .A(n6695), .ZN(n5155) );
  NAND2_X1 U3598 ( .A1(n5232), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n3000) );
  NOR2_X1 U3599 ( .A1(n5254), .A2(n4291), .ZN(n3001) );
  NAND2_X1 U3600 ( .A1(n3524), .A2(n3523), .ZN(n3537) );
  XNOR2_X1 U3601 ( .A(n3525), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3534)
         );
  NAND2_X1 U3602 ( .A1(n3402), .A2(n3046), .ZN(n3463) );
  OR2_X1 U3603 ( .A1(n3384), .A2(n3383), .ZN(n3464) );
  NAND4_X1 U3604 ( .A1(n3247), .A2(n3256), .A3(n3223), .A4(n3558), .ZN(n3224)
         );
  AOI22_X1 U3605 ( .A1(n4123), .A2(n3209), .B1(n3215), .B2(n3218), .ZN(n3223)
         );
  NAND2_X1 U3606 ( .A1(n3211), .A2(n2950), .ZN(n3219) );
  AOI22_X1 U3607 ( .A1(n3292), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3168), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3105) );
  NAND2_X1 U3608 ( .A1(n3074), .A2(n3007), .ZN(n3006) );
  AND2_X1 U3609 ( .A1(n3075), .A2(n3530), .ZN(n3074) );
  NAND2_X1 U3610 ( .A1(n3008), .A2(n3519), .ZN(n3007) );
  INV_X1 U3611 ( .A(n3004), .ZN(n3003) );
  INV_X1 U3612 ( .A(n3541), .ZN(n3011) );
  AND2_X1 U3613 ( .A1(n3503), .A2(n3514), .ZN(n4108) );
  NAND2_X1 U3614 ( .A1(n4239), .A2(n4150), .ZN(n4152) );
  NOR2_X1 U3615 ( .A1(n5216), .A2(n3022), .ZN(n3021) );
  INV_X1 U3616 ( .A(n4095), .ZN(n4066) );
  NAND2_X1 U3617 ( .A1(n3821), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3823)
         );
  INV_X1 U3618 ( .A(n3877), .ZN(n3821) );
  NOR2_X1 U3619 ( .A1(n5103), .A2(n5129), .ZN(n4095) );
  OAI211_X1 U3620 ( .C1(n2953), .C2(n2987), .A(n3045), .B(n3044), .ZN(n3609)
         );
  OR2_X1 U3621 ( .A1(n3046), .A2(n2987), .ZN(n3045) );
  NAND2_X1 U3622 ( .A1(n2953), .A2(n2974), .ZN(n3044) );
  NOR2_X1 U3623 ( .A1(n3053), .A2(n5240), .ZN(n3052) );
  INV_X1 U3624 ( .A(n5205), .ZN(n3053) );
  AND2_X1 U3625 ( .A1(n5469), .A2(n4207), .ZN(n5438) );
  INV_X1 U3626 ( .A(n4231), .ZN(n4225) );
  INV_X1 U3627 ( .A(n4236), .ZN(n4224) );
  NAND2_X1 U3628 ( .A1(n4209), .A2(n4145), .ZN(n4231) );
  OR2_X1 U3629 ( .A1(n3299), .A2(n3298), .ZN(n3439) );
  XNOR2_X1 U3630 ( .A(n3343), .B(n3342), .ZN(n3414) );
  AOI21_X1 U3631 ( .B1(n3214), .B2(n4638), .A(n2949), .ZN(n3180) );
  NAND2_X1 U3632 ( .A1(n4545), .A2(n5129), .ZN(n3036) );
  OAI21_X1 U3633 ( .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n4652), .ZN(n6022) );
  AND2_X1 U3634 ( .A1(n4571), .A2(n5129), .ZN(n5060) );
  NAND2_X1 U3635 ( .A1(n6283), .A2(n4570), .ZN(n4571) );
  INV_X1 U3636 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5112) );
  XNOR2_X1 U3637 ( .A(n2954), .B(n4610), .ZN(n4545) );
  NAND2_X1 U3638 ( .A1(n4459), .A2(n4620), .ZN(n4723) );
  INV_X2 U3639 ( .A(n4092), .ZN(n5280) );
  AND2_X1 U3640 ( .A1(n6768), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5279) );
  OR2_X1 U3641 ( .A1(n4047), .A2(n4046), .ZN(n5157) );
  NAND2_X1 U3642 ( .A1(n3965), .A2(n3021), .ZN(n4045) );
  NAND2_X1 U3643 ( .A1(n3035), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4018)
         );
  NOR2_X1 U3644 ( .A1(n3964), .A2(n3963), .ZN(n3035) );
  NAND2_X1 U3645 ( .A1(n3907), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3964)
         );
  INV_X1 U3646 ( .A(n4322), .ZN(n3936) );
  OR2_X1 U3647 ( .A1(n3845), .A2(n6841), .ZN(n3906) );
  AND2_X1 U3648 ( .A1(n3688), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3689)
         );
  AND2_X1 U3649 ( .A1(n3694), .A2(n3693), .ZN(n5611) );
  INV_X1 U3650 ( .A(n5134), .ZN(n3629) );
  INV_X1 U3651 ( .A(n5133), .ZN(n3630) );
  NAND2_X1 U3652 ( .A1(n3612), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3632)
         );
  INV_X1 U3653 ( .A(n4792), .ZN(n3605) );
  OR3_X1 U3654 ( .A1(n3017), .A2(n5808), .A3(n5730), .ZN(n5746) );
  OAI211_X1 U3655 ( .C1(n3448), .C2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n3447), 
        .B(n6503), .ZN(n3451) );
  NAND3_X1 U3656 ( .A1(n3415), .A2(n3414), .A3(n3057), .ZN(n3408) );
  AND2_X1 U3657 ( .A1(n4862), .A2(n6588), .ZN(n4864) );
  INV_X1 U3658 ( .A(n6099), .ZN(n5986) );
  AND2_X1 U3659 ( .A1(n6213), .A2(n6216), .ZN(n6029) );
  AND2_X1 U3660 ( .A1(n4653), .A2(n6631), .ZN(n4654) );
  OR2_X1 U3661 ( .A1(n5975), .A2(n4580), .ZN(n4905) );
  AND2_X1 U3662 ( .A1(n5972), .A2(n5986), .ZN(n4869) );
  INV_X1 U3663 ( .A(n5060), .ZN(n4668) );
  NAND2_X1 U3664 ( .A1(n3553), .A2(n4111), .ZN(n3554) );
  NAND2_X1 U3665 ( .A1(n3551), .A2(n4111), .ZN(n3552) );
  AND2_X1 U3666 ( .A1(n5215), .A2(n3077), .ZN(n3076) );
  NOR2_X1 U3667 ( .A1(n5286), .A2(REIP_REG_29__SCAN_IN), .ZN(n3077) );
  AOI21_X1 U3668 ( .B1(n5329), .B2(REIP_REG_29__SCAN_IN), .A(n3025), .ZN(n3024) );
  OAI21_X1 U3669 ( .B1(n6327), .B2(n5575), .A(n3026), .ZN(n3025) );
  NAND2_X1 U3670 ( .A1(n6394), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n3026)
         );
  AND2_X1 U3671 ( .A1(n6409), .A2(n5158), .ZN(n6346) );
  NOR2_X1 U3672 ( .A1(n5678), .A2(n5301), .ZN(n5158) );
  AND2_X1 U3673 ( .A1(n5549), .A2(n5164), .ZN(n6399) );
  NOR2_X1 U3674 ( .A1(n3033), .A2(n5301), .ZN(n3032) );
  XNOR2_X1 U3675 ( .A(n3034), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5678)
         );
  NOR2_X1 U3676 ( .A1(n5157), .A2(n5156), .ZN(n3034) );
  OR2_X1 U3677 ( .A1(n5646), .A2(n5816), .ZN(n3957) );
  OR2_X1 U3678 ( .A1(n5652), .A2(n5816), .ZN(n4343) );
  NAND2_X1 U3679 ( .A1(n6298), .A2(n3731), .ZN(n5762) );
  OR2_X1 U3680 ( .A1(n4714), .A2(n5121), .ZN(n6298) );
  OR2_X1 U3681 ( .A1(n4312), .A2(n4354), .ZN(n5583) );
  OR2_X1 U3682 ( .A1(n6692), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6524) );
  INV_X1 U3683 ( .A(n6520), .ZN(n6579) );
  NAND2_X1 U3684 ( .A1(n4268), .A2(n4139), .ZN(n6520) );
  AND2_X1 U3685 ( .A1(n5128), .A2(n4245), .ZN(n4246) );
  INV_X1 U3686 ( .A(n5055), .ZN(n5972) );
  CLKBUF_X1 U3687 ( .A(n4577), .Z(n5975) );
  INV_X1 U3688 ( .A(n4858), .ZN(n5976) );
  NAND2_X1 U3689 ( .A1(n3249), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3496) );
  NAND2_X1 U3690 ( .A1(n3208), .A2(n3234), .ZN(n3247) );
  AND2_X1 U3691 ( .A1(n3214), .A2(n3249), .ZN(n4123) );
  INV_X1 U3692 ( .A(n3512), .ZN(n3008) );
  NAND2_X1 U3693 ( .A1(n3519), .A2(n2984), .ZN(n3075) );
  AND2_X1 U3694 ( .A1(n3523), .A2(n3516), .ZN(n3521) );
  NOR2_X1 U3695 ( .A1(n3048), .A2(n3047), .ZN(n3046) );
  INV_X1 U3696 ( .A(n3455), .ZN(n3048) );
  INV_X1 U3697 ( .A(n3403), .ZN(n3047) );
  OR2_X1 U3698 ( .A1(n3372), .A2(n3371), .ZN(n3465) );
  OAI211_X1 U3700 ( .C1(n3309), .C2(n3351), .A(n3308), .B(n3307), .ZN(n3422)
         );
  OR2_X1 U3701 ( .A1(n3339), .A2(n3338), .ZN(n3340) );
  OR2_X1 U3702 ( .A1(n3214), .A2(n3209), .ZN(n3213) );
  OR2_X1 U3703 ( .A1(n3361), .A2(n3360), .ZN(n3409) );
  AOI22_X1 U3704 ( .A1(n3258), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3104) );
  AOI22_X1 U3705 ( .A1(n3183), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3117) );
  OR2_X1 U3706 ( .A1(n3209), .A2(n5129), .ZN(n3350) );
  NAND2_X1 U3707 ( .A1(n3234), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3351) );
  NAND2_X1 U3708 ( .A1(n3540), .A2(n3399), .ZN(n3543) );
  INV_X1 U3709 ( .A(n3534), .ZN(n3536) );
  NAND2_X1 U3710 ( .A1(n3071), .A2(n3069), .ZN(n4336) );
  AND2_X1 U3711 ( .A1(n3889), .A2(n3070), .ZN(n3069) );
  INV_X1 U3712 ( .A(n3072), .ZN(n3070) );
  NOR2_X1 U3713 ( .A1(n3019), .A2(n3018), .ZN(n3844) );
  NOR2_X1 U3714 ( .A1(n3823), .A2(n5749), .ZN(n3020) );
  OR2_X1 U3715 ( .A1(n5510), .A2(n3073), .ZN(n3072) );
  INV_X1 U3716 ( .A(n5619), .ZN(n3073) );
  XNOR2_X1 U3717 ( .A(n3408), .B(n3403), .ZN(n3560) );
  NAND2_X1 U3718 ( .A1(n3575), .A2(n3726), .ZN(n3576) );
  INV_X1 U3719 ( .A(n3726), .ZN(n3882) );
  OR2_X1 U3720 ( .A1(n3756), .A2(n2994), .ZN(n3092) );
  AND2_X1 U3721 ( .A1(n4198), .A2(n5166), .ZN(n5469) );
  OR2_X1 U3722 ( .A1(n5502), .A2(n5612), .ZN(n3054) );
  NAND2_X1 U3723 ( .A1(n3013), .A2(n3460), .ZN(n3461) );
  OAI21_X1 U3724 ( .B1(n4236), .B2(INSTADDRPOINTER_REG_1__SCAN_IN), .A(n4145), 
        .ZN(n4144) );
  NAND2_X1 U3725 ( .A1(n4239), .A2(n4142), .ZN(n4143) );
  NOR2_X1 U3726 ( .A1(n3228), .A2(n3235), .ZN(n3229) );
  OR2_X1 U3727 ( .A1(n3581), .A2(n3556), .ZN(n5103) );
  AND2_X2 U3728 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4537) );
  AND2_X1 U3729 ( .A1(n3345), .A2(n4604), .ZN(n4956) );
  INV_X1 U3730 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6101) );
  INV_X1 U3731 ( .A(n4868), .ZN(n4735) );
  INV_X1 U3732 ( .A(n3543), .ZN(n3551) );
  NAND2_X1 U3733 ( .A1(n3012), .A2(n3010), .ZN(n3009) );
  NAND2_X1 U3734 ( .A1(n2980), .A2(n3005), .ZN(n3012) );
  CLKBUF_X1 U3735 ( .A(n4396), .Z(n4457) );
  AND2_X1 U3736 ( .A1(n4113), .A2(n4112), .ZN(n4406) );
  NOR2_X1 U3737 ( .A1(n3906), .A2(n4340), .ZN(n3907) );
  AND2_X1 U3738 ( .A1(n4220), .A2(n4219), .ZN(n4313) );
  NOR2_X2 U3739 ( .A1(n4840), .A2(n4162), .ZN(n4895) );
  NAND2_X1 U3740 ( .A1(n4236), .A2(EBX_REG_2__SCAN_IN), .ZN(n4151) );
  NOR2_X1 U3741 ( .A1(n4133), .A2(n4717), .ZN(n4720) );
  NAND2_X1 U3742 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .ZN(n4496) );
  AND2_X1 U3743 ( .A1(n4495), .A2(n5159), .ZN(n6421) );
  OAI21_X1 U3744 ( .B1(n4714), .B2(n4494), .A(n6473), .ZN(n4495) );
  NOR2_X1 U3745 ( .A1(n4714), .A2(n4458), .ZN(n4459) );
  OR2_X1 U3746 ( .A1(n4457), .A2(READY_N), .ZN(n4458) );
  INV_X1 U3747 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5156) );
  NAND2_X1 U3748 ( .A1(n3965), .A2(n2978), .ZN(n4047) );
  OR2_X1 U3749 ( .A1(n5381), .A2(n5412), .ZN(n3935) );
  INV_X1 U3750 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4340) );
  NAND2_X1 U3751 ( .A1(n3844), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3845)
         );
  INV_X1 U3752 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6841) );
  INV_X1 U3753 ( .A(n3020), .ZN(n3826) );
  NAND2_X1 U3754 ( .A1(n3697), .A2(n3030), .ZN(n3877) );
  NOR2_X1 U3755 ( .A1(n2990), .A2(n3031), .ZN(n3030) );
  INV_X1 U3756 ( .A(n3696), .ZN(n3697) );
  NAND2_X1 U3757 ( .A1(n3697), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3876)
         );
  NAND2_X1 U3758 ( .A1(n5403), .A2(n3695), .ZN(n5608) );
  AND2_X1 U3759 ( .A1(PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n3658), .ZN(n3688)
         );
  NOR2_X1 U3760 ( .A1(n3632), .A2(n3631), .ZN(n3657) );
  AND3_X1 U3761 ( .A1(n3628), .A2(n3627), .A3(n3626), .ZN(n5134) );
  NOR2_X1 U3762 ( .A1(n3611), .A2(n3610), .ZN(n3612) );
  AND2_X1 U3763 ( .A1(n3615), .A2(n3062), .ZN(n3061) );
  NAND2_X1 U3764 ( .A1(n6483), .A2(n3063), .ZN(n3062) );
  NAND2_X1 U3765 ( .A1(n3029), .A2(n3027), .ZN(n3611) );
  NOR2_X1 U3766 ( .A1(n6783), .A2(n3028), .ZN(n3027) );
  NOR2_X1 U3767 ( .A1(n3568), .A2(n6783), .ZN(n3601) );
  INV_X1 U3768 ( .A(n3591), .ZN(n3569) );
  NAND2_X1 U3769 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3591) );
  XNOR2_X1 U3770 ( .A(n4244), .B(n4243), .ZN(n5277) );
  INV_X1 U3771 ( .A(n4241), .ZN(n4244) );
  INV_X1 U3772 ( .A(n5677), .ZN(n2999) );
  NOR3_X1 U3773 ( .A1(n5808), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n5244), 
        .ZN(n4101) );
  NAND2_X1 U3774 ( .A1(n5342), .A2(n3050), .ZN(n5228) );
  NOR2_X1 U3775 ( .A1(n3051), .A2(n5262), .ZN(n3050) );
  INV_X1 U3776 ( .A(n3052), .ZN(n3051) );
  AND2_X1 U3777 ( .A1(n4234), .A2(n4233), .ZN(n5205) );
  NAND2_X1 U3778 ( .A1(n5342), .A2(n5205), .ZN(n5241) );
  INV_X1 U3779 ( .A(n5690), .ZN(n5189) );
  AND2_X1 U3780 ( .A1(n5363), .A2(n5344), .ZN(n5342) );
  NOR2_X2 U3781 ( .A1(n5374), .A2(n5362), .ZN(n5363) );
  XNOR2_X1 U3782 ( .A(n5808), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5698)
         );
  NAND2_X1 U3783 ( .A1(n4312), .A2(n4313), .ZN(n5376) );
  AND2_X1 U3784 ( .A1(n5942), .A2(n4286), .ZN(n4347) );
  OR2_X1 U3785 ( .A1(n5964), .A2(n4285), .ZN(n4286) );
  OAI21_X1 U3786 ( .B1(n3758), .B2(n3757), .A(n5808), .ZN(n3043) );
  AND2_X1 U3787 ( .A1(n5165), .A2(n5438), .ZN(n5472) );
  INV_X1 U3788 ( .A(n5729), .ZN(n3014) );
  NOR2_X1 U3789 ( .A1(n5728), .A2(n3016), .ZN(n3015) );
  INV_X1 U3790 ( .A(n5798), .ZN(n3016) );
  AND2_X1 U3791 ( .A1(n4186), .A2(n4185), .ZN(n5604) );
  NAND2_X1 U3792 ( .A1(n5800), .A2(n5798), .ZN(n5789) );
  NAND2_X1 U3793 ( .A1(n5306), .A2(n5129), .ZN(n6692) );
  OR2_X1 U3794 ( .A1(n4893), .A2(n5047), .ZN(n5136) );
  OAI211_X1 U3795 ( .C1(n3042), .C2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n3038), 
        .B(n3037), .ZN(n6477) );
  INV_X1 U3796 ( .A(n3482), .ZN(n3039) );
  INV_X1 U3797 ( .A(n3462), .ZN(n3088) );
  INV_X1 U3798 ( .A(n3086), .ZN(n4989) );
  NAND2_X1 U3799 ( .A1(n4832), .A2(n3454), .ZN(n6485) );
  XNOR2_X1 U3800 ( .A(n3461), .B(n6546), .ZN(n6484) );
  CLKBUF_X1 U3801 ( .A(n4115), .Z(n4116) );
  INV_X1 U3802 ( .A(n4268), .ZN(n4276) );
  XNOR2_X1 U3803 ( .A(n3316), .B(n3317), .ZN(n4434) );
  AND2_X1 U3804 ( .A1(n2962), .A2(n4128), .ZN(n4407) );
  INV_X1 U3805 ( .A(n5270), .ZN(n4494) );
  INV_X1 U3806 ( .A(n4435), .ZN(n6400) );
  CLKBUF_X1 U3807 ( .A(n4537), .Z(n4538) );
  CLKBUF_X1 U3808 ( .A(n4136), .Z(n4137) );
  AND2_X1 U3809 ( .A1(n4947), .A2(n5055), .ZN(n5987) );
  NOR2_X1 U3810 ( .A1(n4736), .A2(n4735), .ZN(n6059) );
  AND3_X1 U3811 ( .A1(n5116), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6062) );
  AND2_X1 U3812 ( .A1(n4732), .A2(n6203), .ZN(n4738) );
  AND2_X1 U3813 ( .A1(n5056), .A2(n5055), .ZN(n6150) );
  AND2_X1 U3814 ( .A1(n4579), .A2(n5975), .ZN(n5056) );
  OR2_X1 U3815 ( .A1(n4534), .A2(n6400), .ZN(n4899) );
  AND2_X1 U3816 ( .A1(n5060), .A2(n5059), .ZN(n6213) );
  AND2_X1 U3817 ( .A1(n5060), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4642) );
  NOR2_X1 U3818 ( .A1(n4905), .A2(n4735), .ZN(n6202) );
  INV_X1 U3819 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6103) );
  AND2_X1 U3820 ( .A1(n5301), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3555) );
  INV_X1 U3821 ( .A(n4496), .ZN(n4573) );
  OR2_X1 U3822 ( .A1(n4116), .A2(n3411), .ZN(n5128) );
  INV_X1 U3823 ( .A(n6436), .ZN(n6693) );
  NAND2_X1 U3824 ( .A1(n4401), .A2(n3080), .ZN(n5149) );
  AND2_X1 U3825 ( .A1(n3079), .A2(n3078), .ZN(n5319) );
  INV_X1 U3826 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6783) );
  AND2_X1 U3827 ( .A1(n6409), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6394) );
  AND2_X1 U3828 ( .A1(n6371), .A2(n5550), .ZN(n6404) );
  INV_X1 U3829 ( .A(n6394), .ZN(n6376) );
  INV_X1 U3830 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6794) );
  INV_X1 U3831 ( .A(n5624), .ZN(n5628) );
  INV_X1 U3832 ( .A(n5626), .ZN(n5627) );
  NAND2_X1 U3833 ( .A1(n4421), .A2(n4420), .ZN(n5626) );
  AND2_X1 U3834 ( .A1(n6420), .A2(n4726), .ZN(n6410) );
  AND2_X1 U3835 ( .A1(n6420), .A2(n4725), .ZN(n6417) );
  INV_X1 U3836 ( .A(n6420), .ZN(n6412) );
  OR2_X1 U3837 ( .A1(n6410), .A2(n6413), .ZN(n6416) );
  INV_X1 U3838 ( .A(n6416), .ZN(n5670) );
  INV_X2 U3839 ( .A(n6417), .ZN(n5675) );
  INV_X1 U3841 ( .A(n6693), .ZN(n6449) );
  CLKBUF_X1 U3842 ( .A(n6471), .Z(n6464) );
  OR2_X1 U3843 ( .A1(n4714), .A2(n5128), .ZN(n6473) );
  NOR2_X1 U3844 ( .A1(n6467), .A2(n4459), .ZN(n6471) );
  INV_X1 U3845 ( .A(n4723), .ZN(n6470) );
  XNOR2_X1 U3846 ( .A(n5324), .B(n5281), .ZN(n5633) );
  NAND2_X1 U3847 ( .A1(n3965), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3966)
         );
  OAI21_X1 U3848 ( .B1(n5345), .B2(n5195), .A(n5347), .ZN(n5696) );
  INV_X1 U3849 ( .A(n3035), .ZN(n4016) );
  NAND2_X1 U3850 ( .A1(n3065), .A2(n3605), .ZN(n4889) );
  OR2_X1 U3851 ( .A1(n5425), .A2(n2981), .ZN(n5418) );
  INV_X1 U3852 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6838) );
  NAND2_X1 U3853 ( .A1(n5742), .A2(n5741), .ZN(n5748) );
  NOR2_X1 U3854 ( .A1(n5740), .A2(n5739), .ZN(n5741) );
  NAND2_X2 U3855 ( .A1(n3437), .A2(n3436), .ZN(n6099) );
  NAND2_X1 U3856 ( .A1(n3435), .A2(n3434), .ZN(n3436) );
  BUF_X1 U3857 ( .A(n3431), .Z(n3437) );
  CLKBUF_X1 U3858 ( .A(n4434), .Z(n4435) );
  NAND2_X1 U3859 ( .A1(n3326), .A2(n2954), .ZN(n4534) );
  INV_X1 U3860 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5116) );
  NAND2_X1 U3861 ( .A1(n3417), .A2(n4580), .ZN(n3058) );
  INV_X1 U3862 ( .A(n6218), .ZN(n6206) );
  NAND2_X1 U3863 ( .A1(n4572), .A2(n4668), .ZN(n6584) );
  AND2_X1 U3864 ( .A1(n4407), .A2(n4620), .ZN(n5270) );
  INV_X1 U3865 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5275) );
  INV_X1 U3866 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3100) );
  INV_X1 U3867 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5300) );
  NOR2_X1 U3868 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n5306) );
  OAI21_X1 U3869 ( .B1(n4867), .B2(n4864), .A(n4863), .ZN(n6591) );
  NAND2_X1 U3870 ( .A1(n4947), .A2(n4868), .ZN(n6595) );
  INV_X1 U3871 ( .A(n6591), .ZN(n4888) );
  INV_X1 U3872 ( .A(n5039), .ZN(n4646) );
  INV_X1 U3873 ( .A(n6143), .ZN(n4765) );
  AOI22_X1 U3874 ( .A1(n6158), .A2(n6155), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6156), .ZN(n6201) );
  INV_X1 U3875 ( .A(n6641), .ZN(n5094) );
  INV_X1 U3876 ( .A(n6226), .ZN(n6071) );
  INV_X1 U3877 ( .A(n6234), .ZN(n6075) );
  INV_X1 U3878 ( .A(n6249), .ZN(n6610) );
  INV_X1 U3879 ( .A(n6256), .ZN(n6617) );
  INV_X1 U3880 ( .A(n6263), .ZN(n6624) );
  INV_X1 U3881 ( .A(n6272), .ZN(n6632) );
  OAI21_X1 U3882 ( .B1(n4657), .B2(n4656), .A(n4655), .ZN(n6638) );
  NAND2_X1 U3883 ( .A1(n5056), .A2(n4869), .ZN(n6634) );
  INV_X1 U3884 ( .A(n4680), .ZN(n4707) );
  AND2_X1 U3885 ( .A1(n5795), .A2(DATAI_17_), .ZN(n6170) );
  AND2_X1 U3886 ( .A1(n5795), .A2(DATAI_18_), .ZN(n6175) );
  AND2_X1 U3887 ( .A1(n5795), .A2(DATAI_19_), .ZN(n6179) );
  AND2_X1 U3888 ( .A1(n5795), .A2(DATAI_21_), .ZN(n6187) );
  AND2_X1 U3889 ( .A1(n5795), .A2(DATAI_22_), .ZN(n6191) );
  AND2_X1 U3890 ( .A1(n5795), .A2(DATAI_23_), .ZN(n6198) );
  INV_X1 U3891 ( .A(n6599), .ZN(n6220) );
  INV_X1 U3892 ( .A(n6170), .ZN(n6233) );
  INV_X1 U3893 ( .A(n6114), .ZN(n6228) );
  INV_X1 U3894 ( .A(n6179), .ZN(n6604) );
  INV_X1 U3895 ( .A(n6606), .ZN(n6244) );
  INV_X1 U3896 ( .A(n6183), .ZN(n6611) );
  INV_X1 U3897 ( .A(n6187), .ZN(n6618) );
  INV_X1 U3898 ( .A(n6620), .ZN(n6258) );
  INV_X1 U3899 ( .A(n6191), .ZN(n6625) );
  INV_X1 U3900 ( .A(n6627), .ZN(n6265) );
  NOR2_X2 U3901 ( .A1(n4905), .A2(n4904), .ZN(n6278) );
  INV_X1 U3902 ( .A(n6637), .ZN(n6274) );
  NAND2_X1 U3903 ( .A1(n5795), .A2(DATAI_24_), .ZN(n6602) );
  INV_X1 U3904 ( .A(n6162), .ZN(n6596) );
  AND2_X1 U3905 ( .A1(n5795), .A2(DATAI_16_), .ZN(n6165) );
  NOR2_X1 U3906 ( .A1(n4728), .A2(n4668), .ZN(n6114) );
  NOR2_X1 U3907 ( .A1(n4729), .A2(n4668), .ZN(n6119) );
  AND2_X1 U3908 ( .A1(n4642), .A2(n4638), .ZN(n6242) );
  NOR2_X1 U3909 ( .A1(n4790), .A2(n4668), .ZN(n6606) );
  AND2_X1 U3910 ( .A1(n5795), .A2(DATAI_20_), .ZN(n6183) );
  NOR2_X2 U3911 ( .A1(n4905), .A2(n4598), .ZN(n4983) );
  NOR2_X1 U3912 ( .A1(n6764), .A2(n4668), .ZN(n6620) );
  NOR2_X1 U3913 ( .A1(n6726), .A2(n4668), .ZN(n6627) );
  NOR2_X1 U3914 ( .A1(n5046), .A2(n4668), .ZN(n6637) );
  INV_X1 U3915 ( .A(n6202), .ZN(n6281) );
  OR2_X1 U3916 ( .A1(n4445), .A2(n6103), .ZN(n6283) );
  INV_X2 U3917 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6768) );
  NOR2_X1 U3918 ( .A1(n5151), .A2(n6297), .ZN(n4369) );
  INV_X1 U3919 ( .A(n6680), .ZN(n6677) );
  INV_X1 U3920 ( .A(STATE_REG_1__SCAN_IN), .ZN(n4378) );
  INV_X2 U3921 ( .A(n6702), .ZN(n6855) );
  AND2_X1 U3922 ( .A1(STATE_REG_1__SCAN_IN), .A2(n6710), .ZN(n6702) );
  INV_X1 U3923 ( .A(n3023), .ZN(n5327) );
  OAI211_X1 U3924 ( .C1(n5330), .C2(n5685), .A(n3079), .B(n3024), .ZN(n3023)
         );
  AND2_X1 U3925 ( .A1(n3957), .A2(n3956), .ZN(n3958) );
  INV_X1 U3926 ( .A(n4327), .ZN(n4328) );
  OAI21_X1 U3927 ( .B1(n5649), .B2(n5816), .A(n4326), .ZN(n4327) );
  AND2_X1 U3928 ( .A1(n4343), .A2(n4342), .ZN(n4344) );
  NAND2_X1 U3929 ( .A1(n3736), .A2(n3735), .ZN(n3737) );
  NAND2_X1 U3930 ( .A1(n4293), .A2(n2996), .ZN(U2987) );
  NOR2_X1 U3931 ( .A1(n5235), .A2(n4292), .ZN(n3002) );
  OAI211_X1 U3932 ( .C1(n5267), .C2(n5266), .A(n5265), .B(n3093), .ZN(n5268)
         );
  AND2_X1 U3933 ( .A1(n4356), .A2(n4355), .ZN(n4357) );
  AND2_X1 U3934 ( .A1(n3092), .A2(n5808), .ZN(n2972) );
  OAI211_X1 U3935 ( .C1(n3452), .C2(n6492), .A(n3450), .B(n3451), .ZN(n4830)
         );
  INV_X1 U3936 ( .A(n4209), .ZN(n4141) );
  AND2_X1 U3937 ( .A1(n3756), .A2(n3757), .ZN(n2973) );
  INV_X1 U3938 ( .A(n4445), .ZN(n3081) );
  AND2_X1 U3939 ( .A1(n3046), .A2(n2987), .ZN(n2974) );
  OR2_X1 U3940 ( .A1(n2981), .A2(n5417), .ZN(n2975) );
  AND2_X1 U3941 ( .A1(n3482), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n2976)
         );
  AND2_X1 U3942 ( .A1(n2973), .A2(n2995), .ZN(n2977) );
  NAND2_X1 U3943 ( .A1(n3020), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3019)
         );
  AND2_X1 U3944 ( .A1(n3021), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n2978)
         );
  BUF_X1 U3945 ( .A(n3137), .Z(n3183) );
  NAND2_X1 U3946 ( .A1(n5720), .A2(n3043), .ZN(n4306) );
  INV_X1 U3947 ( .A(n3399), .ZN(n3526) );
  NOR2_X1 U3948 ( .A1(n5511), .A2(n5510), .ZN(n5512) );
  AND2_X1 U3949 ( .A1(n4321), .A2(n3936), .ZN(n3953) );
  AND2_X1 U3950 ( .A1(n4296), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n2979)
         );
  AND2_X1 U3951 ( .A1(n3006), .A2(n3533), .ZN(n2980) );
  OR2_X1 U3952 ( .A1(n4213), .A2(n4212), .ZN(n2981) );
  AND2_X1 U3953 ( .A1(n3758), .A2(n3756), .ZN(n2982) );
  AOI21_X1 U3954 ( .B1(n3344), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3320), 
        .ZN(n3322) );
  NAND2_X1 U3955 ( .A1(n5767), .A2(n5768), .ZN(n3017) );
  INV_X1 U3956 ( .A(n6409), .ZN(n3033) );
  OR2_X1 U3957 ( .A1(n4837), .A2(n4588), .ZN(n2983) );
  AND3_X1 U3958 ( .A1(n3511), .A2(STATE2_REG_0__SCAN_IN), .A3(n4108), .ZN(
        n2984) );
  AOI21_X1 U3959 ( .B1(n3538), .B2(n3399), .A(n4112), .ZN(n3542) );
  INV_X1 U3960 ( .A(n3542), .ZN(n3005) );
  NOR2_X1 U3961 ( .A1(n5511), .A2(n3072), .ZN(n3890) );
  AND2_X1 U3962 ( .A1(n5342), .A2(n3052), .ZN(n4240) );
  INV_X1 U3963 ( .A(n3057), .ZN(n4580) );
  NAND2_X1 U3964 ( .A1(n3036), .A2(n3362), .ZN(n3057) );
  NAND2_X1 U3965 ( .A1(n3630), .A2(n3629), .ZN(n5511) );
  INV_X1 U3966 ( .A(n5511), .ZN(n3071) );
  OR2_X1 U3967 ( .A1(n2975), .A2(n3049), .ZN(n2985) );
  NAND2_X1 U3968 ( .A1(n5369), .A2(n3076), .ZN(n3079) );
  AND2_X2 U3969 ( .A1(n4548), .A2(n4537), .ZN(n3199) );
  OR2_X1 U3970 ( .A1(n3418), .A2(n3350), .ZN(n2986) );
  INV_X1 U3971 ( .A(n5412), .ZN(n3063) );
  INV_X1 U3972 ( .A(n4791), .ZN(n3065) );
  OR2_X1 U3973 ( .A1(n5623), .A2(n5502), .ZN(n5501) );
  NAND2_X1 U3974 ( .A1(n4830), .A2(n4831), .ZN(n4832) );
  AND2_X1 U3975 ( .A1(n3398), .A2(n3397), .ZN(n2987) );
  NAND2_X1 U3976 ( .A1(n3408), .A2(n3058), .ZN(n3567) );
  OR2_X1 U3977 ( .A1(n4296), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n2988)
         );
  NOR2_X1 U3978 ( .A1(n5425), .A2(n2975), .ZN(n2989) );
  NAND2_X1 U3979 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n2990) );
  NOR2_X1 U3980 ( .A1(n4893), .A2(n3056), .ZN(n2991) );
  XOR2_X1 U3981 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3632), .Z(n2992) );
  INV_X1 U3982 ( .A(n6644), .ZN(n3080) );
  INV_X1 U3983 ( .A(n3568), .ZN(n3029) );
  NAND2_X1 U3984 ( .A1(n4172), .A2(n4171), .ZN(n2993) );
  INV_X1 U3985 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n5129) );
  INV_X1 U3986 ( .A(n6691), .ZN(n6203) );
  NAND2_X1 U3987 ( .A1(n6768), .A2(n6103), .ZN(n6691) );
  INV_X1 U3988 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3031) );
  NAND3_X1 U3989 ( .A1(n4288), .A2(n5863), .A3(n4349), .ZN(n2994) );
  AND3_X1 U3990 ( .A1(n4350), .A2(n5845), .A3(n6838), .ZN(n2995) );
  INV_X1 U3991 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3018) );
  INV_X1 U3992 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5301) );
  INV_X1 U3993 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3022) );
  INV_X1 U3994 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3028) );
  NOR2_X2 U3995 ( .A1(n5958), .A2(n5938), .ZN(n5964) );
  OAI21_X1 U3996 ( .B1(n3006), .B2(n3005), .A(n3003), .ZN(n3010) );
  OAI21_X1 U3997 ( .B1(n3005), .B2(n3533), .A(n3011), .ZN(n3004) );
  NAND2_X1 U3998 ( .A1(n3009), .A2(n3552), .ZN(n3082) );
  NAND2_X1 U3999 ( .A1(n3604), .A2(n3399), .ZN(n3013) );
  NAND2_X2 U4000 ( .A1(n6485), .A2(n6484), .ZN(n6487) );
  INV_X1 U4001 ( .A(n3017), .ZN(n5769) );
  OAI21_X2 U4002 ( .B1(n4577), .B2(n3526), .A(n3420), .ZN(n3449) );
  NAND2_X2 U4003 ( .A1(n5678), .A2(n3032), .ZN(n5330) );
  NAND2_X1 U4004 ( .A1(n3472), .A2(n3086), .ZN(n3040) );
  NAND2_X1 U4005 ( .A1(n3085), .A2(n6487), .ZN(n3041) );
  NAND2_X1 U4006 ( .A1(n3042), .A2(n3482), .ZN(n3483) );
  NAND3_X1 U4007 ( .A1(n3041), .A2(n3040), .A3(n6477), .ZN(n6476) );
  NAND2_X1 U4008 ( .A1(n3042), .A2(n2976), .ZN(n3037) );
  NAND2_X1 U4009 ( .A1(n3039), .A2(n6536), .ZN(n3038) );
  NAND2_X1 U4010 ( .A1(n3614), .A2(n3399), .ZN(n3042) );
  OAI22_X2 U4011 ( .A1(n4306), .A2(n5712), .B1(n5808), .B2(n6838), .ZN(n5705)
         );
  NAND2_X1 U4012 ( .A1(n3402), .A2(n3403), .ZN(n3456) );
  AND2_X2 U4013 ( .A1(n4209), .A2(n5439), .ZN(n4239) );
  NAND2_X1 U4014 ( .A1(n3415), .A2(n3414), .ZN(n3417) );
  INV_X1 U4015 ( .A(n4890), .ZN(n3059) );
  NAND2_X1 U4016 ( .A1(n3059), .A2(n3605), .ZN(n3060) );
  NOR2_X2 U4017 ( .A1(n4791), .A2(n3060), .ZN(n4891) );
  NAND2_X1 U4018 ( .A1(n3614), .A2(n3726), .ZN(n3064) );
  INV_X1 U4019 ( .A(n5194), .ZN(n5358) );
  NOR2_X2 U4020 ( .A1(n4336), .A2(n4337), .ZN(n4321) );
  NOR2_X2 U4021 ( .A1(n6319), .A2(n5212), .ZN(n5460) );
  NAND2_X2 U4022 ( .A1(n5549), .A2(n5161), .ZN(n6333) );
  AND2_X2 U4023 ( .A1(n6409), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5549) );
  INV_X1 U4024 ( .A(n5329), .ZN(n3078) );
  AND2_X2 U4025 ( .A1(n5392), .A2(n5213), .ZN(n5369) );
  NAND2_X1 U4026 ( .A1(n3497), .A2(n4717), .ZN(n3528) );
  NAND2_X2 U4027 ( .A1(n3082), .A2(n3554), .ZN(n4445) );
  NAND2_X1 U4028 ( .A1(n3083), .A2(n2986), .ZN(n3343) );
  NAND3_X1 U4029 ( .A1(n3326), .A2(n4530), .A3(n5129), .ZN(n3083) );
  OAI211_X1 U4030 ( .C1(n3086), .C2(n6487), .A(n3472), .B(n3084), .ZN(n6475)
         );
  NAND2_X1 U4031 ( .A1(n4989), .A2(n3088), .ZN(n3084) );
  NOR2_X1 U4032 ( .A1(n3087), .A2(n3088), .ZN(n3085) );
  INV_X1 U4033 ( .A(n3472), .ZN(n3087) );
  NAND2_X1 U4034 ( .A1(n4987), .A2(n4989), .ZN(n4988) );
  NAND2_X1 U4035 ( .A1(n6487), .A2(n3462), .ZN(n4987) );
  NAND2_X1 U4036 ( .A1(n3758), .A2(n3091), .ZN(n3090) );
  NAND2_X1 U4037 ( .A1(n3758), .A2(n2973), .ZN(n5720) );
  INV_X1 U4038 ( .A(n4321), .ZN(n4338) );
  AOI21_X1 U4039 ( .B1(n4299), .B2(n5190), .A(n4298), .ZN(n4300) );
  NAND2_X1 U4040 ( .A1(n5189), .A2(n4294), .ZN(n4299) );
  NOR3_X2 U4041 ( .A1(n5333), .A2(n5286), .A3(n5285), .ZN(n5316) );
  INV_X1 U4042 ( .A(n3567), .ZN(n4579) );
  AOI22_X1 U4043 ( .A1(n3263), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3173), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3121) );
  OR2_X1 U4044 ( .A1(n5574), .A2(n5966), .ZN(n3093) );
  INV_X1 U4045 ( .A(n5630), .ZN(n5617) );
  INV_X1 U4046 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3525) );
  OR2_X1 U4047 ( .A1(n3242), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3094)
         );
  NOR2_X2 U4048 ( .A1(n4276), .A2(n4246), .ZN(n6541) );
  OAI21_X1 U4049 ( .B1(n3095), .B2(n4144), .A(n4143), .ZN(n4147) );
  INV_X1 U4050 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3545) );
  AND2_X1 U4051 ( .A1(n4209), .A2(n4142), .ZN(n3095) );
  INV_X1 U4052 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6710) );
  INV_X1 U4053 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6293) );
  INV_X1 U4054 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3631) );
  INV_X2 U4055 ( .A(n5816), .ZN(n5795) );
  INV_X1 U4056 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3515) );
  AND3_X1 U4057 ( .A1(n3151), .A2(n3150), .A3(n3149), .ZN(n3096) );
  OR3_X1 U4058 ( .A1(n6292), .A2(n6291), .A3(STATE2_REG_3__SCAN_IN), .ZN(n3097) );
  NOR2_X1 U4059 ( .A1(n6025), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3098)
         );
  INV_X1 U4060 ( .A(n5346), .ZN(n5195) );
  AND2_X1 U4061 ( .A1(n6207), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3502)
         );
  NOR2_X1 U4062 ( .A1(n3525), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3535)
         );
  INV_X1 U4063 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3099) );
  AOI21_X1 U4064 ( .B1(n3537), .B2(n3536), .A(n3535), .ZN(n3547) );
  AOI22_X1 U4065 ( .A1(n4027), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3119) );
  AND2_X1 U4066 ( .A1(n3227), .A2(n3226), .ZN(n3241) );
  AND2_X1 U4067 ( .A1(n3547), .A2(n6293), .ZN(n3544) );
  INV_X1 U4068 ( .A(n3480), .ZN(n3485) );
  OR2_X1 U4069 ( .A1(n3396), .A2(n3395), .ZN(n3478) );
  OR2_X1 U4070 ( .A1(n3269), .A2(n3268), .ZN(n3425) );
  NAND2_X1 U4071 ( .A1(n3544), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4112) );
  NOR2_X1 U4072 ( .A1(READY_N), .A2(n4406), .ZN(n4715) );
  INV_X1 U4073 ( .A(n5611), .ZN(n3695) );
  NAND2_X1 U4074 ( .A1(n2949), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4092) );
  NOR2_X1 U4075 ( .A1(n3400), .A2(n3526), .ZN(n3401) );
  OR2_X1 U4076 ( .A1(n6697), .A2(n4573), .ZN(n4570) );
  INV_X1 U4077 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3963) );
  INV_X1 U4078 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3825) );
  OR2_X1 U4079 ( .A1(n3885), .A2(n5611), .ZN(n5484) );
  INV_X1 U4080 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3610) );
  AND2_X1 U4081 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4349) );
  AND2_X1 U4082 ( .A1(n5808), .A2(n4330), .ZN(n4331) );
  AND2_X1 U4083 ( .A1(n5989), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6016)
         );
  AND2_X1 U4084 ( .A1(n5972), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4858) );
  AND2_X1 U4085 ( .A1(n6156), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6194)
         );
  AND2_X1 U4086 ( .A1(n4642), .A2(n4724), .ZN(n6272) );
  INV_X1 U4087 ( .A(STATE_REG_2__SCAN_IN), .ZN(n3216) );
  AND2_X1 U4088 ( .A1(n4407), .A2(n4397), .ZN(n4401) );
  NOR2_X1 U4089 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n5410) );
  INV_X1 U4090 ( .A(n5410), .ZN(n5412) );
  INV_X1 U4091 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5749) );
  INV_X1 U4092 ( .A(n3734), .ZN(n3735) );
  INV_X1 U4093 ( .A(n4240), .ZN(n5261) );
  INV_X1 U4094 ( .A(n5966), .ZN(n4314) );
  OR2_X1 U4095 ( .A1(n5897), .A2(n4272), .ZN(n5888) );
  AND2_X1 U4096 ( .A1(n4282), .A2(n4281), .ZN(n5942) );
  INV_X1 U4097 ( .A(n5938), .ZN(n6577) );
  INV_X1 U4098 ( .A(n4578), .ZN(n5055) );
  NAND2_X1 U4099 ( .A1(n4947), .A2(n4869), .ZN(n6589) );
  NOR2_X1 U4100 ( .A1(n5975), .A2(n3057), .ZN(n4734) );
  AOI21_X1 U4101 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4955), .A(n4668), .ZN(
        n4951) );
  NAND2_X1 U4102 ( .A1(n6150), .A2(n6099), .ZN(n6196) );
  INV_X1 U4103 ( .A(n6199), .ZN(n5096) );
  INV_X1 U4104 ( .A(n6242), .ZN(n6603) );
  NAND2_X1 U4105 ( .A1(n4666), .A2(n4665), .ZN(n4942) );
  OR2_X1 U4106 ( .A1(n5972), .A2(n6099), .ZN(n4904) );
  INV_X1 U4107 ( .A(n4902), .ZN(n6161) );
  AND2_X1 U4108 ( .A1(n4667), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6208)
         );
  AND2_X1 U4109 ( .A1(n5567), .A2(n5209), .ZN(n5383) );
  NAND2_X1 U4110 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n3689), .ZN(n3696)
         );
  INV_X1 U4111 ( .A(n6365), .ZN(n6378) );
  AND3_X1 U4112 ( .A1(n6524), .A2(n6647), .A3(n6288), .ZN(n5154) );
  NAND2_X1 U4113 ( .A1(n4419), .A2(n4209), .ZN(n4420) );
  AND2_X1 U4114 ( .A1(n6420), .A2(n4727), .ZN(n6413) );
  AOI21_X1 U4115 ( .B1(n4721), .B2(n4720), .A(n4719), .ZN(n4722) );
  NOR2_X1 U4116 ( .A1(n4496), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6436) );
  INV_X1 U4117 ( .A(n6473), .ZN(n6467) );
  OR2_X1 U4118 ( .A1(n5633), .A2(n5816), .ZN(n4099) );
  INV_X1 U4119 ( .A(n6298), .ZN(n6505) );
  AND2_X1 U4120 ( .A1(n5261), .A2(n5242), .ZN(n5576) );
  INV_X1 U4121 ( .A(n6524), .ZN(n6573) );
  AND2_X1 U4122 ( .A1(n5987), .A2(n6099), .ZN(n6019) );
  INV_X1 U4123 ( .A(n6595), .ZN(n6056) );
  NOR2_X1 U4124 ( .A1(n4579), .A2(n3575), .ZN(n4947) );
  OAI21_X1 U4125 ( .B1(n4867), .B2(n4866), .A(n4865), .ZN(n6592) );
  INV_X1 U4126 ( .A(n6589), .ZN(n5041) );
  OAI211_X1 U4127 ( .C1(n6203), .C2(n5000), .A(n4617), .B(n6161), .ZN(n4647)
         );
  NOR2_X1 U4128 ( .A1(n4736), .A2(n4904), .ZN(n6095) );
  NAND4_X1 U4129 ( .A1(n6064), .A2(n6213), .A3(n6063), .A4(n6211), .ZN(n6091)
         );
  OAI21_X1 U4130 ( .B1(n4742), .B2(n4741), .A(n4740), .ZN(n4766) );
  INV_X1 U4131 ( .A(n6196), .ZN(n6145) );
  AND2_X1 U4132 ( .A1(n6150), .A2(n5986), .ZN(n6199) );
  OAI22_X1 U4133 ( .A1(n5064), .A2(n5063), .B1(n6215), .B2(n6211), .ZN(n5098)
         );
  NOR2_X1 U4134 ( .A1(n4731), .A2(n4668), .ZN(n6599) );
  NOR2_X1 U4135 ( .A1(n4787), .A2(n4668), .ZN(n6613) );
  AND2_X1 U4136 ( .A1(n5972), .A2(n6099), .ZN(n4868) );
  INV_X1 U4137 ( .A(n6634), .ZN(n4710) );
  OAI21_X1 U4138 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6103), .A(n5060), 
        .ZN(n4902) );
  INV_X1 U4139 ( .A(n6602), .ZN(n6222) );
  INV_X1 U4140 ( .A(n6616), .ZN(n6253) );
  NAND4_X1 U4141 ( .A1(n6214), .A2(n6213), .A3(n6212), .A4(n6211), .ZN(n6270)
         );
  OAI211_X1 U4142 ( .C1(n6208), .C2(n6203), .A(n4597), .B(n6161), .ZN(n4822)
         );
  NOR2_X1 U4143 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6697) );
  AND3_X1 U4144 ( .A1(n4106), .A2(n6710), .A3(n4364), .ZN(n5159) );
  INV_X1 U4145 ( .A(n6653), .ZN(n6857) );
  INV_X1 U4146 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6297) );
  INV_X1 U4147 ( .A(n5277), .ZN(n5295) );
  NAND2_X1 U4148 ( .A1(n5626), .A2(n2949), .ZN(n5624) );
  INV_X1 U4149 ( .A(DATAI_7_), .ZN(n5046) );
  NAND2_X1 U4150 ( .A1(n4723), .A2(n4722), .ZN(n6420) );
  NAND2_X1 U4151 ( .A1(n6421), .A2(n2967), .ZN(n4856) );
  INV_X1 U4152 ( .A(n6421), .ZN(n6451) );
  INV_X1 U4153 ( .A(n6471), .ZN(n4493) );
  AND2_X1 U4154 ( .A1(n4099), .A2(n4098), .ZN(n4100) );
  OAI21_X1 U4155 ( .B1(n5594), .B2(n5468), .A(n5467), .ZN(n5754) );
  NAND2_X1 U4156 ( .A1(n4369), .A2(n6203), .ZN(n5816) );
  AND2_X1 U4157 ( .A1(n4317), .A2(n4316), .ZN(n4318) );
  INV_X1 U4158 ( .A(n6541), .ZN(n5966) );
  INV_X1 U4159 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6789) );
  INV_X1 U4160 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6207) );
  INV_X1 U4161 ( .A(n6019), .ZN(n4986) );
  AOI22_X1 U4162 ( .A1(n5991), .A2(n5988), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5989), .ZN(n6021) );
  NAND2_X1 U4163 ( .A1(n5987), .A2(n5986), .ZN(n6058) );
  AOI22_X1 U4164 ( .A1(n4616), .A2(n4613), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5000), .ZN(n4650) );
  INV_X1 U4165 ( .A(n6059), .ZN(n6098) );
  AOI22_X1 U4166 ( .A1(n4738), .A2(n4741), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6062), .ZN(n4769) );
  INV_X1 U4167 ( .A(n6613), .ZN(n6251) );
  AOI21_X1 U4168 ( .B1(n5062), .B2(n5063), .A(n5061), .ZN(n5101) );
  INV_X1 U4169 ( .A(n6119), .ZN(n6236) );
  NAND2_X1 U4170 ( .A1(n5056), .A2(n4868), .ZN(n6641) );
  INV_X1 U4171 ( .A(n4679), .ZN(n4713) );
  AOI211_X2 U4172 ( .C1(n6691), .C2(n4903), .A(n4902), .B(n4901), .ZN(n4946)
         );
  INV_X1 U4173 ( .A(n6175), .ZN(n6241) );
  INV_X1 U4174 ( .A(n6198), .ZN(n6633) );
  NAND2_X1 U4175 ( .A1(n3555), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6644) );
  AND2_X1 U4176 ( .A1(n4379), .A2(n6855), .ZN(n6680) );
  INV_X1 U4177 ( .A(READY_N), .ZN(n6824) );
  INV_X1 U4178 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6661) );
  INV_X1 U4179 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6799) );
  NAND2_X1 U4180 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6702), .ZN(n6653) );
  OAI21_X1 U4181 ( .B1(n5928), .B2(n6298), .A(n3739), .ZN(U2972) );
  AND2_X2 U4182 ( .A1(n3099), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3101)
         );
  AND2_X2 U4183 ( .A1(n3101), .A2(n4440), .ZN(n3292) );
  AND2_X2 U4184 ( .A1(n3101), .A2(n4441), .ZN(n3168) );
  NOR2_X4 U4185 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4547) );
  AND2_X2 U4186 ( .A1(n3101), .A2(n4537), .ZN(n4027) );
  AOI22_X1 U4187 ( .A1(n4027), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3103) );
  NOR2_X4 U4188 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4565) );
  AND2_X2 U4189 ( .A1(n3101), .A2(n4565), .ZN(n3137) );
  AND2_X2 U4190 ( .A1(n4565), .A2(n4548), .ZN(n3184) );
  AOI22_X1 U4191 ( .A1(n3137), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3102) );
  AND2_X2 U4192 ( .A1(n4547), .A2(n4565), .ZN(n3198) );
  AOI22_X1 U4193 ( .A1(n4077), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3111) );
  INV_X1 U4194 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3106) );
  AOI22_X1 U4195 ( .A1(n3327), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n2969), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3110) );
  AOI22_X1 U4196 ( .A1(n3328), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3154), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3109) );
  AND2_X2 U4197 ( .A1(n4440), .A2(n3107), .ZN(n3263) );
  AOI22_X1 U4198 ( .A1(n3263), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3108) );
  AOI22_X1 U4199 ( .A1(n3327), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3168), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3116) );
  AOI22_X1 U4200 ( .A1(n3154), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3115) );
  AOI22_X1 U4201 ( .A1(n3258), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3114) );
  AOI22_X1 U4202 ( .A1(n4077), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3120) );
  AOI22_X1 U4203 ( .A1(n3292), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3118) );
  AOI22_X1 U4204 ( .A1(n3183), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3127) );
  AOI22_X1 U4205 ( .A1(n3154), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3126) );
  AOI22_X1 U4206 ( .A1(n3258), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3125) );
  AOI22_X1 U4207 ( .A1(n3327), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3168), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3124) );
  AOI22_X1 U4208 ( .A1(n4077), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3131) );
  AOI22_X1 U4209 ( .A1(n3263), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3173), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3130) );
  AOI22_X1 U4210 ( .A1(n4027), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3129) );
  AOI22_X1 U4211 ( .A1(n3292), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3128) );
  INV_X1 U4212 ( .A(n3219), .ZN(n3144) );
  AOI22_X1 U4213 ( .A1(n4027), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3134) );
  AOI22_X1 U4214 ( .A1(n3292), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3133) );
  AOI22_X1 U4215 ( .A1(n3263), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n2969), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3132) );
  AOI22_X1 U4216 ( .A1(n4077), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3135) );
  CLKBUF_X3 U4217 ( .A(n3137), .Z(n4069) );
  AOI22_X1 U4218 ( .A1(n4069), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3141) );
  AOI22_X1 U4219 ( .A1(n3327), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3168), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3140) );
  AOI22_X1 U4220 ( .A1(n3154), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3139) );
  AOI22_X1 U4221 ( .A1(n3258), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3138) );
  NAND2_X1 U4222 ( .A1(n3144), .A2(n3581), .ZN(n3232) );
  AOI22_X1 U4223 ( .A1(n3154), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3148) );
  AOI22_X1 U4224 ( .A1(n3263), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3292), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3147) );
  AOI22_X1 U4225 ( .A1(n4027), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4077), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3146) );
  AOI22_X1 U4226 ( .A1(n3327), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3145) );
  AOI22_X1 U4227 ( .A1(n3198), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3152) );
  AOI22_X1 U4228 ( .A1(n3168), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3151) );
  AOI22_X1 U4229 ( .A1(n3173), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3150) );
  AOI22_X1 U4230 ( .A1(n3328), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3258), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3149) );
  NAND3_X1 U4231 ( .A1(n3153), .A2(n3152), .A3(n3096), .ZN(n3165) );
  AOI22_X1 U4232 ( .A1(n3183), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3158) );
  AOI22_X1 U4233 ( .A1(n3154), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3157) );
  AOI22_X1 U4234 ( .A1(n3258), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3156) );
  AOI22_X1 U4235 ( .A1(n3327), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3168), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3155) );
  AOI22_X1 U4236 ( .A1(n3263), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n2968), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3162) );
  AOI22_X1 U4237 ( .A1(n4077), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3161) );
  AOI22_X1 U4238 ( .A1(n4027), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3160) );
  AOI22_X1 U4239 ( .A1(n3292), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3159) );
  NAND2_X4 U4240 ( .A1(n3164), .A2(n3163), .ZN(n4620) );
  AOI21_X1 U4241 ( .B1(n3232), .B2(n4624), .A(n4620), .ZN(n3182) );
  MUX2_X1 U4242 ( .A(n2950), .B(n3221), .S(n3237), .Z(n3166) );
  NAND2_X1 U4243 ( .A1(n3166), .A2(n3246), .ZN(n3181) );
  AOI22_X1 U4244 ( .A1(n3327), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3168), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3172) );
  AOI22_X1 U4245 ( .A1(n4069), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3171) );
  AOI22_X1 U4246 ( .A1(n3154), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3170) );
  AOI22_X1 U4247 ( .A1(n3258), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3169) );
  NAND4_X1 U4248 ( .A1(n3172), .A2(n3171), .A3(n3170), .A4(n3169), .ZN(n3179)
         );
  AOI22_X1 U4249 ( .A1(n3263), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3173), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3177) );
  AOI22_X1 U4250 ( .A1(n4077), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3176) );
  AOI22_X1 U4251 ( .A1(n4027), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3175) );
  AOI22_X1 U4252 ( .A1(n3292), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3174) );
  NAND4_X1 U4253 ( .A1(n3177), .A2(n3176), .A3(n3175), .A4(n3174), .ZN(n3178)
         );
  NAND2_X1 U4254 ( .A1(n3231), .A2(n3182), .ZN(n3208) );
  NAND2_X1 U4255 ( .A1(n4069), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3188) );
  NAND2_X1 U4256 ( .A1(n3263), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3187) );
  NAND2_X1 U4257 ( .A1(n3328), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3186) );
  NAND2_X1 U4258 ( .A1(n3184), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3185)
         );
  AND4_X2 U4259 ( .A1(n3188), .A2(n3187), .A3(n3186), .A4(n3185), .ZN(n3207)
         );
  NAND2_X1 U4260 ( .A1(n3258), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3193) );
  NAND2_X1 U4261 ( .A1(n3168), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3192) );
  NAND2_X1 U4262 ( .A1(n3154), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3191) );
  NAND2_X1 U4263 ( .A1(n3189), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3190)
         );
  NAND2_X1 U4264 ( .A1(n3292), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3197)
         );
  NAND2_X1 U4265 ( .A1(n3327), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3196) );
  NAND2_X1 U4266 ( .A1(n3173), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3195) );
  NAND2_X1 U4267 ( .A1(n3333), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3194) );
  NAND2_X1 U4268 ( .A1(n4027), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3203)
         );
  NAND2_X1 U4269 ( .A1(n4077), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3202)
         );
  NAND2_X1 U4270 ( .A1(n3198), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3201) );
  NAND2_X1 U4271 ( .A1(n3199), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3200)
         );
  NAND4_X4 U4272 ( .A1(n3207), .A2(n3206), .A3(n3205), .A4(n3204), .ZN(n3249)
         );
  AND2_X1 U4273 ( .A1(n3211), .A2(n4724), .ZN(n3212) );
  NAND2_X2 U4274 ( .A1(n3213), .A2(n3212), .ZN(n4248) );
  NAND2_X1 U4275 ( .A1(n3216), .A2(n4378), .ZN(n4106) );
  NAND2_X1 U4276 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), .ZN(
        n4364) );
  AND2_X1 U4277 ( .A1(n4106), .A2(n4364), .ZN(n3217) );
  NOR2_X1 U4278 ( .A1(n4620), .A2(n3217), .ZN(n3238) );
  INV_X1 U4279 ( .A(n3238), .ZN(n3218) );
  NOR2_X2 U4280 ( .A1(n3219), .A2(n2949), .ZN(n4125) );
  INV_X1 U4281 ( .A(n4125), .ZN(n3220) );
  NAND2_X1 U4282 ( .A1(n3220), .A2(n3404), .ZN(n3222) );
  NAND2_X1 U4283 ( .A1(n2950), .A2(n3235), .ZN(n3559) );
  OR2_X2 U4284 ( .A1(n3559), .A2(n4158), .ZN(n4437) );
  AND2_X2 U4285 ( .A1(n4437), .A2(n3222), .ZN(n3256) );
  NAND2_X2 U4286 ( .A1(n3224), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3319) );
  NAND2_X1 U4287 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4652) );
  OR2_X1 U4288 ( .A1(n6692), .A2(n6022), .ZN(n3227) );
  INV_X1 U4289 ( .A(n3555), .ZN(n3346) );
  NAND2_X1 U4290 ( .A1(n3346), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3226) );
  NAND2_X1 U4291 ( .A1(n3229), .A2(n4125), .ZN(n4115) );
  INV_X1 U4292 ( .A(n4115), .ZN(n3230) );
  NAND2_X1 U4293 ( .A1(n3230), .A2(n3249), .ZN(n4396) );
  NOR2_X1 U4294 ( .A1(n2959), .A2(n4717), .ZN(n3233) );
  NAND2_X1 U4295 ( .A1(n2962), .A2(n3233), .ZN(n4136) );
  AND3_X2 U4296 ( .A1(n3234), .A2(n3246), .A3(n2945), .ZN(n4258) );
  NOR2_X1 U4297 ( .A1(n4620), .A2(n3235), .ZN(n3236) );
  OAI211_X1 U4298 ( .C1(n4396), .C2(n3238), .A(n4136), .B(n4134), .ZN(n3239)
         );
  NAND2_X1 U4299 ( .A1(n3239), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3240) );
  OAI211_X2 U4300 ( .C1(n3319), .C2(n3225), .A(n3241), .B(n3240), .ZN(n3318)
         );
  INV_X1 U4301 ( .A(n3241), .ZN(n3242) );
  NAND2_X1 U4302 ( .A1(n2965), .A2(n3094), .ZN(n3243) );
  MUX2_X1 U4303 ( .A(n3555), .B(n6692), .S(n6207), .Z(n3244) );
  OAI21_X2 U4304 ( .B1(n3319), .B2(n5275), .A(n3244), .ZN(n3272) );
  AND2_X1 U4305 ( .A1(n3399), .A2(n3245), .ZN(n4255) );
  OAI22_X1 U4306 ( .A1(n3247), .A2(n4255), .B1(n3234), .B2(n3246), .ZN(n4253)
         );
  INV_X1 U4307 ( .A(n4253), .ZN(n3257) );
  NAND2_X1 U4308 ( .A1(n3214), .A2(n3209), .ZN(n3248) );
  NAND2_X1 U4309 ( .A1(n3248), .A2(n4638), .ZN(n3250) );
  AND2_X2 U4310 ( .A1(n2945), .A2(n3249), .ZN(n4236) );
  OAI22_X1 U4311 ( .A1(n4248), .A2(n3250), .B1(n4236), .B2(n4620), .ZN(n3254)
         );
  OR2_X1 U4312 ( .A1(n3214), .A2(n3411), .ZN(n4126) );
  INV_X1 U4313 ( .A(n4258), .ZN(n3251) );
  OR2_X1 U4314 ( .A1(n3251), .A2(n3581), .ZN(n3253) );
  INV_X1 U4315 ( .A(n5306), .ZN(n6646) );
  NOR2_X1 U4316 ( .A1(n6646), .A2(n5129), .ZN(n3252) );
  AND4_X2 U4317 ( .A1(n3254), .A2(n4126), .A3(n3253), .A4(n3252), .ZN(n3255)
         );
  INV_X1 U4318 ( .A(n3350), .ZN(n4418) );
  AOI22_X1 U4319 ( .A1(n2970), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3262) );
  AOI22_X1 U4320 ( .A1(n4069), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3261) );
  AOI22_X1 U4321 ( .A1(n4057), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3260) );
  AOI22_X1 U4322 ( .A1(n4072), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3259) );
  NAND4_X1 U4323 ( .A1(n3262), .A2(n3261), .A3(n3260), .A4(n3259), .ZN(n3269)
         );
  AOI22_X1 U4324 ( .A1(n4051), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3267) );
  AOI22_X1 U4325 ( .A1(n2971), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n2946), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3266) );
  AOI22_X1 U4326 ( .A1(n4078), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3265) );
  AOI22_X1 U4327 ( .A1(n4079), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3264) );
  NAND4_X1 U4328 ( .A1(n3267), .A2(n3266), .A3(n3265), .A4(n3264), .ZN(n3268)
         );
  NAND2_X1 U4329 ( .A1(n4418), .A2(n3425), .ZN(n3270) );
  INV_X1 U4330 ( .A(n3271), .ZN(n3311) );
  INV_X1 U4331 ( .A(n3272), .ZN(n3275) );
  INV_X1 U4332 ( .A(n3273), .ZN(n3274) );
  NAND2_X1 U4333 ( .A1(n3275), .A2(n3274), .ZN(n3276) );
  NAND2_X1 U4334 ( .A1(n3276), .A2(n3317), .ZN(n3582) );
  AOI22_X1 U4335 ( .A1(n3327), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3280) );
  AOI22_X1 U4336 ( .A1(n4069), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3279) );
  AOI22_X1 U4337 ( .A1(n4057), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3278) );
  AOI22_X1 U4338 ( .A1(n4072), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3277) );
  NAND4_X1 U4339 ( .A1(n3280), .A2(n3279), .A3(n3278), .A4(n3277), .ZN(n3287)
         );
  AOI22_X1 U4340 ( .A1(n4051), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3285) );
  AOI22_X1 U4341 ( .A1(n4077), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n2946), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3284) );
  AOI22_X1 U4342 ( .A1(n4078), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3283) );
  AOI22_X1 U4343 ( .A1(n4079), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3282) );
  NAND4_X1 U4344 ( .A1(n3285), .A2(n3284), .A3(n3283), .A4(n3282), .ZN(n3286)
         );
  NOR2_X1 U4345 ( .A1(n3485), .A2(n3350), .ZN(n3305) );
  NOR2_X1 U4346 ( .A1(n3350), .A2(n3480), .ZN(n3306) );
  AOI22_X1 U4347 ( .A1(n4051), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3291) );
  AOI22_X1 U4348 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n3327), .B1(n4072), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3290) );
  AOI22_X1 U4349 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n4070), .B1(n4057), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3289) );
  AOI22_X1 U4350 ( .A1(n4077), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3288) );
  NAND4_X1 U4351 ( .A1(n3291), .A2(n3290), .A3(n3289), .A4(n3288), .ZN(n3299)
         );
  AOI22_X1 U4352 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n4052), .B1(n3983), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3297) );
  AOI22_X1 U4353 ( .A1(n4078), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3296) );
  AOI22_X1 U4354 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n4079), .B1(n2946), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3295) );
  AOI22_X1 U4355 ( .A1(n3293), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3294) );
  NAND4_X1 U4356 ( .A1(n3297), .A2(n3296), .A3(n3295), .A4(n3294), .ZN(n3298)
         );
  MUX2_X1 U4357 ( .A(n3305), .B(n3306), .S(n3439), .Z(n3432) );
  INV_X1 U4358 ( .A(n3439), .ZN(n3302) );
  NAND2_X1 U4359 ( .A1(n3540), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3301) );
  AOI21_X1 U4360 ( .B1(n3245), .B2(n3480), .A(n5129), .ZN(n3300) );
  OAI211_X1 U4361 ( .C1(n3302), .C2(n3249), .A(n3301), .B(n3300), .ZN(n3433)
         );
  NAND2_X1 U4362 ( .A1(n3432), .A2(n3433), .ZN(n3303) );
  OAI21_X2 U4363 ( .B1(n3582), .B2(STATE2_REG_0__SCAN_IN), .A(n3303), .ZN(
        n3304) );
  INV_X1 U4364 ( .A(n3304), .ZN(n3431) );
  INV_X1 U4365 ( .A(n3305), .ZN(n3400) );
  NAND2_X1 U4366 ( .A1(n3431), .A2(n3400), .ZN(n3310) );
  XNOR2_X1 U4367 ( .A(n3311), .B(n3310), .ZN(n3421) );
  INV_X1 U4368 ( .A(n3425), .ZN(n3309) );
  NAND2_X1 U4369 ( .A1(n3540), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3308) );
  INV_X1 U4370 ( .A(n3306), .ZN(n3307) );
  NAND2_X1 U4371 ( .A1(n3421), .A2(n3422), .ZN(n3315) );
  INV_X1 U4372 ( .A(n3312), .ZN(n3313) );
  NAND2_X1 U4373 ( .A1(n3310), .A2(n3313), .ZN(n3314) );
  NAND2_X1 U4374 ( .A1(n2964), .A2(n3317), .ZN(n3325) );
  NAND2_X1 U4375 ( .A1(n3325), .A2(n2956), .ZN(n3321) );
  INV_X1 U4376 ( .A(n3319), .ZN(n3344) );
  XNOR2_X1 U4377 ( .A(n4652), .B(n5112), .ZN(n4672) );
  OAI22_X1 U4378 ( .A1(n4672), .A2(n6692), .B1(n3555), .B2(n5112), .ZN(n3320)
         );
  NAND2_X1 U4379 ( .A1(n3321), .A2(n3322), .ZN(n3326) );
  INV_X1 U4380 ( .A(n3322), .ZN(n3323) );
  AOI22_X1 U4381 ( .A1(n2970), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3332) );
  AOI22_X1 U4382 ( .A1(n4069), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3331) );
  AOI22_X1 U4383 ( .A1(n4057), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3330) );
  AOI22_X1 U4384 ( .A1(n4072), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3329) );
  NAND4_X1 U4385 ( .A1(n3332), .A2(n3331), .A3(n3330), .A4(n3329), .ZN(n3339)
         );
  AOI22_X1 U4386 ( .A1(n4051), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3337) );
  AOI22_X1 U4387 ( .A1(n2971), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n2946), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3336) );
  AOI22_X1 U4388 ( .A1(n4078), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3335) );
  AOI22_X1 U4389 ( .A1(n4079), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3334) );
  NAND4_X1 U4390 ( .A1(n3337), .A2(n3336), .A3(n3335), .A4(n3334), .ZN(n3338)
         );
  INV_X1 U4391 ( .A(n3351), .ZN(n3341) );
  AOI22_X1 U4392 ( .A1(n3540), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3341), 
        .B2(n3340), .ZN(n3342) );
  NAND2_X1 U4393 ( .A1(n3344), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3349) );
  NAND2_X1 U4394 ( .A1(n6062), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4763) );
  NAND2_X1 U4395 ( .A1(n4763), .A2(n5116), .ZN(n3345) );
  AND2_X1 U4396 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4667) );
  NAND2_X1 U4397 ( .A1(n6208), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4604) );
  INV_X1 U4398 ( .A(n6692), .ZN(n3347) );
  AOI22_X1 U4399 ( .A1(n4956), .A2(n3347), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3346), .ZN(n3348) );
  AOI22_X1 U4400 ( .A1(n4051), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3355) );
  AOI22_X1 U4401 ( .A1(n4069), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3354) );
  AOI22_X1 U4402 ( .A1(n4079), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n2946), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4403 ( .A1(n4078), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3352) );
  NAND4_X1 U4404 ( .A1(n3355), .A2(n3354), .A3(n3353), .A4(n3352), .ZN(n3361)
         );
  AOI22_X1 U4405 ( .A1(n2970), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4406 ( .A1(n4072), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4407 ( .A1(n2971), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3357) );
  AOI22_X1 U4408 ( .A1(n3293), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3356) );
  NAND4_X1 U4409 ( .A1(n3359), .A2(n3358), .A3(n3357), .A4(n3356), .ZN(n3360)
         );
  AOI22_X1 U4410 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(n3540), .B1(n3553), 
        .B2(n3409), .ZN(n3362) );
  NAND2_X1 U4411 ( .A1(n3540), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4412 ( .A1(n2970), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4413 ( .A1(n4069), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3365) );
  AOI22_X1 U4414 ( .A1(n4057), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3364) );
  AOI22_X1 U4415 ( .A1(n4072), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3363) );
  NAND4_X1 U4416 ( .A1(n3366), .A2(n3365), .A3(n3364), .A4(n3363), .ZN(n3372)
         );
  AOI22_X1 U4417 ( .A1(n4051), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3370) );
  AOI22_X1 U4418 ( .A1(n2971), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n2946), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4419 ( .A1(n4078), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4420 ( .A1(n4079), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3367) );
  NAND4_X1 U4421 ( .A1(n3370), .A2(n3369), .A3(n3368), .A4(n3367), .ZN(n3371)
         );
  NAND2_X1 U4422 ( .A1(n3553), .A2(n3465), .ZN(n3373) );
  NAND2_X1 U4423 ( .A1(n3374), .A2(n3373), .ZN(n3403) );
  NAND2_X1 U4424 ( .A1(n3540), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3386) );
  AOI22_X1 U4425 ( .A1(n4078), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4426 ( .A1(n2970), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3983), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3377) );
  AOI22_X1 U4427 ( .A1(n4057), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3376) );
  AOI22_X1 U4428 ( .A1(n4051), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3375) );
  NAND4_X1 U4429 ( .A1(n3378), .A2(n3377), .A3(n3376), .A4(n3375), .ZN(n3384)
         );
  AOI22_X1 U4430 ( .A1(n4079), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4431 ( .A1(n4052), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3381) );
  AOI22_X1 U4432 ( .A1(n2946), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3380) );
  AOI22_X1 U4433 ( .A1(n4072), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3379) );
  NAND4_X1 U4434 ( .A1(n3382), .A2(n3381), .A3(n3380), .A4(n3379), .ZN(n3383)
         );
  NAND2_X1 U4435 ( .A1(n3553), .A2(n3464), .ZN(n3385) );
  NAND2_X1 U4436 ( .A1(n3386), .A2(n3385), .ZN(n3455) );
  NAND2_X1 U4437 ( .A1(n3540), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3398) );
  AOI22_X1 U4438 ( .A1(n2970), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3390) );
  AOI22_X1 U4439 ( .A1(n3983), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3389) );
  AOI22_X1 U4440 ( .A1(n4057), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3388) );
  AOI22_X1 U4441 ( .A1(n4072), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3387) );
  NAND4_X1 U4442 ( .A1(n3390), .A2(n3389), .A3(n3388), .A4(n3387), .ZN(n3396)
         );
  AOI22_X1 U4443 ( .A1(n4051), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4444 ( .A1(n2971), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n2946), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3393) );
  AOI22_X1 U4445 ( .A1(n4078), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3392) );
  AOI22_X1 U4446 ( .A1(n4079), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3391) );
  NAND4_X1 U4447 ( .A1(n3394), .A2(n3393), .A3(n3392), .A4(n3391), .ZN(n3395)
         );
  NAND2_X1 U4448 ( .A1(n3553), .A2(n3478), .ZN(n3397) );
  INV_X1 U4449 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6802) );
  NAND2_X1 U4450 ( .A1(n3560), .A2(n3399), .ZN(n3407) );
  NAND2_X1 U4451 ( .A1(n3425), .A2(n3439), .ZN(n3424) );
  NAND2_X1 U4452 ( .A1(n3424), .A2(n3418), .ZN(n3410) );
  NAND2_X1 U4453 ( .A1(n3410), .A2(n3409), .ZN(n3467) );
  XNOR2_X1 U4454 ( .A(n3467), .B(n3465), .ZN(n3405) );
  NAND2_X1 U4455 ( .A1(n3405), .A2(n5174), .ZN(n3406) );
  NAND2_X1 U4456 ( .A1(n3407), .A2(n3406), .ZN(n3453) );
  INV_X1 U4457 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4263) );
  XNOR2_X1 U4458 ( .A(n3453), .B(n4263), .ZN(n4831) );
  XNOR2_X1 U4459 ( .A(n3410), .B(n3409), .ZN(n3412) );
  OR2_X1 U4460 ( .A1(n3412), .A2(n3411), .ZN(n3413) );
  OAI21_X2 U4461 ( .B1(n3567), .B2(n3526), .A(n3413), .ZN(n3448) );
  INV_X1 U4462 ( .A(n3448), .ZN(n6492) );
  OR2_X2 U4463 ( .A1(n3415), .A2(n3414), .ZN(n3416) );
  XNOR2_X1 U4464 ( .A(n3424), .B(n3418), .ZN(n3419) );
  AND2_X1 U4465 ( .A1(n3234), .A2(n4638), .ZN(n4254) );
  AOI21_X1 U4466 ( .B1(n3419), .B2(n5174), .A(n4254), .ZN(n3420) );
  AOI21_X1 U4467 ( .B1(n3449), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3452) );
  INV_X1 U4468 ( .A(n3421), .ZN(n3423) );
  NAND2_X1 U4469 ( .A1(n4578), .A2(n3399), .ZN(n3430) );
  OAI21_X1 U4470 ( .B1(n3439), .B2(n3425), .A(n3424), .ZN(n3427) );
  INV_X1 U4471 ( .A(n2961), .ZN(n3426) );
  OAI211_X1 U4472 ( .C1(n3427), .C2(n3411), .A(n3426), .B(n3235), .ZN(n3428)
         );
  INV_X1 U4473 ( .A(n3428), .ZN(n3429) );
  NAND2_X1 U4474 ( .A1(n3430), .A2(n3429), .ZN(n4514) );
  INV_X1 U4475 ( .A(n3432), .ZN(n3435) );
  INV_X1 U4476 ( .A(n3433), .ZN(n3434) );
  INV_X1 U4477 ( .A(n4254), .ZN(n3438) );
  OAI21_X1 U4478 ( .B1(n3411), .B2(n3439), .A(n3438), .ZN(n3440) );
  INV_X1 U4479 ( .A(n3440), .ZN(n3441) );
  OAI21_X1 U4480 ( .B1(n6099), .B2(n3526), .A(n3441), .ZN(n4463) );
  NAND2_X1 U4481 ( .A1(n4463), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3442)
         );
  INV_X1 U4482 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4518) );
  NAND2_X1 U4483 ( .A1(n3442), .A2(n4518), .ZN(n3444) );
  AND2_X1 U4484 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3443) );
  NAND2_X1 U4485 ( .A1(n4463), .A2(n3443), .ZN(n3445) );
  AND2_X1 U4486 ( .A1(n3444), .A2(n3445), .ZN(n4513) );
  NAND2_X1 U4487 ( .A1(n4514), .A2(n4513), .ZN(n3446) );
  NAND2_X2 U4488 ( .A1(n3446), .A2(n3445), .ZN(n6503) );
  NAND2_X1 U4489 ( .A1(n6502), .A2(n6789), .ZN(n3447) );
  NAND3_X1 U4490 ( .A1(n2957), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3450) );
  NAND2_X1 U4491 ( .A1(n3453), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3454)
         );
  INV_X1 U4492 ( .A(n3465), .ZN(n3457) );
  OR2_X1 U4493 ( .A1(n3467), .A2(n3457), .ZN(n3458) );
  XNOR2_X1 U4494 ( .A(n3458), .B(n3464), .ZN(n3459) );
  NAND2_X1 U4495 ( .A1(n3459), .A2(n5174), .ZN(n3460) );
  INV_X1 U4496 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U4497 ( .A1(n3461), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3462)
         );
  NAND2_X1 U4498 ( .A1(n3609), .A2(n3399), .ZN(n3470) );
  NAND2_X1 U4499 ( .A1(n3465), .A2(n3464), .ZN(n3466) );
  OR2_X1 U4500 ( .A1(n3467), .A2(n3466), .ZN(n3477) );
  XNOR2_X1 U4501 ( .A(n3477), .B(n3478), .ZN(n3468) );
  NAND2_X1 U4502 ( .A1(n3468), .A2(n5174), .ZN(n3469) );
  INV_X1 U4503 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4991) );
  NAND2_X1 U4504 ( .A1(n3471), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3472)
         );
  NAND2_X1 U4505 ( .A1(n3553), .A2(n3480), .ZN(n3474) );
  NAND2_X1 U4506 ( .A1(n3540), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3473) );
  NAND2_X1 U4507 ( .A1(n3474), .A2(n3473), .ZN(n3475) );
  INV_X1 U4508 ( .A(n3477), .ZN(n3479) );
  NAND2_X1 U4509 ( .A1(n3479), .A2(n3478), .ZN(n3486) );
  XNOR2_X1 U4510 ( .A(n3486), .B(n3480), .ZN(n3481) );
  NAND2_X1 U4511 ( .A1(n3481), .A2(n5174), .ZN(n3482) );
  INV_X1 U4512 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6536) );
  NAND2_X1 U4513 ( .A1(n3483), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3484)
         );
  NAND2_X1 U4514 ( .A1(n6476), .A2(n3484), .ZN(n5142) );
  OR3_X1 U4515 ( .A1(n3486), .A2(n3485), .A3(n3411), .ZN(n3487) );
  NAND2_X1 U4516 ( .A1(n3492), .A2(n3487), .ZN(n3488) );
  INV_X1 U4517 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6530) );
  XNOR2_X1 U4518 ( .A(n3488), .B(n6530), .ZN(n5141) );
  NAND2_X1 U4519 ( .A1(n5142), .A2(n5141), .ZN(n5140) );
  NAND2_X1 U4520 ( .A1(n3488), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3489)
         );
  NAND2_X1 U4521 ( .A1(n5140), .A2(n3489), .ZN(n5806) );
  INV_X1 U4522 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5807) );
  NAND2_X1 U4523 ( .A1(n3492), .A2(n5807), .ZN(n3490) );
  NAND2_X1 U4524 ( .A1(n5806), .A2(n3490), .ZN(n3745) );
  NAND2_X1 U4525 ( .A1(n4296), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3743)
         );
  NAND2_X1 U4526 ( .A1(n3745), .A2(n3743), .ZN(n5800) );
  INV_X1 U4527 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3491) );
  NAND2_X1 U4528 ( .A1(n3492), .A2(n3491), .ZN(n5798) );
  AND2_X1 U4529 ( .A1(n3492), .A2(n6802), .ZN(n3750) );
  OR2_X1 U4530 ( .A1(n5789), .A2(n3750), .ZN(n3493) );
  NAND2_X1 U4531 ( .A1(n4296), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5799) );
  OAI211_X1 U4532 ( .C1(n5808), .C2(n6802), .A(n3493), .B(n5799), .ZN(n5784)
         );
  INV_X1 U4533 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3740) );
  XNOR2_X1 U4534 ( .A(n5808), .B(n3740), .ZN(n5785) );
  NAND2_X1 U4535 ( .A1(n3492), .A2(n3740), .ZN(n3748) );
  OAI21_X1 U4536 ( .B1(n5784), .B2(n5785), .A(n3748), .ZN(n5779) );
  XNOR2_X1 U4537 ( .A(n5808), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5778)
         );
  NAND2_X1 U4538 ( .A1(n5779), .A2(n5778), .ZN(n5777) );
  OAI21_X1 U4539 ( .B1(n4296), .B2(INSTADDRPOINTER_REG_13__SCAN_IN), .A(n5777), 
        .ZN(n3495) );
  INV_X1 U4540 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5914) );
  XNOR2_X1 U4541 ( .A(n5808), .B(n5914), .ZN(n3494) );
  XNOR2_X1 U4542 ( .A(n3495), .B(n3494), .ZN(n5928) );
  XNOR2_X1 U4543 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3505) );
  AOI21_X1 U4544 ( .B1(n3559), .B2(n3505), .A(n3496), .ZN(n3498) );
  NAND2_X1 U4545 ( .A1(n4121), .A2(n3235), .ZN(n3497) );
  OR2_X1 U4546 ( .A1(n3498), .A2(n3528), .ZN(n3510) );
  INV_X1 U4547 ( .A(n3502), .ZN(n3500) );
  XNOR2_X1 U4548 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3501) );
  INV_X1 U4549 ( .A(n3501), .ZN(n3499) );
  NAND2_X1 U4550 ( .A1(n3500), .A2(n3499), .ZN(n3503) );
  NAND2_X1 U4551 ( .A1(n3502), .A2(n3501), .ZN(n3514) );
  INV_X1 U4552 ( .A(n4108), .ZN(n3509) );
  NAND2_X1 U4553 ( .A1(n3553), .A2(n4620), .ZN(n3504) );
  NAND2_X1 U4554 ( .A1(n3504), .A2(n3235), .ZN(n3511) );
  AND2_X1 U4555 ( .A1(n3553), .A2(n3505), .ZN(n3506) );
  OAI211_X1 U4556 ( .C1(n3511), .C2(n4108), .A(n3506), .B(n3510), .ZN(n3507)
         );
  NAND2_X1 U4557 ( .A1(n3507), .A2(n3543), .ZN(n3508) );
  OAI21_X1 U4558 ( .B1(n3510), .B2(n3509), .A(n3508), .ZN(n3512) );
  NAND2_X1 U4559 ( .A1(n6101), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3513) );
  NAND2_X1 U4560 ( .A1(n3514), .A2(n3513), .ZN(n3522) );
  NAND2_X1 U4561 ( .A1(n5112), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3523) );
  NAND2_X1 U4562 ( .A1(n3515), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3516) );
  INV_X1 U4563 ( .A(n3521), .ZN(n3517) );
  XNOR2_X1 U4564 ( .A(n3522), .B(n3517), .ZN(n4109) );
  NAND2_X1 U4565 ( .A1(n3553), .A2(n4109), .ZN(n3520) );
  INV_X1 U4566 ( .A(n3528), .ZN(n3518) );
  OAI211_X1 U4567 ( .C1(n4109), .C2(n3532), .A(n3520), .B(n3518), .ZN(n3519)
         );
  INV_X1 U4568 ( .A(n3520), .ZN(n3529) );
  NAND2_X1 U4569 ( .A1(n3522), .A2(n3521), .ZN(n3524) );
  XNOR2_X1 U4570 ( .A(n3537), .B(n3534), .ZN(n4107) );
  NOR2_X1 U4571 ( .A1(n3526), .A2(n4107), .ZN(n3527) );
  AOI21_X1 U4572 ( .B1(n3529), .B2(n3528), .A(n3527), .ZN(n3530) );
  INV_X1 U4573 ( .A(n4107), .ZN(n3531) );
  NAND2_X1 U4574 ( .A1(n3532), .A2(n3531), .ZN(n3533) );
  INV_X1 U4575 ( .A(n3553), .ZN(n3538) );
  INV_X1 U4576 ( .A(n4112), .ZN(n3539) );
  AOI22_X1 U4577 ( .A1(n3540), .A2(n3539), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n5129), .ZN(n3541) );
  INV_X1 U4578 ( .A(n3544), .ZN(n3546) );
  NAND2_X1 U4579 ( .A1(n3546), .A2(n3545), .ZN(n3550) );
  INV_X1 U4580 ( .A(n3547), .ZN(n3548) );
  NAND2_X1 U4581 ( .A1(n3548), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3549) );
  NAND2_X1 U4582 ( .A1(n3209), .A2(n3235), .ZN(n3556) );
  NAND2_X1 U4583 ( .A1(n5103), .A2(n3234), .ZN(n3557) );
  NAND2_X1 U4584 ( .A1(n3558), .A2(n3557), .ZN(n4133) );
  NAND2_X1 U4585 ( .A1(n3560), .A2(n3726), .ZN(n3566) );
  NAND2_X1 U4586 ( .A1(n3569), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3568)
         );
  INV_X1 U4587 ( .A(n3601), .ZN(n3561) );
  OAI21_X1 U4588 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n3029), .A(n3561), 
        .ZN(n5551) );
  NAND2_X1 U4589 ( .A1(n4726), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3594) );
  NAND2_X1 U4590 ( .A1(n5280), .A2(EAX_REG_4__SCAN_IN), .ZN(n3563) );
  OAI21_X1 U4591 ( .B1(n6297), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6768), 
        .ZN(n3562) );
  OAI211_X1 U4592 ( .C1(n3594), .C2(n6293), .A(n3563), .B(n3562), .ZN(n3564)
         );
  OAI21_X1 U4593 ( .B1(n5412), .B2(n5551), .A(n3564), .ZN(n3565) );
  NAND2_X1 U4594 ( .A1(n3566), .A2(n3565), .ZN(n4591) );
  NAND2_X1 U4595 ( .A1(n4579), .A2(n3726), .ZN(n3574) );
  OAI21_X1 U4596 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3569), .A(n3568), 
        .ZN(n6500) );
  AOI22_X1 U4597 ( .A1(n3063), .A2(n6500), .B1(n5279), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3571) );
  NAND2_X1 U4598 ( .A1(n5280), .A2(EAX_REG_3__SCAN_IN), .ZN(n3570) );
  OAI211_X1 U4599 ( .C1(n3594), .C2(n3525), .A(n3571), .B(n3570), .ZN(n3572)
         );
  INV_X1 U4600 ( .A(n3572), .ZN(n3573) );
  NAND2_X1 U4601 ( .A1(n3574), .A2(n3573), .ZN(n4789) );
  AND2_X1 U4602 ( .A1(n4591), .A2(n4789), .ZN(n3600) );
  INV_X1 U4603 ( .A(n4577), .ZN(n3575) );
  INV_X1 U4604 ( .A(n5279), .ZN(n3862) );
  NAND2_X1 U4605 ( .A1(n4578), .A2(n3726), .ZN(n3580) );
  AOI22_X1 U4606 ( .A1(n5280), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6768), .ZN(n3578) );
  INV_X1 U4607 ( .A(n3594), .ZN(n3584) );
  NAND2_X1 U4608 ( .A1(n3584), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3577) );
  AND2_X1 U4609 ( .A1(n3578), .A2(n3577), .ZN(n3579) );
  NAND2_X1 U4610 ( .A1(n3580), .A2(n3579), .ZN(n4452) );
  INV_X1 U4611 ( .A(n3581), .ZN(n4257) );
  AOI21_X1 U4612 ( .B1(n6099), .B2(n4257), .A(n6768), .ZN(n4414) );
  OR2_X1 U4614 ( .A1(n3583), .A2(n3882), .ZN(n3588) );
  AOI22_X1 U4615 ( .A1(n5280), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6768), .ZN(n3586) );
  NAND2_X1 U4616 ( .A1(n3584), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3585) );
  AND2_X1 U4617 ( .A1(n3586), .A2(n3585), .ZN(n3587) );
  NAND2_X1 U4618 ( .A1(n3588), .A2(n3587), .ZN(n4413) );
  NAND2_X1 U4619 ( .A1(n4414), .A2(n4413), .ZN(n4412) );
  INV_X1 U4620 ( .A(n4413), .ZN(n3589) );
  NAND2_X1 U4621 ( .A1(n3589), .A2(n5410), .ZN(n3590) );
  NAND2_X1 U4622 ( .A1(n4412), .A2(n3590), .ZN(n4451) );
  NAND2_X1 U4623 ( .A1(n4452), .A2(n4451), .ZN(n4454) );
  OAI21_X1 U4624 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3591), .ZN(n6509) );
  AOI22_X1 U4625 ( .A1(n3063), .A2(n6509), .B1(n5279), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3593) );
  NAND2_X1 U4626 ( .A1(n5280), .A2(EAX_REG_2__SCAN_IN), .ZN(n3592) );
  OAI211_X1 U4627 ( .C1(n3594), .C2(n3515), .A(n3593), .B(n3592), .ZN(n4584)
         );
  NAND2_X1 U4628 ( .A1(n4585), .A2(n4584), .ZN(n3599) );
  INV_X1 U4629 ( .A(n3595), .ZN(n3597) );
  INV_X1 U4630 ( .A(n4454), .ZN(n3596) );
  NAND2_X1 U4631 ( .A1(n3597), .A2(n3596), .ZN(n3598) );
  NAND2_X2 U4632 ( .A1(n3599), .A2(n3598), .ZN(n4788) );
  NAND2_X1 U4633 ( .A1(n3600), .A2(n4788), .ZN(n4791) );
  INV_X1 U4634 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4784) );
  OAI21_X1 U4635 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n3601), .A(n3611), 
        .ZN(n6491) );
  AOI22_X1 U4636 ( .A1(n3063), .A2(n6491), .B1(n5279), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3602) );
  OAI21_X1 U4637 ( .B1(n4092), .B2(n4784), .A(n3602), .ZN(n3603) );
  AOI21_X1 U4638 ( .B1(n3604), .B2(n3726), .A(n3603), .ZN(n4792) );
  INV_X1 U4639 ( .A(n3611), .ZN(n3606) );
  XNOR2_X1 U4640 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .B(n3606), .ZN(n5536) );
  INV_X1 U4641 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4776) );
  OAI22_X1 U4642 ( .A1(n4092), .A2(n4776), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3610), .ZN(n3607) );
  MUX2_X1 U4643 ( .A(n5536), .B(n3607), .S(n5412), .Z(n3608) );
  AOI21_X1 U4644 ( .B1(n3609), .B2(n3726), .A(n3608), .ZN(n4890) );
  OR2_X1 U4645 ( .A1(n3612), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3613) );
  NAND2_X1 U4646 ( .A1(n3613), .A2(n3632), .ZN(n6483) );
  AOI22_X1 U4647 ( .A1(n5280), .A2(EAX_REG_7__SCAN_IN), .B1(n5279), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4648 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n2971), .B1(n4078), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3619) );
  AOI22_X1 U4649 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n4079), .B1(n4551), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4650 ( .A1(n3983), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3617) );
  AOI22_X1 U4651 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(n4057), .B1(n4071), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3616) );
  NAND4_X1 U4652 ( .A1(n3619), .A2(n3618), .A3(n3617), .A4(n3616), .ZN(n3625)
         );
  AOI22_X1 U4653 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n4052), .B1(n2970), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3623) );
  AOI22_X1 U4654 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n4070), .B1(n4072), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3622) );
  AOI22_X1 U4655 ( .A1(n2946), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3621) );
  AOI22_X1 U4656 ( .A1(n4051), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3620) );
  NAND4_X1 U4657 ( .A1(n3623), .A2(n3622), .A3(n3621), .A4(n3620), .ZN(n3624)
         );
  OAI21_X1 U4658 ( .B1(n3625), .B2(n3624), .A(n3726), .ZN(n3628) );
  AOI22_X1 U4659 ( .A1(n5279), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n5410), 
        .B2(n2992), .ZN(n3627) );
  NAND2_X1 U4660 ( .A1(n5280), .A2(EAX_REG_8__SCAN_IN), .ZN(n3626) );
  XNOR2_X1 U4661 ( .A(n3657), .B(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5811) );
  AOI22_X1 U4662 ( .A1(n2970), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3636) );
  AOI22_X1 U4663 ( .A1(n2946), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3635) );
  AOI22_X1 U4664 ( .A1(n3983), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3634) );
  AOI22_X1 U4665 ( .A1(n4051), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3633) );
  NAND4_X1 U4666 ( .A1(n3636), .A2(n3635), .A3(n3634), .A4(n3633), .ZN(n3642)
         );
  AOI22_X1 U4667 ( .A1(n4078), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4668 ( .A1(n4079), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4669 ( .A1(n3293), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4072), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3638) );
  AOI22_X1 U4670 ( .A1(n4057), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3637) );
  NAND4_X1 U4671 ( .A1(n3640), .A2(n3639), .A3(n3638), .A4(n3637), .ZN(n3641)
         );
  OAI21_X1 U4672 ( .B1(n3642), .B2(n3641), .A(n3726), .ZN(n3645) );
  NAND2_X1 U4673 ( .A1(n5280), .A2(EAX_REG_9__SCAN_IN), .ZN(n3644) );
  NAND2_X1 U4674 ( .A1(n5279), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3643)
         );
  NAND3_X1 U4675 ( .A1(n3645), .A2(n3644), .A3(n3643), .ZN(n3646) );
  AOI21_X1 U4676 ( .B1(n5811), .B2(n3063), .A(n3646), .ZN(n5510) );
  AOI22_X1 U4677 ( .A1(n4078), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3650) );
  AOI22_X1 U4678 ( .A1(n2970), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3649) );
  AOI22_X1 U4679 ( .A1(n4079), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3648) );
  AOI22_X1 U4680 ( .A1(n3328), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3647) );
  NAND4_X1 U4681 ( .A1(n3650), .A2(n3649), .A3(n3648), .A4(n3647), .ZN(n3656)
         );
  AOI22_X1 U4682 ( .A1(n3983), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4072), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3654) );
  AOI22_X1 U4683 ( .A1(n4057), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3653) );
  AOI22_X1 U4684 ( .A1(n2946), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3652) );
  AOI22_X1 U4685 ( .A1(n4051), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3651) );
  NAND4_X1 U4686 ( .A1(n3654), .A2(n3653), .A3(n3652), .A4(n3651), .ZN(n3655)
         );
  NOR2_X1 U4687 ( .A1(n3656), .A2(n3655), .ZN(n3664) );
  NAND2_X1 U4688 ( .A1(n3657), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3659)
         );
  INV_X1 U4689 ( .A(n3659), .ZN(n3658) );
  INV_X1 U4690 ( .A(n3688), .ZN(n3661) );
  INV_X1 U4691 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6743) );
  NAND2_X1 U4692 ( .A1(n6743), .A2(n3659), .ZN(n3660) );
  NAND2_X1 U4693 ( .A1(n3661), .A2(n3660), .ZN(n6353) );
  AOI22_X1 U4694 ( .A1(n6353), .A2(n3063), .B1(n5279), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3663) );
  NAND2_X1 U4695 ( .A1(n5280), .A2(EAX_REG_10__SCAN_IN), .ZN(n3662) );
  OAI211_X1 U4696 ( .C1(n3882), .C2(n3664), .A(n3663), .B(n3662), .ZN(n5619)
         );
  AOI22_X1 U4697 ( .A1(n4079), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4698 ( .A1(n4052), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4699 ( .A1(n4057), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3666) );
  AOI22_X1 U4700 ( .A1(n2946), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3665) );
  NAND4_X1 U4701 ( .A1(n3668), .A2(n3667), .A3(n3666), .A4(n3665), .ZN(n3674)
         );
  AOI22_X1 U4702 ( .A1(n4051), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U4703 ( .A1(n2970), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3983), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4704 ( .A1(n4078), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4705 ( .A1(n4072), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3669) );
  NAND4_X1 U4706 ( .A1(n3672), .A2(n3671), .A3(n3670), .A4(n3669), .ZN(n3673)
         );
  NOR2_X1 U4707 ( .A1(n3674), .A2(n3673), .ZN(n3677) );
  XNOR2_X1 U4708 ( .A(n3688), .B(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5793)
         );
  AOI22_X1 U4709 ( .A1(n5793), .A2(n3063), .B1(n5279), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3676) );
  NAND2_X1 U4710 ( .A1(n5280), .A2(EAX_REG_11__SCAN_IN), .ZN(n3675) );
  OAI211_X1 U4711 ( .C1(n3882), .C2(n3677), .A(n3676), .B(n3675), .ZN(n5497)
         );
  AND2_X1 U4712 ( .A1(n3890), .A2(n5497), .ZN(n5403) );
  INV_X1 U4713 ( .A(n5403), .ZN(n5610) );
  AOI22_X1 U4714 ( .A1(n4051), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n2970), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3681) );
  AOI22_X1 U4715 ( .A1(n4052), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3983), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3680) );
  AOI22_X1 U4716 ( .A1(n4079), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n2946), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3679) );
  AOI22_X1 U4717 ( .A1(n4070), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3678) );
  NAND4_X1 U4718 ( .A1(n3681), .A2(n3680), .A3(n3679), .A4(n3678), .ZN(n3687)
         );
  AOI22_X1 U4719 ( .A1(n3293), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4720 ( .A1(n4072), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3684) );
  AOI22_X1 U4721 ( .A1(n4078), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4722 ( .A1(n2971), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3682) );
  NAND4_X1 U4723 ( .A1(n3685), .A2(n3684), .A3(n3683), .A4(n3682), .ZN(n3686)
         );
  OAI21_X1 U4724 ( .B1(n3687), .B2(n3686), .A(n3726), .ZN(n3694) );
  INV_X1 U4725 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6791) );
  OAI21_X1 U4726 ( .B1(n4724), .B2(n6791), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n3692) );
  OAI21_X1 U4727 ( .B1(n3689), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n3696), 
        .ZN(n6349) );
  OAI22_X1 U4728 ( .A1(n6349), .A2(n5412), .B1(PHYADDRPOINTER_REG_12__SCAN_IN), 
        .B2(n3862), .ZN(n3690) );
  INV_X1 U4729 ( .A(n3690), .ZN(n3691) );
  NAND2_X1 U4730 ( .A1(n3692), .A2(n3691), .ZN(n3693) );
  NAND2_X1 U4731 ( .A1(n5280), .A2(EAX_REG_13__SCAN_IN), .ZN(n3699) );
  OAI21_X1 U4732 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3697), .A(n3876), 
        .ZN(n6329) );
  AOI22_X1 U4733 ( .A1(n5410), .A2(n6329), .B1(n5279), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3698) );
  NAND2_X1 U4734 ( .A1(n3699), .A2(n3698), .ZN(n3884) );
  INV_X1 U4735 ( .A(n3884), .ZN(n3711) );
  AOI22_X1 U4736 ( .A1(n2970), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4737 ( .A1(n3983), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3702) );
  AOI22_X1 U4738 ( .A1(n4057), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3701) );
  AOI22_X1 U4739 ( .A1(n4072), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3700) );
  NAND4_X1 U4740 ( .A1(n3703), .A2(n3702), .A3(n3701), .A4(n3700), .ZN(n3709)
         );
  AOI22_X1 U4741 ( .A1(n4051), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3707) );
  AOI22_X1 U4742 ( .A1(n2971), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n2946), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4743 ( .A1(n4078), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4744 ( .A1(n4079), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3704) );
  NAND4_X1 U4745 ( .A1(n3707), .A2(n3706), .A3(n3705), .A4(n3704), .ZN(n3708)
         );
  OR2_X1 U4746 ( .A1(n3709), .A2(n3708), .ZN(n3710) );
  AND2_X1 U4747 ( .A1(n3726), .A2(n3710), .ZN(n5601) );
  INV_X1 U4748 ( .A(n5601), .ZN(n3712) );
  INV_X1 U4749 ( .A(EAX_REG_14__SCAN_IN), .ZN(n5186) );
  INV_X1 U4750 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5168) );
  OAI22_X1 U4751 ( .A1(n4092), .A2(n5186), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5168), .ZN(n3713) );
  NAND2_X1 U4752 ( .A1(n3713), .A2(n5412), .ZN(n3728) );
  AOI22_X1 U4753 ( .A1(n4051), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4079), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4754 ( .A1(n2970), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3983), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4755 ( .A1(n4072), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3715) );
  AOI22_X1 U4756 ( .A1(n4078), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3714) );
  NAND4_X1 U4757 ( .A1(n3717), .A2(n3716), .A3(n3715), .A4(n3714), .ZN(n3723)
         );
  AOI22_X1 U4758 ( .A1(n2971), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4759 ( .A1(n4052), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4760 ( .A1(n2946), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4761 ( .A1(n4057), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3718) );
  NAND4_X1 U4762 ( .A1(n3721), .A2(n3720), .A3(n3719), .A4(n3718), .ZN(n3722)
         );
  OR2_X1 U4763 ( .A1(n3723), .A2(n3722), .ZN(n3725) );
  XNOR2_X1 U4764 ( .A(n3876), .B(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5162)
         );
  NOR2_X1 U4765 ( .A1(n5162), .A2(n5412), .ZN(n3724) );
  AOI21_X1 U4766 ( .B1(n3726), .B2(n3725), .A(n3724), .ZN(n3727) );
  NAND2_X1 U4767 ( .A1(n3728), .A2(n3727), .ZN(n3883) );
  NAND2_X1 U4768 ( .A1(n3729), .A2(n3883), .ZN(n5486) );
  OAI21_X1 U4769 ( .B1(n3729), .B2(n3883), .A(n5486), .ZN(n5148) );
  NAND2_X1 U4770 ( .A1(n5129), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5151) );
  NOR2_X1 U4771 ( .A1(n5148), .A2(n5816), .ZN(n3738) );
  NAND2_X1 U4772 ( .A1(n6692), .A2(n6691), .ZN(n3730) );
  NAND2_X1 U4773 ( .A1(n3730), .A2(n5129), .ZN(n3731) );
  NAND2_X1 U4774 ( .A1(n5129), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3733) );
  NAND2_X1 U4775 ( .A1(n6297), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3732) );
  NAND2_X1 U4776 ( .A1(n3733), .A2(n3732), .ZN(n4465) );
  NAND2_X1 U4777 ( .A1(n5764), .A2(n5162), .ZN(n3736) );
  NAND2_X1 U4778 ( .A1(n6573), .A2(REIP_REG_14__SCAN_IN), .ZN(n5916) );
  OAI21_X1 U4779 ( .B1(n5762), .B2(n5168), .A(n5916), .ZN(n3734) );
  NOR2_X1 U4780 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3741) );
  INV_X1 U4781 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5929) );
  NAND4_X1 U4782 ( .A1(n3741), .A2(n5914), .A3(n5929), .A4(n3740), .ZN(n3742)
         );
  NAND2_X1 U4783 ( .A1(n4296), .A2(n3742), .ZN(n5729) );
  AND2_X1 U4784 ( .A1(n3743), .A2(n5729), .ZN(n3744) );
  NAND2_X1 U4785 ( .A1(n3745), .A2(n3744), .ZN(n3755) );
  NAND2_X1 U4786 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3746) );
  NAND2_X1 U4787 ( .A1(n3492), .A2(n3746), .ZN(n3747) );
  NAND2_X1 U4788 ( .A1(n3748), .A2(n3747), .ZN(n3749) );
  AND2_X1 U4789 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4271) );
  AND2_X1 U4790 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4283) );
  NAND2_X1 U4791 ( .A1(n4271), .A2(n4283), .ZN(n3751) );
  AND2_X1 U4792 ( .A1(n3492), .A2(n3751), .ZN(n3752) );
  NOR2_X1 U4793 ( .A1(n5728), .A2(n3752), .ZN(n3753) );
  AND2_X1 U4794 ( .A1(n5798), .A2(n3753), .ZN(n3754) );
  AOI21_X2 U4795 ( .B1(n3755), .B2(n3754), .A(n2979), .ZN(n3758) );
  INV_X1 U4796 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5889) );
  INV_X1 U4797 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U4798 ( .A1(n5889), .A2(n5899), .ZN(n5730) );
  OAI21_X1 U4799 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5730), .A(n4296), 
        .ZN(n3756) );
  INV_X1 U4800 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3757) );
  XNOR2_X1 U4801 ( .A(n5808), .B(n6838), .ZN(n5712) );
  XNOR2_X1 U4802 ( .A(n4296), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5706)
         );
  NOR2_X2 U4803 ( .A1(n5705), .A2(n5706), .ZN(n4332) );
  INV_X1 U4804 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3760) );
  NAND2_X1 U4805 ( .A1(n5808), .A2(n4349), .ZN(n4307) );
  NOR3_X1 U4806 ( .A1(n4307), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n3760), 
        .ZN(n3759) );
  AOI21_X1 U4807 ( .B1(INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n3760), .A(n3759), 
        .ZN(n3766) );
  NOR2_X1 U4808 ( .A1(n5808), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4333)
         );
  NAND2_X1 U4809 ( .A1(n4333), .A2(n3760), .ZN(n3762) );
  NAND3_X1 U4810 ( .A1(n5808), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n4349), .ZN(n3761) );
  NAND3_X1 U4811 ( .A1(n3762), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n3761), .ZN(n3765) );
  AND2_X1 U4812 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4288) );
  INV_X1 U4813 ( .A(n4288), .ZN(n4275) );
  OAI21_X1 U4814 ( .B1(n3762), .B2(INSTADDRPOINTER_REG_24__SCAN_IN), .A(n4275), 
        .ZN(n3763) );
  NAND2_X1 U4815 ( .A1(n4332), .A2(n3763), .ZN(n3764) );
  OAI211_X1 U4816 ( .C1(n4332), .C2(n3766), .A(n3765), .B(n3764), .ZN(n5842)
         );
  NAND2_X1 U4817 ( .A1(n5842), .A2(n6505), .ZN(n3959) );
  AOI22_X1 U4818 ( .A1(n4079), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4819 ( .A1(n4051), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3769) );
  AOI22_X1 U4820 ( .A1(n4052), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4821 ( .A1(n2946), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3767) );
  NAND4_X1 U4822 ( .A1(n3770), .A2(n3769), .A3(n3768), .A4(n3767), .ZN(n3776)
         );
  AOI22_X1 U4823 ( .A1(n2970), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3983), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4824 ( .A1(n4072), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4825 ( .A1(n4078), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4826 ( .A1(n3293), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3771) );
  NAND4_X1 U4827 ( .A1(n3774), .A2(n3773), .A3(n3772), .A4(n3771), .ZN(n3775)
         );
  OR2_X1 U4828 ( .A1(n3776), .A2(n3775), .ZN(n3777) );
  NAND2_X1 U4829 ( .A1(n4095), .A2(n3777), .ZN(n3779) );
  AOI22_X1 U4830 ( .A1(n5280), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6768), .ZN(n3778) );
  NAND2_X1 U4831 ( .A1(n3779), .A2(n3778), .ZN(n5413) );
  AOI22_X1 U4832 ( .A1(n4052), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3983), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4833 ( .A1(n3293), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4072), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4834 ( .A1(n4057), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4835 ( .A1(n4551), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n2946), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3780) );
  NAND4_X1 U4836 ( .A1(n3783), .A2(n3782), .A3(n3781), .A4(n3780), .ZN(n3789)
         );
  AOI22_X1 U4837 ( .A1(n4051), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4079), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4838 ( .A1(n4078), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4839 ( .A1(n2970), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4840 ( .A1(n2971), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3784) );
  NAND4_X1 U4841 ( .A1(n3787), .A2(n3786), .A3(n3785), .A4(n3784), .ZN(n3788)
         );
  OR2_X1 U4842 ( .A1(n3789), .A2(n3788), .ZN(n3790) );
  NAND2_X1 U4843 ( .A1(n4095), .A2(n3790), .ZN(n3792) );
  AOI22_X1 U4844 ( .A1(n5280), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6768), .ZN(n3791) );
  NAND2_X1 U4845 ( .A1(n3792), .A2(n3791), .ZN(n5411) );
  NAND3_X1 U4846 ( .A1(n5413), .A2(n5411), .A3(n5412), .ZN(n3820) );
  AOI22_X1 U4847 ( .A1(n4051), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4848 ( .A1(n2970), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4849 ( .A1(n4057), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4850 ( .A1(n4078), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3793) );
  NAND4_X1 U4851 ( .A1(n3796), .A2(n3795), .A3(n3794), .A4(n3793), .ZN(n3802)
         );
  AOI22_X1 U4852 ( .A1(n4079), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3800) );
  AOI22_X1 U4853 ( .A1(n3983), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3799) );
  AOI22_X1 U4854 ( .A1(n2946), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4855 ( .A1(n4072), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3797) );
  NAND4_X1 U4856 ( .A1(n3800), .A2(n3799), .A3(n3798), .A4(n3797), .ZN(n3801)
         );
  OR2_X1 U4857 ( .A1(n3802), .A2(n3801), .ZN(n3803) );
  NAND2_X1 U4858 ( .A1(n4095), .A2(n3803), .ZN(n3805) );
  AOI22_X1 U4859 ( .A1(n5280), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6768), .ZN(n3804) );
  NAND2_X1 U4860 ( .A1(n3805), .A2(n3804), .ZN(n5405) );
  AOI22_X1 U4861 ( .A1(n4079), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n2970), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4862 ( .A1(n4052), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3983), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4863 ( .A1(n4057), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4864 ( .A1(n2946), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3806) );
  NAND4_X1 U4865 ( .A1(n3809), .A2(n3808), .A3(n3807), .A4(n3806), .ZN(n3815)
         );
  AOI22_X1 U4866 ( .A1(n4051), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3813) );
  AOI22_X1 U4867 ( .A1(n3293), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4868 ( .A1(n4078), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4869 ( .A1(n4072), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3810) );
  NAND4_X1 U4870 ( .A1(n3813), .A2(n3812), .A3(n3811), .A4(n3810), .ZN(n3814)
         );
  OR2_X1 U4871 ( .A1(n3815), .A2(n3814), .ZN(n3816) );
  NAND2_X1 U4872 ( .A1(n4095), .A2(n3816), .ZN(n3818) );
  AOI22_X1 U4873 ( .A1(n5280), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6768), .ZN(n3817) );
  NAND2_X1 U4874 ( .A1(n3818), .A2(n3817), .ZN(n5407) );
  NAND2_X1 U4875 ( .A1(n5405), .A2(n5407), .ZN(n3819) );
  OR2_X1 U4876 ( .A1(n3820), .A2(n3819), .ZN(n3850) );
  INV_X1 U4877 ( .A(n3844), .ZN(n3828) );
  INV_X1 U4878 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3822) );
  XNOR2_X1 U4879 ( .A(n3828), .B(n3822), .ZN(n5716) );
  NAND2_X1 U4880 ( .A1(n3823), .A2(n5749), .ZN(n3824) );
  NAND2_X1 U4881 ( .A1(n3826), .A2(n3824), .ZN(n5476) );
  AND2_X1 U4882 ( .A1(n5476), .A2(n5410), .ZN(n3829) );
  XNOR2_X1 U4883 ( .A(n3826), .B(n3825), .ZN(n5735) );
  NAND2_X1 U4884 ( .A1(n3019), .A2(n3018), .ZN(n3827) );
  NAND2_X1 U4885 ( .A1(n3828), .A2(n3827), .ZN(n5724) );
  NAND4_X1 U4886 ( .A1(n5716), .A2(n3829), .A3(n5735), .A4(n5724), .ZN(n3849)
         );
  AOI22_X1 U4887 ( .A1(n4051), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4888 ( .A1(n2970), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4889 ( .A1(n4072), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4890 ( .A1(n4052), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3830) );
  NAND4_X1 U4891 ( .A1(n3833), .A2(n3832), .A3(n3831), .A4(n3830), .ZN(n3839)
         );
  AOI22_X1 U4892 ( .A1(n4079), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3983), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4893 ( .A1(n3293), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4894 ( .A1(n4078), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4895 ( .A1(n2946), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3834) );
  NAND4_X1 U4896 ( .A1(n3837), .A2(n3836), .A3(n3835), .A4(n3834), .ZN(n3838)
         );
  NOR2_X1 U4897 ( .A1(n3839), .A2(n3838), .ZN(n3843) );
  OAI21_X1 U4898 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6297), .A(n6768), 
        .ZN(n3840) );
  INV_X1 U4899 ( .A(n3840), .ZN(n3841) );
  AOI21_X1 U4900 ( .B1(n5280), .B2(EAX_REG_21__SCAN_IN), .A(n3841), .ZN(n3842)
         );
  OAI21_X1 U4901 ( .B1(n4066), .B2(n3843), .A(n3842), .ZN(n3848) );
  NAND2_X1 U4902 ( .A1(n3845), .A2(n6841), .ZN(n3846) );
  NAND2_X1 U4903 ( .A1(n3906), .A2(n3846), .ZN(n5708) );
  OR2_X1 U4904 ( .A1(n5708), .A2(n5412), .ZN(n3847) );
  NAND2_X1 U4905 ( .A1(n3848), .A2(n3847), .ZN(n5415) );
  AOI21_X1 U4906 ( .B1(n3850), .B2(n3849), .A(n5415), .ZN(n3887) );
  AOI22_X1 U4907 ( .A1(n4078), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4908 ( .A1(n3328), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4072), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3853) );
  AOI22_X1 U4909 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n4070), .B1(n4057), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3852) );
  AOI22_X1 U4910 ( .A1(n4051), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3851) );
  NAND4_X1 U4911 ( .A1(n3854), .A2(n3853), .A3(n3852), .A4(n3851), .ZN(n3860)
         );
  AOI22_X1 U4912 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n2970), .B1(n4052), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4913 ( .A1(n4079), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4914 ( .A1(n2946), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4915 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n3983), .B1(n4071), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3855) );
  NAND4_X1 U4916 ( .A1(n3858), .A2(n3857), .A3(n3856), .A4(n3855), .ZN(n3859)
         );
  OR2_X1 U4917 ( .A1(n3860), .A2(n3859), .ZN(n3861) );
  NAND2_X1 U4918 ( .A1(n4095), .A2(n3861), .ZN(n3865) );
  XNOR2_X1 U4919 ( .A(n3877), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6322)
         );
  INV_X1 U4920 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5761) );
  OAI22_X1 U4921 ( .A1(n6322), .A2(n5412), .B1(n5761), .B2(n3862), .ZN(n3863)
         );
  AOI21_X1 U4922 ( .B1(n5280), .B2(EAX_REG_16__SCAN_IN), .A(n3863), .ZN(n3864)
         );
  NAND2_X1 U4923 ( .A1(n3865), .A2(n3864), .ZN(n5591) );
  INV_X1 U4924 ( .A(n5591), .ZN(n3886) );
  AOI22_X1 U4925 ( .A1(n4078), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3869) );
  AOI22_X1 U4926 ( .A1(n2970), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4927 ( .A1(n4072), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3867) );
  AOI22_X1 U4928 ( .A1(n3293), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3866) );
  NAND4_X1 U4929 ( .A1(n3869), .A2(n3868), .A3(n3867), .A4(n3866), .ZN(n3875)
         );
  AOI22_X1 U4930 ( .A1(n4051), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4931 ( .A1(n3983), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4932 ( .A1(n2946), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4933 ( .A1(n4079), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3870) );
  NAND4_X1 U4934 ( .A1(n3873), .A2(n3872), .A3(n3871), .A4(n3870), .ZN(n3874)
         );
  NOR2_X1 U4935 ( .A1(n3875), .A2(n3874), .ZN(n3881) );
  INV_X1 U4936 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6756) );
  OAI21_X1 U4937 ( .B1(n3876), .B2(n5168), .A(n6756), .ZN(n3878) );
  NAND2_X1 U4938 ( .A1(n3878), .A2(n3877), .ZN(n5773) );
  AOI22_X1 U4939 ( .A1(n5773), .A2(n3063), .B1(PHYADDRPOINTER_REG_15__SCAN_IN), 
        .B2(n5279), .ZN(n3880) );
  NAND2_X1 U4940 ( .A1(n5280), .A2(EAX_REG_15__SCAN_IN), .ZN(n3879) );
  OAI211_X1 U4941 ( .C1(n3882), .C2(n3881), .A(n3880), .B(n3879), .ZN(n5483)
         );
  OAI211_X1 U4942 ( .C1(n5601), .C2(n3884), .A(n3883), .B(n5483), .ZN(n3885)
         );
  NOR2_X1 U4943 ( .A1(n3886), .A2(n5484), .ZN(n5402) );
  AND2_X1 U4944 ( .A1(n3887), .A2(n5402), .ZN(n3888) );
  AND2_X1 U4945 ( .A1(n3888), .A2(n5497), .ZN(n3889) );
  AOI22_X1 U4946 ( .A1(n2970), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4947 ( .A1(n3983), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4948 ( .A1(n4057), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4949 ( .A1(n4072), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3891) );
  NAND4_X1 U4950 ( .A1(n3894), .A2(n3893), .A3(n3892), .A4(n3891), .ZN(n3900)
         );
  AOI22_X1 U4951 ( .A1(n4051), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3898) );
  AOI22_X1 U4952 ( .A1(n2971), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n2946), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4953 ( .A1(n4078), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4954 ( .A1(n4079), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3895) );
  NAND4_X1 U4955 ( .A1(n3898), .A2(n3897), .A3(n3896), .A4(n3895), .ZN(n3899)
         );
  NOR2_X1 U4956 ( .A1(n3900), .A2(n3899), .ZN(n3903) );
  AOI21_X1 U4957 ( .B1(n4340), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3901) );
  AOI21_X1 U4958 ( .B1(n5280), .B2(EAX_REG_22__SCAN_IN), .A(n3901), .ZN(n3902)
         );
  OAI21_X1 U4959 ( .B1(n4066), .B2(n3903), .A(n3902), .ZN(n3905) );
  XNOR2_X1 U4960 ( .A(n3906), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5391)
         );
  NAND2_X1 U4961 ( .A1(n5391), .A2(n5410), .ZN(n3904) );
  NAND2_X1 U4962 ( .A1(n3905), .A2(n3904), .ZN(n4337) );
  INV_X1 U4963 ( .A(n3907), .ZN(n3908) );
  INV_X1 U4964 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5382) );
  NAND2_X1 U4965 ( .A1(n3908), .A2(n5382), .ZN(n3909) );
  NAND2_X1 U4966 ( .A1(n3964), .A2(n3909), .ZN(n5381) );
  AOI22_X1 U4967 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n4079), .B1(n4051), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4968 ( .A1(n2970), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4969 ( .A1(n4052), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4970 ( .A1(n3281), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3910) );
  NAND4_X1 U4971 ( .A1(n3913), .A2(n3912), .A3(n3911), .A4(n3910), .ZN(n3919)
         );
  AOI22_X1 U4972 ( .A1(n2971), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3983), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4973 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n4072), .B1(n4070), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4974 ( .A1(n4078), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n2946), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4975 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n3293), .B1(n4071), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3914) );
  NAND4_X1 U4976 ( .A1(n3917), .A2(n3916), .A3(n3915), .A4(n3914), .ZN(n3918)
         );
  NOR2_X1 U4977 ( .A1(n3919), .A2(n3918), .ZN(n3937) );
  AOI22_X1 U4978 ( .A1(n2970), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4979 ( .A1(n3983), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4980 ( .A1(n4078), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n2946), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3921) );
  AOI22_X1 U4981 ( .A1(n4079), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3920) );
  NAND4_X1 U4982 ( .A1(n3923), .A2(n3922), .A3(n3921), .A4(n3920), .ZN(n3929)
         );
  AOI22_X1 U4983 ( .A1(n4051), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4984 ( .A1(n4072), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3926) );
  AOI22_X1 U4985 ( .A1(n2971), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3925) );
  AOI22_X1 U4986 ( .A1(n3293), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3924) );
  NAND4_X1 U4987 ( .A1(n3927), .A2(n3926), .A3(n3925), .A4(n3924), .ZN(n3928)
         );
  NOR2_X1 U4988 ( .A1(n3929), .A2(n3928), .ZN(n3938) );
  XNOR2_X1 U4989 ( .A(n3937), .B(n3938), .ZN(n3933) );
  NAND2_X1 U4990 ( .A1(n6768), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3930)
         );
  NAND2_X1 U4991 ( .A1(n5412), .A2(n3930), .ZN(n3931) );
  AOI21_X1 U4992 ( .B1(n5280), .B2(EAX_REG_23__SCAN_IN), .A(n3931), .ZN(n3932)
         );
  OAI21_X1 U4993 ( .B1(n4066), .B2(n3933), .A(n3932), .ZN(n3934) );
  NAND2_X1 U4994 ( .A1(n3935), .A2(n3934), .ZN(n4322) );
  XNOR2_X1 U4995 ( .A(n3964), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5368)
         );
  NOR2_X1 U4996 ( .A1(n3938), .A2(n3937), .ZN(n3991) );
  AOI22_X1 U4997 ( .A1(n2970), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4998 ( .A1(n3983), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4999 ( .A1(n4057), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3940) );
  AOI22_X1 U5000 ( .A1(n4072), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3939) );
  NAND4_X1 U5001 ( .A1(n3942), .A2(n3941), .A3(n3940), .A4(n3939), .ZN(n3948)
         );
  AOI22_X1 U5002 ( .A1(n4051), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U5003 ( .A1(n2971), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n2946), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U5004 ( .A1(n4078), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U5005 ( .A1(n4079), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3943) );
  NAND4_X1 U5006 ( .A1(n3946), .A2(n3945), .A3(n3944), .A4(n3943), .ZN(n3947)
         );
  OR2_X1 U5007 ( .A1(n3948), .A2(n3947), .ZN(n3990) );
  INV_X1 U5008 ( .A(n3990), .ZN(n3949) );
  XNOR2_X1 U5009 ( .A(n3991), .B(n3949), .ZN(n3950) );
  NAND2_X1 U5010 ( .A1(n3950), .A2(n4095), .ZN(n3952) );
  AOI22_X1 U5011 ( .A1(n5280), .A2(EAX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n5279), .ZN(n3951) );
  OAI211_X1 U5012 ( .C1(n5368), .C2(n5412), .A(n3952), .B(n3951), .ZN(n3954)
         );
  NAND2_X2 U5013 ( .A1(n3953), .A2(n3954), .ZN(n5194) );
  OAI21_X1 U5014 ( .B1(n3953), .B2(n3954), .A(n5194), .ZN(n5646) );
  NAND2_X1 U5015 ( .A1(n6573), .A2(REIP_REG_24__SCAN_IN), .ZN(n5843) );
  OAI21_X1 U5016 ( .B1(n5762), .B2(n3963), .A(n5843), .ZN(n3955) );
  AOI21_X1 U5017 ( .B1(n5764), .B2(n5368), .A(n3955), .ZN(n3956) );
  NAND2_X1 U5018 ( .A1(n3959), .A2(n3958), .ZN(U2962) );
  NOR2_X1 U5019 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4350) );
  NOR2_X1 U5020 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5845) );
  AND2_X1 U5021 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5863) );
  INV_X1 U5022 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5822) );
  INV_X1 U5023 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5247) );
  NAND2_X1 U5024 ( .A1(n5822), .A2(n5247), .ZN(n5244) );
  NAND2_X1 U5025 ( .A1(n5690), .A2(n4101), .ZN(n5252) );
  AND2_X1 U5026 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5828) );
  AND2_X1 U5027 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5243) );
  NAND3_X1 U5028 ( .A1(n5808), .A2(n5828), .A3(n5243), .ZN(n3960) );
  NAND2_X1 U5029 ( .A1(n4102), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3961) );
  XNOR2_X1 U5030 ( .A(n3962), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5239)
         );
  INV_X1 U5031 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4015) );
  INV_X1 U5032 ( .A(n4018), .ZN(n3965) );
  INV_X1 U5033 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5216) );
  NAND2_X1 U5034 ( .A1(n3966), .A2(n5216), .ZN(n3967) );
  NAND2_X1 U5035 ( .A1(n4045), .A2(n3967), .ZN(n5210) );
  AOI22_X1 U5036 ( .A1(n4078), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3971) );
  AOI22_X1 U5037 ( .A1(n4051), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3983), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3970) );
  AOI22_X1 U5038 ( .A1(n4079), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3969) );
  AOI22_X1 U5039 ( .A1(n4057), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3968) );
  NAND4_X1 U5040 ( .A1(n3971), .A2(n3970), .A3(n3969), .A4(n3968), .ZN(n3977)
         );
  AOI22_X1 U5041 ( .A1(n2970), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U5042 ( .A1(n4052), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U5043 ( .A1(n4072), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U5044 ( .A1(n2946), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3972) );
  NAND4_X1 U5045 ( .A1(n3975), .A2(n3974), .A3(n3973), .A4(n3972), .ZN(n3976)
         );
  NOR2_X1 U5046 ( .A1(n3977), .A2(n3976), .ZN(n4039) );
  AOI22_X1 U5047 ( .A1(n4051), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U5048 ( .A1(n2971), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n2946), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U5049 ( .A1(n4078), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U5050 ( .A1(n4079), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3979) );
  NAND4_X1 U5051 ( .A1(n3982), .A2(n3981), .A3(n3980), .A4(n3979), .ZN(n3989)
         );
  AOI22_X1 U5052 ( .A1(n2970), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3987) );
  AOI22_X1 U5053 ( .A1(n3983), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3986) );
  AOI22_X1 U5054 ( .A1(n4057), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U5055 ( .A1(n4072), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3984) );
  NAND4_X1 U5056 ( .A1(n3987), .A2(n3986), .A3(n3985), .A4(n3984), .ZN(n3988)
         );
  NOR2_X1 U5057 ( .A1(n3989), .A2(n3988), .ZN(n4020) );
  NAND2_X1 U5058 ( .A1(n3991), .A2(n3990), .ZN(n4019) );
  NOR2_X1 U5059 ( .A1(n4020), .A2(n4019), .ZN(n4008) );
  AOI22_X1 U5060 ( .A1(n2970), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U5061 ( .A1(n3983), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U5062 ( .A1(n4057), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U5063 ( .A1(n4072), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3992) );
  NAND4_X1 U5064 ( .A1(n3995), .A2(n3994), .A3(n3993), .A4(n3992), .ZN(n4001)
         );
  AOI22_X1 U5065 ( .A1(n4051), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U5066 ( .A1(n2971), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n2946), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U5067 ( .A1(n4078), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U5068 ( .A1(n4079), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3996) );
  NAND4_X1 U5069 ( .A1(n3999), .A2(n3998), .A3(n3997), .A4(n3996), .ZN(n4000)
         );
  OR2_X1 U5070 ( .A1(n4001), .A2(n4000), .ZN(n4007) );
  NAND2_X1 U5071 ( .A1(n4008), .A2(n4007), .ZN(n4038) );
  XNOR2_X1 U5072 ( .A(n4039), .B(n4038), .ZN(n4005) );
  NAND2_X1 U5073 ( .A1(n6768), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4002)
         );
  NAND2_X1 U5074 ( .A1(n5412), .A2(n4002), .ZN(n4003) );
  AOI21_X1 U5075 ( .B1(n5280), .B2(EAX_REG_27__SCAN_IN), .A(n4003), .ZN(n4004)
         );
  OAI21_X1 U5076 ( .B1(n4005), .B2(n4066), .A(n4004), .ZN(n4006) );
  OAI21_X1 U5077 ( .B1(n5210), .B2(n5412), .A(n4006), .ZN(n5196) );
  XNOR2_X1 U5078 ( .A(n4008), .B(n4007), .ZN(n4012) );
  NAND2_X1 U5079 ( .A1(n6768), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4009)
         );
  NAND2_X1 U5080 ( .A1(n5412), .A2(n4009), .ZN(n4010) );
  AOI21_X1 U5081 ( .B1(n5280), .B2(EAX_REG_26__SCAN_IN), .A(n4010), .ZN(n4011)
         );
  OAI21_X1 U5082 ( .B1(n4012), .B2(n4066), .A(n4011), .ZN(n4014) );
  XNOR2_X1 U5083 ( .A(n4018), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5693)
         );
  NAND2_X1 U5084 ( .A1(n5693), .A2(n3063), .ZN(n4013) );
  NAND2_X1 U5085 ( .A1(n4014), .A2(n4013), .ZN(n5346) );
  NOR2_X1 U5086 ( .A1(n5196), .A2(n5346), .ZN(n4026) );
  NAND2_X1 U5087 ( .A1(n4016), .A2(n4015), .ZN(n4017) );
  NAND2_X1 U5088 ( .A1(n4018), .A2(n4017), .ZN(n5700) );
  XNOR2_X1 U5089 ( .A(n4020), .B(n4019), .ZN(n4024) );
  NAND2_X1 U5090 ( .A1(n6768), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4021)
         );
  NAND2_X1 U5091 ( .A1(n5412), .A2(n4021), .ZN(n4022) );
  AOI21_X1 U5092 ( .B1(n5280), .B2(EAX_REG_25__SCAN_IN), .A(n4022), .ZN(n4023)
         );
  OAI21_X1 U5093 ( .B1(n4024), .B2(n4066), .A(n4023), .ZN(n4025) );
  OAI21_X1 U5094 ( .B1(n5700), .B2(n5412), .A(n4025), .ZN(n5193) );
  INV_X1 U5095 ( .A(n5193), .ZN(n5357) );
  AND2_X1 U5096 ( .A1(n4026), .A2(n5357), .ZN(n4301) );
  AOI22_X1 U5097 ( .A1(n4051), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U5098 ( .A1(n2971), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n2946), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U5099 ( .A1(n4027), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U5100 ( .A1(n4079), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4028) );
  NAND4_X1 U5101 ( .A1(n4031), .A2(n4030), .A3(n4029), .A4(n4028), .ZN(n4037)
         );
  AOI22_X1 U5102 ( .A1(n2970), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U5103 ( .A1(n4069), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4034) );
  AOI22_X1 U5104 ( .A1(n4057), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U5105 ( .A1(n4072), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4032) );
  NAND4_X1 U5106 ( .A1(n4035), .A2(n4034), .A3(n4033), .A4(n4032), .ZN(n4036)
         );
  OR2_X1 U5107 ( .A1(n4037), .A2(n4036), .ZN(n4049) );
  NOR2_X1 U5108 ( .A1(n4039), .A2(n4038), .ZN(n4050) );
  XOR2_X1 U5109 ( .A(n4049), .B(n4050), .Z(n4040) );
  NAND2_X1 U5110 ( .A1(n4040), .A2(n4095), .ZN(n4043) );
  INV_X1 U5111 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5334) );
  NOR2_X1 U5112 ( .A1(n5334), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4041) );
  AOI211_X1 U5113 ( .C1(n5280), .C2(EAX_REG_28__SCAN_IN), .A(n3063), .B(n4041), 
        .ZN(n4042) );
  XNOR2_X1 U5114 ( .A(n4045), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5336)
         );
  AOI22_X1 U5115 ( .A1(n4043), .A2(n4042), .B1(n3063), .B2(n5336), .ZN(n4302)
         );
  AND2_X1 U5116 ( .A1(n4301), .A2(n4302), .ZN(n4044) );
  INV_X1 U5117 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4046) );
  NAND2_X1 U5118 ( .A1(n4047), .A2(n4046), .ZN(n4048) );
  NAND2_X1 U5119 ( .A1(n5157), .A2(n4048), .ZN(n5685) );
  NAND2_X1 U5120 ( .A1(n4050), .A2(n4049), .ZN(n4086) );
  AOI22_X1 U5121 ( .A1(n4078), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n2971), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U5122 ( .A1(n4051), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n2970), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4055) );
  AOI22_X1 U5123 ( .A1(n4052), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4054) );
  AOI22_X1 U5124 ( .A1(n4072), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4053) );
  NAND4_X1 U5125 ( .A1(n4056), .A2(n4055), .A3(n4054), .A4(n4053), .ZN(n4063)
         );
  AOI22_X1 U5126 ( .A1(n4069), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U5127 ( .A1(n2946), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U5128 ( .A1(n4057), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U5129 ( .A1(n4079), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4058) );
  NAND4_X1 U5130 ( .A1(n4061), .A2(n4060), .A3(n4059), .A4(n4058), .ZN(n4062)
         );
  NOR2_X1 U5131 ( .A1(n4063), .A2(n4062), .ZN(n4087) );
  XNOR2_X1 U5132 ( .A(n4086), .B(n4087), .ZN(n4067) );
  OAI21_X1 U5133 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6297), .A(n6768), 
        .ZN(n4065) );
  NAND2_X1 U5134 ( .A1(n5280), .A2(EAX_REG_29__SCAN_IN), .ZN(n4064) );
  OAI211_X1 U5135 ( .C1(n4067), .C2(n4066), .A(n4065), .B(n4064), .ZN(n4068)
         );
  OAI21_X1 U5136 ( .B1(n5685), .B2(n5412), .A(n4068), .ZN(n5326) );
  XNOR2_X1 U5137 ( .A(n5157), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5315)
         );
  AOI22_X1 U5138 ( .A1(n2970), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4052), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U5139 ( .A1(n4069), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3328), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4075) );
  AOI22_X1 U5140 ( .A1(n4057), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4074) );
  AOI22_X1 U5141 ( .A1(n4072), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4071), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4073) );
  NAND4_X1 U5142 ( .A1(n4076), .A2(n4075), .A3(n4074), .A4(n4073), .ZN(n4085)
         );
  AOI22_X1 U5143 ( .A1(n4051), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4551), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U5144 ( .A1(n2971), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n2946), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4082) );
  AOI22_X1 U5145 ( .A1(n4078), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4081) );
  AOI22_X1 U5146 ( .A1(n4079), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3978), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4080) );
  NAND4_X1 U5147 ( .A1(n4083), .A2(n4082), .A3(n4081), .A4(n4080), .ZN(n4084)
         );
  OR2_X1 U5148 ( .A1(n4085), .A2(n4084), .ZN(n4089) );
  OR2_X1 U5149 ( .A1(n4087), .A2(n4086), .ZN(n4088) );
  XNOR2_X1 U5150 ( .A(n4089), .B(n4088), .ZN(n4094) );
  INV_X1 U5151 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4091) );
  NAND2_X1 U5152 ( .A1(n6768), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4090)
         );
  OAI211_X1 U5153 ( .C1(n4092), .C2(n4091), .A(n4090), .B(n5412), .ZN(n4093)
         );
  AOI21_X1 U5154 ( .B1(n4095), .B2(n4094), .A(n4093), .ZN(n4096) );
  AOI21_X1 U5155 ( .B1(n5315), .B2(n5410), .A(n4096), .ZN(n5281) );
  NAND2_X1 U5156 ( .A1(n6573), .A2(REIP_REG_30__SCAN_IN), .ZN(n5233) );
  OAI21_X1 U5157 ( .B1(n5762), .B2(n5156), .A(n5233), .ZN(n4097) );
  AOI21_X1 U5158 ( .B1(n5764), .B2(n5315), .A(n4097), .ZN(n4098) );
  OAI21_X1 U5159 ( .B1(n5239), .B2(n6298), .A(n4100), .ZN(U2956) );
  INV_X1 U5160 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4291) );
  INV_X1 U5161 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5255) );
  NAND3_X1 U5162 ( .A1(n4101), .A2(n4291), .A3(n5255), .ZN(n4104) );
  NAND3_X1 U5163 ( .A1(n4102), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4103) );
  OAI21_X1 U5164 ( .B1(n5697), .B2(n4104), .A(n4103), .ZN(n4105) );
  XNOR2_X1 U5165 ( .A(n4105), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5682)
         );
  INV_X1 U5166 ( .A(n5159), .ZN(n5102) );
  AND3_X1 U5167 ( .A1(n4109), .A2(n4108), .A3(n4107), .ZN(n4110) );
  OR2_X1 U5168 ( .A1(n4111), .A2(n4110), .ZN(n4113) );
  INV_X1 U5169 ( .A(n4715), .ZN(n4114) );
  AOI21_X1 U5170 ( .B1(n4620), .B2(n5102), .A(n4114), .ZN(n4120) );
  OAI21_X1 U5171 ( .B1(n4620), .B2(n5159), .A(n6824), .ZN(n4427) );
  INV_X1 U5172 ( .A(n4726), .ZN(n4247) );
  OAI211_X1 U5173 ( .C1(n4116), .C2(n4427), .A(n3249), .B(n4247), .ZN(n4117)
         );
  INV_X1 U5174 ( .A(n4117), .ZN(n4118) );
  NOR2_X1 U5175 ( .A1(n4445), .A2(n4118), .ZN(n4119) );
  MUX2_X1 U5176 ( .A(n4120), .B(n4119), .S(n3246), .Z(n4131) );
  NOR2_X1 U5177 ( .A1(n5103), .A2(n4121), .ZN(n4122) );
  NAND2_X1 U5178 ( .A1(n4445), .A2(n4122), .ZN(n4130) );
  INV_X1 U5179 ( .A(n4123), .ZN(n4124) );
  OR2_X1 U5180 ( .A1(n4125), .A2(n4124), .ZN(n4127) );
  NAND2_X1 U5181 ( .A1(n4127), .A2(n4126), .ZN(n4252) );
  NOR2_X1 U5182 ( .A1(n4133), .A2(n4252), .ZN(n4266) );
  NOR2_X1 U5183 ( .A1(n2959), .A2(n3249), .ZN(n4128) );
  OR2_X1 U5184 ( .A1(n4266), .A2(n4407), .ZN(n4129) );
  NAND2_X1 U5185 ( .A1(n4130), .A2(n4129), .ZN(n4432) );
  INV_X1 U5186 ( .A(n4720), .ZN(n4536) );
  OAI22_X1 U5187 ( .A1(n4116), .A2(n4141), .B1(n4134), .B2(n3245), .ZN(n4135)
         );
  INV_X1 U5188 ( .A(n4135), .ZN(n4138) );
  NAND4_X1 U5189 ( .A1(n4536), .A2(n4138), .A3(n4137), .A4(n5121), .ZN(n4139)
         );
  AND2_X1 U5190 ( .A1(n4141), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4140)
         );
  AOI21_X1 U5191 ( .B1(n4423), .B2(EBX_REG_30__SCAN_IN), .A(n4140), .ZN(n5227)
         );
  INV_X1 U5192 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4142) );
  INV_X1 U5193 ( .A(EBX_REG_0__SCAN_IN), .ZN(n6754) );
  NAND2_X1 U5194 ( .A1(n4145), .A2(n6754), .ZN(n4146) );
  OAI21_X1 U5195 ( .B1(n4236), .B2(n6754), .A(n4146), .ZN(n4422) );
  XNOR2_X1 U5196 ( .A(n4147), .B(n4422), .ZN(n4455) );
  NAND2_X1 U5197 ( .A1(n4455), .A2(n4209), .ZN(n4148) );
  NAND2_X1 U5198 ( .A1(n4148), .A2(n4147), .ZN(n4587) );
  MUX2_X1 U5199 ( .A(n4231), .B(n4145), .S(EBX_REG_3__SCAN_IN), .Z(n4149) );
  OAI21_X1 U5200 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n4423), .A(n4149), 
        .ZN(n4837) );
  INV_X1 U5201 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4150) );
  NAND2_X1 U5202 ( .A1(n4152), .A2(n4151), .ZN(n4155) );
  NAND2_X1 U5203 ( .A1(n4236), .A2(n2947), .ZN(n4200) );
  NAND2_X1 U5204 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n2947), .ZN(n4153)
         );
  NAND2_X1 U5205 ( .A1(n4200), .A2(n4153), .ZN(n4154) );
  NOR2_X1 U5206 ( .A1(n4155), .A2(n4154), .ZN(n4588) );
  MUX2_X1 U5207 ( .A(n4231), .B(n4145), .S(EBX_REG_5__SCAN_IN), .Z(n4156) );
  OAI21_X1 U5208 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4423), .A(n4156), 
        .ZN(n4157) );
  INV_X1 U5209 ( .A(n4157), .ZN(n4824) );
  INV_X1 U5210 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6839) );
  NAND2_X1 U5211 ( .A1(n4209), .A2(n6839), .ZN(n4159) );
  OAI211_X1 U5212 ( .C1(n4236), .C2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4145), 
        .B(n4159), .ZN(n4161) );
  NAND2_X1 U5213 ( .A1(n4239), .A2(n6839), .ZN(n4160) );
  NAND2_X1 U5214 ( .A1(n4161), .A2(n4160), .ZN(n4825) );
  NAND2_X1 U5215 ( .A1(n4824), .A2(n4825), .ZN(n4162) );
  INV_X1 U5216 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U5217 ( .A1(n4209), .A2(n5531), .ZN(n4163) );
  OAI211_X1 U5218 ( .C1(n4236), .C2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n4145), 
        .B(n4163), .ZN(n4165) );
  NAND2_X1 U5219 ( .A1(n4239), .A2(n5531), .ZN(n4164) );
  NAND2_X1 U5220 ( .A1(n4165), .A2(n4164), .ZN(n4894) );
  MUX2_X1 U5221 ( .A(n4231), .B(n4145), .S(EBX_REG_7__SCAN_IN), .Z(n4166) );
  OAI21_X1 U5222 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n4423), .A(n4166), 
        .ZN(n5047) );
  INV_X1 U5223 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5523) );
  NAND2_X1 U5224 ( .A1(n4209), .A2(n5523), .ZN(n4167) );
  OAI211_X1 U5225 ( .C1(n4236), .C2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n4145), 
        .B(n4167), .ZN(n4169) );
  NAND2_X1 U5226 ( .A1(n4239), .A2(n5523), .ZN(n4168) );
  AND2_X1 U5227 ( .A1(n4169), .A2(n4168), .ZN(n5135) );
  INV_X1 U5228 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6818) );
  NAND2_X1 U5229 ( .A1(n4209), .A2(n6818), .ZN(n4170) );
  OAI211_X1 U5230 ( .C1(n5439), .C2(n5807), .A(n4224), .B(n4170), .ZN(n4172)
         );
  NAND2_X1 U5231 ( .A1(n4225), .A2(n6818), .ZN(n4171) );
  INV_X1 U5232 ( .A(n4239), .ZN(n4215) );
  MUX2_X1 U5233 ( .A(n4215), .B(n4224), .S(EBX_REG_10__SCAN_IN), .Z(n4175) );
  NAND2_X1 U5234 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n4141), .ZN(n4173) );
  AND2_X1 U5235 ( .A1(n4200), .A2(n4173), .ZN(n4174) );
  NAND2_X1 U5236 ( .A1(n4175), .A2(n4174), .ZN(n5621) );
  NAND2_X1 U5237 ( .A1(n5514), .A2(n5621), .ZN(n5623) );
  INV_X1 U5238 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5615) );
  NAND2_X1 U5239 ( .A1(n4209), .A2(n5615), .ZN(n4177) );
  NAND2_X1 U5240 ( .A1(n4145), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4176) );
  NAND3_X1 U5241 ( .A1(n4224), .A2(n4177), .A3(n4176), .ZN(n4179) );
  NAND2_X1 U5242 ( .A1(n4225), .A2(n5615), .ZN(n4178) );
  NAND2_X1 U5243 ( .A1(n4179), .A2(n4178), .ZN(n5502) );
  MUX2_X1 U5244 ( .A(n4239), .B(n4236), .S(EBX_REG_12__SCAN_IN), .Z(n4182) );
  NAND2_X1 U5245 ( .A1(n4141), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4180) );
  NAND2_X1 U5246 ( .A1(n4200), .A2(n4180), .ZN(n4181) );
  NOR2_X1 U5247 ( .A1(n4182), .A2(n4181), .ZN(n5612) );
  NAND2_X1 U5248 ( .A1(n4209), .A2(n6794), .ZN(n4184) );
  NAND2_X1 U5249 ( .A1(n4145), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4183) );
  NAND3_X1 U5250 ( .A1(n4224), .A2(n4184), .A3(n4183), .ZN(n4186) );
  NAND2_X1 U5251 ( .A1(n4225), .A2(n6794), .ZN(n4185) );
  INV_X1 U5252 ( .A(EBX_REG_19__SCAN_IN), .ZN(n4188) );
  NAND2_X1 U5253 ( .A1(n4209), .A2(n4188), .ZN(n4187) );
  OAI211_X1 U5254 ( .C1(n4236), .C2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n4145), .B(n4187), .ZN(n4190) );
  NAND2_X1 U5255 ( .A1(n4239), .A2(n4188), .ZN(n4189) );
  NAND2_X1 U5256 ( .A1(n4190), .A2(n4189), .ZN(n5443) );
  INV_X1 U5257 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6793) );
  NAND2_X1 U5258 ( .A1(n4209), .A2(n6793), .ZN(n4192) );
  NAND2_X1 U5259 ( .A1(n4145), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4191) );
  NAND3_X1 U5260 ( .A1(n4224), .A2(n4192), .A3(n4191), .ZN(n4194) );
  NAND2_X1 U5261 ( .A1(n4225), .A2(n6793), .ZN(n4193) );
  NAND2_X1 U5262 ( .A1(n4194), .A2(n4193), .ZN(n5487) );
  INV_X1 U5263 ( .A(n5487), .ZN(n4198) );
  MUX2_X1 U5264 ( .A(n4215), .B(n4224), .S(EBX_REG_14__SCAN_IN), .Z(n4197) );
  NAND2_X1 U5265 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n4141), .ZN(n4195) );
  AND2_X1 U5266 ( .A1(n4200), .A2(n4195), .ZN(n4196) );
  NAND2_X1 U5267 ( .A1(n4197), .A2(n4196), .ZN(n5166) );
  MUX2_X1 U5268 ( .A(n4215), .B(n4224), .S(EBX_REG_16__SCAN_IN), .Z(n4202) );
  NAND2_X1 U5269 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n4141), .ZN(n4199) );
  AND2_X1 U5270 ( .A1(n4200), .A2(n4199), .ZN(n4201) );
  NAND2_X1 U5271 ( .A1(n4202), .A2(n4201), .ZN(n5595) );
  NAND2_X1 U5272 ( .A1(n4145), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4203) );
  OAI211_X1 U5273 ( .C1(EBX_REG_17__SCAN_IN), .C2(n4141), .A(n4224), .B(n4203), 
        .ZN(n4206) );
  INV_X1 U5274 ( .A(EBX_REG_17__SCAN_IN), .ZN(n4204) );
  NAND2_X1 U5275 ( .A1(n4225), .A2(n4204), .ZN(n4205) );
  AND2_X1 U5276 ( .A1(n4206), .A2(n4205), .ZN(n5470) );
  AND2_X1 U5277 ( .A1(n5595), .A2(n5470), .ZN(n4207) );
  NAND2_X1 U5278 ( .A1(n5165), .A2(n4208), .ZN(n5425) );
  INV_X1 U5279 ( .A(n4423), .ZN(n4232) );
  NOR2_X1 U5280 ( .A1(n4141), .A2(EBX_REG_20__SCAN_IN), .ZN(n4210) );
  AOI21_X1 U5281 ( .B1(n4232), .B2(n6838), .A(n4210), .ZN(n5426) );
  INV_X1 U5282 ( .A(EBX_REG_18__SCAN_IN), .ZN(n4211) );
  NAND2_X1 U5283 ( .A1(n4209), .A2(n4211), .ZN(n5440) );
  OAI21_X1 U5284 ( .B1(n4423), .B2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n5440), 
        .ZN(n5441) );
  INV_X1 U5285 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5587) );
  OAI22_X1 U5286 ( .A1(n5426), .A2(n5441), .B1(n4145), .B2(n5587), .ZN(n4213)
         );
  AND2_X1 U5287 ( .A1(n5441), .A2(n4145), .ZN(n4212) );
  MUX2_X1 U5288 ( .A(n4231), .B(n4145), .S(EBX_REG_21__SCAN_IN), .Z(n4214) );
  OAI21_X1 U5289 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n4423), .A(n4214), 
        .ZN(n5417) );
  MUX2_X1 U5290 ( .A(n4215), .B(n4224), .S(EBX_REG_22__SCAN_IN), .Z(n4217) );
  NAND2_X1 U5291 ( .A1(n4141), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4216) );
  NAND2_X1 U5292 ( .A1(n4217), .A2(n4216), .ZN(n4353) );
  NAND2_X1 U5293 ( .A1(n4145), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4218) );
  OAI211_X1 U5294 ( .C1(EBX_REG_23__SCAN_IN), .C2(n4141), .A(n4224), .B(n4218), 
        .ZN(n4220) );
  INV_X1 U5295 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U5296 ( .A1(n4225), .A2(n5582), .ZN(n4219) );
  MUX2_X1 U5297 ( .A(n4239), .B(n4236), .S(EBX_REG_24__SCAN_IN), .Z(n4222) );
  AND2_X1 U5298 ( .A1(n4141), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4221)
         );
  NOR2_X1 U5299 ( .A1(n4222), .A2(n4221), .ZN(n5377) );
  NAND2_X1 U5300 ( .A1(n4145), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4223) );
  OAI211_X1 U5301 ( .C1(EBX_REG_25__SCAN_IN), .C2(n4141), .A(n4224), .B(n4223), 
        .ZN(n4227) );
  INV_X1 U5302 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U5303 ( .A1(n4225), .A2(n5579), .ZN(n4226) );
  NAND2_X1 U5304 ( .A1(n4227), .A2(n4226), .ZN(n5362) );
  INV_X1 U5305 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U5306 ( .A1(n4209), .A2(n5578), .ZN(n4228) );
  OAI211_X1 U5307 ( .C1(n4236), .C2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n4145), .B(n4228), .ZN(n4230) );
  NAND2_X1 U5308 ( .A1(n4239), .A2(n5578), .ZN(n4229) );
  NAND2_X1 U5309 ( .A1(n4230), .A2(n4229), .ZN(n5344) );
  MUX2_X1 U5310 ( .A(n4231), .B(n4145), .S(EBX_REG_27__SCAN_IN), .Z(n4234) );
  NAND2_X1 U5311 ( .A1(n4232), .A2(n5822), .ZN(n4233) );
  INV_X1 U5312 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U5313 ( .A1(n4209), .A2(n5339), .ZN(n4235) );
  OAI211_X1 U5314 ( .C1(n4236), .C2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n4145), .B(n4235), .ZN(n4238) );
  NAND2_X1 U5315 ( .A1(n4239), .A2(n5339), .ZN(n4237) );
  AND2_X1 U5316 ( .A1(n4238), .A2(n4237), .ZN(n5240) );
  OAI22_X1 U5317 ( .A1(n4423), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        EBX_REG_29__SCAN_IN), .B2(n4141), .ZN(n5262) );
  INV_X1 U5318 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5575) );
  NAND2_X1 U5319 ( .A1(n4239), .A2(n5575), .ZN(n5260) );
  OAI22_X2 U5320 ( .A1(n5228), .A2(n5439), .B1(n5260), .B2(n5261), .ZN(n5259)
         );
  NOR2_X1 U5321 ( .A1(n5226), .A2(n5439), .ZN(n5231) );
  AOI21_X1 U5322 ( .B1(n5227), .B2(n5259), .A(n5231), .ZN(n4241) );
  OAI22_X1 U5323 ( .A1(n4423), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4141), .ZN(n4242) );
  INV_X1 U5324 ( .A(n4242), .ZN(n4243) );
  OR2_X1 U5325 ( .A1(n4134), .A2(n3209), .ZN(n4245) );
  AOI22_X1 U5326 ( .A1(n4248), .A2(n5439), .B1(n4624), .B2(n4247), .ZN(n4250)
         );
  NAND2_X1 U5327 ( .A1(n3234), .A2(n4620), .ZN(n5542) );
  NOR2_X1 U5328 ( .A1(n5542), .A2(n4624), .ZN(n4424) );
  OAI21_X1 U5329 ( .B1(n4424), .B2(n4423), .A(n2961), .ZN(n4249) );
  NAND2_X1 U5330 ( .A1(n4250), .A2(n4249), .ZN(n4251) );
  OR3_X1 U5331 ( .A1(n4253), .A2(n4252), .A3(n4251), .ZN(n4439) );
  INV_X1 U5332 ( .A(n4439), .ZN(n4261) );
  NAND2_X1 U5333 ( .A1(n4255), .A2(n4254), .ZN(n4260) );
  NAND2_X1 U5334 ( .A1(n4256), .A2(n4257), .ZN(n4259) );
  INV_X1 U5335 ( .A(n5103), .ZN(n4442) );
  NAND2_X1 U5336 ( .A1(n4442), .A2(n4258), .ZN(n4555) );
  NAND4_X1 U5337 ( .A1(n4261), .A2(n4260), .A3(n4259), .A4(n4555), .ZN(n4262)
         );
  NAND2_X1 U5338 ( .A1(n5300), .A2(n5921), .ZN(n4517) );
  NAND2_X1 U5339 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5957) );
  NAND2_X1 U5340 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5956) );
  NOR2_X1 U5341 ( .A1(n5957), .A2(n5956), .ZN(n4270) );
  INV_X1 U5342 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6568) );
  NOR2_X1 U5343 ( .A1(n6568), .A2(n4263), .ZN(n6548) );
  INV_X1 U5344 ( .A(n6548), .ZN(n6557) );
  NAND2_X1 U5345 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4269) );
  NAND2_X1 U5346 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4992) );
  NOR3_X1 U5347 ( .A1(n6557), .A2(n4269), .A3(n4992), .ZN(n5959) );
  NAND2_X1 U5348 ( .A1(n4270), .A2(n5959), .ZN(n4280) );
  INV_X1 U5349 ( .A(n4280), .ZN(n4264) );
  NAND2_X1 U5350 ( .A1(n6570), .A2(n4264), .ZN(n5861) );
  NOR2_X1 U5351 ( .A1(n5103), .A2(n4141), .ZN(n4265) );
  NAND2_X1 U5352 ( .A1(n4266), .A2(n4265), .ZN(n4535) );
  INV_X1 U5353 ( .A(n4535), .ZN(n4267) );
  NAND2_X1 U5354 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6571) );
  NAND2_X1 U5355 ( .A1(n6789), .A2(n6571), .ZN(n6555) );
  NAND2_X1 U5356 ( .A1(n6548), .A2(n6555), .ZN(n6542) );
  NOR2_X1 U5357 ( .A1(n6542), .A2(n4269), .ZN(n5961) );
  AND2_X1 U5358 ( .A1(n5961), .A2(n4270), .ZN(n4277) );
  NAND2_X1 U5359 ( .A1(n5938), .A2(n4277), .ZN(n5924) );
  NAND2_X1 U5360 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5937) );
  NOR2_X1 U5361 ( .A1(n5937), .A2(n5929), .ZN(n5922) );
  NAND2_X1 U5362 ( .A1(n5922), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5897) );
  INV_X1 U5363 ( .A(n4271), .ZN(n4272) );
  NOR2_X1 U5364 ( .A1(n5888), .A2(n5889), .ZN(n4273) );
  NAND2_X1 U5365 ( .A1(n5952), .A2(n4273), .ZN(n5881) );
  INV_X1 U5366 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6784) );
  INV_X1 U5367 ( .A(n5863), .ZN(n4274) );
  NOR2_X1 U5368 ( .A1(n5873), .A2(n4274), .ZN(n4348) );
  NAND2_X1 U5369 ( .A1(n4348), .A2(n4349), .ZN(n5846) );
  INV_X1 U5370 ( .A(n5828), .ZN(n4290) );
  NOR2_X1 U5371 ( .A1(n5835), .A2(n4290), .ZN(n5823) );
  NAND3_X1 U5372 ( .A1(n5823), .A2(n5243), .A3(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5235) );
  INV_X1 U5373 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4446) );
  NAND2_X1 U5374 ( .A1(n4446), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4292) );
  NAND2_X1 U5375 ( .A1(n6573), .A2(REIP_REG_31__SCAN_IN), .ZN(n5677) );
  INV_X1 U5376 ( .A(n5964), .ZN(n5896) );
  NAND2_X1 U5377 ( .A1(n4276), .A2(n6524), .ZN(n4515) );
  OAI21_X1 U5378 ( .B1(n5923), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4515), 
        .ZN(n5963) );
  INV_X1 U5379 ( .A(n4277), .ZN(n4278) );
  AND2_X1 U5380 ( .A1(n5938), .A2(n4278), .ZN(n4279) );
  NOR2_X1 U5381 ( .A1(n5963), .A2(n4279), .ZN(n4282) );
  NAND2_X1 U5382 ( .A1(n5958), .A2(n4280), .ZN(n4281) );
  NAND2_X1 U5383 ( .A1(n5863), .A2(n4283), .ZN(n4284) );
  NOR2_X1 U5384 ( .A1(n5888), .A2(n4284), .ZN(n4285) );
  OR2_X1 U5385 ( .A1(n5964), .A2(n4349), .ZN(n4287) );
  NAND2_X1 U5386 ( .A1(n4347), .A2(n4287), .ZN(n4311) );
  INV_X1 U5387 ( .A(n6570), .ZN(n4990) );
  AOI21_X1 U5388 ( .B1(n4990), .B2(n6577), .A(n4288), .ZN(n4289) );
  AOI21_X1 U5389 ( .B1(n4290), .B2(n5896), .A(n5838), .ZN(n5818) );
  OAI211_X1 U5390 ( .C1(n5243), .C2(n5964), .A(n5818), .B(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5254) );
  INV_X1 U5391 ( .A(n5838), .ZN(n5844) );
  NAND2_X1 U5392 ( .A1(n5844), .A2(n5964), .ZN(n5232) );
  AND2_X1 U5393 ( .A1(n5808), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4294)
         );
  NOR2_X1 U5394 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5827) );
  NAND3_X1 U5395 ( .A1(n4295), .A2(n4296), .A3(n5827), .ZN(n5190) );
  INV_X1 U5396 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4297) );
  AND2_X1 U5397 ( .A1(n4297), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4298)
         );
  XNOR2_X1 U5398 ( .A(n4300), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5250)
         );
  NAND2_X1 U5399 ( .A1(n6573), .A2(REIP_REG_28__SCAN_IN), .ZN(n5245) );
  OAI21_X1 U5400 ( .B1(n5762), .B2(n5334), .A(n5245), .ZN(n4304) );
  OAI21_X1 U5401 ( .B1(n5197), .B2(n4302), .A(n5325), .ZN(n5639) );
  NOR2_X1 U5402 ( .A1(n5639), .A2(n5816), .ZN(n4303) );
  OAI21_X1 U5403 ( .B1(n5250), .B2(n6298), .A(n4305), .ZN(U2958) );
  NOR3_X1 U5404 ( .A1(n4306), .A2(n6838), .A3(n4307), .ZN(n4308) );
  AOI21_X2 U5405 ( .B1(n4332), .B2(n4333), .A(n4308), .ZN(n4309) );
  XNOR2_X2 U5406 ( .A(n4309), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4320)
         );
  NAND2_X1 U5407 ( .A1(n4320), .A2(n6579), .ZN(n4319) );
  INV_X1 U5408 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6781) );
  NOR2_X1 U5409 ( .A1(n6524), .A2(n6781), .ZN(n4325) );
  NOR2_X1 U5410 ( .A1(n5846), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4310)
         );
  AOI211_X1 U5411 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n4311), .A(n4325), .B(n4310), .ZN(n4317) );
  OAI21_X1 U5412 ( .B1(n4312), .B2(n4313), .A(n5376), .ZN(n5581) );
  INV_X1 U5413 ( .A(n5581), .ZN(n4315) );
  NAND2_X1 U5414 ( .A1(n4315), .A2(n4314), .ZN(n4316) );
  NAND2_X1 U5415 ( .A1(n4319), .A2(n4318), .ZN(U2995) );
  NAND2_X1 U5416 ( .A1(n4320), .A2(n6505), .ZN(n4329) );
  AND2_X1 U5417 ( .A1(n4338), .A2(n4322), .ZN(n4323) );
  OR2_X1 U5418 ( .A1(n3953), .A2(n4323), .ZN(n5649) );
  NOR2_X1 U5419 ( .A1(n6510), .A2(n5381), .ZN(n4324) );
  AOI211_X1 U5420 ( .C1(n6501), .C2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n4325), 
        .B(n4324), .ZN(n4326) );
  NAND2_X1 U5421 ( .A1(n4329), .A2(n4328), .ZN(U2963) );
  INV_X1 U5422 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4330) );
  NOR2_X1 U5423 ( .A1(n4332), .A2(n4331), .ZN(n4335) );
  AOI21_X1 U5424 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5808), .A(n4333), 
        .ZN(n4334) );
  XNOR2_X1 U5425 ( .A(n4335), .B(n4334), .ZN(n4346) );
  NAND2_X1 U5426 ( .A1(n4346), .A2(n6505), .ZN(n4345) );
  INV_X1 U5427 ( .A(n4336), .ZN(n5414) );
  INV_X1 U5428 ( .A(n4337), .ZN(n4339) );
  OAI21_X1 U5429 ( .B1(n5414), .B2(n4339), .A(n4338), .ZN(n5652) );
  INV_X1 U5430 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6704) );
  NOR2_X1 U5431 ( .A1(n6524), .A2(n6704), .ZN(n4352) );
  NOR2_X1 U5432 ( .A1(n5762), .A2(n4340), .ZN(n4341) );
  AOI211_X1 U5433 ( .C1(n5764), .C2(n5391), .A(n4352), .B(n4341), .ZN(n4342)
         );
  NAND2_X1 U5434 ( .A1(n4345), .A2(n4344), .ZN(U2964) );
  NAND2_X1 U5435 ( .A1(n4346), .A2(n6579), .ZN(n4358) );
  INV_X1 U5436 ( .A(n4347), .ZN(n5854) );
  INV_X1 U5437 ( .A(n4348), .ZN(n5856) );
  NOR3_X1 U5438 ( .A1(n5856), .A2(n4350), .A3(n4349), .ZN(n4351) );
  AOI211_X1 U5439 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5854), .A(n4352), .B(n4351), .ZN(n4356) );
  NOR2_X1 U5440 ( .A1(n2989), .A2(n4353), .ZN(n4354) );
  OR2_X1 U5441 ( .A1(n5583), .A2(n5966), .ZN(n4355) );
  NAND2_X1 U5442 ( .A1(n4358), .A2(n4357), .ZN(U2996) );
  INV_X1 U5443 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n4371) );
  NOR2_X1 U5444 ( .A1(n6710), .A2(n4371), .ZN(n4365) );
  AND2_X1 U5445 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n4372) );
  NAND2_X1 U5446 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n4359) );
  OAI21_X1 U5447 ( .B1(n4365), .B2(n4372), .A(n4359), .ZN(n4360) );
  OAI211_X1 U5448 ( .C1(n4378), .C2(n6824), .A(n4360), .B(n5102), .ZN(U3182)
         );
  AOI221_X1 U5449 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6824), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n4361) );
  AOI221_X1 U5450 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n4361), .C2(HOLD), .A(n6710), .ZN(n4368) );
  AND2_X1 U5451 ( .A1(n4364), .A2(n6710), .ZN(n4363) );
  INV_X1 U5452 ( .A(NA_N), .ZN(n4366) );
  NAND2_X1 U5453 ( .A1(n4366), .A2(STATE_REG_2__SCAN_IN), .ZN(n4362) );
  AND2_X1 U5454 ( .A1(n4363), .A2(n4362), .ZN(n4373) );
  AOI22_X1 U5455 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n4377) );
  INV_X1 U5456 ( .A(n4364), .ZN(n4376) );
  AOI21_X1 U5457 ( .B1(n4366), .B2(n4365), .A(n4376), .ZN(n4367) );
  OAI22_X1 U5458 ( .A1(n4368), .A2(n4373), .B1(n4377), .B2(n4367), .ZN(U3183)
         );
  NAND2_X1 U5459 ( .A1(n6824), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6645) );
  NAND2_X1 U5460 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4573), .ZN(n5131) );
  INV_X1 U5461 ( .A(n5131), .ZN(n4568) );
  AOI211_X1 U5462 ( .C1(n6768), .C2(n6645), .A(n4568), .B(n6697), .ZN(n4370)
         );
  OR2_X1 U5463 ( .A1(n4370), .A2(n4369), .ZN(U3150) );
  OAI21_X1 U5464 ( .B1(n4372), .B2(n4371), .A(n6855), .ZN(n4375) );
  INV_X1 U5465 ( .A(n4373), .ZN(n4374) );
  OAI211_X1 U5466 ( .C1(n4377), .C2(n4376), .A(n4375), .B(n4374), .ZN(U3181)
         );
  INV_X1 U5467 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6734) );
  OAI21_X1 U5468 ( .B1(n4378), .B2(STATE_REG_2__SCAN_IN), .A(
        STATE_REG_0__SCAN_IN), .ZN(n4379) );
  OAI21_X1 U5469 ( .B1(n6702), .B2(n6734), .A(n6677), .ZN(U2789) );
  INV_X1 U5470 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5490) );
  NOR2_X2 U5471 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6855), .ZN(n6856) );
  AOI22_X1 U5472 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6856), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6855), .ZN(n4380) );
  OAI21_X1 U5473 ( .B1(n5490), .B2(n6653), .A(n4380), .ZN(U3198) );
  INV_X1 U5474 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6525) );
  AOI22_X1 U5475 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6856), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6855), .ZN(n4381) );
  OAI21_X1 U5476 ( .B1(n6525), .B2(n6653), .A(n4381), .ZN(U3191) );
  AOI22_X1 U5477 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6856), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6855), .ZN(n4382) );
  OAI21_X1 U5478 ( .B1(n6799), .B2(n6653), .A(n4382), .ZN(U3209) );
  AOI22_X1 U5479 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6856), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6855), .ZN(n4383) );
  OAI21_X1 U5480 ( .B1(n5810), .B2(n6653), .A(n4383), .ZN(U3192) );
  INV_X1 U5481 ( .A(REIP_REG_10__SCAN_IN), .ZN(n5965) );
  AOI22_X1 U5482 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6856), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6855), .ZN(n4384) );
  OAI21_X1 U5483 ( .B1(n5965), .B2(n6653), .A(n4384), .ZN(U3193) );
  AOI22_X1 U5484 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6856), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6855), .ZN(n4385) );
  OAI21_X1 U5485 ( .B1(n6661), .B2(n6653), .A(n4385), .ZN(U3190) );
  AOI22_X1 U5486 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6856), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6855), .ZN(n4386) );
  OAI21_X1 U5487 ( .B1(n5220), .B2(n6653), .A(n4386), .ZN(U3210) );
  INV_X1 U5488 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6670) );
  AOI22_X1 U5489 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6856), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6855), .ZN(n4387) );
  OAI21_X1 U5490 ( .B1(n6670), .B2(n6653), .A(n4387), .ZN(U3204) );
  INV_X1 U5491 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6657) );
  AOI22_X1 U5492 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6856), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6855), .ZN(n4388) );
  OAI21_X1 U5493 ( .B1(n6657), .B2(n6653), .A(n4388), .ZN(U3187) );
  INV_X1 U5494 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6800) );
  AOI22_X1 U5495 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6856), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6855), .ZN(n4389) );
  OAI21_X1 U5496 ( .B1(n6800), .B2(n6653), .A(n4389), .ZN(U3207) );
  INV_X1 U5497 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6655) );
  AOI22_X1 U5498 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6856), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6855), .ZN(n4390) );
  OAI21_X1 U5499 ( .B1(n6655), .B2(n6653), .A(n4390), .ZN(U3185) );
  INV_X1 U5500 ( .A(REIP_REG_17__SCAN_IN), .ZN(n4395) );
  AOI22_X1 U5501 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6856), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6855), .ZN(n4391) );
  OAI21_X1 U5502 ( .B1(n4395), .B2(n6653), .A(n4391), .ZN(U3200) );
  INV_X1 U5503 ( .A(REIP_REG_29__SCAN_IN), .ZN(n5285) );
  AOI22_X1 U5504 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6856), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6855), .ZN(n4392) );
  OAI21_X1 U5505 ( .B1(n5285), .B2(n6653), .A(n4392), .ZN(U3212) );
  INV_X1 U5506 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6665) );
  AOI22_X1 U5507 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6856), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6855), .ZN(n4393) );
  OAI21_X1 U5508 ( .B1(n6665), .B2(n6653), .A(n4393), .ZN(U3196) );
  INV_X1 U5509 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6767) );
  AOI22_X1 U5510 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6856), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6855), .ZN(n4394) );
  OAI21_X1 U5511 ( .B1(n6767), .B2(n6653), .A(n4394), .ZN(U3197) );
  INV_X1 U5512 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5759) );
  INV_X1 U5513 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n6723) );
  INV_X1 U5514 ( .A(n6856), .ZN(n6674) );
  OAI222_X1 U5515 ( .A1(n6653), .A2(n5759), .B1(n6702), .B2(n6723), .C1(n4395), 
        .C2(n6674), .ZN(U3199) );
  INV_X1 U5516 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6834) );
  OAI222_X1 U5517 ( .A1(n6653), .A2(n6704), .B1(n6702), .B2(n6834), .C1(n6781), 
        .C2(n6674), .ZN(U3205) );
  INV_X1 U5518 ( .A(n4717), .ZN(n5548) );
  INV_X1 U5519 ( .A(n4457), .ZN(n4398) );
  INV_X1 U5520 ( .A(n4406), .ZN(n4397) );
  OAI22_X1 U5521 ( .A1(n3081), .A2(n5548), .B1(n4398), .B2(n4401), .ZN(n4403)
         );
  OAI21_X1 U5522 ( .B1(n4403), .B2(n6644), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n4400) );
  NAND3_X1 U5523 ( .A1(n5306), .A2(STATE2_REG_0__SCAN_IN), .A3(n6768), .ZN(
        n4399) );
  NAND2_X1 U5524 ( .A1(n4400), .A2(n4399), .ZN(U2790) );
  NOR2_X1 U5525 ( .A1(n6691), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5310) );
  AOI21_X1 U5526 ( .B1(n5149), .B2(MEMORYFETCH_REG_SCAN_IN), .A(n5310), .ZN(
        n4402) );
  NAND2_X1 U5527 ( .A1(n5150), .A2(n4402), .ZN(U2788) );
  NAND2_X1 U5528 ( .A1(n3411), .A2(n5542), .ZN(n5311) );
  AOI21_X1 U5529 ( .B1(n5311), .B2(n5102), .A(READY_N), .ZN(n6696) );
  NOR2_X1 U5530 ( .A1(n4403), .A2(n6696), .ZN(n5120) );
  NOR2_X1 U5531 ( .A1(n5120), .A2(n6644), .ZN(n6300) );
  INV_X1 U5532 ( .A(MORE_REG_SCAN_IN), .ZN(n4411) );
  NAND2_X1 U5533 ( .A1(n5121), .A2(n4457), .ZN(n4404) );
  NOR2_X1 U5534 ( .A1(n4720), .A2(n4404), .ZN(n4405) );
  MUX2_X1 U5535 ( .A(n4535), .B(n4405), .S(n4445), .Z(n4409) );
  NAND2_X1 U5536 ( .A1(n4407), .A2(n4406), .ZN(n4408) );
  NAND2_X1 U5537 ( .A1(n4409), .A2(n4408), .ZN(n5124) );
  NAND2_X1 U5538 ( .A1(n6300), .A2(n5124), .ZN(n4410) );
  OAI21_X1 U5539 ( .B1(n6300), .B2(n4411), .A(n4410), .ZN(U3471) );
  OAI21_X1 U5540 ( .B1(n4414), .B2(n4413), .A(n4412), .ZN(n5571) );
  NOR2_X1 U5541 ( .A1(n4535), .A2(n6644), .ZN(n4415) );
  NAND2_X1 U5542 ( .A1(n4445), .A2(n4415), .ZN(n4421) );
  AND2_X1 U5543 ( .A1(n2945), .A2(n4631), .ZN(n4417) );
  AND3_X1 U5544 ( .A1(n3246), .A2(n3215), .A3(n5301), .ZN(n4416) );
  NAND4_X1 U5545 ( .A1(n5280), .A2(n4418), .A3(n4417), .A4(n4416), .ZN(n4716)
         );
  INV_X1 U5546 ( .A(n4716), .ZN(n4419) );
  NAND2_X2 U5547 ( .A1(n5626), .A2(n4724), .ZN(n5630) );
  OAI21_X1 U5548 ( .B1(n4423), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4422), 
        .ZN(n5565) );
  OAI222_X1 U5549 ( .A1(n5571), .A2(n5630), .B1(n5626), .B2(n6754), .C1(n5565), 
        .C2(n5624), .ZN(U2859) );
  INV_X1 U5550 ( .A(n4137), .ZN(n4425) );
  AOI21_X1 U5551 ( .B1(n4425), .B2(n4715), .A(n4424), .ZN(n4426) );
  OAI21_X1 U5552 ( .B1(n4445), .B2(n4536), .A(n4426), .ZN(n4431) );
  AOI21_X1 U5553 ( .B1(n4457), .B2(n5102), .A(n4427), .ZN(n4428) );
  OAI21_X1 U5554 ( .B1(n5270), .B2(n3230), .A(n4428), .ZN(n4429) );
  NOR2_X1 U5555 ( .A1(n4445), .A2(n4429), .ZN(n4430) );
  NAND2_X1 U5556 ( .A1(n4561), .A2(n3080), .ZN(n6291) );
  NAND2_X1 U5557 ( .A1(n4568), .A2(FLUSH_REG_SCAN_IN), .ZN(n4433) );
  OAI211_X1 U5558 ( .C1(STATE2_REG_0__SCAN_IN), .C2(n6103), .A(n6291), .B(
        n4433), .ZN(n6294) );
  INV_X1 U5559 ( .A(n4256), .ZN(n4436) );
  NAND4_X1 U5560 ( .A1(n4437), .A2(n4137), .A3(n4436), .A4(n4116), .ZN(n4438)
         );
  NOR2_X1 U5561 ( .A1(n4439), .A2(n4438), .ZN(n5104) );
  INV_X1 U5562 ( .A(n5104), .ZN(n4546) );
  OAI21_X1 U5563 ( .B1(n4440), .B2(n4441), .A(n4442), .ZN(n4443) );
  OAI21_X1 U5564 ( .B1(n4494), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n4443), 
        .ZN(n4444) );
  AOI21_X1 U5565 ( .B1(n6400), .B2(n4546), .A(n4444), .ZN(n5106) );
  INV_X1 U5566 ( .A(n6283), .ZN(n5298) );
  NAND2_X1 U5567 ( .A1(n5298), .A2(n4441), .ZN(n4448) );
  AOI22_X1 U5568 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4446), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4518), .ZN(n5299) );
  NAND3_X1 U5569 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5299), .A3(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4447) );
  OAI211_X1 U5570 ( .C1(n5106), .C2(n6646), .A(n4448), .B(n4447), .ZN(n4449)
         );
  AOI22_X1 U5571 ( .A1(n4449), .A2(n6294), .B1(n4440), .B2(n5298), .ZN(n4450)
         );
  OAI21_X1 U5572 ( .B1(n3225), .B2(n6294), .A(n4450), .ZN(U3460) );
  OR2_X1 U5573 ( .A1(n4452), .A2(n4451), .ZN(n4453) );
  NAND2_X1 U5574 ( .A1(n4454), .A2(n4453), .ZN(n6405) );
  XNOR2_X1 U5575 ( .A(n4455), .B(n4209), .ZN(n4521) );
  AOI22_X1 U5576 ( .A1(n5628), .A2(n4521), .B1(n5627), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4456) );
  OAI21_X1 U5577 ( .B1(n6405), .B2(n5630), .A(n4456), .ZN(U2858) );
  INV_X1 U5578 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4461) );
  NAND2_X1 U5579 ( .A1(n6471), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4460) );
  NAND2_X1 U5580 ( .A1(n6470), .A2(DATAI_1_), .ZN(n4785) );
  OAI211_X1 U5581 ( .C1(n6473), .C2(n4461), .A(n4460), .B(n4785), .ZN(U2925)
         );
  INV_X1 U5582 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6425) );
  NAND2_X1 U5583 ( .A1(n6471), .A2(LWORD_REG_13__SCAN_IN), .ZN(n4462) );
  INV_X1 U5584 ( .A(DATAI_13_), .ZN(n5669) );
  OR2_X1 U5585 ( .A1(n4723), .A2(n5669), .ZN(n4770) );
  OAI211_X1 U5586 ( .C1(n6473), .C2(n6425), .A(n4462), .B(n4770), .ZN(U2952)
         );
  XNOR2_X1 U5587 ( .A(n4463), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4512)
         );
  INV_X1 U5588 ( .A(n5571), .ZN(n4464) );
  NAND2_X1 U5589 ( .A1(n4464), .A2(n5795), .ZN(n4468) );
  OR2_X1 U5590 ( .A1(n6501), .A2(n4465), .ZN(n4466) );
  AOI22_X1 U5591 ( .A1(n4466), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .B1(n6573), 
        .B2(REIP_REG_0__SCAN_IN), .ZN(n4467) );
  OAI211_X1 U5592 ( .C1(n4512), .C2(n6298), .A(n4468), .B(n4467), .ZN(U2986)
         );
  INV_X1 U5593 ( .A(LWORD_REG_8__SCAN_IN), .ZN(n4470) );
  INV_X1 U5594 ( .A(DATAI_8_), .ZN(n5139) );
  NOR2_X1 U5595 ( .A1(n4723), .A2(n5139), .ZN(n4490) );
  AOI21_X1 U5596 ( .B1(n6467), .B2(EAX_REG_8__SCAN_IN), .A(n4490), .ZN(n4469)
         );
  OAI21_X1 U5597 ( .B1(n4493), .B2(n4470), .A(n4469), .ZN(U2947) );
  INV_X1 U5598 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n4472) );
  INV_X1 U5599 ( .A(DATAI_4_), .ZN(n4787) );
  NOR2_X1 U5600 ( .A1(n4723), .A2(n4787), .ZN(n4479) );
  AOI21_X1 U5601 ( .B1(n6467), .B2(EAX_REG_20__SCAN_IN), .A(n4479), .ZN(n4471)
         );
  OAI21_X1 U5602 ( .B1(n4493), .B2(n4472), .A(n4471), .ZN(U2928) );
  INV_X1 U5603 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n6803) );
  NOR2_X1 U5604 ( .A1(n4723), .A2(n5046), .ZN(n4476) );
  AOI21_X1 U5605 ( .B1(n6467), .B2(EAX_REG_7__SCAN_IN), .A(n4476), .ZN(n4473)
         );
  OAI21_X1 U5606 ( .B1(n4493), .B2(n6803), .A(n4473), .ZN(U2946) );
  INV_X1 U5607 ( .A(UWORD_REG_2__SCAN_IN), .ZN(n4475) );
  INV_X1 U5608 ( .A(DATAI_2_), .ZN(n4729) );
  NOR2_X1 U5609 ( .A1(n4723), .A2(n4729), .ZN(n4484) );
  AOI21_X1 U5610 ( .B1(n6467), .B2(EAX_REG_18__SCAN_IN), .A(n4484), .ZN(n4474)
         );
  OAI21_X1 U5611 ( .B1(n4493), .B2(n4475), .A(n4474), .ZN(U2926) );
  INV_X1 U5612 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n4478) );
  AOI21_X1 U5613 ( .B1(n6467), .B2(EAX_REG_23__SCAN_IN), .A(n4476), .ZN(n4477)
         );
  OAI21_X1 U5614 ( .B1(n4493), .B2(n4478), .A(n4477), .ZN(U2931) );
  INV_X1 U5615 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n4481) );
  AOI21_X1 U5616 ( .B1(n6467), .B2(EAX_REG_4__SCAN_IN), .A(n4479), .ZN(n4480)
         );
  OAI21_X1 U5617 ( .B1(n4493), .B2(n4481), .A(n4480), .ZN(U2943) );
  INV_X1 U5618 ( .A(LWORD_REG_3__SCAN_IN), .ZN(n4483) );
  INV_X1 U5619 ( .A(DATAI_3_), .ZN(n4790) );
  NOR2_X1 U5620 ( .A1(n4723), .A2(n4790), .ZN(n4487) );
  AOI21_X1 U5621 ( .B1(n6467), .B2(EAX_REG_3__SCAN_IN), .A(n4487), .ZN(n4482)
         );
  OAI21_X1 U5622 ( .B1(n4493), .B2(n4483), .A(n4482), .ZN(U2942) );
  INV_X1 U5623 ( .A(LWORD_REG_2__SCAN_IN), .ZN(n4486) );
  AOI21_X1 U5624 ( .B1(n6467), .B2(EAX_REG_2__SCAN_IN), .A(n4484), .ZN(n4485)
         );
  OAI21_X1 U5625 ( .B1(n4493), .B2(n4486), .A(n4485), .ZN(U2941) );
  INV_X1 U5626 ( .A(UWORD_REG_3__SCAN_IN), .ZN(n4489) );
  AOI21_X1 U5627 ( .B1(n6467), .B2(EAX_REG_19__SCAN_IN), .A(n4487), .ZN(n4488)
         );
  OAI21_X1 U5628 ( .B1(n4493), .B2(n4489), .A(n4488), .ZN(U2927) );
  INV_X1 U5629 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n4492) );
  AOI21_X1 U5630 ( .B1(n6467), .B2(EAX_REG_24__SCAN_IN), .A(n4490), .ZN(n4491)
         );
  OAI21_X1 U5631 ( .B1(n4493), .B2(n4492), .A(n4491), .ZN(U2932) );
  INV_X1 U5632 ( .A(EAX_REG_24__SCAN_IN), .ZN(n6731) );
  AOI22_X1 U5633 ( .A1(n6449), .A2(UWORD_REG_8__SCAN_IN), .B1(n6448), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4497) );
  OAI21_X1 U5634 ( .B1(n6731), .B2(n4856), .A(n4497), .ZN(U2899) );
  INV_X1 U5635 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4499) );
  AOI22_X1 U5636 ( .A1(n6449), .A2(UWORD_REG_9__SCAN_IN), .B1(n6448), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4498) );
  OAI21_X1 U5637 ( .B1(n4499), .B2(n4856), .A(n4498), .ZN(U2898) );
  INV_X1 U5638 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4501) );
  AOI22_X1 U5639 ( .A1(n6449), .A2(UWORD_REG_10__SCAN_IN), .B1(n6448), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4500) );
  OAI21_X1 U5640 ( .B1(n4501), .B2(n4856), .A(n4500), .ZN(U2897) );
  AOI22_X1 U5641 ( .A1(n6449), .A2(UWORD_REG_14__SCAN_IN), .B1(n6448), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4502) );
  OAI21_X1 U5642 ( .B1(n4091), .B2(n4856), .A(n4502), .ZN(U2893) );
  INV_X1 U5643 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4504) );
  AOI22_X1 U5644 ( .A1(n6449), .A2(UWORD_REG_11__SCAN_IN), .B1(n6448), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4503) );
  OAI21_X1 U5645 ( .B1(n4504), .B2(n4856), .A(n4503), .ZN(U2896) );
  INV_X1 U5646 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4506) );
  AOI22_X1 U5647 ( .A1(n6449), .A2(UWORD_REG_12__SCAN_IN), .B1(n6448), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4505) );
  OAI21_X1 U5648 ( .B1(n4506), .B2(n4856), .A(n4505), .ZN(U2895) );
  INV_X1 U5649 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4772) );
  AOI22_X1 U5650 ( .A1(n6449), .A2(UWORD_REG_13__SCAN_IN), .B1(n6448), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4507) );
  OAI21_X1 U5651 ( .B1(n4772), .B2(n4856), .A(n4507), .ZN(U2894) );
  NAND2_X1 U5652 ( .A1(n6577), .A2(n5923), .ZN(n5919) );
  AOI21_X1 U5653 ( .B1(n4515), .B2(n5921), .A(n5300), .ZN(n4508) );
  AOI21_X1 U5654 ( .B1(n5300), .B2(n5919), .A(n4508), .ZN(n4511) );
  INV_X1 U5655 ( .A(n5565), .ZN(n4509) );
  AOI22_X1 U5656 ( .A1(n6541), .A2(n4509), .B1(n6573), .B2(REIP_REG_0__SCAN_IN), .ZN(n4510) );
  OAI211_X1 U5657 ( .C1(n4512), .C2(n6520), .A(n4511), .B(n4510), .ZN(U3018)
         );
  XNOR2_X1 U5658 ( .A(n4514), .B(n4513), .ZN(n4529) );
  INV_X1 U5659 ( .A(n4515), .ZN(n4516) );
  AOI21_X1 U5660 ( .B1(n5919), .B2(n5300), .A(n4516), .ZN(n4520) );
  NAND2_X1 U5661 ( .A1(n5896), .A2(n4517), .ZN(n4519) );
  MUX2_X1 U5662 ( .A(n4520), .B(n4519), .S(n4518), .Z(n4523) );
  INV_X1 U5663 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6681) );
  NOR2_X1 U5664 ( .A1(n6524), .A2(n6681), .ZN(n4524) );
  AOI21_X1 U5665 ( .B1(n6541), .B2(n4521), .A(n4524), .ZN(n4522) );
  OAI211_X1 U5666 ( .C1(n4529), .C2(n6520), .A(n4523), .B(n4522), .ZN(U3017)
         );
  INV_X1 U5667 ( .A(n4524), .ZN(n4525) );
  OAI21_X1 U5668 ( .B1(n5762), .B2(n6821), .A(n4525), .ZN(n4527) );
  NOR2_X1 U5669 ( .A1(n6405), .A2(n5816), .ZN(n4526) );
  AOI211_X1 U5670 ( .C1(n5764), .C2(n6821), .A(n4527), .B(n4526), .ZN(n4528)
         );
  OAI21_X1 U5671 ( .B1(n4529), .B2(n6298), .A(n4528), .ZN(U2985) );
  INV_X1 U5672 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6299) );
  NAND2_X1 U5673 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6299), .ZN(n4564) );
  INV_X1 U5674 ( .A(n4548), .ZN(n4563) );
  MUX2_X1 U5675 ( .A(n4561), .B(FLUSH_REG_SCAN_IN), .S(STATE2_REG_1__SCAN_IN), 
        .Z(n4532) );
  INV_X1 U5676 ( .A(n4610), .ZN(n4998) );
  NOR2_X1 U5677 ( .A1(n2954), .A2(n4998), .ZN(n4531) );
  XNOR2_X1 U5678 ( .A(n4531), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5547)
         );
  OR3_X1 U5679 ( .A1(n5547), .A2(STATE2_REG_1__SCAN_IN), .A3(n4137), .ZN(n6292) );
  OAI21_X1 U5680 ( .B1(n6293), .B2(n4532), .A(n6292), .ZN(n4533) );
  INV_X1 U5681 ( .A(n4533), .ZN(n4566) );
  OR2_X1 U5682 ( .A1(n4534), .A2(n5104), .ZN(n4544) );
  NAND2_X1 U5683 ( .A1(n4536), .A2(n4535), .ZN(n4558) );
  XNOR2_X1 U5684 ( .A(n4538), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4542)
         );
  XNOR2_X1 U5685 ( .A(n3515), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4539)
         );
  NAND2_X1 U5686 ( .A1(n5270), .A2(n4539), .ZN(n4540) );
  OAI21_X1 U5687 ( .B1(n4542), .B2(n4555), .A(n4540), .ZN(n4541) );
  AOI21_X1 U5688 ( .B1(n4558), .B2(n4542), .A(n4541), .ZN(n4543) );
  NAND2_X1 U5689 ( .A1(n4544), .A2(n4543), .ZN(n5305) );
  INV_X1 U5690 ( .A(n4561), .ZN(n5105) );
  MUX2_X1 U5691 ( .A(n5305), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(n5105), 
        .Z(n5111) );
  NAND2_X1 U5692 ( .A1(n6218), .A2(n4546), .ZN(n4560) );
  MUX2_X1 U5693 ( .A(n4547), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4538), 
        .Z(n4549) );
  NOR2_X1 U5694 ( .A1(n4549), .A2(n4548), .ZN(n4557) );
  AOI21_X1 U5695 ( .B1(n4538), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3525), 
        .ZN(n4550) );
  NOR2_X1 U5696 ( .A1(n4551), .A2(n4550), .ZN(n5981) );
  NAND2_X1 U5697 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4552) );
  XNOR2_X1 U5698 ( .A(n4552), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4553)
         );
  NAND2_X1 U5699 ( .A1(n5270), .A2(n4553), .ZN(n4554) );
  OAI21_X1 U5700 ( .B1(n5981), .B2(n4555), .A(n4554), .ZN(n4556) );
  AOI21_X1 U5701 ( .B1(n4558), .B2(n4557), .A(n4556), .ZN(n4559) );
  NAND2_X1 U5702 ( .A1(n4560), .A2(n4559), .ZN(n5980) );
  MUX2_X1 U5703 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5980), .S(n4561), 
        .Z(n5117) );
  NAND3_X1 U5704 ( .A1(n5111), .A2(n5117), .A3(n5301), .ZN(n4562) );
  OAI211_X1 U5705 ( .C1(n4564), .C2(n4563), .A(n4566), .B(n4562), .ZN(n5125)
         );
  NAND2_X1 U5706 ( .A1(n4566), .A2(n4565), .ZN(n4567) );
  NAND2_X1 U5707 ( .A1(n5125), .A2(n4567), .ZN(n4574) );
  NAND2_X1 U5708 ( .A1(n4574), .A2(n6299), .ZN(n4569) );
  NAND2_X1 U5709 ( .A1(n4569), .A2(n4568), .ZN(n4572) );
  AND2_X1 U5710 ( .A1(n4574), .A2(n4573), .ZN(n6285) );
  AND2_X1 U5711 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6103), .ZN(n5977) );
  OAI22_X1 U5712 ( .A1(n6099), .A2(n6691), .B1(n3583), .B2(n5977), .ZN(n4575)
         );
  OAI21_X1 U5713 ( .B1(n6285), .B2(n4575), .A(n6584), .ZN(n4576) );
  OAI21_X1 U5714 ( .B1(n6584), .B2(n6207), .A(n4576), .ZN(U3465) );
  OR2_X1 U5715 ( .A1(n5972), .A2(n6297), .ZN(n4608) );
  NOR2_X1 U5716 ( .A1(n4905), .A2(n4608), .ZN(n4900) );
  NOR2_X1 U5717 ( .A1(n4900), .A2(n5056), .ZN(n4859) );
  NAND2_X1 U5718 ( .A1(n4734), .A2(n4858), .ZN(n4732) );
  AOI21_X1 U5719 ( .B1(n4859), .B2(n4732), .A(n6691), .ZN(n4582) );
  NAND2_X1 U5720 ( .A1(n6203), .A2(n6297), .ZN(n6149) );
  OAI22_X1 U5721 ( .A1(n3567), .A2(n6149), .B1(n6206), .B2(n5977), .ZN(n4581)
         );
  OAI21_X1 U5722 ( .B1(n4582), .B2(n4581), .A(n6584), .ZN(n4583) );
  OAI21_X1 U5723 ( .B1(n6584), .B2(n5116), .A(n4583), .ZN(U3462) );
  NOR2_X1 U5724 ( .A1(n4585), .A2(n4584), .ZN(n4586) );
  NOR2_X1 U5725 ( .A1(n4788), .A2(n4586), .ZN(n6506) );
  INV_X1 U5726 ( .A(n6506), .ZN(n4730) );
  OR2_X1 U5727 ( .A1(n4587), .A2(n4588), .ZN(n4838) );
  NAND2_X1 U5728 ( .A1(n4587), .A2(n4588), .ZN(n4589) );
  AND2_X1 U5729 ( .A1(n4838), .A2(n4589), .ZN(n6574) );
  AOI22_X1 U5730 ( .A1(n5628), .A2(n6574), .B1(EBX_REG_2__SCAN_IN), .B2(n5627), 
        .ZN(n4590) );
  OAI21_X1 U5731 ( .B1(n4730), .B2(n5630), .A(n4590), .ZN(U2857) );
  AND2_X1 U5732 ( .A1(n4788), .A2(n4789), .ZN(n4592) );
  OAI21_X1 U5733 ( .B1(n4592), .B2(n4591), .A(n4791), .ZN(n5552) );
  XNOR2_X1 U5734 ( .A(n4840), .B(n4825), .ZN(n6553) );
  AOI22_X1 U5735 ( .A1(n5628), .A2(n6553), .B1(n5627), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4593) );
  OAI21_X1 U5736 ( .B1(n5552), .B2(n5630), .A(n4593), .ZN(U2855) );
  INV_X1 U5737 ( .A(n4905), .ZN(n4666) );
  AOI21_X1 U5738 ( .B1(n4666), .B2(n5972), .A(n5816), .ZN(n4596) );
  INV_X1 U5739 ( .A(n6149), .ZN(n4948) );
  INV_X1 U5740 ( .A(n3583), .ZN(n4594) );
  NAND2_X1 U5741 ( .A1(n6218), .A2(n4594), .ZN(n6152) );
  INV_X1 U5742 ( .A(n6152), .ZN(n4595) );
  NOR2_X1 U5743 ( .A1(n4534), .A2(n4435), .ZN(n6065) );
  INV_X1 U5744 ( .A(n4604), .ZN(n4817) );
  AOI21_X1 U5745 ( .B1(n4595), .B2(n6065), .A(n4817), .ZN(n4599) );
  OAI21_X1 U5746 ( .B1(n4596), .B2(n4948), .A(n4599), .ZN(n4597) );
  NAND2_X1 U5747 ( .A1(n4822), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4607)
         );
  INV_X1 U5748 ( .A(n4869), .ZN(n4598) );
  AND2_X1 U5749 ( .A1(n4642), .A2(n2967), .ZN(n6162) );
  INV_X1 U5750 ( .A(n4599), .ZN(n4600) );
  NAND2_X1 U5751 ( .A1(n4600), .A2(n6203), .ZN(n4602) );
  NAND2_X1 U5752 ( .A1(n6208), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4601) );
  NAND2_X1 U5753 ( .A1(n4602), .A2(n4601), .ZN(n4818) );
  INV_X1 U5754 ( .A(DATAI_0_), .ZN(n4731) );
  NAND2_X1 U5755 ( .A1(n4818), .A2(n6599), .ZN(n4603) );
  OAI21_X1 U5756 ( .B1(n6596), .B2(n4604), .A(n4603), .ZN(n4605) );
  AOI21_X1 U5757 ( .B1(n4983), .B2(n6165), .A(n4605), .ZN(n4606) );
  OAI211_X1 U5758 ( .C1(n6281), .C2(n6602), .A(n4607), .B(n4606), .ZN(U3140)
         );
  INV_X1 U5759 ( .A(n4608), .ZN(n4609) );
  AOI21_X1 U5760 ( .B1(n4734), .B2(n4609), .A(n6691), .ZN(n4616) );
  INV_X1 U5761 ( .A(n4899), .ZN(n4997) );
  NOR2_X1 U5762 ( .A1(n3583), .A2(n4610), .ZN(n4612) );
  AND3_X1 U5763 ( .A1(n6101), .A2(n5116), .A3(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), 
        .ZN(n5000) );
  NAND2_X1 U5764 ( .A1(n5000), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4643) );
  INV_X1 U5765 ( .A(n4643), .ZN(n4611) );
  AOI21_X1 U5766 ( .B1(n4997), .B2(n4612), .A(n4611), .ZN(n4615) );
  INV_X1 U5767 ( .A(n4615), .ZN(n4613) );
  NOR2_X1 U5768 ( .A1(n5972), .A2(n5986), .ZN(n4665) );
  NAND2_X1 U5769 ( .A1(n4734), .A2(n4665), .ZN(n5039) );
  INV_X1 U5770 ( .A(n4734), .ZN(n4736) );
  INV_X1 U5771 ( .A(n6095), .ZN(n4644) );
  INV_X1 U5772 ( .A(n6165), .ZN(n6597) );
  OAI22_X1 U5773 ( .A1(n4644), .A2(n6597), .B1(n6596), .B2(n4643), .ZN(n4614)
         );
  AOI21_X1 U5774 ( .B1(n6222), .B2(n4646), .A(n4614), .ZN(n4619) );
  NAND2_X1 U5775 ( .A1(n4616), .A2(n4615), .ZN(n4617) );
  NAND2_X1 U5776 ( .A1(n4647), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4618) );
  OAI211_X1 U5777 ( .C1(n4650), .C2(n6220), .A(n4619), .B(n4618), .ZN(U3060)
         );
  INV_X1 U5778 ( .A(DATAI_1_), .ZN(n4728) );
  NAND2_X1 U5779 ( .A1(n5795), .A2(DATAI_25_), .ZN(n6168) );
  INV_X1 U5780 ( .A(n6168), .ZN(n6230) );
  AND2_X1 U5781 ( .A1(n4642), .A2(n4620), .ZN(n6226) );
  OAI22_X1 U5782 ( .A1(n4644), .A2(n6233), .B1(n6071), .B2(n4643), .ZN(n4621)
         );
  AOI21_X1 U5783 ( .B1(n6230), .B2(n4646), .A(n4621), .ZN(n4623) );
  NAND2_X1 U5784 ( .A1(n4647), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4622) );
  OAI211_X1 U5785 ( .C1(n4650), .C2(n6228), .A(n4623), .B(n4622), .ZN(U3061)
         );
  NAND2_X1 U5786 ( .A1(n5795), .A2(DATAI_26_), .ZN(n6173) );
  INV_X1 U5787 ( .A(n6173), .ZN(n6238) );
  AND2_X1 U5788 ( .A1(n4642), .A2(n4624), .ZN(n6234) );
  OAI22_X1 U5789 ( .A1(n4644), .A2(n6241), .B1(n6075), .B2(n4643), .ZN(n4625)
         );
  AOI21_X1 U5790 ( .B1(n6238), .B2(n4646), .A(n4625), .ZN(n4627) );
  NAND2_X1 U5791 ( .A1(n4647), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4626) );
  OAI211_X1 U5792 ( .C1(n4650), .C2(n6236), .A(n4627), .B(n4626), .ZN(U3062)
         );
  INV_X1 U5793 ( .A(DATAI_5_), .ZN(n6764) );
  NAND2_X1 U5794 ( .A1(n5795), .A2(DATAI_29_), .ZN(n6623) );
  INV_X1 U5795 ( .A(n6623), .ZN(n6260) );
  AND2_X1 U5796 ( .A1(n4642), .A2(n3235), .ZN(n6256) );
  OAI22_X1 U5797 ( .A1(n4644), .A2(n6618), .B1(n6617), .B2(n4643), .ZN(n4628)
         );
  AOI21_X1 U5798 ( .B1(n6260), .B2(n4646), .A(n4628), .ZN(n4630) );
  NAND2_X1 U5799 ( .A1(n4647), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4629) );
  OAI211_X1 U5800 ( .C1(n4650), .C2(n6258), .A(n4630), .B(n4629), .ZN(U3065)
         );
  INV_X1 U5801 ( .A(DATAI_6_), .ZN(n6726) );
  NAND2_X1 U5802 ( .A1(n5795), .A2(DATAI_30_), .ZN(n6630) );
  INV_X1 U5803 ( .A(n6630), .ZN(n6267) );
  AND2_X1 U5804 ( .A1(n4642), .A2(n4631), .ZN(n6263) );
  OAI22_X1 U5805 ( .A1(n4644), .A2(n6625), .B1(n6624), .B2(n4643), .ZN(n4632)
         );
  AOI21_X1 U5806 ( .B1(n6267), .B2(n4646), .A(n4632), .ZN(n4634) );
  NAND2_X1 U5807 ( .A1(n4647), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4633) );
  OAI211_X1 U5808 ( .C1(n4650), .C2(n6265), .A(n4634), .B(n4633), .ZN(U3066)
         );
  NAND2_X1 U5809 ( .A1(n5795), .A2(DATAI_31_), .ZN(n6642) );
  INV_X1 U5810 ( .A(n6642), .ZN(n6277) );
  OAI22_X1 U5811 ( .A1(n4644), .A2(n6633), .B1(n6632), .B2(n4643), .ZN(n4635)
         );
  AOI21_X1 U5812 ( .B1(n6277), .B2(n4646), .A(n4635), .ZN(n4637) );
  NAND2_X1 U5813 ( .A1(n4647), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4636) );
  OAI211_X1 U5814 ( .C1(n4650), .C2(n6274), .A(n4637), .B(n4636), .ZN(U3067)
         );
  NAND2_X1 U5815 ( .A1(n5795), .A2(DATAI_27_), .ZN(n6609) );
  INV_X1 U5816 ( .A(n6609), .ZN(n6246) );
  OAI22_X1 U5817 ( .A1(n4644), .A2(n6604), .B1(n6603), .B2(n4643), .ZN(n4639)
         );
  AOI21_X1 U5818 ( .B1(n6246), .B2(n4646), .A(n4639), .ZN(n4641) );
  NAND2_X1 U5819 ( .A1(n4647), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4640) );
  OAI211_X1 U5820 ( .C1(n4650), .C2(n6244), .A(n4641), .B(n4640), .ZN(U3063)
         );
  NAND2_X1 U5821 ( .A1(n5795), .A2(DATAI_28_), .ZN(n6616) );
  AND2_X1 U5822 ( .A1(n4642), .A2(n3209), .ZN(n6249) );
  OAI22_X1 U5823 ( .A1(n4644), .A2(n6611), .B1(n6610), .B2(n4643), .ZN(n4645)
         );
  AOI21_X1 U5824 ( .B1(n6253), .B2(n4646), .A(n4645), .ZN(n4649) );
  NAND2_X1 U5825 ( .A1(n4647), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4648) );
  OAI211_X1 U5826 ( .C1(n4650), .C2(n6251), .A(n4649), .B(n4648), .ZN(U3064)
         );
  INV_X1 U5827 ( .A(n5056), .ZN(n4651) );
  OAI21_X1 U5828 ( .B1(n4651), .B2(n5976), .A(n6203), .ZN(n4657) );
  AND2_X1 U5829 ( .A1(n4534), .A2(n6400), .ZN(n4861) );
  NAND2_X1 U5830 ( .A1(n4861), .A2(n6218), .ZN(n5063) );
  OR2_X1 U5831 ( .A1(n5063), .A2(n3583), .ZN(n4653) );
  AND2_X1 U5832 ( .A1(n5112), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6102)
         );
  INV_X1 U5833 ( .A(n4652), .ZN(n5108) );
  NAND2_X1 U5834 ( .A1(n6102), .A2(n5108), .ZN(n6631) );
  NAND3_X1 U5835 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n5112), .ZN(n5058) );
  OAI22_X1 U5836 ( .A1(n4657), .A2(n4654), .B1(n5058), .B2(n6768), .ZN(n6636)
         );
  INV_X1 U5837 ( .A(n6636), .ZN(n4664) );
  INV_X1 U5838 ( .A(n4654), .ZN(n4656) );
  AOI21_X1 U5839 ( .B1(n6691), .B2(n5058), .A(n4902), .ZN(n4655) );
  NOR2_X1 U5840 ( .A1(n6641), .A2(n6168), .ZN(n4659) );
  OAI22_X1 U5841 ( .A1(n6634), .A2(n6233), .B1(n6071), .B2(n6631), .ZN(n4658)
         );
  AOI211_X1 U5842 ( .C1(n6638), .C2(INSTQUEUE_REG_11__1__SCAN_IN), .A(n4659), 
        .B(n4658), .ZN(n4660) );
  OAI21_X1 U5843 ( .B1(n4664), .B2(n6228), .A(n4660), .ZN(U3109) );
  NOR2_X1 U5844 ( .A1(n6641), .A2(n6173), .ZN(n4662) );
  OAI22_X1 U5845 ( .A1(n6634), .A2(n6241), .B1(n6075), .B2(n6631), .ZN(n4661)
         );
  AOI211_X1 U5846 ( .C1(n6638), .C2(INSTQUEUE_REG_11__2__SCAN_IN), .A(n4662), 
        .B(n4661), .ZN(n4663) );
  OAI21_X1 U5847 ( .B1(n4664), .B2(n6236), .A(n4663), .ZN(U3110) );
  AOI21_X1 U5848 ( .B1(n6634), .B2(n4942), .A(n6297), .ZN(n4671) );
  OAI21_X1 U5849 ( .B1(n4899), .B2(n4998), .A(n6203), .ZN(n4670) );
  AND2_X1 U5850 ( .A1(n4667), .A2(n6101), .ZN(n4907) );
  NAND2_X1 U5851 ( .A1(n4907), .A2(n6207), .ZN(n4681) );
  NAND2_X1 U5852 ( .A1(n4672), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6211) );
  INV_X1 U5853 ( .A(n6211), .ZN(n6023) );
  INV_X1 U5854 ( .A(n6022), .ZN(n4955) );
  OAI21_X1 U5855 ( .B1(n4956), .B2(n6768), .A(n4951), .ZN(n6105) );
  AOI211_X1 U5856 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4681), .A(n6023), .B(
        n6105), .ZN(n4669) );
  OAI21_X1 U5857 ( .B1(n4671), .B2(n4670), .A(n4669), .ZN(n4679) );
  NAND2_X1 U5858 ( .A1(n4679), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4678)
         );
  INV_X1 U5859 ( .A(n4942), .ZN(n4676) );
  NOR2_X1 U5860 ( .A1(n4899), .A2(n6691), .ZN(n5004) );
  NAND2_X1 U5861 ( .A1(n5004), .A2(n6218), .ZN(n4674) );
  NAND2_X1 U5862 ( .A1(n4956), .A2(n6022), .ZN(n6108) );
  OR2_X1 U5863 ( .A1(n4672), .A2(n6768), .ZN(n6216) );
  OR2_X1 U5864 ( .A1(n6108), .A2(n6216), .ZN(n4673) );
  AND2_X1 U5865 ( .A1(n4674), .A2(n4673), .ZN(n4680) );
  OAI22_X1 U5866 ( .A1(n6596), .A2(n4681), .B1(n4680), .B2(n6220), .ZN(n4675)
         );
  AOI21_X1 U5867 ( .B1(n4676), .B2(n6165), .A(n4675), .ZN(n4677) );
  OAI211_X1 U5868 ( .C1(n6634), .C2(n6602), .A(n4678), .B(n4677), .ZN(U3116)
         );
  INV_X1 U5869 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4685) );
  INV_X1 U5870 ( .A(n4681), .ZN(n4706) );
  AOI22_X1 U5871 ( .A1(n4707), .A2(n6637), .B1(n6272), .B2(n4706), .ZN(n4682)
         );
  OAI21_X1 U5872 ( .B1(n4942), .B2(n6633), .A(n4682), .ZN(n4683) );
  AOI21_X1 U5873 ( .B1(n6277), .B2(n4710), .A(n4683), .ZN(n4684) );
  OAI21_X1 U5874 ( .B1(n4713), .B2(n4685), .A(n4684), .ZN(U3123) );
  INV_X1 U5875 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4689) );
  AOI22_X1 U5876 ( .A1(n4707), .A2(n6627), .B1(n6263), .B2(n4706), .ZN(n4686)
         );
  OAI21_X1 U5877 ( .B1(n4942), .B2(n6625), .A(n4686), .ZN(n4687) );
  AOI21_X1 U5878 ( .B1(n6267), .B2(n4710), .A(n4687), .ZN(n4688) );
  OAI21_X1 U5879 ( .B1(n4713), .B2(n4689), .A(n4688), .ZN(U3122) );
  INV_X1 U5880 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4693) );
  AOI22_X1 U5881 ( .A1(n4707), .A2(n6119), .B1(n6234), .B2(n4706), .ZN(n4690)
         );
  OAI21_X1 U5882 ( .B1(n4942), .B2(n6241), .A(n4690), .ZN(n4691) );
  AOI21_X1 U5883 ( .B1(n6238), .B2(n4710), .A(n4691), .ZN(n4692) );
  OAI21_X1 U5884 ( .B1(n4713), .B2(n4693), .A(n4692), .ZN(U3118) );
  INV_X1 U5885 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4697) );
  AOI22_X1 U5886 ( .A1(n4707), .A2(n6613), .B1(n6249), .B2(n4706), .ZN(n4694)
         );
  OAI21_X1 U5887 ( .B1(n4942), .B2(n6611), .A(n4694), .ZN(n4695) );
  AOI21_X1 U5888 ( .B1(n6253), .B2(n4710), .A(n4695), .ZN(n4696) );
  OAI21_X1 U5889 ( .B1(n4713), .B2(n4697), .A(n4696), .ZN(U3120) );
  INV_X1 U5890 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4701) );
  AOI22_X1 U5891 ( .A1(n4707), .A2(n6114), .B1(n6226), .B2(n4706), .ZN(n4698)
         );
  OAI21_X1 U5892 ( .B1(n4942), .B2(n6233), .A(n4698), .ZN(n4699) );
  AOI21_X1 U5893 ( .B1(n6230), .B2(n4710), .A(n4699), .ZN(n4700) );
  OAI21_X1 U5894 ( .B1(n4713), .B2(n4701), .A(n4700), .ZN(U3117) );
  INV_X1 U5895 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4705) );
  AOI22_X1 U5896 ( .A1(n4707), .A2(n6606), .B1(n6242), .B2(n4706), .ZN(n4702)
         );
  OAI21_X1 U5897 ( .B1(n4942), .B2(n6604), .A(n4702), .ZN(n4703) );
  AOI21_X1 U5898 ( .B1(n6246), .B2(n4710), .A(n4703), .ZN(n4704) );
  OAI21_X1 U5899 ( .B1(n4713), .B2(n4705), .A(n4704), .ZN(U3119) );
  INV_X1 U5900 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4712) );
  AOI22_X1 U5901 ( .A1(n4707), .A2(n6620), .B1(n6256), .B2(n4706), .ZN(n4708)
         );
  OAI21_X1 U5902 ( .B1(n4942), .B2(n6618), .A(n4708), .ZN(n4709) );
  AOI21_X1 U5903 ( .B1(n6260), .B2(n4710), .A(n4709), .ZN(n4711) );
  OAI21_X1 U5904 ( .B1(n4713), .B2(n4712), .A(n4711), .ZN(U3121) );
  INV_X1 U5905 ( .A(n4714), .ZN(n4721) );
  NAND2_X1 U5906 ( .A1(n3080), .A2(n4715), .ZN(n4718) );
  OAI22_X1 U5907 ( .A1(n4137), .A2(n4718), .B1(n4717), .B2(n4716), .ZN(n4719)
         );
  AND2_X1 U5908 ( .A1(n3215), .A2(n4724), .ZN(n4727) );
  NOR2_X1 U5909 ( .A1(n4727), .A2(n4726), .ZN(n4725) );
  INV_X1 U5910 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6447) );
  OAI222_X1 U5911 ( .A1(n6405), .A2(n5675), .B1(n5670), .B2(n4728), .C1(n6420), 
        .C2(n6447), .ZN(U2890) );
  INV_X1 U5912 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6445) );
  OAI222_X1 U5913 ( .A1(n4730), .A2(n5675), .B1(n5670), .B2(n4729), .C1(n6420), 
        .C2(n6445), .ZN(U2889) );
  INV_X1 U5914 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6452) );
  OAI222_X1 U5915 ( .A1(n5571), .A2(n5675), .B1(n5670), .B2(n4731), .C1(n6420), 
        .C2(n6452), .ZN(U2891) );
  NAND2_X1 U5916 ( .A1(n6065), .A2(n4998), .ZN(n6060) );
  OR2_X1 U5917 ( .A1(n6060), .A2(n3583), .ZN(n4733) );
  NAND2_X1 U5918 ( .A1(n4733), .A2(n4763), .ZN(n4741) );
  NAND2_X1 U5919 ( .A1(n4734), .A2(n4869), .ZN(n6143) );
  OAI22_X1 U5920 ( .A1(n6098), .A2(n6623), .B1(n4763), .B2(n6617), .ZN(n4737)
         );
  AOI21_X1 U5921 ( .B1(n6187), .B2(n4765), .A(n4737), .ZN(n4744) );
  INV_X1 U5922 ( .A(n4738), .ZN(n4742) );
  INV_X1 U5923 ( .A(n6062), .ZN(n4739) );
  AOI21_X1 U5924 ( .B1(n4739), .B2(n6691), .A(n4902), .ZN(n4740) );
  NAND2_X1 U5925 ( .A1(n4766), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4743) );
  OAI211_X1 U5926 ( .C1(n4769), .C2(n6258), .A(n4744), .B(n4743), .ZN(U3081)
         );
  OAI22_X1 U5927 ( .A1(n6098), .A2(n6602), .B1(n4763), .B2(n6596), .ZN(n4745)
         );
  AOI21_X1 U5928 ( .B1(n6165), .B2(n4765), .A(n4745), .ZN(n4747) );
  NAND2_X1 U5929 ( .A1(n4766), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4746) );
  OAI211_X1 U5930 ( .C1(n4769), .C2(n6220), .A(n4747), .B(n4746), .ZN(U3076)
         );
  OAI22_X1 U5931 ( .A1(n6098), .A2(n6616), .B1(n4763), .B2(n6610), .ZN(n4748)
         );
  AOI21_X1 U5932 ( .B1(n6183), .B2(n4765), .A(n4748), .ZN(n4750) );
  NAND2_X1 U5933 ( .A1(n4766), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4749) );
  OAI211_X1 U5934 ( .C1(n4769), .C2(n6251), .A(n4750), .B(n4749), .ZN(U3080)
         );
  OAI22_X1 U5935 ( .A1(n6098), .A2(n6609), .B1(n4763), .B2(n6603), .ZN(n4751)
         );
  AOI21_X1 U5936 ( .B1(n6179), .B2(n4765), .A(n4751), .ZN(n4753) );
  NAND2_X1 U5937 ( .A1(n4766), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4752) );
  OAI211_X1 U5938 ( .C1(n4769), .C2(n6244), .A(n4753), .B(n4752), .ZN(U3079)
         );
  OAI22_X1 U5939 ( .A1(n6098), .A2(n6173), .B1(n4763), .B2(n6075), .ZN(n4754)
         );
  AOI21_X1 U5940 ( .B1(n6175), .B2(n4765), .A(n4754), .ZN(n4756) );
  NAND2_X1 U5941 ( .A1(n4766), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4755) );
  OAI211_X1 U5942 ( .C1(n4769), .C2(n6236), .A(n4756), .B(n4755), .ZN(U3078)
         );
  OAI22_X1 U5943 ( .A1(n6098), .A2(n6642), .B1(n4763), .B2(n6632), .ZN(n4757)
         );
  AOI21_X1 U5944 ( .B1(n6198), .B2(n4765), .A(n4757), .ZN(n4759) );
  NAND2_X1 U5945 ( .A1(n4766), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4758) );
  OAI211_X1 U5946 ( .C1(n4769), .C2(n6274), .A(n4759), .B(n4758), .ZN(U3083)
         );
  OAI22_X1 U5947 ( .A1(n6098), .A2(n6630), .B1(n4763), .B2(n6624), .ZN(n4760)
         );
  AOI21_X1 U5948 ( .B1(n6191), .B2(n4765), .A(n4760), .ZN(n4762) );
  NAND2_X1 U5949 ( .A1(n4766), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4761) );
  OAI211_X1 U5950 ( .C1(n4769), .C2(n6265), .A(n4762), .B(n4761), .ZN(U3082)
         );
  OAI22_X1 U5951 ( .A1(n6098), .A2(n6168), .B1(n4763), .B2(n6071), .ZN(n4764)
         );
  AOI21_X1 U5952 ( .B1(n6170), .B2(n4765), .A(n4764), .ZN(n4768) );
  NAND2_X1 U5953 ( .A1(n4766), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4767) );
  OAI211_X1 U5954 ( .C1(n4769), .C2(n6228), .A(n4768), .B(n4767), .ZN(U3077)
         );
  NAND2_X1 U5955 ( .A1(n6464), .A2(UWORD_REG_13__SCAN_IN), .ZN(n4771) );
  OAI211_X1 U5956 ( .C1(n6473), .C2(n4772), .A(n4771), .B(n4770), .ZN(U2937)
         );
  INV_X1 U5957 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4774) );
  NAND2_X1 U5958 ( .A1(n6464), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4773) );
  NAND2_X1 U5959 ( .A1(n6470), .A2(DATAI_0_), .ZN(n4780) );
  OAI211_X1 U5960 ( .C1(n6473), .C2(n4774), .A(n4773), .B(n4780), .ZN(U2924)
         );
  NAND2_X1 U5961 ( .A1(n6464), .A2(LWORD_REG_6__SCAN_IN), .ZN(n4775) );
  NAND2_X1 U5962 ( .A1(n6470), .A2(DATAI_6_), .ZN(n4778) );
  OAI211_X1 U5963 ( .C1(n6473), .C2(n4776), .A(n4775), .B(n4778), .ZN(U2945)
         );
  INV_X1 U5964 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4852) );
  NAND2_X1 U5965 ( .A1(n6464), .A2(UWORD_REG_5__SCAN_IN), .ZN(n4777) );
  NAND2_X1 U5966 ( .A1(n6470), .A2(DATAI_5_), .ZN(n4782) );
  OAI211_X1 U5967 ( .C1(n6473), .C2(n4852), .A(n4777), .B(n4782), .ZN(U2929)
         );
  NAND2_X1 U5968 ( .A1(n6464), .A2(UWORD_REG_6__SCAN_IN), .ZN(n4779) );
  OAI211_X1 U5969 ( .C1(n6473), .C2(n4848), .A(n4779), .B(n4778), .ZN(U2930)
         );
  NAND2_X1 U5970 ( .A1(n6464), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4781) );
  OAI211_X1 U5971 ( .C1(n6473), .C2(n6452), .A(n4781), .B(n4780), .ZN(U2939)
         );
  NAND2_X1 U5972 ( .A1(n6464), .A2(LWORD_REG_5__SCAN_IN), .ZN(n4783) );
  OAI211_X1 U5973 ( .C1(n6473), .C2(n4784), .A(n4783), .B(n4782), .ZN(U2944)
         );
  NAND2_X1 U5974 ( .A1(n6464), .A2(LWORD_REG_1__SCAN_IN), .ZN(n4786) );
  OAI211_X1 U5975 ( .C1(n6473), .C2(n6447), .A(n4786), .B(n4785), .ZN(U2940)
         );
  INV_X1 U5976 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6441) );
  OAI222_X1 U5977 ( .A1(n5552), .A2(n5675), .B1(n5670), .B2(n4787), .C1(n6420), 
        .C2(n6441), .ZN(U2887) );
  XOR2_X1 U5978 ( .A(n4789), .B(n4788), .Z(n6497) );
  INV_X1 U5979 ( .A(n6497), .ZN(n4841) );
  INV_X1 U5980 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6443) );
  OAI222_X1 U5981 ( .A1(n4841), .A2(n5675), .B1(n5670), .B2(n4790), .C1(n6420), 
        .C2(n6443), .ZN(U2888) );
  XNOR2_X1 U5982 ( .A(n3065), .B(n4792), .ZN(n6488) );
  INV_X1 U5983 ( .A(n6488), .ZN(n4829) );
  OAI222_X1 U5984 ( .A1(n5675), .A2(n4829), .B1(n6420), .B2(n4784), .C1(n6764), 
        .C2(n5670), .ZN(U2886) );
  AOI22_X1 U5985 ( .A1(n4818), .A2(n6606), .B1(n4817), .B2(n6242), .ZN(n4794)
         );
  NAND2_X1 U5986 ( .A1(n4983), .A2(n6179), .ZN(n4793) );
  OAI211_X1 U5987 ( .C1(n6281), .C2(n6609), .A(n4794), .B(n4793), .ZN(n4795)
         );
  AOI21_X1 U5988 ( .B1(n4822), .B2(INSTQUEUE_REG_15__3__SCAN_IN), .A(n4795), 
        .ZN(n4796) );
  INV_X1 U5989 ( .A(n4796), .ZN(U3143) );
  AOI22_X1 U5990 ( .A1(n4818), .A2(n6613), .B1(n4817), .B2(n6249), .ZN(n4798)
         );
  NAND2_X1 U5991 ( .A1(n4983), .A2(n6183), .ZN(n4797) );
  OAI211_X1 U5992 ( .C1(n6281), .C2(n6616), .A(n4798), .B(n4797), .ZN(n4799)
         );
  AOI21_X1 U5993 ( .B1(n4822), .B2(INSTQUEUE_REG_15__4__SCAN_IN), .A(n4799), 
        .ZN(n4800) );
  INV_X1 U5994 ( .A(n4800), .ZN(U3144) );
  AOI22_X1 U5995 ( .A1(n4818), .A2(n6114), .B1(n4817), .B2(n6226), .ZN(n4802)
         );
  NAND2_X1 U5996 ( .A1(n4983), .A2(n6170), .ZN(n4801) );
  OAI211_X1 U5997 ( .C1(n6281), .C2(n6168), .A(n4802), .B(n4801), .ZN(n4803)
         );
  AOI21_X1 U5998 ( .B1(n4822), .B2(INSTQUEUE_REG_15__1__SCAN_IN), .A(n4803), 
        .ZN(n4804) );
  INV_X1 U5999 ( .A(n4804), .ZN(U3141) );
  AOI22_X1 U6000 ( .A1(n4818), .A2(n6119), .B1(n4817), .B2(n6234), .ZN(n4806)
         );
  NAND2_X1 U6001 ( .A1(n4983), .A2(n6175), .ZN(n4805) );
  OAI211_X1 U6002 ( .C1(n6281), .C2(n6173), .A(n4806), .B(n4805), .ZN(n4807)
         );
  AOI21_X1 U6003 ( .B1(n4822), .B2(INSTQUEUE_REG_15__2__SCAN_IN), .A(n4807), 
        .ZN(n4808) );
  INV_X1 U6004 ( .A(n4808), .ZN(U3142) );
  AOI22_X1 U6005 ( .A1(n4818), .A2(n6620), .B1(n4817), .B2(n6256), .ZN(n4810)
         );
  NAND2_X1 U6006 ( .A1(n4983), .A2(n6187), .ZN(n4809) );
  OAI211_X1 U6007 ( .C1(n6281), .C2(n6623), .A(n4810), .B(n4809), .ZN(n4811)
         );
  AOI21_X1 U6008 ( .B1(n4822), .B2(INSTQUEUE_REG_15__5__SCAN_IN), .A(n4811), 
        .ZN(n4812) );
  INV_X1 U6009 ( .A(n4812), .ZN(U3145) );
  AOI22_X1 U6010 ( .A1(n4818), .A2(n6637), .B1(n4817), .B2(n6272), .ZN(n4814)
         );
  NAND2_X1 U6011 ( .A1(n4983), .A2(n6198), .ZN(n4813) );
  OAI211_X1 U6012 ( .C1(n6281), .C2(n6642), .A(n4814), .B(n4813), .ZN(n4815)
         );
  AOI21_X1 U6013 ( .B1(n4822), .B2(INSTQUEUE_REG_15__7__SCAN_IN), .A(n4815), 
        .ZN(n4816) );
  INV_X1 U6014 ( .A(n4816), .ZN(U3147) );
  AOI22_X1 U6015 ( .A1(n4818), .A2(n6627), .B1(n4817), .B2(n6263), .ZN(n4820)
         );
  NAND2_X1 U6016 ( .A1(n4983), .A2(n6191), .ZN(n4819) );
  OAI211_X1 U6017 ( .C1(n6281), .C2(n6630), .A(n4820), .B(n4819), .ZN(n4821)
         );
  AOI21_X1 U6018 ( .B1(n4822), .B2(INSTQUEUE_REG_15__6__SCAN_IN), .A(n4821), 
        .ZN(n4823) );
  INV_X1 U6019 ( .A(n4823), .ZN(U3146) );
  INV_X1 U6020 ( .A(n4840), .ZN(n4826) );
  AOI21_X1 U6021 ( .B1(n4826), .B2(n4825), .A(n4824), .ZN(n4827) );
  OR2_X1 U6022 ( .A1(n4827), .A2(n4895), .ZN(n6538) );
  INV_X1 U6023 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4828) );
  OAI222_X1 U6024 ( .A1(n6538), .A2(n5624), .B1(n5630), .B2(n4829), .C1(n4828), 
        .C2(n5626), .ZN(U2854) );
  OAI21_X1 U6025 ( .B1(n4831), .B2(n4830), .A(n4832), .ZN(n4833) );
  INV_X1 U6026 ( .A(n4833), .ZN(n6554) );
  NAND2_X1 U6027 ( .A1(n6554), .A2(n6505), .ZN(n4836) );
  NOR2_X1 U6028 ( .A1(n6524), .A2(n6657), .ZN(n6552) );
  NOR2_X1 U6029 ( .A1(n6510), .A2(n5551), .ZN(n4834) );
  AOI211_X1 U6030 ( .C1(n6501), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6552), 
        .B(n4834), .ZN(n4835) );
  OAI211_X1 U6031 ( .C1(n5552), .C2(n5816), .A(n4836), .B(n4835), .ZN(U2982)
         );
  NAND2_X1 U6032 ( .A1(n4838), .A2(n4837), .ZN(n4839) );
  NAND2_X1 U6033 ( .A1(n4840), .A2(n4839), .ZN(n5558) );
  INV_X1 U6034 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4842) );
  OAI222_X1 U6035 ( .A1(n5558), .A2(n5624), .B1(n4842), .B2(n5626), .C1(n5630), 
        .C2(n4841), .ZN(U2856) );
  AOI22_X1 U6036 ( .A1(n6436), .A2(UWORD_REG_1__SCAN_IN), .B1(n6439), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4843) );
  OAI21_X1 U6037 ( .B1(n4461), .B2(n4856), .A(n4843), .ZN(U2906) );
  INV_X1 U6038 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4845) );
  AOI22_X1 U6039 ( .A1(n6436), .A2(UWORD_REG_2__SCAN_IN), .B1(n6439), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4844) );
  OAI21_X1 U6040 ( .B1(n4845), .B2(n4856), .A(n4844), .ZN(U2905) );
  AOI22_X1 U6041 ( .A1(n6436), .A2(UWORD_REG_0__SCAN_IN), .B1(n6439), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4846) );
  OAI21_X1 U6042 ( .B1(n4774), .B2(n4856), .A(n4846), .ZN(U2907) );
  INV_X1 U6043 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4848) );
  AOI22_X1 U6044 ( .A1(n6449), .A2(UWORD_REG_6__SCAN_IN), .B1(n6439), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4847) );
  OAI21_X1 U6045 ( .B1(n4848), .B2(n4856), .A(n4847), .ZN(U2901) );
  INV_X1 U6046 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4850) );
  AOI22_X1 U6047 ( .A1(n6449), .A2(UWORD_REG_4__SCAN_IN), .B1(n6439), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4849) );
  OAI21_X1 U6048 ( .B1(n4850), .B2(n4856), .A(n4849), .ZN(U2903) );
  AOI22_X1 U6049 ( .A1(n6449), .A2(UWORD_REG_5__SCAN_IN), .B1(n6439), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4851) );
  OAI21_X1 U6050 ( .B1(n4852), .B2(n4856), .A(n4851), .ZN(U2902) );
  INV_X1 U6051 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4854) );
  AOI22_X1 U6052 ( .A1(n6449), .A2(UWORD_REG_7__SCAN_IN), .B1(n6439), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4853) );
  OAI21_X1 U6053 ( .B1(n4854), .B2(n4856), .A(n4853), .ZN(U2900) );
  INV_X1 U6054 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4857) );
  AOI22_X1 U6055 ( .A1(n6449), .A2(UWORD_REG_3__SCAN_IN), .B1(n6439), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4855) );
  OAI21_X1 U6056 ( .B1(n4857), .B2(n4856), .A(n4855), .ZN(U2904) );
  NAND3_X1 U6057 ( .A1(n4859), .A2(n4858), .A3(n5975), .ZN(n4860) );
  NAND2_X1 U6058 ( .A1(n4860), .A2(n6203), .ZN(n4867) );
  NAND2_X1 U6059 ( .A1(n6206), .A2(n4861), .ZN(n6028) );
  OR2_X1 U6060 ( .A1(n6028), .A2(n3583), .ZN(n4862) );
  NOR2_X1 U6061 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4950) );
  NAND2_X1 U6062 ( .A1(n4950), .A2(n5108), .ZN(n6588) );
  NAND3_X1 U6063 ( .A1(n4950), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        STATE2_REG_2__SCAN_IN), .ZN(n4863) );
  INV_X1 U6064 ( .A(n4864), .ZN(n4866) );
  NAND2_X1 U6065 ( .A1(n4950), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6025) );
  AOI21_X1 U6066 ( .B1(n6025), .B2(n6691), .A(n4902), .ZN(n4865) );
  NOR2_X1 U6067 ( .A1(n6595), .A2(n6602), .ZN(n4871) );
  OAI22_X1 U6068 ( .A1(n6589), .A2(n6597), .B1(n6596), .B2(n6588), .ZN(n4870)
         );
  AOI211_X1 U6069 ( .C1(n6592), .C2(INSTQUEUE_REG_3__0__SCAN_IN), .A(n4871), 
        .B(n4870), .ZN(n4872) );
  OAI21_X1 U6070 ( .B1(n4888), .B2(n6220), .A(n4872), .ZN(U3044) );
  NOR2_X1 U6071 ( .A1(n6595), .A2(n6642), .ZN(n4874) );
  OAI22_X1 U6072 ( .A1(n6589), .A2(n6633), .B1(n6632), .B2(n6588), .ZN(n4873)
         );
  AOI211_X1 U6073 ( .C1(n6592), .C2(INSTQUEUE_REG_3__7__SCAN_IN), .A(n4874), 
        .B(n4873), .ZN(n4875) );
  OAI21_X1 U6074 ( .B1(n4888), .B2(n6274), .A(n4875), .ZN(U3051) );
  NOR2_X1 U6075 ( .A1(n6595), .A2(n6173), .ZN(n4877) );
  OAI22_X1 U6076 ( .A1(n6589), .A2(n6241), .B1(n6075), .B2(n6588), .ZN(n4876)
         );
  AOI211_X1 U6077 ( .C1(n6592), .C2(INSTQUEUE_REG_3__2__SCAN_IN), .A(n4877), 
        .B(n4876), .ZN(n4878) );
  OAI21_X1 U6078 ( .B1(n4888), .B2(n6236), .A(n4878), .ZN(U3046) );
  NOR2_X1 U6079 ( .A1(n6595), .A2(n6623), .ZN(n4880) );
  OAI22_X1 U6080 ( .A1(n6589), .A2(n6618), .B1(n6617), .B2(n6588), .ZN(n4879)
         );
  AOI211_X1 U6081 ( .C1(n6592), .C2(INSTQUEUE_REG_3__5__SCAN_IN), .A(n4880), 
        .B(n4879), .ZN(n4881) );
  OAI21_X1 U6082 ( .B1(n4888), .B2(n6258), .A(n4881), .ZN(U3049) );
  NOR2_X1 U6083 ( .A1(n6595), .A2(n6609), .ZN(n4883) );
  OAI22_X1 U6084 ( .A1(n6589), .A2(n6604), .B1(n6603), .B2(n6588), .ZN(n4882)
         );
  AOI211_X1 U6085 ( .C1(n6592), .C2(INSTQUEUE_REG_3__3__SCAN_IN), .A(n4883), 
        .B(n4882), .ZN(n4884) );
  OAI21_X1 U6086 ( .B1(n4888), .B2(n6244), .A(n4884), .ZN(U3047) );
  NOR2_X1 U6087 ( .A1(n6595), .A2(n6168), .ZN(n4886) );
  OAI22_X1 U6088 ( .A1(n6589), .A2(n6233), .B1(n6071), .B2(n6588), .ZN(n4885)
         );
  AOI211_X1 U6089 ( .C1(n6592), .C2(INSTQUEUE_REG_3__1__SCAN_IN), .A(n4886), 
        .B(n4885), .ZN(n4887) );
  OAI21_X1 U6090 ( .B1(n4888), .B2(n6228), .A(n4887), .ZN(U3045) );
  AND2_X1 U6091 ( .A1(n4890), .A2(n4889), .ZN(n4892) );
  OR2_X1 U6092 ( .A1(n4892), .A2(n4891), .ZN(n5537) );
  OR2_X1 U6093 ( .A1(n4895), .A2(n4894), .ZN(n4896) );
  NAND2_X1 U6094 ( .A1(n4893), .A2(n4896), .ZN(n5535) );
  INV_X1 U6095 ( .A(n5535), .ZN(n4897) );
  AOI22_X1 U6096 ( .A1(n5628), .A2(n4897), .B1(n5627), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4898) );
  OAI21_X1 U6097 ( .B1(n5537), .B2(n5630), .A(n4898), .ZN(U2853) );
  INV_X1 U6098 ( .A(n4907), .ZN(n4903) );
  NAND2_X1 U6099 ( .A1(n4907), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4910) );
  OAI21_X1 U6100 ( .B1(n6152), .B2(n4899), .A(n4910), .ZN(n4906) );
  NOR3_X1 U6101 ( .A1(n4900), .A2(n6691), .A3(n4906), .ZN(n4901) );
  INV_X1 U6102 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4914) );
  NAND2_X1 U6103 ( .A1(n4906), .A2(n6203), .ZN(n4909) );
  NAND2_X1 U6104 ( .A1(n4907), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4908) );
  NAND2_X1 U6105 ( .A1(n4909), .A2(n4908), .ZN(n4940) );
  INV_X1 U6106 ( .A(n4910), .ZN(n4939) );
  AOI22_X1 U6107 ( .A1(n4940), .A2(n6627), .B1(n6263), .B2(n4939), .ZN(n4911)
         );
  OAI21_X1 U6108 ( .B1(n4942), .B2(n6630), .A(n4911), .ZN(n4912) );
  AOI21_X1 U6109 ( .B1(n6191), .B2(n6278), .A(n4912), .ZN(n4913) );
  OAI21_X1 U6110 ( .B1(n4946), .B2(n4914), .A(n4913), .ZN(U3130) );
  INV_X1 U6111 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4918) );
  AOI22_X1 U6112 ( .A1(n4940), .A2(n6606), .B1(n6242), .B2(n4939), .ZN(n4915)
         );
  OAI21_X1 U6113 ( .B1(n4942), .B2(n6609), .A(n4915), .ZN(n4916) );
  AOI21_X1 U6114 ( .B1(n6179), .B2(n6278), .A(n4916), .ZN(n4917) );
  OAI21_X1 U6115 ( .B1(n4946), .B2(n4918), .A(n4917), .ZN(U3127) );
  INV_X1 U6116 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4922) );
  AOI22_X1 U6117 ( .A1(n4940), .A2(n6637), .B1(n6272), .B2(n4939), .ZN(n4919)
         );
  OAI21_X1 U6118 ( .B1(n4942), .B2(n6642), .A(n4919), .ZN(n4920) );
  AOI21_X1 U6119 ( .B1(n6198), .B2(n6278), .A(n4920), .ZN(n4921) );
  OAI21_X1 U6120 ( .B1(n4946), .B2(n4922), .A(n4921), .ZN(U3131) );
  INV_X1 U6121 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4926) );
  AOI22_X1 U6122 ( .A1(n4940), .A2(n6599), .B1(n6162), .B2(n4939), .ZN(n4923)
         );
  OAI21_X1 U6123 ( .B1(n4942), .B2(n6602), .A(n4923), .ZN(n4924) );
  AOI21_X1 U6124 ( .B1(n6165), .B2(n6278), .A(n4924), .ZN(n4925) );
  OAI21_X1 U6125 ( .B1(n4946), .B2(n4926), .A(n4925), .ZN(U3124) );
  INV_X1 U6126 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4930) );
  AOI22_X1 U6127 ( .A1(n4940), .A2(n6114), .B1(n6226), .B2(n4939), .ZN(n4927)
         );
  OAI21_X1 U6128 ( .B1(n4942), .B2(n6168), .A(n4927), .ZN(n4928) );
  AOI21_X1 U6129 ( .B1(n6170), .B2(n6278), .A(n4928), .ZN(n4929) );
  OAI21_X1 U6130 ( .B1(n4946), .B2(n4930), .A(n4929), .ZN(U3125) );
  INV_X1 U6131 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4934) );
  AOI22_X1 U6132 ( .A1(n4940), .A2(n6613), .B1(n6249), .B2(n4939), .ZN(n4931)
         );
  OAI21_X1 U6133 ( .B1(n4942), .B2(n6616), .A(n4931), .ZN(n4932) );
  AOI21_X1 U6134 ( .B1(n6183), .B2(n6278), .A(n4932), .ZN(n4933) );
  OAI21_X1 U6135 ( .B1(n4946), .B2(n4934), .A(n4933), .ZN(U3128) );
  INV_X1 U6136 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4938) );
  AOI22_X1 U6137 ( .A1(n4940), .A2(n6620), .B1(n6256), .B2(n4939), .ZN(n4935)
         );
  OAI21_X1 U6138 ( .B1(n4942), .B2(n6623), .A(n4935), .ZN(n4936) );
  AOI21_X1 U6139 ( .B1(n6187), .B2(n6278), .A(n4936), .ZN(n4937) );
  OAI21_X1 U6140 ( .B1(n4946), .B2(n4938), .A(n4937), .ZN(U3129) );
  INV_X1 U6141 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4945) );
  AOI22_X1 U6142 ( .A1(n4940), .A2(n6119), .B1(n6234), .B2(n4939), .ZN(n4941)
         );
  OAI21_X1 U6143 ( .B1(n4942), .B2(n6173), .A(n4941), .ZN(n4943) );
  AOI21_X1 U6144 ( .B1(n6175), .B2(n6278), .A(n4943), .ZN(n4944) );
  OAI21_X1 U6145 ( .B1(n4946), .B2(n4945), .A(n4944), .ZN(U3126) );
  NOR3_X1 U6146 ( .A1(n6019), .A2(n4983), .A3(n6691), .ZN(n4949) );
  NAND2_X1 U6147 ( .A1(n4534), .A2(n4435), .ZN(n6151) );
  OR2_X1 U6148 ( .A1(n6218), .A2(n6151), .ZN(n5985) );
  OAI21_X1 U6149 ( .B1(n4949), .B2(n4948), .A(n5985), .ZN(n4954) );
  AND2_X1 U6150 ( .A1(n4950), .A2(n6101), .ZN(n5989) );
  NAND2_X1 U6151 ( .A1(n5989), .A2(n6207), .ZN(n4980) );
  INV_X1 U6152 ( .A(n6216), .ZN(n6067) );
  INV_X1 U6153 ( .A(n4956), .ZN(n4952) );
  OAI21_X1 U6154 ( .B1(n6768), .B2(n4952), .A(n4951), .ZN(n5002) );
  AOI211_X1 U6155 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4980), .A(n6067), .B(
        n5002), .ZN(n4953) );
  NAND2_X1 U6156 ( .A1(n4954), .A2(n4953), .ZN(n4979) );
  NAND2_X1 U6157 ( .A1(n4979), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4960) );
  INV_X1 U6158 ( .A(n5985), .ZN(n4957) );
  NOR2_X1 U6159 ( .A1(n4956), .A2(n4955), .ZN(n5005) );
  AOI22_X1 U6160 ( .A1(n4957), .A2(n6203), .B1(n6023), .B2(n5005), .ZN(n4981)
         );
  OAI22_X1 U6161 ( .A1(n4981), .A2(n6251), .B1(n6610), .B2(n4980), .ZN(n4958)
         );
  AOI21_X1 U6162 ( .B1(n4983), .B2(n6253), .A(n4958), .ZN(n4959) );
  OAI211_X1 U6163 ( .C1(n4986), .C2(n6611), .A(n4960), .B(n4959), .ZN(U3024)
         );
  NAND2_X1 U6164 ( .A1(n4979), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4963) );
  OAI22_X1 U6165 ( .A1(n4981), .A2(n6274), .B1(n6632), .B2(n4980), .ZN(n4961)
         );
  AOI21_X1 U6166 ( .B1(n4983), .B2(n6277), .A(n4961), .ZN(n4962) );
  OAI211_X1 U6167 ( .C1(n4986), .C2(n6633), .A(n4963), .B(n4962), .ZN(U3027)
         );
  NAND2_X1 U6168 ( .A1(n4979), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4966) );
  OAI22_X1 U6169 ( .A1(n4981), .A2(n6265), .B1(n6624), .B2(n4980), .ZN(n4964)
         );
  AOI21_X1 U6170 ( .B1(n4983), .B2(n6267), .A(n4964), .ZN(n4965) );
  OAI211_X1 U6171 ( .C1(n4986), .C2(n6625), .A(n4966), .B(n4965), .ZN(U3026)
         );
  NAND2_X1 U6172 ( .A1(n4979), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4969) );
  OAI22_X1 U6173 ( .A1(n4981), .A2(n6244), .B1(n6603), .B2(n4980), .ZN(n4967)
         );
  AOI21_X1 U6174 ( .B1(n4983), .B2(n6246), .A(n4967), .ZN(n4968) );
  OAI211_X1 U6175 ( .C1(n4986), .C2(n6604), .A(n4969), .B(n4968), .ZN(U3023)
         );
  NAND2_X1 U6176 ( .A1(n4979), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4972) );
  OAI22_X1 U6177 ( .A1(n4981), .A2(n6236), .B1(n6075), .B2(n4980), .ZN(n4970)
         );
  AOI21_X1 U6178 ( .B1(n4983), .B2(n6238), .A(n4970), .ZN(n4971) );
  OAI211_X1 U6179 ( .C1(n4986), .C2(n6241), .A(n4972), .B(n4971), .ZN(U3022)
         );
  NAND2_X1 U6180 ( .A1(n4979), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4975) );
  OAI22_X1 U6181 ( .A1(n4981), .A2(n6258), .B1(n6617), .B2(n4980), .ZN(n4973)
         );
  AOI21_X1 U6182 ( .B1(n4983), .B2(n6260), .A(n4973), .ZN(n4974) );
  OAI211_X1 U6183 ( .C1(n4986), .C2(n6618), .A(n4975), .B(n4974), .ZN(U3025)
         );
  NAND2_X1 U6184 ( .A1(n4979), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4978) );
  OAI22_X1 U6185 ( .A1(n4981), .A2(n6220), .B1(n6596), .B2(n4980), .ZN(n4976)
         );
  AOI21_X1 U6186 ( .B1(n4983), .B2(n6222), .A(n4976), .ZN(n4977) );
  OAI211_X1 U6187 ( .C1(n4986), .C2(n6597), .A(n4978), .B(n4977), .ZN(U3020)
         );
  NAND2_X1 U6188 ( .A1(n4979), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4985) );
  OAI22_X1 U6189 ( .A1(n4981), .A2(n6228), .B1(n6071), .B2(n4980), .ZN(n4982)
         );
  AOI21_X1 U6190 ( .B1(n4983), .B2(n6230), .A(n4982), .ZN(n4984) );
  OAI211_X1 U6191 ( .C1(n4986), .C2(n6233), .A(n4985), .B(n4984), .ZN(U3021)
         );
  OAI21_X1 U6192 ( .B1(n4987), .B2(n4989), .A(n4988), .ZN(n5054) );
  NOR2_X1 U6193 ( .A1(n4990), .A2(n4992), .ZN(n6547) );
  NOR2_X1 U6194 ( .A1(n5938), .A2(n6547), .ZN(n6556) );
  NOR3_X1 U6195 ( .A1(n6556), .A2(n6542), .A3(n6546), .ZN(n5955) );
  NAND2_X1 U6196 ( .A1(n5955), .A2(n4991), .ZN(n4996) );
  NOR2_X1 U6197 ( .A1(n6546), .A2(n6542), .ZN(n4993) );
  AOI21_X1 U6198 ( .B1(n5958), .B2(n4992), .A(n5963), .ZN(n6582) );
  OAI21_X1 U6199 ( .B1(n5964), .B2(n4993), .A(n6582), .ZN(n6545) );
  INV_X1 U6200 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6659) );
  OAI22_X1 U6201 ( .A1(n5966), .A2(n5535), .B1(n6659), .B2(n6524), .ZN(n4994)
         );
  AOI21_X1 U6202 ( .B1(n6545), .B2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n4994), 
        .ZN(n4995) );
  OAI211_X1 U6203 ( .C1(n5054), .C2(n6520), .A(n4996), .B(n4995), .ZN(U3012)
         );
  OAI222_X1 U6204 ( .A1(n5537), .A2(n5675), .B1(n5670), .B2(n6726), .C1(n6420), 
        .C2(n4776), .ZN(U2885) );
  NAND3_X1 U6205 ( .A1(n6589), .A2(n6203), .A3(n5039), .ZN(n4999) );
  AOI22_X1 U6206 ( .A1(n4999), .A2(n6149), .B1(n4998), .B2(n4997), .ZN(n5003)
         );
  AND2_X1 U6207 ( .A1(n5000), .A2(n6207), .ZN(n5036) );
  OAI21_X1 U6208 ( .B1(n5036), .B2(n6103), .A(n6211), .ZN(n5001) );
  NOR3_X2 U6209 ( .A1(n5003), .A2(n5002), .A3(n5001), .ZN(n5044) );
  INV_X1 U6210 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5011) );
  NAND2_X1 U6211 ( .A1(n5004), .A2(n6206), .ZN(n5007) );
  NAND2_X1 U6212 ( .A1(n5005), .A2(n6067), .ZN(n5006) );
  NAND2_X1 U6213 ( .A1(n5007), .A2(n5006), .ZN(n5037) );
  AOI22_X1 U6214 ( .A1(n5037), .A2(n6599), .B1(n6162), .B2(n5036), .ZN(n5008)
         );
  OAI21_X1 U6215 ( .B1(n5039), .B2(n6597), .A(n5008), .ZN(n5009) );
  AOI21_X1 U6216 ( .B1(n5041), .B2(n6222), .A(n5009), .ZN(n5010) );
  OAI21_X1 U6217 ( .B1(n5044), .B2(n5011), .A(n5010), .ZN(U3052) );
  INV_X1 U6218 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5015) );
  AOI22_X1 U6219 ( .A1(n5037), .A2(n6114), .B1(n6226), .B2(n5036), .ZN(n5012)
         );
  OAI21_X1 U6220 ( .B1(n5039), .B2(n6233), .A(n5012), .ZN(n5013) );
  AOI21_X1 U6221 ( .B1(n5041), .B2(n6230), .A(n5013), .ZN(n5014) );
  OAI21_X1 U6222 ( .B1(n5044), .B2(n5015), .A(n5014), .ZN(U3053) );
  INV_X1 U6223 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5019) );
  AOI22_X1 U6224 ( .A1(n5037), .A2(n6637), .B1(n6272), .B2(n5036), .ZN(n5016)
         );
  OAI21_X1 U6225 ( .B1(n5039), .B2(n6633), .A(n5016), .ZN(n5017) );
  AOI21_X1 U6226 ( .B1(n5041), .B2(n6277), .A(n5017), .ZN(n5018) );
  OAI21_X1 U6227 ( .B1(n5044), .B2(n5019), .A(n5018), .ZN(U3059) );
  INV_X1 U6228 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5023) );
  AOI22_X1 U6229 ( .A1(n5037), .A2(n6627), .B1(n6263), .B2(n5036), .ZN(n5020)
         );
  OAI21_X1 U6230 ( .B1(n5039), .B2(n6625), .A(n5020), .ZN(n5021) );
  AOI21_X1 U6231 ( .B1(n5041), .B2(n6267), .A(n5021), .ZN(n5022) );
  OAI21_X1 U6232 ( .B1(n5044), .B2(n5023), .A(n5022), .ZN(U3058) );
  INV_X1 U6233 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5027) );
  AOI22_X1 U6234 ( .A1(n5037), .A2(n6620), .B1(n6256), .B2(n5036), .ZN(n5024)
         );
  OAI21_X1 U6235 ( .B1(n5039), .B2(n6618), .A(n5024), .ZN(n5025) );
  AOI21_X1 U6236 ( .B1(n5041), .B2(n6260), .A(n5025), .ZN(n5026) );
  OAI21_X1 U6237 ( .B1(n5044), .B2(n5027), .A(n5026), .ZN(U3057) );
  INV_X1 U6238 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5031) );
  AOI22_X1 U6239 ( .A1(n5037), .A2(n6613), .B1(n6249), .B2(n5036), .ZN(n5028)
         );
  OAI21_X1 U6240 ( .B1(n5039), .B2(n6611), .A(n5028), .ZN(n5029) );
  AOI21_X1 U6241 ( .B1(n5041), .B2(n6253), .A(n5029), .ZN(n5030) );
  OAI21_X1 U6242 ( .B1(n5044), .B2(n5031), .A(n5030), .ZN(U3056) );
  INV_X1 U6243 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5035) );
  AOI22_X1 U6244 ( .A1(n5037), .A2(n6606), .B1(n6242), .B2(n5036), .ZN(n5032)
         );
  OAI21_X1 U6245 ( .B1(n5039), .B2(n6604), .A(n5032), .ZN(n5033) );
  AOI21_X1 U6246 ( .B1(n5041), .B2(n6246), .A(n5033), .ZN(n5034) );
  OAI21_X1 U6247 ( .B1(n5044), .B2(n5035), .A(n5034), .ZN(U3055) );
  INV_X1 U6248 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5043) );
  AOI22_X1 U6249 ( .A1(n5037), .A2(n6119), .B1(n6234), .B2(n5036), .ZN(n5038)
         );
  OAI21_X1 U6250 ( .B1(n5039), .B2(n6241), .A(n5038), .ZN(n5040) );
  AOI21_X1 U6251 ( .B1(n5041), .B2(n6238), .A(n5040), .ZN(n5042) );
  OAI21_X1 U6252 ( .B1(n5044), .B2(n5043), .A(n5042), .ZN(U3054) );
  XNOR2_X1 U6253 ( .A(n4891), .B(n5045), .ZN(n6479) );
  INV_X1 U6254 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6435) );
  OAI222_X1 U6255 ( .A1(n5675), .A2(n6479), .B1(n6420), .B2(n6435), .C1(n5046), 
        .C2(n5670), .ZN(U2884) );
  NAND2_X1 U6256 ( .A1(n4893), .A2(n5047), .ZN(n5048) );
  NAND2_X1 U6257 ( .A1(n5136), .A2(n5048), .ZN(n6531) );
  INV_X1 U6258 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5049) );
  OAI222_X1 U6259 ( .A1(n6531), .A2(n5624), .B1(n5630), .B2(n6479), .C1(n5049), 
        .C2(n5626), .ZN(U2852) );
  INV_X1 U6260 ( .A(n5537), .ZN(n5052) );
  AOI22_X1 U6261 ( .A1(n6501), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .B1(n6573), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n5050) );
  OAI21_X1 U6262 ( .B1(n5536), .B2(n6510), .A(n5050), .ZN(n5051) );
  AOI21_X1 U6263 ( .B1(n5052), .B2(n5795), .A(n5051), .ZN(n5053) );
  OAI21_X1 U6264 ( .B1(n5054), .B2(n6298), .A(n5053), .ZN(U2980) );
  OAI21_X1 U6265 ( .B1(n6199), .B2(n5094), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5057) );
  NAND2_X1 U6266 ( .A1(n5057), .A2(n6203), .ZN(n5064) );
  INV_X1 U6267 ( .A(n5064), .ZN(n5062) );
  NOR2_X1 U6268 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5058), .ZN(n5093)
         );
  NAND2_X1 U6269 ( .A1(n6022), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5059) );
  NAND2_X1 U6270 ( .A1(n5116), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6209) );
  OAI211_X1 U6271 ( .C1(n5093), .C2(n6103), .A(n6029), .B(n6209), .ZN(n5061)
         );
  INV_X1 U6272 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5068) );
  OR2_X1 U6273 ( .A1(n6022), .A2(n5116), .ZN(n6215) );
  AOI22_X1 U6274 ( .A1(n5094), .A2(n6165), .B1(n5093), .B2(n6162), .ZN(n5065)
         );
  OAI21_X1 U6275 ( .B1(n5096), .B2(n6602), .A(n5065), .ZN(n5066) );
  AOI21_X1 U6276 ( .B1(n5098), .B2(n6599), .A(n5066), .ZN(n5067) );
  OAI21_X1 U6277 ( .B1(n5101), .B2(n5068), .A(n5067), .ZN(U3100) );
  INV_X1 U6278 ( .A(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5072) );
  AOI22_X1 U6279 ( .A1(n5094), .A2(n6198), .B1(n5093), .B2(n6272), .ZN(n5069)
         );
  OAI21_X1 U6280 ( .B1(n5096), .B2(n6642), .A(n5069), .ZN(n5070) );
  AOI21_X1 U6281 ( .B1(n5098), .B2(n6637), .A(n5070), .ZN(n5071) );
  OAI21_X1 U6282 ( .B1(n5101), .B2(n5072), .A(n5071), .ZN(U3107) );
  INV_X1 U6283 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5076) );
  AOI22_X1 U6284 ( .A1(n5094), .A2(n6175), .B1(n5093), .B2(n6234), .ZN(n5073)
         );
  OAI21_X1 U6285 ( .B1(n5096), .B2(n6173), .A(n5073), .ZN(n5074) );
  AOI21_X1 U6286 ( .B1(n5098), .B2(n6119), .A(n5074), .ZN(n5075) );
  OAI21_X1 U6287 ( .B1(n5101), .B2(n5076), .A(n5075), .ZN(U3102) );
  INV_X1 U6288 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5080) );
  AOI22_X1 U6289 ( .A1(n5094), .A2(n6191), .B1(n5093), .B2(n6263), .ZN(n5077)
         );
  OAI21_X1 U6290 ( .B1(n5096), .B2(n6630), .A(n5077), .ZN(n5078) );
  AOI21_X1 U6291 ( .B1(n5098), .B2(n6627), .A(n5078), .ZN(n5079) );
  OAI21_X1 U6292 ( .B1(n5101), .B2(n5080), .A(n5079), .ZN(U3106) );
  INV_X1 U6293 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5084) );
  AOI22_X1 U6294 ( .A1(n5094), .A2(n6183), .B1(n5093), .B2(n6249), .ZN(n5081)
         );
  OAI21_X1 U6295 ( .B1(n5096), .B2(n6616), .A(n5081), .ZN(n5082) );
  AOI21_X1 U6296 ( .B1(n5098), .B2(n6613), .A(n5082), .ZN(n5083) );
  OAI21_X1 U6297 ( .B1(n5101), .B2(n5084), .A(n5083), .ZN(U3104) );
  INV_X1 U6298 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5088) );
  AOI22_X1 U6299 ( .A1(n5094), .A2(n6187), .B1(n5093), .B2(n6256), .ZN(n5085)
         );
  OAI21_X1 U6300 ( .B1(n5096), .B2(n6623), .A(n5085), .ZN(n5086) );
  AOI21_X1 U6301 ( .B1(n5098), .B2(n6620), .A(n5086), .ZN(n5087) );
  OAI21_X1 U6302 ( .B1(n5101), .B2(n5088), .A(n5087), .ZN(U3105) );
  INV_X1 U6303 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5092) );
  AOI22_X1 U6304 ( .A1(n5094), .A2(n6179), .B1(n5093), .B2(n6242), .ZN(n5089)
         );
  OAI21_X1 U6305 ( .B1(n5096), .B2(n6609), .A(n5089), .ZN(n5090) );
  AOI21_X1 U6306 ( .B1(n5098), .B2(n6606), .A(n5090), .ZN(n5091) );
  OAI21_X1 U6307 ( .B1(n5101), .B2(n5092), .A(n5091), .ZN(U3103) );
  INV_X1 U6308 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5100) );
  AOI22_X1 U6309 ( .A1(n5094), .A2(n6170), .B1(n5093), .B2(n6226), .ZN(n5095)
         );
  OAI21_X1 U6310 ( .B1(n5096), .B2(n6168), .A(n5095), .ZN(n5097) );
  AOI21_X1 U6311 ( .B1(n5098), .B2(n6114), .A(n5097), .ZN(n5099) );
  OAI21_X1 U6312 ( .B1(n5101), .B2(n5100), .A(n5099), .ZN(U3101) );
  NAND2_X1 U6313 ( .A1(n6824), .A2(n6297), .ZN(n5175) );
  OR2_X1 U6314 ( .A1(n5102), .A2(n5175), .ZN(n5173) );
  INV_X1 U6315 ( .A(n5117), .ZN(n5119) );
  INV_X1 U6316 ( .A(n5111), .ZN(n5114) );
  OAI22_X1 U6317 ( .A1(n3583), .A2(n5104), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5103), .ZN(n5271) );
  AOI21_X1 U6318 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5270), .A(n5271), 
        .ZN(n5107) );
  AOI21_X1 U6319 ( .B1(n5107), .B2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5110) );
  AOI211_X1 U6320 ( .C1(n5108), .C2(n5107), .A(n5106), .B(n5105), .ZN(n5109)
         );
  AOI211_X1 U6321 ( .C1(n5112), .C2(n5111), .A(n5110), .B(n5109), .ZN(n5113)
         );
  AOI21_X1 U6322 ( .B1(n5114), .B2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(n5113), 
        .ZN(n5115) );
  AOI21_X1 U6323 ( .B1(n5117), .B2(n5116), .A(n5115), .ZN(n5118) );
  AOI211_X1 U6324 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n5119), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n5118), .ZN(n5126) );
  OAI21_X1 U6325 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n5120), 
        .ZN(n5122) );
  NAND2_X1 U6326 ( .A1(n5122), .A2(n5121), .ZN(n5123) );
  OAI22_X1 U6327 ( .A1(n6282), .A2(n6644), .B1(n6824), .B2(n6693), .ZN(n5127)
         );
  OAI21_X1 U6328 ( .B1(n5173), .B2(n5128), .A(n5127), .ZN(n6650) );
  INV_X1 U6329 ( .A(n6650), .ZN(n5130) );
  OAI21_X1 U6330 ( .B1(n5130), .B2(n5129), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n5132) );
  NAND2_X1 U6331 ( .A1(n5132), .A2(n5131), .ZN(U3453) );
  AOI21_X1 U6332 ( .B1(n5134), .B2(n5133), .A(n3071), .ZN(n5146) );
  INV_X1 U6333 ( .A(n5146), .ZN(n5529) );
  AND2_X1 U6334 ( .A1(n5136), .A2(n5135), .ZN(n5137) );
  OR2_X1 U6335 ( .A1(n5137), .A2(n2991), .ZN(n5522) );
  INV_X1 U6336 ( .A(n5522), .ZN(n6522) );
  AOI22_X1 U6337 ( .A1(n6522), .A2(n5628), .B1(n5627), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n5138) );
  OAI21_X1 U6338 ( .B1(n5529), .B2(n5630), .A(n5138), .ZN(U2851) );
  INV_X1 U6339 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6717) );
  OAI222_X1 U6340 ( .A1(n5529), .A2(n5675), .B1(n5670), .B2(n5139), .C1(n6420), 
        .C2(n6717), .ZN(U2883) );
  OR2_X1 U6341 ( .A1(n5142), .A2(n5141), .ZN(n5143) );
  NAND2_X1 U6342 ( .A1(n5140), .A2(n5143), .ZN(n6521) );
  AOI22_X1 U6343 ( .A1(n6501), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6573), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n5144) );
  OAI21_X1 U6344 ( .B1(n6510), .B2(n2992), .A(n5144), .ZN(n5145) );
  AOI21_X1 U6345 ( .B1(n5146), .B2(n5795), .A(n5145), .ZN(n5147) );
  OAI21_X1 U6346 ( .B1(n6298), .B2(n6521), .A(n5147), .ZN(U2978) );
  INV_X1 U6347 ( .A(n5151), .ZN(n5152) );
  NAND2_X1 U6348 ( .A1(n5152), .A2(n5410), .ZN(n6647) );
  AND2_X1 U6349 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5153) );
  NAND2_X1 U6350 ( .A1(n6697), .A2(n5153), .ZN(n6288) );
  NAND2_X1 U6351 ( .A1(n3249), .A2(n5159), .ZN(n5160) );
  AOI21_X1 U6352 ( .B1(n4141), .B2(n5160), .A(n5175), .ZN(n5161) );
  INV_X1 U6353 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6663) );
  NAND2_X1 U6354 ( .A1(REIP_REG_3__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .ZN(
        n5540) );
  NOR2_X1 U6355 ( .A1(n6681), .A2(n5540), .ZN(n5544) );
  NAND3_X1 U6356 ( .A1(REIP_REG_5__SCAN_IN), .A2(REIP_REG_4__SCAN_IN), .A3(
        n5544), .ZN(n5530) );
  NOR4_X1 U6357 ( .A1(n6525), .A2(n6661), .A3(n6659), .A4(n5530), .ZN(n5517)
         );
  NAND4_X1 U6358 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5517), .A3(
        REIP_REG_10__SCAN_IN), .A4(REIP_REG_9__SCAN_IN), .ZN(n6332) );
  NOR2_X1 U6359 ( .A1(n6663), .A2(n6332), .ZN(n6335) );
  NAND2_X1 U6360 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6335), .ZN(n5181) );
  NOR2_X1 U6361 ( .A1(n6767), .A2(n5181), .ZN(n5491) );
  OR2_X1 U6362 ( .A1(n6333), .A2(n5491), .ZN(n5182) );
  AND2_X1 U6363 ( .A1(n5182), .A2(n6409), .ZN(n6316) );
  INV_X1 U6364 ( .A(n6316), .ZN(n5184) );
  INV_X1 U6365 ( .A(n5162), .ZN(n5171) );
  NAND2_X1 U6366 ( .A1(n6409), .A2(n5310), .ZN(n6365) );
  NAND2_X1 U6367 ( .A1(n5175), .A2(EBX_REG_31__SCAN_IN), .ZN(n5163) );
  NOR2_X1 U6368 ( .A1(n4141), .A2(n5163), .ZN(n5164) );
  NAND2_X1 U6369 ( .A1(n5165), .A2(n5166), .ZN(n5488) );
  OR2_X1 U6370 ( .A1(n5165), .A2(n5166), .ZN(n5167) );
  NAND2_X1 U6371 ( .A1(n5488), .A2(n5167), .ZN(n5917) );
  OAI22_X1 U6372 ( .A1(n5168), .A2(n6376), .B1(n6375), .B2(n5917), .ZN(n5169)
         );
  INV_X1 U6373 ( .A(n5169), .ZN(n5170) );
  OAI211_X1 U6374 ( .C1(n5330), .C2(n5171), .A(n6365), .B(n5170), .ZN(n5172)
         );
  INV_X1 U6375 ( .A(n5172), .ZN(n5180) );
  AND2_X1 U6376 ( .A1(n5174), .A2(n5173), .ZN(n5287) );
  INV_X1 U6377 ( .A(n5287), .ZN(n5177) );
  INV_X1 U6378 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5278) );
  NAND3_X1 U6379 ( .A1(n3249), .A2(n5278), .A3(n5175), .ZN(n5176) );
  NAND2_X1 U6380 ( .A1(n5177), .A2(n5176), .ZN(n5178) );
  NAND2_X1 U6381 ( .A1(n6398), .A2(EBX_REG_14__SCAN_IN), .ZN(n5179) );
  OAI211_X1 U6382 ( .C1(n5182), .C2(n5181), .A(n5180), .B(n5179), .ZN(n5183)
         );
  AOI21_X1 U6383 ( .B1(n5184), .B2(REIP_REG_14__SCAN_IN), .A(n5183), .ZN(n5185) );
  OAI21_X1 U6384 ( .B1(n5148), .B2(n6371), .A(n5185), .ZN(U2813) );
  INV_X1 U6385 ( .A(DATAI_14_), .ZN(n5187) );
  OAI222_X1 U6386 ( .A1(n5675), .A2(n5148), .B1(n5187), .B2(n5670), .C1(n5186), 
        .C2(n6420), .ZN(U2877) );
  INV_X1 U6387 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5188) );
  OAI222_X1 U6388 ( .A1(n5630), .A2(n5148), .B1(n5626), .B2(n5188), .C1(n5917), 
        .C2(n5624), .ZN(U2845) );
  NAND3_X1 U6389 ( .A1(n5189), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n5808), .ZN(n5191) );
  NAND2_X1 U6390 ( .A1(n5191), .A2(n5190), .ZN(n5192) );
  XNOR2_X1 U6391 ( .A(n5192), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5825)
         );
  NOR2_X1 U6392 ( .A1(n5194), .A2(n5193), .ZN(n5345) );
  NAND2_X1 U6393 ( .A1(n5345), .A2(n5195), .ZN(n5347) );
  AND2_X1 U6394 ( .A1(n5347), .A2(n5196), .ZN(n5198) );
  NOR2_X1 U6395 ( .A1(n5198), .A2(n5197), .ZN(n5202) );
  NAND2_X1 U6396 ( .A1(n6573), .A2(REIP_REG_27__SCAN_IN), .ZN(n5817) );
  NAND2_X1 U6397 ( .A1(n6501), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5199)
         );
  OAI211_X1 U6398 ( .C1(n6510), .C2(n5210), .A(n5817), .B(n5199), .ZN(n5200)
         );
  AOI21_X1 U6399 ( .B1(n5202), .B2(n5795), .A(n5200), .ZN(n5201) );
  OAI21_X1 U6400 ( .B1(n5825), .B2(n6298), .A(n5201), .ZN(U2959) );
  INV_X1 U6401 ( .A(n5202), .ZN(n5224) );
  AOI22_X1 U6402 ( .A1(n6410), .A2(DATAI_27_), .B1(n6412), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5204) );
  NAND2_X1 U6403 ( .A1(n6413), .A2(DATAI_11_), .ZN(n5203) );
  OAI211_X1 U6404 ( .C1(n5224), .C2(n5675), .A(n5204), .B(n5203), .ZN(U2864)
         );
  INV_X1 U6405 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5206) );
  OAI21_X1 U6406 ( .B1(n5342), .B2(n5205), .A(n5241), .ZN(n5819) );
  OAI222_X1 U6407 ( .A1(n5206), .A2(n5626), .B1(n5624), .B2(n5819), .C1(n5224), 
        .C2(n5630), .ZN(U2832) );
  INV_X1 U6408 ( .A(n5819), .ZN(n5222) );
  NAND3_X1 U6409 ( .A1(REIP_REG_26__SCAN_IN), .A2(REIP_REG_24__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5214) );
  NAND2_X1 U6410 ( .A1(n6333), .A2(n6409), .ZN(n5567) );
  NAND2_X1 U6411 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5491), .ZN(n5211) );
  NAND2_X1 U6412 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .ZN(
        n5212) );
  NOR2_X1 U6413 ( .A1(n5211), .A2(n5212), .ZN(n5207) );
  AND2_X1 U6414 ( .A1(n6409), .A2(n5207), .ZN(n5395) );
  AND3_X1 U6415 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n5396) );
  AND2_X1 U6416 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5208) );
  NAND4_X1 U6417 ( .A1(n5395), .A2(REIP_REG_23__SCAN_IN), .A3(n5396), .A4(
        n5208), .ZN(n5209) );
  AOI21_X1 U6418 ( .B1(n5214), .B2(n5567), .A(n5383), .ZN(n5350) );
  INV_X1 U6419 ( .A(REIP_REG_27__SCAN_IN), .ZN(n5220) );
  NOR2_X1 U6420 ( .A1(n5330), .A2(n5210), .ZN(n5218) );
  AND2_X1 U6421 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .ZN(
        n5213) );
  INV_X1 U6422 ( .A(n5214), .ZN(n5215) );
  OAI22_X1 U6423 ( .A1(n6376), .A2(n5216), .B1(REIP_REG_27__SCAN_IN), .B2(
        n5333), .ZN(n5217) );
  AOI211_X1 U6424 ( .C1(EBX_REG_27__SCAN_IN), .C2(n6398), .A(n5218), .B(n5217), 
        .ZN(n5219) );
  OAI21_X1 U6425 ( .B1(n5350), .B2(n5220), .A(n5219), .ZN(n5221) );
  AOI21_X1 U6426 ( .B1(n5222), .B2(n6399), .A(n5221), .ZN(n5223) );
  OAI21_X1 U6427 ( .B1(n5224), .B2(n6371), .A(n5223), .ZN(U2800) );
  INV_X1 U6428 ( .A(n5227), .ZN(n5225) );
  OAI21_X1 U6429 ( .B1(n5226), .B2(n5261), .A(n5225), .ZN(n5230) );
  OAI211_X1 U6430 ( .C1(n4240), .C2(n4145), .A(n5228), .B(n5227), .ZN(n5229)
         );
  OAI21_X1 U6431 ( .B1(n5231), .B2(n5230), .A(n5229), .ZN(n5572) );
  INV_X1 U6432 ( .A(n5572), .ZN(n5237) );
  NAND3_X1 U6433 ( .A1(n5254), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5232), .ZN(n5234) );
  OAI211_X1 U6434 ( .C1(n5235), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5234), .B(n5233), .ZN(n5236) );
  AOI21_X1 U6435 ( .B1(n5237), .B2(n6541), .A(n5236), .ZN(n5238) );
  OAI21_X1 U6436 ( .B1(n5239), .B2(n6520), .A(n5238), .ZN(U2988) );
  NAND2_X1 U6437 ( .A1(n5241), .A2(n5240), .ZN(n5242) );
  INV_X1 U6438 ( .A(n5243), .ZN(n5256) );
  NAND3_X1 U6439 ( .A1(n5823), .A2(n5244), .A3(n5256), .ZN(n5246) );
  OAI211_X1 U6440 ( .C1(n5818), .C2(n5247), .A(n5246), .B(n5245), .ZN(n5248)
         );
  AOI21_X1 U6441 ( .B1(n5576), .B2(n4314), .A(n5248), .ZN(n5249) );
  OAI21_X1 U6442 ( .B1(n5250), .B2(n6520), .A(n5249), .ZN(U2990) );
  INV_X1 U6443 ( .A(n4102), .ZN(n5251) );
  NAND2_X1 U6444 ( .A1(n5252), .A2(n5251), .ZN(n5253) );
  XNOR2_X1 U6445 ( .A(n5253), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5689)
         );
  INV_X1 U6446 ( .A(n5254), .ZN(n5267) );
  INV_X1 U6447 ( .A(n5823), .ZN(n5257) );
  OAI21_X1 U6448 ( .B1(n5257), .B2(n5256), .A(n5255), .ZN(n5258) );
  INV_X1 U6449 ( .A(n5258), .ZN(n5266) );
  NOR2_X1 U6450 ( .A1(n6524), .A2(n5285), .ZN(n5683) );
  INV_X1 U6451 ( .A(n5683), .ZN(n5265) );
  INV_X1 U6452 ( .A(n5259), .ZN(n5264) );
  OAI211_X1 U6453 ( .C1(n5439), .C2(n5262), .A(n5261), .B(n5260), .ZN(n5263)
         );
  INV_X1 U6454 ( .A(n5268), .ZN(n5269) );
  OAI21_X1 U6455 ( .B1(n5689), .B2(n6520), .A(n5269), .ZN(U2989) );
  INV_X1 U6456 ( .A(n6294), .ZN(n5307) );
  AOI21_X1 U6457 ( .B1(n5270), .B2(n5306), .A(n5307), .ZN(n5276) );
  INV_X1 U6458 ( .A(n5271), .ZN(n5272) );
  OAI22_X1 U6459 ( .A1(n5272), .A2(n6646), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n5301), .ZN(n5273) );
  AOI21_X1 U6460 ( .B1(n5298), .B2(n5275), .A(n5273), .ZN(n5274) );
  OAI22_X1 U6461 ( .A1(n5276), .A2(n5275), .B1(n5307), .B2(n5274), .ZN(U3461)
         );
  OAI22_X1 U6462 ( .A1(n5295), .A2(n5624), .B1(n5278), .B2(n5626), .ZN(U2828)
         );
  AOI22_X1 U6463 ( .A1(n5280), .A2(EAX_REG_31__SCAN_IN), .B1(n5279), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5283) );
  AND2_X1 U6464 ( .A1(n5324), .A2(n5281), .ZN(n5282) );
  XNOR2_X1 U6465 ( .A(n5283), .B(n5282), .ZN(n5680) );
  NAND2_X1 U6466 ( .A1(n5680), .A2(n6346), .ZN(n5294) );
  NAND2_X1 U6467 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5286) );
  INV_X1 U6468 ( .A(n5286), .ZN(n5284) );
  OAI21_X1 U6469 ( .B1(n6333), .B2(n5284), .A(n5350), .ZN(n5329) );
  OAI21_X1 U6470 ( .B1(REIP_REG_30__SCAN_IN), .B2(n6333), .A(n5319), .ZN(n5292) );
  INV_X1 U6471 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5290) );
  INV_X1 U6472 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6675) );
  NAND3_X1 U6473 ( .A1(n5316), .A2(REIP_REG_30__SCAN_IN), .A3(n6675), .ZN(
        n5289) );
  NAND3_X1 U6474 ( .A1(n5549), .A2(EBX_REG_31__SCAN_IN), .A3(n5287), .ZN(n5288) );
  OAI211_X1 U6475 ( .C1(n6376), .C2(n5290), .A(n5289), .B(n5288), .ZN(n5291)
         );
  AOI21_X1 U6476 ( .B1(n5292), .B2(REIP_REG_31__SCAN_IN), .A(n5291), .ZN(n5293) );
  OAI211_X1 U6477 ( .C1(n5295), .C2(n6375), .A(n5294), .B(n5293), .ZN(U2796)
         );
  NAND3_X1 U6478 ( .A1(n5680), .A2(n2949), .A3(n6420), .ZN(n5297) );
  AOI22_X1 U6479 ( .A1(n6410), .A2(DATAI_31_), .B1(n6412), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5296) );
  NAND2_X1 U6480 ( .A1(n5297), .A2(n5296), .ZN(U2860) );
  INV_X1 U6481 ( .A(n4538), .ZN(n5302) );
  AOI21_X1 U6482 ( .B1(n5298), .B2(n5302), .A(n5307), .ZN(n5309) );
  NOR3_X1 U6483 ( .A1(n5301), .A2(n5300), .A3(n5299), .ZN(n5304) );
  NOR3_X1 U6484 ( .A1(n6283), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n5302), 
        .ZN(n5303) );
  AOI211_X1 U6485 ( .C1(n5306), .C2(n5305), .A(n5304), .B(n5303), .ZN(n5308)
         );
  OAI22_X1 U6486 ( .A1(n5309), .A2(n3515), .B1(n5308), .B2(n5307), .ZN(U3459)
         );
  OR2_X1 U6487 ( .A1(n5310), .A2(READREQUEST_REG_SCAN_IN), .ZN(n5313) );
  INV_X1 U6488 ( .A(n5311), .ZN(n5312) );
  MUX2_X1 U6489 ( .A(n5313), .B(n5312), .S(n6695), .Z(U3474) );
  INV_X1 U6490 ( .A(n5633), .ZN(n5314) );
  NAND2_X1 U6491 ( .A1(n5314), .A2(n6346), .ZN(n5323) );
  INV_X1 U6492 ( .A(n5315), .ZN(n5318) );
  INV_X1 U6493 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6792) );
  AOI22_X1 U6494 ( .A1(n6394), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .B1(n5316), 
        .B2(n6792), .ZN(n5317) );
  OAI21_X1 U6495 ( .B1(n5318), .B2(n5330), .A(n5317), .ZN(n5321) );
  NOR2_X1 U6496 ( .A1(n5319), .A2(n6792), .ZN(n5320) );
  AOI211_X1 U6497 ( .C1(EBX_REG_30__SCAN_IN), .C2(n6398), .A(n5321), .B(n5320), 
        .ZN(n5322) );
  OAI211_X1 U6498 ( .C1(n6375), .C2(n5572), .A(n5323), .B(n5322), .ZN(U2797)
         );
  AOI21_X1 U6499 ( .B1(n5326), .B2(n5325), .A(n5324), .ZN(n5687) );
  NAND2_X1 U6500 ( .A1(n5687), .A2(n6346), .ZN(n5328) );
  OAI211_X1 U6501 ( .C1(n6375), .C2(n5574), .A(n5328), .B(n5327), .ZN(U2798)
         );
  NAND2_X1 U6502 ( .A1(n5329), .A2(REIP_REG_28__SCAN_IN), .ZN(n5338) );
  INV_X1 U6503 ( .A(REIP_REG_28__SCAN_IN), .ZN(n5331) );
  NAND2_X1 U6504 ( .A1(n5331), .A2(REIP_REG_27__SCAN_IN), .ZN(n5332) );
  OAI22_X1 U6505 ( .A1(n6376), .A2(n5334), .B1(n5333), .B2(n5332), .ZN(n5335)
         );
  AOI21_X1 U6506 ( .B1(n5336), .B2(n6397), .A(n5335), .ZN(n5337) );
  OAI211_X1 U6507 ( .C1(n5339), .C2(n6327), .A(n5338), .B(n5337), .ZN(n5340)
         );
  AOI21_X1 U6508 ( .B1(n5576), .B2(n6399), .A(n5340), .ZN(n5341) );
  OAI21_X1 U6509 ( .B1(n5639), .B2(n6371), .A(n5341), .ZN(U2799) );
  INV_X1 U6510 ( .A(n5342), .ZN(n5343) );
  OAI21_X1 U6511 ( .B1(n5363), .B2(n5344), .A(n5343), .ZN(n5833) );
  INV_X1 U6512 ( .A(n5345), .ZN(n5356) );
  INV_X1 U6513 ( .A(n5696), .ZN(n5348) );
  NAND2_X1 U6514 ( .A1(n5348), .A2(n6346), .ZN(n5355) );
  INV_X1 U6515 ( .A(n5693), .ZN(n5349) );
  OAI22_X1 U6516 ( .A1(n6376), .A2(n3022), .B1(n5349), .B2(n5330), .ZN(n5353)
         );
  NAND3_X1 U6517 ( .A1(n5369), .A2(REIP_REG_24__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5351) );
  AOI21_X1 U6518 ( .B1(n6799), .B2(n5351), .A(n5350), .ZN(n5352) );
  AOI211_X1 U6519 ( .C1(n6398), .C2(EBX_REG_26__SCAN_IN), .A(n5353), .B(n5352), 
        .ZN(n5354) );
  OAI211_X1 U6520 ( .C1(n6375), .C2(n5833), .A(n5355), .B(n5354), .ZN(U2801)
         );
  OAI21_X1 U6521 ( .B1(n5358), .B2(n5357), .A(n5356), .ZN(n5704) );
  NAND2_X1 U6522 ( .A1(n6398), .A2(EBX_REG_25__SCAN_IN), .ZN(n5361) );
  XOR2_X1 U6523 ( .A(REIP_REG_24__SCAN_IN), .B(REIP_REG_25__SCAN_IN), .Z(n5359) );
  AOI22_X1 U6524 ( .A1(n6394), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .B1(n5369), 
        .B2(n5359), .ZN(n5360) );
  OAI211_X1 U6525 ( .C1(n5330), .C2(n5700), .A(n5361), .B(n5360), .ZN(n5366)
         );
  AND2_X1 U6526 ( .A1(n5374), .A2(n5362), .ZN(n5364) );
  OR2_X1 U6527 ( .A1(n5364), .A2(n5363), .ZN(n5841) );
  NOR2_X1 U6528 ( .A1(n5841), .A2(n6375), .ZN(n5365) );
  AOI211_X1 U6529 ( .C1(n5383), .C2(REIP_REG_25__SCAN_IN), .A(n5366), .B(n5365), .ZN(n5367) );
  OAI21_X1 U6530 ( .B1(n5704), .B2(n6371), .A(n5367), .ZN(U2802) );
  INV_X1 U6531 ( .A(n5368), .ZN(n5372) );
  NAND2_X1 U6532 ( .A1(n6398), .A2(EBX_REG_24__SCAN_IN), .ZN(n5371) );
  AOI22_X1 U6533 ( .A1(n6394), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .B1(n5369), 
        .B2(n6800), .ZN(n5370) );
  OAI211_X1 U6534 ( .C1(n5330), .C2(n5372), .A(n5371), .B(n5370), .ZN(n5373)
         );
  AOI21_X1 U6535 ( .B1(REIP_REG_24__SCAN_IN), .B2(n5383), .A(n5373), .ZN(n5379) );
  INV_X1 U6536 ( .A(n5374), .ZN(n5375) );
  AOI21_X1 U6537 ( .B1(n5377), .B2(n5376), .A(n5375), .ZN(n5850) );
  NAND2_X1 U6538 ( .A1(n5850), .A2(n6399), .ZN(n5378) );
  OAI211_X1 U6539 ( .C1(n5646), .C2(n6371), .A(n5379), .B(n5378), .ZN(U2803)
         );
  INV_X1 U6540 ( .A(n5649), .ZN(n5380) );
  NAND2_X1 U6541 ( .A1(n5380), .A2(n6346), .ZN(n5389) );
  OAI22_X1 U6542 ( .A1(n6376), .A2(n5382), .B1(n5381), .B2(n5330), .ZN(n5387)
         );
  INV_X1 U6543 ( .A(n5383), .ZN(n5385) );
  AOI21_X1 U6544 ( .B1(n5392), .B2(REIP_REG_22__SCAN_IN), .A(
        REIP_REG_23__SCAN_IN), .ZN(n5384) );
  NOR2_X1 U6545 ( .A1(n5385), .A2(n5384), .ZN(n5386) );
  AOI211_X1 U6546 ( .C1(n6398), .C2(EBX_REG_23__SCAN_IN), .A(n5387), .B(n5386), 
        .ZN(n5388) );
  OAI211_X1 U6547 ( .C1(n6375), .C2(n5581), .A(n5389), .B(n5388), .ZN(U2804)
         );
  INV_X1 U6548 ( .A(n5652), .ZN(n5390) );
  NAND2_X1 U6549 ( .A1(n5390), .A2(n6346), .ZN(n5401) );
  INV_X1 U6550 ( .A(n5391), .ZN(n5394) );
  AOI22_X1 U6551 ( .A1(n6394), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .B1(n5392), 
        .B2(n6704), .ZN(n5393) );
  OAI21_X1 U6552 ( .B1(n5394), .B2(n5330), .A(n5393), .ZN(n5399) );
  INV_X1 U6553 ( .A(n5395), .ZN(n5444) );
  INV_X1 U6554 ( .A(n5396), .ZN(n5397) );
  OAI21_X1 U6555 ( .B1(n5444), .B2(n5397), .A(n5567), .ZN(n5428) );
  NAND3_X1 U6556 ( .A1(n6670), .A2(REIP_REG_20__SCAN_IN), .A3(n5430), .ZN(
        n5419) );
  AOI21_X1 U6557 ( .B1(n5428), .B2(n5419), .A(n6704), .ZN(n5398) );
  AOI211_X1 U6558 ( .C1(EBX_REG_22__SCAN_IN), .C2(n6398), .A(n5399), .B(n5398), 
        .ZN(n5400) );
  OAI211_X1 U6559 ( .C1(n6375), .C2(n5583), .A(n5401), .B(n5400), .ZN(U2805)
         );
  AND2_X2 U6560 ( .A1(n5403), .A2(n5402), .ZN(n5594) );
  INV_X1 U6561 ( .A(n5594), .ZN(n5406) );
  INV_X1 U6562 ( .A(n5476), .ZN(n5751) );
  NAND2_X1 U6563 ( .A1(n5751), .A2(n3063), .ZN(n5404) );
  OAI21_X1 U6564 ( .B1(n5405), .B2(n3063), .A(n5404), .ZN(n5465) );
  NOR2_X2 U6565 ( .A1(n5406), .A2(n5465), .ZN(n5466) );
  MUX2_X1 U6566 ( .A(n5407), .B(n5735), .S(n5410), .Z(n5453) );
  NAND2_X1 U6567 ( .A1(n5466), .A2(n5453), .ZN(n5452) );
  INV_X1 U6568 ( .A(n5724), .ZN(n5408) );
  NAND2_X1 U6569 ( .A1(n5408), .A2(n5410), .ZN(n5409) );
  OAI21_X1 U6570 ( .B1(n5411), .B2(n5410), .A(n5409), .ZN(n5436) );
  NOR2_X2 U6571 ( .A1(n5452), .A2(n5436), .ZN(n5713) );
  MUX2_X1 U6572 ( .A(n5716), .B(n5413), .S(n5412), .Z(n5714) );
  NAND2_X1 U6573 ( .A1(n5713), .A2(n5714), .ZN(n5416) );
  AOI21_X2 U6574 ( .B1(n5416), .B2(n5415), .A(n5414), .ZN(n5710) );
  INV_X1 U6575 ( .A(n5710), .ZN(n5655) );
  XOR2_X1 U6576 ( .A(n5418), .B(n5417), .Z(n5858) );
  NAND2_X1 U6577 ( .A1(n6394), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5420)
         );
  OAI211_X1 U6578 ( .C1(n5330), .C2(n5708), .A(n5420), .B(n5419), .ZN(n5421)
         );
  AOI21_X1 U6579 ( .B1(n6398), .B2(EBX_REG_21__SCAN_IN), .A(n5421), .ZN(n5422)
         );
  OAI21_X1 U6580 ( .B1(n5428), .B2(n6670), .A(n5422), .ZN(n5423) );
  AOI21_X1 U6581 ( .B1(n5858), .B2(n6399), .A(n5423), .ZN(n5424) );
  OAI21_X1 U6582 ( .B1(n5655), .B2(n6371), .A(n5424), .ZN(U2806) );
  XNOR2_X1 U6583 ( .A(n5714), .B(n5713), .ZN(n5658) );
  MUX2_X1 U6584 ( .A(n5441), .B(n4145), .S(n5425), .Z(n5427) );
  XNOR2_X1 U6585 ( .A(n5427), .B(n5426), .ZN(n5866) );
  INV_X1 U6586 ( .A(n5428), .ZN(n5429) );
  OAI21_X1 U6587 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5430), .A(n5429), .ZN(n5433) );
  INV_X1 U6588 ( .A(n5716), .ZN(n5431) );
  AOI22_X1 U6589 ( .A1(n6397), .A2(n5431), .B1(n6394), .B2(
        PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5432) );
  OAI211_X1 U6590 ( .C1(n6327), .C2(n5587), .A(n5433), .B(n5432), .ZN(n5434)
         );
  AOI21_X1 U6591 ( .B1(n5866), .B2(n6399), .A(n5434), .ZN(n5435) );
  OAI21_X1 U6592 ( .B1(n5658), .B2(n6371), .A(n5435), .ZN(U2807) );
  AOI21_X1 U6593 ( .B1(n5436), .B2(n5452), .A(n5713), .ZN(n5726) );
  INV_X1 U6594 ( .A(n5726), .ZN(n5661) );
  NAND2_X1 U6595 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5437) );
  OAI211_X1 U6596 ( .C1(REIP_REG_19__SCAN_IN), .C2(REIP_REG_18__SCAN_IN), .A(
        n5460), .B(n5437), .ZN(n5451) );
  MUX2_X1 U6597 ( .A(n5441), .B(n5440), .S(n5439), .Z(n5456) );
  INV_X1 U6598 ( .A(n5456), .ZN(n5442) );
  NAND2_X1 U6599 ( .A1(n5472), .A2(n5442), .ZN(n5454) );
  XNOR2_X1 U6600 ( .A(n5454), .B(n5443), .ZN(n5875) );
  INV_X1 U6601 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5448) );
  NAND2_X1 U6602 ( .A1(n5567), .A2(n5444), .ZN(n5479) );
  NAND2_X1 U6603 ( .A1(n6394), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5445)
         );
  OAI211_X1 U6604 ( .C1(n5330), .C2(n5724), .A(n5445), .B(n6365), .ZN(n5446)
         );
  AOI21_X1 U6605 ( .B1(n6398), .B2(EBX_REG_19__SCAN_IN), .A(n5446), .ZN(n5447)
         );
  OAI21_X1 U6606 ( .B1(n5448), .B2(n5479), .A(n5447), .ZN(n5449) );
  AOI21_X1 U6607 ( .B1(n5875), .B2(n6399), .A(n5449), .ZN(n5450) );
  OAI211_X1 U6608 ( .C1(n5661), .C2(n6371), .A(n5451), .B(n5450), .ZN(U2808)
         );
  OAI21_X1 U6609 ( .B1(n5466), .B2(n5453), .A(n5452), .ZN(n5732) );
  INV_X1 U6610 ( .A(n5472), .ZN(n5457) );
  INV_X1 U6611 ( .A(n5454), .ZN(n5455) );
  AOI21_X1 U6612 ( .B1(n5457), .B2(n5456), .A(n5455), .ZN(n5879) );
  INV_X1 U6613 ( .A(REIP_REG_18__SCAN_IN), .ZN(n5733) );
  AOI21_X1 U6614 ( .B1(n6394), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6378), 
        .ZN(n5458) );
  OAI21_X1 U6615 ( .B1(n5735), .B2(n5330), .A(n5458), .ZN(n5459) );
  AOI21_X1 U6616 ( .B1(EBX_REG_18__SCAN_IN), .B2(n6398), .A(n5459), .ZN(n5462)
         );
  NAND2_X1 U6617 ( .A1(n5460), .A2(n5733), .ZN(n5461) );
  OAI211_X1 U6618 ( .C1(n5479), .C2(n5733), .A(n5462), .B(n5461), .ZN(n5463)
         );
  AOI21_X1 U6619 ( .B1(n5879), .B2(n6399), .A(n5463), .ZN(n5464) );
  OAI21_X1 U6620 ( .B1(n5732), .B2(n6371), .A(n5464), .ZN(U2809) );
  INV_X1 U6621 ( .A(n5465), .ZN(n5468) );
  INV_X1 U6622 ( .A(n5466), .ZN(n5467) );
  NAND2_X1 U6623 ( .A1(n5165), .A2(n5469), .ZN(n5597) );
  INV_X1 U6624 ( .A(n5597), .ZN(n5471) );
  AOI21_X1 U6625 ( .B1(n5471), .B2(n5595), .A(n5470), .ZN(n5473) );
  NOR2_X1 U6626 ( .A1(n5473), .A2(n5472), .ZN(n5887) );
  INV_X1 U6627 ( .A(n6319), .ZN(n5474) );
  AOI21_X1 U6628 ( .B1(n5474), .B2(REIP_REG_16__SCAN_IN), .A(
        REIP_REG_17__SCAN_IN), .ZN(n5480) );
  AOI21_X1 U6629 ( .B1(n6394), .B2(PHYADDRPOINTER_REG_17__SCAN_IN), .A(n6378), 
        .ZN(n5475) );
  OAI21_X1 U6630 ( .B1(n5476), .B2(n5330), .A(n5475), .ZN(n5477) );
  AOI21_X1 U6631 ( .B1(n6398), .B2(EBX_REG_17__SCAN_IN), .A(n5477), .ZN(n5478)
         );
  OAI21_X1 U6632 ( .B1(n5480), .B2(n5479), .A(n5478), .ZN(n5481) );
  AOI21_X1 U6633 ( .B1(n5887), .B2(n6399), .A(n5481), .ZN(n5482) );
  OAI21_X1 U6634 ( .B1(n5754), .B2(n6371), .A(n5482), .ZN(U2810) );
  INV_X1 U6635 ( .A(n5483), .ZN(n5485) );
  NOR2_X1 U6636 ( .A1(n5610), .A2(n5484), .ZN(n5592) );
  AOI21_X1 U6637 ( .B1(n5486), .B2(n5485), .A(n5592), .ZN(n5775) );
  INV_X1 U6638 ( .A(n5775), .ZN(n5667) );
  NAND2_X1 U6639 ( .A1(n5488), .A2(n5487), .ZN(n5489) );
  AND2_X1 U6640 ( .A1(n5597), .A2(n5489), .ZN(n5910) );
  OAI22_X1 U6641 ( .A1(n6316), .A2(n5490), .B1(n5773), .B2(n5330), .ZN(n5495)
         );
  AOI21_X1 U6642 ( .B1(n6394), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6378), 
        .ZN(n5493) );
  INV_X1 U6643 ( .A(n6333), .ZN(n6384) );
  NAND3_X1 U6644 ( .A1(n6384), .A2(n5491), .A3(n5490), .ZN(n5492) );
  OAI211_X1 U6645 ( .C1(n6327), .C2(n6793), .A(n5493), .B(n5492), .ZN(n5494)
         );
  AOI211_X1 U6646 ( .C1(n5910), .C2(n6399), .A(n5495), .B(n5494), .ZN(n5496)
         );
  OAI21_X1 U6647 ( .B1(n5667), .B2(n6371), .A(n5496), .ZN(U2812) );
  OAI21_X1 U6648 ( .B1(n3890), .B2(n5497), .A(n5610), .ZN(n5672) );
  INV_X1 U6649 ( .A(n5672), .ZN(n5796) );
  INV_X1 U6650 ( .A(n6332), .ZN(n5498) );
  OR2_X1 U6651 ( .A1(n6333), .A2(n5498), .ZN(n5499) );
  AND2_X1 U6652 ( .A1(n5499), .A2(n6409), .ZN(n6340) );
  INV_X1 U6653 ( .A(n6340), .ZN(n6334) );
  AOI22_X1 U6654 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n6394), .B1(
        REIP_REG_11__SCAN_IN), .B2(n6334), .ZN(n5500) );
  OAI21_X1 U6655 ( .B1(n5615), .B2(n6327), .A(n5500), .ZN(n5508) );
  NAND2_X1 U6656 ( .A1(n5623), .A2(n5502), .ZN(n5503) );
  NAND2_X1 U6657 ( .A1(n5501), .A2(n5503), .ZN(n5950) );
  INV_X1 U6658 ( .A(n5793), .ZN(n5505) );
  NAND2_X1 U6659 ( .A1(n6384), .A2(n5517), .ZN(n6351) );
  NOR4_X1 U6660 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5965), .A3(n5810), .A4(n6351), .ZN(n5504) );
  AOI211_X1 U6661 ( .C1(n6397), .C2(n5505), .A(n5504), .B(n6378), .ZN(n5506)
         );
  OAI21_X1 U6662 ( .B1(n6375), .B2(n5950), .A(n5506), .ZN(n5507) );
  AOI211_X1 U6663 ( .C1(n5796), .C2(n6346), .A(n5508), .B(n5507), .ZN(n5509)
         );
  INV_X1 U6664 ( .A(n5509), .ZN(U2816) );
  AND2_X1 U6665 ( .A1(n5511), .A2(n5510), .ZN(n5513) );
  OR2_X1 U6666 ( .A1(n5513), .A2(n5512), .ZN(n5815) );
  INV_X1 U6667 ( .A(n2991), .ZN(n5515) );
  AOI21_X1 U6668 ( .B1(n5515), .B2(n2993), .A(n5514), .ZN(n6513) );
  NOR2_X1 U6669 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6351), .ZN(n6357) );
  INV_X1 U6670 ( .A(n6357), .ZN(n5516) );
  OAI211_X1 U6671 ( .C1(n5330), .C2(n5811), .A(n6365), .B(n5516), .ZN(n5520)
         );
  OAI21_X1 U6672 ( .B1(n6333), .B2(n5517), .A(n6409), .ZN(n6356) );
  AOI22_X1 U6673 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n6394), .B1(
        REIP_REG_9__SCAN_IN), .B2(n6356), .ZN(n5518) );
  OAI21_X1 U6674 ( .B1(n6818), .B2(n6327), .A(n5518), .ZN(n5519) );
  AOI211_X1 U6675 ( .C1(n6513), .C2(n6399), .A(n5520), .B(n5519), .ZN(n5521)
         );
  OAI21_X1 U6676 ( .B1(n6371), .B2(n5815), .A(n5521), .ZN(U2818) );
  OAI22_X1 U6677 ( .A1(n6376), .A2(n3631), .B1(n5330), .B2(n2992), .ZN(n5525)
         );
  OAI22_X1 U6678 ( .A1(n5523), .A2(n6327), .B1(n6375), .B2(n5522), .ZN(n5524)
         );
  NOR3_X1 U6679 ( .A1(n5525), .A2(n6378), .A3(n5524), .ZN(n5528) );
  NOR2_X1 U6680 ( .A1(n6333), .A2(n5530), .ZN(n5533) );
  NAND2_X1 U6681 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5533), .ZN(n6362) );
  OAI21_X1 U6682 ( .B1(n6661), .B2(n6362), .A(n6525), .ZN(n5526) );
  NAND2_X1 U6683 ( .A1(n5526), .A2(n6356), .ZN(n5527) );
  OAI211_X1 U6684 ( .C1(n5529), .C2(n6371), .A(n5528), .B(n5527), .ZN(U2819)
         );
  OAI21_X1 U6685 ( .B1(n3033), .B2(n5530), .A(n5567), .ZN(n6383) );
  OAI22_X1 U6686 ( .A1(n6383), .A2(n6659), .B1(n5531), .B2(n6327), .ZN(n5532)
         );
  AOI211_X1 U6687 ( .C1(n6394), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6378), 
        .B(n5532), .ZN(n5534) );
  NAND2_X1 U6688 ( .A1(n5533), .A2(n6659), .ZN(n6364) );
  OAI211_X1 U6689 ( .C1(n5535), .C2(n6375), .A(n5534), .B(n6364), .ZN(n5539)
         );
  OAI22_X1 U6690 ( .A1(n5537), .A2(n6371), .B1(n5536), .B2(n5330), .ZN(n5538)
         );
  OR2_X1 U6691 ( .A1(n5539), .A2(n5538), .ZN(U2821) );
  NOR3_X1 U6692 ( .A1(n6333), .A2(n6681), .A3(n5540), .ZN(n6374) );
  AOI22_X1 U6693 ( .A1(n6399), .A2(n6553), .B1(n6374), .B2(n6657), .ZN(n5541)
         );
  OAI211_X1 U6694 ( .C1(n6376), .C2(n6783), .A(n5541), .B(n6365), .ZN(n5555)
         );
  INV_X1 U6695 ( .A(n5542), .ZN(n5543) );
  NAND2_X1 U6696 ( .A1(n5549), .A2(n5543), .ZN(n6389) );
  OR2_X1 U6697 ( .A1(n6333), .A2(n5544), .ZN(n5545) );
  NAND2_X1 U6698 ( .A1(n5545), .A2(n6409), .ZN(n5556) );
  AOI22_X1 U6699 ( .A1(EBX_REG_4__SCAN_IN), .A2(n6398), .B1(
        REIP_REG_4__SCAN_IN), .B2(n5556), .ZN(n5546) );
  OAI21_X1 U6700 ( .B1(n5547), .B2(n6389), .A(n5546), .ZN(n5554) );
  NAND2_X1 U6701 ( .A1(n5549), .A2(n5548), .ZN(n5550) );
  OAI22_X1 U6702 ( .A1(n5552), .A2(n6404), .B1(n5551), .B2(n5330), .ZN(n5553)
         );
  OR3_X1 U6703 ( .A1(n5555), .A2(n5554), .A3(n5553), .ZN(U2823) );
  INV_X1 U6704 ( .A(n6404), .ZN(n6392) );
  OR2_X1 U6705 ( .A1(n6333), .A2(REIP_REG_1__SCAN_IN), .ZN(n6396) );
  AND3_X1 U6706 ( .A1(n6396), .A2(n6409), .A3(REIP_REG_2__SCAN_IN), .ZN(n6385)
         );
  OAI21_X1 U6707 ( .B1(n6385), .B2(REIP_REG_3__SCAN_IN), .A(n5556), .ZN(n5562)
         );
  INV_X1 U6708 ( .A(n6500), .ZN(n5557) );
  AOI22_X1 U6709 ( .A1(n6397), .A2(n5557), .B1(n6394), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5561) );
  INV_X1 U6710 ( .A(n6389), .ZN(n6401) );
  INV_X1 U6711 ( .A(n5558), .ZN(n6563) );
  AOI22_X1 U6712 ( .A1(n6401), .A2(n6218), .B1(n6399), .B2(n6563), .ZN(n5560)
         );
  NAND2_X1 U6713 ( .A1(n6398), .A2(EBX_REG_3__SCAN_IN), .ZN(n5559) );
  NAND4_X1 U6714 ( .A1(n5562), .A2(n5561), .A3(n5560), .A4(n5559), .ZN(n5563)
         );
  AOI21_X1 U6715 ( .B1(n6497), .B2(n6392), .A(n5563), .ZN(n5564) );
  INV_X1 U6716 ( .A(n5564), .ZN(U2824) );
  OAI22_X1 U6717 ( .A1(n6375), .A2(n5565), .B1(n3583), .B2(n6389), .ZN(n5566)
         );
  AOI21_X1 U6718 ( .B1(REIP_REG_0__SCAN_IN), .B2(n5567), .A(n5566), .ZN(n5570)
         );
  NAND2_X1 U6719 ( .A1(n6376), .A2(n5330), .ZN(n5568) );
  AOI22_X1 U6720 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n5568), .B1(n6398), 
        .B2(EBX_REG_0__SCAN_IN), .ZN(n5569) );
  OAI211_X1 U6721 ( .C1(n6404), .C2(n5571), .A(n5570), .B(n5569), .ZN(U2827)
         );
  INV_X1 U6722 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5573) );
  OAI222_X1 U6723 ( .A1(n5630), .A2(n5633), .B1(n5626), .B2(n5573), .C1(n5572), 
        .C2(n5624), .ZN(U2829) );
  INV_X1 U6724 ( .A(n5687), .ZN(n5636) );
  OAI222_X1 U6725 ( .A1(n5575), .A2(n5626), .B1(n5624), .B2(n5574), .C1(n5636), 
        .C2(n5630), .ZN(U2830) );
  AOI22_X1 U6726 ( .A1(n5576), .A2(n5628), .B1(n5627), .B2(EBX_REG_28__SCAN_IN), .ZN(n5577) );
  OAI21_X1 U6727 ( .B1(n5639), .B2(n5630), .A(n5577), .ZN(U2831) );
  OAI222_X1 U6728 ( .A1(n5578), .A2(n5626), .B1(n5624), .B2(n5833), .C1(n5696), 
        .C2(n5630), .ZN(U2833) );
  OAI222_X1 U6729 ( .A1(n5579), .A2(n5626), .B1(n5624), .B2(n5841), .C1(n5704), 
        .C2(n5630), .ZN(U2834) );
  AOI22_X1 U6730 ( .A1(n5850), .A2(n5628), .B1(n5627), .B2(EBX_REG_24__SCAN_IN), .ZN(n5580) );
  OAI21_X1 U6731 ( .B1(n5646), .B2(n5630), .A(n5580), .ZN(U2835) );
  OAI222_X1 U6732 ( .A1(n5582), .A2(n5626), .B1(n5624), .B2(n5581), .C1(n5649), 
        .C2(n5630), .ZN(U2836) );
  INV_X1 U6733 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5584) );
  OAI222_X1 U6734 ( .A1(n5584), .A2(n5626), .B1(n5624), .B2(n5583), .C1(n5652), 
        .C2(n5630), .ZN(U2837) );
  AOI22_X1 U6735 ( .A1(n5858), .A2(n5628), .B1(n5627), .B2(EBX_REG_21__SCAN_IN), .ZN(n5585) );
  OAI21_X1 U6736 ( .B1(n5655), .B2(n5630), .A(n5585), .ZN(U2838) );
  INV_X1 U6737 ( .A(n5866), .ZN(n5586) );
  OAI222_X1 U6738 ( .A1(n5630), .A2(n5658), .B1(n5626), .B2(n5587), .C1(n5586), 
        .C2(n5624), .ZN(U2839) );
  AOI22_X1 U6739 ( .A1(n5875), .A2(n5628), .B1(EBX_REG_19__SCAN_IN), .B2(n5627), .ZN(n5588) );
  OAI21_X1 U6740 ( .B1(n5661), .B2(n5630), .A(n5588), .ZN(U2840) );
  INV_X1 U6741 ( .A(n5879), .ZN(n5589) );
  OAI222_X1 U6742 ( .A1(n5630), .A2(n5732), .B1(n5626), .B2(n4211), .C1(n5589), 
        .C2(n5624), .ZN(U2841) );
  AOI22_X1 U6743 ( .A1(n5887), .A2(n5628), .B1(n5627), .B2(EBX_REG_17__SCAN_IN), .ZN(n5590) );
  OAI21_X1 U6744 ( .B1(n5754), .B2(n5630), .A(n5590), .ZN(U2842) );
  NOR2_X1 U6745 ( .A1(n5592), .A2(n5591), .ZN(n5593) );
  INV_X1 U6746 ( .A(n5595), .ZN(n5596) );
  XNOR2_X1 U6747 ( .A(n5597), .B(n5596), .ZN(n6325) );
  INV_X1 U6748 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5598) );
  OAI222_X1 U6749 ( .A1(n6321), .A2(n5630), .B1(n5624), .B2(n6325), .C1(n5626), 
        .C2(n5598), .ZN(U2843) );
  NOR2_X1 U6750 ( .A1(n5626), .A2(n6793), .ZN(n5599) );
  AOI21_X1 U6751 ( .B1(n5910), .B2(n5628), .A(n5599), .ZN(n5600) );
  OAI21_X1 U6752 ( .B1(n5667), .B2(n5630), .A(n5600), .ZN(U2844) );
  XNOR2_X1 U6753 ( .A(n5602), .B(n5601), .ZN(n6331) );
  NOR2_X1 U6754 ( .A1(n5603), .A2(n5604), .ZN(n5605) );
  OR2_X1 U6755 ( .A1(n5165), .A2(n5605), .ZN(n6326) );
  OAI22_X1 U6756 ( .A1(n6326), .A2(n5624), .B1(n6794), .B2(n5626), .ZN(n5606)
         );
  AOI21_X1 U6757 ( .B1(n6331), .B2(n5617), .A(n5606), .ZN(n5607) );
  INV_X1 U6758 ( .A(n5607), .ZN(U2846) );
  INV_X1 U6759 ( .A(n5608), .ZN(n5609) );
  AOI21_X1 U6760 ( .B1(n5611), .B2(n5610), .A(n5609), .ZN(n6418) );
  INV_X1 U6761 ( .A(n6418), .ZN(n5614) );
  AOI21_X1 U6762 ( .B1(n5612), .B2(n5501), .A(n5603), .ZN(n6343) );
  AOI22_X1 U6763 ( .A1(n6343), .A2(n5628), .B1(EBX_REG_12__SCAN_IN), .B2(n5627), .ZN(n5613) );
  OAI21_X1 U6764 ( .B1(n5614), .B2(n5630), .A(n5613), .ZN(U2847) );
  OAI22_X1 U6765 ( .A1(n5950), .A2(n5624), .B1(n5615), .B2(n5626), .ZN(n5616)
         );
  AOI21_X1 U6766 ( .B1(n5796), .B2(n5617), .A(n5616), .ZN(n5618) );
  INV_X1 U6767 ( .A(n5618), .ZN(U2848) );
  NOR2_X1 U6768 ( .A1(n5512), .A2(n5619), .ZN(n5620) );
  OR2_X1 U6769 ( .A1(n3890), .A2(n5620), .ZN(n6354) );
  INV_X1 U6770 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5625) );
  OR2_X1 U6771 ( .A1(n5514), .A2(n5621), .ZN(n5622) );
  AND2_X1 U6772 ( .A1(n5623), .A2(n5622), .ZN(n6350) );
  INV_X1 U6773 ( .A(n6350), .ZN(n5967) );
  OAI222_X1 U6774 ( .A1(n6354), .A2(n5630), .B1(n5626), .B2(n5625), .C1(n5624), 
        .C2(n5967), .ZN(U2849) );
  AOI22_X1 U6775 ( .A1(n6513), .A2(n5628), .B1(n5627), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n5629) );
  OAI21_X1 U6776 ( .B1(n5815), .B2(n5630), .A(n5629), .ZN(U2850) );
  AOI22_X1 U6777 ( .A1(n6410), .A2(DATAI_30_), .B1(n6412), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U6778 ( .A1(n6413), .A2(DATAI_14_), .ZN(n5631) );
  OAI211_X1 U6779 ( .C1(n5633), .C2(n5675), .A(n5632), .B(n5631), .ZN(U2861)
         );
  AOI22_X1 U6780 ( .A1(n6410), .A2(DATAI_29_), .B1(n6412), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U6781 ( .A1(n6413), .A2(DATAI_13_), .ZN(n5634) );
  OAI211_X1 U6782 ( .C1(n5636), .C2(n5675), .A(n5635), .B(n5634), .ZN(U2862)
         );
  AOI22_X1 U6783 ( .A1(n6410), .A2(DATAI_28_), .B1(n6412), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U6784 ( .A1(n6413), .A2(DATAI_12_), .ZN(n5637) );
  OAI211_X1 U6785 ( .C1(n5639), .C2(n5675), .A(n5638), .B(n5637), .ZN(U2863)
         );
  AOI22_X1 U6786 ( .A1(n6410), .A2(DATAI_26_), .B1(n6412), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U6787 ( .A1(n6413), .A2(DATAI_10_), .ZN(n5640) );
  OAI211_X1 U6788 ( .C1(n5696), .C2(n5675), .A(n5641), .B(n5640), .ZN(U2865)
         );
  AOI22_X1 U6789 ( .A1(n6410), .A2(DATAI_25_), .B1(n6412), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5643) );
  NAND2_X1 U6790 ( .A1(n6413), .A2(DATAI_9_), .ZN(n5642) );
  OAI211_X1 U6791 ( .C1(n5704), .C2(n5675), .A(n5643), .B(n5642), .ZN(U2866)
         );
  AOI22_X1 U6792 ( .A1(n6410), .A2(DATAI_24_), .B1(n6412), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U6793 ( .A1(n6413), .A2(DATAI_8_), .ZN(n5644) );
  OAI211_X1 U6794 ( .C1(n5646), .C2(n5675), .A(n5645), .B(n5644), .ZN(U2867)
         );
  AOI22_X1 U6795 ( .A1(n6410), .A2(DATAI_23_), .B1(n6412), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U6796 ( .A1(n6413), .A2(DATAI_7_), .ZN(n5647) );
  OAI211_X1 U6797 ( .C1(n5649), .C2(n5675), .A(n5648), .B(n5647), .ZN(U2868)
         );
  AOI22_X1 U6798 ( .A1(n6410), .A2(DATAI_22_), .B1(n6412), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5651) );
  NAND2_X1 U6799 ( .A1(n6413), .A2(DATAI_6_), .ZN(n5650) );
  OAI211_X1 U6800 ( .C1(n5652), .C2(n5675), .A(n5651), .B(n5650), .ZN(U2869)
         );
  AOI22_X1 U6801 ( .A1(n6410), .A2(DATAI_21_), .B1(n6412), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U6802 ( .A1(n6413), .A2(DATAI_5_), .ZN(n5653) );
  OAI211_X1 U6803 ( .C1(n5655), .C2(n5675), .A(n5654), .B(n5653), .ZN(U2870)
         );
  AOI22_X1 U6804 ( .A1(n6410), .A2(DATAI_20_), .B1(n6412), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U6805 ( .A1(n6413), .A2(DATAI_4_), .ZN(n5656) );
  OAI211_X1 U6806 ( .C1(n5658), .C2(n5675), .A(n5657), .B(n5656), .ZN(U2871)
         );
  AOI22_X1 U6807 ( .A1(n6410), .A2(DATAI_19_), .B1(n6412), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5660) );
  NAND2_X1 U6808 ( .A1(n6413), .A2(DATAI_3_), .ZN(n5659) );
  OAI211_X1 U6809 ( .C1(n5661), .C2(n5675), .A(n5660), .B(n5659), .ZN(U2872)
         );
  AOI22_X1 U6810 ( .A1(n6410), .A2(DATAI_18_), .B1(n6412), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U6811 ( .A1(n6413), .A2(DATAI_2_), .ZN(n5662) );
  OAI211_X1 U6812 ( .C1(n5732), .C2(n5675), .A(n5663), .B(n5662), .ZN(U2873)
         );
  AOI22_X1 U6813 ( .A1(n6410), .A2(DATAI_17_), .B1(n6412), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U6814 ( .A1(n6413), .A2(DATAI_1_), .ZN(n5664) );
  OAI211_X1 U6815 ( .C1(n5754), .C2(n5675), .A(n5665), .B(n5664), .ZN(U2874)
         );
  AOI22_X1 U6816 ( .A1(n6416), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n6412), .ZN(n5666) );
  OAI21_X1 U6817 ( .B1(n5667), .B2(n5675), .A(n5666), .ZN(U2876) );
  INV_X1 U6818 ( .A(n6331), .ZN(n5668) );
  OAI222_X1 U6819 ( .A1(n6420), .A2(n6425), .B1(n5670), .B2(n5669), .C1(n5675), 
        .C2(n5668), .ZN(U2878) );
  AOI22_X1 U6820 ( .A1(n6416), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n6412), .ZN(n5671) );
  OAI21_X1 U6821 ( .B1(n5672), .B2(n5675), .A(n5671), .ZN(U2880) );
  AOI22_X1 U6822 ( .A1(n6416), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n6412), .ZN(n5673) );
  OAI21_X1 U6823 ( .B1(n6354), .B2(n5675), .A(n5673), .ZN(U2881) );
  AOI22_X1 U6824 ( .A1(n6416), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n6412), .ZN(n5674) );
  OAI21_X1 U6825 ( .B1(n5815), .B2(n5675), .A(n5674), .ZN(U2882) );
  NAND2_X1 U6826 ( .A1(n6501), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5676)
         );
  OAI211_X1 U6827 ( .C1(n6510), .C2(n5678), .A(n5677), .B(n5676), .ZN(n5679)
         );
  AOI21_X1 U6828 ( .B1(n5680), .B2(n5795), .A(n5679), .ZN(n5681) );
  OAI21_X1 U6829 ( .B1(n5682), .B2(n6298), .A(n5681), .ZN(U2955) );
  AOI21_X1 U6830 ( .B1(n6501), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5683), 
        .ZN(n5684) );
  OAI21_X1 U6831 ( .B1(n5685), .B2(n6510), .A(n5684), .ZN(n5686) );
  AOI21_X1 U6832 ( .B1(n5687), .B2(n5795), .A(n5686), .ZN(n5688) );
  OAI21_X1 U6833 ( .B1(n5689), .B2(n6298), .A(n5688), .ZN(U2957) );
  XNOR2_X1 U6834 ( .A(n5808), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5691)
         );
  NAND2_X1 U6835 ( .A1(n5826), .A2(n6505), .ZN(n5695) );
  NOR2_X1 U6836 ( .A1(n6524), .A2(n6799), .ZN(n5830) );
  NOR2_X1 U6837 ( .A1(n5762), .A2(n3022), .ZN(n5692) );
  AOI211_X1 U6838 ( .C1(n5764), .C2(n5693), .A(n5830), .B(n5692), .ZN(n5694)
         );
  OAI211_X1 U6839 ( .C1(n5816), .C2(n5696), .A(n5695), .B(n5694), .ZN(U2960)
         );
  OAI21_X1 U6840 ( .B1(n4295), .B2(n5698), .A(n5697), .ZN(n5834) );
  NAND2_X1 U6841 ( .A1(n5834), .A2(n6505), .ZN(n5703) );
  INV_X1 U6842 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5699) );
  NOR2_X1 U6843 ( .A1(n6524), .A2(n5699), .ZN(n5837) );
  NOR2_X1 U6844 ( .A1(n6510), .A2(n5700), .ZN(n5701) );
  AOI211_X1 U6845 ( .C1(n6501), .C2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n5837), 
        .B(n5701), .ZN(n5702) );
  OAI211_X1 U6846 ( .C1(n5816), .C2(n5704), .A(n5703), .B(n5702), .ZN(U2961)
         );
  AOI21_X1 U6847 ( .B1(n5705), .B2(n5706), .A(n2958), .ZN(n5860) );
  NOR2_X1 U6848 ( .A1(n6524), .A2(n6670), .ZN(n5853) );
  AOI21_X1 U6849 ( .B1(n6501), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5853), 
        .ZN(n5707) );
  OAI21_X1 U6850 ( .B1(n5708), .B2(n6510), .A(n5707), .ZN(n5709) );
  AOI21_X1 U6851 ( .B1(n5710), .B2(n5795), .A(n5709), .ZN(n5711) );
  OAI21_X1 U6852 ( .B1(n5860), .B2(n6298), .A(n5711), .ZN(U2965) );
  XNOR2_X1 U6853 ( .A(n4306), .B(n5712), .ZN(n5869) );
  XOR2_X1 U6854 ( .A(n5714), .B(n5713), .Z(n5718) );
  INV_X1 U6855 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6668) );
  NOR2_X1 U6856 ( .A1(n6524), .A2(n6668), .ZN(n5865) );
  AOI21_X1 U6857 ( .B1(n6501), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5865), 
        .ZN(n5715) );
  OAI21_X1 U6858 ( .B1(n5716), .B2(n6510), .A(n5715), .ZN(n5717) );
  AOI21_X1 U6859 ( .B1(n5718), .B2(n5795), .A(n5717), .ZN(n5719) );
  OAI21_X1 U6860 ( .B1(n6298), .B2(n5869), .A(n5719), .ZN(U2966) );
  BUF_X1 U6861 ( .A(n5720), .Z(n5721) );
  OAI21_X1 U6862 ( .B1(n2982), .B2(n3757), .A(n5721), .ZN(n5722) );
  XNOR2_X1 U6863 ( .A(n5722), .B(n5808), .ZN(n5877) );
  NAND2_X1 U6864 ( .A1(n6573), .A2(REIP_REG_19__SCAN_IN), .ZN(n5871) );
  NAND2_X1 U6865 ( .A1(n6501), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5723)
         );
  OAI211_X1 U6866 ( .C1(n6510), .C2(n5724), .A(n5871), .B(n5723), .ZN(n5725)
         );
  AOI21_X1 U6867 ( .B1(n5726), .B2(n5795), .A(n5725), .ZN(n5727) );
  OAI21_X1 U6868 ( .B1(n6298), .B2(n5877), .A(n5727), .ZN(U2967) );
  INV_X1 U6869 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5906) );
  XNOR2_X1 U6870 ( .A(n5808), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5768)
         );
  NAND2_X1 U6871 ( .A1(n5808), .A2(n5899), .ZN(n5755) );
  NAND2_X1 U6872 ( .A1(n5758), .A2(n5755), .ZN(n5743) );
  NAND2_X1 U6873 ( .A1(n5808), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5744) );
  XNOR2_X1 U6874 ( .A(n5731), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5884)
         );
  INV_X1 U6875 ( .A(n5732), .ZN(n5737) );
  NOR2_X1 U6876 ( .A1(n6524), .A2(n5733), .ZN(n5878) );
  AOI21_X1 U6877 ( .B1(n6501), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5878), 
        .ZN(n5734) );
  OAI21_X1 U6878 ( .B1(n5735), .B2(n6510), .A(n5734), .ZN(n5736) );
  AOI21_X1 U6879 ( .B1(n5737), .B2(n5795), .A(n5736), .ZN(n5738) );
  OAI21_X1 U6880 ( .B1(n5884), .B2(n6298), .A(n5738), .ZN(U2968) );
  NAND2_X1 U6881 ( .A1(n4296), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U6882 ( .A1(n5743), .A2(n5756), .ZN(n5742) );
  NOR2_X1 U6883 ( .A1(n5808), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5740)
         );
  INV_X1 U6884 ( .A(n5744), .ZN(n5739) );
  INV_X1 U6885 ( .A(n5743), .ZN(n5745) );
  NAND3_X1 U6886 ( .A1(n5748), .A2(n5747), .A3(n5746), .ZN(n5885) );
  NAND2_X1 U6887 ( .A1(n5885), .A2(n6505), .ZN(n5753) );
  NAND2_X1 U6888 ( .A1(n6573), .A2(REIP_REG_17__SCAN_IN), .ZN(n5892) );
  OAI21_X1 U6889 ( .B1(n5762), .B2(n5749), .A(n5892), .ZN(n5750) );
  AOI21_X1 U6890 ( .B1(n5764), .B2(n5751), .A(n5750), .ZN(n5752) );
  OAI211_X1 U6891 ( .C1(n5816), .C2(n5754), .A(n5753), .B(n5752), .ZN(U2969)
         );
  NAND2_X1 U6892 ( .A1(n5756), .A2(n5755), .ZN(n5757) );
  XNOR2_X1 U6893 ( .A(n5758), .B(n5757), .ZN(n5895) );
  NAND2_X1 U6894 ( .A1(n5895), .A2(n6505), .ZN(n5766) );
  NOR2_X1 U6895 ( .A1(n6524), .A2(n5759), .ZN(n5901) );
  INV_X1 U6896 ( .A(n5901), .ZN(n5760) );
  OAI21_X1 U6897 ( .B1(n5762), .B2(n5761), .A(n5760), .ZN(n5763) );
  AOI21_X1 U6898 ( .B1(n5764), .B2(n6322), .A(n5763), .ZN(n5765) );
  OAI211_X1 U6899 ( .C1(n5816), .C2(n6321), .A(n5766), .B(n5765), .ZN(U2970)
         );
  INV_X1 U6900 ( .A(n5767), .ZN(n5771) );
  INV_X1 U6901 ( .A(n5768), .ZN(n5770) );
  AOI21_X1 U6902 ( .B1(n5771), .B2(n5770), .A(n5769), .ZN(n5913) );
  NAND2_X1 U6903 ( .A1(n6573), .A2(REIP_REG_15__SCAN_IN), .ZN(n5905) );
  NAND2_X1 U6904 ( .A1(n6501), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5772)
         );
  OAI211_X1 U6905 ( .C1(n6510), .C2(n5773), .A(n5905), .B(n5772), .ZN(n5774)
         );
  AOI21_X1 U6906 ( .B1(n5775), .B2(n5795), .A(n5774), .ZN(n5776) );
  OAI21_X1 U6907 ( .B1(n5913), .B2(n6298), .A(n5776), .ZN(U2971) );
  OAI21_X1 U6908 ( .B1(n5779), .B2(n5778), .A(n5777), .ZN(n5780) );
  INV_X1 U6909 ( .A(n5780), .ZN(n5936) );
  NAND2_X1 U6910 ( .A1(n6573), .A2(REIP_REG_13__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U6911 ( .A1(n6501), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5781)
         );
  OAI211_X1 U6912 ( .C1(n6510), .C2(n6329), .A(n5931), .B(n5781), .ZN(n5782)
         );
  AOI21_X1 U6913 ( .B1(n6331), .B2(n5795), .A(n5782), .ZN(n5783) );
  OAI21_X1 U6914 ( .B1(n5936), .B2(n6298), .A(n5783), .ZN(U2973) );
  XOR2_X1 U6915 ( .A(n5785), .B(n5784), .Z(n5946) );
  NOR2_X1 U6916 ( .A1(n6524), .A2(n6663), .ZN(n5944) );
  AOI21_X1 U6917 ( .B1(n6501), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n5944), 
        .ZN(n5786) );
  OAI21_X1 U6918 ( .B1(n6349), .B2(n6510), .A(n5786), .ZN(n5787) );
  AOI21_X1 U6919 ( .B1(n6418), .B2(n5795), .A(n5787), .ZN(n5788) );
  OAI21_X1 U6920 ( .B1(n5946), .B2(n6298), .A(n5788), .ZN(U2974) );
  NAND2_X1 U6921 ( .A1(n5789), .A2(n5799), .ZN(n5791) );
  XNOR2_X1 U6922 ( .A(n5808), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5790)
         );
  XNOR2_X1 U6923 ( .A(n5791), .B(n5790), .ZN(n5954) );
  NAND2_X1 U6924 ( .A1(n6573), .A2(REIP_REG_11__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U6925 ( .A1(n6501), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5792)
         );
  OAI211_X1 U6926 ( .C1(n6510), .C2(n5793), .A(n5948), .B(n5792), .ZN(n5794)
         );
  AOI21_X1 U6927 ( .B1(n5796), .B2(n5795), .A(n5794), .ZN(n5797) );
  OAI21_X1 U6928 ( .B1(n5954), .B2(n6298), .A(n5797), .ZN(U2975) );
  NAND2_X1 U6929 ( .A1(n5799), .A2(n5798), .ZN(n5801) );
  XOR2_X1 U6930 ( .A(n5801), .B(n5800), .Z(n5971) );
  INV_X1 U6931 ( .A(n6354), .ZN(n5804) );
  AOI22_X1 U6932 ( .A1(n6501), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6573), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5802) );
  OAI21_X1 U6933 ( .B1(n6353), .B2(n6510), .A(n5802), .ZN(n5803) );
  AOI21_X1 U6934 ( .B1(n5804), .B2(n5795), .A(n5803), .ZN(n5805) );
  OAI21_X1 U6935 ( .B1(n5971), .B2(n6298), .A(n5805), .ZN(U2976) );
  XNOR2_X1 U6936 ( .A(n5808), .B(n5807), .ZN(n5809) );
  XNOR2_X1 U6937 ( .A(n5806), .B(n5809), .ZN(n6515) );
  NAND2_X1 U6938 ( .A1(n6515), .A2(n6505), .ZN(n5814) );
  INV_X1 U6939 ( .A(REIP_REG_9__SCAN_IN), .ZN(n5810) );
  NOR2_X1 U6940 ( .A1(n6524), .A2(n5810), .ZN(n6512) );
  NOR2_X1 U6941 ( .A1(n6510), .A2(n5811), .ZN(n5812) );
  AOI211_X1 U6942 ( .C1(n6501), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6512), 
        .B(n5812), .ZN(n5813) );
  OAI211_X1 U6943 ( .C1(n5816), .C2(n5815), .A(n5814), .B(n5813), .ZN(U2977)
         );
  OAI21_X1 U6944 ( .B1(n5818), .B2(n5822), .A(n5817), .ZN(n5821) );
  NOR2_X1 U6945 ( .A1(n5819), .A2(n5966), .ZN(n5820) );
  AOI211_X1 U6946 ( .C1(n5823), .C2(n5822), .A(n5821), .B(n5820), .ZN(n5824)
         );
  OAI21_X1 U6947 ( .B1(n5825), .B2(n6520), .A(n5824), .ZN(U2991) );
  NAND2_X1 U6948 ( .A1(n5826), .A2(n6579), .ZN(n5832) );
  NOR3_X1 U6949 ( .A1(n5835), .A2(n5828), .A3(n5827), .ZN(n5829) );
  AOI211_X1 U6950 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n5838), .A(n5830), .B(n5829), .ZN(n5831) );
  OAI211_X1 U6951 ( .C1(n5966), .C2(n5833), .A(n5832), .B(n5831), .ZN(U2992)
         );
  NAND2_X1 U6952 ( .A1(n5834), .A2(n6579), .ZN(n5840) );
  NOR2_X1 U6953 ( .A1(n5835), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5836)
         );
  AOI211_X1 U6954 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5838), .A(n5837), .B(n5836), .ZN(n5839) );
  OAI211_X1 U6955 ( .C1(n5966), .C2(n5841), .A(n5840), .B(n5839), .ZN(U2993)
         );
  INV_X1 U6956 ( .A(n5842), .ZN(n5852) );
  INV_X1 U6957 ( .A(n5843), .ZN(n5849) );
  INV_X1 U6958 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5847) );
  AOI211_X1 U6959 ( .C1(n5847), .C2(n5846), .A(n5845), .B(n5844), .ZN(n5848)
         );
  AOI211_X1 U6960 ( .C1(n5850), .C2(n6541), .A(n5849), .B(n5848), .ZN(n5851)
         );
  OAI21_X1 U6961 ( .B1(n5852), .B2(n6520), .A(n5851), .ZN(U2994) );
  AOI21_X1 U6962 ( .B1(n5854), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5853), 
        .ZN(n5855) );
  OAI21_X1 U6963 ( .B1(n5856), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5855), 
        .ZN(n5857) );
  AOI21_X1 U6964 ( .B1(n5858), .B2(n6541), .A(n5857), .ZN(n5859) );
  OAI21_X1 U6965 ( .B1(n5860), .B2(n6520), .A(n5859), .ZN(U2997) );
  INV_X1 U6966 ( .A(n5861), .ZN(n5939) );
  AOI22_X1 U6967 ( .A1(n5896), .A2(n5888), .B1(n5938), .B2(n5889), .ZN(n5862)
         );
  NAND2_X1 U6968 ( .A1(n5862), .A2(n5942), .ZN(n5886) );
  AOI21_X1 U6969 ( .B1(n5939), .B2(n5889), .A(n5886), .ZN(n5880) );
  OAI21_X1 U6970 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5964), .A(n5880), 
        .ZN(n5870) );
  AOI211_X1 U6971 ( .C1(n3757), .C2(n6838), .A(n5863), .B(n5873), .ZN(n5864)
         );
  AOI211_X1 U6972 ( .C1(INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n5870), .A(n5865), .B(n5864), .ZN(n5868) );
  NAND2_X1 U6973 ( .A1(n5866), .A2(n6541), .ZN(n5867) );
  OAI211_X1 U6974 ( .C1(n5869), .C2(n6520), .A(n5868), .B(n5867), .ZN(U2998)
         );
  NAND2_X1 U6975 ( .A1(n5870), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5872) );
  OAI211_X1 U6976 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n5873), .A(n5872), .B(n5871), .ZN(n5874) );
  AOI21_X1 U6977 ( .B1(n6541), .B2(n5875), .A(n5874), .ZN(n5876) );
  OAI21_X1 U6978 ( .B1(n5877), .B2(n6520), .A(n5876), .ZN(U2999) );
  AOI21_X1 U6979 ( .B1(n5879), .B2(n4314), .A(n5878), .ZN(n5883) );
  MUX2_X1 U6980 ( .A(n5881), .B(n5880), .S(INSTADDRPOINTER_REG_18__SCAN_IN), 
        .Z(n5882) );
  OAI211_X1 U6981 ( .C1(n5884), .C2(n6520), .A(n5883), .B(n5882), .ZN(U3000)
         );
  NAND2_X1 U6982 ( .A1(n5885), .A2(n6579), .ZN(n5894) );
  AOI22_X1 U6983 ( .A1(n5887), .A2(n6541), .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5886), .ZN(n5893) );
  INV_X1 U6984 ( .A(n5888), .ZN(n5890) );
  NAND3_X1 U6985 ( .A1(n5952), .A2(n5890), .A3(n5889), .ZN(n5891) );
  NAND4_X1 U6986 ( .A1(n5894), .A2(n5893), .A3(n5892), .A4(n5891), .ZN(U3001)
         );
  NAND2_X1 U6987 ( .A1(n5895), .A2(n6579), .ZN(n5904) );
  NOR3_X1 U6988 ( .A1(n5897), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5906), 
        .ZN(n5902) );
  INV_X1 U6989 ( .A(n5942), .ZN(n5947) );
  AOI21_X1 U6990 ( .B1(n5897), .B2(n5896), .A(n5947), .ZN(n5907) );
  INV_X1 U6991 ( .A(n5897), .ZN(n5898) );
  NAND3_X1 U6992 ( .A1(n5952), .A2(n5898), .A3(n5906), .ZN(n5911) );
  AOI21_X1 U6993 ( .B1(n5907), .B2(n5911), .A(n5899), .ZN(n5900) );
  AOI211_X1 U6994 ( .C1(n5902), .C2(n5952), .A(n5901), .B(n5900), .ZN(n5903)
         );
  OAI211_X1 U6995 ( .C1(n6325), .C2(n5966), .A(n5904), .B(n5903), .ZN(U3002)
         );
  INV_X1 U6996 ( .A(n5905), .ZN(n5909) );
  NOR2_X1 U6997 ( .A1(n5907), .A2(n5906), .ZN(n5908) );
  AOI211_X1 U6998 ( .C1(n6541), .C2(n5910), .A(n5909), .B(n5908), .ZN(n5912)
         );
  OAI211_X1 U6999 ( .C1(n5913), .C2(n6520), .A(n5912), .B(n5911), .ZN(U3003)
         );
  NAND3_X1 U7000 ( .A1(n5952), .A2(n5922), .A3(n5914), .ZN(n5915) );
  OAI211_X1 U7001 ( .C1(n5917), .C2(n5966), .A(n5916), .B(n5915), .ZN(n5918)
         );
  INV_X1 U7002 ( .A(n5918), .ZN(n5927) );
  NAND2_X1 U7003 ( .A1(n5919), .A2(n5937), .ZN(n5920) );
  OAI211_X1 U7004 ( .C1(n5922), .C2(n5921), .A(n5942), .B(n5920), .ZN(n5934)
         );
  AOI21_X1 U7005 ( .B1(n5924), .B2(n5923), .A(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5925) );
  OAI21_X1 U7006 ( .B1(n5934), .B2(n5925), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5926) );
  OAI211_X1 U7007 ( .C1(n5928), .C2(n6520), .A(n5927), .B(n5926), .ZN(U3004)
         );
  INV_X1 U7008 ( .A(n5937), .ZN(n5930) );
  NAND3_X1 U7009 ( .A1(n5952), .A2(n5930), .A3(n5929), .ZN(n5932) );
  OAI211_X1 U7010 ( .C1(n6326), .C2(n5966), .A(n5932), .B(n5931), .ZN(n5933)
         );
  AOI21_X1 U7011 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5934), .A(n5933), 
        .ZN(n5935) );
  OAI21_X1 U7012 ( .B1(n5936), .B2(n6520), .A(n5935), .ZN(U3005) );
  OAI21_X1 U7013 ( .B1(n5939), .B2(n5938), .A(n5937), .ZN(n5941) );
  AOI21_X1 U7014 ( .B1(n5952), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5940) );
  AOI21_X1 U7015 ( .B1(n5942), .B2(n5941), .A(n5940), .ZN(n5943) );
  AOI211_X1 U7016 ( .C1(n6541), .C2(n6343), .A(n5944), .B(n5943), .ZN(n5945)
         );
  OAI21_X1 U7017 ( .B1(n5946), .B2(n6520), .A(n5945), .ZN(U3006) );
  NAND2_X1 U7018 ( .A1(n5947), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5949) );
  OAI211_X1 U7019 ( .C1(n5966), .C2(n5950), .A(n5949), .B(n5948), .ZN(n5951)
         );
  AOI21_X1 U7020 ( .B1(n6802), .B2(n5952), .A(n5951), .ZN(n5953) );
  OAI21_X1 U7021 ( .B1(n5954), .B2(n6520), .A(n5953), .ZN(U3007) );
  NAND2_X1 U7022 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n5955), .ZN(n6537)
         );
  NOR2_X1 U7023 ( .A1(n5957), .A2(n6537), .ZN(n6514) );
  OAI211_X1 U7024 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6514), .B(n5956), .ZN(n5970) );
  INV_X1 U7025 ( .A(n5957), .ZN(n6519) );
  INV_X1 U7026 ( .A(n5958), .ZN(n5960) );
  OAI22_X1 U7027 ( .A1(n5961), .A2(n6577), .B1(n5960), .B2(n5959), .ZN(n5962)
         );
  NOR2_X1 U7028 ( .A1(n5963), .A2(n5962), .ZN(n6535) );
  OAI21_X1 U7029 ( .B1(n6519), .B2(n5964), .A(n6535), .ZN(n6511) );
  OAI22_X1 U7030 ( .A1(n5967), .A2(n5966), .B1(n5965), .B2(n6524), .ZN(n5968)
         );
  AOI21_X1 U7031 ( .B1(n6511), .B2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n5968), 
        .ZN(n5969) );
  OAI211_X1 U7032 ( .C1(n5971), .C2(n6520), .A(n5970), .B(n5969), .ZN(U3008)
         );
  OAI211_X1 U7033 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n5972), .A(n5976), .B(
        n6203), .ZN(n5973) );
  OAI21_X1 U7034 ( .B1(n5977), .B2(n4435), .A(n5973), .ZN(n5974) );
  MUX2_X1 U7035 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5974), .S(n6584), 
        .Z(U3464) );
  XNOR2_X1 U7036 ( .A(n5976), .B(n5975), .ZN(n5978) );
  OAI22_X1 U7037 ( .A1(n5978), .A2(n6691), .B1(n4534), .B2(n5977), .ZN(n5979)
         );
  MUX2_X1 U7038 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5979), .S(n6584), 
        .Z(U3463) );
  INV_X1 U7039 ( .A(n5980), .ZN(n5982) );
  OAI22_X1 U7040 ( .A1(n5982), .A2(n6646), .B1(n5981), .B2(n6283), .ZN(n5983)
         );
  MUX2_X1 U7041 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5983), .S(n6294), 
        .Z(U3456) );
  OAI21_X1 U7042 ( .B1(n5987), .B2(n6691), .A(n6149), .ZN(n5991) );
  INV_X1 U7043 ( .A(n6016), .ZN(n5984) );
  OAI21_X1 U7044 ( .B1(n5985), .B2(n3583), .A(n5984), .ZN(n5988) );
  INV_X1 U7045 ( .A(n5988), .ZN(n5992) );
  INV_X1 U7046 ( .A(n5989), .ZN(n5990) );
  AOI22_X1 U7047 ( .A1(n5992), .A2(n5991), .B1(n6691), .B2(n5990), .ZN(n5993)
         );
  NAND2_X1 U7048 ( .A1(n6161), .A2(n5993), .ZN(n6015) );
  AOI22_X1 U7049 ( .A1(n6162), .A2(n6016), .B1(INSTQUEUE_REG_1__0__SCAN_IN), 
        .B2(n6015), .ZN(n5994) );
  OAI21_X1 U7050 ( .B1(n6058), .B2(n6597), .A(n5994), .ZN(n5995) );
  AOI21_X1 U7051 ( .B1(n6222), .B2(n6019), .A(n5995), .ZN(n5996) );
  OAI21_X1 U7052 ( .B1(n6021), .B2(n6220), .A(n5996), .ZN(U3028) );
  AOI22_X1 U7053 ( .A1(n6226), .A2(n6016), .B1(INSTQUEUE_REG_1__1__SCAN_IN), 
        .B2(n6015), .ZN(n5997) );
  OAI21_X1 U7054 ( .B1(n6058), .B2(n6233), .A(n5997), .ZN(n5998) );
  AOI21_X1 U7055 ( .B1(n6230), .B2(n6019), .A(n5998), .ZN(n5999) );
  OAI21_X1 U7056 ( .B1(n6021), .B2(n6228), .A(n5999), .ZN(U3029) );
  AOI22_X1 U7057 ( .A1(n6234), .A2(n6016), .B1(INSTQUEUE_REG_1__2__SCAN_IN), 
        .B2(n6015), .ZN(n6000) );
  OAI21_X1 U7058 ( .B1(n6058), .B2(n6241), .A(n6000), .ZN(n6001) );
  AOI21_X1 U7059 ( .B1(n6238), .B2(n6019), .A(n6001), .ZN(n6002) );
  OAI21_X1 U7060 ( .B1(n6021), .B2(n6236), .A(n6002), .ZN(U3030) );
  AOI22_X1 U7061 ( .A1(n6242), .A2(n6016), .B1(INSTQUEUE_REG_1__3__SCAN_IN), 
        .B2(n6015), .ZN(n6003) );
  OAI21_X1 U7062 ( .B1(n6058), .B2(n6604), .A(n6003), .ZN(n6004) );
  AOI21_X1 U7063 ( .B1(n6246), .B2(n6019), .A(n6004), .ZN(n6005) );
  OAI21_X1 U7064 ( .B1(n6021), .B2(n6244), .A(n6005), .ZN(U3031) );
  AOI22_X1 U7065 ( .A1(n6249), .A2(n6016), .B1(INSTQUEUE_REG_1__4__SCAN_IN), 
        .B2(n6015), .ZN(n6006) );
  OAI21_X1 U7066 ( .B1(n6058), .B2(n6611), .A(n6006), .ZN(n6007) );
  AOI21_X1 U7067 ( .B1(n6253), .B2(n6019), .A(n6007), .ZN(n6008) );
  OAI21_X1 U7068 ( .B1(n6021), .B2(n6251), .A(n6008), .ZN(U3032) );
  AOI22_X1 U7069 ( .A1(n6256), .A2(n6016), .B1(INSTQUEUE_REG_1__5__SCAN_IN), 
        .B2(n6015), .ZN(n6009) );
  OAI21_X1 U7070 ( .B1(n6058), .B2(n6618), .A(n6009), .ZN(n6010) );
  AOI21_X1 U7071 ( .B1(n6260), .B2(n6019), .A(n6010), .ZN(n6011) );
  OAI21_X1 U7072 ( .B1(n6021), .B2(n6258), .A(n6011), .ZN(U3033) );
  AOI22_X1 U7073 ( .A1(n6263), .A2(n6016), .B1(INSTQUEUE_REG_1__6__SCAN_IN), 
        .B2(n6015), .ZN(n6012) );
  OAI21_X1 U7074 ( .B1(n6058), .B2(n6625), .A(n6012), .ZN(n6013) );
  AOI21_X1 U7075 ( .B1(n6267), .B2(n6019), .A(n6013), .ZN(n6014) );
  OAI21_X1 U7076 ( .B1(n6021), .B2(n6265), .A(n6014), .ZN(U3034) );
  AOI22_X1 U7077 ( .A1(n6272), .A2(n6016), .B1(INSTQUEUE_REG_1__7__SCAN_IN), 
        .B2(n6015), .ZN(n6017) );
  OAI21_X1 U7078 ( .B1(n6058), .B2(n6633), .A(n6017), .ZN(n6018) );
  AOI21_X1 U7079 ( .B1(n6277), .B2(n6019), .A(n6018), .ZN(n6020) );
  OAI21_X1 U7080 ( .B1(n6021), .B2(n6274), .A(n6020), .ZN(U3035) );
  INV_X1 U7081 ( .A(n6028), .ZN(n6024) );
  NOR2_X1 U7082 ( .A1(n6022), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6066)
         );
  AOI22_X1 U7083 ( .A1(n6024), .A2(n6203), .B1(n6023), .B2(n6066), .ZN(n6054)
         );
  INV_X1 U7084 ( .A(n6058), .ZN(n6026) );
  OAI21_X1 U7085 ( .B1(n6056), .B2(n6026), .A(n6149), .ZN(n6027) );
  NAND2_X1 U7086 ( .A1(n6028), .A2(n6027), .ZN(n6030) );
  OAI221_X1 U7087 ( .B1(n3098), .B2(n6103), .C1(n3098), .C2(n6030), .A(n6029), 
        .ZN(n6052) );
  AOI22_X1 U7088 ( .A1(n6162), .A2(n3098), .B1(INSTQUEUE_REG_2__0__SCAN_IN), 
        .B2(n6052), .ZN(n6031) );
  OAI21_X1 U7089 ( .B1(n6054), .B2(n6220), .A(n6031), .ZN(n6032) );
  AOI21_X1 U7090 ( .B1(n6056), .B2(n6165), .A(n6032), .ZN(n6033) );
  OAI21_X1 U7091 ( .B1(n6602), .B2(n6058), .A(n6033), .ZN(U3036) );
  AOI22_X1 U7092 ( .A1(n6226), .A2(n3098), .B1(INSTQUEUE_REG_2__1__SCAN_IN), 
        .B2(n6052), .ZN(n6034) );
  OAI21_X1 U7093 ( .B1(n6054), .B2(n6228), .A(n6034), .ZN(n6035) );
  AOI21_X1 U7094 ( .B1(n6056), .B2(n6170), .A(n6035), .ZN(n6036) );
  OAI21_X1 U7095 ( .B1(n6168), .B2(n6058), .A(n6036), .ZN(U3037) );
  AOI22_X1 U7096 ( .A1(n6234), .A2(n3098), .B1(INSTQUEUE_REG_2__2__SCAN_IN), 
        .B2(n6052), .ZN(n6037) );
  OAI21_X1 U7097 ( .B1(n6054), .B2(n6236), .A(n6037), .ZN(n6038) );
  AOI21_X1 U7098 ( .B1(n6056), .B2(n6175), .A(n6038), .ZN(n6039) );
  OAI21_X1 U7099 ( .B1(n6173), .B2(n6058), .A(n6039), .ZN(U3038) );
  AOI22_X1 U7100 ( .A1(n6242), .A2(n3098), .B1(INSTQUEUE_REG_2__3__SCAN_IN), 
        .B2(n6052), .ZN(n6040) );
  OAI21_X1 U7101 ( .B1(n6054), .B2(n6244), .A(n6040), .ZN(n6041) );
  AOI21_X1 U7102 ( .B1(n6056), .B2(n6179), .A(n6041), .ZN(n6042) );
  OAI21_X1 U7103 ( .B1(n6609), .B2(n6058), .A(n6042), .ZN(U3039) );
  AOI22_X1 U7104 ( .A1(n6249), .A2(n3098), .B1(INSTQUEUE_REG_2__4__SCAN_IN), 
        .B2(n6052), .ZN(n6043) );
  OAI21_X1 U7105 ( .B1(n6054), .B2(n6251), .A(n6043), .ZN(n6044) );
  AOI21_X1 U7106 ( .B1(n6056), .B2(n6183), .A(n6044), .ZN(n6045) );
  OAI21_X1 U7107 ( .B1(n6616), .B2(n6058), .A(n6045), .ZN(U3040) );
  AOI22_X1 U7108 ( .A1(n6256), .A2(n3098), .B1(INSTQUEUE_REG_2__5__SCAN_IN), 
        .B2(n6052), .ZN(n6046) );
  OAI21_X1 U7109 ( .B1(n6054), .B2(n6258), .A(n6046), .ZN(n6047) );
  AOI21_X1 U7110 ( .B1(n6056), .B2(n6187), .A(n6047), .ZN(n6048) );
  OAI21_X1 U7111 ( .B1(n6623), .B2(n6058), .A(n6048), .ZN(U3041) );
  AOI22_X1 U7112 ( .A1(n6263), .A2(n3098), .B1(INSTQUEUE_REG_2__6__SCAN_IN), 
        .B2(n6052), .ZN(n6049) );
  OAI21_X1 U7113 ( .B1(n6054), .B2(n6265), .A(n6049), .ZN(n6050) );
  AOI21_X1 U7114 ( .B1(n6056), .B2(n6191), .A(n6050), .ZN(n6051) );
  OAI21_X1 U7115 ( .B1(n6630), .B2(n6058), .A(n6051), .ZN(U3042) );
  AOI22_X1 U7116 ( .A1(n6272), .A2(n3098), .B1(INSTQUEUE_REG_2__7__SCAN_IN), 
        .B2(n6052), .ZN(n6053) );
  OAI21_X1 U7117 ( .B1(n6054), .B2(n6274), .A(n6053), .ZN(n6055) );
  AOI21_X1 U7118 ( .B1(n6056), .B2(n6198), .A(n6055), .ZN(n6057) );
  OAI21_X1 U7119 ( .B1(n6642), .B2(n6058), .A(n6057), .ZN(U3043) );
  OAI21_X1 U7120 ( .B1(n6059), .B2(n6095), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6061) );
  NAND3_X1 U7121 ( .A1(n6061), .A2(n6203), .A3(n6060), .ZN(n6064) );
  NAND2_X1 U7122 ( .A1(n6062), .A2(n6207), .ZN(n6092) );
  AOI21_X1 U7123 ( .B1(n6092), .B2(STATE2_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U7124 ( .A1(n6091), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n6070) );
  INV_X1 U7125 ( .A(n6065), .ZN(n6205) );
  NOR2_X1 U7126 ( .A1(n6205), .A2(n6691), .ZN(n6219) );
  AOI22_X1 U7127 ( .A1(n6219), .A2(n6206), .B1(n6067), .B2(n6066), .ZN(n6093)
         );
  OAI22_X1 U7128 ( .A1(n6093), .A2(n6220), .B1(n6596), .B2(n6092), .ZN(n6068)
         );
  AOI21_X1 U7129 ( .B1(n6095), .B2(n6222), .A(n6068), .ZN(n6069) );
  OAI211_X1 U7130 ( .C1(n6098), .C2(n6597), .A(n6070), .B(n6069), .ZN(U3068)
         );
  NAND2_X1 U7131 ( .A1(n6091), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n6074) );
  OAI22_X1 U7132 ( .A1(n6093), .A2(n6228), .B1(n6071), .B2(n6092), .ZN(n6072)
         );
  AOI21_X1 U7133 ( .B1(n6095), .B2(n6230), .A(n6072), .ZN(n6073) );
  OAI211_X1 U7134 ( .C1(n6098), .C2(n6233), .A(n6074), .B(n6073), .ZN(U3069)
         );
  NAND2_X1 U7135 ( .A1(n6091), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n6078) );
  OAI22_X1 U7136 ( .A1(n6093), .A2(n6236), .B1(n6075), .B2(n6092), .ZN(n6076)
         );
  AOI21_X1 U7137 ( .B1(n6095), .B2(n6238), .A(n6076), .ZN(n6077) );
  OAI211_X1 U7138 ( .C1(n6098), .C2(n6241), .A(n6078), .B(n6077), .ZN(U3070)
         );
  NAND2_X1 U7139 ( .A1(n6091), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n6081) );
  OAI22_X1 U7140 ( .A1(n6093), .A2(n6244), .B1(n6603), .B2(n6092), .ZN(n6079)
         );
  AOI21_X1 U7141 ( .B1(n6095), .B2(n6246), .A(n6079), .ZN(n6080) );
  OAI211_X1 U7142 ( .C1(n6098), .C2(n6604), .A(n6081), .B(n6080), .ZN(U3071)
         );
  NAND2_X1 U7143 ( .A1(n6091), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n6084) );
  OAI22_X1 U7144 ( .A1(n6093), .A2(n6251), .B1(n6610), .B2(n6092), .ZN(n6082)
         );
  AOI21_X1 U7145 ( .B1(n6095), .B2(n6253), .A(n6082), .ZN(n6083) );
  OAI211_X1 U7146 ( .C1(n6098), .C2(n6611), .A(n6084), .B(n6083), .ZN(U3072)
         );
  NAND2_X1 U7147 ( .A1(n6091), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n6087) );
  OAI22_X1 U7148 ( .A1(n6093), .A2(n6258), .B1(n6617), .B2(n6092), .ZN(n6085)
         );
  AOI21_X1 U7149 ( .B1(n6095), .B2(n6260), .A(n6085), .ZN(n6086) );
  OAI211_X1 U7150 ( .C1(n6098), .C2(n6618), .A(n6087), .B(n6086), .ZN(U3073)
         );
  NAND2_X1 U7151 ( .A1(n6091), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n6090) );
  OAI22_X1 U7152 ( .A1(n6093), .A2(n6265), .B1(n6624), .B2(n6092), .ZN(n6088)
         );
  AOI21_X1 U7153 ( .B1(n6095), .B2(n6267), .A(n6088), .ZN(n6089) );
  OAI211_X1 U7154 ( .C1(n6098), .C2(n6625), .A(n6090), .B(n6089), .ZN(U3074)
         );
  NAND2_X1 U7155 ( .A1(n6091), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n6097) );
  OAI22_X1 U7156 ( .A1(n6093), .A2(n6274), .B1(n6632), .B2(n6092), .ZN(n6094)
         );
  AOI21_X1 U7157 ( .B1(n6095), .B2(n6277), .A(n6094), .ZN(n6096) );
  OAI211_X1 U7158 ( .C1(n6098), .C2(n6633), .A(n6097), .B(n6096), .ZN(U3075)
         );
  NAND3_X1 U7159 ( .A1(n6196), .A2(n6203), .A3(n6143), .ZN(n6100) );
  NOR2_X1 U7160 ( .A1(n6206), .A2(n6151), .ZN(n6107) );
  AOI21_X1 U7161 ( .B1(n6100), .B2(n6149), .A(n6107), .ZN(n6106) );
  AND2_X1 U7162 ( .A1(n6102), .A2(n6101), .ZN(n6156) );
  AND2_X1 U7163 ( .A1(n6156), .A2(n6207), .ZN(n6140) );
  OAI21_X1 U7164 ( .B1(n6140), .B2(n6103), .A(n6216), .ZN(n6104) );
  NOR3_X2 U7165 ( .A1(n6106), .A2(n6105), .A3(n6104), .ZN(n6148) );
  INV_X1 U7166 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n6113) );
  INV_X1 U7167 ( .A(n6107), .ZN(n6109) );
  OAI22_X1 U7168 ( .A1(n6109), .A2(n6691), .B1(n6211), .B2(n6108), .ZN(n6141)
         );
  AOI22_X1 U7169 ( .A1(n6141), .A2(n6599), .B1(n6162), .B2(n6140), .ZN(n6110)
         );
  OAI21_X1 U7170 ( .B1(n6143), .B2(n6602), .A(n6110), .ZN(n6111) );
  AOI21_X1 U7171 ( .B1(n6145), .B2(n6165), .A(n6111), .ZN(n6112) );
  OAI21_X1 U7172 ( .B1(n6148), .B2(n6113), .A(n6112), .ZN(U3084) );
  INV_X1 U7173 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n6118) );
  AOI22_X1 U7174 ( .A1(n6141), .A2(n6114), .B1(n6226), .B2(n6140), .ZN(n6115)
         );
  OAI21_X1 U7175 ( .B1(n6143), .B2(n6168), .A(n6115), .ZN(n6116) );
  AOI21_X1 U7176 ( .B1(n6145), .B2(n6170), .A(n6116), .ZN(n6117) );
  OAI21_X1 U7177 ( .B1(n6148), .B2(n6118), .A(n6117), .ZN(U3085) );
  INV_X1 U7178 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n6123) );
  AOI22_X1 U7179 ( .A1(n6141), .A2(n6119), .B1(n6234), .B2(n6140), .ZN(n6120)
         );
  OAI21_X1 U7180 ( .B1(n6143), .B2(n6173), .A(n6120), .ZN(n6121) );
  AOI21_X1 U7181 ( .B1(n6145), .B2(n6175), .A(n6121), .ZN(n6122) );
  OAI21_X1 U7182 ( .B1(n6148), .B2(n6123), .A(n6122), .ZN(U3086) );
  INV_X1 U7183 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n6127) );
  AOI22_X1 U7184 ( .A1(n6141), .A2(n6606), .B1(n6242), .B2(n6140), .ZN(n6124)
         );
  OAI21_X1 U7185 ( .B1(n6143), .B2(n6609), .A(n6124), .ZN(n6125) );
  AOI21_X1 U7186 ( .B1(n6145), .B2(n6179), .A(n6125), .ZN(n6126) );
  OAI21_X1 U7187 ( .B1(n6148), .B2(n6127), .A(n6126), .ZN(U3087) );
  INV_X1 U7188 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n6131) );
  AOI22_X1 U7189 ( .A1(n6141), .A2(n6613), .B1(n6249), .B2(n6140), .ZN(n6128)
         );
  OAI21_X1 U7190 ( .B1(n6143), .B2(n6616), .A(n6128), .ZN(n6129) );
  AOI21_X1 U7191 ( .B1(n6145), .B2(n6183), .A(n6129), .ZN(n6130) );
  OAI21_X1 U7192 ( .B1(n6148), .B2(n6131), .A(n6130), .ZN(U3088) );
  INV_X1 U7193 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n6135) );
  AOI22_X1 U7194 ( .A1(n6141), .A2(n6620), .B1(n6256), .B2(n6140), .ZN(n6132)
         );
  OAI21_X1 U7195 ( .B1(n6143), .B2(n6623), .A(n6132), .ZN(n6133) );
  AOI21_X1 U7196 ( .B1(n6145), .B2(n6187), .A(n6133), .ZN(n6134) );
  OAI21_X1 U7197 ( .B1(n6148), .B2(n6135), .A(n6134), .ZN(U3089) );
  INV_X1 U7198 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n6139) );
  AOI22_X1 U7199 ( .A1(n6141), .A2(n6627), .B1(n6263), .B2(n6140), .ZN(n6136)
         );
  OAI21_X1 U7200 ( .B1(n6143), .B2(n6630), .A(n6136), .ZN(n6137) );
  AOI21_X1 U7201 ( .B1(n6145), .B2(n6191), .A(n6137), .ZN(n6138) );
  OAI21_X1 U7202 ( .B1(n6148), .B2(n6139), .A(n6138), .ZN(U3090) );
  INV_X1 U7203 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n6147) );
  AOI22_X1 U7204 ( .A1(n6141), .A2(n6637), .B1(n6272), .B2(n6140), .ZN(n6142)
         );
  OAI21_X1 U7205 ( .B1(n6143), .B2(n6642), .A(n6142), .ZN(n6144) );
  AOI21_X1 U7206 ( .B1(n6145), .B2(n6198), .A(n6144), .ZN(n6146) );
  OAI21_X1 U7207 ( .B1(n6148), .B2(n6147), .A(n6146), .ZN(U3091) );
  OAI21_X1 U7208 ( .B1(n6150), .B2(n6691), .A(n6149), .ZN(n6158) );
  OR2_X1 U7209 ( .A1(n6152), .A2(n6151), .ZN(n6154) );
  INV_X1 U7210 ( .A(n6194), .ZN(n6153) );
  NAND2_X1 U7211 ( .A1(n6154), .A2(n6153), .ZN(n6155) );
  INV_X1 U7212 ( .A(n6155), .ZN(n6159) );
  INV_X1 U7213 ( .A(n6156), .ZN(n6157) );
  AOI22_X1 U7214 ( .A1(n6159), .A2(n6158), .B1(n6691), .B2(n6157), .ZN(n6160)
         );
  NAND2_X1 U7215 ( .A1(n6161), .A2(n6160), .ZN(n6193) );
  AOI22_X1 U7216 ( .A1(n6162), .A2(n6194), .B1(INSTQUEUE_REG_9__0__SCAN_IN), 
        .B2(n6193), .ZN(n6163) );
  OAI21_X1 U7217 ( .B1(n6196), .B2(n6602), .A(n6163), .ZN(n6164) );
  AOI21_X1 U7218 ( .B1(n6199), .B2(n6165), .A(n6164), .ZN(n6166) );
  OAI21_X1 U7219 ( .B1(n6201), .B2(n6220), .A(n6166), .ZN(U3092) );
  AOI22_X1 U7220 ( .A1(n6226), .A2(n6194), .B1(INSTQUEUE_REG_9__1__SCAN_IN), 
        .B2(n6193), .ZN(n6167) );
  OAI21_X1 U7221 ( .B1(n6196), .B2(n6168), .A(n6167), .ZN(n6169) );
  AOI21_X1 U7222 ( .B1(n6199), .B2(n6170), .A(n6169), .ZN(n6171) );
  OAI21_X1 U7223 ( .B1(n6201), .B2(n6228), .A(n6171), .ZN(U3093) );
  AOI22_X1 U7224 ( .A1(n6234), .A2(n6194), .B1(INSTQUEUE_REG_9__2__SCAN_IN), 
        .B2(n6193), .ZN(n6172) );
  OAI21_X1 U7225 ( .B1(n6196), .B2(n6173), .A(n6172), .ZN(n6174) );
  AOI21_X1 U7226 ( .B1(n6199), .B2(n6175), .A(n6174), .ZN(n6176) );
  OAI21_X1 U7227 ( .B1(n6201), .B2(n6236), .A(n6176), .ZN(U3094) );
  AOI22_X1 U7228 ( .A1(n6242), .A2(n6194), .B1(INSTQUEUE_REG_9__3__SCAN_IN), 
        .B2(n6193), .ZN(n6177) );
  OAI21_X1 U7229 ( .B1(n6196), .B2(n6609), .A(n6177), .ZN(n6178) );
  AOI21_X1 U7230 ( .B1(n6199), .B2(n6179), .A(n6178), .ZN(n6180) );
  OAI21_X1 U7231 ( .B1(n6201), .B2(n6244), .A(n6180), .ZN(U3095) );
  AOI22_X1 U7232 ( .A1(n6249), .A2(n6194), .B1(INSTQUEUE_REG_9__4__SCAN_IN), 
        .B2(n6193), .ZN(n6181) );
  OAI21_X1 U7233 ( .B1(n6196), .B2(n6616), .A(n6181), .ZN(n6182) );
  AOI21_X1 U7234 ( .B1(n6199), .B2(n6183), .A(n6182), .ZN(n6184) );
  OAI21_X1 U7235 ( .B1(n6201), .B2(n6251), .A(n6184), .ZN(U3096) );
  AOI22_X1 U7236 ( .A1(n6256), .A2(n6194), .B1(INSTQUEUE_REG_9__5__SCAN_IN), 
        .B2(n6193), .ZN(n6185) );
  OAI21_X1 U7237 ( .B1(n6196), .B2(n6623), .A(n6185), .ZN(n6186) );
  AOI21_X1 U7238 ( .B1(n6199), .B2(n6187), .A(n6186), .ZN(n6188) );
  OAI21_X1 U7239 ( .B1(n6201), .B2(n6258), .A(n6188), .ZN(U3097) );
  AOI22_X1 U7240 ( .A1(n6263), .A2(n6194), .B1(INSTQUEUE_REG_9__6__SCAN_IN), 
        .B2(n6193), .ZN(n6189) );
  OAI21_X1 U7241 ( .B1(n6196), .B2(n6630), .A(n6189), .ZN(n6190) );
  AOI21_X1 U7242 ( .B1(n6199), .B2(n6191), .A(n6190), .ZN(n6192) );
  OAI21_X1 U7243 ( .B1(n6201), .B2(n6265), .A(n6192), .ZN(U3098) );
  AOI22_X1 U7244 ( .A1(n6272), .A2(n6194), .B1(INSTQUEUE_REG_9__7__SCAN_IN), 
        .B2(n6193), .ZN(n6195) );
  OAI21_X1 U7245 ( .B1(n6196), .B2(n6642), .A(n6195), .ZN(n6197) );
  AOI21_X1 U7246 ( .B1(n6199), .B2(n6198), .A(n6197), .ZN(n6200) );
  OAI21_X1 U7247 ( .B1(n6201), .B2(n6274), .A(n6200), .ZN(U3099) );
  OAI21_X1 U7248 ( .B1(n6202), .B2(n6278), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6204) );
  OAI211_X1 U7249 ( .C1(n6206), .C2(n6205), .A(n6204), .B(n6203), .ZN(n6214)
         );
  NAND2_X1 U7250 ( .A1(n6208), .A2(n6207), .ZN(n6225) );
  INV_X1 U7251 ( .A(n6209), .ZN(n6210) );
  AOI21_X1 U7252 ( .B1(n6225), .B2(STATE2_REG_3__SCAN_IN), .A(n6210), .ZN(
        n6212) );
  NAND2_X1 U7253 ( .A1(n6270), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n6224)
         );
  NOR2_X1 U7254 ( .A1(n6216), .A2(n6215), .ZN(n6217) );
  AOI21_X1 U7255 ( .B1(n6219), .B2(n6218), .A(n6217), .ZN(n6275) );
  OAI22_X1 U7256 ( .A1(n6275), .A2(n6220), .B1(n6596), .B2(n6225), .ZN(n6221)
         );
  AOI21_X1 U7257 ( .B1(n6278), .B2(n6222), .A(n6221), .ZN(n6223) );
  OAI211_X1 U7258 ( .C1(n6281), .C2(n6597), .A(n6224), .B(n6223), .ZN(U3132)
         );
  NAND2_X1 U7259 ( .A1(n6270), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n6232)
         );
  INV_X1 U7260 ( .A(n6225), .ZN(n6271) );
  NAND2_X1 U7261 ( .A1(n6226), .A2(n6271), .ZN(n6227) );
  OAI21_X1 U7262 ( .B1(n6275), .B2(n6228), .A(n6227), .ZN(n6229) );
  AOI21_X1 U7263 ( .B1(n6278), .B2(n6230), .A(n6229), .ZN(n6231) );
  OAI211_X1 U7264 ( .C1(n6281), .C2(n6233), .A(n6232), .B(n6231), .ZN(U3133)
         );
  NAND2_X1 U7265 ( .A1(n6270), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n6240)
         );
  NAND2_X1 U7266 ( .A1(n6234), .A2(n6271), .ZN(n6235) );
  OAI21_X1 U7267 ( .B1(n6275), .B2(n6236), .A(n6235), .ZN(n6237) );
  AOI21_X1 U7268 ( .B1(n6278), .B2(n6238), .A(n6237), .ZN(n6239) );
  OAI211_X1 U7269 ( .C1(n6281), .C2(n6241), .A(n6240), .B(n6239), .ZN(U3134)
         );
  NAND2_X1 U7270 ( .A1(n6270), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n6248)
         );
  NAND2_X1 U7271 ( .A1(n6242), .A2(n6271), .ZN(n6243) );
  OAI21_X1 U7272 ( .B1(n6275), .B2(n6244), .A(n6243), .ZN(n6245) );
  AOI21_X1 U7273 ( .B1(n6278), .B2(n6246), .A(n6245), .ZN(n6247) );
  OAI211_X1 U7274 ( .C1(n6281), .C2(n6604), .A(n6248), .B(n6247), .ZN(U3135)
         );
  NAND2_X1 U7275 ( .A1(n6270), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n6255)
         );
  NAND2_X1 U7276 ( .A1(n6249), .A2(n6271), .ZN(n6250) );
  OAI21_X1 U7277 ( .B1(n6275), .B2(n6251), .A(n6250), .ZN(n6252) );
  AOI21_X1 U7278 ( .B1(n6278), .B2(n6253), .A(n6252), .ZN(n6254) );
  OAI211_X1 U7279 ( .C1(n6281), .C2(n6611), .A(n6255), .B(n6254), .ZN(U3136)
         );
  NAND2_X1 U7280 ( .A1(n6270), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n6262)
         );
  NAND2_X1 U7281 ( .A1(n6256), .A2(n6271), .ZN(n6257) );
  OAI21_X1 U7282 ( .B1(n6275), .B2(n6258), .A(n6257), .ZN(n6259) );
  AOI21_X1 U7283 ( .B1(n6278), .B2(n6260), .A(n6259), .ZN(n6261) );
  OAI211_X1 U7284 ( .C1(n6281), .C2(n6618), .A(n6262), .B(n6261), .ZN(U3137)
         );
  NAND2_X1 U7285 ( .A1(n6270), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n6269)
         );
  NAND2_X1 U7286 ( .A1(n6263), .A2(n6271), .ZN(n6264) );
  OAI21_X1 U7287 ( .B1(n6275), .B2(n6265), .A(n6264), .ZN(n6266) );
  AOI21_X1 U7288 ( .B1(n6278), .B2(n6267), .A(n6266), .ZN(n6268) );
  OAI211_X1 U7289 ( .C1(n6281), .C2(n6625), .A(n6269), .B(n6268), .ZN(U3138)
         );
  NAND2_X1 U7290 ( .A1(n6270), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n6280)
         );
  NAND2_X1 U7291 ( .A1(n6272), .A2(n6271), .ZN(n6273) );
  OAI21_X1 U7292 ( .B1(n6275), .B2(n6274), .A(n6273), .ZN(n6276) );
  AOI21_X1 U7293 ( .B1(n6278), .B2(n6277), .A(n6276), .ZN(n6279) );
  OAI211_X1 U7294 ( .C1(n6281), .C2(n6633), .A(n6280), .B(n6279), .ZN(U3139)
         );
  INV_X1 U7295 ( .A(n6282), .ZN(n6290) );
  INV_X1 U7296 ( .A(n6697), .ZN(n6284) );
  OAI21_X1 U7297 ( .B1(n6284), .B2(n6283), .A(n6650), .ZN(n6287) );
  OAI21_X1 U7298 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6824), .A(n6650), .ZN(
        n6643) );
  NOR2_X1 U7299 ( .A1(n6643), .A2(n6285), .ZN(n6286) );
  MUX2_X1 U7300 ( .A(n6287), .B(n6286), .S(STATE2_REG_0__SCAN_IN), .Z(n6289)
         );
  OAI211_X1 U7301 ( .C1(n6290), .C2(n6644), .A(n6289), .B(n6288), .ZN(U3148)
         );
  AND2_X1 U7302 ( .A1(n6439), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  OAI21_X1 U7303 ( .B1(n6294), .B2(n6293), .A(n3097), .ZN(U3455) );
  NOR2_X1 U7304 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6296) );
  OAI21_X1 U7305 ( .B1(n6296), .B2(D_C_N_REG_SCAN_IN), .A(n6855), .ZN(n6295)
         );
  OAI21_X1 U7306 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6855), .A(n6295), .ZN(
        U2791) );
  OAI21_X1 U7307 ( .B1(BS16_N), .B2(n6296), .A(n6680), .ZN(n6679) );
  OAI21_X1 U7308 ( .B1(n6680), .B2(n6297), .A(n6679), .ZN(U2792) );
  OAI21_X1 U7309 ( .B1(n6300), .B2(n6299), .A(n6298), .ZN(U2793) );
  NOR4_X1 U7310 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n6304) );
  NOR4_X1 U7311 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_17__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n6303) );
  NOR4_X1 U7312 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6302) );
  NOR4_X1 U7313 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6301) );
  NAND4_X1 U7314 ( .A1(n6304), .A2(n6303), .A3(n6302), .A4(n6301), .ZN(n6310)
         );
  NOR4_X1 U7315 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_5__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(
        n6308) );
  INV_X1 U7316 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6716) );
  INV_X1 U7317 ( .A(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6708) );
  NAND2_X1 U7318 ( .A1(n6716), .A2(n6708), .ZN(n6798) );
  AOI21_X1 U7319 ( .B1(DATAWIDTH_REG_1__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), .A(n6798), .ZN(n6307) );
  NOR4_X1 U7320 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n6306) );
  NOR4_X1 U7321 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_9__SCAN_IN), .A4(DATAWIDTH_REG_10__SCAN_IN), .ZN(
        n6305) );
  NAND4_X1 U7322 ( .A1(n6308), .A2(n6307), .A3(n6306), .A4(n6305), .ZN(n6309)
         );
  NOR2_X1 U7323 ( .A1(n6310), .A2(n6309), .ZN(n6685) );
  INV_X1 U7324 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6312) );
  NOR3_X1 U7325 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6313) );
  OAI21_X1 U7326 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6313), .A(n6685), .ZN(n6311)
         );
  OAI21_X1 U7327 ( .B1(n6685), .B2(n6312), .A(n6311), .ZN(U2794) );
  INV_X1 U7328 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6819) );
  AOI21_X1 U7329 ( .B1(n6681), .B2(n6819), .A(n6313), .ZN(n6315) );
  INV_X1 U7330 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6314) );
  INV_X1 U7331 ( .A(n6685), .ZN(n6688) );
  AOI22_X1 U7332 ( .A1(n6685), .A2(n6315), .B1(n6314), .B2(n6688), .ZN(U2795)
         );
  OAI21_X1 U7333 ( .B1(REIP_REG_15__SCAN_IN), .B2(n6333), .A(n6316), .ZN(n6317) );
  AOI22_X1 U7334 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6398), .B1(
        REIP_REG_16__SCAN_IN), .B2(n6317), .ZN(n6318) );
  OAI21_X1 U7335 ( .B1(REIP_REG_16__SCAN_IN), .B2(n6319), .A(n6318), .ZN(n6320) );
  AOI211_X1 U7336 ( .C1(n6394), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6378), 
        .B(n6320), .ZN(n6324) );
  INV_X1 U7337 ( .A(n6321), .ZN(n6411) );
  AOI22_X1 U7338 ( .A1(n6411), .A2(n6346), .B1(n6322), .B2(n6397), .ZN(n6323)
         );
  OAI211_X1 U7339 ( .C1(n6375), .C2(n6325), .A(n6324), .B(n6323), .ZN(U2811)
         );
  OAI22_X1 U7340 ( .A1(n6794), .A2(n6327), .B1(n6375), .B2(n6326), .ZN(n6328)
         );
  AOI211_X1 U7341 ( .C1(n6394), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6378), 
        .B(n6328), .ZN(n6339) );
  INV_X1 U7342 ( .A(n6329), .ZN(n6330) );
  AOI22_X1 U7343 ( .A1(n6331), .A2(n6346), .B1(n6330), .B2(n6397), .ZN(n6338)
         );
  NOR3_X1 U7344 ( .A1(n6333), .A2(REIP_REG_12__SCAN_IN), .A3(n6332), .ZN(n6342) );
  OAI21_X1 U7345 ( .B1(n6342), .B2(n6334), .A(REIP_REG_13__SCAN_IN), .ZN(n6337) );
  NAND3_X1 U7346 ( .A1(n6384), .A2(n6665), .A3(n6335), .ZN(n6336) );
  NAND4_X1 U7347 ( .A1(n6339), .A2(n6338), .A3(n6337), .A4(n6336), .ZN(U2814)
         );
  NOR2_X1 U7348 ( .A1(n6340), .A2(n6663), .ZN(n6341) );
  AOI211_X1 U7349 ( .C1(n6398), .C2(EBX_REG_12__SCAN_IN), .A(n6342), .B(n6341), 
        .ZN(n6348) );
  INV_X1 U7350 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6836) );
  NAND2_X1 U7351 ( .A1(n6343), .A2(n6399), .ZN(n6344) );
  OAI211_X1 U7352 ( .C1(n6836), .C2(n6376), .A(n6344), .B(n6365), .ZN(n6345)
         );
  AOI21_X1 U7353 ( .B1(n6418), .B2(n6346), .A(n6345), .ZN(n6347) );
  OAI211_X1 U7354 ( .C1(n6349), .C2(n5330), .A(n6348), .B(n6347), .ZN(U2815)
         );
  AOI22_X1 U7355 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6398), .B1(n6399), .B2(n6350), .ZN(n6361) );
  NOR3_X1 U7356 ( .A1(REIP_REG_10__SCAN_IN), .A2(n5810), .A3(n6351), .ZN(n6352) );
  AOI211_X1 U7357 ( .C1(n6394), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6378), 
        .B(n6352), .ZN(n6360) );
  OAI22_X1 U7358 ( .A1(n6354), .A2(n6371), .B1(n6353), .B2(n5330), .ZN(n6355)
         );
  INV_X1 U7359 ( .A(n6355), .ZN(n6359) );
  OAI21_X1 U7360 ( .B1(n6357), .B2(n6356), .A(REIP_REG_10__SCAN_IN), .ZN(n6358) );
  NAND4_X1 U7361 ( .A1(n6361), .A2(n6360), .A3(n6359), .A4(n6358), .ZN(U2817)
         );
  OAI22_X1 U7362 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6362), .B1(n6375), .B2(n6531), .ZN(n6363) );
  AOI21_X1 U7363 ( .B1(EBX_REG_7__SCAN_IN), .B2(n6398), .A(n6363), .ZN(n6370)
         );
  AOI21_X1 U7364 ( .B1(n6383), .B2(n6364), .A(n6661), .ZN(n6368) );
  INV_X1 U7365 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6366) );
  OAI21_X1 U7366 ( .B1(n6376), .B2(n6366), .A(n6365), .ZN(n6367) );
  NOR2_X1 U7367 ( .A1(n6368), .A2(n6367), .ZN(n6369) );
  OAI211_X1 U7368 ( .C1(n6479), .C2(n6371), .A(n6370), .B(n6369), .ZN(n6372)
         );
  INV_X1 U7369 ( .A(n6372), .ZN(n6373) );
  OAI21_X1 U7370 ( .B1(n6483), .B2(n5330), .A(n6373), .ZN(U2820) );
  AOI21_X1 U7371 ( .B1(REIP_REG_4__SCAN_IN), .B2(n6374), .A(
        REIP_REG_5__SCAN_IN), .ZN(n6382) );
  OAI22_X1 U7372 ( .A1(n3028), .A2(n6376), .B1(n6375), .B2(n6538), .ZN(n6377)
         );
  AOI211_X1 U7373 ( .C1(n6398), .C2(EBX_REG_5__SCAN_IN), .A(n6378), .B(n6377), 
        .ZN(n6381) );
  NOR2_X1 U7374 ( .A1(n5330), .A2(n6491), .ZN(n6379) );
  AOI21_X1 U7375 ( .B1(n6488), .B2(n6392), .A(n6379), .ZN(n6380) );
  OAI211_X1 U7376 ( .C1(n6383), .C2(n6382), .A(n6381), .B(n6380), .ZN(U2822)
         );
  NAND2_X1 U7377 ( .A1(n6384), .A2(REIP_REG_1__SCAN_IN), .ZN(n6386) );
  AOI21_X1 U7378 ( .B1(n6655), .B2(n6386), .A(n6385), .ZN(n6391) );
  NAND2_X1 U7379 ( .A1(n6399), .A2(n6574), .ZN(n6388) );
  AOI22_X1 U7380 ( .A1(EBX_REG_2__SCAN_IN), .A2(n6398), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n6394), .ZN(n6387) );
  OAI211_X1 U7381 ( .C1(n6389), .C2(n4534), .A(n6388), .B(n6387), .ZN(n6390)
         );
  AOI211_X1 U7382 ( .C1(n6506), .C2(n6392), .A(n6391), .B(n6390), .ZN(n6393)
         );
  OAI21_X1 U7383 ( .B1(n6509), .B2(n5330), .A(n6393), .ZN(U2825) );
  NAND2_X1 U7384 ( .A1(n6394), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6395)
         );
  AND2_X1 U7385 ( .A1(n6396), .A2(n6395), .ZN(n6408) );
  AOI22_X1 U7386 ( .A1(n6398), .A2(EBX_REG_1__SCAN_IN), .B1(n6397), .B2(n6821), 
        .ZN(n6403) );
  AOI22_X1 U7387 ( .A1(n6401), .A2(n6400), .B1(n6399), .B2(n4455), .ZN(n6402)
         );
  OAI211_X1 U7388 ( .C1(n6405), .C2(n6404), .A(n6403), .B(n6402), .ZN(n6406)
         );
  INV_X1 U7389 ( .A(n6406), .ZN(n6407) );
  OAI211_X1 U7390 ( .C1(n6409), .C2(n6681), .A(n6408), .B(n6407), .ZN(U2826)
         );
  AOI22_X1 U7391 ( .A1(n6411), .A2(n6417), .B1(n6410), .B2(DATAI_16_), .ZN(
        n6415) );
  AOI22_X1 U7392 ( .A1(n6413), .A2(DATAI_0_), .B1(n6412), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6414) );
  NAND2_X1 U7393 ( .A1(n6415), .A2(n6414), .ZN(U2875) );
  AOI22_X1 U7394 ( .A1(n6418), .A2(n6417), .B1(DATAI_12_), .B2(n6416), .ZN(
        n6419) );
  OAI21_X1 U7395 ( .B1(n6791), .B2(n6420), .A(n6419), .ZN(U2879) );
  INV_X1 U7396 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6474) );
  AOI22_X1 U7397 ( .A1(n6449), .A2(LWORD_REG_15__SCAN_IN), .B1(n6439), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6422) );
  OAI21_X1 U7398 ( .B1(n6474), .B2(n6451), .A(n6422), .ZN(U2908) );
  AOI22_X1 U7399 ( .A1(n6449), .A2(LWORD_REG_14__SCAN_IN), .B1(n6439), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6423) );
  OAI21_X1 U7400 ( .B1(n5186), .B2(n6451), .A(n6423), .ZN(U2909) );
  AOI22_X1 U7401 ( .A1(n6449), .A2(LWORD_REG_13__SCAN_IN), .B1(n6439), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6424) );
  OAI21_X1 U7402 ( .B1(n6425), .B2(n6451), .A(n6424), .ZN(U2910) );
  AOI22_X1 U7403 ( .A1(n6449), .A2(LWORD_REG_12__SCAN_IN), .B1(n6439), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6426) );
  OAI21_X1 U7404 ( .B1(n6791), .B2(n6451), .A(n6426), .ZN(U2911) );
  INV_X1 U7405 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6428) );
  AOI22_X1 U7406 ( .A1(n6436), .A2(LWORD_REG_11__SCAN_IN), .B1(n6439), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6427) );
  OAI21_X1 U7407 ( .B1(n6428), .B2(n6451), .A(n6427), .ZN(U2912) );
  INV_X1 U7408 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6430) );
  AOI22_X1 U7409 ( .A1(n6436), .A2(LWORD_REG_10__SCAN_IN), .B1(n6439), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6429) );
  OAI21_X1 U7410 ( .B1(n6430), .B2(n6451), .A(n6429), .ZN(U2913) );
  INV_X1 U7411 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6432) );
  AOI22_X1 U7412 ( .A1(n6436), .A2(LWORD_REG_9__SCAN_IN), .B1(n6439), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6431) );
  OAI21_X1 U7413 ( .B1(n6432), .B2(n6451), .A(n6431), .ZN(U2914) );
  AOI22_X1 U7414 ( .A1(n6436), .A2(LWORD_REG_8__SCAN_IN), .B1(n6439), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6433) );
  OAI21_X1 U7415 ( .B1(n6717), .B2(n6451), .A(n6433), .ZN(U2915) );
  AOI22_X1 U7416 ( .A1(n6436), .A2(LWORD_REG_7__SCAN_IN), .B1(n6439), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6434) );
  OAI21_X1 U7417 ( .B1(n6435), .B2(n6451), .A(n6434), .ZN(U2916) );
  AOI22_X1 U7418 ( .A1(n6436), .A2(LWORD_REG_6__SCAN_IN), .B1(n6439), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6437) );
  OAI21_X1 U7419 ( .B1(n4776), .B2(n6451), .A(n6437), .ZN(U2917) );
  AOI22_X1 U7420 ( .A1(n6449), .A2(LWORD_REG_5__SCAN_IN), .B1(n6439), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6438) );
  OAI21_X1 U7421 ( .B1(n4784), .B2(n6451), .A(n6438), .ZN(U2918) );
  AOI22_X1 U7422 ( .A1(n6449), .A2(LWORD_REG_4__SCAN_IN), .B1(n6439), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6440) );
  OAI21_X1 U7423 ( .B1(n6441), .B2(n6451), .A(n6440), .ZN(U2919) );
  AOI22_X1 U7424 ( .A1(n6449), .A2(LWORD_REG_3__SCAN_IN), .B1(n6448), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6442) );
  OAI21_X1 U7425 ( .B1(n6443), .B2(n6451), .A(n6442), .ZN(U2920) );
  AOI22_X1 U7426 ( .A1(n6449), .A2(LWORD_REG_2__SCAN_IN), .B1(n6448), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6444) );
  OAI21_X1 U7427 ( .B1(n6445), .B2(n6451), .A(n6444), .ZN(U2921) );
  AOI22_X1 U7428 ( .A1(n6449), .A2(LWORD_REG_1__SCAN_IN), .B1(n6448), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6446) );
  OAI21_X1 U7429 ( .B1(n6447), .B2(n6451), .A(n6446), .ZN(U2922) );
  AOI22_X1 U7430 ( .A1(n6449), .A2(LWORD_REG_0__SCAN_IN), .B1(n6448), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6450) );
  OAI21_X1 U7431 ( .B1(n6452), .B2(n6451), .A(n6450), .ZN(U2923) );
  AOI22_X1 U7432 ( .A1(EAX_REG_25__SCAN_IN), .A2(n6467), .B1(n6471), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n6453) );
  NAND2_X1 U7433 ( .A1(n6470), .A2(DATAI_9_), .ZN(n6458) );
  NAND2_X1 U7434 ( .A1(n6453), .A2(n6458), .ZN(U2933) );
  AOI22_X1 U7435 ( .A1(EAX_REG_26__SCAN_IN), .A2(n6467), .B1(n6464), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n6454) );
  NAND2_X1 U7436 ( .A1(n6470), .A2(DATAI_10_), .ZN(n6460) );
  NAND2_X1 U7437 ( .A1(n6454), .A2(n6460), .ZN(U2934) );
  AOI22_X1 U7438 ( .A1(EAX_REG_27__SCAN_IN), .A2(n6467), .B1(n6464), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n6455) );
  NAND2_X1 U7439 ( .A1(n6470), .A2(DATAI_11_), .ZN(n6462) );
  NAND2_X1 U7440 ( .A1(n6455), .A2(n6462), .ZN(U2935) );
  AOI22_X1 U7441 ( .A1(EAX_REG_28__SCAN_IN), .A2(n6467), .B1(n6464), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n6456) );
  NAND2_X1 U7442 ( .A1(n6470), .A2(DATAI_12_), .ZN(n6465) );
  NAND2_X1 U7443 ( .A1(n6456), .A2(n6465), .ZN(U2936) );
  AOI22_X1 U7444 ( .A1(EAX_REG_30__SCAN_IN), .A2(n6467), .B1(n6464), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n6457) );
  NAND2_X1 U7445 ( .A1(n6470), .A2(DATAI_14_), .ZN(n6468) );
  NAND2_X1 U7446 ( .A1(n6457), .A2(n6468), .ZN(U2938) );
  AOI22_X1 U7447 ( .A1(EAX_REG_9__SCAN_IN), .A2(n6467), .B1(n6471), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n6459) );
  NAND2_X1 U7448 ( .A1(n6459), .A2(n6458), .ZN(U2948) );
  AOI22_X1 U7449 ( .A1(EAX_REG_10__SCAN_IN), .A2(n6467), .B1(n6464), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n6461) );
  NAND2_X1 U7450 ( .A1(n6461), .A2(n6460), .ZN(U2949) );
  AOI22_X1 U7451 ( .A1(EAX_REG_11__SCAN_IN), .A2(n6467), .B1(n6464), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U7452 ( .A1(n6463), .A2(n6462), .ZN(U2950) );
  AOI22_X1 U7453 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6467), .B1(n6464), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n6466) );
  NAND2_X1 U7454 ( .A1(n6466), .A2(n6465), .ZN(U2951) );
  AOI22_X1 U7455 ( .A1(EAX_REG_14__SCAN_IN), .A2(n6467), .B1(n6471), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n6469) );
  NAND2_X1 U7456 ( .A1(n6469), .A2(n6468), .ZN(U2953) );
  AOI22_X1 U7457 ( .A1(n6471), .A2(LWORD_REG_15__SCAN_IN), .B1(n6470), .B2(
        DATAI_15_), .ZN(n6472) );
  OAI21_X1 U7458 ( .B1(n6474), .B2(n6473), .A(n6472), .ZN(U2954) );
  AOI22_X1 U7459 ( .A1(n6501), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .B1(n6573), 
        .B2(REIP_REG_7__SCAN_IN), .ZN(n6482) );
  OAI21_X1 U7460 ( .B1(n6475), .B2(n6477), .A(n2955), .ZN(n6478) );
  INV_X1 U7461 ( .A(n6478), .ZN(n6532) );
  INV_X1 U7462 ( .A(n6479), .ZN(n6480) );
  AOI22_X1 U7463 ( .A1(n6532), .A2(n6505), .B1(n5795), .B2(n6480), .ZN(n6481)
         );
  OAI211_X1 U7464 ( .C1(n6510), .C2(n6483), .A(n6482), .B(n6481), .ZN(U2979)
         );
  AND2_X1 U7465 ( .A1(n6573), .A2(REIP_REG_5__SCAN_IN), .ZN(n6539) );
  AOI21_X1 U7466 ( .B1(n6501), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n6539), 
        .ZN(n6490) );
  OR2_X1 U7467 ( .A1(n6485), .A2(n6484), .ZN(n6486) );
  AND2_X1 U7468 ( .A1(n6487), .A2(n6486), .ZN(n6543) );
  AOI22_X1 U7469 ( .A1(n6543), .A2(n6505), .B1(n5795), .B2(n6488), .ZN(n6489)
         );
  OAI211_X1 U7470 ( .C1(n6510), .C2(n6491), .A(n6490), .B(n6489), .ZN(U2981)
         );
  AND2_X1 U7471 ( .A1(n6573), .A2(REIP_REG_3__SCAN_IN), .ZN(n6562) );
  AOI21_X1 U7472 ( .B1(n6501), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n6562), 
        .ZN(n6499) );
  XNOR2_X1 U7473 ( .A(n6492), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6496)
         );
  INV_X1 U7474 ( .A(n6503), .ZN(n6493) );
  OAI21_X1 U7475 ( .B1(n6493), .B2(n6789), .A(n2963), .ZN(n6494) );
  OAI21_X1 U7476 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6503), .A(n6494), 
        .ZN(n6495) );
  XNOR2_X1 U7477 ( .A(n6496), .B(n6495), .ZN(n6564) );
  AOI22_X1 U7478 ( .A1(n6497), .A2(n5795), .B1(n6505), .B2(n6564), .ZN(n6498)
         );
  OAI211_X1 U7479 ( .C1(n6510), .C2(n6500), .A(n6499), .B(n6498), .ZN(U2983)
         );
  AOI22_X1 U7480 ( .A1(n6501), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n6573), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6508) );
  XNOR2_X1 U7481 ( .A(n2963), .B(n6789), .ZN(n6504) );
  XNOR2_X1 U7482 ( .A(n6504), .B(n6503), .ZN(n6580) );
  AOI22_X1 U7483 ( .A1(n6506), .A2(n5795), .B1(n6580), .B2(n6505), .ZN(n6507)
         );
  OAI211_X1 U7484 ( .C1(n6510), .C2(n6509), .A(n6508), .B(n6507), .ZN(U2984)
         );
  INV_X1 U7485 ( .A(n6511), .ZN(n6518) );
  AOI21_X1 U7486 ( .B1(n6513), .B2(n4314), .A(n6512), .ZN(n6517) );
  AOI22_X1 U7487 ( .A1(n6515), .A2(n6579), .B1(n6514), .B2(n5807), .ZN(n6516)
         );
  OAI211_X1 U7488 ( .C1(n6518), .C2(n5807), .A(n6517), .B(n6516), .ZN(U3009)
         );
  AOI211_X1 U7489 ( .C1(n6536), .C2(n6530), .A(n6519), .B(n6537), .ZN(n6528)
         );
  NOR2_X1 U7490 ( .A1(n6521), .A2(n6520), .ZN(n6527) );
  NAND2_X1 U7491 ( .A1(n6541), .A2(n6522), .ZN(n6523) );
  OAI21_X1 U7492 ( .B1(n6525), .B2(n6524), .A(n6523), .ZN(n6526) );
  NOR3_X1 U7493 ( .A1(n6528), .A2(n6527), .A3(n6526), .ZN(n6529) );
  OAI21_X1 U7494 ( .B1(n6535), .B2(n6530), .A(n6529), .ZN(U3010) );
  INV_X1 U7495 ( .A(n6531), .ZN(n6533) );
  AOI222_X1 U7496 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6573), .B1(n6541), .B2(
        n6533), .C1(n6579), .C2(n6532), .ZN(n6534) );
  OAI221_X1 U7497 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n6537), .C1(n6536), .C2(n6535), .A(n6534), .ZN(U3011) );
  INV_X1 U7498 ( .A(n6538), .ZN(n6540) );
  AOI21_X1 U7499 ( .B1(n6541), .B2(n6540), .A(n6539), .ZN(n6551) );
  OAI21_X1 U7500 ( .B1(n6577), .B2(n6542), .A(n6546), .ZN(n6544) );
  AOI22_X1 U7501 ( .A1(n6545), .A2(n6544), .B1(n6579), .B2(n6543), .ZN(n6550)
         );
  NAND3_X1 U7502 ( .A1(n6548), .A2(n6547), .A3(n6546), .ZN(n6549) );
  NAND3_X1 U7503 ( .A1(n6551), .A2(n6550), .A3(n6549), .ZN(U3013) );
  AOI21_X1 U7504 ( .B1(n6541), .B2(n6553), .A(n6552), .ZN(n6560) );
  OAI21_X1 U7505 ( .B1(n6555), .B2(n6577), .A(n6582), .ZN(n6561) );
  AOI22_X1 U7506 ( .A1(n6561), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .B1(n6579), 
        .B2(n6554), .ZN(n6559) );
  INV_X1 U7507 ( .A(n6555), .ZN(n6572) );
  NOR2_X1 U7508 ( .A1(n6572), .A2(n6556), .ZN(n6565) );
  OAI211_X1 U7509 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6565), .B(n6557), .ZN(n6558) );
  NAND3_X1 U7510 ( .A1(n6560), .A2(n6559), .A3(n6558), .ZN(U3014) );
  INV_X1 U7511 ( .A(n6561), .ZN(n6569) );
  AOI21_X1 U7512 ( .B1(n4314), .B2(n6563), .A(n6562), .ZN(n6567) );
  AOI22_X1 U7513 ( .A1(n6565), .A2(n6568), .B1(n6579), .B2(n6564), .ZN(n6566)
         );
  OAI211_X1 U7514 ( .C1(n6569), .C2(n6568), .A(n6567), .B(n6566), .ZN(U3015)
         );
  NAND2_X1 U7515 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6570), .ZN(n6583)
         );
  AOI21_X1 U7516 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n3443), .A(n6572), 
        .ZN(n6576) );
  AOI22_X1 U7517 ( .A1(n6541), .A2(n6574), .B1(n6573), .B2(REIP_REG_2__SCAN_IN), .ZN(n6575) );
  OAI21_X1 U7518 ( .B1(n6577), .B2(n6576), .A(n6575), .ZN(n6578) );
  AOI21_X1 U7519 ( .B1(n6580), .B2(n6579), .A(n6578), .ZN(n6581) );
  OAI221_X1 U7520 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6583), .C1(n6789), .C2(n6582), .A(n6581), .ZN(U3016) );
  NOR2_X1 U7521 ( .A1(n3545), .A2(n6584), .ZN(U3019) );
  OAI22_X1 U7522 ( .A1(n6589), .A2(n6611), .B1(n6610), .B2(n6588), .ZN(n6585)
         );
  INV_X1 U7523 ( .A(n6585), .ZN(n6587) );
  AOI22_X1 U7524 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6592), .B1(n6613), 
        .B2(n6591), .ZN(n6586) );
  OAI211_X1 U7525 ( .C1(n6595), .C2(n6616), .A(n6587), .B(n6586), .ZN(U3048)
         );
  OAI22_X1 U7526 ( .A1(n6589), .A2(n6625), .B1(n6624), .B2(n6588), .ZN(n6590)
         );
  INV_X1 U7527 ( .A(n6590), .ZN(n6594) );
  AOI22_X1 U7528 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6592), .B1(n6627), 
        .B2(n6591), .ZN(n6593) );
  OAI211_X1 U7529 ( .C1(n6595), .C2(n6630), .A(n6594), .B(n6593), .ZN(U3050)
         );
  OAI22_X1 U7530 ( .A1(n6634), .A2(n6597), .B1(n6596), .B2(n6631), .ZN(n6598)
         );
  INV_X1 U7531 ( .A(n6598), .ZN(n6601) );
  AOI22_X1 U7532 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6638), .B1(n6599), 
        .B2(n6636), .ZN(n6600) );
  OAI211_X1 U7533 ( .C1(n6602), .C2(n6641), .A(n6601), .B(n6600), .ZN(U3108)
         );
  OAI22_X1 U7534 ( .A1(n6634), .A2(n6604), .B1(n6603), .B2(n6631), .ZN(n6605)
         );
  INV_X1 U7535 ( .A(n6605), .ZN(n6608) );
  AOI22_X1 U7536 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6638), .B1(n6606), 
        .B2(n6636), .ZN(n6607) );
  OAI211_X1 U7537 ( .C1(n6609), .C2(n6641), .A(n6608), .B(n6607), .ZN(U3111)
         );
  OAI22_X1 U7538 ( .A1(n6634), .A2(n6611), .B1(n6610), .B2(n6631), .ZN(n6612)
         );
  INV_X1 U7539 ( .A(n6612), .ZN(n6615) );
  AOI22_X1 U7540 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6638), .B1(n6613), 
        .B2(n6636), .ZN(n6614) );
  OAI211_X1 U7541 ( .C1(n6616), .C2(n6641), .A(n6615), .B(n6614), .ZN(U3112)
         );
  OAI22_X1 U7542 ( .A1(n6634), .A2(n6618), .B1(n6617), .B2(n6631), .ZN(n6619)
         );
  INV_X1 U7543 ( .A(n6619), .ZN(n6622) );
  AOI22_X1 U7544 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6638), .B1(n6620), 
        .B2(n6636), .ZN(n6621) );
  OAI211_X1 U7545 ( .C1(n6623), .C2(n6641), .A(n6622), .B(n6621), .ZN(U3113)
         );
  OAI22_X1 U7546 ( .A1(n6634), .A2(n6625), .B1(n6624), .B2(n6631), .ZN(n6626)
         );
  INV_X1 U7547 ( .A(n6626), .ZN(n6629) );
  AOI22_X1 U7548 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6638), .B1(n6627), 
        .B2(n6636), .ZN(n6628) );
  OAI211_X1 U7549 ( .C1(n6630), .C2(n6641), .A(n6629), .B(n6628), .ZN(U3114)
         );
  OAI22_X1 U7550 ( .A1(n6634), .A2(n6633), .B1(n6632), .B2(n6631), .ZN(n6635)
         );
  INV_X1 U7551 ( .A(n6635), .ZN(n6640) );
  AOI22_X1 U7552 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6638), .B1(n6637), 
        .B2(n6636), .ZN(n6639) );
  OAI211_X1 U7553 ( .C1(n6642), .C2(n6641), .A(n6640), .B(n6639), .ZN(U3115)
         );
  OAI211_X1 U7554 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(n6643), .B(STATE2_REG_1__SCAN_IN), .ZN(n6652) );
  OAI21_X1 U7555 ( .B1(n6646), .B2(n6645), .A(n6644), .ZN(n6649) );
  INV_X1 U7556 ( .A(n6647), .ZN(n6648) );
  AOI21_X1 U7557 ( .B1(n6650), .B2(n6649), .A(n6648), .ZN(n6651) );
  NAND2_X1 U7558 ( .A1(n6652), .A2(n6651), .ZN(U3149) );
  AND2_X1 U7559 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6677), .ZN(U3151) );
  AND2_X1 U7560 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6677), .ZN(U3152) );
  AND2_X1 U7561 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6677), .ZN(U3153) );
  AND2_X1 U7562 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6677), .ZN(U3154) );
  AND2_X1 U7563 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6677), .ZN(U3155) );
  AND2_X1 U7564 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6677), .ZN(U3156) );
  AND2_X1 U7565 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6677), .ZN(U3157) );
  AND2_X1 U7566 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6677), .ZN(U3158) );
  AND2_X1 U7567 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6677), .ZN(U3159) );
  AND2_X1 U7568 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6677), .ZN(U3160) );
  AND2_X1 U7569 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6677), .ZN(U3161) );
  AND2_X1 U7570 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6677), .ZN(U3162) );
  AND2_X1 U7571 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6677), .ZN(U3163) );
  AND2_X1 U7572 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6677), .ZN(U3164) );
  AND2_X1 U7573 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6677), .ZN(U3165) );
  AND2_X1 U7574 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6677), .ZN(U3166) );
  AND2_X1 U7575 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6677), .ZN(U3167) );
  AND2_X1 U7576 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6677), .ZN(U3168) );
  AND2_X1 U7577 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6677), .ZN(U3169) );
  NOR2_X1 U7578 ( .A1(n6680), .A2(n6716), .ZN(U3170) );
  AND2_X1 U7579 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6677), .ZN(U3171) );
  AND2_X1 U7580 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6677), .ZN(U3172) );
  AND2_X1 U7581 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6677), .ZN(U3173) );
  AND2_X1 U7582 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6677), .ZN(U3174) );
  AND2_X1 U7583 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6677), .ZN(U3175) );
  AND2_X1 U7584 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6677), .ZN(U3176) );
  AND2_X1 U7585 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6677), .ZN(U3177) );
  AND2_X1 U7586 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6677), .ZN(U3178) );
  NOR2_X1 U7587 ( .A1(n6680), .A2(n6708), .ZN(U3179) );
  AND2_X1 U7588 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6677), .ZN(U3180) );
  AOI22_X1 U7589 ( .A1(n6857), .A2(REIP_REG_1__SCAN_IN), .B1(n6855), .B2(
        ADDRESS_REG_0__SCAN_IN), .ZN(n6654) );
  OAI21_X1 U7590 ( .B1(n6655), .B2(n6674), .A(n6654), .ZN(U3184) );
  AOI22_X1 U7591 ( .A1(n6857), .A2(REIP_REG_3__SCAN_IN), .B1(n6855), .B2(
        ADDRESS_REG_2__SCAN_IN), .ZN(n6656) );
  OAI21_X1 U7592 ( .B1(n6657), .B2(n6674), .A(n6656), .ZN(U3186) );
  AOI22_X1 U7593 ( .A1(n6857), .A2(REIP_REG_5__SCAN_IN), .B1(n6855), .B2(
        ADDRESS_REG_4__SCAN_IN), .ZN(n6658) );
  OAI21_X1 U7594 ( .B1(n6659), .B2(n6674), .A(n6658), .ZN(U3188) );
  AOI22_X1 U7595 ( .A1(n6857), .A2(REIP_REG_6__SCAN_IN), .B1(n6855), .B2(
        ADDRESS_REG_5__SCAN_IN), .ZN(n6660) );
  OAI21_X1 U7596 ( .B1(n6661), .B2(n6674), .A(n6660), .ZN(U3189) );
  AOI22_X1 U7597 ( .A1(n6857), .A2(REIP_REG_11__SCAN_IN), .B1(n6855), .B2(
        ADDRESS_REG_10__SCAN_IN), .ZN(n6662) );
  OAI21_X1 U7598 ( .B1(n6663), .B2(n6674), .A(n6662), .ZN(U3194) );
  AOI22_X1 U7599 ( .A1(n6857), .A2(REIP_REG_12__SCAN_IN), .B1(n6855), .B2(
        ADDRESS_REG_11__SCAN_IN), .ZN(n6664) );
  OAI21_X1 U7600 ( .B1(n6665), .B2(n6674), .A(n6664), .ZN(U3195) );
  AOI22_X1 U7601 ( .A1(n6857), .A2(REIP_REG_18__SCAN_IN), .B1(n6855), .B2(
        ADDRESS_REG_17__SCAN_IN), .ZN(n6666) );
  OAI21_X1 U7602 ( .B1(n5448), .B2(n6674), .A(n6666), .ZN(U3201) );
  AOI22_X1 U7603 ( .A1(n6857), .A2(REIP_REG_19__SCAN_IN), .B1(n6855), .B2(
        ADDRESS_REG_18__SCAN_IN), .ZN(n6667) );
  OAI21_X1 U7604 ( .B1(n6668), .B2(n6674), .A(n6667), .ZN(U3202) );
  AOI22_X1 U7605 ( .A1(n6857), .A2(REIP_REG_20__SCAN_IN), .B1(n6855), .B2(
        ADDRESS_REG_19__SCAN_IN), .ZN(n6669) );
  OAI21_X1 U7606 ( .B1(n6670), .B2(n6674), .A(n6669), .ZN(U3203) );
  AOI22_X1 U7607 ( .A1(n6857), .A2(REIP_REG_23__SCAN_IN), .B1(n6855), .B2(
        ADDRESS_REG_22__SCAN_IN), .ZN(n6671) );
  OAI21_X1 U7608 ( .B1(n6800), .B2(n6674), .A(n6671), .ZN(U3206) );
  AOI22_X1 U7609 ( .A1(n6857), .A2(REIP_REG_25__SCAN_IN), .B1(n6855), .B2(
        ADDRESS_REG_24__SCAN_IN), .ZN(n6672) );
  OAI21_X1 U7610 ( .B1(n6799), .B2(n6674), .A(n6672), .ZN(U3208) );
  AOI22_X1 U7611 ( .A1(n6857), .A2(REIP_REG_30__SCAN_IN), .B1(n6855), .B2(
        ADDRESS_REG_29__SCAN_IN), .ZN(n6673) );
  OAI21_X1 U7612 ( .B1(n6675), .B2(n6674), .A(n6673), .ZN(U3213) );
  MUX2_X1 U7613 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6702), .Z(U3445) );
  MUX2_X1 U7614 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6702), .Z(U3446) );
  MUX2_X1 U7615 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6702), .Z(U3447) );
  MUX2_X1 U7616 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6702), .Z(U3448) );
  INV_X1 U7617 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6678) );
  INV_X1 U7618 ( .A(n6679), .ZN(n6676) );
  AOI21_X1 U7619 ( .B1(n6678), .B2(n6677), .A(n6676), .ZN(U3451) );
  OAI21_X1 U7620 ( .B1(n6680), .B2(n6819), .A(n6679), .ZN(U3452) );
  AOI21_X1 U7621 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6682) );
  AOI22_X1 U7622 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6682), .B2(n6681), .ZN(n6684) );
  INV_X1 U7623 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6683) );
  AOI22_X1 U7624 ( .A1(n6685), .A2(n6684), .B1(n6683), .B2(n6688), .ZN(U3468)
         );
  INV_X1 U7625 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6689) );
  INV_X1 U7626 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6687) );
  NOR2_X1 U7627 ( .A1(n6688), .A2(REIP_REG_1__SCAN_IN), .ZN(n6686) );
  AOI22_X1 U7628 ( .A1(n6689), .A2(n6688), .B1(n6687), .B2(n6686), .ZN(U3469)
         );
  NAND2_X1 U7629 ( .A1(n6855), .A2(W_R_N_REG_SCAN_IN), .ZN(n6690) );
  OAI21_X1 U7630 ( .B1(n6855), .B2(READREQUEST_REG_SCAN_IN), .A(n6690), .ZN(
        U3470) );
  OAI211_X1 U7631 ( .C1(READY_N), .C2(n6693), .A(n6692), .B(n6691), .ZN(n6694)
         );
  NOR2_X1 U7632 ( .A1(n6695), .A2(n6694), .ZN(n6701) );
  OAI211_X1 U7633 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n3411), .A(n6696), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6698) );
  AOI21_X1 U7634 ( .B1(n6698), .B2(STATE2_REG_0__SCAN_IN), .A(n6697), .ZN(
        n6700) );
  NAND2_X1 U7635 ( .A1(n6701), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6699) );
  OAI21_X1 U7636 ( .B1(n6701), .B2(n6700), .A(n6699), .ZN(U3472) );
  MUX2_X1 U7637 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6702), .Z(U3473) );
  OAI22_X1 U7638 ( .A1(n3031), .A2(keyinput58), .B1(n6704), .B2(keyinput22), 
        .ZN(n6703) );
  AOI221_X1 U7639 ( .B1(n3031), .B2(keyinput58), .C1(keyinput22), .C2(n6704), 
        .A(n6703), .ZN(n6715) );
  INV_X1 U7640 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n6706) );
  OAI22_X1 U7641 ( .A1(n5448), .A2(keyinput42), .B1(n6706), .B2(keyinput56), 
        .ZN(n6705) );
  AOI221_X1 U7642 ( .B1(n5448), .B2(keyinput42), .C1(keyinput56), .C2(n6706), 
        .A(n6705), .ZN(n6714) );
  OAI22_X1 U7643 ( .A1(n6800), .A2(keyinput48), .B1(n6708), .B2(keyinput44), 
        .ZN(n6707) );
  AOI221_X1 U7644 ( .B1(n6800), .B2(keyinput48), .C1(keyinput44), .C2(n6708), 
        .A(n6707), .ZN(n6713) );
  INV_X1 U7645 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n6711) );
  OAI22_X1 U7646 ( .A1(n6711), .A2(keyinput47), .B1(n6710), .B2(keyinput57), 
        .ZN(n6709) );
  AOI221_X1 U7647 ( .B1(n6711), .B2(keyinput47), .C1(keyinput57), .C2(n6710), 
        .A(n6709), .ZN(n6712) );
  NAND4_X1 U7648 ( .A1(n6715), .A2(n6714), .A3(n6713), .A4(n6712), .ZN(n6854)
         );
  XNOR2_X1 U7649 ( .A(n6716), .B(keyinput62), .ZN(n6721) );
  XOR2_X1 U7650 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .B(keyinput8), .Z(n6720) );
  XNOR2_X1 U7651 ( .A(n3515), .B(keyinput28), .ZN(n6719) );
  XNOR2_X1 U7652 ( .A(keyinput39), .B(n6717), .ZN(n6718) );
  NOR4_X1 U7653 ( .A1(n6721), .A2(n6720), .A3(n6719), .A4(n6718), .ZN(n6729)
         );
  OAI22_X1 U7654 ( .A1(n6799), .A2(keyinput18), .B1(n6723), .B2(keyinput53), 
        .ZN(n6722) );
  AOI221_X1 U7655 ( .B1(n6799), .B2(keyinput18), .C1(keyinput53), .C2(n6723), 
        .A(n6722), .ZN(n6728) );
  INV_X1 U7656 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n6725) );
  OAI22_X1 U7657 ( .A1(n6726), .A2(keyinput54), .B1(n6725), .B2(keyinput29), 
        .ZN(n6724) );
  AOI221_X1 U7658 ( .B1(n6726), .B2(keyinput54), .C1(keyinput29), .C2(n6725), 
        .A(n6724), .ZN(n6727) );
  NAND3_X1 U7659 ( .A1(n6729), .A2(n6728), .A3(n6727), .ZN(n6853) );
  INV_X1 U7660 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n6732) );
  AOI22_X1 U7661 ( .A1(n6732), .A2(keyinput60), .B1(n6731), .B2(keyinput51), 
        .ZN(n6730) );
  OAI221_X1 U7662 ( .B1(n6732), .B2(keyinput60), .C1(n6731), .C2(keyinput51), 
        .A(n6730), .ZN(n6740) );
  INV_X1 U7663 ( .A(EAX_REG_31__SCAN_IN), .ZN(n6795) );
  AOI22_X1 U7664 ( .A1(n6795), .A2(keyinput24), .B1(keyinput23), .B2(n6734), 
        .ZN(n6733) );
  OAI221_X1 U7665 ( .B1(n6795), .B2(keyinput24), .C1(n6734), .C2(keyinput23), 
        .A(n6733), .ZN(n6739) );
  INV_X1 U7666 ( .A(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n6796) );
  AOI22_X1 U7667 ( .A1(n6796), .A2(keyinput46), .B1(keyinput19), .B2(n5100), 
        .ZN(n6735) );
  OAI221_X1 U7668 ( .B1(n6796), .B2(keyinput46), .C1(n5100), .C2(keyinput19), 
        .A(n6735), .ZN(n6738) );
  AOI22_X1 U7669 ( .A1(n4475), .A2(keyinput1), .B1(n6789), .B2(keyinput43), 
        .ZN(n6736) );
  OAI221_X1 U7670 ( .B1(n4475), .B2(keyinput1), .C1(n6789), .C2(keyinput43), 
        .A(n6736), .ZN(n6737) );
  NOR4_X1 U7671 ( .A1(n6740), .A2(n6739), .A3(n6738), .A4(n6737), .ZN(n6778)
         );
  INV_X1 U7672 ( .A(UWORD_REG_13__SCAN_IN), .ZN(n6742) );
  AOI22_X1 U7673 ( .A1(n6743), .A2(keyinput2), .B1(keyinput34), .B2(n6742), 
        .ZN(n6741) );
  OAI221_X1 U7674 ( .B1(n6743), .B2(keyinput2), .C1(n6742), .C2(keyinput34), 
        .A(n6741), .ZN(n6751) );
  AOI22_X1 U7675 ( .A1(n6794), .A2(keyinput32), .B1(keyinput16), .B2(n6792), 
        .ZN(n6744) );
  OAI221_X1 U7676 ( .B1(n6794), .B2(keyinput32), .C1(n6792), .C2(keyinput16), 
        .A(n6744), .ZN(n6750) );
  AOI22_X1 U7677 ( .A1(n6793), .A2(keyinput9), .B1(keyinput14), .B2(n6791), 
        .ZN(n6745) );
  OAI221_X1 U7678 ( .B1(n6793), .B2(keyinput9), .C1(n6791), .C2(keyinput14), 
        .A(n6745), .ZN(n6749) );
  XNOR2_X1 U7679 ( .A(INSTQUEUE_REG_9__2__SCAN_IN), .B(keyinput33), .ZN(n6747)
         );
  XNOR2_X1 U7680 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .B(keyinput61), .ZN(n6746) );
  NAND2_X1 U7681 ( .A1(n6747), .A2(n6746), .ZN(n6748) );
  NOR4_X1 U7682 ( .A1(n6751), .A2(n6750), .A3(n6749), .A4(n6748), .ZN(n6777)
         );
  INV_X1 U7683 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n6782) );
  AOI22_X1 U7684 ( .A1(n6782), .A2(keyinput50), .B1(keyinput31), .B2(n6781), 
        .ZN(n6752) );
  OAI221_X1 U7685 ( .B1(n6782), .B2(keyinput50), .C1(n6781), .C2(keyinput31), 
        .A(n6752), .ZN(n6762) );
  AOI22_X1 U7686 ( .A1(n6754), .A2(keyinput26), .B1(n4712), .B2(keyinput7), 
        .ZN(n6753) );
  OAI221_X1 U7687 ( .B1(n6754), .B2(keyinput26), .C1(n4712), .C2(keyinput7), 
        .A(n6753), .ZN(n6761) );
  AOI22_X1 U7688 ( .A1(n6756), .A2(keyinput25), .B1(keyinput40), .B2(n6783), 
        .ZN(n6755) );
  OAI221_X1 U7689 ( .B1(n6756), .B2(keyinput25), .C1(n6783), .C2(keyinput40), 
        .A(n6755), .ZN(n6760) );
  XNOR2_X1 U7690 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .B(keyinput36), .ZN(
        n6758) );
  XNOR2_X1 U7691 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .B(keyinput5), .ZN(n6757)
         );
  NAND2_X1 U7692 ( .A1(n6758), .A2(n6757), .ZN(n6759) );
  NOR4_X1 U7693 ( .A1(n6762), .A2(n6761), .A3(n6760), .A4(n6759), .ZN(n6776)
         );
  INV_X1 U7694 ( .A(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n6780) );
  AOI22_X1 U7695 ( .A1(n6780), .A2(keyinput55), .B1(keyinput12), .B2(n6764), 
        .ZN(n6763) );
  OAI221_X1 U7696 ( .B1(n6780), .B2(keyinput55), .C1(n6764), .C2(keyinput12), 
        .A(n6763), .ZN(n6774) );
  AOI22_X1 U7697 ( .A1(n6803), .A2(keyinput10), .B1(n6802), .B2(keyinput49), 
        .ZN(n6765) );
  OAI221_X1 U7698 ( .B1(n6803), .B2(keyinput10), .C1(n6802), .C2(keyinput49), 
        .A(n6765), .ZN(n6773) );
  AOI22_X1 U7699 ( .A1(n6768), .A2(keyinput3), .B1(keyinput6), .B2(n6767), 
        .ZN(n6766) );
  OAI221_X1 U7700 ( .B1(n6768), .B2(keyinput3), .C1(n6767), .C2(keyinput6), 
        .A(n6766), .ZN(n6772) );
  XNOR2_X1 U7701 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .B(keyinput59), .ZN(n6770) );
  XNOR2_X1 U7702 ( .A(keyinput37), .B(DATAI_21_), .ZN(n6769) );
  NAND2_X1 U7703 ( .A1(n6770), .A2(n6769), .ZN(n6771) );
  NOR4_X1 U7704 ( .A1(n6774), .A2(n6773), .A3(n6772), .A4(n6771), .ZN(n6775)
         );
  NAND4_X1 U7705 ( .A1(n6778), .A2(n6777), .A3(n6776), .A4(n6775), .ZN(n6852)
         );
  NOR4_X1 U7706 ( .A1(PHYADDRPOINTER_REG_10__SCAN_IN), .A2(EBX_REG_0__SCAN_IN), 
        .A3(UWORD_REG_13__SCAN_IN), .A4(n4712), .ZN(n6788) );
  INV_X1 U7707 ( .A(DATAI_21_), .ZN(n6779) );
  NOR4_X1 U7708 ( .A1(DATAI_5_), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .A3(n6780), 
        .A4(n6779), .ZN(n6787) );
  NOR4_X1 U7709 ( .A1(STATE2_REG_2__SCAN_IN), .A2(REIP_REG_14__SCAN_IN), .A3(
        n6782), .A4(n6781), .ZN(n6786) );
  AND4_X1 U7710 ( .A1(n6784), .A2(n6783), .A3(INSTQUEUE_REG_8__3__SCAN_IN), 
        .A4(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6785) );
  NAND4_X1 U7711 ( .A1(n6788), .A2(n6787), .A3(n6786), .A4(n6785), .ZN(n6850)
         );
  INV_X1 U7712 ( .A(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n6790) );
  NOR4_X1 U7713 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(UWORD_REG_2__SCAN_IN), 
        .A3(n6790), .A4(n6789), .ZN(n6816) );
  NOR4_X1 U7714 ( .A1(n6794), .A2(n6793), .A3(n6792), .A4(n6791), .ZN(n6815)
         );
  NAND4_X1 U7715 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(ADS_N_REG_SCAN_IN), 
        .A3(n6796), .A4(n6795), .ZN(n6797) );
  NOR4_X1 U7716 ( .A1(EAX_REG_24__SCAN_IN), .A2(DATAO_REG_27__SCAN_IN), .A3(
        n6798), .A4(n6797), .ZN(n6814) );
  NAND4_X1 U7717 ( .A1(EAX_REG_8__SCAN_IN), .A2(DATAI_6_), .A3(
        DATAO_REG_14__SCAN_IN), .A4(n6799), .ZN(n6812) );
  NOR3_X1 U7718 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        DATAO_REG_13__SCAN_IN), .A3(n5448), .ZN(n6805) );
  NOR4_X1 U7719 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), 
        .A3(REIP_REG_22__SCAN_IN), .A4(n6800), .ZN(n6801) );
  AND4_X1 U7720 ( .A1(n6802), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .A3(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A4(n6801), .ZN(n6804) );
  NAND4_X1 U7721 ( .A1(n6805), .A2(ADDRESS_REG_15__SCAN_IN), .A3(n6804), .A4(
        n6803), .ZN(n6811) );
  NAND4_X1 U7722 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(
        INSTQUEUE_REG_10__6__SCAN_IN), .A3(ADDRESS_REG_21__SCAN_IN), .A4(n6836), .ZN(n6810) );
  NOR4_X1 U7723 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(READY_N), .A3(
        DATAWIDTH_REG_1__SCAN_IN), .A4(n6818), .ZN(n6808) );
  NOR4_X1 U7724 ( .A1(EBX_REG_4__SCAN_IN), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .A3(LWORD_REG_13__SCAN_IN), .A4(n6841), .ZN(n6807) );
  AND4_X1 U7725 ( .A1(n6821), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        INSTQUEUE_REG_14__7__SCAN_IN), .A4(LWORD_REG_10__SCAN_IN), .ZN(n6806)
         );
  NAND3_X1 U7726 ( .A1(n6808), .A2(n6807), .A3(n6806), .ZN(n6809) );
  NOR4_X1 U7727 ( .A1(n6812), .A2(n6811), .A3(n6810), .A4(n6809), .ZN(n6813)
         );
  NAND4_X1 U7728 ( .A1(n6816), .A2(n6815), .A3(n6814), .A4(n6813), .ZN(n6849)
         );
  AOI22_X1 U7729 ( .A1(n6819), .A2(keyinput15), .B1(n6818), .B2(keyinput11), 
        .ZN(n6817) );
  OAI221_X1 U7730 ( .B1(n6819), .B2(keyinput15), .C1(n6818), .C2(keyinput11), 
        .A(n6817), .ZN(n6831) );
  INV_X1 U7731 ( .A(LWORD_REG_10__SCAN_IN), .ZN(n6822) );
  INV_X1 U7732 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6821) );
  AOI22_X1 U7733 ( .A1(n6822), .A2(keyinput0), .B1(n6821), .B2(keyinput35), 
        .ZN(n6820) );
  OAI221_X1 U7734 ( .B1(n6822), .B2(keyinput0), .C1(n6821), .C2(keyinput35), 
        .A(n6820), .ZN(n6830) );
  INV_X1 U7735 ( .A(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n6825) );
  AOI22_X1 U7736 ( .A1(n6825), .A2(keyinput38), .B1(keyinput13), .B2(n6824), 
        .ZN(n6823) );
  OAI221_X1 U7737 ( .B1(n6825), .B2(keyinput38), .C1(n6824), .C2(keyinput13), 
        .A(n6823), .ZN(n6829) );
  XNOR2_X1 U7738 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .B(keyinput20), .ZN(
        n6827) );
  XNOR2_X1 U7739 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .B(keyinput21), .ZN(n6826) );
  NAND2_X1 U7740 ( .A1(n6827), .A2(n6826), .ZN(n6828) );
  NOR4_X1 U7741 ( .A1(n6831), .A2(n6830), .A3(n6829), .A4(n6828), .ZN(n6848)
         );
  INV_X1 U7742 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n6833) );
  AOI22_X1 U7743 ( .A1(n6834), .A2(keyinput17), .B1(n6833), .B2(keyinput63), 
        .ZN(n6832) );
  OAI221_X1 U7744 ( .B1(n6834), .B2(keyinput17), .C1(n6833), .C2(keyinput63), 
        .A(n6832), .ZN(n6846) );
  AOI22_X1 U7745 ( .A1(n6836), .A2(keyinput27), .B1(n5080), .B2(keyinput4), 
        .ZN(n6835) );
  OAI221_X1 U7746 ( .B1(n6836), .B2(keyinput27), .C1(n5080), .C2(keyinput4), 
        .A(n6835), .ZN(n6845) );
  AOI22_X1 U7747 ( .A1(n6839), .A2(keyinput41), .B1(keyinput45), .B2(n6838), 
        .ZN(n6837) );
  OAI221_X1 U7748 ( .B1(n6839), .B2(keyinput41), .C1(n6838), .C2(keyinput45), 
        .A(n6837), .ZN(n6844) );
  INV_X1 U7749 ( .A(LWORD_REG_13__SCAN_IN), .ZN(n6842) );
  AOI22_X1 U7750 ( .A1(n6842), .A2(keyinput30), .B1(n6841), .B2(keyinput52), 
        .ZN(n6840) );
  OAI221_X1 U7751 ( .B1(n6842), .B2(keyinput30), .C1(n6841), .C2(keyinput52), 
        .A(n6840), .ZN(n6843) );
  NOR4_X1 U7752 ( .A1(n6846), .A2(n6845), .A3(n6844), .A4(n6843), .ZN(n6847)
         );
  OAI211_X1 U7753 ( .C1(n6850), .C2(n6849), .A(n6848), .B(n6847), .ZN(n6851)
         );
  NOR4_X1 U7754 ( .A1(n6854), .A2(n6853), .A3(n6852), .A4(n6851), .ZN(n6859)
         );
  AOI222_X1 U7755 ( .A1(n6857), .A2(REIP_REG_28__SCAN_IN), .B1(
        REIP_REG_29__SCAN_IN), .B2(n6856), .C1(ADDRESS_REG_27__SCAN_IN), .C2(
        n6855), .ZN(n6858) );
  XNOR2_X1 U7756 ( .A(n6859), .B(n6858), .ZN(U3211) );
  CLKBUF_X1 U3415 ( .A(n3311), .Z(n3312) );
  INV_X1 U3434 ( .A(n3237), .ZN(n3167) );
  INV_X1 U3538 ( .A(n3165), .ZN(n3246) );
  CLKBUF_X1 U3557 ( .A(n3318), .Z(n2956) );
  INV_X2 U3567 ( .A(n3249), .ZN(n3234) );
  CLKBUF_X1 U3576 ( .A(n3237), .Z(n4631) );
  AND2_X1 U3580 ( .A1(n3107), .A2(n4537), .ZN(n3173) );
  CLKBUF_X1 U3699 ( .A(n3582), .Z(n3583) );
  CLKBUF_X2 U3840 ( .A(n3210), .Z(n4724) );
  CLKBUF_X1 U4613 ( .A(n6448), .Z(n6439) );
endmodule

