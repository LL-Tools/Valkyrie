

module b20_C_gen_AntiSAT_k_256_2 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, 
        keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, 
        keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, 
        keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, 
        keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, 
        keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, 
        keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, 
        keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, 
        keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104, 
        keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108, 
        keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112, 
        keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116, 
        keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120, 
        keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124, 
        keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, 
        keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, 
        keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, 
        keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, 
        keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, 
        keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, 
        keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, 
        keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541;

  CLKBUF_X2 U5016 ( .A(n6546), .Z(n7534) );
  CLKBUF_X1 U5017 ( .A(n6544), .Z(n7504) );
  INV_X2 U5018 ( .A(n7768), .ZN(n7775) );
  NAND2_X1 U5019 ( .A1(n8295), .A2(n7998), .ZN(n4892) );
  INV_X2 U5020 ( .A(n6625), .ZN(n5711) );
  CLKBUF_X1 U5021 ( .A(n5190), .Z(n5861) );
  OR2_X1 U5022 ( .A1(n5214), .A2(n8803), .ZN(n5178) );
  NAND2_X1 U5023 ( .A1(n5719), .A2(n5720), .ZN(n5190) );
  CLKBUF_X1 U5024 ( .A(n8760), .Z(n4510) );
  CLKBUF_X1 U5025 ( .A(n6933), .Z(n4511) );
  INV_X1 U5026 ( .A(n6541), .ZN(n7307) );
  INV_X1 U5027 ( .A(n7998), .ZN(n8292) );
  INV_X1 U5028 ( .A(n8295), .ZN(n7959) );
  INV_X1 U5029 ( .A(n9386), .ZN(n9626) );
  INV_X1 U5030 ( .A(n4602), .ZN(n7989) );
  INV_X1 U5031 ( .A(n7534), .ZN(n7526) );
  AND3_X1 U5032 ( .A1(n6731), .A2(n6730), .A3(n6729), .ZN(n6844) );
  AOI21_X1 U5033 ( .B1(n8452), .B2(n6809), .A(n8451), .ZN(n8457) );
  XNOR2_X1 U5034 ( .A(n4835), .B(n4834), .ZN(n8477) );
  INV_X1 U5035 ( .A(n8802), .ZN(n8728) );
  INV_X1 U5036 ( .A(n5222), .ZN(n7579) );
  AND3_X2 U5037 ( .A1(n6447), .A2(n6446), .A3(n6445), .ZN(n8077) );
  AOI211_X1 U5038 ( .C1(n8572), .C2(n9877), .A(n8571), .B(n8570), .ZN(n8573)
         );
  INV_X1 U5039 ( .A(n9598), .ZN(n9585) );
  AND2_X2 U5040 ( .A1(n6423), .A2(n8788), .ZN(n8802) );
  CLKBUF_X3 U5041 ( .A(n5153), .Z(n6178) );
  OAI211_X2 U5042 ( .C1(n7662), .C2(n7661), .A(n7660), .B(n7659), .ZN(n7665)
         );
  NAND4_X2 U5043 ( .A1(n6575), .A2(n6574), .A3(n6573), .A4(n6572), .ZN(n9172)
         );
  OAI22_X2 U5044 ( .A1(n6783), .A2(n5053), .B1(n6789), .B2(n10044), .ZN(n6968)
         );
  AOI21_X2 U5045 ( .B1(n6999), .B2(n5732), .A(n4538), .ZN(n6783) );
  CLKBUF_X3 U5046 ( .A(n6676), .Z(n9175) );
  NAND4_X1 U5047 ( .A1(n6453), .A2(n6452), .A3(n6451), .A4(n6450), .ZN(n6676)
         );
  NAND4_X2 U5048 ( .A1(n6556), .A2(n6555), .A3(n6554), .A4(n6553), .ZN(n9173)
         );
  NAND2_X1 U5049 ( .A1(n5967), .A2(n5966), .ZN(n4512) );
  NAND4_X4 U5050 ( .A1(n6405), .A2(n6404), .A3(n6403), .A4(n6402), .ZN(n9177)
         );
  XNOR2_X2 U5051 ( .A(n5949), .B(n5948), .ZN(n5967) );
  NAND2_X2 U5052 ( .A1(n5155), .A2(n5154), .ZN(n9860) );
  XNOR2_X2 U5053 ( .A(n5781), .B(n5780), .ZN(n5791) );
  NAND2_X2 U5054 ( .A1(n5779), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5781) );
  OAI21_X2 U5056 ( .B1(n6981), .B2(n5380), .A(n7678), .ZN(n7183) );
  BUF_X4 U5057 ( .A(n7978), .Z(n4513) );
  NOR2_X2 U5058 ( .A1(n5950), .A2(n5947), .ZN(n5949) );
  NAND2_X2 U5059 ( .A1(n6507), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8452) );
  NOR2_X2 U5060 ( .A1(n6241), .A2(n6337), .ZN(n6342) );
  XNOR2_X2 U5061 ( .A(n8535), .B(n8536), .ZN(n8504) );
  NOR2_X2 U5062 ( .A1(n4544), .A2(n8503), .ZN(n8535) );
  AOI21_X1 U5063 ( .B1(n4807), .B2(n7617), .A(n4576), .ZN(n4779) );
  NAND2_X1 U5064 ( .A1(n9503), .A2(n4760), .ZN(n9474) );
  INV_X1 U5065 ( .A(n8650), .ZN(n8826) );
  NAND2_X1 U5066 ( .A1(n9575), .A2(n8239), .ZN(n9578) );
  NAND2_X1 U5067 ( .A1(n5735), .A2(n5734), .ZN(n6982) );
  OR2_X1 U5068 ( .A1(n6504), .A2(n4670), .ZN(n4669) );
  XNOR2_X2 U5069 ( .A(n6722), .B(n9174), .ZN(n6684) );
  NOR2_X1 U5070 ( .A1(n9178), .A2(n6917), .ZN(n6672) );
  INV_X1 U5071 ( .A(n5868), .ZN(n8790) );
  NAND2_X2 U5072 ( .A1(n5793), .A2(n6083), .ZN(n6073) );
  CLKBUF_X2 U5073 ( .A(n6551), .Z(n7988) );
  CLKBUF_X2 U5075 ( .A(n5213), .Z(n5484) );
  XNOR2_X1 U5077 ( .A(n5170), .B(n8977), .ZN(n7554) );
  INV_X1 U5078 ( .A(n5928), .ZN(n7550) );
  AND2_X1 U5079 ( .A1(n9872), .A2(n9873), .ZN(n9870) );
  CLKBUF_X2 U5080 ( .A(n5158), .Z(n7468) );
  AOI21_X1 U5081 ( .B1(n4781), .B2(n4780), .A(n4778), .ZN(n7785) );
  OAI21_X1 U5082 ( .B1(n5039), .B2(n10070), .A(n5038), .ZN(n5836) );
  INV_X1 U5083 ( .A(n4779), .ZN(n4778) );
  NOR2_X1 U5084 ( .A1(n7779), .A2(n5824), .ZN(n4780) );
  NOR2_X1 U5085 ( .A1(n7765), .A2(n7764), .ZN(n7776) );
  OAI21_X1 U5086 ( .B1(n5761), .B2(n4535), .A(n5045), .ZN(n8589) );
  NAND2_X1 U5087 ( .A1(n5044), .A2(n5755), .ZN(n8648) );
  AOI21_X1 U5088 ( .B1(n9063), .B2(n4859), .A(n4856), .ZN(n4855) );
  OAI21_X1 U5089 ( .B1(n9453), .B2(n4750), .A(n4748), .ZN(n9299) );
  OAI21_X1 U5090 ( .B1(n9959), .B2(n4906), .A(n4905), .ZN(n8555) );
  NAND2_X1 U5091 ( .A1(n9116), .A2(n9117), .ZN(n9115) );
  NAND2_X1 U5092 ( .A1(n4857), .A2(n7931), .ZN(n4856) );
  XNOR2_X1 U5093 ( .A(n8542), .B(n8541), .ZN(n9959) );
  INV_X1 U5094 ( .A(n4749), .ZN(n4748) );
  OAI21_X1 U5095 ( .B1(n4516), .B2(n4750), .A(n9415), .ZN(n4749) );
  NOR2_X1 U5096 ( .A1(n9941), .A2(n8540), .ZN(n8542) );
  NAND2_X1 U5097 ( .A1(n8424), .A2(n8026), .ZN(n8353) );
  OAI21_X1 U5098 ( .B1(n9578), .B2(n4757), .A(n4755), .ZN(n8243) );
  NAND2_X1 U5099 ( .A1(n4673), .A2(n4545), .ZN(n4672) );
  NOR2_X1 U5100 ( .A1(n9913), .A2(n8474), .ZN(n9932) );
  NAND2_X1 U5101 ( .A1(n4743), .A2(n8127), .ZN(n8237) );
  NOR2_X1 U5102 ( .A1(n4607), .A2(n10041), .ZN(n4606) );
  AND2_X1 U5103 ( .A1(n5013), .A2(n8737), .ZN(n5012) );
  NOR2_X1 U5104 ( .A1(n9892), .A2(n4596), .ZN(n8473) );
  NAND2_X1 U5105 ( .A1(n6847), .A2(n4887), .ZN(n7106) );
  INV_X1 U5106 ( .A(n9811), .ZN(n7318) );
  NOR2_X1 U5107 ( .A1(n4669), .A2(n6816), .ZN(n4668) );
  OAI211_X1 U5108 ( .C1(n5861), .C2(n6164), .A(n5233), .B(n5232), .ZN(n9997)
         );
  INV_X4 U5109 ( .A(n8048), .ZN(n8051) );
  NOR2_X1 U5110 ( .A1(n6909), .A2(n9327), .ZN(n9538) );
  AND4_X1 U5111 ( .A1(n5242), .A2(n5241), .A3(n5240), .A4(n5239), .ZN(n10001)
         );
  NAND2_X1 U5112 ( .A1(n5246), .A2(n5245), .ZN(n5252) );
  INV_X1 U5113 ( .A(n5721), .ZN(n8796) );
  AND4_X1 U5114 ( .A1(n5187), .A2(n5186), .A3(n5185), .A4(n5184), .ZN(n5721)
         );
  NAND2_X2 U5115 ( .A1(n5958), .A2(n5957), .ZN(n8295) );
  NAND4_X2 U5116 ( .A1(n6492), .A2(n6491), .A3(n6490), .A4(n6489), .ZN(n9174)
         );
  NAND4_X2 U5117 ( .A1(n5209), .A2(n5208), .A3(n5207), .A4(n5206), .ZN(n9998)
         );
  NAND2_X1 U5118 ( .A1(n5139), .A2(n7782), .ZN(n5867) );
  NAND4_X1 U5119 ( .A1(n5935), .A2(n5934), .A3(n5933), .A4(n5932), .ZN(n9178)
         );
  NAND2_X1 U5120 ( .A1(n5230), .A2(n5229), .ZN(n5246) );
  OAI211_X1 U5121 ( .C1(n7577), .C2(n6070), .A(n5113), .B(n5166), .ZN(n5868)
         );
  XNOR2_X1 U5122 ( .A(n5126), .B(n5128), .ZN(n5139) );
  AND2_X2 U5123 ( .A1(n7551), .A2(n5928), .ZN(n7978) );
  AND2_X4 U5124 ( .A1(n5958), .A2(n5940), .ZN(n6541) );
  NAND2_X1 U5125 ( .A1(n6181), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6280) );
  AOI21_X1 U5126 ( .B1(n6275), .B2(n4530), .A(n6274), .ZN(n6277) );
  BUF_X2 U5127 ( .A(n5927), .Z(n7551) );
  OR3_X2 U5128 ( .A1(n7558), .A2(n9794), .A3(n7452), .ZN(n5958) );
  NAND2_X2 U5129 ( .A1(n5190), .A2(n6433), .ZN(n7577) );
  XNOR2_X1 U5130 ( .A(n5784), .B(n5783), .ZN(n5794) );
  XNOR2_X1 U5131 ( .A(n5849), .B(n5848), .ZN(n7558) );
  INV_X1 U5132 ( .A(n5175), .ZN(n8287) );
  NAND2_X1 U5133 ( .A1(n5782), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5784) );
  XNOR2_X1 U5134 ( .A(n5923), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U5135 ( .A1(n8979), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5170) );
  XNOR2_X1 U5136 ( .A(n5146), .B(n5145), .ZN(n5720) );
  XNOR2_X1 U5137 ( .A(n5172), .B(n5144), .ZN(n5719) );
  NOR2_X1 U5138 ( .A1(n5922), .A2(n4536), .ZN(n5925) );
  NAND2_X1 U5139 ( .A1(n5788), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5146) );
  INV_X2 U5140 ( .A(n9790), .ZN(n7300) );
  OR2_X1 U5141 ( .A1(n9851), .A2(n6155), .ZN(n9853) );
  INV_X1 U5142 ( .A(n5778), .ZN(n5143) );
  AND3_X2 U5143 ( .A1(n5844), .A2(n4762), .A3(n5996), .ZN(n5846) );
  NOR2_X1 U5144 ( .A1(n4565), .A2(n5090), .ZN(n5089) );
  NAND2_X1 U5145 ( .A1(n5150), .A2(n5151), .ZN(n5158) );
  NAND2_X1 U5146 ( .A1(n5149), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5150) );
  OR2_X1 U5147 ( .A1(n6178), .A2(n4909), .ZN(n4908) );
  NAND2_X1 U5148 ( .A1(n5153), .A2(n5117), .ZN(n5257) );
  OAI21_X1 U5149 ( .B1(P1_RD_REG_SCAN_IN), .B2(P1_ADDR_REG_19__SCAN_IN), .A(
        n5147), .ZN(n5151) );
  AND2_X1 U5150 ( .A1(n5838), .A2(n6024), .ZN(n5839) );
  AND3_X1 U5151 ( .A1(n5991), .A2(n5972), .A3(n5056), .ZN(n5996) );
  NOR2_X2 U5152 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5972) );
  NOR2_X1 U5153 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5118) );
  INV_X1 U5154 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5258) );
  NOR2_X1 U5155 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5119) );
  INV_X1 U5156 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5130) );
  INV_X1 U5157 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5128) );
  NOR2_X1 U5158 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5117) );
  INV_X1 U5159 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5479) );
  INV_X1 U5160 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5147) );
  INV_X1 U5161 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5438) );
  INV_X4 U5162 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U5163 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5441) );
  INV_X4 U5164 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5165 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6056) );
  NOR2_X1 U5166 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5838) );
  INV_X1 U5167 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5069) );
  INV_X1 U5168 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U5169 ( .A1(n5177), .A2(n5175), .ZN(n5213) );
  NOR2_X1 U5170 ( .A1(n6810), .A2(n5352), .ZN(n6878) );
  AOI21_X2 U5171 ( .B1(n8340), .B2(n8339), .A(n8037), .ZN(n8399) );
  INV_X4 U5172 ( .A(n5211), .ZN(n5182) );
  NOR2_X2 U5173 ( .A1(n4709), .A2(n7449), .ZN(n7384) );
  NOR2_X2 U5174 ( .A1(n8353), .A2(n8354), .ZN(n8364) );
  OAI21_X2 U5175 ( .B1(n7005), .B2(n6737), .A(n8079), .ZN(n7046) );
  OAI21_X2 U5176 ( .B1(n4611), .B2(n4610), .A(n4608), .ZN(n7005) );
  OAI21_X2 U5177 ( .B1(n8364), .B2(n8363), .A(n8362), .ZN(n8361) );
  NAND2_X2 U5178 ( .A1(n8647), .A2(n7746), .ZN(n8641) );
  AOI21_X2 U5179 ( .B1(n8657), .B2(n7742), .A(n7744), .ZN(n8647) );
  INV_X1 U5180 ( .A(n7504), .ZN(n4514) );
  NAND2_X1 U5181 ( .A1(n4512), .A2(n6433), .ZN(n6544) );
  NOR2_X2 U5182 ( .A1(n9431), .A2(n9445), .ZN(n9434) );
  OR2_X1 U5183 ( .A1(n7206), .A2(n6664), .ZN(n6706) );
  XNOR2_X1 U5184 ( .A(n9177), .B(n7206), .ZN(n6673) );
  OAI211_X4 U5185 ( .C1(n6544), .C2(n6434), .A(n5055), .B(n5054), .ZN(n7206)
         );
  AND2_X1 U5186 ( .A1(n5089), .A2(n10342), .ZN(n5088) );
  OAI21_X1 U5187 ( .B1(n5549), .B2(n5548), .A(n5547), .ZN(n5562) );
  AOI21_X1 U5188 ( .B1(n4787), .B2(n7768), .A(n4786), .ZN(n4785) );
  NAND2_X1 U5189 ( .A1(n8042), .A2(n8838), .ZN(n4942) );
  INV_X1 U5190 ( .A(n7618), .ZN(n7626) );
  OAI21_X1 U5191 ( .B1(n5533), .B2(n5532), .A(n5531), .ZN(n5549) );
  AND2_X1 U5192 ( .A1(n5839), .A2(n5067), .ZN(n4762) );
  AND2_X1 U5193 ( .A1(n5069), .A2(n5845), .ZN(n5067) );
  INV_X1 U5194 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U5195 ( .A1(n7644), .A2(n4551), .ZN(n4783) );
  AOI21_X1 U5196 ( .B1(n4619), .B2(n8142), .A(n4618), .ZN(n4617) );
  OAI21_X1 U5197 ( .B1(n7753), .B2(n7775), .A(n8622), .ZN(n4771) );
  NAND2_X1 U5198 ( .A1(n8175), .A2(n4701), .ZN(n8069) );
  NAND2_X1 U5199 ( .A1(n4703), .A2(n4702), .ZN(n4701) );
  NAND2_X1 U5200 ( .A1(n4704), .A2(n9303), .ZN(n4703) );
  AND2_X1 U5201 ( .A1(n9940), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8503) );
  AOI21_X1 U5202 ( .B1(n5017), .B2(n5015), .A(n4566), .ZN(n5014) );
  INV_X1 U5203 ( .A(n5022), .ZN(n5015) );
  INV_X1 U5204 ( .A(n7690), .ZN(n4806) );
  NAND2_X1 U5205 ( .A1(n5167), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5172) );
  NAND2_X1 U5206 ( .A1(n5143), .A2(n5049), .ZN(n5788) );
  AND2_X1 U5207 ( .A1(n5142), .A2(n5050), .ZN(n5049) );
  INV_X1 U5208 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5050) );
  MUX2_X1 U5209 ( .A(n8277), .B(n8189), .S(n9265), .Z(n8190) );
  NOR2_X1 U5210 ( .A1(n9376), .A2(n9355), .ZN(n4718) );
  AND2_X1 U5211 ( .A1(n5081), .A2(n9278), .ZN(n5080) );
  OR2_X1 U5212 ( .A1(n9681), .A2(n9485), .ZN(n9278) );
  NAND2_X1 U5213 ( .A1(n5085), .A2(n5083), .ZN(n5081) );
  INV_X1 U5214 ( .A(n5083), .ZN(n5082) );
  AND2_X1 U5215 ( .A1(n9552), .A2(n8240), .ZN(n4759) );
  OR2_X1 U5216 ( .A1(n7422), .A2(n9167), .ZN(n7337) );
  AND2_X1 U5217 ( .A1(n5636), .A2(n5621), .ZN(n5634) );
  NAND2_X1 U5218 ( .A1(n5856), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5953) );
  OAI21_X1 U5219 ( .B1(n5473), .B2(SI_15_), .A(n5475), .ZN(n5491) );
  AND2_X1 U5220 ( .A1(n4997), .A2(n4996), .ZN(n5473) );
  INV_X1 U5221 ( .A(n4998), .ZN(n4996) );
  AND2_X1 U5222 ( .A1(n5365), .A2(n4543), .ZN(n4699) );
  INV_X1 U5223 ( .A(n7616), .ZN(n7617) );
  NAND2_X1 U5224 ( .A1(n4667), .A2(n4666), .ZN(n4665) );
  INV_X1 U5225 ( .A(n6880), .ZN(n4666) );
  AOI21_X1 U5226 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n9940), .A(n9930), .ZN(
        n8511) );
  AND2_X1 U5227 ( .A1(n7573), .A2(n5717), .ZN(n7613) );
  INV_X1 U5228 ( .A(n5008), .ZN(n5007) );
  OAI21_X1 U5229 ( .B1(n8648), .B2(n5756), .A(n5757), .ZN(n8634) );
  NAND2_X1 U5230 ( .A1(n8736), .A2(n7625), .ZN(n4810) );
  INV_X1 U5231 ( .A(n5861), .ZN(n5537) );
  INV_X1 U5232 ( .A(n7577), .ZN(n5538) );
  NAND2_X1 U5233 ( .A1(n5025), .A2(n5024), .ZN(n8772) );
  AOI21_X1 U5234 ( .B1(n5027), .B2(n5029), .A(n4564), .ZN(n5024) );
  OR2_X1 U5235 ( .A1(n5909), .A2(n7768), .ZN(n10027) );
  AND2_X1 U5236 ( .A1(n7296), .A2(n7618), .ZN(n10060) );
  NOR2_X1 U5237 ( .A1(n8105), .A2(n8252), .ZN(n8273) );
  INV_X1 U5238 ( .A(n4513), .ZN(n7992) );
  INV_X1 U5239 ( .A(n7798), .ZN(n7907) );
  NAND2_X1 U5240 ( .A1(n8068), .A2(n9607), .ZN(n9307) );
  NAND2_X1 U5241 ( .A1(n9284), .A2(n9283), .ZN(n9397) );
  NOR2_X1 U5242 ( .A1(n4588), .A2(n5058), .ZN(n5057) );
  OR2_X1 U5243 ( .A1(n9676), .A2(n9437), .ZN(n9296) );
  NAND2_X1 U5244 ( .A1(n9519), .A2(n8245), .ZN(n9503) );
  AND2_X1 U5245 ( .A1(n7520), .A2(n7519), .ZN(n9495) );
  NAND2_X1 U5247 ( .A1(n6675), .A2(n6674), .ZN(n6700) );
  NAND2_X1 U5248 ( .A1(n6680), .A2(n6679), .ZN(n6703) );
  NAND2_X1 U5249 ( .A1(n5929), .A2(n5928), .ZN(n6551) );
  INV_X1 U5250 ( .A(n7504), .ZN(n7533) );
  NAND2_X1 U5251 ( .A1(n7298), .A2(n8267), .ZN(n6912) );
  XNOR2_X1 U5252 ( .A(n7453), .B(SI_29_), .ZN(n7549) );
  INV_X1 U5253 ( .A(n4977), .ZN(n5576) );
  AOI21_X1 U5254 ( .B1(n5562), .B2(n4978), .A(n4979), .ZN(n4977) );
  NAND2_X1 U5255 ( .A1(n5846), .A2(n10261), .ZN(n5937) );
  NOR2_X1 U5256 ( .A1(n4885), .A2(n6115), .ZN(n4884) );
  NAND2_X1 U5257 ( .A1(n4689), .A2(n4694), .ZN(n5436) );
  INV_X1 U5258 ( .A(n4695), .ZN(n4694) );
  NAND2_X1 U5259 ( .A1(n5361), .A2(n4690), .ZN(n4689) );
  OAI21_X1 U5260 ( .B1(n4697), .B2(n4696), .A(n5421), .ZN(n4695) );
  NAND2_X1 U5261 ( .A1(n4692), .A2(n4699), .ZN(n5382) );
  OAI21_X1 U5262 ( .B1(n4938), .B2(n4936), .A(n4592), .ZN(n4934) );
  NOR2_X1 U5263 ( .A1(n4937), .A2(n4936), .ZN(n4935) );
  AND2_X1 U5264 ( .A1(n4872), .A2(n4871), .ZN(n8307) );
  NOR2_X1 U5265 ( .A1(n8011), .A2(n8009), .ZN(n4871) );
  NAND2_X1 U5266 ( .A1(n4783), .A2(n4782), .ZN(n7639) );
  NOR2_X1 U5267 ( .A1(n4634), .A2(n8194), .ZN(n4633) );
  INV_X1 U5268 ( .A(n8207), .ZN(n4634) );
  AOI21_X1 U5269 ( .B1(n4621), .B2(n4620), .A(n8238), .ZN(n4619) );
  INV_X1 U5270 ( .A(n8143), .ZN(n4620) );
  AOI21_X1 U5271 ( .B1(n4614), .B2(n4616), .A(n4575), .ZN(n4613) );
  AND2_X1 U5272 ( .A1(n8166), .A2(n4625), .ZN(n4624) );
  NOR2_X1 U5273 ( .A1(n9382), .A2(n8161), .ZN(n4625) );
  OR3_X1 U5274 ( .A1(n8160), .A2(n4750), .A3(n8194), .ZN(n8167) );
  NOR2_X1 U5275 ( .A1(n7752), .A2(n7768), .ZN(n4770) );
  INV_X1 U5276 ( .A(n5690), .ZN(n4985) );
  INV_X1 U5277 ( .A(n4984), .ZN(n4983) );
  OAI21_X1 U5278 ( .B1(n5688), .B2(n4985), .A(n5703), .ZN(n4984) );
  NOR2_X1 U5279 ( .A1(n4979), .A2(n4976), .ZN(n4975) );
  INV_X1 U5280 ( .A(n5547), .ZN(n4976) );
  NAND2_X1 U5281 ( .A1(n4765), .A2(n4549), .ZN(n7765) );
  NAND2_X1 U5282 ( .A1(n4766), .A2(n4562), .ZN(n4765) );
  NAND2_X1 U5283 ( .A1(n7622), .A2(n4764), .ZN(n4763) );
  NOR2_X1 U5284 ( .A1(n5739), .A2(n5018), .ZN(n5017) );
  INV_X1 U5285 ( .A(n5020), .ZN(n5018) );
  AOI21_X1 U5286 ( .B1(n5548), .B2(n4975), .A(n4974), .ZN(n4973) );
  INV_X1 U5287 ( .A(n4978), .ZN(n4974) );
  INV_X1 U5288 ( .A(n5577), .ZN(n5578) );
  AOI21_X1 U5289 ( .B1(n4929), .B2(n4932), .A(n8388), .ZN(n4927) );
  INV_X1 U5290 ( .A(n4929), .ZN(n4928) );
  NOR2_X1 U5291 ( .A1(n4557), .A2(n7618), .ZN(n4808) );
  AND2_X1 U5292 ( .A1(n8581), .A2(n8591), .ZN(n7773) );
  OR2_X1 U5293 ( .A1(n9870), .A2(n4578), .ZN(n4663) );
  AND2_X1 U5294 ( .A1(n4663), .A2(n6164), .ZN(n6244) );
  NOR2_X1 U5295 ( .A1(n7134), .A2(n4605), .ZN(n8469) );
  NOR2_X1 U5296 ( .A1(n6895), .A2(n6896), .ZN(n4605) );
  AND3_X1 U5297 ( .A1(n4897), .A2(n4895), .A3(n4899), .ZN(n8501) );
  INV_X1 U5298 ( .A(n5709), .ZN(n7796) );
  NOR2_X1 U5299 ( .A1(n4815), .A2(n4521), .ZN(n4813) );
  INV_X1 U5300 ( .A(n7730), .ZN(n4815) );
  NAND2_X1 U5301 ( .A1(n5746), .A2(n4532), .ZN(n5037) );
  OAI211_X1 U5302 ( .C1(n5861), .C2(n9880), .A(n5204), .B(n5203), .ZN(n5873)
         );
  OR2_X1 U5303 ( .A1(n7577), .A2(n5195), .ZN(n5203) );
  INV_X1 U5304 ( .A(n5762), .ZN(n5047) );
  NOR2_X1 U5305 ( .A1(n8598), .A2(n4791), .ZN(n4790) );
  INV_X1 U5306 ( .A(n4793), .ZN(n4791) );
  INV_X1 U5307 ( .A(n5017), .ZN(n5016) );
  OAI21_X1 U5308 ( .B1(n7684), .B2(n4806), .A(n5434), .ZN(n4805) );
  OR2_X1 U5309 ( .A1(n8964), .A2(n8023), .ZN(n7698) );
  AND2_X1 U5310 ( .A1(n7589), .A2(n7588), .ZN(n7691) );
  OAI21_X1 U5311 ( .B1(n5912), .B2(n5892), .A(n6073), .ZN(n5828) );
  NAND2_X1 U5312 ( .A1(n4950), .A2(n4949), .ZN(n5125) );
  AND2_X1 U5313 ( .A1(n5479), .A2(n5130), .ZN(n4949) );
  INV_X1 U5314 ( .A(n5478), .ZN(n4950) );
  NOR2_X2 U5315 ( .A1(n4951), .A2(n5257), .ZN(n5383) );
  NAND2_X1 U5316 ( .A1(n4881), .A2(n4879), .ZN(n4878) );
  INV_X1 U5317 ( .A(n4883), .ZN(n4879) );
  NAND2_X1 U5318 ( .A1(n7417), .A2(n7416), .ZN(n7434) );
  NOR2_X1 U5319 ( .A1(n7890), .A2(n4868), .ZN(n4867) );
  NAND2_X1 U5320 ( .A1(n4865), .A2(n7889), .ZN(n4864) );
  OR2_X1 U5321 ( .A1(n7890), .A2(n4866), .ZN(n4865) );
  INV_X1 U5322 ( .A(n4685), .ZN(n8256) );
  OAI21_X1 U5323 ( .B1(n8254), .B2(n8253), .A(n4686), .ZN(n4685) );
  NOR2_X1 U5324 ( .A1(n8255), .A2(n4556), .ZN(n4686) );
  OR2_X1 U5325 ( .A1(n7985), .A2(n9146), .ZN(n7987) );
  OR2_X1 U5326 ( .A1(n9376), .A2(n9626), .ZN(n8198) );
  AND2_X1 U5327 ( .A1(n4520), .A2(n9751), .ZN(n4716) );
  AND2_X1 U5328 ( .A1(n6477), .A2(n9343), .ZN(n6469) );
  NAND2_X1 U5329 ( .A1(n5671), .A2(n5670), .ZN(n5689) );
  AOI21_X1 U5330 ( .B1(n4969), .B2(n4971), .A(n4968), .ZN(n4967) );
  INV_X1 U5331 ( .A(n5636), .ZN(n4968) );
  NAND2_X1 U5332 ( .A1(n4626), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5936) );
  NAND2_X1 U5333 ( .A1(n4700), .A2(n5513), .ZN(n5533) );
  NAND2_X1 U5334 ( .A1(n4995), .A2(n4587), .ZN(n4700) );
  NAND2_X1 U5335 ( .A1(n4955), .A2(n4956), .ZN(n5361) );
  NAND2_X1 U5336 ( .A1(n5303), .A2(n4515), .ZN(n4955) );
  AOI21_X1 U5337 ( .B1(n4515), .B2(n4957), .A(n4571), .ZN(n4956) );
  AOI21_X1 U5338 ( .B1(n5308), .B2(n4963), .A(n4962), .ZN(n4961) );
  INV_X1 U5339 ( .A(n5323), .ZN(n4962) );
  INV_X1 U5340 ( .A(n5302), .ZN(n4963) );
  NAND2_X1 U5341 ( .A1(n8413), .A2(n8414), .ZN(n4918) );
  INV_X1 U5342 ( .A(n5872), .ZN(n4915) );
  AND2_X1 U5343 ( .A1(n4931), .A2(n4930), .ZN(n4929) );
  INV_X1 U5344 ( .A(n7289), .ZN(n4930) );
  NOR2_X1 U5345 ( .A1(n4941), .A2(n4940), .ZN(n4939) );
  INV_X1 U5346 ( .A(n8041), .ZN(n4940) );
  INV_X1 U5347 ( .A(n4942), .ZN(n4941) );
  NAND2_X1 U5348 ( .A1(n4593), .A2(n4942), .ZN(n4938) );
  NOR2_X1 U5349 ( .A1(n8380), .A2(n4948), .ZN(n4947) );
  INV_X1 U5350 ( .A(n8033), .ZN(n4948) );
  INV_X1 U5351 ( .A(n6307), .ZN(n4921) );
  INV_X1 U5352 ( .A(n5885), .ZN(n4923) );
  OR2_X1 U5353 ( .A1(n7770), .A2(n7769), .ZN(n7771) );
  NOR2_X1 U5354 ( .A1(n9883), .A2(n9884), .ZN(n9882) );
  AOI21_X1 U5355 ( .B1(n6350), .B2(n4529), .A(n6349), .ZN(n6504) );
  NAND2_X1 U5356 ( .A1(n6246), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6350) );
  NAND2_X1 U5357 ( .A1(n7140), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4664) );
  OR2_X1 U5358 ( .A1(n7132), .A2(n4898), .ZN(n4897) );
  OR2_X1 U5359 ( .A1(n9891), .A2(n5387), .ZN(n4898) );
  NAND2_X1 U5360 ( .A1(n8498), .A2(n4896), .ZN(n4895) );
  INV_X1 U5361 ( .A(n9891), .ZN(n4896) );
  OAI21_X1 U5362 ( .B1(n7135), .B2(n4847), .A(n4846), .ZN(n9892) );
  NAND2_X1 U5363 ( .A1(n4850), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4847) );
  NAND2_X1 U5364 ( .A1(n8471), .A2(n4850), .ZN(n4846) );
  INV_X1 U5365 ( .A(n9893), .ZN(n4850) );
  OR2_X1 U5366 ( .A1(n7135), .A2(n7188), .ZN(n4849) );
  XNOR2_X1 U5367 ( .A(n8501), .B(n8500), .ZN(n9907) );
  INV_X1 U5368 ( .A(n9924), .ZN(n4671) );
  OAI21_X1 U5369 ( .B1(n8477), .B2(n4832), .A(n4831), .ZN(n9943) );
  NAND2_X1 U5370 ( .A1(n4833), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4832) );
  NAND2_X1 U5371 ( .A1(n8513), .A2(n4833), .ZN(n4831) );
  XNOR2_X1 U5372 ( .A(n5766), .B(n7613), .ZN(n5042) );
  NAND2_X1 U5373 ( .A1(n4797), .A2(n7757), .ZN(n4796) );
  INV_X1 U5374 ( .A(n8600), .ZN(n8598) );
  AND2_X1 U5375 ( .A1(n5759), .A2(n4800), .ZN(n8622) );
  INV_X1 U5376 ( .A(n5484), .ZN(n5710) );
  NAND2_X1 U5377 ( .A1(n5624), .A2(n10479), .ZN(n5644) );
  INV_X1 U5378 ( .A(n5625), .ZN(n5624) );
  OR2_X1 U5379 ( .A1(n8863), .A2(n8869), .ZN(n7723) );
  AND2_X1 U5380 ( .A1(n5749), .A2(n8668), .ZN(n8681) );
  AND2_X1 U5381 ( .A1(n7167), .A2(n5736), .ZN(n5032) );
  NAND2_X1 U5382 ( .A1(n5031), .A2(n7167), .ZN(n5030) );
  INV_X1 U5383 ( .A(n5033), .ZN(n5031) );
  AOI21_X1 U5384 ( .B1(n4537), .B2(n5736), .A(n5034), .ZN(n5033) );
  INV_X1 U5385 ( .A(n7166), .ZN(n5034) );
  NAND2_X1 U5386 ( .A1(n5733), .A2(n5116), .ZN(n5735) );
  AND2_X1 U5387 ( .A1(n7659), .A2(n7645), .ZN(n7642) );
  NAND2_X1 U5388 ( .A1(n6167), .A2(n6083), .ZN(n5912) );
  NAND2_X1 U5389 ( .A1(n7576), .A2(n7575), .ZN(n7783) );
  INV_X1 U5390 ( .A(n4799), .ZN(n4798) );
  OAI21_X1 U5391 ( .B1(n7586), .B2(n5633), .A(n4800), .ZN(n4799) );
  AOI21_X1 U5392 ( .B1(n4798), .B2(n7586), .A(n7754), .ZN(n4797) );
  INV_X1 U5393 ( .A(n8613), .ZN(n8636) );
  NAND2_X1 U5394 ( .A1(n8658), .A2(n8659), .ZN(n5044) );
  NOR2_X1 U5395 ( .A1(n8725), .A2(n7713), .ZN(n4809) );
  OAI21_X1 U5396 ( .B1(n5737), .B2(n5016), .A(n5014), .ZN(n8738) );
  NOR2_X1 U5397 ( .A1(n5738), .A2(n5023), .ZN(n5022) );
  INV_X1 U5398 ( .A(n7588), .ZN(n5023) );
  NAND2_X1 U5399 ( .A1(n5021), .A2(n8023), .ZN(n5020) );
  AND2_X1 U5400 ( .A1(n7703), .A2(n7715), .ZN(n8748) );
  INV_X1 U5401 ( .A(n7691), .ZN(n8773) );
  NAND2_X1 U5402 ( .A1(n7153), .A2(n7684), .ZN(n7157) );
  NAND2_X1 U5403 ( .A1(n5909), .A2(n7775), .ZN(n10025) );
  INV_X1 U5404 ( .A(n10027), .ZN(n10043) );
  INV_X1 U5405 ( .A(n10025), .ZN(n10042) );
  AND2_X1 U5406 ( .A1(n5142), .A2(n5052), .ZN(n5051) );
  NOR2_X1 U5407 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n5052) );
  AND2_X1 U5408 ( .A1(n5789), .A2(n5788), .ZN(n5798) );
  INV_X1 U5409 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5780) );
  INV_X1 U5410 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5141) );
  AND2_X1 U5411 ( .A1(n9007), .A2(n4882), .ZN(n4881) );
  NAND2_X1 U5412 ( .A1(n7957), .A2(n9129), .ZN(n4882) );
  OAI22_X1 U5413 ( .A1(n9035), .A2(n9036), .B1(n7943), .B2(n7942), .ZN(n7958)
         );
  NAND2_X1 U5414 ( .A1(n6664), .A2(n4892), .ZN(n5959) );
  AND2_X1 U5415 ( .A1(n7437), .A2(n5112), .ZN(n4851) );
  OR2_X1 U5416 ( .A1(n7958), .A2(n7957), .ZN(n9127) );
  NAND2_X1 U5417 ( .A1(n7958), .A2(n7957), .ZN(n9128) );
  NAND2_X1 U5418 ( .A1(n6616), .A2(n6440), .ZN(n4875) );
  NAND2_X1 U5419 ( .A1(n6617), .A2(n6442), .ZN(n4874) );
  NAND2_X1 U5420 ( .A1(n6843), .A2(n9069), .ZN(n4887) );
  OR2_X1 U5421 ( .A1(n6842), .A2(n6841), .ZN(n6847) );
  NAND2_X1 U5422 ( .A1(n7551), .A2(n7550), .ZN(n7933) );
  XNOR2_X1 U5423 ( .A(n7572), .B(n4739), .ZN(n7566) );
  OR2_X1 U5424 ( .A1(n6004), .A2(n6003), .ZN(n4724) );
  AND2_X1 U5425 ( .A1(n4724), .A2(n4723), .ZN(n6017) );
  NAND2_X1 U5426 ( .A1(n6015), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4723) );
  OR2_X1 U5427 ( .A1(n6017), .A2(n6016), .ZN(n4722) );
  OR2_X1 U5428 ( .A1(n6048), .A2(n6047), .ZN(n4728) );
  AND2_X1 U5429 ( .A1(n4728), .A2(n4727), .ZN(n6063) );
  NAND2_X1 U5430 ( .A1(n6061), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4727) );
  OR2_X1 U5431 ( .A1(n6063), .A2(n6062), .ZN(n4726) );
  NOR2_X1 U5432 ( .A1(n9179), .A2(n4660), .ZN(n9192) );
  AND2_X1 U5433 ( .A1(n9187), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n4660) );
  XNOR2_X1 U5434 ( .A(n9250), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n4736) );
  AND2_X1 U5435 ( .A1(n8184), .A2(n8185), .ZN(n9289) );
  AND2_X1 U5436 ( .A1(n8195), .A2(n9307), .ZN(n9322) );
  OR2_X1 U5437 ( .A1(n9323), .A2(n9322), .ZN(n9325) );
  AND2_X1 U5438 ( .A1(n8196), .A2(n9306), .ZN(n9344) );
  INV_X1 U5439 ( .A(n4745), .ZN(n4744) );
  OAI21_X1 U5440 ( .B1(n4518), .B2(n4746), .A(n9351), .ZN(n4745) );
  INV_X1 U5441 ( .A(n9303), .ZN(n4746) );
  OR2_X1 U5442 ( .A1(n9390), .A2(n9374), .ZN(n9302) );
  NAND2_X1 U5443 ( .A1(n9384), .A2(n4518), .ZN(n9368) );
  NOR2_X1 U5444 ( .A1(n9286), .A2(n5103), .ZN(n5102) );
  INV_X1 U5445 ( .A(n5104), .ZN(n5103) );
  INV_X1 U5446 ( .A(n5100), .ZN(n5099) );
  OAI22_X1 U5447 ( .A1(n9286), .A2(n5101), .B1(n9390), .B2(n9649), .ZN(n5100)
         );
  NAND2_X1 U5448 ( .A1(n5104), .A2(n4534), .ZN(n5101) );
  NAND2_X1 U5449 ( .A1(n9408), .A2(n9658), .ZN(n5104) );
  NAND2_X1 U5450 ( .A1(n9302), .A2(n8169), .ZN(n9382) );
  NAND2_X1 U5451 ( .A1(n9428), .A2(n9282), .ZN(n5059) );
  NAND2_X1 U5452 ( .A1(n9453), .A2(n4516), .ZN(n9429) );
  AND2_X1 U5453 ( .A1(n9296), .A2(n8200), .ZN(n9454) );
  NAND2_X1 U5454 ( .A1(n4577), .A2(n4519), .ZN(n5083) );
  NOR2_X1 U5455 ( .A1(n9476), .A2(n4761), .ZN(n4760) );
  INV_X1 U5456 ( .A(n4756), .ZN(n4755) );
  OAI21_X1 U5457 ( .B1(n4759), .B2(n4757), .A(n9534), .ZN(n4756) );
  AND2_X1 U5458 ( .A1(n8205), .A2(n8242), .ZN(n9534) );
  AND2_X1 U5459 ( .A1(n8145), .A2(n8241), .ZN(n9552) );
  NAND2_X1 U5460 ( .A1(n9578), .A2(n4759), .ZN(n9550) );
  NAND2_X1 U5461 ( .A1(n5060), .A2(n5063), .ZN(n9573) );
  AOI21_X1 U5462 ( .B1(n8236), .B2(n5064), .A(n4568), .ZN(n5063) );
  OR2_X1 U5463 ( .A1(n7346), .A2(n7345), .ZN(n7371) );
  OR2_X1 U5464 ( .A1(n7449), .A2(n9166), .ZN(n7380) );
  NAND2_X1 U5465 ( .A1(n7343), .A2(n8223), .ZN(n7381) );
  OR2_X1 U5466 ( .A1(n7241), .A2(n7240), .ZN(n7266) );
  AND4_X1 U5467 ( .A1(n7271), .A2(n7270), .A3(n7269), .A4(n7268), .ZN(n9046)
         );
  AND2_X1 U5468 ( .A1(n8084), .A2(n8219), .ZN(n4740) );
  INV_X1 U5469 ( .A(n5076), .ZN(n5075) );
  OAI22_X1 U5470 ( .A1(n7235), .A2(n7032), .B1(n7318), .B2(n9169), .ZN(n5076)
         );
  AOI21_X1 U5471 ( .B1(n5075), .B2(n7235), .A(n5074), .ZN(n5073) );
  INV_X1 U5472 ( .A(n7237), .ZN(n5074) );
  AND2_X1 U5473 ( .A1(n8123), .A2(n8121), .ZN(n7235) );
  NAND2_X1 U5474 ( .A1(n6724), .A2(n6723), .ZN(n7010) );
  NAND2_X1 U5475 ( .A1(n6700), .A2(n8213), .ZN(n4611) );
  OR2_X1 U5476 ( .A1(n6912), .A2(n8268), .ZN(n9494) );
  NAND2_X1 U5477 ( .A1(n7474), .A2(n7473), .ZN(n8105) );
  NAND2_X1 U5478 ( .A1(n7480), .A2(n7479), .ZN(n9265) );
  NAND2_X1 U5479 ( .A1(n7508), .A2(n7507), .ZN(n9272) );
  AND4_X1 U5480 ( .A1(n7839), .A2(n7838), .A3(n7837), .A4(n7836), .ZN(n9732)
         );
  AND3_X1 U5481 ( .A1(n7037), .A2(n7036), .A3(n7035), .ZN(n9811) );
  NAND2_X1 U5482 ( .A1(n6663), .A2(n8259), .ZN(n9708) );
  OR2_X1 U5483 ( .A1(n7229), .A2(n7572), .ZN(n5054) );
  NAND2_X1 U5484 ( .A1(n5968), .A2(n8259), .ZN(n9731) );
  INV_X1 U5485 ( .A(n9693), .ZN(n9713) );
  NAND2_X1 U5486 ( .A1(n5958), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6097) );
  AND2_X1 U5487 ( .A1(n6101), .A2(n6100), .ZN(n6395) );
  OR2_X1 U5488 ( .A1(n5925), .A2(n5854), .ZN(n5923) );
  XNOR2_X1 U5489 ( .A(n5704), .B(n5703), .ZN(n8308) );
  NAND2_X1 U5490 ( .A1(n4982), .A2(n5690), .ZN(n5704) );
  NAND2_X1 U5491 ( .A1(n5689), .A2(n5688), .ZN(n4982) );
  INV_X1 U5492 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5850) );
  INV_X1 U5493 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5847) );
  XNOR2_X1 U5494 ( .A(n5635), .B(n5634), .ZN(n7490) );
  NAND2_X1 U5495 ( .A1(n5606), .A2(n5605), .ZN(n5618) );
  XNOR2_X1 U5496 ( .A(n5858), .B(P1_IR_REG_23__SCAN_IN), .ZN(n6480) );
  XNOR2_X1 U5497 ( .A(n5936), .B(P1_IR_REG_21__SCAN_IN), .ZN(n8075) );
  NAND2_X1 U5498 ( .A1(n5844), .A2(n5068), .ZN(n6597) );
  INV_X1 U5499 ( .A(n6055), .ZN(n5068) );
  NAND2_X1 U5500 ( .A1(n4995), .A2(n5494), .ZN(n5510) );
  XNOR2_X1 U5501 ( .A(n5491), .B(n5477), .ZN(n7515) );
  OR2_X1 U5502 ( .A1(n6266), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n6267) );
  NAND2_X1 U5503 ( .A1(n5436), .A2(n5435), .ZN(n5455) );
  AND2_X1 U5504 ( .A1(n5435), .A2(n5420), .ZN(n5421) );
  INV_X1 U5505 ( .A(n4986), .ZN(n4696) );
  AOI21_X1 U5506 ( .B1(n4992), .B2(n4989), .A(n4987), .ZN(n4986) );
  INV_X1 U5507 ( .A(n5416), .ZN(n4987) );
  NOR2_X1 U5508 ( .A1(n4698), .A2(n4988), .ZN(n4697) );
  INV_X1 U5509 ( .A(n4699), .ZN(n4698) );
  INV_X1 U5510 ( .A(n4989), .ZN(n4988) );
  AND2_X1 U5511 ( .A1(n4994), .A2(n4542), .ZN(n4989) );
  INV_X1 U5512 ( .A(n5400), .ZN(n4994) );
  NAND2_X1 U5513 ( .A1(n5382), .A2(n4991), .ZN(n4990) );
  NAND2_X1 U5514 ( .A1(n4953), .A2(n5285), .ZN(n4682) );
  NAND2_X1 U5515 ( .A1(n5246), .A2(n4683), .ZN(n4681) );
  AND2_X1 U5516 ( .A1(n5260), .A2(n4684), .ZN(n4683) );
  AND2_X1 U5517 ( .A1(n5245), .A2(n5285), .ZN(n4684) );
  NAND3_X1 U5518 ( .A1(n4681), .A2(n5290), .A3(n4682), .ZN(n5303) );
  NOR2_X1 U5519 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5056) );
  OR2_X1 U5520 ( .A1(n8025), .A2(n8357), .ZN(n8026) );
  NAND2_X1 U5521 ( .A1(n5915), .A2(n8788), .ZN(n8419) );
  INV_X1 U5522 ( .A(n5139), .ZN(n7784) );
  INV_X1 U5523 ( .A(n7296), .ZN(n7789) );
  NAND2_X1 U5524 ( .A1(n9867), .A2(n4603), .ZN(n6162) );
  OR2_X1 U5525 ( .A1(n6160), .A2(n6161), .ZN(n4603) );
  OR2_X1 U5526 ( .A1(n6878), .A2(n6879), .ZN(n4667) );
  INV_X1 U5527 ( .A(n4665), .ZN(n7131) );
  INV_X1 U5528 ( .A(n8546), .ZN(n4676) );
  NAND2_X1 U5529 ( .A1(n8547), .A2(n8558), .ZN(n4675) );
  NOR2_X1 U5530 ( .A1(n8518), .A2(n8517), .ZN(n8552) );
  OAI21_X1 U5531 ( .B1(n9958), .B2(n4679), .A(n4678), .ZN(n4677) );
  NAND2_X1 U5532 ( .A1(n4680), .A2(n8545), .ZN(n4679) );
  INV_X1 U5533 ( .A(n8555), .ZN(n4678) );
  INV_X1 U5534 ( .A(n8543), .ZN(n4680) );
  NOR2_X1 U5535 ( .A1(n8555), .A2(n8554), .ZN(n8556) );
  OAI21_X1 U5536 ( .B1(n8559), .B2(n8558), .A(n8557), .ZN(n8565) );
  NAND2_X1 U5537 ( .A1(n4827), .A2(n4826), .ZN(n4830) );
  AOI21_X1 U5538 ( .B1(n8516), .B2(n4828), .A(n8551), .ZN(n4826) );
  NAND2_X1 U5539 ( .A1(n9961), .A2(n4828), .ZN(n4827) );
  INV_X1 U5540 ( .A(n8788), .ZN(n8756) );
  NAND2_X1 U5541 ( .A1(n5408), .A2(n5407), .ZN(n7688) );
  OR2_X1 U5542 ( .A1(n7252), .A2(n5222), .ZN(n5372) );
  INV_X1 U5543 ( .A(n8793), .ZN(n8784) );
  AOI21_X1 U5544 ( .B1(n7549), .B2(n7579), .A(n5708), .ZN(n7619) );
  NAND2_X1 U5545 ( .A1(n5043), .A2(n5040), .ZN(n5039) );
  NAND2_X1 U5546 ( .A1(n8582), .A2(n10019), .ZN(n5043) );
  NOR2_X1 U5547 ( .A1(n8577), .A2(n5777), .ZN(n5040) );
  OR2_X1 U5548 ( .A1(n10070), .A2(n10062), .ZN(n8933) );
  NAND2_X1 U5549 ( .A1(n5426), .A2(n5425), .ZN(n8971) );
  AND2_X1 U5550 ( .A1(n8298), .A2(n9143), .ZN(n4870) );
  NAND2_X1 U5551 ( .A1(n7503), .A2(n7502), .ZN(n9431) );
  AND4_X1 U5552 ( .A1(n7869), .A2(n7868), .A3(n7867), .A4(n7866), .ZN(n9707)
         );
  INV_X1 U5553 ( .A(n9495), .ZN(n9696) );
  NAND2_X1 U5554 ( .A1(n7532), .A2(n7531), .ZN(n9676) );
  AND2_X1 U5555 ( .A1(n9144), .A2(n9145), .ZN(n4873) );
  INV_X1 U5556 ( .A(n9164), .ZN(n9143) );
  OAI21_X2 U5557 ( .B1(n6476), .B2(n6475), .A(n9557), .ZN(n9162) );
  AOI21_X1 U5558 ( .B1(n9328), .B2(n7962), .A(n6361), .ZN(n9607) );
  XNOR2_X1 U5559 ( .A(n7572), .B(n4644), .ZN(n7563) );
  NOR2_X1 U5560 ( .A1(n6958), .A2(n6957), .ZN(n9179) );
  XNOR2_X1 U5561 ( .A(n9192), .B(n9201), .ZN(n9181) );
  NOR2_X1 U5562 ( .A1(n9212), .A2(n4729), .ZN(n9213) );
  AND2_X1 U5563 ( .A1(n9217), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4729) );
  NAND2_X1 U5564 ( .A1(n9213), .A2(n9214), .ZN(n9228) );
  NAND2_X1 U5565 ( .A1(n7483), .A2(n7482), .ZN(n8101) );
  INV_X1 U5566 ( .A(n9661), .ZN(n9422) );
  INV_X1 U5567 ( .A(n9776), .ZN(n9568) );
  NAND2_X1 U5568 ( .A1(n7255), .A2(n7254), .ZN(n7422) );
  NAND2_X2 U5569 ( .A1(n8271), .A2(n6474), .ZN(n9557) );
  INV_X1 U5570 ( .A(n6473), .ZN(n6474) );
  OAI21_X1 U5571 ( .B1(n7071), .B2(n8113), .A(n4633), .ZN(n4632) );
  NAND2_X1 U5572 ( .A1(n7704), .A2(n7703), .ZN(n4784) );
  NAND2_X1 U5573 ( .A1(n7724), .A2(n4777), .ZN(n4776) );
  AND2_X1 U5574 ( .A1(n7723), .A2(n7722), .ZN(n4777) );
  INV_X1 U5575 ( .A(n4617), .ZN(n4616) );
  AOI21_X1 U5576 ( .B1(n4617), .B2(n4615), .A(n4573), .ZN(n4614) );
  INV_X1 U5577 ( .A(n4619), .ZN(n4615) );
  NAND2_X1 U5578 ( .A1(n4775), .A2(n4773), .ZN(n4772) );
  NOR2_X1 U5579 ( .A1(n7728), .A2(n4774), .ZN(n4773) );
  NAND2_X1 U5580 ( .A1(n4776), .A2(n7775), .ZN(n4775) );
  AND2_X1 U5581 ( .A1(n7726), .A2(n7768), .ZN(n4774) );
  AOI21_X1 U5582 ( .B1(n8147), .B2(n8204), .A(n4643), .ZN(n4642) );
  NAND2_X1 U5583 ( .A1(n8244), .A2(n8277), .ZN(n4643) );
  AND2_X1 U5584 ( .A1(n7744), .A2(n7775), .ZN(n4786) );
  OAI21_X1 U5585 ( .B1(n4623), .B2(n4622), .A(n8170), .ZN(n8176) );
  AOI21_X1 U5586 ( .B1(n8159), .B2(n8158), .A(n4541), .ZN(n4622) );
  AOI21_X1 U5587 ( .B1(n8182), .B2(n8181), .A(n4639), .ZN(n4638) );
  OAI21_X1 U5588 ( .B1(n8175), .B2(n8194), .A(n8195), .ZN(n4639) );
  INV_X1 U5589 ( .A(n7760), .ZN(n4764) );
  INV_X1 U5590 ( .A(n8184), .ZN(n5004) );
  NAND2_X1 U5591 ( .A1(n5141), .A2(n5036), .ZN(n5035) );
  INV_X1 U5592 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5036) );
  AND2_X1 U5593 ( .A1(n7406), .A2(n7306), .ZN(n4888) );
  NAND2_X1 U5594 ( .A1(n9061), .A2(n9060), .ZN(n4866) );
  NAND2_X1 U5595 ( .A1(n4635), .A2(n5002), .ZN(n8189) );
  AOI21_X1 U5596 ( .B1(n5004), .B2(n8277), .A(n5003), .ZN(n5002) );
  NAND2_X1 U5597 ( .A1(n4636), .A2(n9289), .ZN(n4635) );
  NOR2_X1 U5598 ( .A1(n8185), .A2(n8277), .ZN(n5003) );
  NAND2_X1 U5599 ( .A1(n4981), .A2(n4980), .ZN(n7455) );
  AOI21_X1 U5600 ( .B1(n4983), .B2(n4985), .A(n4599), .ZN(n4980) );
  INV_X1 U5601 ( .A(n4970), .ZN(n4969) );
  OAI21_X1 U5602 ( .B1(n5605), .B2(n4971), .A(n5634), .ZN(n4970) );
  INV_X1 U5603 ( .A(n5617), .ZN(n4971) );
  NOR2_X1 U5604 ( .A1(n5454), .A2(SI_14_), .ZN(n4998) );
  AND2_X1 U5605 ( .A1(n5435), .A2(n5000), .ZN(n4999) );
  NAND2_X1 U5606 ( .A1(n5454), .A2(SI_14_), .ZN(n5000) );
  INV_X1 U5607 ( .A(n5339), .ZN(n4958) );
  INV_X1 U5608 ( .A(n5308), .ZN(n4957) );
  INV_X1 U5609 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5148) );
  INV_X1 U5610 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10463) );
  NAND2_X1 U5611 ( .A1(n7582), .A2(n7581), .ZN(n7583) );
  OAI21_X1 U5612 ( .B1(n7615), .B2(n7626), .A(n5824), .ZN(n7616) );
  NAND2_X1 U5613 ( .A1(n4574), .A2(n6242), .ZN(n4843) );
  NAND2_X1 U5614 ( .A1(n4840), .A2(n4843), .ZN(n6510) );
  AND2_X1 U5615 ( .A1(n4844), .A2(n4841), .ZN(n4840) );
  NAND2_X1 U5616 ( .A1(n6505), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4841) );
  AOI21_X1 U5617 ( .B1(n8527), .B2(n8541), .A(n8526), .ZN(n8529) );
  INV_X1 U5618 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10479) );
  OAI21_X1 U5619 ( .B1(n5750), .B2(n5009), .A(n8676), .ZN(n5008) );
  OR2_X1 U5620 ( .A1(n5554), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U5621 ( .A1(n5014), .A2(n5016), .ZN(n5013) );
  OR2_X1 U5622 ( .A1(n10059), .A2(n7186), .ZN(n7679) );
  OR2_X1 U5623 ( .A1(n10045), .A2(n6947), .ZN(n7655) );
  NAND2_X1 U5624 ( .A1(n10008), .A2(n6296), .ZN(n7644) );
  NAND2_X1 U5625 ( .A1(n6936), .A2(n9997), .ZN(n7658) );
  NAND2_X1 U5626 ( .A1(n8790), .A2(n5870), .ZN(n7633) );
  AOI21_X1 U5627 ( .B1(n5028), .B2(n5030), .A(n4567), .ZN(n5027) );
  INV_X1 U5628 ( .A(n5032), .ZN(n5028) );
  INV_X1 U5629 ( .A(n5030), .ZN(n5029) );
  INV_X1 U5630 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5802) );
  INV_X1 U5631 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5515) );
  NAND2_X1 U5632 ( .A1(n7302), .A2(n7301), .ZN(n4889) );
  INV_X1 U5633 ( .A(n7883), .ZN(n8289) );
  INV_X1 U5634 ( .A(n8276), .ZN(n8260) );
  INV_X1 U5635 ( .A(n8070), .ZN(n4688) );
  NAND2_X1 U5636 ( .A1(n8251), .A2(n8071), .ZN(n4687) );
  NOR2_X1 U5637 ( .A1(n8069), .A2(n8178), .ZN(n8251) );
  OAI21_X1 U5638 ( .B1(n8189), .B2(n9265), .A(n5001), .ZN(n8186) );
  NAND2_X1 U5639 ( .A1(n9265), .A2(n8277), .ZN(n5001) );
  NAND2_X1 U5640 ( .A1(n9408), .A2(n9285), .ZN(n9381) );
  INV_X1 U5641 ( .A(n5109), .ZN(n5058) );
  NOR2_X1 U5642 ( .A1(n9689), .A2(n4713), .ZN(n4712) );
  INV_X1 U5643 ( .A(n4714), .ZN(n4713) );
  NOR2_X1 U5644 ( .A1(n9696), .A2(n9528), .ZN(n4714) );
  INV_X1 U5645 ( .A(n8241), .ZN(n4757) );
  INV_X1 U5646 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7370) );
  NOR2_X1 U5647 ( .A1(n5065), .A2(n5062), .ZN(n5061) );
  INV_X1 U5648 ( .A(n8223), .ZN(n5062) );
  INV_X1 U5649 ( .A(n8236), .ZN(n5065) );
  INV_X1 U5650 ( .A(n7380), .ZN(n5064) );
  INV_X1 U5651 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7240) );
  NOR2_X1 U5652 ( .A1(n7318), .A2(n7113), .ZN(n4708) );
  NOR2_X1 U5653 ( .A1(n9592), .A2(n9568), .ZN(n9565) );
  NOR2_X1 U5654 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5943) );
  XNOR2_X1 U5655 ( .A(n7455), .B(n7456), .ZN(n7453) );
  AND2_X1 U5656 ( .A1(n5690), .A2(n5674), .ZN(n5688) );
  AND2_X1 U5657 ( .A1(n5670), .A2(n5657), .ZN(n5668) );
  AND2_X1 U5658 ( .A1(n5653), .A2(n5639), .ZN(n5651) );
  AOI21_X1 U5659 ( .B1(n5579), .B2(n5115), .A(n5114), .ZN(n5584) );
  AND2_X1 U5660 ( .A1(n5560), .A2(n5561), .ZN(n4979) );
  OR2_X1 U5661 ( .A1(n5560), .A2(n5561), .ZN(n4978) );
  INV_X1 U5662 ( .A(SI_20_), .ZN(n5561) );
  INV_X1 U5663 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6092) );
  INV_X1 U5664 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5841) );
  INV_X1 U5665 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5842) );
  INV_X1 U5666 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5843) );
  NAND2_X1 U5667 ( .A1(n5492), .A2(n5107), .ZN(n4995) );
  INV_X1 U5668 ( .A(SI_13_), .ZN(n10246) );
  NOR2_X1 U5669 ( .A1(n4696), .A2(n4691), .ZN(n4690) );
  INV_X1 U5670 ( .A(n5360), .ZN(n4691) );
  INV_X1 U5671 ( .A(n5397), .ZN(n4993) );
  INV_X1 U5672 ( .A(SI_6_), .ZN(n10338) );
  OAI21_X1 U5673 ( .B1(n7468), .B2(n4707), .A(n4706), .ZN(n5247) );
  NAND2_X1 U5674 ( .A1(n7468), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n4706) );
  OAI22_X1 U5675 ( .A1(n7468), .A2(n5196), .B1(n6433), .B2(n5195), .ZN(n5197)
         );
  NAND2_X1 U5676 ( .A1(n5541), .A2(n10463), .ZN(n5554) );
  INV_X1 U5677 ( .A(n5542), .ZN(n5541) );
  INV_X1 U5678 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10476) );
  NAND2_X1 U5679 ( .A1(n4932), .A2(n8437), .ZN(n4931) );
  INV_X1 U5680 ( .A(n4939), .ZN(n4937) );
  INV_X1 U5681 ( .A(n8372), .ZN(n4936) );
  NAND2_X1 U5682 ( .A1(n5503), .A2(n5502), .ZN(n5521) );
  INV_X1 U5683 ( .A(n5504), .ZN(n5503) );
  AOI21_X1 U5684 ( .B1(n4927), .B2(n4928), .A(n4926), .ZN(n4925) );
  INV_X1 U5685 ( .A(n8387), .ZN(n4926) );
  INV_X1 U5686 ( .A(n5720), .ZN(n6154) );
  NAND2_X1 U5687 ( .A1(n9869), .A2(n9868), .ZN(n9867) );
  OAI211_X1 U5688 ( .C1(n9882), .C2(n4823), .A(n4821), .B(n4820), .ZN(n6174)
         );
  NOR2_X1 U5689 ( .A1(n4663), .A2(n6164), .ZN(n4662) );
  NAND2_X1 U5690 ( .A1(n6174), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6275) );
  NAND2_X1 U5691 ( .A1(n6241), .A2(n6337), .ZN(n4845) );
  NOR2_X1 U5692 ( .A1(n4842), .A2(n6342), .ZN(n6340) );
  NAND2_X1 U5693 ( .A1(n4845), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4842) );
  NOR2_X1 U5694 ( .A1(n6509), .A2(n6348), .ZN(n4670) );
  OR2_X1 U5695 ( .A1(n5325), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U5696 ( .A1(n6510), .A2(n6816), .ZN(n8458) );
  NOR2_X1 U5697 ( .A1(n6511), .A2(n6500), .ZN(n8461) );
  OAI21_X1 U5698 ( .B1(n6807), .B2(n4838), .A(n4837), .ZN(n7134) );
  NAND2_X1 U5699 ( .A1(n4839), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4838) );
  NAND2_X1 U5700 ( .A1(n6894), .A2(n4839), .ZN(n4837) );
  INV_X1 U5701 ( .A(n6897), .ZN(n4839) );
  INV_X1 U5702 ( .A(n4849), .ZN(n8470) );
  NAND2_X1 U5703 ( .A1(n8490), .A2(n8491), .ZN(n8523) );
  NAND2_X1 U5704 ( .A1(n4904), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4903) );
  NAND2_X1 U5705 ( .A1(n8537), .A2(n4904), .ZN(n4902) );
  INV_X1 U5706 ( .A(n9942), .ZN(n4904) );
  NAND2_X1 U5707 ( .A1(n4907), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4906) );
  INV_X1 U5708 ( .A(n8545), .ZN(n4907) );
  INV_X1 U5709 ( .A(n8517), .ZN(n4828) );
  OR2_X1 U5710 ( .A1(n5694), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5709) );
  AOI21_X1 U5711 ( .B1(n4797), .B2(n4795), .A(n4794), .ZN(n4793) );
  INV_X1 U5712 ( .A(n7758), .ZN(n4794) );
  NOR2_X1 U5713 ( .A1(n4798), .A2(n5667), .ZN(n4795) );
  OR2_X1 U5714 ( .A1(n5590), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5610) );
  AND2_X1 U5715 ( .A1(n5754), .A2(n7742), .ZN(n8656) );
  AOI21_X1 U5716 ( .B1(n4813), .B2(n4816), .A(n7735), .ZN(n4812) );
  INV_X1 U5717 ( .A(n4817), .ZN(n4816) );
  INV_X1 U5718 ( .A(n8656), .ZN(n8659) );
  NOR2_X1 U5719 ( .A1(n7734), .A2(n4818), .ZN(n4817) );
  INV_X1 U5720 ( .A(n7723), .ZN(n4818) );
  NAND2_X1 U5721 ( .A1(n5010), .A2(n5750), .ZN(n8680) );
  INV_X1 U5722 ( .A(n8682), .ZN(n5010) );
  NAND2_X1 U5723 ( .A1(n5037), .A2(n5747), .ZN(n8691) );
  NAND2_X1 U5724 ( .A1(n5462), .A2(n5461), .ZN(n5485) );
  INV_X1 U5725 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5461) );
  OR2_X1 U5726 ( .A1(n5447), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5463) );
  OR2_X1 U5727 ( .A1(n5388), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5410) );
  OR2_X1 U5728 ( .A1(n5374), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5388) );
  NOR2_X1 U5729 ( .A1(n10026), .A2(n10037), .ZN(n5053) );
  OR2_X1 U5730 ( .A1(n5330), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5350) );
  OR2_X1 U5731 ( .A1(n5295), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5316) );
  OAI21_X1 U5732 ( .B1(n6414), .B2(n5730), .A(n5729), .ZN(n6757) );
  NAND2_X1 U5733 ( .A1(n7644), .A2(n7658), .ZN(n6920) );
  OR2_X1 U5734 ( .A1(n5214), .A2(n6778), .ZN(n5206) );
  AND2_X1 U5735 ( .A1(n5828), .A2(n5898), .ZN(n6420) );
  OR2_X1 U5736 ( .A1(n7794), .A2(n7793), .ZN(n8807) );
  INV_X1 U5737 ( .A(n5046), .ZN(n5045) );
  OAI21_X1 U5738 ( .B1(n4517), .B2(n4535), .A(n7622), .ZN(n5046) );
  NAND2_X1 U5739 ( .A1(n4789), .A2(n4788), .ZN(n8587) );
  AOI21_X1 U5740 ( .B1(n4790), .B2(n4796), .A(n4522), .ZN(n4788) );
  AND2_X1 U5741 ( .A1(n7746), .A2(n8640), .ZN(n8649) );
  AOI21_X1 U5742 ( .B1(n4804), .B2(n4806), .A(n7694), .ZN(n4803) );
  INV_X1 U5743 ( .A(n4805), .ZN(n4804) );
  NOR2_X1 U5744 ( .A1(n5897), .A2(n5823), .ZN(n5911) );
  INV_X1 U5745 ( .A(n10019), .ZN(n10064) );
  XNOR2_X1 U5746 ( .A(n5801), .B(n5802), .ZN(n6166) );
  INV_X1 U5747 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5173) );
  INV_X1 U5748 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5144) );
  NAND2_X1 U5749 ( .A1(n5124), .A2(n5123), .ZN(n5478) );
  NOR2_X1 U5750 ( .A1(n5122), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n5123) );
  INV_X1 U5751 ( .A(n5424), .ZN(n5124) );
  NAND2_X1 U5752 ( .A1(n4950), .A2(n5479), .ZN(n5498) );
  AND2_X1 U5753 ( .A1(n5383), .A2(n5129), .ZN(n5404) );
  OR2_X1 U5754 ( .A1(n7371), .A2(n7370), .ZN(n7834) );
  NAND2_X1 U5755 ( .A1(n9115), .A2(n4890), .ZN(n8998) );
  NOR2_X1 U5756 ( .A1(n7843), .A2(n4891), .ZN(n4890) );
  INV_X1 U5757 ( .A(n7832), .ZN(n4891) );
  OR2_X1 U5758 ( .A1(n7957), .A2(n9129), .ZN(n4883) );
  AND2_X1 U5759 ( .A1(n8007), .A2(n8006), .ZN(n8009) );
  NAND2_X1 U5760 ( .A1(n6912), .A2(n4561), .ZN(n4893) );
  OR2_X1 U5761 ( .A1(n8075), .A2(n9343), .ZN(n4894) );
  AND2_X1 U5762 ( .A1(n7928), .A2(n4860), .ZN(n4859) );
  NAND2_X1 U5763 ( .A1(n4539), .A2(n4861), .ZN(n4860) );
  NOR2_X1 U5764 ( .A1(n4864), .A2(n4867), .ZN(n4861) );
  NAND2_X1 U5765 ( .A1(n4859), .A2(n4862), .ZN(n4857) );
  NAND2_X1 U5766 ( .A1(n4539), .A2(n4863), .ZN(n4862) );
  INV_X1 U5767 ( .A(n4864), .ZN(n4863) );
  NAND2_X1 U5768 ( .A1(n4854), .A2(n4852), .ZN(n9042) );
  NOR2_X1 U5769 ( .A1(n4853), .A2(n7816), .ZN(n4852) );
  INV_X1 U5770 ( .A(n9043), .ZN(n4853) );
  AND2_X1 U5771 ( .A1(n7886), .A2(n7885), .ZN(n9082) );
  INV_X1 U5772 ( .A(n4881), .ZN(n4880) );
  AND2_X1 U5773 ( .A1(n7972), .A2(n4878), .ZN(n4877) );
  OR2_X1 U5774 ( .A1(n6430), .A2(n5961), .ZN(n5965) );
  NAND2_X1 U5775 ( .A1(n5965), .A2(n5964), .ZN(n6432) );
  INV_X1 U5776 ( .A(n4858), .ZN(n9024) );
  AOI21_X1 U5777 ( .B1(n9063), .B2(n4867), .A(n4864), .ZN(n4858) );
  NOR2_X1 U5778 ( .A1(n6479), .A2(n6468), .ZN(n6486) );
  OR2_X1 U5779 ( .A1(n6222), .A2(n6221), .ZN(n4656) );
  AND2_X1 U5780 ( .A1(n4722), .A2(n4721), .ZN(n6031) );
  NAND2_X1 U5781 ( .A1(n6029), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4721) );
  OR2_X1 U5782 ( .A1(n6044), .A2(n6043), .ZN(n4654) );
  OR2_X1 U5783 ( .A1(n6059), .A2(n6058), .ZN(n4652) );
  AND2_X1 U5784 ( .A1(n4726), .A2(n4725), .ZN(n6206) );
  NAND2_X1 U5785 ( .A1(n6202), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4725) );
  AND2_X1 U5786 ( .A1(n4652), .A2(n4651), .ZN(n6196) );
  NAND2_X1 U5787 ( .A1(n6202), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n4651) );
  NOR2_X1 U5788 ( .A1(n4731), .A2(n6641), .ZN(n6642) );
  AND2_X1 U5789 ( .A1(n7340), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4731) );
  NAND2_X1 U5790 ( .A1(n6642), .A2(n6643), .ZN(n6796) );
  NOR2_X1 U5791 ( .A1(n9186), .A2(n4737), .ZN(n9202) );
  AND2_X1 U5792 ( .A1(n9187), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4737) );
  NAND2_X1 U5793 ( .A1(n9216), .A2(n4650), .ZN(n9218) );
  OR2_X1 U5794 ( .A1(n9217), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n4650) );
  NAND2_X1 U5795 ( .A1(n9218), .A2(n9219), .ZN(n9240) );
  INV_X1 U5796 ( .A(n9289), .ZN(n9308) );
  AND3_X1 U5797 ( .A1(n6121), .A2(n6120), .A3(n6119), .ZN(n9311) );
  OR2_X1 U5798 ( .A1(n7987), .A2(n6234), .ZN(n9294) );
  AND2_X1 U5799 ( .A1(n7995), .A2(n7994), .ZN(n9341) );
  OR2_X1 U5800 ( .A1(n9356), .A2(n7988), .ZN(n7995) );
  NAND2_X1 U5801 ( .A1(n9389), .A2(n4718), .ZN(n9353) );
  AOI21_X1 U5802 ( .B1(n5096), .B2(n5095), .A(n4548), .ZN(n5094) );
  INV_X1 U5803 ( .A(n5102), .ZN(n5095) );
  AND3_X1 U5804 ( .A1(n7965), .A2(n7964), .A3(n7963), .ZN(n9374) );
  NAND2_X1 U5805 ( .A1(n9389), .A2(n9639), .ZN(n9369) );
  OR2_X1 U5806 ( .A1(n9408), .A2(n9417), .ZN(n9401) );
  OR2_X1 U5807 ( .A1(n7906), .A2(n7892), .ZN(n7934) );
  AND2_X1 U5808 ( .A1(n9536), .A2(n4710), .ZN(n9468) );
  AND2_X1 U5809 ( .A1(n4712), .A2(n4711), .ZN(n4710) );
  NAND2_X1 U5810 ( .A1(n5078), .A2(n5077), .ZN(n9444) );
  AOI21_X1 U5811 ( .B1(n5080), .B2(n5082), .A(n4591), .ZN(n5077) );
  NAND2_X1 U5812 ( .A1(n9536), .A2(n4712), .ZN(n9479) );
  OR2_X1 U5813 ( .A1(n7864), .A2(n7863), .ZN(n9087) );
  NAND2_X1 U5814 ( .A1(n9536), .A2(n9702), .ZN(n9522) );
  AND2_X1 U5815 ( .A1(n9565), .A2(n9546), .ZN(n9536) );
  INV_X1 U5816 ( .A(n9719), .ZN(n9525) );
  NAND2_X1 U5817 ( .A1(n9572), .A2(n9273), .ZN(n9555) );
  NAND2_X1 U5818 ( .A1(n9779), .A2(n9562), .ZN(n9273) );
  INV_X1 U5819 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7345) );
  NAND2_X1 U5820 ( .A1(n7364), .A2(n7363), .ZN(n4743) );
  AND4_X1 U5821 ( .A1(n7246), .A2(n7245), .A3(n7244), .A4(n7243), .ZN(n7446)
         );
  AND4_X1 U5822 ( .A1(n7351), .A2(n7350), .A3(n7349), .A4(n7348), .ZN(n9580)
         );
  AOI21_X1 U5823 ( .B1(n5073), .B2(n5076), .A(n4572), .ZN(n5071) );
  INV_X1 U5824 ( .A(n5073), .ZN(n5072) );
  NAND2_X1 U5825 ( .A1(n7098), .A2(n4708), .ZN(n7279) );
  NAND2_X1 U5826 ( .A1(n7098), .A2(n7260), .ZN(n7097) );
  NOR2_X1 U5827 ( .A1(n7013), .A2(n9071), .ZN(n7078) );
  INV_X1 U5828 ( .A(n8210), .ZN(n4610) );
  AOI21_X1 U5829 ( .B1(n6703), .B2(n6683), .A(n6682), .ZN(n6724) );
  NOR2_X1 U5830 ( .A1(n6706), .A2(n6707), .ZN(n6705) );
  OAI211_X1 U5831 ( .C1(n6399), .C2(n6469), .A(n6485), .B(n6912), .ZN(n7355)
         );
  OR2_X1 U5832 ( .A1(n6673), .A2(n6662), .ZN(n6680) );
  AND2_X1 U5833 ( .A1(n7803), .A2(n7802), .ZN(n9627) );
  NAND2_X1 U5834 ( .A1(n4705), .A2(n7492), .ZN(n9390) );
  NAND2_X1 U5835 ( .A1(n7490), .A2(n7533), .ZN(n4705) );
  AND2_X1 U5836 ( .A1(n7500), .A2(n7499), .ZN(n9661) );
  INV_X1 U5837 ( .A(n9485), .ZN(n9686) );
  AND3_X1 U5838 ( .A1(n6853), .A2(n6852), .A3(n6851), .ZN(n9806) );
  AND3_X1 U5839 ( .A1(n6550), .A2(n6549), .A3(n6548), .ZN(n9801) );
  OR2_X1 U5840 ( .A1(n6912), .A2(n6469), .ZN(n9831) );
  AND3_X1 U5841 ( .A1(n6466), .A2(n6473), .A3(n6905), .ZN(n6408) );
  INV_X1 U5842 ( .A(n9708), .ZN(n9721) );
  INV_X1 U5843 ( .A(n9731), .ZN(n9720) );
  INV_X1 U5844 ( .A(n9834), .ZN(n9717) );
  XNOR2_X1 U5845 ( .A(n5926), .B(n9786), .ZN(n5927) );
  NAND2_X1 U5846 ( .A1(n9788), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5926) );
  XNOR2_X1 U5847 ( .A(n5689), .B(n5688), .ZN(n8986) );
  NAND2_X1 U5848 ( .A1(n5382), .A2(n5381), .ZN(n5398) );
  NAND2_X1 U5849 ( .A1(n4959), .A2(n4961), .ZN(n5340) );
  NAND2_X1 U5850 ( .A1(n4960), .A2(n5308), .ZN(n4959) );
  INV_X1 U5851 ( .A(n5303), .ZN(n4960) );
  OR2_X1 U5852 ( .A1(n6025), .A2(n5854), .ZN(n6039) );
  INV_X1 U5853 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6024) );
  OR2_X1 U5854 ( .A1(n5156), .A2(SI_1_), .ZN(n5157) );
  NAND2_X1 U5855 ( .A1(n6433), .A2(n5941), .ZN(n5159) );
  NAND2_X1 U5856 ( .A1(n5800), .A2(n5799), .ZN(n6167) );
  NAND2_X1 U5857 ( .A1(n6585), .A2(n6584), .ZN(n6588) );
  NOR2_X1 U5858 ( .A1(n8310), .A2(n4917), .ZN(n4916) );
  INV_X1 U5859 ( .A(n8047), .ZN(n4917) );
  NAND2_X1 U5860 ( .A1(n4918), .A2(n8047), .ZN(n8309) );
  NAND2_X1 U5861 ( .A1(n8397), .A2(n8041), .ZN(n4943) );
  NAND2_X1 U5862 ( .A1(n4915), .A2(n6316), .ZN(n4912) );
  NAND2_X1 U5863 ( .A1(n8333), .A2(n8332), .ZN(n8331) );
  AND2_X1 U5864 ( .A1(n6632), .A2(n5716), .ZN(n8591) );
  AOI21_X1 U5865 ( .B1(n4947), .B2(n4945), .A(n4590), .ZN(n4944) );
  INV_X1 U5866 ( .A(n4947), .ZN(n4946) );
  INV_X1 U5867 ( .A(n8332), .ZN(n4945) );
  NAND2_X1 U5868 ( .A1(n5641), .A2(n5640), .ZN(n8830) );
  INV_X1 U5869 ( .A(n8764), .ZN(n8357) );
  NAND2_X1 U5870 ( .A1(n6308), .A2(n6307), .ZN(n6365) );
  NAND2_X1 U5871 ( .A1(n8397), .A2(n4939), .ZN(n4933) );
  NAND2_X1 U5872 ( .A1(n5623), .A2(n5622), .ZN(n8376) );
  INV_X1 U5873 ( .A(n8427), .ZN(n8406) );
  NAND2_X1 U5874 ( .A1(n8331), .A2(n8033), .ZN(n8379) );
  NAND2_X1 U5875 ( .A1(n7168), .A2(n7287), .ZN(n7286) );
  NAND2_X1 U5876 ( .A1(n6300), .A2(n6301), .ZN(n4914) );
  AOI21_X1 U5877 ( .B1(n4923), .B2(n4922), .A(n4920), .ZN(n6367) );
  AND2_X1 U5878 ( .A1(n6364), .A2(n5883), .ZN(n4922) );
  NAND2_X1 U5879 ( .A1(n6367), .A2(n6366), .ZN(n6585) );
  INV_X1 U5880 ( .A(n8439), .ZN(n6785) );
  AOI22_X1 U5881 ( .A1(n8318), .A2(n8319), .B1(n8024), .B2(n8023), .ZN(n8426)
         );
  INV_X1 U5882 ( .A(n8409), .ZN(n8431) );
  NAND2_X1 U5883 ( .A1(n5650), .A2(n5649), .ZN(n8613) );
  NAND2_X1 U5884 ( .A1(n5632), .A2(n5631), .ZN(n8650) );
  NAND2_X1 U5885 ( .A1(n5616), .A2(n5615), .ZN(n8838) );
  NAND2_X1 U5886 ( .A1(n5575), .A2(n5574), .ZN(n8856) );
  OAI21_X1 U5887 ( .B1(n9860), .B2(n6171), .A(n6172), .ZN(n9863) );
  AOI21_X1 U5888 ( .B1(n6255), .B2(n6254), .A(n6253), .ZN(n6273) );
  AOI21_X1 U5889 ( .B1(n6509), .B2(n6503), .A(n6502), .ZN(n6819) );
  NOR2_X1 U5890 ( .A1(n6807), .A2(n6971), .ZN(n6893) );
  NAND2_X1 U5891 ( .A1(n4895), .A2(n4897), .ZN(n9890) );
  INV_X1 U5892 ( .A(n8471), .ZN(n4848) );
  INV_X1 U5893 ( .A(n4673), .ZN(n9906) );
  INV_X1 U5894 ( .A(n4672), .ZN(n9925) );
  INV_X1 U5895 ( .A(n8511), .ZN(n4835) );
  NOR2_X1 U5896 ( .A1(n8477), .A2(n8476), .ZN(n8512) );
  OAI21_X1 U5897 ( .B1(n9961), .B2(n4604), .A(n8462), .ZN(n9970) );
  AND2_X1 U5898 ( .A1(n9962), .A2(n8519), .ZN(n4604) );
  INV_X1 U5899 ( .A(n7574), .ZN(n5718) );
  NAND2_X1 U5900 ( .A1(n5041), .A2(n4589), .ZN(n8577) );
  NAND2_X1 U5901 ( .A1(n5042), .A2(n10005), .ZN(n5041) );
  NAND2_X1 U5902 ( .A1(n5048), .A2(n5762), .ZN(n8601) );
  NAND2_X1 U5903 ( .A1(n5761), .A2(n4517), .ZN(n5048) );
  NAND2_X1 U5904 ( .A1(n5666), .A2(n5665), .ZN(n8631) );
  INV_X1 U5905 ( .A(n8856), .ZN(n8663) );
  NAND2_X1 U5906 ( .A1(n5589), .A2(n5588), .ZN(n8665) );
  NAND2_X1 U5907 ( .A1(n5565), .A2(n5564), .ZN(n8845) );
  NAND2_X1 U5908 ( .A1(n8703), .A2(n7723), .ZN(n8679) );
  NAND2_X1 U5909 ( .A1(n5540), .A2(n5539), .ZN(n8863) );
  NAND2_X1 U5910 ( .A1(n5520), .A2(n5519), .ZN(n8873) );
  INV_X1 U5911 ( .A(n8694), .ZN(n8876) );
  NAND2_X1 U5912 ( .A1(n5501), .A2(n5500), .ZN(n8733) );
  NAND2_X1 U5913 ( .A1(n5026), .A2(n5030), .ZN(n7152) );
  NAND2_X1 U5914 ( .A1(n6982), .A2(n5032), .ZN(n5026) );
  OAI21_X1 U5915 ( .B1(n6982), .B2(n4537), .A(n5736), .ZN(n7184) );
  NOR2_X1 U5916 ( .A1(n6423), .A2(n8778), .ZN(n8757) );
  NOR2_X1 U5917 ( .A1(n8802), .A2(n9979), .ZN(n8684) );
  NOR2_X1 U5918 ( .A1(n8802), .A2(n10025), .ZN(n8795) );
  NOR2_X1 U5919 ( .A1(n8802), .A2(n6764), .ZN(n8793) );
  NAND2_X1 U5920 ( .A1(n5914), .A2(n5913), .ZN(n8788) );
  INV_X1 U5921 ( .A(n7783), .ZN(n7582) );
  NAND2_X1 U5922 ( .A1(n5693), .A2(n5692), .ZN(n8898) );
  NAND2_X1 U5923 ( .A1(n5659), .A2(n5658), .ZN(n8907) );
  NAND2_X1 U5924 ( .A1(n4792), .A2(n4797), .ZN(n8610) );
  NAND2_X1 U5925 ( .A1(n8641), .A2(n4798), .ZN(n4792) );
  AOI21_X1 U5926 ( .B1(n8641), .B2(n5633), .A(n7586), .ZN(n8621) );
  INV_X1 U5927 ( .A(n8376), .ZN(n8916) );
  NAND2_X1 U5928 ( .A1(n5609), .A2(n5608), .ZN(n8922) );
  NAND2_X1 U5929 ( .A1(n5553), .A2(n5552), .ZN(n8937) );
  NAND2_X1 U5930 ( .A1(n4810), .A2(n5740), .ZN(n8723) );
  NAND2_X1 U5931 ( .A1(n5483), .A2(n5482), .ZN(n5741) );
  AND2_X1 U5932 ( .A1(n8742), .A2(n8741), .ZN(n8951) );
  NAND2_X1 U5933 ( .A1(n5460), .A2(n5459), .ZN(n8958) );
  NAND2_X1 U5934 ( .A1(n5019), .A2(n5020), .ZN(n8751) );
  NAND2_X1 U5935 ( .A1(n5737), .A2(n5022), .ZN(n5019) );
  NAND2_X1 U5936 ( .A1(n5737), .A2(n7588), .ZN(n8761) );
  INV_X1 U5937 ( .A(n8933), .ZN(n8970) );
  NAND2_X1 U5938 ( .A1(n7157), .A2(n7690), .ZN(n8771) );
  AND2_X1 U5939 ( .A1(n6166), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6083) );
  INV_X1 U5940 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8977) );
  INV_X1 U5941 ( .A(n5798), .ZN(n8993) );
  XNOR2_X1 U5942 ( .A(n5134), .B(n5141), .ZN(n7296) );
  INV_X1 U5943 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7215) );
  NAND2_X1 U5944 ( .A1(n5136), .A2(n4550), .ZN(n7618) );
  INV_X1 U5945 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6831) );
  INV_X1 U5946 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6601) );
  AND2_X1 U5947 ( .A1(n6433), .A2(P2_U3151), .ZN(n8988) );
  NAND2_X1 U5948 ( .A1(n9127), .A2(n9129), .ZN(n9006) );
  NAND2_X1 U5949 ( .A1(n4876), .A2(n4881), .ZN(n9098) );
  NAND2_X1 U5950 ( .A1(n7958), .A2(n4883), .ZN(n4876) );
  NAND2_X1 U5951 ( .A1(n4886), .A2(n6847), .ZN(n9068) );
  INV_X1 U5952 ( .A(n4887), .ZN(n4886) );
  NAND2_X1 U5953 ( .A1(n7438), .A2(n7437), .ZN(n7810) );
  NAND2_X1 U5954 ( .A1(n4875), .A2(n4874), .ZN(n6464) );
  OR2_X1 U5955 ( .A1(n6487), .A2(n5968), .ZN(n9159) );
  OR2_X1 U5956 ( .A1(n6487), .A2(n6663), .ZN(n9158) );
  NAND2_X1 U5957 ( .A1(n7487), .A2(n7486), .ZN(n9355) );
  NAND2_X1 U5958 ( .A1(n9088), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9157) );
  NAND2_X1 U5959 ( .A1(n7514), .A2(n7513), .ZN(n9711) );
  OAI21_X1 U5960 ( .B1(n4631), .B2(n8267), .A(n8266), .ZN(n4630) );
  AOI21_X1 U5961 ( .B1(n8269), .B2(n6477), .A(n8285), .ZN(n4628) );
  INV_X1 U5962 ( .A(n9341), .ZN(n9636) );
  INV_X1 U5963 ( .A(n9374), .ZN(n9649) );
  OR2_X1 U5964 ( .A1(n5958), .A2(n5859), .ZN(n9176) );
  NOR2_X1 U5965 ( .A1(n5993), .A2(n4657), .ZN(n6222) );
  AND2_X1 U5966 ( .A1(n6002), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4657) );
  INV_X1 U5967 ( .A(n4656), .ZN(n6220) );
  INV_X1 U5968 ( .A(n4724), .ZN(n6014) );
  NOR2_X1 U5969 ( .A1(n6000), .A2(n5999), .ZN(n6010) );
  AND2_X1 U5970 ( .A1(n4656), .A2(n4655), .ZN(n6000) );
  NAND2_X1 U5971 ( .A1(n6217), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4655) );
  INV_X1 U5972 ( .A(n4722), .ZN(n6028) );
  INV_X1 U5973 ( .A(n4654), .ZN(n6054) );
  INV_X1 U5974 ( .A(n4728), .ZN(n6060) );
  AND2_X1 U5975 ( .A1(n4654), .A2(n4653), .ZN(n6059) );
  NAND2_X1 U5976 ( .A1(n6061), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n4653) );
  INV_X1 U5977 ( .A(n4652), .ZN(n6194) );
  INV_X1 U5978 ( .A(n4726), .ZN(n6201) );
  NOR2_X1 U5979 ( .A1(n6521), .A2(n4730), .ZN(n6524) );
  AND2_X1 U5980 ( .A1(n7253), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4730) );
  NOR2_X1 U5981 ( .A1(n6524), .A2(n6523), .ZN(n6641) );
  NOR2_X1 U5982 ( .A1(n6525), .A2(n4658), .ZN(n6527) );
  AND2_X1 U5983 ( .A1(n7253), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4658) );
  NOR2_X1 U5984 ( .A1(n6527), .A2(n6526), .ZN(n6637) );
  NOR2_X1 U5985 ( .A1(n4659), .A2(n6637), .ZN(n6639) );
  AND2_X1 U5986 ( .A1(n7340), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4659) );
  NAND2_X1 U5987 ( .A1(n6639), .A2(n6638), .ZN(n6792) );
  NOR2_X1 U5988 ( .A1(n6959), .A2(n4738), .ZN(n6963) );
  AND2_X1 U5989 ( .A1(n7506), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4738) );
  NOR2_X1 U5990 ( .A1(n6963), .A2(n6962), .ZN(n9186) );
  NOR2_X1 U5991 ( .A1(n6956), .A2(n4661), .ZN(n6958) );
  AND2_X1 U5992 ( .A1(n7506), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n4661) );
  XNOR2_X1 U5993 ( .A(n9202), .B(n9201), .ZN(n9188) );
  NAND2_X1 U5994 ( .A1(n6107), .A2(n9793), .ZN(n9254) );
  NOR2_X1 U5995 ( .A1(n9193), .A2(n9194), .ZN(n9197) );
  NAND2_X1 U5996 ( .A1(n9197), .A2(n9196), .ZN(n9216) );
  AND2_X1 U5997 ( .A1(n9228), .A2(n9227), .ZN(n9232) );
  NAND2_X1 U5998 ( .A1(n9232), .A2(n9231), .ZN(n9249) );
  NAND2_X1 U5999 ( .A1(n9261), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4735) );
  INV_X1 U6000 ( .A(n9260), .ZN(n4734) );
  NAND2_X1 U6001 ( .A1(n9257), .A2(n4553), .ZN(n4647) );
  NAND2_X1 U6002 ( .A1(n4736), .A2(n9230), .ZN(n4732) );
  OAI22_X1 U6003 ( .A1(n9256), .A2(n9254), .B1(n4736), .B2(n9259), .ZN(n4649)
         );
  NOR2_X1 U6004 ( .A1(n7537), .A2(n9494), .ZN(n7545) );
  AND2_X1 U6005 ( .A1(n9325), .A2(n9324), .ZN(n9617) );
  NAND2_X1 U6006 ( .A1(n9368), .A2(n9303), .ZN(n9352) );
  NAND2_X1 U6007 ( .A1(n5098), .A2(n5099), .ZN(n9366) );
  NAND2_X1 U6008 ( .A1(n9397), .A2(n5102), .ZN(n5098) );
  OAI21_X1 U6009 ( .B1(n9397), .B2(n4534), .A(n5104), .ZN(n9380) );
  NAND2_X1 U6010 ( .A1(n9429), .A2(n9297), .ZN(n9416) );
  NAND2_X1 U6011 ( .A1(n5059), .A2(n5109), .ZN(n9414) );
  INV_X1 U6012 ( .A(n9405), .ZN(n9667) );
  NOR2_X1 U6013 ( .A1(n4752), .A2(n4751), .ZN(n5106) );
  INV_X1 U6014 ( .A(n9296), .ZN(n4751) );
  INV_X1 U6015 ( .A(n9453), .ZN(n4752) );
  NAND2_X1 U6016 ( .A1(n5079), .A2(n5083), .ZN(n9461) );
  NAND2_X1 U6017 ( .A1(n9493), .A2(n5084), .ZN(n5079) );
  AND2_X1 U6018 ( .A1(n5086), .A2(n5087), .ZN(n9477) );
  NAND2_X1 U6019 ( .A1(n9493), .A2(n9276), .ZN(n5086) );
  NAND2_X1 U6020 ( .A1(n9503), .A2(n8246), .ZN(n9475) );
  NAND2_X1 U6021 ( .A1(n9550), .A2(n8241), .ZN(n9535) );
  NOR2_X1 U6022 ( .A1(n9585), .A2(n9693), .ZN(n9548) );
  NOR2_X1 U6023 ( .A1(n4758), .A2(n4618), .ZN(n9551) );
  INV_X1 U6024 ( .A(n9578), .ZN(n4758) );
  NAND2_X1 U6025 ( .A1(n7382), .A2(n8236), .ZN(n9271) );
  NAND2_X1 U6026 ( .A1(n7381), .A2(n7380), .ZN(n7382) );
  NOR2_X1 U6027 ( .A1(n4742), .A2(n4741), .ZN(n7263) );
  NAND2_X1 U6028 ( .A1(n5070), .A2(n5073), .ZN(n7275) );
  NAND2_X1 U6029 ( .A1(n7088), .A2(n5075), .ZN(n5070) );
  AND2_X1 U6030 ( .A1(n7088), .A2(n7032), .ZN(n7236) );
  NAND2_X1 U6031 ( .A1(n4611), .A2(n6678), .ZN(n6735) );
  INV_X1 U6032 ( .A(n9538), .ZN(n9595) );
  INV_X1 U6033 ( .A(n9494), .ZN(n9593) );
  AND2_X1 U6034 ( .A1(n9598), .A2(n6910), .ZN(n9569) );
  NAND2_X1 U6035 ( .A1(n6401), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6402) );
  AND2_X1 U6036 ( .A1(n9598), .A2(n9720), .ZN(n9587) );
  INV_X2 U6037 ( .A(n9847), .ZN(n9850) );
  INV_X1 U6038 ( .A(n8105), .ZN(n8188) );
  INV_X1 U6039 ( .A(n9265), .ZN(n9746) );
  INV_X1 U6040 ( .A(n9612), .ZN(n4720) );
  INV_X1 U6041 ( .A(n9390), .ZN(n9763) );
  AND2_X1 U6042 ( .A1(n7511), .A2(n7510), .ZN(n9776) );
  INV_X2 U6043 ( .A(n9836), .ZN(n9838) );
  NAND2_X1 U6044 ( .A1(n8271), .A2(n6102), .ZN(n9797) );
  INV_X1 U6045 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9786) );
  XNOR2_X1 U6046 ( .A(n7472), .B(n7471), .ZN(n8976) );
  CLKBUF_X1 U6047 ( .A(n5967), .Z(n5968) );
  CLKBUF_X1 U6048 ( .A(n5966), .Z(n9793) );
  NAND2_X1 U6049 ( .A1(n5852), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U6050 ( .A1(n5852), .A2(n5851), .ZN(n9794) );
  XNOR2_X1 U6051 ( .A(n5853), .B(n10342), .ZN(n7452) );
  NAND2_X1 U6052 ( .A1(n4540), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5853) );
  INV_X1 U6053 ( .A(n5954), .ZN(n7298) );
  INV_X1 U6054 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10416) );
  INV_X1 U6055 ( .A(n8075), .ZN(n8267) );
  INV_X1 U6056 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10247) );
  NAND2_X1 U6057 ( .A1(n5844), .A2(n5069), .ZN(n5066) );
  INV_X1 U6058 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6599) );
  INV_X1 U6059 ( .A(n4693), .ZN(n5422) );
  AOI21_X1 U6060 ( .B1(n4692), .B2(n4697), .A(n4696), .ZN(n4693) );
  NAND2_X1 U6061 ( .A1(n4990), .A2(n4989), .ZN(n5417) );
  NAND2_X1 U6062 ( .A1(n4990), .A2(n4542), .ZN(n5401) );
  NAND2_X1 U6063 ( .A1(n4692), .A2(n4543), .ZN(n5367) );
  NAND2_X1 U6064 ( .A1(n5309), .A2(n5308), .ZN(n5324) );
  NAND2_X1 U6065 ( .A1(n5303), .A2(n5302), .ZN(n5309) );
  INV_X1 U6066 ( .A(n4953), .ZN(n4952) );
  XNOR2_X1 U6067 ( .A(n10141), .B(n4645), .ZN(n7572) );
  NAND2_X1 U6068 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4645) );
  INV_X1 U6069 ( .A(n4667), .ZN(n6881) );
  AOI21_X1 U6070 ( .B1(n4677), .B2(n9877), .A(n4674), .ZN(n8548) );
  NAND2_X1 U6071 ( .A1(n4676), .A2(n4675), .ZN(n4674) );
  XNOR2_X1 U6072 ( .A(n4830), .B(n4829), .ZN(n8574) );
  INV_X1 U6073 ( .A(n8563), .ZN(n4829) );
  INV_X1 U6074 ( .A(n5039), .ZN(n5834) );
  NAND2_X1 U6075 ( .A1(n10070), .A2(n5835), .ZN(n5038) );
  OAI211_X1 U6076 ( .C1(n8307), .C2(n8306), .A(n8305), .B(n4869), .ZN(P1_U3220) );
  NAND2_X1 U6077 ( .A1(n8307), .A2(n4870), .ZN(n4869) );
  NAND2_X1 U6078 ( .A1(n4648), .A2(n4646), .ZN(P1_U3262) );
  AOI21_X1 U6079 ( .B1(n4649), .B2(n9343), .A(n4733), .ZN(n4648) );
  NAND2_X1 U6080 ( .A1(n4647), .A2(n9327), .ZN(n4646) );
  NAND2_X1 U6081 ( .A1(n4735), .A2(n4734), .ZN(n4733) );
  NAND2_X1 U6082 ( .A1(n7485), .A2(n7484), .ZN(n8068) );
  INV_X1 U6083 ( .A(n7287), .ZN(n4932) );
  INV_X1 U6084 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5403) );
  AND2_X1 U6085 ( .A1(n4961), .A2(n4958), .ZN(n4515) );
  AND2_X1 U6086 ( .A1(n9430), .A2(n9296), .ZN(n4516) );
  AND2_X1 U6087 ( .A1(n5760), .A2(n4533), .ZN(n4517) );
  AND2_X1 U6088 ( .A1(n4747), .A2(n9302), .ZN(n4518) );
  INV_X1 U6089 ( .A(n7815), .ZN(n7816) );
  OR2_X1 U6090 ( .A1(n9689), .A2(n9505), .ZN(n4519) );
  OR3_X1 U6091 ( .A1(n6146), .A2(n6145), .A3(n6144), .ZN(n9658) );
  AND2_X1 U6092 ( .A1(n4718), .A2(n4717), .ZN(n4520) );
  NAND2_X1 U6093 ( .A1(n5687), .A2(n5686), .ZN(n8614) );
  INV_X1 U6094 ( .A(n8142), .ZN(n4621) );
  AND2_X1 U6095 ( .A1(n4817), .A2(n4814), .ZN(n4521) );
  INV_X1 U6096 ( .A(n5097), .ZN(n5096) );
  NAND2_X1 U6097 ( .A1(n4546), .A2(n5099), .ZN(n5097) );
  AND2_X1 U6098 ( .A1(n7718), .A2(n7708), .ZN(n7706) );
  INV_X1 U6099 ( .A(n7706), .ZN(n8725) );
  AND2_X1 U6100 ( .A1(n4801), .A2(n8614), .ZN(n4522) );
  NOR2_X1 U6101 ( .A1(n7422), .A2(n9817), .ZN(n4523) );
  AND2_X1 U6102 ( .A1(n9696), .A2(n9699), .ZN(n9275) );
  AND2_X1 U6103 ( .A1(n5357), .A2(n7670), .ZN(n4524) );
  AND2_X1 U6104 ( .A1(n6586), .A2(n6584), .ZN(n4525) );
  INV_X1 U6105 ( .A(n7667), .ZN(n7596) );
  AND2_X1 U6106 ( .A1(n6781), .A2(n7669), .ZN(n7667) );
  AND2_X1 U6107 ( .A1(n6341), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4526) );
  AND2_X1 U6108 ( .A1(n4854), .A2(n7815), .ZN(n4527) );
  NOR2_X1 U6109 ( .A1(n8073), .A2(n6672), .ZN(n4528) );
  OR2_X1 U6110 ( .A1(n6245), .A2(n6337), .ZN(n4529) );
  NAND2_X1 U6111 ( .A1(n4824), .A2(n6164), .ZN(n4530) );
  XNOR2_X1 U6112 ( .A(n5953), .B(P1_IR_REG_22__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U6113 ( .A1(n5972), .A2(n5837), .ZN(n5975) );
  OR2_X1 U6114 ( .A1(n4642), .A2(n4641), .ZN(n4531) );
  NAND2_X1 U6115 ( .A1(n9052), .A2(n4873), .ZN(n4872) );
  NAND2_X1 U6116 ( .A1(n8873), .A2(n8694), .ZN(n4532) );
  OR2_X1 U6117 ( .A1(n8907), .A2(n8631), .ZN(n4533) );
  NOR2_X1 U6118 ( .A1(n9408), .A2(n9658), .ZN(n4534) );
  OR2_X1 U6119 ( .A1(n5764), .A2(n5047), .ZN(n4535) );
  NAND2_X1 U6120 ( .A1(n5943), .A2(n5921), .ZN(n4536) );
  AND2_X1 U6121 ( .A1(n10059), .A2(n10041), .ZN(n4537) );
  NOR2_X1 U6122 ( .A1(n10030), .A2(n8439), .ZN(n4538) );
  AND2_X1 U6123 ( .A1(n7918), .A2(n7917), .ZN(n4539) );
  NAND2_X1 U6124 ( .A1(n5846), .A2(n5089), .ZN(n4540) );
  AOI21_X1 U6125 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n6289), .A(n6277), .ZN(
        n6241) );
  OR3_X1 U6126 ( .A1(n8162), .A2(n8155), .A3(n8277), .ZN(n4541) );
  NAND2_X1 U6127 ( .A1(n4933), .A2(n4938), .ZN(n8371) );
  OR2_X1 U6128 ( .A1(n5396), .A2(SI_11_), .ZN(n4542) );
  OR2_X1 U6129 ( .A1(n5359), .A2(SI_9_), .ZN(n4543) );
  INV_X1 U6130 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n10261) );
  XNOR2_X1 U6131 ( .A(n4943), .B(n8042), .ZN(n8325) );
  AND2_X1 U6132 ( .A1(n4672), .A2(n4671), .ZN(n4544) );
  OAI21_X1 U6133 ( .B1(n9063), .B2(n9061), .A(n9060), .ZN(n9081) );
  NAND2_X1 U6134 ( .A1(n8680), .A2(n5751), .ZN(n8675) );
  INV_X1 U6135 ( .A(n9297), .ZN(n4750) );
  NAND2_X1 U6136 ( .A1(n7489), .A2(n7488), .ZN(n9376) );
  OR2_X1 U6137 ( .A1(n8500), .A2(n8501), .ZN(n4545) );
  AND4_X1 U6138 ( .A1(n5335), .A2(n5334), .A3(n5333), .A4(n5332), .ZN(n10026)
         );
  OR2_X1 U6139 ( .A1(n9376), .A2(n9386), .ZN(n4546) );
  AND2_X1 U6140 ( .A1(n4665), .A2(n4664), .ZN(n4547) );
  AND3_X1 U6141 ( .A1(n7031), .A2(n7030), .A3(n7029), .ZN(n7260) );
  AND2_X1 U6142 ( .A1(n9376), .A2(n9386), .ZN(n4548) );
  AND2_X1 U6143 ( .A1(n7763), .A2(n4763), .ZN(n4549) );
  OR3_X1 U6144 ( .A1(n5137), .A2(P2_IR_REG_20__SCAN_IN), .A3(
        P2_IR_REG_21__SCAN_IN), .ZN(n4550) );
  AND2_X1 U6145 ( .A1(n7638), .A2(n7775), .ZN(n4551) );
  INV_X1 U6146 ( .A(n8181), .ZN(n4702) );
  AND2_X1 U6147 ( .A1(n8703), .A2(n4817), .ZN(n4552) );
  AND2_X1 U6148 ( .A1(n4732), .A2(n9258), .ZN(n4553) );
  AND2_X1 U6149 ( .A1(n9384), .A2(n9302), .ZN(n4554) );
  NAND2_X1 U6150 ( .A1(n5383), .A2(n5133), .ZN(n5137) );
  AND2_X1 U6151 ( .A1(n9689), .A2(n9505), .ZN(n4555) );
  AND2_X1 U6152 ( .A1(n9265), .A2(n8252), .ZN(n4556) );
  NOR2_X1 U6153 ( .A1(n7611), .A2(n7582), .ZN(n4557) );
  OR2_X1 U6154 ( .A1(n9696), .A2(n9685), .ZN(n8246) );
  INV_X1 U6155 ( .A(n8246), .ZN(n4761) );
  OR2_X1 U6156 ( .A1(n5137), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n4558) );
  NAND2_X1 U6157 ( .A1(n7523), .A2(n7522), .ZN(n9689) );
  NOR2_X1 U6158 ( .A1(n8538), .A2(n8537), .ZN(n4559) );
  NOR2_X1 U6159 ( .A1(n8512), .A2(n8513), .ZN(n4560) );
  AND2_X1 U6160 ( .A1(n8278), .A2(n4894), .ZN(n4561) );
  AND2_X1 U6161 ( .A1(n7759), .A2(n8600), .ZN(n4562) );
  AND2_X1 U6162 ( .A1(n8331), .A2(n4947), .ZN(n4563) );
  INV_X1 U6163 ( .A(n9528), .ZN(n9702) );
  NAND2_X1 U6164 ( .A1(n7517), .A2(n7516), .ZN(n9528) );
  AND2_X1 U6165 ( .A1(n7688), .A2(n8775), .ZN(n4564) );
  NAND3_X1 U6166 ( .A1(n5847), .A2(n10232), .A3(n5855), .ZN(n4565) );
  INV_X1 U6167 ( .A(n7449), .ZN(n9784) );
  NAND2_X1 U6168 ( .A1(n7342), .A2(n7341), .ZN(n7449) );
  AND2_X1 U6169 ( .A1(n8958), .A2(n8764), .ZN(n4566) );
  OR2_X1 U6170 ( .A1(n8907), .A2(n8827), .ZN(n7757) );
  AND4_X1 U6171 ( .A1(n7059), .A2(n7058), .A3(n7057), .A4(n7056), .ZN(n7428)
         );
  OR2_X1 U6172 ( .A1(n8845), .A2(n8663), .ZN(n7740) );
  NOR2_X1 U6173 ( .A1(n7688), .A2(n8775), .ZN(n4567) );
  OR2_X1 U6174 ( .A1(n8958), .A2(n8357), .ZN(n7703) );
  NOR2_X1 U6175 ( .A1(n9270), .A2(n9269), .ZN(n4568) );
  NAND2_X1 U6176 ( .A1(n7496), .A2(n7495), .ZN(n9408) );
  AND2_X1 U6177 ( .A1(n8076), .A2(n9016), .ZN(n4569) );
  INV_X1 U6178 ( .A(n6664), .ZN(n6917) );
  AND4_X1 U6179 ( .A1(n6372), .A2(n10283), .A3(n5843), .A4(n6190), .ZN(n4570)
         );
  AND2_X1 U6180 ( .A1(n8830), .A2(n8636), .ZN(n7755) );
  INV_X1 U6181 ( .A(n7755), .ZN(n4800) );
  AND2_X1 U6182 ( .A1(n5338), .A2(n10417), .ZN(n4571) );
  AND2_X1 U6183 ( .A1(n7428), .A2(n7274), .ZN(n4572) );
  AND2_X1 U6184 ( .A1(n7723), .A2(n7727), .ZN(n8700) );
  INV_X1 U6185 ( .A(n8700), .ZN(n4814) );
  INV_X1 U6186 ( .A(n4992), .ZN(n4991) );
  NAND2_X1 U6187 ( .A1(n4993), .A2(n5381), .ZN(n4992) );
  NAND2_X1 U6188 ( .A1(n9552), .A2(n8206), .ZN(n4573) );
  AND2_X1 U6189 ( .A1(n4845), .A2(n4526), .ZN(n4574) );
  NAND2_X1 U6190 ( .A1(n8145), .A2(n8205), .ZN(n4575) );
  AND2_X1 U6191 ( .A1(n7783), .A2(n7794), .ZN(n4576) );
  AND2_X1 U6192 ( .A1(n9307), .A2(n9306), .ZN(n8175) );
  OR2_X1 U6193 ( .A1(n8607), .A2(n8614), .ZN(n7622) );
  INV_X1 U6194 ( .A(n5085), .ZN(n5084) );
  NAND2_X1 U6195 ( .A1(n4519), .A2(n9276), .ZN(n5085) );
  OR2_X1 U6196 ( .A1(n9275), .A2(n4555), .ZN(n4577) );
  AND2_X1 U6197 ( .A1(n9880), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4578) );
  NOR2_X1 U6198 ( .A1(n4998), .A2(n5474), .ZN(n4579) );
  NAND2_X1 U6199 ( .A1(n9389), .A2(n4520), .ZN(n4719) );
  INV_X1 U6200 ( .A(n5751), .ZN(n5009) );
  NAND2_X1 U6201 ( .A1(n5247), .A2(SI_4_), .ZN(n5260) );
  AND2_X1 U6202 ( .A1(n4814), .A2(n5747), .ZN(n4580) );
  INV_X1 U6203 ( .A(n8068), .ZN(n9751) );
  NAND2_X1 U6204 ( .A1(n6363), .A2(n10011), .ZN(n4581) );
  NAND2_X1 U6205 ( .A1(n8183), .A2(n8277), .ZN(n4582) );
  AND2_X1 U6206 ( .A1(n10261), .A2(n5938), .ZN(n5091) );
  INV_X1 U6207 ( .A(n5091), .ZN(n5090) );
  NOR2_X1 U6208 ( .A1(n5035), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n4583) );
  INV_X1 U6209 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4911) );
  AND2_X1 U6210 ( .A1(n4682), .A2(n4681), .ZN(n4584) );
  NAND2_X1 U6211 ( .A1(n7528), .A2(n7527), .ZN(n9681) );
  INV_X1 U6212 ( .A(n9681), .ZN(n4711) );
  NAND2_X1 U6213 ( .A1(n5677), .A2(n5676), .ZN(n8607) );
  INV_X1 U6214 ( .A(n8607), .ZN(n4801) );
  NAND2_X1 U6215 ( .A1(n4889), .A2(n7306), .ZN(n7404) );
  NAND2_X1 U6216 ( .A1(n7298), .A2(n9327), .ZN(n8277) );
  NAND2_X1 U6217 ( .A1(n7536), .A2(n7535), .ZN(n9620) );
  INV_X1 U6218 ( .A(n9620), .ZN(n4717) );
  AND2_X1 U6219 ( .A1(n7286), .A2(n4929), .ZN(n4585) );
  INV_X1 U6220 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4965) );
  AND4_X1 U6221 ( .A1(n7377), .A2(n7376), .A3(n7375), .A4(n7374), .ZN(n9562)
         );
  INV_X1 U6222 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n4707) );
  INV_X1 U6223 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n4739) );
  INV_X1 U6224 ( .A(n6895), .ZN(n7140) );
  INV_X1 U6225 ( .A(n9367), .ZN(n4747) );
  AND2_X1 U6226 ( .A1(n5345), .A2(n5369), .ZN(n6892) );
  INV_X1 U6227 ( .A(n10041), .ZN(n7186) );
  OR2_X1 U6228 ( .A1(n9676), .A2(n9666), .ZN(n4586) );
  NAND2_X1 U6229 ( .A1(n5597), .A2(n5596), .ZN(n8846) );
  OR2_X1 U6230 ( .A1(n5741), .A2(n8726), .ZN(n5740) );
  NAND2_X1 U6231 ( .A1(n9536), .A2(n4714), .ZN(n4715) );
  AND2_X1 U6232 ( .A1(n5512), .A2(n5494), .ZN(n4587) );
  NOR2_X1 U6233 ( .A1(n9661), .A2(n9405), .ZN(n4588) );
  OR2_X1 U6234 ( .A1(n5776), .A2(n7793), .ZN(n4589) );
  NOR2_X1 U6235 ( .A1(n8035), .A2(n8862), .ZN(n4590) );
  NOR2_X1 U6236 ( .A1(n4711), .A2(n9686), .ZN(n4591) );
  NAND2_X1 U6237 ( .A1(n8043), .A2(n8826), .ZN(n4592) );
  NOR2_X1 U6238 ( .A1(n8042), .A2(n8838), .ZN(n4593) );
  AND2_X1 U6239 ( .A1(n4901), .A2(n4900), .ZN(n4594) );
  AND2_X1 U6240 ( .A1(n4849), .A2(n4848), .ZN(n4595) );
  AND2_X2 U6241 ( .A1(n5833), .A2(n5832), .ZN(n10070) );
  AND2_X1 U6242 ( .A1(n9905), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4596) );
  XNOR2_X1 U6243 ( .A(n4836), .B(n6882), .ZN(n6807) );
  INV_X1 U6244 ( .A(n9060), .ZN(n4868) );
  INV_X1 U6245 ( .A(n8240), .ZN(n4618) );
  NAND2_X1 U6246 ( .A1(n4923), .A2(n5883), .ZN(n6308) );
  NAND2_X1 U6247 ( .A1(n5336), .A2(n7670), .ZN(n6975) );
  NOR2_X1 U6248 ( .A1(n6893), .A2(n6894), .ZN(n4597) );
  NAND2_X1 U6249 ( .A1(n5996), .A2(n5839), .ZN(n6055) );
  OR2_X1 U6250 ( .A1(n6055), .A2(n5066), .ZN(n4598) );
  AND2_X1 U6251 ( .A1(n5707), .A2(n5706), .ZN(n4599) );
  AND2_X1 U6252 ( .A1(n6847), .A2(n6843), .ZN(n4600) );
  INV_X1 U6253 ( .A(n9275), .ZN(n5087) );
  AND2_X1 U6254 ( .A1(n6176), .A2(n8561), .ZN(n9877) );
  NAND2_X1 U6255 ( .A1(n4914), .A2(n5872), .ZN(n6315) );
  NAND2_X1 U6256 ( .A1(n5445), .A2(n5444), .ZN(n8964) );
  INV_X1 U6257 ( .A(n8964), .ZN(n5021) );
  NAND2_X1 U6258 ( .A1(n4844), .A2(n4843), .ZN(n4601) );
  INV_X1 U6259 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n10141) );
  INV_X1 U6260 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5837) );
  INV_X1 U6261 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5855) );
  INV_X1 U6262 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5848) );
  XNOR2_X1 U6263 ( .A(n5939), .B(n5938), .ZN(n6477) );
  INV_X1 U6264 ( .A(n5824), .ZN(n7782) );
  XNOR2_X1 U6265 ( .A(n5138), .B(P2_IR_REG_20__SCAN_IN), .ZN(n5824) );
  INV_X1 U6266 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n10513) );
  INV_X1 U6267 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n4644) );
  NOR2_X1 U6268 ( .A1(n8504), .A2(n8884), .ZN(n8538) );
  OR2_X1 U6269 ( .A1(n7132), .A2(n5387), .ZN(n4901) );
  OAI21_X1 U6270 ( .B1(n8504), .B2(n4903), .A(n4902), .ZN(n9941) );
  INV_X1 U6271 ( .A(n8536), .ZN(n4834) );
  NAND2_X1 U6272 ( .A1(n7047), .A2(n8108), .ZN(n7071) );
  NAND2_X1 U6273 ( .A1(n4637), .A2(n4582), .ZN(n4636) );
  OAI21_X1 U6274 ( .B1(n8148), .B2(n8277), .A(n8203), .ZN(n4641) );
  INV_X1 U6275 ( .A(n8180), .ZN(n4640) );
  OAI21_X1 U6276 ( .B1(n8168), .B2(n8167), .A(n4624), .ZN(n4623) );
  AOI21_X1 U6277 ( .B1(n8274), .B2(n9327), .A(n8194), .ZN(n4631) );
  OAI211_X1 U6278 ( .C1(n8114), .C2(n8277), .A(n8116), .B(n4632), .ZN(n8120)
         );
  NAND2_X1 U6279 ( .A1(n4630), .A2(n8268), .ZN(n4629) );
  NAND2_X1 U6280 ( .A1(n4629), .A2(n4628), .ZN(n4627) );
  NAND3_X1 U6281 ( .A1(n5383), .A2(n5133), .A3(n4583), .ZN(n5778) );
  NAND2_X1 U6282 ( .A1(n7711), .A2(n7710), .ZN(n7724) );
  AOI21_X1 U6283 ( .B1(n7739), .B2(n8656), .A(n7738), .ZN(n7745) );
  NAND2_X1 U6284 ( .A1(n4768), .A2(n4767), .ZN(n4766) );
  OAI21_X1 U6285 ( .B1(n7712), .B2(n4784), .A(n7705), .ZN(n7707) );
  NAND2_X1 U6286 ( .A1(n7781), .A2(n7780), .ZN(n4781) );
  NOR2_X1 U6287 ( .A1(n7729), .A2(n4772), .ZN(n7731) );
  AOI21_X2 U6288 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n9956), .A(n9943), .ZN(
        n8515) );
  OR2_X1 U6289 ( .A1(n5793), .A2(P2_D_REG_0__SCAN_IN), .ZN(n5792) );
  OAI21_X1 U6290 ( .B1(n8030), .B2(n8740), .A(n8361), .ZN(n8404) );
  NAND2_X1 U6291 ( .A1(n6605), .A2(n6604), .ZN(n6653) );
  OAI22_X1 U6292 ( .A1(n8346), .A2(n8347), .B1(n8045), .B2(n8613), .ZN(n8413)
         );
  NAND2_X2 U6293 ( .A1(n6946), .A2(n6945), .ZN(n4607) );
  AOI21_X2 U6294 ( .B1(n7165), .B2(n7164), .A(n4606), .ZN(n7168) );
  XNOR2_X2 U6295 ( .A(n4607), .B(n7186), .ZN(n7165) );
  OAI21_X2 U6296 ( .B1(n6653), .B2(n6652), .A(n6651), .ZN(n6655) );
  NAND2_X1 U6297 ( .A1(n5261), .A2(n5260), .ZN(n5267) );
  NAND2_X2 U6298 ( .A1(n8399), .A2(n8398), .ZN(n8397) );
  NAND2_X1 U6299 ( .A1(n6364), .A2(n4921), .ZN(n4919) );
  OAI211_X2 U6300 ( .C1(n5861), .C2(n6261), .A(n5270), .B(n5269), .ZN(n6427)
         );
  INV_X1 U6301 ( .A(n6678), .ZN(n4609) );
  AOI21_X2 U6302 ( .B1(n4609), .B2(n8210), .A(n4569), .ZN(n4608) );
  NAND2_X1 U6303 ( .A1(n4612), .A2(n4613), .ZN(n8146) );
  NAND2_X1 U6304 ( .A1(n8144), .A2(n4614), .ZN(n4612) );
  INV_X1 U6305 ( .A(n5846), .ZN(n5951) );
  NAND2_X1 U6306 ( .A1(n5846), .A2(n5091), .ZN(n4626) );
  NAND3_X1 U6307 ( .A1(n8283), .A2(n8284), .A3(n4627), .ZN(P1_U3242) );
  NAND3_X1 U6308 ( .A1(n4640), .A2(n8174), .A3(n4638), .ZN(n4637) );
  OR2_X1 U6309 ( .A1(n6544), .A2(n6443), .ZN(n6446) );
  NAND2_X2 U6310 ( .A1(n5967), .A2(n5966), .ZN(n7229) );
  XNOR2_X1 U6311 ( .A(n5950), .B(P1_IR_REG_27__SCAN_IN), .ZN(n5966) );
  NOR2_X2 U6312 ( .A1(n6244), .A2(n4662), .ZN(n6181) );
  NOR2_X2 U6313 ( .A1(n8455), .A2(n4668), .ZN(n6507) );
  AND2_X2 U6314 ( .A1(n4669), .A2(n6816), .ZN(n8455) );
  OR2_X2 U6315 ( .A1(n9907), .A2(n9908), .ZN(n4673) );
  NAND3_X1 U6316 ( .A1(n4688), .A2(n8184), .A3(n4687), .ZN(n8254) );
  NAND2_X1 U6317 ( .A1(n5361), .A2(n5360), .ZN(n4692) );
  NAND3_X1 U6318 ( .A1(n8067), .A2(n8064), .A3(n8198), .ZN(n4704) );
  INV_X4 U6319 ( .A(n5158), .ZN(n6433) );
  NAND3_X1 U6320 ( .A1(n4523), .A2(n4708), .A3(n7098), .ZN(n4709) );
  INV_X1 U6321 ( .A(n4715), .ZN(n9478) );
  NAND2_X2 U6322 ( .A1(n9389), .A2(n4716), .ZN(n9326) );
  INV_X1 U6323 ( .A(n4719), .ZN(n9334) );
  NAND3_X1 U6324 ( .A1(n9613), .A2(n9611), .A3(n4720), .ZN(n9747) );
  NAND2_X1 U6325 ( .A1(n7262), .A2(n4740), .ZN(n7364) );
  INV_X1 U6326 ( .A(n8084), .ZN(n4741) );
  INV_X1 U6327 ( .A(n7262), .ZN(n4742) );
  OAI21_X2 U6328 ( .B1(n9384), .B2(n4746), .A(n4744), .ZN(n9350) );
  NAND2_X1 U6329 ( .A1(n4754), .A2(n4753), .ZN(P1_U3551) );
  OR2_X1 U6330 ( .A1(n9850), .A2(n6237), .ZN(n4753) );
  NAND2_X1 U6331 ( .A1(n9747), .A2(n9850), .ZN(n4754) );
  OAI22_X1 U6332 ( .A1(n9312), .A2(n9693), .B1(n9311), .B2(n9310), .ZN(n9612)
         );
  INV_X1 U6333 ( .A(n9474), .ZN(n8247) );
  AND2_X2 U6334 ( .A1(n4570), .A2(n4884), .ZN(n5844) );
  INV_X1 U6335 ( .A(n8611), .ZN(n4767) );
  OAI21_X1 U6336 ( .B1(n4771), .B2(n4770), .A(n4769), .ZN(n4768) );
  INV_X1 U6337 ( .A(n7756), .ZN(n4769) );
  NAND3_X1 U6338 ( .A1(n7658), .A2(n7637), .A3(n7768), .ZN(n4782) );
  AND2_X1 U6339 ( .A1(n7702), .A2(n8748), .ZN(n7712) );
  AND2_X1 U6340 ( .A1(n7745), .A2(n4785), .ZN(n7751) );
  NAND3_X1 U6341 ( .A1(n7743), .A2(n8640), .A3(n7742), .ZN(n4787) );
  NAND2_X1 U6342 ( .A1(n8641), .A2(n4790), .ZN(n4789) );
  OAI21_X1 U6343 ( .B1(n8641), .B2(n4796), .A(n4793), .ZN(n8599) );
  NAND2_X1 U6344 ( .A1(n7153), .A2(n4804), .ZN(n4802) );
  NAND2_X1 U6345 ( .A1(n4802), .A2(n4803), .ZN(n8760) );
  OAI21_X2 U6346 ( .B1(n7585), .B2(n7584), .A(n4808), .ZN(n4807) );
  NAND2_X1 U6347 ( .A1(n4810), .A2(n4809), .ZN(n8721) );
  NAND2_X1 U6348 ( .A1(n8701), .A2(n4813), .ZN(n4811) );
  NAND2_X1 U6349 ( .A1(n4811), .A2(n4812), .ZN(n8657) );
  NAND2_X1 U6350 ( .A1(n8701), .A2(n8700), .ZN(n8703) );
  NAND2_X1 U6351 ( .A1(n5336), .A2(n4524), .ZN(n6974) );
  NAND2_X1 U6352 ( .A1(n6974), .A2(n7655), .ZN(n6981) );
  NAND2_X2 U6353 ( .A1(n7629), .A2(n7633), .ZN(n8799) );
  NAND2_X2 U6354 ( .A1(n5005), .A2(n5868), .ZN(n7629) );
  NAND2_X1 U6355 ( .A1(n4819), .A2(n4825), .ZN(n4824) );
  INV_X1 U6356 ( .A(n9882), .ZN(n4819) );
  NAND2_X1 U6357 ( .A1(n9882), .A2(n6255), .ZN(n4820) );
  NAND2_X1 U6358 ( .A1(n6255), .A2(n4822), .ZN(n4821) );
  INV_X1 U6359 ( .A(n4825), .ZN(n4822) );
  NAND2_X1 U6360 ( .A1(n6164), .A2(n4825), .ZN(n4823) );
  NAND2_X1 U6361 ( .A1(n9880), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4825) );
  NOR2_X1 U6362 ( .A1(n9961), .A2(n8516), .ZN(n8518) );
  INV_X1 U6363 ( .A(n9944), .ZN(n4833) );
  INV_X1 U6364 ( .A(n6891), .ZN(n4836) );
  NAND2_X1 U6365 ( .A1(n6342), .A2(n6341), .ZN(n4844) );
  NAND2_X1 U6366 ( .A1(n6242), .A2(n4845), .ZN(n6243) );
  NOR2_X1 U6367 ( .A1(n9863), .A2(n8803), .ZN(n9862) );
  NAND2_X1 U6368 ( .A1(n5322), .A2(n7667), .ZN(n6993) );
  NAND2_X1 U6369 ( .A1(n5256), .A2(n7645), .ZN(n6413) );
  NAND2_X1 U6370 ( .A1(n5210), .A2(n7637), .ZN(n6922) );
  NOR2_X1 U6371 ( .A1(n7766), .A2(n7574), .ZN(n7585) );
  INV_X1 U6372 ( .A(n5528), .ZN(n8714) );
  NAND2_X1 U6373 ( .A1(n5702), .A2(n5701), .ZN(n7574) );
  NAND2_X1 U6374 ( .A1(n7593), .A2(n5192), .ZN(n8785) );
  NAND3_X2 U6375 ( .A1(n5219), .A2(n4910), .A3(n4908), .ZN(n9880) );
  NAND2_X1 U6376 ( .A1(n7438), .A2(n4851), .ZN(n4854) );
  INV_X1 U6377 ( .A(n4855), .ZN(n9035) );
  NAND3_X1 U6378 ( .A1(n4875), .A2(n6463), .A3(n4874), .ZN(n6532) );
  OAI21_X1 U6379 ( .B1(n7958), .B2(n4880), .A(n4877), .ZN(n9095) );
  NAND3_X1 U6380 ( .A1(n5842), .A2(n5841), .A3(n6056), .ZN(n4885) );
  NAND2_X1 U6381 ( .A1(n7106), .A2(n7105), .ZN(n7108) );
  NAND2_X1 U6382 ( .A1(n4889), .A2(n4888), .ZN(n7417) );
  NAND2_X1 U6383 ( .A1(n9115), .A2(n7832), .ZN(n7844) );
  INV_X2 U6384 ( .A(n4892), .ZN(n7883) );
  NAND2_X4 U6385 ( .A1(n4893), .A2(n5958), .ZN(n7998) );
  NOR2_X2 U6386 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5153) );
  XNOR2_X1 U6387 ( .A(n6245), .B(n6261), .ZN(n6246) );
  INV_X1 U6388 ( .A(n4901), .ZN(n8497) );
  NAND2_X1 U6389 ( .A1(n9905), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4899) );
  INV_X1 U6390 ( .A(n8498), .ZN(n4900) );
  NOR2_X1 U6391 ( .A1(n9959), .A2(n9960), .ZN(n9958) );
  NAND2_X1 U6392 ( .A1(n8543), .A2(n4907), .ZN(n4905) );
  NAND2_X1 U6393 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4909) );
  NAND2_X1 U6394 ( .A1(n5403), .A2(n4911), .ZN(n4910) );
  INV_X2 U6395 ( .A(n5874), .ZN(n8048) );
  OAI211_X2 U6396 ( .C1(n5864), .C2(n5865), .A(n5866), .B(n5867), .ZN(n5874)
         );
  NAND3_X1 U6397 ( .A1(n6300), .A2(n6316), .A3(n6301), .ZN(n4913) );
  NAND3_X1 U6398 ( .A1(n4913), .A2(n5877), .A3(n4912), .ZN(n6292) );
  NAND2_X1 U6399 ( .A1(n4918), .A2(n4916), .ZN(n8311) );
  NAND2_X1 U6400 ( .A1(n4581), .A2(n4919), .ZN(n4920) );
  NAND2_X1 U6401 ( .A1(n6585), .A2(n4525), .ZN(n6605) );
  NAND2_X1 U6402 ( .A1(n4924), .A2(n4925), .ZN(n8386) );
  NAND2_X1 U6403 ( .A1(n7168), .A2(n4927), .ZN(n4924) );
  NAND2_X1 U6404 ( .A1(n7286), .A2(n4931), .ZN(n7288) );
  AOI21_X2 U6405 ( .B1(n8397), .B2(n4935), .A(n4934), .ZN(n8346) );
  OAI21_X1 U6406 ( .B1(n8333), .B2(n4946), .A(n4944), .ZN(n8340) );
  NAND4_X1 U6407 ( .A1(n5120), .A2(n5119), .A3(n5118), .A4(n5258), .ZN(n4951)
         );
  OAI21_X1 U6408 ( .B1(n5251), .B2(n4954), .A(n5266), .ZN(n4953) );
  INV_X1 U6409 ( .A(n5260), .ZN(n4954) );
  OAI21_X1 U6410 ( .B1(n5252), .B2(n4954), .A(n4952), .ZN(n5286) );
  NAND2_X1 U6411 ( .A1(n5252), .A2(n5251), .ZN(n5261) );
  OAI21_X1 U6412 ( .B1(n5158), .B2(n4965), .A(n4964), .ZN(n5156) );
  NAND2_X1 U6413 ( .A1(n5158), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4964) );
  NAND2_X1 U6414 ( .A1(n4966), .A2(n4967), .ZN(n5652) );
  NAND2_X1 U6415 ( .A1(n5606), .A2(n4969), .ZN(n4966) );
  NAND2_X1 U6416 ( .A1(n5618), .A2(n5617), .ZN(n5635) );
  NAND2_X1 U6417 ( .A1(n4972), .A2(n4973), .ZN(n5579) );
  NAND2_X1 U6418 ( .A1(n5549), .A2(n4975), .ZN(n4972) );
  NAND2_X1 U6419 ( .A1(n5689), .A2(n4983), .ZN(n4981) );
  NAND2_X1 U6420 ( .A1(n5436), .A2(n4999), .ZN(n4997) );
  NAND2_X1 U6421 ( .A1(n4997), .A2(n4579), .ZN(n5472) );
  NAND4_X4 U6422 ( .A1(n5179), .A2(n5181), .A3(n5178), .A4(n5180), .ZN(n5870)
         );
  INV_X1 U6423 ( .A(n5870), .ZN(n5005) );
  NAND2_X1 U6424 ( .A1(n5006), .A2(n5007), .ZN(n5753) );
  NAND2_X1 U6425 ( .A1(n8682), .A2(n5751), .ZN(n5006) );
  NAND2_X1 U6426 ( .A1(n5011), .A2(n5012), .ZN(n5743) );
  NAND2_X1 U6427 ( .A1(n5737), .A2(n5014), .ZN(n5011) );
  NAND2_X1 U6428 ( .A1(n6982), .A2(n5027), .ZN(n5025) );
  NAND2_X1 U6429 ( .A1(n5037), .A2(n4580), .ZN(n8693) );
  NAND2_X1 U6430 ( .A1(n5761), .A2(n5760), .ZN(n8612) );
  NAND2_X1 U6431 ( .A1(n5143), .A2(n5142), .ZN(n5786) );
  NAND2_X1 U6432 ( .A1(n5143), .A2(n5051), .ZN(n5167) );
  INV_X1 U6433 ( .A(n6968), .ZN(n5733) );
  OR2_X2 U6434 ( .A1(n6546), .A2(n4965), .ZN(n5055) );
  NAND2_X2 U6435 ( .A1(n7229), .A2(n7468), .ZN(n6546) );
  NAND3_X1 U6436 ( .A1(n5991), .A2(n5972), .A3(n5837), .ZN(n5994) );
  NAND2_X1 U6437 ( .A1(n5059), .A2(n5057), .ZN(n9284) );
  NAND2_X1 U6438 ( .A1(n7343), .A2(n5061), .ZN(n5060) );
  OAI21_X1 U6439 ( .B1(n7088), .B2(n5072), .A(n5071), .ZN(n7277) );
  OAI21_X1 U6440 ( .B1(n7088), .B2(n7235), .A(n5075), .ZN(n7238) );
  NAND2_X1 U6441 ( .A1(n9493), .A2(n5080), .ZN(n5078) );
  NAND2_X1 U6442 ( .A1(n5846), .A2(n5088), .ZN(n5922) );
  NAND2_X1 U6443 ( .A1(n9397), .A2(n5094), .ZN(n5093) );
  OAI21_X1 U6444 ( .B1(n9397), .B2(n5097), .A(n5094), .ZN(n9349) );
  NAND2_X1 U6445 ( .A1(n5093), .A2(n5092), .ZN(n9288) );
  AOI21_X1 U6446 ( .B1(n5094), .B2(n5097), .A(n9351), .ZN(n5092) );
  NAND2_X1 U6447 ( .A1(n6532), .A2(n6531), .ZN(n9013) );
  OAI21_X1 U6448 ( .B1(n9318), .B2(n9317), .A(n9307), .ZN(n9309) );
  INV_X1 U6449 ( .A(n5200), .ZN(n5198) );
  INV_X1 U6450 ( .A(n8799), .ZN(n7593) );
  INV_X1 U6451 ( .A(n5927), .ZN(n5929) );
  NAND2_X1 U6452 ( .A1(n5922), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5946) );
  AOI22_X2 U6453 ( .A1(n8404), .A2(n8405), .B1(n8876), .B2(n8031), .ZN(n8333)
         );
  AND2_X1 U6454 ( .A1(n9676), .A2(n9666), .ZN(n5105) );
  INV_X1 U6455 ( .A(n8681), .ZN(n5750) );
  NAND2_X2 U6456 ( .A1(n6909), .A2(n9557), .ZN(n9598) );
  INV_X1 U6457 ( .A(n8541), .ZN(n9976) );
  INV_X1 U6458 ( .A(n9505), .ZN(n9277) );
  INV_X1 U6459 ( .A(P2_U3893), .ZN(n8531) );
  OR2_X1 U6460 ( .A1(n5493), .A2(SI_16_), .ZN(n5107) );
  INV_X1 U6461 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7494) );
  NAND2_X1 U6462 ( .A1(n8799), .A2(n8800), .ZN(n8798) );
  OR2_X1 U6463 ( .A1(n9751), .A2(n9607), .ZN(n5108) );
  OR2_X1 U6464 ( .A1(n9281), .A2(n9280), .ZN(n5109) );
  NOR2_X1 U6465 ( .A1(n5968), .A2(n9793), .ZN(n5110) );
  INV_X1 U6466 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7335) );
  INV_X1 U6467 ( .A(SI_18_), .ZN(n5514) );
  INV_X1 U6468 ( .A(n9666), .ZN(n9437) );
  INV_X1 U6469 ( .A(n8737), .ZN(n7704) );
  INV_X1 U6470 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5195) );
  AOI21_X1 U6471 ( .B1(n7580), .B2(n7579), .A(n7578), .ZN(n8809) );
  INV_X1 U6472 ( .A(n9272), .ZN(n9779) );
  AND3_X1 U6473 ( .A1(n6126), .A2(n6125), .A3(n6124), .ZN(n8252) );
  OR2_X1 U6474 ( .A1(n7619), .A2(n8933), .ZN(n5111) );
  NAND2_X1 U6475 ( .A1(n7811), .A2(n7812), .ZN(n5112) );
  OR2_X1 U6476 ( .A1(n5190), .A2(n9860), .ZN(n5113) );
  AND3_X2 U6477 ( .A1(n5818), .A2(n6420), .A3(n6422), .ZN(n10087) );
  AND2_X1 U6478 ( .A1(n5578), .A2(SI_21_), .ZN(n5114) );
  OR2_X1 U6479 ( .A1(n5578), .A2(SI_21_), .ZN(n5115) );
  INV_X1 U6480 ( .A(n9431), .ZN(n9281) );
  INV_X1 U6481 ( .A(n9817), .ZN(n7274) );
  OR2_X1 U6482 ( .A1(n10045), .A2(n8438), .ZN(n5116) );
  NAND2_X1 U6483 ( .A1(n7709), .A2(n7775), .ZN(n7710) );
  OAI21_X1 U6484 ( .B1(n7751), .B2(n7748), .A(n7747), .ZN(n7753) );
  NAND2_X1 U6485 ( .A1(n8196), .A2(n8197), .ZN(n8181) );
  INV_X1 U6486 ( .A(n8809), .ZN(n7581) );
  NOR4_X1 U6487 ( .A1(n7776), .A2(n7775), .A3(n7774), .A4(n7773), .ZN(n7777)
         );
  NAND2_X1 U6488 ( .A1(n7772), .A2(n7771), .ZN(n7781) );
  AND2_X1 U6489 ( .A1(n9956), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8540) );
  NAND2_X1 U6490 ( .A1(n8798), .A2(n5722), .ZN(n6774) );
  NOR3_X1 U6491 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .A3(
        P2_IR_REG_24__SCAN_IN), .ZN(n5142) );
  NOR2_X1 U6492 ( .A1(n8260), .A2(n6470), .ZN(n8261) );
  INV_X1 U6493 ( .A(SI_22_), .ZN(n10260) );
  INV_X1 U6494 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U6495 ( .A1(n8040), .A2(n8846), .ZN(n8041) );
  INV_X1 U6496 ( .A(n5568), .ZN(n5567) );
  INV_X1 U6497 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5145) );
  NAND2_X1 U6498 ( .A1(n7621), .A2(n8602), .ZN(n5701) );
  NAND2_X1 U6499 ( .A1(n5778), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U6500 ( .A1(n9023), .A2(n9138), .ZN(n7917) );
  OAI21_X1 U6501 ( .B1(n8262), .B2(n8273), .A(n8261), .ZN(n8263) );
  INV_X1 U6502 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7039) );
  INV_X1 U6503 ( .A(n9657), .ZN(n9280) );
  INV_X1 U6504 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5948) );
  INV_X1 U6505 ( .A(SI_27_), .ZN(n10406) );
  INV_X1 U6506 ( .A(SI_24_), .ZN(n10293) );
  INV_X1 U6507 ( .A(SI_17_), .ZN(n10434) );
  INV_X1 U6508 ( .A(n8763), .ZN(n8021) );
  NAND2_X1 U6509 ( .A1(n5567), .A2(n5566), .ZN(n5590) );
  OR2_X1 U6510 ( .A1(n5212), .A2(n5183), .ZN(n5184) );
  NAND2_X1 U6511 ( .A1(n5190), .A2(n7468), .ZN(n5222) );
  OR2_X1 U6512 ( .A1(n5812), .A2(n5866), .ZN(n5906) );
  INV_X1 U6513 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5129) );
  INV_X1 U6514 ( .A(n9087), .ZN(n9085) );
  AND2_X1 U6515 ( .A1(n9096), .A2(n9097), .ZN(n7972) );
  OR2_X1 U6516 ( .A1(n7945), .A2(n9131), .ZN(n7947) );
  OR2_X1 U6517 ( .A1(n7040), .A2(n7039), .ZN(n7054) );
  NOR2_X1 U6518 ( .A1(n9610), .A2(n9609), .ZN(n9611) );
  INV_X1 U6519 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5924) );
  INV_X1 U6520 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5938) );
  INV_X1 U6521 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6372) );
  OR2_X1 U6522 ( .A1(n6086), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n6116) );
  OAI21_X1 U6523 ( .B1(n6433), .B2(P1_DATAO_REG_0__SCAN_IN), .A(n5159), .ZN(
        n5160) );
  OR2_X1 U6524 ( .A1(n8032), .A2(n8869), .ZN(n8033) );
  INV_X1 U6525 ( .A(n5894), .ZN(n5888) );
  AND2_X1 U6526 ( .A1(n6632), .A2(n6631), .ZN(n7794) );
  INV_X1 U6527 ( .A(n8631), .ZN(n8827) );
  OR2_X1 U6528 ( .A1(n5610), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5625) );
  INV_X1 U6529 ( .A(n8740), .ZN(n8868) );
  INV_X1 U6530 ( .A(n6920), .ZN(n7592) );
  OR2_X1 U6531 ( .A1(n10087), .A2(n5819), .ZN(n5820) );
  OR2_X1 U6532 ( .A1(n5827), .A2(n5815), .ZN(n5816) );
  OR2_X1 U6533 ( .A1(n5864), .A2(n5827), .ZN(n5897) );
  INV_X1 U6534 ( .A(n8437), .ZN(n7321) );
  INV_X1 U6535 ( .A(n8438), .ZN(n6947) );
  AND2_X1 U6536 ( .A1(n5768), .A2(n5767), .ZN(n9979) );
  INV_X1 U6537 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U6538 ( .A1(n7929), .A2(n7930), .ZN(n7931) );
  OR2_X1 U6539 ( .A1(n7960), .A2(n9101), .ZN(n7976) );
  INV_X1 U6540 ( .A(n9658), .ZN(n9285) );
  INV_X1 U6541 ( .A(n5968), .ZN(n6663) );
  OR2_X1 U6542 ( .A1(n9731), .A2(n7539), .ZN(n9310) );
  INV_X1 U6543 ( .A(n9304), .ZN(n9351) );
  INV_X1 U6544 ( .A(n9676), .ZN(n9448) );
  INV_X1 U6545 ( .A(n8077), .ZN(n6707) );
  NAND2_X1 U6546 ( .A1(n8986), .A2(n7533), .ZN(n7536) );
  INV_X1 U6547 ( .A(n7229), .ZN(n7525) );
  OR2_X1 U6548 ( .A1(n8277), .A2(n8268), .ZN(n9737) );
  OR2_X1 U6549 ( .A1(n9494), .A2(n9343), .ZN(n6473) );
  NAND2_X1 U6550 ( .A1(n5925), .A2(n5924), .ZN(n9788) );
  NAND2_X1 U6551 ( .A1(n5857), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5858) );
  AND2_X1 U6552 ( .A1(n5798), .A2(n5797), .ZN(n5799) );
  INV_X1 U6553 ( .A(n8838), .ZN(n8637) );
  NAND2_X1 U6554 ( .A1(n5910), .A2(n5908), .ZN(n8409) );
  INV_X1 U6555 ( .A(n8428), .ZN(n8415) );
  INV_X1 U6556 ( .A(n8421), .ZN(n8423) );
  OR2_X1 U6557 ( .A1(n5211), .A2(n5205), .ZN(n5207) );
  INV_X1 U6558 ( .A(n8566), .ZN(n9967) );
  INV_X1 U6559 ( .A(n9888), .ZN(n9957) );
  OR2_X1 U6560 ( .A1(n6422), .A2(n6421), .ZN(n6423) );
  CLKBUF_X1 U6561 ( .A(n8757), .Z(n8745) );
  OAI21_X1 U6562 ( .B1(n7619), .B2(n8853), .A(n5820), .ZN(n5821) );
  INV_X1 U6563 ( .A(n8853), .ZN(n8890) );
  NAND2_X1 U6564 ( .A1(n5817), .A2(n5816), .ZN(n6422) );
  INV_X1 U6565 ( .A(n8622), .ZN(n8620) );
  INV_X1 U6566 ( .A(n10060), .ZN(n10062) );
  AND2_X1 U6567 ( .A1(n7698), .A2(n7699), .ZN(n8762) );
  NAND2_X1 U6568 ( .A1(n9988), .A2(n10055), .ZN(n10019) );
  INV_X1 U6569 ( .A(n9979), .ZN(n10005) );
  OR2_X1 U6570 ( .A1(n5907), .A2(n5831), .ZN(n5832) );
  INV_X1 U6571 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5405) );
  INV_X1 U6572 ( .A(n6477), .ZN(n8268) );
  AND2_X1 U6573 ( .A1(n9294), .A2(n6358), .ZN(n9328) );
  AND4_X1 U6574 ( .A1(n7951), .A2(n7950), .A3(n7949), .A4(n7948), .ZN(n9405)
         );
  AND4_X1 U6575 ( .A1(n7882), .A2(n7881), .A3(n7880), .A4(n7879), .ZN(n9685)
         );
  OR2_X1 U6576 ( .A1(n6480), .A2(P1_U3086), .ZN(n5859) );
  AND2_X1 U6577 ( .A1(n5985), .A2(n5978), .ZN(n6107) );
  NAND2_X1 U6578 ( .A1(n6107), .A2(n5110), .ZN(n9259) );
  INV_X1 U6579 ( .A(n9254), .ZN(n9255) );
  AND2_X1 U6580 ( .A1(n9335), .A2(n4719), .ZN(n9622) );
  AND2_X1 U6581 ( .A1(n8199), .A2(n9381), .ZN(n9399) );
  INV_X1 U6582 ( .A(n9600), .ZN(n9556) );
  AND2_X1 U6583 ( .A1(n6397), .A2(n6396), .ZN(n6467) );
  AND2_X1 U6584 ( .A1(n6400), .A2(n8278), .ZN(n9693) );
  NAND2_X1 U6585 ( .A1(n7355), .A2(n9737), .ZN(n9834) );
  AND2_X1 U6586 ( .A1(n8271), .A2(n6904), .ZN(n6409) );
  INV_X1 U6587 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n10342) );
  INV_X1 U6588 ( .A(n6083), .ZN(n5863) );
  AND2_X1 U6589 ( .A1(n8787), .A2(n7627), .ZN(n9978) );
  AND2_X1 U6590 ( .A1(n5905), .A2(n5904), .ZN(n8428) );
  AND2_X1 U6591 ( .A1(n5890), .A2(n5889), .ZN(n8421) );
  NAND2_X1 U6592 ( .A1(n5700), .A2(n5699), .ZN(n8602) );
  INV_X1 U6593 ( .A(n10026), .ZN(n10044) );
  INV_X1 U6594 ( .A(n6936), .ZN(n10008) );
  OR2_X1 U6595 ( .A1(P2_U3150), .A2(n6168), .ZN(n9888) );
  INV_X1 U6596 ( .A(n9877), .ZN(n9971) );
  MUX2_X1 U6597 ( .A(n6165), .B(n8531), .S(n7786), .Z(n9977) );
  OR2_X1 U6598 ( .A1(n6226), .A2(n8561), .ZN(n9963) );
  INV_X1 U6599 ( .A(n8795), .ZN(n8731) );
  NAND2_X1 U6600 ( .A1(n10087), .A2(n10019), .ZN(n8893) );
  INV_X1 U6601 ( .A(n10087), .ZN(n10085) );
  INV_X1 U6602 ( .A(n8665), .ZN(n8929) );
  OR2_X1 U6603 ( .A1(n10070), .A2(n10064), .ZN(n8974) );
  INV_X2 U6604 ( .A(n10070), .ZN(n10068) );
  INV_X1 U6605 ( .A(n8500), .ZN(n9923) );
  INV_X1 U6606 ( .A(n9408), .ZN(n9652) );
  INV_X1 U6607 ( .A(n9376), .ZN(n9639) );
  INV_X1 U6608 ( .A(n9162), .ZN(n9126) );
  NAND2_X1 U6609 ( .A1(n6486), .A2(n6471), .ZN(n9164) );
  NAND2_X1 U6610 ( .A1(n6107), .A2(n5968), .ZN(n9258) );
  INV_X1 U6611 ( .A(n9569), .ZN(n9590) );
  NAND2_X1 U6612 ( .A1(n9598), .A2(n7011), .ZN(n9600) );
  NAND2_X1 U6613 ( .A1(n9850), .A2(n9712), .ZN(n9742) );
  NAND3_X1 U6614 ( .A1(n6409), .A2(n6408), .A3(n6467), .ZN(n9847) );
  NAND2_X1 U6615 ( .A1(n9838), .A2(n9712), .ZN(n9783) );
  NAND3_X1 U6616 ( .A1(n6409), .A2(n6408), .A3(n6908), .ZN(n9836) );
  INV_X1 U6617 ( .A(n9797), .ZN(n9799) );
  NOR2_X1 U6618 ( .A1(n6097), .A2(n6480), .ZN(n8271) );
  INV_X1 U6619 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7498) );
  INV_X2 U6620 ( .A(n9176), .ZN(P1_U3973) );
  NOR2_X1 U6621 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5120) );
  NAND2_X1 U6622 ( .A1(n5404), .A2(n5405), .ZN(n5424) );
  INV_X1 U6623 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5121) );
  NAND2_X1 U6624 ( .A1(n5441), .A2(n5121), .ZN(n5122) );
  NAND2_X1 U6625 ( .A1(n5125), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U6626 ( .A1(n5516), .A2(n5515), .ZN(n5518) );
  NAND2_X1 U6627 ( .A1(n5518), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5126) );
  NOR2_X1 U6628 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5127) );
  NAND4_X1 U6629 ( .A1(n5127), .A2(n5405), .A3(n5438), .A4(n5441), .ZN(n5132)
         );
  NAND4_X1 U6630 ( .A1(n5130), .A2(n5479), .A3(n5129), .A4(n5128), .ZN(n5131)
         );
  NOR2_X1 U6631 ( .A1(n5132), .A2(n5131), .ZN(n5133) );
  NAND2_X1 U6632 ( .A1(n4550), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5134) );
  NAND2_X1 U6633 ( .A1(n5139), .A2(n7789), .ZN(n5812) );
  NAND2_X1 U6634 ( .A1(n4558), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5135) );
  MUX2_X1 U6635 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5135), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n5136) );
  NAND2_X1 U6636 ( .A1(n5137), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5138) );
  NAND2_X1 U6637 ( .A1(n7626), .A2(n7782), .ZN(n5866) );
  NAND2_X1 U6638 ( .A1(n5906), .A2(n10062), .ZN(n6718) );
  AND2_X1 U6639 ( .A1(n5867), .A2(n5812), .ZN(n5140) );
  OR2_X1 U6640 ( .A1(n6718), .A2(n5140), .ZN(n9988) );
  NAND2_X1 U6641 ( .A1(n7784), .A2(n7782), .ZN(n6412) );
  OR2_X1 U6642 ( .A1(n6412), .A2(n7789), .ZN(n10055) );
  NAND2_X1 U6643 ( .A1(n5148), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5149) );
  INV_X1 U6644 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U6645 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5152) );
  MUX2_X1 U6646 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5152), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5155) );
  INV_X1 U6647 ( .A(n6178), .ZN(n5154) );
  NAND2_X1 U6648 ( .A1(n5156), .A2(SI_1_), .ZN(n5193) );
  INV_X1 U6649 ( .A(SI_1_), .ZN(n10343) );
  NAND2_X1 U6650 ( .A1(n5193), .A2(n5157), .ZN(n5164) );
  INV_X1 U6651 ( .A(n5164), .ZN(n5161) );
  INV_X1 U6652 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5188) );
  INV_X1 U6653 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5941) );
  NOR2_X1 U6654 ( .A1(n5160), .A2(n10450), .ZN(n5162) );
  NAND2_X1 U6655 ( .A1(n5161), .A2(n5162), .ZN(n5194) );
  INV_X1 U6656 ( .A(n5162), .ZN(n5163) );
  NAND2_X1 U6657 ( .A1(n5164), .A2(n5163), .ZN(n5165) );
  NAND2_X1 U6658 ( .A1(n5194), .A2(n5165), .ZN(n6434) );
  OR2_X1 U6659 ( .A1(n5222), .A2(n6434), .ZN(n5166) );
  INV_X1 U6660 ( .A(n5167), .ZN(n5169) );
  NOR2_X1 U6661 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n5168) );
  NAND2_X1 U6662 ( .A1(n5169), .A2(n5168), .ZN(n8979) );
  NAND2_X1 U6663 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), 
        .ZN(n5171) );
  NAND2_X1 U6664 ( .A1(n5172), .A2(n5171), .ZN(n5174) );
  XNOR2_X2 U6665 ( .A(n5174), .B(n5173), .ZN(n5175) );
  NAND2_X1 U6666 ( .A1(n7554), .A2(n5175), .ZN(n5212) );
  INV_X1 U6667 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6155) );
  OR2_X1 U6668 ( .A1(n5212), .A2(n6155), .ZN(n5181) );
  INV_X1 U6669 ( .A(n7554), .ZN(n5177) );
  INV_X1 U6670 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n8789) );
  OR2_X1 U6671 ( .A1(n5213), .A2(n8789), .ZN(n5180) );
  NAND2_X2 U6672 ( .A1(n7554), .A2(n8287), .ZN(n5211) );
  INV_X1 U6673 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5176) );
  OR2_X1 U6674 ( .A1(n5211), .A2(n5176), .ZN(n5179) );
  NAND2_X2 U6675 ( .A1(n5177), .A2(n8287), .ZN(n5214) );
  INV_X1 U6676 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n8803) );
  INV_X1 U6677 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6717) );
  OR2_X1 U6678 ( .A1(n5213), .A2(n6717), .ZN(n5187) );
  INV_X1 U6679 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6170) );
  OR2_X1 U6680 ( .A1(n5214), .A2(n6170), .ZN(n5186) );
  NAND2_X1 U6681 ( .A1(n5182), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5185) );
  INV_X1 U6682 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5183) );
  INV_X1 U6683 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U6684 ( .A1(n7468), .A2(SI_0_), .ZN(n5189) );
  XNOR2_X1 U6685 ( .A(n5189), .B(n5188), .ZN(n8995) );
  MUX2_X1 U6686 ( .A(n6177), .B(n8995), .S(n5861), .Z(n6211) );
  INV_X1 U6687 ( .A(n6211), .ZN(n5191) );
  NAND2_X1 U6688 ( .A1(n5721), .A2(n5191), .ZN(n8787) );
  INV_X1 U6689 ( .A(n8787), .ZN(n5192) );
  NAND2_X1 U6690 ( .A1(n8785), .A2(n7629), .ZN(n6773) );
  NAND2_X1 U6691 ( .A1(n6178), .A2(n4911), .ZN(n5219) );
  NAND2_X1 U6692 ( .A1(n5194), .A2(n5193), .ZN(n5200) );
  INV_X1 U6693 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5196) );
  NAND2_X1 U6694 ( .A1(n5197), .A2(SI_2_), .ZN(n5223) );
  OAI21_X1 U6695 ( .B1(n5197), .B2(SI_2_), .A(n5223), .ZN(n5199) );
  NAND2_X1 U6696 ( .A1(n5198), .A2(n5199), .ZN(n5202) );
  INV_X1 U6697 ( .A(n5199), .ZN(n5201) );
  NAND2_X1 U6698 ( .A1(n5201), .A2(n5200), .ZN(n5224) );
  NAND2_X1 U6699 ( .A1(n5202), .A2(n5224), .ZN(n6443) );
  OR2_X1 U6700 ( .A1(n5222), .A2(n6443), .ZN(n5204) );
  INV_X1 U6701 ( .A(n5873), .ZN(n9989) );
  INV_X1 U6702 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9874) );
  OR2_X1 U6703 ( .A1(n5213), .A2(n9874), .ZN(n5209) );
  OR2_X1 U6704 ( .A1(n5212), .A2(n10073), .ZN(n5208) );
  INV_X1 U6705 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5205) );
  INV_X1 U6706 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6778) );
  OR2_X1 U6707 ( .A1(n9989), .A2(n9998), .ZN(n7637) );
  NAND2_X1 U6708 ( .A1(n9989), .A2(n9998), .ZN(n7638) );
  NAND2_X1 U6709 ( .A1(n7637), .A2(n7638), .ZN(n7590) );
  INV_X1 U6710 ( .A(n7590), .ZN(n7635) );
  NAND2_X1 U6711 ( .A1(n6773), .A2(n7635), .ZN(n5210) );
  NAND2_X1 U6712 ( .A1(n5182), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5218) );
  OR2_X1 U6713 ( .A1(n6625), .A2(n10075), .ZN(n5217) );
  OR2_X1 U6714 ( .A1(n5484), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5216) );
  INV_X1 U6715 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6926) );
  OR2_X1 U6716 ( .A1(n5214), .A2(n6926), .ZN(n5215) );
  AND4_X2 U6717 ( .A1(n5218), .A2(n5217), .A3(n5216), .A4(n5215), .ZN(n6936)
         );
  NAND2_X1 U6718 ( .A1(n5219), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5220) );
  MUX2_X1 U6719 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5220), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5221) );
  NAND2_X1 U6720 ( .A1(n5221), .A2(n5257), .ZN(n6164) );
  NAND2_X1 U6721 ( .A1(n5224), .A2(n5223), .ZN(n5230) );
  MUX2_X1 U6722 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n6433), .Z(n5225) );
  NAND2_X1 U6723 ( .A1(n5225), .A2(SI_3_), .ZN(n5245) );
  INV_X1 U6724 ( .A(n5225), .ZN(n5227) );
  INV_X1 U6725 ( .A(SI_3_), .ZN(n5226) );
  NAND2_X1 U6726 ( .A1(n5227), .A2(n5226), .ZN(n5228) );
  AND2_X1 U6727 ( .A1(n5245), .A2(n5228), .ZN(n5229) );
  OR2_X1 U6728 ( .A1(n5230), .A2(n5229), .ZN(n5231) );
  NAND2_X1 U6729 ( .A1(n5246), .A2(n5231), .ZN(n6534) );
  OR2_X1 U6730 ( .A1(n5222), .A2(n6534), .ZN(n5233) );
  INV_X1 U6731 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6069) );
  OR2_X1 U6732 ( .A1(n7577), .A2(n6069), .ZN(n5232) );
  NAND2_X1 U6733 ( .A1(n6922), .A2(n7592), .ZN(n6921) );
  NAND2_X1 U6734 ( .A1(n6921), .A2(n7658), .ZN(n6933) );
  NAND2_X1 U6735 ( .A1(n5711), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5242) );
  INV_X1 U6736 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5234) );
  OR2_X1 U6737 ( .A1(n5211), .A2(n5234), .ZN(n5241) );
  INV_X1 U6738 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5236) );
  INV_X1 U6739 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5235) );
  NAND2_X1 U6740 ( .A1(n5236), .A2(n5235), .ZN(n5272) );
  NAND2_X1 U6741 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5237) );
  AND2_X1 U6742 ( .A1(n5272), .A2(n5237), .ZN(n6934) );
  OR2_X1 U6743 ( .A1(n5484), .A2(n6934), .ZN(n5240) );
  INV_X1 U6744 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5238) );
  OR2_X1 U6745 ( .A1(n5214), .A2(n5238), .ZN(n5239) );
  NAND2_X1 U6746 ( .A1(n5257), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5244) );
  INV_X1 U6747 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5243) );
  XNOR2_X1 U6748 ( .A(n5244), .B(n5243), .ZN(n6289) );
  INV_X1 U6749 ( .A(n5247), .ZN(n5249) );
  INV_X1 U6750 ( .A(SI_4_), .ZN(n5248) );
  NAND2_X1 U6751 ( .A1(n5249), .A2(n5248), .ZN(n5250) );
  AND2_X1 U6752 ( .A1(n5260), .A2(n5250), .ZN(n5251) );
  OR2_X1 U6753 ( .A1(n5252), .A2(n5251), .ZN(n5253) );
  NAND2_X1 U6754 ( .A1(n5261), .A2(n5253), .ZN(n6545) );
  OR2_X1 U6755 ( .A1(n5222), .A2(n6545), .ZN(n5255) );
  INV_X1 U6756 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6071) );
  OR2_X1 U6757 ( .A1(n7577), .A2(n6071), .ZN(n5254) );
  OAI211_X1 U6758 ( .C1(n5861), .C2(n6289), .A(n5255), .B(n5254), .ZN(n10007)
         );
  OR2_X1 U6759 ( .A1(n10001), .A2(n10007), .ZN(n7659) );
  NAND2_X1 U6760 ( .A1(n10001), .A2(n10007), .ZN(n7645) );
  NAND2_X1 U6761 ( .A1(n6933), .A2(n7642), .ZN(n5256) );
  OR2_X1 U6762 ( .A1(n5257), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5279) );
  NAND2_X1 U6763 ( .A1(n5279), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5259) );
  XNOR2_X1 U6764 ( .A(n5259), .B(n5258), .ZN(n6261) );
  MUX2_X1 U6765 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n6433), .Z(n5262) );
  NAND2_X1 U6766 ( .A1(n5262), .A2(SI_5_), .ZN(n5285) );
  INV_X1 U6767 ( .A(n5262), .ZN(n5264) );
  INV_X1 U6768 ( .A(SI_5_), .ZN(n5263) );
  NAND2_X1 U6769 ( .A1(n5264), .A2(n5263), .ZN(n5265) );
  AND2_X1 U6770 ( .A1(n5285), .A2(n5265), .ZN(n5266) );
  OR2_X1 U6771 ( .A1(n5267), .A2(n5266), .ZN(n5268) );
  NAND2_X1 U6772 ( .A1(n5286), .A2(n5268), .ZN(n6727) );
  OR2_X1 U6773 ( .A1(n5222), .A2(n6727), .ZN(n5270) );
  INV_X1 U6774 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6072) );
  OR2_X1 U6775 ( .A1(n7577), .A2(n6072), .ZN(n5269) );
  INV_X1 U6776 ( .A(n6427), .ZN(n10014) );
  NAND2_X1 U6777 ( .A1(n5182), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5277) );
  INV_X1 U6778 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6259) );
  OR2_X1 U6779 ( .A1(n6625), .A2(n6259), .ZN(n5276) );
  INV_X1 U6780 ( .A(n5272), .ZN(n5271) );
  NAND2_X1 U6781 ( .A1(n5271), .A2(n10404), .ZN(n5295) );
  NAND2_X1 U6782 ( .A1(n5272), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5273) );
  AND2_X1 U6783 ( .A1(n5295), .A2(n5273), .ZN(n6424) );
  OR2_X1 U6784 ( .A1(n5484), .A2(n6424), .ZN(n5275) );
  INV_X1 U6785 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6260) );
  OR2_X1 U6786 ( .A1(n6628), .A2(n6260), .ZN(n5274) );
  NAND4_X1 U6787 ( .A1(n5277), .A2(n5276), .A3(n5275), .A4(n5274), .ZN(n8441)
         );
  OR2_X1 U6788 ( .A1(n10014), .A2(n8441), .ZN(n7664) );
  INV_X1 U6789 ( .A(n7664), .ZN(n5278) );
  OR2_X2 U6790 ( .A1(n6413), .A2(n5278), .ZN(n6761) );
  NOR2_X1 U6791 ( .A1(n5279), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5283) );
  INV_X1 U6792 ( .A(n5283), .ZN(n5280) );
  NAND2_X1 U6793 ( .A1(n5280), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5281) );
  MUX2_X1 U6794 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5281), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5284) );
  INV_X1 U6795 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5282) );
  NAND2_X1 U6796 ( .A1(n5283), .A2(n5282), .ZN(n5325) );
  NAND2_X1 U6797 ( .A1(n5284), .A2(n5325), .ZN(n6505) );
  MUX2_X1 U6798 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6433), .Z(n5287) );
  NAND2_X1 U6799 ( .A1(n5287), .A2(SI_6_), .ZN(n5302) );
  INV_X1 U6800 ( .A(n5287), .ZN(n5288) );
  NAND2_X1 U6801 ( .A1(n5288), .A2(n10338), .ZN(n5289) );
  AND2_X1 U6802 ( .A1(n5302), .A2(n5289), .ZN(n5290) );
  OR2_X1 U6803 ( .A1(n4584), .A2(n5290), .ZN(n5291) );
  NAND2_X1 U6804 ( .A1(n5303), .A2(n5291), .ZN(n6848) );
  OR2_X1 U6805 ( .A1(n6848), .A2(n5222), .ZN(n5293) );
  INV_X1 U6806 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6074) );
  OR2_X1 U6807 ( .A1(n7577), .A2(n6074), .ZN(n5292) );
  OAI211_X1 U6808 ( .C1(n5861), .C2(n6505), .A(n5293), .B(n5292), .ZN(n10021)
         );
  INV_X1 U6809 ( .A(n10021), .ZN(n6766) );
  NAND2_X1 U6810 ( .A1(n5711), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5300) );
  INV_X1 U6811 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5294) );
  OR2_X1 U6812 ( .A1(n5211), .A2(n5294), .ZN(n5299) );
  NAND2_X1 U6813 ( .A1(n5295), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5296) );
  AND2_X1 U6814 ( .A1(n5316), .A2(n5296), .ZN(n6765) );
  OR2_X1 U6815 ( .A1(n5484), .A2(n6765), .ZN(n5298) );
  INV_X1 U6816 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6508) );
  OR2_X1 U6817 ( .A1(n6628), .A2(n6508), .ZN(n5297) );
  NAND4_X1 U6818 ( .A1(n5300), .A2(n5299), .A3(n5298), .A4(n5297), .ZN(n8440)
         );
  NAND2_X1 U6819 ( .A1(n6766), .A2(n8440), .ZN(n7666) );
  NAND2_X1 U6820 ( .A1(n10014), .A2(n8441), .ZN(n7660) );
  AND2_X1 U6821 ( .A1(n7666), .A2(n7660), .ZN(n7647) );
  NAND2_X1 U6822 ( .A1(n6761), .A2(n7647), .ZN(n5301) );
  INV_X1 U6823 ( .A(n8440), .ZN(n10028) );
  NAND2_X1 U6824 ( .A1(n10028), .A2(n10021), .ZN(n7663) );
  NAND2_X1 U6825 ( .A1(n5301), .A2(n7663), .ZN(n6992) );
  INV_X1 U6826 ( .A(n6992), .ZN(n5322) );
  MUX2_X1 U6827 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6433), .Z(n5304) );
  NAND2_X1 U6828 ( .A1(n5304), .A2(SI_7_), .ZN(n5323) );
  INV_X1 U6829 ( .A(n5304), .ZN(n5306) );
  INV_X1 U6830 ( .A(SI_7_), .ZN(n5305) );
  NAND2_X1 U6831 ( .A1(n5306), .A2(n5305), .ZN(n5307) );
  AND2_X1 U6832 ( .A1(n5323), .A2(n5307), .ZN(n5308) );
  OR2_X1 U6833 ( .A1(n5309), .A2(n5308), .ZN(n5310) );
  NAND2_X1 U6834 ( .A1(n5324), .A2(n5310), .ZN(n7026) );
  OR2_X1 U6835 ( .A1(n7026), .A2(n5222), .ZN(n5313) );
  NAND2_X1 U6836 ( .A1(n5325), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5311) );
  XNOR2_X1 U6837 ( .A(n5311), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6506) );
  AOI22_X1 U6838 ( .A1(n5538), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5537), .B2(
        n6506), .ZN(n5312) );
  NAND2_X1 U6839 ( .A1(n5313), .A2(n5312), .ZN(n10030) );
  NAND2_X1 U6840 ( .A1(n5182), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5321) );
  INV_X1 U6841 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6499) );
  OR2_X1 U6842 ( .A1(n6625), .A2(n6499), .ZN(n5320) );
  INV_X1 U6843 ( .A(n5316), .ZN(n5315) );
  INV_X1 U6844 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5314) );
  NAND2_X1 U6845 ( .A1(n5315), .A2(n5314), .ZN(n5330) );
  NAND2_X1 U6846 ( .A1(n5316), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5317) );
  AND2_X1 U6847 ( .A1(n5330), .A2(n5317), .ZN(n6995) );
  OR2_X1 U6848 ( .A1(n5484), .A2(n6995), .ZN(n5319) );
  INV_X1 U6849 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6500) );
  OR2_X1 U6850 ( .A1(n5214), .A2(n6500), .ZN(n5318) );
  NAND4_X1 U6851 ( .A1(n5321), .A2(n5320), .A3(n5319), .A4(n5318), .ZN(n8439)
         );
  OR2_X1 U6852 ( .A1(n10030), .A2(n6785), .ZN(n6781) );
  NAND2_X1 U6853 ( .A1(n10030), .A2(n6785), .ZN(n7669) );
  MUX2_X1 U6854 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n6433), .Z(n5337) );
  XNOR2_X1 U6855 ( .A(n5337), .B(SI_8_), .ZN(n5339) );
  XNOR2_X1 U6856 ( .A(n5340), .B(n5339), .ZN(n7033) );
  NAND2_X1 U6857 ( .A1(n7033), .A2(n7579), .ZN(n5328) );
  NAND2_X1 U6858 ( .A1(n5342), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5326) );
  XNOR2_X1 U6859 ( .A(n5326), .B(P2_IR_REG_8__SCAN_IN), .ZN(n8450) );
  AOI22_X1 U6860 ( .A1(n5538), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5537), .B2(
        n8450), .ZN(n5327) );
  NAND2_X1 U6861 ( .A1(n5328), .A2(n5327), .ZN(n6789) );
  NAND2_X1 U6862 ( .A1(n5711), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5335) );
  INV_X1 U6863 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5329) );
  OR2_X1 U6864 ( .A1(n5211), .A2(n5329), .ZN(n5334) );
  NAND2_X1 U6865 ( .A1(n5330), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5331) );
  AND2_X1 U6866 ( .A1(n5350), .A2(n5331), .ZN(n6786) );
  OR2_X1 U6867 ( .A1(n5484), .A2(n6786), .ZN(n5333) );
  INV_X1 U6868 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6787) );
  OR2_X1 U6869 ( .A1(n6628), .A2(n6787), .ZN(n5332) );
  OR2_X1 U6870 ( .A1(n6789), .A2(n10026), .ZN(n7652) );
  AND2_X1 U6871 ( .A1(n7652), .A2(n6781), .ZN(n7650) );
  NAND2_X1 U6872 ( .A1(n6993), .A2(n7650), .ZN(n5336) );
  NAND2_X1 U6873 ( .A1(n6789), .A2(n10026), .ZN(n7670) );
  INV_X1 U6874 ( .A(n5337), .ZN(n5338) );
  INV_X1 U6875 ( .A(SI_8_), .ZN(n10417) );
  INV_X1 U6876 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6090) );
  INV_X1 U6877 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5341) );
  MUX2_X1 U6878 ( .A(n6090), .B(n5341), .S(n6433), .Z(n5358) );
  XNOR2_X1 U6879 ( .A(n5358), .B(SI_9_), .ZN(n5360) );
  XNOR2_X1 U6880 ( .A(n5361), .B(n5360), .ZN(n7228) );
  NAND2_X1 U6881 ( .A1(n7228), .A2(n7579), .ZN(n5347) );
  OAI21_X1 U6882 ( .B1(n5342), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5344) );
  INV_X1 U6883 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5343) );
  OR2_X1 U6884 ( .A1(n5344), .A2(n5343), .ZN(n5345) );
  NAND2_X1 U6885 ( .A1(n5344), .A2(n5343), .ZN(n5369) );
  AOI22_X1 U6886 ( .A1(n5538), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5537), .B2(
        n6892), .ZN(n5346) );
  NAND2_X1 U6887 ( .A1(n5347), .A2(n5346), .ZN(n10045) );
  NAND2_X1 U6888 ( .A1(n5182), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5356) );
  INV_X1 U6889 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6971) );
  OR2_X1 U6890 ( .A1(n5214), .A2(n6971), .ZN(n5355) );
  INV_X1 U6891 ( .A(n5350), .ZN(n5349) );
  INV_X1 U6892 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U6893 ( .A1(n5349), .A2(n5348), .ZN(n5374) );
  NAND2_X1 U6894 ( .A1(n5350), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5351) );
  AND2_X1 U6895 ( .A1(n5374), .A2(n5351), .ZN(n6970) );
  OR2_X1 U6896 ( .A1(n5484), .A2(n6970), .ZN(n5354) );
  INV_X1 U6897 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5352) );
  OR2_X1 U6898 ( .A1(n6625), .A2(n5352), .ZN(n5353) );
  NAND4_X1 U6899 ( .A1(n5356), .A2(n5355), .A3(n5354), .A4(n5353), .ZN(n8438)
         );
  NAND2_X1 U6900 ( .A1(n10045), .A2(n6947), .ZN(n7672) );
  NAND2_X1 U6901 ( .A1(n7655), .A2(n7672), .ZN(n7601) );
  INV_X1 U6902 ( .A(n7601), .ZN(n5357) );
  INV_X1 U6903 ( .A(n5358), .ZN(n5359) );
  MUX2_X1 U6904 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6433), .Z(n5362) );
  NAND2_X1 U6905 ( .A1(n5362), .A2(SI_10_), .ZN(n5381) );
  INV_X1 U6906 ( .A(n5362), .ZN(n5363) );
  INV_X1 U6907 ( .A(SI_10_), .ZN(n10451) );
  NAND2_X1 U6908 ( .A1(n5363), .A2(n10451), .ZN(n5364) );
  NAND2_X1 U6909 ( .A1(n5381), .A2(n5364), .ZN(n5366) );
  INV_X1 U6910 ( .A(n5366), .ZN(n5365) );
  NAND2_X1 U6911 ( .A1(n5367), .A2(n5366), .ZN(n5368) );
  NAND2_X1 U6912 ( .A1(n5382), .A2(n5368), .ZN(n7252) );
  NAND2_X1 U6913 ( .A1(n5369), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5370) );
  XNOR2_X1 U6914 ( .A(n5370), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6895) );
  AOI22_X1 U6915 ( .A1(n5538), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5537), .B2(
        n6895), .ZN(n5371) );
  NAND2_X1 U6916 ( .A1(n5372), .A2(n5371), .ZN(n10059) );
  NAND2_X1 U6917 ( .A1(n5182), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5379) );
  INV_X1 U6918 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5373) );
  OR2_X1 U6919 ( .A1(n6625), .A2(n5373), .ZN(n5378) );
  NAND2_X1 U6920 ( .A1(n5374), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5375) );
  AND2_X1 U6921 ( .A1(n5388), .A2(n5375), .ZN(n6988) );
  OR2_X1 U6922 ( .A1(n5484), .A2(n6988), .ZN(n5377) );
  INV_X1 U6923 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6896) );
  OR2_X1 U6924 ( .A1(n6628), .A2(n6896), .ZN(n5376) );
  NAND4_X1 U6925 ( .A1(n5379), .A2(n5378), .A3(n5377), .A4(n5376), .ZN(n10041)
         );
  INV_X1 U6926 ( .A(n7679), .ZN(n5380) );
  NAND2_X1 U6927 ( .A1(n10059), .A2(n7186), .ZN(n7678) );
  MUX2_X1 U6928 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6433), .Z(n5396) );
  XNOR2_X1 U6929 ( .A(n5396), .B(SI_11_), .ZN(n5397) );
  XNOR2_X1 U6930 ( .A(n5398), .B(n5397), .ZN(n7339) );
  NAND2_X1 U6931 ( .A1(n7339), .A2(n7579), .ZN(n5386) );
  OR2_X1 U6932 ( .A1(n5383), .A2(n5403), .ZN(n5384) );
  XNOR2_X1 U6933 ( .A(n5384), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8496) );
  AOI22_X1 U6934 ( .A1(n5538), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5537), .B2(
        n8496), .ZN(n5385) );
  NAND2_X1 U6935 ( .A1(n5386), .A2(n5385), .ZN(n7190) );
  NAND2_X1 U6936 ( .A1(n5182), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5393) );
  INV_X1 U6937 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5387) );
  OR2_X1 U6938 ( .A1(n6625), .A2(n5387), .ZN(n5392) );
  NAND2_X1 U6939 ( .A1(n5388), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5389) );
  AND2_X1 U6940 ( .A1(n5410), .A2(n5389), .ZN(n7187) );
  OR2_X1 U6941 ( .A1(n5484), .A2(n7187), .ZN(n5391) );
  INV_X1 U6942 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7188) );
  OR2_X1 U6943 ( .A1(n6628), .A2(n7188), .ZN(n5390) );
  NAND4_X1 U6944 ( .A1(n5393), .A2(n5392), .A3(n5391), .A4(n5390), .ZN(n8437)
         );
  NAND2_X1 U6945 ( .A1(n7190), .A2(n7321), .ZN(n7683) );
  INV_X1 U6946 ( .A(n7683), .ZN(n5394) );
  OR2_X1 U6947 ( .A1(n7190), .A2(n7321), .ZN(n7682) );
  NAND2_X1 U6948 ( .A1(n5395), .A2(n7682), .ZN(n7153) );
  MUX2_X1 U6949 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6433), .Z(n5399) );
  NAND2_X1 U6950 ( .A1(n5399), .A2(SI_12_), .ZN(n5416) );
  OAI21_X1 U6951 ( .B1(n5399), .B2(SI_12_), .A(n5416), .ZN(n5400) );
  NAND2_X1 U6952 ( .A1(n5401), .A2(n5400), .ZN(n5402) );
  NAND2_X1 U6953 ( .A1(n5402), .A2(n5417), .ZN(n7365) );
  OR2_X1 U6954 ( .A1(n7365), .A2(n5222), .ZN(n5408) );
  OR2_X1 U6955 ( .A1(n5404), .A2(n5403), .ZN(n5406) );
  XNOR2_X1 U6956 ( .A(n5406), .B(n5405), .ZN(n9905) );
  INV_X1 U6957 ( .A(n9905), .ZN(n8481) );
  AOI22_X1 U6958 ( .A1(n5538), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5537), .B2(
        n8481), .ZN(n5407) );
  NAND2_X1 U6959 ( .A1(n5182), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5415) );
  INV_X1 U6960 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7325) );
  OR2_X1 U6961 ( .A1(n6625), .A2(n7325), .ZN(n5414) );
  INV_X1 U6962 ( .A(n5410), .ZN(n5409) );
  NAND2_X1 U6963 ( .A1(n5409), .A2(n10476), .ZN(n5428) );
  NAND2_X1 U6964 ( .A1(n5410), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5411) );
  AND2_X1 U6965 ( .A1(n5428), .A2(n5411), .ZN(n7292) );
  OR2_X1 U6966 ( .A1(n5484), .A2(n7292), .ZN(n5413) );
  INV_X1 U6967 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7158) );
  OR2_X1 U6968 ( .A1(n6628), .A2(n7158), .ZN(n5412) );
  NAND4_X1 U6969 ( .A1(n5415), .A2(n5414), .A3(n5413), .A4(n5412), .ZN(n8775)
         );
  XNOR2_X1 U6970 ( .A(n7688), .B(n8775), .ZN(n7684) );
  INV_X1 U6971 ( .A(n8775), .ZN(n8392) );
  OR2_X1 U6972 ( .A1(n7688), .A2(n8392), .ZN(n7690) );
  MUX2_X1 U6973 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6433), .Z(n5418) );
  NAND2_X1 U6974 ( .A1(n5418), .A2(SI_13_), .ZN(n5435) );
  INV_X1 U6975 ( .A(n5418), .ZN(n5419) );
  NAND2_X1 U6976 ( .A1(n5419), .A2(n10246), .ZN(n5420) );
  OR2_X1 U6977 ( .A1(n5422), .A2(n5421), .ZN(n5423) );
  NAND2_X1 U6978 ( .A1(n5436), .A2(n5423), .ZN(n7505) );
  OR2_X1 U6979 ( .A1(n7505), .A2(n5222), .ZN(n5426) );
  NAND2_X1 U6980 ( .A1(n5424), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5439) );
  XNOR2_X1 U6981 ( .A(n5439), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8500) );
  AOI22_X1 U6982 ( .A1(n5538), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5537), .B2(
        n8500), .ZN(n5425) );
  NAND2_X1 U6983 ( .A1(n5182), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5433) );
  INV_X1 U6984 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9908) );
  OR2_X1 U6985 ( .A1(n6625), .A2(n9908), .ZN(n5432) );
  INV_X1 U6986 ( .A(n5428), .ZN(n5427) );
  NAND2_X1 U6987 ( .A1(n5427), .A2(n10393), .ZN(n5447) );
  NAND2_X1 U6988 ( .A1(n5428), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5429) );
  AND2_X1 U6989 ( .A1(n5447), .A2(n5429), .ZN(n8777) );
  OR2_X1 U6990 ( .A1(n5484), .A2(n8777), .ZN(n5431) );
  INV_X1 U6991 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n9915) );
  OR2_X1 U6992 ( .A1(n6628), .A2(n9915), .ZN(n5430) );
  NAND4_X1 U6993 ( .A1(n5433), .A2(n5432), .A3(n5431), .A4(n5430), .ZN(n8763)
         );
  AND2_X1 U6994 ( .A1(n8971), .A2(n8021), .ZN(n7695) );
  INV_X1 U6995 ( .A(n7695), .ZN(n5434) );
  NOR2_X1 U6996 ( .A1(n8971), .A2(n8021), .ZN(n7694) );
  MUX2_X1 U6997 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6433), .Z(n5454) );
  XNOR2_X1 U6998 ( .A(n5454), .B(SI_14_), .ZN(n5437) );
  XNOR2_X1 U6999 ( .A(n5455), .B(n5437), .ZN(n7509) );
  NAND2_X1 U7000 ( .A1(n7509), .A2(n7579), .ZN(n5445) );
  NAND2_X1 U7001 ( .A1(n5439), .A2(n5438), .ZN(n5440) );
  NAND2_X1 U7002 ( .A1(n5440), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5442) );
  NAND2_X1 U7003 ( .A1(n5442), .A2(n5441), .ZN(n5457) );
  OR2_X1 U7004 ( .A1(n5442), .A2(n5441), .ZN(n5443) );
  NAND2_X1 U7005 ( .A1(n5457), .A2(n5443), .ZN(n9940) );
  INV_X1 U7006 ( .A(n9940), .ZN(n8478) );
  AOI22_X1 U7007 ( .A1(n5538), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5537), .B2(
        n8478), .ZN(n5444) );
  NAND2_X1 U7008 ( .A1(n5182), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5452) );
  INV_X1 U7009 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5446) );
  OR2_X1 U7010 ( .A1(n6628), .A2(n5446), .ZN(n5451) );
  NAND2_X1 U7011 ( .A1(n5447), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5448) );
  AND2_X1 U7012 ( .A1(n5463), .A2(n5448), .ZN(n8766) );
  OR2_X1 U7013 ( .A1(n5484), .A2(n8766), .ZN(n5450) );
  INV_X1 U7014 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8887) );
  OR2_X1 U7015 ( .A1(n6625), .A2(n8887), .ZN(n5449) );
  NAND4_X1 U7016 ( .A1(n5452), .A2(n5451), .A3(n5450), .A4(n5449), .ZN(n8774)
         );
  INV_X1 U7017 ( .A(n8774), .ZN(n8023) );
  NAND2_X1 U7018 ( .A1(n8964), .A2(n8023), .ZN(n7699) );
  NAND2_X1 U7019 ( .A1(n8760), .A2(n7699), .ZN(n5453) );
  NAND2_X1 U7020 ( .A1(n5453), .A2(n7698), .ZN(n8749) );
  MUX2_X1 U7021 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6433), .Z(n5470) );
  XNOR2_X1 U7022 ( .A(n5470), .B(SI_15_), .ZN(n5456) );
  XNOR2_X1 U7023 ( .A(n5473), .B(n5456), .ZN(n7512) );
  NAND2_X1 U7024 ( .A1(n7512), .A2(n7579), .ZN(n5460) );
  NAND2_X1 U7025 ( .A1(n5457), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5458) );
  XNOR2_X1 U7026 ( .A(n5458), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8536) );
  AOI22_X1 U7027 ( .A1(n5538), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5537), .B2(
        n8536), .ZN(n5459) );
  NAND2_X1 U7028 ( .A1(n5182), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5468) );
  INV_X1 U7029 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8884) );
  OR2_X1 U7030 ( .A1(n6625), .A2(n8884), .ZN(n5467) );
  INV_X1 U7031 ( .A(n5463), .ZN(n5462) );
  NAND2_X1 U7032 ( .A1(n5463), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5464) );
  AND2_X1 U7033 ( .A1(n5485), .A2(n5464), .ZN(n8754) );
  OR2_X1 U7034 ( .A1(n5484), .A2(n8754), .ZN(n5466) );
  OR2_X1 U7035 ( .A1(n6628), .A2(n8476), .ZN(n5465) );
  NAND4_X1 U7036 ( .A1(n5468), .A2(n5467), .A3(n5466), .A4(n5465), .ZN(n8764)
         );
  NAND2_X1 U7037 ( .A1(n8958), .A2(n8357), .ZN(n7715) );
  NAND2_X1 U7038 ( .A1(n8749), .A2(n7715), .ZN(n5469) );
  NAND2_X1 U7039 ( .A1(n5469), .A2(n7703), .ZN(n8736) );
  INV_X1 U7040 ( .A(n5470), .ZN(n5471) );
  NAND2_X1 U7041 ( .A1(n5472), .A2(n5471), .ZN(n5475) );
  INV_X1 U7042 ( .A(SI_15_), .ZN(n5474) );
  MUX2_X1 U7043 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n6433), .Z(n5493) );
  INV_X1 U7044 ( .A(SI_16_), .ZN(n5476) );
  XNOR2_X1 U7045 ( .A(n5493), .B(n5476), .ZN(n5477) );
  NAND2_X1 U7046 ( .A1(n7515), .A2(n7579), .ZN(n5483) );
  NAND2_X1 U7047 ( .A1(n5478), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5480) );
  MUX2_X1 U7048 ( .A(n5480), .B(P2_IR_REG_31__SCAN_IN), .S(n5479), .Z(n5481)
         );
  NAND2_X1 U7049 ( .A1(n5481), .A2(n5498), .ZN(n9956) );
  INV_X1 U7050 ( .A(n9956), .ZN(n8539) );
  AOI22_X1 U7051 ( .A1(n5538), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5537), .B2(
        n8539), .ZN(n5482) );
  OR2_X2 U7052 ( .A1(n5485), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5504) );
  NAND2_X1 U7053 ( .A1(n5485), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5486) );
  NAND2_X1 U7054 ( .A1(n5504), .A2(n5486), .ZN(n8744) );
  NAND2_X1 U7055 ( .A1(n5710), .A2(n8744), .ZN(n5490) );
  INV_X1 U7056 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8881) );
  OR2_X1 U7057 ( .A1(n6625), .A2(n8881), .ZN(n5489) );
  INV_X1 U7058 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8952) );
  OR2_X1 U7059 ( .A1(n5211), .A2(n8952), .ZN(n5488) );
  INV_X1 U7060 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8743) );
  OR2_X1 U7061 ( .A1(n6628), .A2(n8743), .ZN(n5487) );
  NAND4_X1 U7062 ( .A1(n5490), .A2(n5489), .A3(n5488), .A4(n5487), .ZN(n8752)
         );
  INV_X1 U7063 ( .A(n8752), .ZN(n8726) );
  NAND2_X1 U7064 ( .A1(n5741), .A2(n8726), .ZN(n7625) );
  INV_X1 U7065 ( .A(n5491), .ZN(n5492) );
  NAND2_X1 U7066 ( .A1(n5493), .A2(SI_16_), .ZN(n5494) );
  MUX2_X1 U7067 ( .A(n6601), .B(n6599), .S(n6433), .Z(n5495) );
  NAND2_X1 U7068 ( .A1(n5495), .A2(n10434), .ZN(n5513) );
  INV_X1 U7069 ( .A(n5495), .ZN(n5496) );
  NAND2_X1 U7070 ( .A1(n5496), .A2(SI_17_), .ZN(n5497) );
  NAND2_X1 U7071 ( .A1(n5513), .A2(n5497), .ZN(n5511) );
  XNOR2_X1 U7072 ( .A(n5510), .B(n5511), .ZN(n7518) );
  NAND2_X1 U7073 ( .A1(n7518), .A2(n7579), .ZN(n5501) );
  NAND2_X1 U7074 ( .A1(n5498), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5499) );
  XNOR2_X1 U7075 ( .A(n5499), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8541) );
  AOI22_X1 U7076 ( .A1(n5538), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5537), .B2(
        n8541), .ZN(n5500) );
  INV_X1 U7077 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5502) );
  NAND2_X1 U7078 ( .A1(n5504), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U7079 ( .A1(n5521), .A2(n5505), .ZN(n8729) );
  NAND2_X1 U7080 ( .A1(n5710), .A2(n8729), .ZN(n5509) );
  INV_X1 U7081 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8948) );
  OR2_X1 U7082 ( .A1(n5211), .A2(n8948), .ZN(n5508) );
  INV_X1 U7083 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8519) );
  OR2_X1 U7084 ( .A1(n6628), .A2(n8519), .ZN(n5507) );
  INV_X1 U7085 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9960) );
  OR2_X1 U7086 ( .A1(n6625), .A2(n9960), .ZN(n5506) );
  NAND4_X1 U7087 ( .A1(n5509), .A2(n5508), .A3(n5507), .A4(n5506), .ZN(n8740)
         );
  OR2_X1 U7088 ( .A1(n8733), .A2(n8868), .ZN(n7718) );
  NAND2_X1 U7089 ( .A1(n8733), .A2(n8868), .ZN(n7708) );
  NAND2_X1 U7090 ( .A1(n8721), .A2(n7708), .ZN(n8713) );
  INV_X1 U7091 ( .A(n5511), .ZN(n5512) );
  MUX2_X1 U7092 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6433), .Z(n5530) );
  XNOR2_X1 U7093 ( .A(n5530), .B(n5514), .ZN(n5529) );
  XNOR2_X1 U7094 ( .A(n5533), .B(n5529), .ZN(n7521) );
  NAND2_X1 U7095 ( .A1(n7521), .A2(n7579), .ZN(n5520) );
  OR2_X1 U7096 ( .A1(n5516), .A2(n5515), .ZN(n5517) );
  AND2_X1 U7097 ( .A1(n5518), .A2(n5517), .ZN(n8558) );
  AOI22_X1 U7098 ( .A1(n5538), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5537), .B2(
        n8558), .ZN(n5519) );
  OR2_X2 U7099 ( .A1(n5521), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5542) );
  NAND2_X1 U7100 ( .A1(n5521), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U7101 ( .A1(n5542), .A2(n5522), .ZN(n8709) );
  NAND2_X1 U7102 ( .A1(n8709), .A2(n5710), .ZN(n5527) );
  NAND2_X1 U7103 ( .A1(n5711), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U7104 ( .A1(n5182), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5525) );
  INV_X1 U7105 ( .A(n5214), .ZN(n5523) );
  NAND2_X1 U7106 ( .A1(n5523), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5524) );
  NAND4_X1 U7107 ( .A1(n5527), .A2(n5526), .A3(n5525), .A4(n5524), .ZN(n8694)
         );
  NOR2_X1 U7108 ( .A1(n8873), .A2(n8876), .ZN(n7719) );
  INV_X1 U7109 ( .A(n7719), .ZN(n7722) );
  NAND2_X1 U7110 ( .A1(n8873), .A2(n8876), .ZN(n7725) );
  NAND2_X1 U7111 ( .A1(n7722), .A2(n7725), .ZN(n8708) );
  NOR2_X1 U7112 ( .A1(n8713), .A2(n8708), .ZN(n5528) );
  NAND2_X1 U7113 ( .A1(n8714), .A2(n7722), .ZN(n8701) );
  INV_X1 U7114 ( .A(n5529), .ZN(n5532) );
  NAND2_X1 U7115 ( .A1(n5530), .A2(SI_18_), .ZN(n5531) );
  MUX2_X1 U7116 ( .A(n6831), .B(n10247), .S(n6433), .Z(n5534) );
  INV_X1 U7117 ( .A(SI_19_), .ZN(n10394) );
  NAND2_X1 U7118 ( .A1(n5534), .A2(n10394), .ZN(n5547) );
  INV_X1 U7119 ( .A(n5534), .ZN(n5535) );
  NAND2_X1 U7120 ( .A1(n5535), .A2(SI_19_), .ZN(n5536) );
  NAND2_X1 U7121 ( .A1(n5547), .A2(n5536), .ZN(n5548) );
  XNOR2_X1 U7122 ( .A(n5549), .B(n5548), .ZN(n7524) );
  NAND2_X1 U7123 ( .A1(n7524), .A2(n7579), .ZN(n5540) );
  AOI22_X1 U7124 ( .A1(n5538), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7784), .B2(
        n5537), .ZN(n5539) );
  INV_X1 U7125 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U7126 ( .A1(n5542), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5543) );
  NAND2_X1 U7127 ( .A1(n5554), .A2(n5543), .ZN(n8697) );
  NAND2_X1 U7128 ( .A1(n8697), .A2(n5710), .ZN(n5545) );
  AOI22_X1 U7129 ( .A1(n5711), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n5182), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n5544) );
  OAI211_X1 U7130 ( .C1(n6628), .C2(n5546), .A(n5545), .B(n5544), .ZN(n8855)
         );
  INV_X1 U7131 ( .A(n8855), .ZN(n8869) );
  NAND2_X1 U7132 ( .A1(n8863), .A2(n8869), .ZN(n7727) );
  MUX2_X1 U7133 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6433), .Z(n5559) );
  XNOR2_X1 U7134 ( .A(n5559), .B(n5561), .ZN(n5550) );
  XNOR2_X1 U7135 ( .A(n5562), .B(n5550), .ZN(n7529) );
  NAND2_X1 U7136 ( .A1(n7529), .A2(n7579), .ZN(n5553) );
  INV_X1 U7137 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n5551) );
  OR2_X1 U7138 ( .A1(n7577), .A2(n5551), .ZN(n5552) );
  INV_X1 U7139 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5558) );
  NAND2_X1 U7140 ( .A1(n5554), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5555) );
  NAND2_X1 U7141 ( .A1(n5568), .A2(n5555), .ZN(n8685) );
  NAND2_X1 U7142 ( .A1(n8685), .A2(n5710), .ZN(n5557) );
  AOI22_X1 U7143 ( .A1(n5711), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n5182), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n5556) );
  OAI211_X1 U7144 ( .C1(n6628), .C2(n5558), .A(n5557), .B(n5556), .ZN(n8862)
         );
  INV_X1 U7145 ( .A(n8862), .ZN(n8699) );
  OR2_X1 U7146 ( .A1(n8937), .A2(n8699), .ZN(n5749) );
  INV_X1 U7147 ( .A(n5749), .ZN(n7734) );
  INV_X1 U7148 ( .A(n5559), .ZN(n5560) );
  MUX2_X1 U7149 ( .A(n7215), .B(n10416), .S(n6433), .Z(n5577) );
  XNOR2_X1 U7150 ( .A(n5577), .B(SI_21_), .ZN(n5563) );
  XNOR2_X1 U7151 ( .A(n5576), .B(n5563), .ZN(n7501) );
  NAND2_X1 U7152 ( .A1(n7501), .A2(n7579), .ZN(n5565) );
  OR2_X1 U7153 ( .A1(n7577), .A2(n7215), .ZN(n5564) );
  INV_X1 U7154 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5566) );
  NAND2_X1 U7155 ( .A1(n5568), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U7156 ( .A1(n5590), .A2(n5569), .ZN(n8671) );
  NAND2_X1 U7157 ( .A1(n8671), .A2(n5710), .ZN(n5575) );
  INV_X1 U7158 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U7159 ( .A1(n5711), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5571) );
  NAND2_X1 U7160 ( .A1(n5182), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5570) );
  OAI211_X1 U7161 ( .C1(n5572), .C2(n6628), .A(n5571), .B(n5570), .ZN(n5573)
         );
  INV_X1 U7162 ( .A(n5573), .ZN(n5574) );
  NAND2_X1 U7163 ( .A1(n8845), .A2(n8663), .ZN(n7733) );
  NAND2_X1 U7164 ( .A1(n8937), .A2(n8699), .ZN(n8668) );
  AND2_X1 U7165 ( .A1(n7733), .A2(n8668), .ZN(n7730) );
  INV_X1 U7166 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7297) );
  MUX2_X1 U7167 ( .A(n7297), .B(n7498), .S(n6433), .Z(n5580) );
  NAND2_X1 U7168 ( .A1(n5580), .A2(n10260), .ZN(n5598) );
  INV_X1 U7169 ( .A(n5580), .ZN(n5581) );
  NAND2_X1 U7170 ( .A1(n5581), .A2(SI_22_), .ZN(n5582) );
  NAND2_X1 U7171 ( .A1(n5598), .A2(n5582), .ZN(n5585) );
  INV_X1 U7172 ( .A(n5585), .ZN(n5583) );
  NAND2_X1 U7173 ( .A1(n5584), .A2(n5583), .ZN(n5599) );
  INV_X1 U7174 ( .A(n5584), .ZN(n5586) );
  NAND2_X1 U7175 ( .A1(n5586), .A2(n5585), .ZN(n5587) );
  NAND2_X1 U7176 ( .A1(n5599), .A2(n5587), .ZN(n7497) );
  NAND2_X1 U7177 ( .A1(n7497), .A2(n7579), .ZN(n5589) );
  OR2_X1 U7178 ( .A1(n7577), .A2(n7297), .ZN(n5588) );
  NAND2_X1 U7179 ( .A1(n5590), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5591) );
  NAND2_X1 U7180 ( .A1(n5610), .A2(n5591), .ZN(n8660) );
  NAND2_X1 U7181 ( .A1(n8660), .A2(n5710), .ZN(n5597) );
  INV_X1 U7182 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U7183 ( .A1(n5711), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U7184 ( .A1(n5182), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5592) );
  OAI211_X1 U7185 ( .C1(n5594), .C2(n6628), .A(n5593), .B(n5592), .ZN(n5595)
         );
  INV_X1 U7186 ( .A(n5595), .ZN(n5596) );
  INV_X1 U7187 ( .A(n8846), .ZN(n8039) );
  NAND2_X1 U7188 ( .A1(n8665), .A2(n8039), .ZN(n7742) );
  OR2_X1 U7189 ( .A1(n8665), .A2(n8039), .ZN(n5754) );
  INV_X1 U7190 ( .A(n5754), .ZN(n7744) );
  NAND2_X1 U7191 ( .A1(n5599), .A2(n5598), .ZN(n5606) );
  INV_X1 U7192 ( .A(n5606), .ZN(n5603) );
  MUX2_X1 U7193 ( .A(n7335), .B(n7494), .S(n6433), .Z(n5600) );
  INV_X1 U7194 ( .A(SI_23_), .ZN(n10473) );
  NAND2_X1 U7195 ( .A1(n5600), .A2(n10473), .ZN(n5617) );
  INV_X1 U7196 ( .A(n5600), .ZN(n5601) );
  NAND2_X1 U7197 ( .A1(n5601), .A2(SI_23_), .ZN(n5602) );
  NAND2_X1 U7198 ( .A1(n5617), .A2(n5602), .ZN(n5604) );
  NAND2_X1 U7199 ( .A1(n5603), .A2(n5604), .ZN(n5607) );
  INV_X1 U7200 ( .A(n5604), .ZN(n5605) );
  NAND2_X1 U7201 ( .A1(n5607), .A2(n5618), .ZN(n7493) );
  NAND2_X1 U7202 ( .A1(n7493), .A2(n7579), .ZN(n5609) );
  OR2_X1 U7203 ( .A1(n7577), .A2(n7335), .ZN(n5608) );
  NAND2_X1 U7204 ( .A1(n5610), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U7205 ( .A1(n5625), .A2(n5611), .ZN(n8653) );
  NAND2_X1 U7206 ( .A1(n8653), .A2(n5710), .ZN(n5616) );
  INV_X1 U7207 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8652) );
  NAND2_X1 U7208 ( .A1(n5711), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U7209 ( .A1(n5182), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5612) );
  OAI211_X1 U7210 ( .C1(n8652), .C2(n6628), .A(n5613), .B(n5612), .ZN(n5614)
         );
  INV_X1 U7211 ( .A(n5614), .ZN(n5615) );
  NOR2_X1 U7212 ( .A1(n8922), .A2(n8637), .ZN(n7738) );
  INV_X1 U7213 ( .A(n7738), .ZN(n7746) );
  INV_X1 U7214 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7560) );
  INV_X1 U7215 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7491) );
  MUX2_X1 U7216 ( .A(n7560), .B(n7491), .S(n6433), .Z(n5619) );
  NAND2_X1 U7217 ( .A1(n5619), .A2(n10293), .ZN(n5636) );
  INV_X1 U7218 ( .A(n5619), .ZN(n5620) );
  NAND2_X1 U7219 ( .A1(n5620), .A2(SI_24_), .ZN(n5621) );
  NAND2_X1 U7220 ( .A1(n7490), .A2(n7579), .ZN(n5623) );
  OR2_X1 U7221 ( .A1(n7577), .A2(n7560), .ZN(n5622) );
  NAND2_X1 U7222 ( .A1(n5625), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U7223 ( .A1(n5644), .A2(n5626), .ZN(n8639) );
  NAND2_X1 U7224 ( .A1(n8639), .A2(n5710), .ZN(n5632) );
  INV_X1 U7225 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n5629) );
  NAND2_X1 U7226 ( .A1(n5182), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5628) );
  NAND2_X1 U7227 ( .A1(n5711), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5627) );
  OAI211_X1 U7228 ( .C1(n5629), .C2(n6628), .A(n5628), .B(n5627), .ZN(n5630)
         );
  INV_X1 U7229 ( .A(n5630), .ZN(n5631) );
  NAND2_X1 U7230 ( .A1(n8376), .A2(n8826), .ZN(n7747) );
  NAND2_X1 U7231 ( .A1(n8922), .A2(n8637), .ZN(n8640) );
  NAND2_X1 U7232 ( .A1(n7747), .A2(n8640), .ZN(n7750) );
  INV_X1 U7233 ( .A(n7750), .ZN(n5633) );
  NAND2_X1 U7234 ( .A1(n8916), .A2(n8650), .ZN(n7749) );
  INV_X1 U7235 ( .A(n7749), .ZN(n7586) );
  INV_X1 U7236 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7556) );
  INV_X1 U7237 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10489) );
  MUX2_X1 U7238 ( .A(n7556), .B(n10489), .S(n6433), .Z(n5637) );
  INV_X1 U7239 ( .A(SI_25_), .ZN(n10243) );
  NAND2_X1 U7240 ( .A1(n5637), .A2(n10243), .ZN(n5653) );
  INV_X1 U7241 ( .A(n5637), .ZN(n5638) );
  NAND2_X1 U7242 ( .A1(n5638), .A2(SI_25_), .ZN(n5639) );
  XNOR2_X1 U7243 ( .A(n5652), .B(n5651), .ZN(n7555) );
  NAND2_X1 U7244 ( .A1(n7555), .A2(n7579), .ZN(n5641) );
  OR2_X1 U7245 ( .A1(n7577), .A2(n7556), .ZN(n5640) );
  INV_X1 U7246 ( .A(n5644), .ZN(n5643) );
  INV_X1 U7247 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U7248 ( .A1(n5643), .A2(n5642), .ZN(n5660) );
  NAND2_X1 U7249 ( .A1(n5644), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U7250 ( .A1(n5660), .A2(n5645), .ZN(n8625) );
  NAND2_X1 U7251 ( .A1(n8625), .A2(n5710), .ZN(n5650) );
  INV_X1 U7252 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8629) );
  NAND2_X1 U7253 ( .A1(n5182), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5647) );
  NAND2_X1 U7254 ( .A1(n5711), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5646) );
  OAI211_X1 U7255 ( .C1(n8629), .C2(n6628), .A(n5647), .B(n5646), .ZN(n5648)
         );
  INV_X1 U7256 ( .A(n5648), .ZN(n5649) );
  NOR2_X1 U7257 ( .A1(n8830), .A2(n8636), .ZN(n7754) );
  INV_X1 U7258 ( .A(n7754), .ZN(n5759) );
  NAND2_X1 U7259 ( .A1(n5652), .A2(n5651), .ZN(n5654) );
  NAND2_X1 U7260 ( .A1(n5654), .A2(n5653), .ZN(n5669) );
  INV_X1 U7261 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8992) );
  INV_X1 U7262 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7559) );
  MUX2_X1 U7263 ( .A(n8992), .B(n7559), .S(n6433), .Z(n5655) );
  INV_X1 U7264 ( .A(SI_26_), .ZN(n10419) );
  NAND2_X1 U7265 ( .A1(n5655), .A2(n10419), .ZN(n5670) );
  INV_X1 U7266 ( .A(n5655), .ZN(n5656) );
  NAND2_X1 U7267 ( .A1(n5656), .A2(SI_26_), .ZN(n5657) );
  XNOR2_X1 U7268 ( .A(n5669), .B(n5668), .ZN(n7557) );
  NAND2_X1 U7269 ( .A1(n7557), .A2(n7579), .ZN(n5659) );
  OR2_X1 U7270 ( .A1(n7577), .A2(n8992), .ZN(n5658) );
  OR2_X2 U7271 ( .A1(n5660), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5680) );
  NAND2_X1 U7272 ( .A1(n5660), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7273 ( .A1(n5680), .A2(n5661), .ZN(n8617) );
  NAND2_X1 U7274 ( .A1(n8617), .A2(n5710), .ZN(n5666) );
  INV_X1 U7275 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8616) );
  NAND2_X1 U7276 ( .A1(n5711), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U7277 ( .A1(n5182), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5662) );
  OAI211_X1 U7278 ( .C1(n8616), .C2(n6628), .A(n5663), .B(n5662), .ZN(n5664)
         );
  INV_X1 U7279 ( .A(n5664), .ZN(n5665) );
  INV_X1 U7280 ( .A(n7757), .ZN(n5667) );
  NAND2_X1 U7281 ( .A1(n8907), .A2(n8827), .ZN(n7758) );
  NAND2_X1 U7282 ( .A1(n5669), .A2(n5668), .ZN(n5671) );
  INV_X1 U7283 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5675) );
  INV_X1 U7284 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10190) );
  MUX2_X1 U7285 ( .A(n5675), .B(n10190), .S(n6433), .Z(n5672) );
  NAND2_X1 U7286 ( .A1(n5672), .A2(n10406), .ZN(n5690) );
  INV_X1 U7287 ( .A(n5672), .ZN(n5673) );
  NAND2_X1 U7288 ( .A1(n5673), .A2(SI_27_), .ZN(n5674) );
  NAND2_X1 U7289 ( .A1(n8986), .A2(n7579), .ZN(n5677) );
  OR2_X1 U7290 ( .A1(n7577), .A2(n5675), .ZN(n5676) );
  INV_X1 U7291 ( .A(n5680), .ZN(n5679) );
  INV_X1 U7292 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U7293 ( .A1(n5679), .A2(n5678), .ZN(n5694) );
  NAND2_X1 U7294 ( .A1(n5680), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5681) );
  NAND2_X1 U7295 ( .A1(n5694), .A2(n5681), .ZN(n8603) );
  NAND2_X1 U7296 ( .A1(n8603), .A2(n5710), .ZN(n5687) );
  INV_X1 U7297 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U7298 ( .A1(n5711), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U7299 ( .A1(n5182), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5682) );
  OAI211_X1 U7300 ( .C1(n5684), .C2(n5214), .A(n5683), .B(n5682), .ZN(n5685)
         );
  INV_X1 U7301 ( .A(n5685), .ZN(n5686) );
  NAND2_X1 U7302 ( .A1(n8607), .A2(n8614), .ZN(n5763) );
  NAND2_X1 U7303 ( .A1(n7622), .A2(n5763), .ZN(n8600) );
  INV_X1 U7304 ( .A(n8614), .ZN(n8590) );
  MUX2_X1 U7305 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6433), .Z(n5705) );
  INV_X1 U7306 ( .A(SI_28_), .ZN(n5706) );
  XNOR2_X1 U7307 ( .A(n5705), .B(n5706), .ZN(n5703) );
  NAND2_X1 U7308 ( .A1(n8308), .A2(n7579), .ZN(n5693) );
  INV_X1 U7309 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5691) );
  OR2_X1 U7310 ( .A1(n7577), .A2(n5691), .ZN(n5692) );
  NAND2_X1 U7311 ( .A1(n5694), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5695) );
  NAND2_X1 U7312 ( .A1(n5709), .A2(n5695), .ZN(n8595) );
  NAND2_X1 U7313 ( .A1(n8595), .A2(n5710), .ZN(n5700) );
  INV_X1 U7314 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8594) );
  NAND2_X1 U7315 ( .A1(n5711), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U7316 ( .A1(n5182), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5696) );
  OAI211_X1 U7317 ( .C1(n8594), .C2(n5214), .A(n5697), .B(n5696), .ZN(n5698)
         );
  INV_X1 U7318 ( .A(n5698), .ZN(n5699) );
  XNOR2_X2 U7319 ( .A(n8898), .B(n8602), .ZN(n8586) );
  NAND2_X1 U7320 ( .A1(n8587), .A2(n8586), .ZN(n5702) );
  INV_X1 U7321 ( .A(n8898), .ZN(n7621) );
  INV_X1 U7322 ( .A(n5705), .ZN(n5707) );
  INV_X1 U7323 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7481) );
  INV_X1 U7324 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8286) );
  MUX2_X1 U7325 ( .A(n7481), .B(n8286), .S(n7468), .Z(n7456) );
  NOR2_X1 U7326 ( .A1(n7577), .A2(n8286), .ZN(n5708) );
  NAND2_X1 U7327 ( .A1(n7796), .A2(n5710), .ZN(n6632) );
  INV_X1 U7328 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n5714) );
  NAND2_X1 U7329 ( .A1(n5182), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5713) );
  NAND2_X1 U7330 ( .A1(n5711), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5712) );
  OAI211_X1 U7331 ( .C1(n5714), .C2(n6628), .A(n5713), .B(n5712), .ZN(n5715)
         );
  INV_X1 U7332 ( .A(n5715), .ZN(n5716) );
  INV_X1 U7333 ( .A(n8591), .ZN(n6635) );
  AND2_X1 U7334 ( .A1(n7619), .A2(n6635), .ZN(n7766) );
  INV_X1 U7335 ( .A(n7766), .ZN(n7573) );
  INV_X1 U7336 ( .A(n7619), .ZN(n8581) );
  INV_X1 U7337 ( .A(n7773), .ZN(n5717) );
  XNOR2_X1 U7338 ( .A(n5718), .B(n7613), .ZN(n8582) );
  INV_X1 U7339 ( .A(n8602), .ZN(n8816) );
  INV_X1 U7340 ( .A(n5719), .ZN(n7786) );
  XNOR2_X1 U7341 ( .A(n7786), .B(n6154), .ZN(n5909) );
  NAND2_X2 U7342 ( .A1(n7789), .A2(n7626), .ZN(n7768) );
  NOR2_X1 U7343 ( .A1(n8816), .A2(n10027), .ZN(n5777) );
  NAND2_X1 U7344 ( .A1(n5191), .A2(n8796), .ZN(n8800) );
  OR2_X1 U7345 ( .A1(n5870), .A2(n5868), .ZN(n5722) );
  NAND2_X1 U7346 ( .A1(n6774), .A2(n7590), .ZN(n5724) );
  OR2_X1 U7347 ( .A1(n9998), .A2(n5873), .ZN(n5723) );
  NAND2_X1 U7348 ( .A1(n5724), .A2(n5723), .ZN(n6919) );
  NAND2_X1 U7349 ( .A1(n6919), .A2(n6920), .ZN(n5726) );
  INV_X1 U7350 ( .A(n9997), .ZN(n6296) );
  NAND2_X1 U7351 ( .A1(n6936), .A2(n6296), .ZN(n5725) );
  NAND2_X1 U7352 ( .A1(n5726), .A2(n5725), .ZN(n6939) );
  INV_X1 U7353 ( .A(n7642), .ZN(n7591) );
  NAND2_X1 U7354 ( .A1(n6939), .A2(n7591), .ZN(n5728) );
  INV_X1 U7355 ( .A(n10007), .ZN(n6935) );
  NAND2_X1 U7356 ( .A1(n10001), .A2(n6935), .ZN(n5727) );
  NAND2_X1 U7357 ( .A1(n5728), .A2(n5727), .ZN(n6414) );
  NOR2_X1 U7358 ( .A1(n8441), .A2(n6427), .ZN(n5730) );
  NAND2_X1 U7359 ( .A1(n8441), .A2(n6427), .ZN(n5729) );
  OR2_X1 U7360 ( .A1(n10021), .A2(n8440), .ZN(n6755) );
  NAND2_X1 U7361 ( .A1(n6757), .A2(n6755), .ZN(n6999) );
  NAND2_X1 U7362 ( .A1(n10021), .A2(n8440), .ZN(n6998) );
  NAND2_X1 U7363 ( .A1(n10030), .A2(n8439), .ZN(n5731) );
  AND2_X1 U7364 ( .A1(n6998), .A2(n5731), .ZN(n5732) );
  INV_X1 U7365 ( .A(n6789), .ZN(n10037) );
  NAND2_X1 U7366 ( .A1(n10045), .A2(n8438), .ZN(n5734) );
  OR2_X1 U7367 ( .A1(n10059), .A2(n10041), .ZN(n5736) );
  NAND2_X1 U7368 ( .A1(n7190), .A2(n8437), .ZN(n7166) );
  OR2_X1 U7369 ( .A1(n7190), .A2(n8437), .ZN(n7167) );
  OR2_X1 U7370 ( .A1(n8971), .A2(n8763), .ZN(n7589) );
  NAND2_X1 U7371 ( .A1(n8772), .A2(n7589), .ZN(n5737) );
  NAND2_X1 U7372 ( .A1(n8971), .A2(n8763), .ZN(n7588) );
  AND2_X1 U7373 ( .A1(n8964), .A2(n8774), .ZN(n5738) );
  NOR2_X1 U7374 ( .A1(n8958), .A2(n8764), .ZN(n5739) );
  NAND2_X1 U7375 ( .A1(n5740), .A2(n7625), .ZN(n8737) );
  NAND2_X1 U7376 ( .A1(n5741), .A2(n8752), .ZN(n5742) );
  NAND2_X1 U7377 ( .A1(n5743), .A2(n5742), .ZN(n8724) );
  NAND2_X1 U7378 ( .A1(n8724), .A2(n8725), .ZN(n5745) );
  NAND2_X1 U7379 ( .A1(n8733), .A2(n8740), .ZN(n5744) );
  NAND2_X1 U7380 ( .A1(n5745), .A2(n5744), .ZN(n8707) );
  INV_X1 U7381 ( .A(n8707), .ZN(n5746) );
  OR2_X1 U7382 ( .A1(n8873), .A2(n8694), .ZN(n5747) );
  NAND2_X1 U7383 ( .A1(n8863), .A2(n8855), .ZN(n5748) );
  NAND2_X1 U7384 ( .A1(n8693), .A2(n5748), .ZN(n8682) );
  OR2_X1 U7385 ( .A1(n8937), .A2(n8862), .ZN(n5751) );
  NAND2_X1 U7386 ( .A1(n7740), .A2(n7733), .ZN(n8676) );
  OR2_X1 U7387 ( .A1(n8845), .A2(n8856), .ZN(n5752) );
  NAND2_X1 U7388 ( .A1(n5753), .A2(n5752), .ZN(n8658) );
  OR2_X1 U7389 ( .A1(n8665), .A2(n8846), .ZN(n5755) );
  NOR2_X1 U7390 ( .A1(n8922), .A2(n8838), .ZN(n5756) );
  NAND2_X1 U7391 ( .A1(n8922), .A2(n8838), .ZN(n5757) );
  AND2_X1 U7392 ( .A1(n8376), .A2(n8650), .ZN(n5758) );
  OAI22_X1 U7393 ( .A1(n8634), .A2(n5758), .B1(n8650), .B2(n8376), .ZN(n8623)
         );
  NAND2_X1 U7394 ( .A1(n8623), .A2(n8620), .ZN(n5761) );
  OR2_X1 U7395 ( .A1(n8830), .A2(n8613), .ZN(n5760) );
  NAND2_X1 U7396 ( .A1(n8907), .A2(n8631), .ZN(n5762) );
  INV_X1 U7397 ( .A(n5763), .ZN(n5764) );
  NOR2_X1 U7398 ( .A1(n8898), .A2(n8602), .ZN(n5765) );
  OAI22_X1 U7399 ( .A1(n8589), .A2(n5765), .B1(n8816), .B2(n7621), .ZN(n5766)
         );
  OR2_X1 U7400 ( .A1(n5139), .A2(n7296), .ZN(n5768) );
  NAND2_X1 U7401 ( .A1(n7626), .A2(n5824), .ZN(n5767) );
  INV_X1 U7402 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n5772) );
  NAND2_X1 U7403 ( .A1(n5182), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5771) );
  INV_X1 U7404 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n5769) );
  OR2_X1 U7405 ( .A1(n6625), .A2(n5769), .ZN(n5770) );
  OAI211_X1 U7406 ( .C1(n5772), .C2(n5214), .A(n5771), .B(n5770), .ZN(n5773)
         );
  INV_X1 U7407 ( .A(n5773), .ZN(n5774) );
  NAND2_X1 U7408 ( .A1(n6632), .A2(n5774), .ZN(n8436) );
  INV_X1 U7409 ( .A(n8436), .ZN(n5776) );
  AND2_X1 U7410 ( .A1(n5861), .A2(P2_B_REG_SCAN_IN), .ZN(n5775) );
  OR2_X1 U7411 ( .A1(n10025), .A2(n5775), .ZN(n7793) );
  NAND2_X1 U7412 ( .A1(n5801), .A2(n5802), .ZN(n5779) );
  XNOR2_X1 U7413 ( .A(n5791), .B(P2_B_REG_SCAN_IN), .ZN(n5785) );
  NAND2_X1 U7414 ( .A1(n5781), .A2(n5780), .ZN(n5782) );
  NAND2_X1 U7415 ( .A1(n5785), .A2(n5794), .ZN(n5790) );
  NAND2_X1 U7416 ( .A1(n5786), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5787) );
  MUX2_X1 U7417 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5787), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5789) );
  NAND2_X1 U7418 ( .A1(n5790), .A2(n5798), .ZN(n5793) );
  NAND2_X1 U7419 ( .A1(n5791), .A2(n8993), .ZN(n6078) );
  NAND2_X1 U7420 ( .A1(n5792), .A2(n6078), .ZN(n5864) );
  OR2_X1 U7421 ( .A1(n5793), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U7422 ( .A1(n5794), .A2(n8993), .ZN(n6081) );
  NAND2_X1 U7423 ( .A1(n5795), .A2(n6081), .ZN(n5827) );
  NOR2_X1 U7424 ( .A1(n10055), .A2(n7626), .ZN(n5914) );
  INV_X1 U7425 ( .A(n5914), .ZN(n5796) );
  AND2_X1 U7426 ( .A1(n5897), .A2(n5796), .ZN(n5818) );
  INV_X1 U7427 ( .A(n5794), .ZN(n5800) );
  INV_X1 U7428 ( .A(n5791), .ZN(n5797) );
  NOR4_X1 U7429 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n5811) );
  OR4_X1 U7430 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5808) );
  NOR4_X1 U7431 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5806) );
  NOR4_X1 U7432 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5805) );
  NOR4_X1 U7433 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5804) );
  NOR4_X1 U7434 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5803) );
  NAND4_X1 U7435 ( .A1(n5806), .A2(n5805), .A3(n5804), .A4(n5803), .ZN(n5807)
         );
  NOR4_X1 U7436 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        n5808), .A4(n5807), .ZN(n5810) );
  NOR4_X1 U7437 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5809) );
  NAND3_X1 U7438 ( .A1(n5811), .A2(n5810), .A3(n5809), .ZN(n5892) );
  NAND2_X1 U7439 ( .A1(n5867), .A2(n7775), .ZN(n5898) );
  OR2_X1 U7440 ( .A1(n5812), .A2(n7782), .ZN(n5813) );
  NAND2_X1 U7441 ( .A1(n5813), .A2(n7768), .ZN(n5814) );
  OR2_X1 U7442 ( .A1(n5864), .A2(n5814), .ZN(n5817) );
  INV_X1 U7443 ( .A(n5814), .ZN(n5815) );
  NAND2_X1 U7444 ( .A1(n10087), .A2(n10060), .ZN(n8853) );
  INV_X1 U7445 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5819) );
  INV_X1 U7446 ( .A(n5821), .ZN(n5822) );
  OAI21_X1 U7447 ( .B1(n5834), .B2(n10085), .A(n5822), .ZN(P2_U3488) );
  INV_X1 U7448 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5835) );
  INV_X1 U7449 ( .A(n5828), .ZN(n5823) );
  NAND2_X1 U7450 ( .A1(n7618), .A2(n5824), .ZN(n5865) );
  NOR2_X1 U7451 ( .A1(n7296), .A2(n5865), .ZN(n5825) );
  AND2_X1 U7452 ( .A1(n7784), .A2(n5825), .ZN(n5894) );
  NAND2_X1 U7453 ( .A1(n5888), .A2(n5906), .ZN(n5826) );
  NAND2_X1 U7454 ( .A1(n5911), .A2(n5826), .ZN(n5833) );
  NAND2_X1 U7455 ( .A1(n5864), .A2(n5827), .ZN(n6419) );
  INV_X1 U7456 ( .A(n6419), .ZN(n5829) );
  NAND2_X1 U7457 ( .A1(n5829), .A2(n5828), .ZN(n5907) );
  NAND2_X1 U7458 ( .A1(n6412), .A2(n10060), .ZN(n8778) );
  AND2_X1 U7459 ( .A1(n7768), .A2(n10062), .ZN(n5830) );
  NAND2_X1 U7460 ( .A1(n5888), .A2(n5830), .ZN(n5886) );
  NAND2_X1 U7461 ( .A1(n8778), .A2(n5886), .ZN(n5895) );
  INV_X1 U7462 ( .A(n5895), .ZN(n5831) );
  NAND2_X1 U7463 ( .A1(n5836), .A2(n5111), .ZN(P2_U3456) );
  NAND2_X1 U7464 ( .A1(n5840), .A2(n6092), .ZN(n6115) );
  NAND2_X1 U7465 ( .A1(n5946), .A2(n5850), .ZN(n5852) );
  OR2_X1 U7466 ( .A1(n5946), .A2(n5850), .ZN(n5851) );
  INV_X1 U7467 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U7468 ( .A1(n5936), .A2(n5855), .ZN(n5856) );
  NAND2_X1 U7469 ( .A1(n5953), .A2(n10232), .ZN(n5857) );
  NAND2_X1 U7470 ( .A1(n6167), .A2(n7768), .ZN(n5860) );
  NAND2_X1 U7471 ( .A1(n5860), .A2(n6166), .ZN(n6169) );
  NAND2_X1 U7472 ( .A1(n6169), .A2(n5861), .ZN(n5862) );
  NAND2_X1 U7473 ( .A1(n5862), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NOR2_X4 U7474 ( .A1(n6167), .A2(n5863), .ZN(P2_U3893) );
  XNOR2_X1 U7475 ( .A(n5868), .B(n5874), .ZN(n5871) );
  NAND2_X1 U7476 ( .A1(n5871), .A2(n5005), .ZN(n5872) );
  INV_X1 U7477 ( .A(n8048), .ZN(n5869) );
  OAI21_X1 U7478 ( .B1(n5869), .B2(n5191), .A(n8787), .ZN(n6300) );
  XNOR2_X1 U7479 ( .A(n5871), .B(n5870), .ZN(n6301) );
  XNOR2_X1 U7480 ( .A(n5874), .B(n5873), .ZN(n5876) );
  XNOR2_X1 U7481 ( .A(n5876), .B(n9998), .ZN(n6316) );
  INV_X1 U7482 ( .A(n9998), .ZN(n5875) );
  NAND2_X1 U7483 ( .A1(n5876), .A2(n5875), .ZN(n5877) );
  INV_X1 U7484 ( .A(n6292), .ZN(n5879) );
  XNOR2_X1 U7485 ( .A(n8051), .B(n9997), .ZN(n5880) );
  XNOR2_X1 U7486 ( .A(n5880), .B(n6936), .ZN(n6293) );
  INV_X1 U7487 ( .A(n6293), .ZN(n5878) );
  NAND2_X1 U7488 ( .A1(n5879), .A2(n5878), .ZN(n6290) );
  INV_X1 U7489 ( .A(n5880), .ZN(n5881) );
  NAND2_X1 U7490 ( .A1(n5881), .A2(n10008), .ZN(n5882) );
  NAND2_X1 U7491 ( .A1(n6290), .A2(n5882), .ZN(n5885) );
  XNOR2_X1 U7492 ( .A(n8051), .B(n10007), .ZN(n6306) );
  XNOR2_X1 U7493 ( .A(n6306), .B(n10001), .ZN(n5884) );
  INV_X1 U7494 ( .A(n5884), .ZN(n5883) );
  NAND2_X1 U7495 ( .A1(n5885), .A2(n5884), .ZN(n5891) );
  INV_X1 U7496 ( .A(n5886), .ZN(n5887) );
  NAND2_X1 U7497 ( .A1(n5911), .A2(n5887), .ZN(n5890) );
  OR2_X1 U7498 ( .A1(n5907), .A2(n5888), .ZN(n5889) );
  AOI21_X1 U7499 ( .B1(n6308), .B2(n5891), .A(n8421), .ZN(n5920) );
  INV_X1 U7500 ( .A(n5793), .ZN(n5893) );
  AND2_X1 U7501 ( .A1(n5893), .A2(n5892), .ZN(n5896) );
  OR2_X1 U7502 ( .A1(n6419), .A2(n5896), .ZN(n5903) );
  NAND2_X1 U7503 ( .A1(n5903), .A2(n5894), .ZN(n5901) );
  AND2_X1 U7504 ( .A1(n6167), .A2(n6166), .ZN(n5900) );
  OAI21_X1 U7505 ( .B1(n5897), .B2(n5896), .A(n5895), .ZN(n5899) );
  NAND4_X1 U7506 ( .A1(n5901), .A2(n5900), .A3(n5899), .A4(n5898), .ZN(n5902)
         );
  NAND2_X1 U7507 ( .A1(n5902), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5905) );
  NOR2_X1 U7508 ( .A1(n5912), .A2(n5906), .ZN(n7787) );
  NAND2_X1 U7509 ( .A1(n5903), .A2(n7787), .ZN(n5904) );
  NOR2_X1 U7510 ( .A1(n8428), .A2(n6934), .ZN(n5919) );
  NOR2_X1 U7511 ( .A1(n5907), .A2(n5906), .ZN(n5910) );
  INV_X1 U7512 ( .A(n5909), .ZN(n5908) );
  NAND2_X1 U7513 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6284) );
  OAI21_X1 U7514 ( .B1(n8409), .B2(n6936), .A(n6284), .ZN(n5918) );
  NAND2_X1 U7515 ( .A1(n5910), .A2(n5909), .ZN(n8427) );
  INV_X1 U7516 ( .A(n8441), .ZN(n10011) );
  NAND2_X1 U7517 ( .A1(n5911), .A2(n10060), .ZN(n5915) );
  INV_X1 U7518 ( .A(n5912), .ZN(n5913) );
  NAND2_X1 U7519 ( .A1(n8419), .A2(n10007), .ZN(n5916) );
  OAI21_X1 U7520 ( .B1(n8427), .B2(n10011), .A(n5916), .ZN(n5917) );
  OR4_X1 U7521 ( .A1(n5920), .A2(n5919), .A3(n5918), .A4(n5917), .ZN(P2_U3170)
         );
  NOR2_X1 U7522 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5921) );
  NAND2_X1 U7523 ( .A1(n4513), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5935) );
  INV_X1 U7524 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6911) );
  OR2_X1 U7525 ( .A1(n6551), .A2(n6911), .ZN(n5934) );
  NAND2_X4 U7526 ( .A1(n5929), .A2(n7550), .ZN(n7981) );
  INV_X1 U7527 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5930) );
  OR2_X1 U7528 ( .A1(n7981), .A2(n5930), .ZN(n5933) );
  INV_X1 U7529 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5931) );
  OR2_X1 U7530 ( .A1(n7933), .A2(n5931), .ZN(n5932) );
  NAND2_X1 U7531 ( .A1(n5937), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5939) );
  AND2_X1 U7532 ( .A1(n8075), .A2(n6477), .ZN(n5940) );
  NAND2_X1 U7533 ( .A1(n9178), .A2(n6541), .ZN(n5960) );
  NOR2_X1 U7534 ( .A1(n7468), .A2(n10450), .ZN(n5942) );
  XNOR2_X1 U7535 ( .A(n5942), .B(n5941), .ZN(n9796) );
  INV_X1 U7536 ( .A(n5943), .ZN(n5944) );
  NAND2_X1 U7537 ( .A1(n5944), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7538 ( .A1(n5946), .A2(n5945), .ZN(n5950) );
  AND2_X1 U7539 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5947) );
  MUX2_X1 U7540 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9796), .S(n7229), .Z(n6664) );
  NAND2_X1 U7541 ( .A1(n5951), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5952) );
  XNOR2_X2 U7542 ( .A(n5952), .B(n10261), .ZN(n9343) );
  NAND2_X1 U7543 ( .A1(n8075), .A2(n8268), .ZN(n8278) );
  INV_X1 U7544 ( .A(n6469), .ZN(n6398) );
  INV_X2 U7545 ( .A(n9343), .ZN(n9327) );
  AND2_X1 U7546 ( .A1(n6477), .A2(n9327), .ZN(n5955) );
  NAND2_X1 U7547 ( .A1(n8075), .A2(n5955), .ZN(n7063) );
  OAI21_X1 U7548 ( .B1(n5954), .B2(n6398), .A(n7063), .ZN(n5956) );
  INV_X1 U7549 ( .A(n5956), .ZN(n5957) );
  NAND2_X1 U7550 ( .A1(n5960), .A2(n5959), .ZN(n6430) );
  INV_X1 U7551 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6105) );
  NOR2_X1 U7552 ( .A1(n5958), .A2(n6105), .ZN(n5961) );
  INV_X1 U7553 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7554 ( .A1(n9178), .A2(n7959), .ZN(n5963) );
  NAND2_X1 U7555 ( .A1(n6664), .A2(n6541), .ZN(n5962) );
  OAI211_X1 U7556 ( .C1(n5958), .C2(n5981), .A(n5963), .B(n5962), .ZN(n5964)
         );
  OAI21_X1 U7557 ( .B1(n5965), .B2(n5964), .A(n6432), .ZN(n6498) );
  NAND3_X1 U7558 ( .A1(n6498), .A2(n9793), .A3(n6663), .ZN(n5971) );
  OAI21_X1 U7559 ( .B1(n9793), .B2(P1_REG2_REG_0__SCAN_IN), .A(n6663), .ZN(
        n6104) );
  NAND2_X1 U7560 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n7567) );
  INV_X1 U7561 ( .A(n7567), .ZN(n5969) );
  AOI22_X1 U7562 ( .A1(n5981), .A2(n6104), .B1(n5110), .B2(n5969), .ZN(n5970)
         );
  AND3_X1 U7563 ( .A1(n5971), .A2(P1_U3973), .A3(n5970), .ZN(n6009) );
  INV_X1 U7564 ( .A(n7572), .ZN(n5982) );
  NOR2_X1 U7565 ( .A1(n7566), .A2(n7567), .ZN(n7565) );
  AOI21_X1 U7566 ( .B1(n5982), .B2(P1_REG2_REG_1__SCAN_IN), .A(n7565), .ZN(
        n5980) );
  NOR2_X1 U7567 ( .A1(n5972), .A2(n5854), .ZN(n5973) );
  MUX2_X1 U7568 ( .A(n5854), .B(n5973), .S(P1_IR_REG_2__SCAN_IN), .Z(n5974) );
  INV_X1 U7569 ( .A(n5974), .ZN(n5976) );
  NAND2_X1 U7570 ( .A1(n5976), .A2(n5975), .ZN(n6444) );
  XOR2_X1 U7571 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6444), .Z(n5979) );
  NOR2_X1 U7572 ( .A1(n5980), .A2(n5979), .ZN(n6001) );
  NAND2_X1 U7573 ( .A1(n5954), .A2(n8075), .ZN(n6470) );
  OR2_X1 U7574 ( .A1(n6480), .A2(n6470), .ZN(n5977) );
  AND2_X1 U7575 ( .A1(n7229), .A2(n5977), .ZN(n5985) );
  NAND2_X1 U7576 ( .A1(n6480), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8285) );
  NAND2_X1 U7577 ( .A1(n6097), .A2(n8285), .ZN(n5978) );
  AOI211_X1 U7578 ( .C1(n5980), .C2(n5979), .A(n6001), .B(n9259), .ZN(n5990)
         );
  NOR3_X1 U7579 ( .A1(n7563), .A2(n6105), .A3(n5981), .ZN(n7562) );
  AOI21_X1 U7580 ( .B1(n5982), .B2(P1_REG1_REG_1__SCAN_IN), .A(n7562), .ZN(
        n5984) );
  XOR2_X1 U7581 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6444), .Z(n5983) );
  NOR2_X1 U7582 ( .A1(n5984), .A2(n5983), .ZN(n5993) );
  AOI211_X1 U7583 ( .C1(n5984), .C2(n5983), .A(n5993), .B(n9254), .ZN(n5989)
         );
  INV_X1 U7584 ( .A(n5985), .ZN(n5986) );
  OAI211_X2 U7585 ( .C1(n5958), .C2(n6480), .A(n5986), .B(P1_STATE_REG_SCAN_IN), .ZN(n9234) );
  INV_X1 U7586 ( .A(n9234), .ZN(n9261) );
  AOI22_X1 U7587 ( .A1(n9261), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n5987) );
  OAI21_X1 U7588 ( .B1(n6444), .B2(n9258), .A(n5987), .ZN(n5988) );
  OR4_X1 U7589 ( .A1(n6009), .A2(n5990), .A3(n5989), .A4(n5988), .ZN(P1_U3245)
         );
  NAND2_X1 U7590 ( .A1(n5975), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5992) );
  INV_X1 U7591 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5991) );
  XNOR2_X1 U7592 ( .A(n5992), .B(n5991), .ZN(n6535) );
  INV_X1 U7593 ( .A(n6535), .ZN(n6217) );
  INV_X1 U7594 ( .A(n6444), .ZN(n6002) );
  XOR2_X1 U7595 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6535), .Z(n6221) );
  NAND2_X1 U7596 ( .A1(n5994), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5995) );
  MUX2_X1 U7597 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5995), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5998) );
  INV_X1 U7598 ( .A(n5996), .ZN(n5997) );
  NAND2_X1 U7599 ( .A1(n5998), .A2(n5997), .ZN(n6547) );
  XOR2_X1 U7600 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6547), .Z(n5999) );
  AOI211_X1 U7601 ( .C1(n6000), .C2(n5999), .A(n6010), .B(n9254), .ZN(n6008)
         );
  AOI21_X1 U7602 ( .B1(n6002), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6001), .ZN(
        n6216) );
  XOR2_X1 U7603 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6535), .Z(n6215) );
  NOR2_X1 U7604 ( .A1(n6216), .A2(n6215), .ZN(n6214) );
  AOI21_X1 U7605 ( .B1(n6217), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6214), .ZN(
        n6004) );
  INV_X1 U7606 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7016) );
  XNOR2_X1 U7607 ( .A(n6547), .B(n7016), .ZN(n6003) );
  AOI211_X1 U7608 ( .C1(n6004), .C2(n6003), .A(n6014), .B(n9259), .ZN(n6007)
         );
  AND2_X1 U7609 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n6577) );
  AOI21_X1 U7610 ( .B1(n9261), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6577), .ZN(
        n6005) );
  OAI21_X1 U7611 ( .B1(n9258), .B2(n6547), .A(n6005), .ZN(n6006) );
  OR4_X1 U7612 ( .A1(n6009), .A2(n6008), .A3(n6007), .A4(n6006), .ZN(P1_U3247)
         );
  INV_X1 U7613 ( .A(n6547), .ZN(n6015) );
  AOI21_X1 U7614 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n6015), .A(n6010), .ZN(
        n6013) );
  OR2_X1 U7615 ( .A1(n5996), .A2(n5854), .ZN(n6011) );
  XNOR2_X1 U7616 ( .A(n6011), .B(n6024), .ZN(n6728) );
  XOR2_X1 U7617 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6728), .Z(n6012) );
  NOR2_X1 U7618 ( .A1(n6013), .A2(n6012), .ZN(n6023) );
  AOI211_X1 U7619 ( .C1(n6013), .C2(n6012), .A(n9254), .B(n6023), .ZN(n6022)
         );
  NOR2_X1 U7620 ( .A1(n9258), .A2(n6728), .ZN(n6021) );
  INV_X1 U7621 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7217) );
  XNOR2_X1 U7622 ( .A(n6728), .B(n7217), .ZN(n6016) );
  AOI211_X1 U7623 ( .C1(n6017), .C2(n6016), .A(n9259), .B(n6028), .ZN(n6020)
         );
  INV_X1 U7624 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7625 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9073) );
  OAI21_X1 U7626 ( .B1(n9234), .B2(n6018), .A(n9073), .ZN(n6019) );
  OR4_X1 U7627 ( .A1(n6022), .A2(n6021), .A3(n6020), .A4(n6019), .ZN(P1_U3248)
         );
  INV_X1 U7628 ( .A(n6728), .ZN(n6029) );
  AOI21_X1 U7629 ( .B1(n6029), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6023), .ZN(
        n6027) );
  AND2_X1 U7630 ( .A1(n5996), .A2(n6024), .ZN(n6025) );
  INV_X1 U7631 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6038) );
  XNOR2_X1 U7632 ( .A(n6039), .B(n6038), .ZN(n6850) );
  XOR2_X1 U7633 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6850), .Z(n6026) );
  NOR2_X1 U7634 ( .A1(n6027), .A2(n6026), .ZN(n6037) );
  AOI211_X1 U7635 ( .C1(n6027), .C2(n6026), .A(n9254), .B(n6037), .ZN(n6036)
         );
  NOR2_X1 U7636 ( .A1(n9258), .A2(n6850), .ZN(n6035) );
  INV_X1 U7637 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7081) );
  XNOR2_X1 U7638 ( .A(n6850), .B(n7081), .ZN(n6030) );
  NOR2_X1 U7639 ( .A1(n6031), .A2(n6030), .ZN(n6045) );
  AOI211_X1 U7640 ( .C1(n6031), .C2(n6030), .A(n9259), .B(n6045), .ZN(n6034)
         );
  INV_X1 U7641 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6032) );
  NAND2_X1 U7642 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6871) );
  OAI21_X1 U7643 ( .B1(n9234), .B2(n6032), .A(n6871), .ZN(n6033) );
  OR4_X1 U7644 ( .A1(n6036), .A2(n6035), .A3(n6034), .A4(n6033), .ZN(P1_U3249)
         );
  INV_X1 U7645 ( .A(n6850), .ZN(n6046) );
  AOI21_X1 U7646 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n6046), .A(n6037), .ZN(
        n6044) );
  NAND2_X1 U7647 ( .A1(n6039), .A2(n6038), .ZN(n6040) );
  NAND2_X1 U7648 ( .A1(n6040), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6042) );
  INV_X1 U7649 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6041) );
  XNOR2_X1 U7650 ( .A(n6042), .B(n6041), .ZN(n7028) );
  XOR2_X1 U7651 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n7028), .Z(n6043) );
  AOI211_X1 U7652 ( .C1(n6044), .C2(n6043), .A(n9254), .B(n6054), .ZN(n6053)
         );
  NOR2_X1 U7653 ( .A1(n9258), .A2(n7028), .ZN(n6052) );
  AOI21_X1 U7654 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6046), .A(n6045), .ZN(
        n6048) );
  INV_X1 U7655 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7099) );
  XNOR2_X1 U7656 ( .A(n7028), .B(n7099), .ZN(n6047) );
  AOI211_X1 U7657 ( .C1(n6048), .C2(n6047), .A(n9259), .B(n6060), .ZN(n6051)
         );
  INV_X1 U7658 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U7659 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7114) );
  OAI21_X1 U7660 ( .B1(n9234), .B2(n6049), .A(n7114), .ZN(n6050) );
  OR4_X1 U7661 ( .A1(n6053), .A2(n6052), .A3(n6051), .A4(n6050), .ZN(P1_U3250)
         );
  INV_X1 U7662 ( .A(n7028), .ZN(n6061) );
  NAND2_X1 U7663 ( .A1(n6055), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6057) );
  XNOR2_X1 U7664 ( .A(n6057), .B(n6056), .ZN(n7034) );
  XOR2_X1 U7665 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n7034), .Z(n6058) );
  AOI211_X1 U7666 ( .C1(n6059), .C2(n6058), .A(n9254), .B(n6194), .ZN(n6068)
         );
  NOR2_X1 U7667 ( .A1(n9258), .A2(n7034), .ZN(n6067) );
  INV_X1 U7668 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7066) );
  XNOR2_X1 U7669 ( .A(n7034), .B(n7066), .ZN(n6062) );
  AOI211_X1 U7670 ( .C1(n6063), .C2(n6062), .A(n9259), .B(n6201), .ZN(n6066)
         );
  INV_X1 U7671 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7672 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n7313) );
  OAI21_X1 U7673 ( .B1(n9234), .B2(n6064), .A(n7313), .ZN(n6065) );
  OR4_X1 U7674 ( .A1(n6068), .A2(n6067), .A3(n6066), .A4(n6065), .ZN(P1_U3251)
         );
  AND2_X1 U7675 ( .A1(n7468), .A2(P1_U3086), .ZN(n6931) );
  INV_X2 U7676 ( .A(n6931), .ZN(n6832) );
  NOR2_X1 U7677 ( .A1(n7468), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9790) );
  OAI222_X1 U7678 ( .A1(n6832), .A2(n5196), .B1(n7300), .B2(n6443), .C1(
        P1_U3086), .C2(n6444), .ZN(P1_U3353) );
  INV_X1 U7679 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6533) );
  OAI222_X1 U7680 ( .A1(n6832), .A2(n6533), .B1(n7300), .B2(n6534), .C1(
        P1_U3086), .C2(n6535), .ZN(P1_U3352) );
  OAI222_X1 U7681 ( .A1(n6832), .A2(n4965), .B1(n7300), .B2(n6434), .C1(
        P1_U3086), .C2(n7572), .ZN(P1_U3354) );
  AND2_X1 U7682 ( .A1(n7468), .A2(P2_U3151), .ZN(n8981) );
  INV_X2 U7683 ( .A(n8988), .ZN(n8991) );
  OAI222_X1 U7684 ( .A1(n8990), .A2(n6534), .B1(n6164), .B2(P2_U3151), .C1(
        n6069), .C2(n8991), .ZN(P2_U3292) );
  INV_X2 U7685 ( .A(n8981), .ZN(n8990) );
  OAI222_X1 U7686 ( .A1(n8990), .A2(n6443), .B1(n9880), .B2(P2_U3151), .C1(
        n5195), .C2(n8991), .ZN(P2_U3293) );
  OAI222_X1 U7687 ( .A1(n8990), .A2(n6434), .B1(n9860), .B2(P2_U3151), .C1(
        n6070), .C2(n8991), .ZN(P2_U3294) );
  OAI222_X1 U7688 ( .A1(n8990), .A2(n6545), .B1(n6289), .B2(P2_U3151), .C1(
        n6071), .C2(n8991), .ZN(P2_U3291) );
  OAI222_X1 U7689 ( .A1(P1_U3086), .A2(n6547), .B1(n7300), .B2(n6545), .C1(
        n4707), .C2(n6832), .ZN(P1_U3351) );
  OAI222_X1 U7690 ( .A1(n8990), .A2(n6727), .B1(n6261), .B2(P2_U3151), .C1(
        n6072), .C2(n8991), .ZN(P2_U3290) );
  INV_X1 U7691 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6726) );
  OAI222_X1 U7692 ( .A1(n6832), .A2(n6726), .B1(n7300), .B2(n6727), .C1(
        P1_U3086), .C2(n6728), .ZN(P1_U3350) );
  AND2_X1 U7693 ( .A1(n6073), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U7694 ( .A1(n6073), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U7695 ( .A1(n6073), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U7696 ( .A1(n6073), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U7697 ( .A1(n6073), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U7698 ( .A1(n6073), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U7699 ( .A1(n6073), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U7700 ( .A1(n6073), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U7701 ( .A1(n6073), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U7702 ( .A1(n6073), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U7703 ( .A1(n6073), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U7704 ( .A1(n6073), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U7705 ( .A1(n6073), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U7706 ( .A1(n6073), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  OAI222_X1 U7707 ( .A1(n8990), .A2(n6848), .B1(n6505), .B2(P2_U3151), .C1(
        n6074), .C2(n8991), .ZN(P2_U3289) );
  INV_X1 U7708 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6849) );
  OAI222_X1 U7709 ( .A1(P1_U3086), .A2(n6850), .B1(n7300), .B2(n6848), .C1(
        n6849), .C2(n6832), .ZN(P1_U3349) );
  INV_X1 U7710 ( .A(n6506), .ZN(n6816) );
  INV_X1 U7711 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6075) );
  OAI222_X1 U7712 ( .A1(n8990), .A2(n7026), .B1(n6816), .B2(P2_U3151), .C1(
        n6075), .C2(n8991), .ZN(P2_U3288) );
  INV_X1 U7713 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7027) );
  OAI222_X1 U7714 ( .A1(P1_U3086), .A2(n7028), .B1(n7300), .B2(n7026), .C1(
        n7027), .C2(n6832), .ZN(P1_U3348) );
  INV_X1 U7715 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6076) );
  INV_X1 U7716 ( .A(n7033), .ZN(n6077) );
  INV_X1 U7717 ( .A(n8450), .ZN(n6814) );
  OAI222_X1 U7718 ( .A1(n8991), .A2(n6076), .B1(n8990), .B2(n6077), .C1(
        P2_U3151), .C2(n6814), .ZN(P2_U3287) );
  INV_X1 U7719 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10478) );
  OAI222_X1 U7720 ( .A1(n7034), .A2(P1_U3086), .B1(n7300), .B2(n6077), .C1(
        n10478), .C2(n6832), .ZN(P1_U3347) );
  INV_X1 U7721 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6080) );
  INV_X1 U7722 ( .A(n6078), .ZN(n6079) );
  AOI22_X1 U7723 ( .A1(n6073), .A2(n6080), .B1(n6083), .B2(n6079), .ZN(
        P2_U3376) );
  INV_X1 U7724 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6084) );
  INV_X1 U7725 ( .A(n6081), .ZN(n6082) );
  AOI22_X1 U7726 ( .A1(n6073), .A2(n6084), .B1(n6083), .B2(n6082), .ZN(
        P2_U3377) );
  AND2_X1 U7727 ( .A1(n6073), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U7728 ( .A1(n6073), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U7729 ( .A1(n6073), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U7730 ( .A1(n6073), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U7731 ( .A1(n6073), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U7732 ( .A1(n6073), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U7733 ( .A1(n6073), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U7734 ( .A1(n6073), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U7735 ( .A1(n6073), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U7736 ( .A1(n6073), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U7737 ( .A1(n6073), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U7738 ( .A1(n6073), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U7739 ( .A1(n6073), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U7740 ( .A1(n6073), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U7741 ( .A1(n6073), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U7742 ( .A1(n6073), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  OR2_X1 U7743 ( .A1(n6055), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7744 ( .A1(n6116), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6093) );
  XNOR2_X1 U7745 ( .A(n6093), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7253) );
  AOI22_X1 U7746 ( .A1(n7253), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n6931), .ZN(n6085) );
  OAI21_X1 U7747 ( .B1(n7252), .B2(n7300), .A(n6085), .ZN(P1_U3345) );
  INV_X1 U7748 ( .A(n7228), .ZN(n6091) );
  NAND2_X1 U7749 ( .A1(n6086), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6087) );
  XNOR2_X1 U7750 ( .A(n6087), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7230) );
  AOI22_X1 U7751 ( .A1(n7230), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n6931), .ZN(n6088) );
  OAI21_X1 U7752 ( .B1(n6091), .B2(n7300), .A(n6088), .ZN(P1_U3346) );
  INV_X1 U7753 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6089) );
  OAI222_X1 U7754 ( .A1(n8990), .A2(n7252), .B1(n7140), .B2(P2_U3151), .C1(
        n6089), .C2(n8991), .ZN(P2_U3285) );
  INV_X1 U7755 ( .A(n6892), .ZN(n6882) );
  OAI222_X1 U7756 ( .A1(n8990), .A2(n6091), .B1(n6882), .B2(P2_U3151), .C1(
        n6090), .C2(n8991), .ZN(P2_U3286) );
  INV_X1 U7757 ( .A(n7339), .ZN(n6111) );
  NAND2_X1 U7758 ( .A1(n6093), .A2(n10490), .ZN(n6094) );
  NAND2_X1 U7759 ( .A1(n6094), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6095) );
  XNOR2_X1 U7760 ( .A(n6095), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7340) );
  AOI22_X1 U7761 ( .A1(n7340), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n6931), .ZN(n6096) );
  OAI21_X1 U7762 ( .B1(n6111), .B2(n7300), .A(n6096), .ZN(P1_U3344) );
  NAND2_X1 U7763 ( .A1(n9794), .A2(P1_B_REG_SCAN_IN), .ZN(n6099) );
  INV_X1 U7764 ( .A(n7452), .ZN(n6098) );
  MUX2_X1 U7765 ( .A(n6099), .B(P1_B_REG_SCAN_IN), .S(n6098), .Z(n6101) );
  INV_X1 U7766 ( .A(n7558), .ZN(n6100) );
  INV_X1 U7767 ( .A(n6395), .ZN(n6102) );
  INV_X1 U7768 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10433) );
  NAND2_X1 U7769 ( .A1(n7558), .A2(n7452), .ZN(n6396) );
  INV_X1 U7770 ( .A(n6396), .ZN(n6103) );
  AOI22_X1 U7771 ( .A1(n9797), .A2(n10433), .B1(n8271), .B2(n6103), .ZN(
        P1_U3439) );
  AOI21_X1 U7772 ( .B1(n9793), .B2(n6105), .A(n6104), .ZN(n6106) );
  XNOR2_X1 U7773 ( .A(n6106), .B(P1_IR_REG_0__SCAN_IN), .ZN(n6110) );
  INV_X1 U7774 ( .A(n6107), .ZN(n6109) );
  AOI22_X1 U7775 ( .A1(n9261), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n6108) );
  OAI21_X1 U7776 ( .B1(n6110), .B2(n6109), .A(n6108), .ZN(P1_U3243) );
  INV_X1 U7777 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6112) );
  INV_X1 U7778 ( .A(n8496), .ZN(n8483) );
  OAI222_X1 U7779 ( .A1(n8991), .A2(n6112), .B1(n8990), .B2(n6111), .C1(
        P2_U3151), .C2(n8483), .ZN(P2_U3284) );
  INV_X1 U7780 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6113) );
  OAI222_X1 U7781 ( .A1(n8990), .A2(n7365), .B1(n9905), .B2(P2_U3151), .C1(
        n6113), .C2(n8991), .ZN(P2_U3283) );
  INV_X1 U7782 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10452) );
  NAND2_X1 U7783 ( .A1(n8763), .A2(P2_U3893), .ZN(n6114) );
  OAI21_X1 U7784 ( .B1(P2_U3893), .B2(n10452), .A(n6114), .ZN(P2_U3504) );
  NOR2_X1 U7785 ( .A1(n6116), .A2(n6115), .ZN(n6191) );
  OR2_X1 U7786 ( .A1(n6191), .A2(n5854), .ZN(n6117) );
  XNOR2_X1 U7787 ( .A(n6117), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7366) );
  INV_X1 U7788 ( .A(n7366), .ZN(n6647) );
  INV_X1 U7789 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10259) );
  OAI222_X1 U7790 ( .A1(P1_U3086), .A2(n6647), .B1(n7300), .B2(n7365), .C1(
        n10259), .C2(n6832), .ZN(P1_U3343) );
  NOR2_X1 U7791 ( .A1(n9261), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U7792 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7552) );
  INV_X1 U7793 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9604) );
  OR2_X1 U7794 ( .A1(n7992), .A2(n9604), .ZN(n6121) );
  INV_X1 U7795 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n6118) );
  OR2_X1 U7796 ( .A1(n7981), .A2(n6118), .ZN(n6120) );
  INV_X1 U7797 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9744) );
  OR2_X1 U7798 ( .A1(n4602), .A2(n9744), .ZN(n6119) );
  INV_X1 U7799 ( .A(n9311), .ZN(n8187) );
  NAND2_X1 U7800 ( .A1(n8187), .A2(P1_U3973), .ZN(n6122) );
  OAI21_X1 U7801 ( .B1(n7552), .B2(P1_U3973), .A(n6122), .ZN(P1_U3584) );
  INV_X1 U7802 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U7803 ( .A1(n4513), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6126) );
  INV_X1 U7804 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6123) );
  OR2_X1 U7805 ( .A1(n7981), .A2(n6123), .ZN(n6125) );
  INV_X1 U7806 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n7540) );
  OR2_X1 U7807 ( .A1(n4602), .A2(n7540), .ZN(n6124) );
  INV_X1 U7808 ( .A(n8252), .ZN(n8257) );
  NAND2_X1 U7809 ( .A1(n8257), .A2(P1_U3973), .ZN(n6127) );
  OAI21_X1 U7810 ( .B1(P1_U3973), .B2(n6128), .A(n6127), .ZN(P1_U3585) );
  NAND2_X1 U7811 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6569) );
  INV_X1 U7812 ( .A(n6569), .ZN(n6129) );
  NAND2_X1 U7813 ( .A1(n6129), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6741) );
  INV_X1 U7814 ( .A(n6741), .ZN(n6130) );
  NAND2_X1 U7815 ( .A1(n6130), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6864) );
  INV_X1 U7816 ( .A(n6864), .ZN(n6131) );
  NAND2_X1 U7817 ( .A1(n6131), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7040) );
  INV_X1 U7818 ( .A(n7054), .ZN(n6132) );
  NAND2_X1 U7819 ( .A1(n6132), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7241) );
  INV_X1 U7820 ( .A(n7266), .ZN(n6133) );
  NAND2_X1 U7821 ( .A1(n6133), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7346) );
  INV_X1 U7822 ( .A(n7834), .ZN(n6134) );
  NAND2_X1 U7823 ( .A1(n6134), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7847) );
  INV_X1 U7824 ( .A(n7847), .ZN(n6135) );
  NAND2_X1 U7825 ( .A1(n6135), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7864) );
  INV_X1 U7826 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7863) );
  AND2_X1 U7827 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n6136) );
  NAND2_X1 U7828 ( .A1(n9085), .A2(n6136), .ZN(n7906) );
  INV_X1 U7829 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7892) );
  INV_X1 U7830 ( .A(n7934), .ZN(n6138) );
  AND2_X1 U7831 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_21__SCAN_IN), 
        .ZN(n6137) );
  NAND2_X1 U7832 ( .A1(n6138), .A2(n6137), .ZN(n7945) );
  INV_X1 U7833 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9131) );
  INV_X1 U7834 ( .A(n7947), .ZN(n6139) );
  NAND2_X1 U7835 ( .A1(n6139), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7960) );
  INV_X1 U7836 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7837 ( .A1(n7947), .A2(n6140), .ZN(n6141) );
  NAND2_X1 U7838 ( .A1(n7960), .A2(n6141), .ZN(n9403) );
  NOR2_X1 U7839 ( .A1(n9403), .A2(n7988), .ZN(n6146) );
  INV_X1 U7840 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9404) );
  NOR2_X1 U7841 ( .A1(n7981), .A2(n9404), .ZN(n6145) );
  INV_X1 U7842 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n6143) );
  NAND2_X1 U7843 ( .A1(n7989), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6142) );
  OAI21_X1 U7844 ( .B1(n6143), .B2(n7992), .A(n6142), .ZN(n6144) );
  NAND2_X1 U7845 ( .A1(n9658), .A2(P1_U3973), .ZN(n6147) );
  OAI21_X1 U7846 ( .B1(P1_U3973), .B2(n7335), .A(n6147), .ZN(P1_U3577) );
  NAND2_X1 U7847 ( .A1(n7989), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6152) );
  INV_X1 U7848 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n6148) );
  OR2_X1 U7849 ( .A1(n7992), .A2(n6148), .ZN(n6151) );
  INV_X1 U7850 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9110) );
  XNOR2_X1 U7851 ( .A(n7934), .B(n9110), .ZN(n9449) );
  OR2_X1 U7852 ( .A1(n7988), .A2(n9449), .ZN(n6150) );
  INV_X1 U7853 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9450) );
  OR2_X1 U7854 ( .A1(n7981), .A2(n9450), .ZN(n6149) );
  NAND4_X1 U7855 ( .A1(n6152), .A2(n6151), .A3(n6150), .A4(n6149), .ZN(n9666)
         );
  NAND2_X1 U7856 ( .A1(n9666), .A2(P1_U3973), .ZN(n6153) );
  OAI21_X1 U7857 ( .B1(n5551), .B2(P1_U3973), .A(n6153), .ZN(P1_U3574) );
  INV_X4 U7858 ( .A(n6154), .ZN(n8561) );
  MUX2_X1 U7859 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8561), .Z(n6252) );
  XNOR2_X1 U7860 ( .A(n6252), .B(n6164), .ZN(n6163) );
  INV_X1 U7861 ( .A(n9880), .ZN(n6161) );
  MUX2_X1 U7862 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8561), .Z(n6159) );
  INV_X1 U7863 ( .A(n6159), .ZN(n6160) );
  MUX2_X1 U7864 ( .A(n8803), .B(n6155), .S(n5720), .Z(n6156) );
  XNOR2_X1 U7865 ( .A(n6156), .B(n9860), .ZN(n9857) );
  MUX2_X1 U7866 ( .A(n6170), .B(n5183), .S(n8561), .Z(n6227) );
  NAND2_X1 U7867 ( .A1(n6227), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n9856) );
  NAND2_X1 U7868 ( .A1(n9857), .A2(n9856), .ZN(n9855) );
  INV_X1 U7869 ( .A(n6156), .ZN(n6157) );
  NAND2_X1 U7870 ( .A1(n6157), .A2(n9860), .ZN(n6158) );
  NAND2_X1 U7871 ( .A1(n9855), .A2(n6158), .ZN(n9869) );
  XNOR2_X1 U7872 ( .A(n6159), .B(n6161), .ZN(n9868) );
  NOR2_X1 U7873 ( .A1(n6162), .A2(n6163), .ZN(n6253) );
  AOI21_X1 U7874 ( .B1(n6163), .B2(n6162), .A(n6253), .ZN(n6188) );
  NAND2_X1 U7875 ( .A1(P2_U3893), .A2(n5719), .ZN(n8566) );
  INV_X1 U7876 ( .A(n6164), .ZN(n6255) );
  NOR2_X1 U7877 ( .A1(n8561), .A2(P2_U3151), .ZN(n8987) );
  NAND2_X1 U7878 ( .A1(n6169), .A2(n8987), .ZN(n6165) );
  INV_X1 U7879 ( .A(n9977), .ZN(n8492) );
  INV_X1 U7880 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6185) );
  INV_X1 U7881 ( .A(n6166), .ZN(n7333) );
  NOR2_X1 U7882 ( .A1(n6167), .A2(n7333), .ZN(n6168) );
  NOR2_X1 U7883 ( .A1(n5719), .A2(P2_U3151), .ZN(n8983) );
  AND2_X1 U7884 ( .A1(n8983), .A2(n6169), .ZN(n6176) );
  INV_X1 U7885 ( .A(n6176), .ZN(n6226) );
  INV_X1 U7886 ( .A(n9963), .ZN(n8462) );
  NOR2_X1 U7887 ( .A1(n6170), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U7888 ( .A1(n6178), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6172) );
  INV_X1 U7889 ( .A(n6172), .ZN(n6173) );
  NOR2_X1 U7890 ( .A1(n9862), .A2(n6173), .ZN(n9883) );
  XNOR2_X1 U7891 ( .A(n9880), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n9884) );
  OAI21_X1 U7892 ( .B1(n6174), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6275), .ZN(
        n6175) );
  AOI22_X1 U7893 ( .A1(n8462), .A2(n6175), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        P2_U3151), .ZN(n6184) );
  XNOR2_X1 U7894 ( .A(n9880), .B(n10073), .ZN(n9873) );
  AND2_X1 U7895 ( .A1(n6177), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6179) );
  NAND2_X1 U7896 ( .A1(n6178), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6180) );
  OAI21_X1 U7897 ( .B1(n9860), .B2(n6179), .A(n6180), .ZN(n9851) );
  NAND2_X1 U7898 ( .A1(n9853), .A2(n6180), .ZN(n9872) );
  OAI21_X1 U7899 ( .B1(n6181), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6280), .ZN(
        n6182) );
  NAND2_X1 U7900 ( .A1(n9877), .A2(n6182), .ZN(n6183) );
  OAI211_X1 U7901 ( .C1(n6185), .C2(n9888), .A(n6184), .B(n6183), .ZN(n6186)
         );
  AOI21_X1 U7902 ( .B1(n6255), .B2(n8492), .A(n6186), .ZN(n6187) );
  OAI21_X1 U7903 ( .B1(n6188), .B2(n8566), .A(n6187), .ZN(P2_U3185) );
  INV_X1 U7904 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6189) );
  OAI222_X1 U7905 ( .A1(n8990), .A2(n7505), .B1(n9923), .B2(P2_U3151), .C1(
        n6189), .C2(n8991), .ZN(P2_U3282) );
  NAND2_X1 U7906 ( .A1(n6191), .A2(n6190), .ZN(n6266) );
  NAND2_X1 U7907 ( .A1(n6266), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6192) );
  XNOR2_X1 U7908 ( .A(n6192), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7506) );
  INV_X1 U7909 ( .A(n7506), .ZN(n6193) );
  OAI222_X1 U7910 ( .A1(n6193), .A2(P1_U3086), .B1(n6832), .B2(n10452), .C1(
        n7505), .C2(n7300), .ZN(P1_U3342) );
  INV_X1 U7911 ( .A(n7034), .ZN(n6202) );
  INV_X1 U7912 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7052) );
  MUX2_X1 U7913 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n7052), .S(n7230), .Z(n6195)
         );
  NAND2_X1 U7914 ( .A1(n6196), .A2(n6195), .ZN(n6322) );
  OAI21_X1 U7915 ( .B1(n6196), .B2(n6195), .A(n6322), .ZN(n6200) );
  INV_X1 U7916 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6198) );
  INV_X1 U7917 ( .A(n9258), .ZN(n9236) );
  NAND2_X1 U7918 ( .A1(n9236), .A2(n7230), .ZN(n6197) );
  NAND2_X1 U7919 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n7397) );
  OAI211_X1 U7920 ( .C1(n6198), .C2(n9234), .A(n6197), .B(n7397), .ZN(n6199)
         );
  AOI21_X1 U7921 ( .B1(n6200), .B2(n9255), .A(n6199), .ZN(n6209) );
  INV_X1 U7922 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6203) );
  MUX2_X1 U7923 ( .A(n6203), .B(P1_REG2_REG_9__SCAN_IN), .S(n7230), .Z(n6204)
         );
  INV_X1 U7924 ( .A(n6204), .ZN(n6205) );
  NAND2_X1 U7925 ( .A1(n6206), .A2(n6205), .ZN(n6326) );
  OAI21_X1 U7926 ( .B1(n6206), .B2(n6205), .A(n6326), .ZN(n6207) );
  INV_X1 U7927 ( .A(n9259), .ZN(n9230) );
  NAND2_X1 U7928 ( .A1(n6207), .A2(n9230), .ZN(n6208) );
  NAND2_X1 U7929 ( .A1(n6209), .A2(n6208), .ZN(P1_U3252) );
  NAND2_X1 U7930 ( .A1(n8838), .A2(P2_U3893), .ZN(n6210) );
  OAI21_X1 U7931 ( .B1(P2_U3893), .B2(n7494), .A(n6210), .ZN(P2_U3514) );
  NAND2_X1 U7932 ( .A1(n8796), .A2(n6211), .ZN(n7627) );
  AOI22_X1 U7933 ( .A1(n8406), .A2(n5870), .B1(n5191), .B2(n8419), .ZN(n6213)
         );
  NAND2_X1 U7934 ( .A1(n8428), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6319) );
  NAND2_X1 U7935 ( .A1(n6319), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6212) );
  OAI211_X1 U7936 ( .C1(n8421), .C2(n9978), .A(n6213), .B(n6212), .ZN(P2_U3172) );
  AOI211_X1 U7937 ( .C1(n6216), .C2(n6215), .A(n6214), .B(n9259), .ZN(n6225)
         );
  INV_X1 U7938 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U7939 ( .A1(n9236), .A2(n6217), .ZN(n6218) );
  NAND2_X1 U7940 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9017) );
  OAI211_X1 U7941 ( .C1(n6219), .C2(n9234), .A(n6218), .B(n9017), .ZN(n6224)
         );
  AOI211_X1 U7942 ( .C1(n6222), .C2(n6221), .A(n6220), .B(n9254), .ZN(n6223)
         );
  OR3_X1 U7943 ( .A1(n6225), .A2(n6224), .A3(n6223), .ZN(P1_U3246) );
  INV_X1 U7944 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U7945 ( .A1(n8492), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6231) );
  NAND2_X1 U7946 ( .A1(n6226), .A2(n8566), .ZN(n6229) );
  OAI21_X1 U7947 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6227), .A(n9856), .ZN(n6228) );
  AOI22_X1 U7948 ( .A1(n6229), .A2(n6228), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        P2_U3151), .ZN(n6230) );
  OAI211_X1 U7949 ( .C1(n9888), .C2(n6232), .A(n6231), .B(n6230), .ZN(P2_U3182) );
  INV_X1 U7950 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9101) );
  INV_X1 U7951 ( .A(n7976), .ZN(n6233) );
  NAND2_X1 U7952 ( .A1(n6233), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n7985) );
  INV_X1 U7953 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9146) );
  NAND2_X1 U7954 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6234) );
  INV_X1 U7955 ( .A(n9294), .ZN(n6239) );
  INV_X1 U7956 ( .A(n6551), .ZN(n7962) );
  INV_X1 U7957 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U7958 ( .A1(n7798), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7959 ( .A1(n7989), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6235) );
  OAI211_X1 U7960 ( .C1(n7992), .C2(n6237), .A(n6236), .B(n6235), .ZN(n6238)
         );
  AOI21_X1 U7961 ( .B1(n6239), .B2(n7962), .A(n6238), .ZN(n9319) );
  NAND2_X1 U7962 ( .A1(n9176), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6240) );
  OAI21_X1 U7963 ( .B1(n9319), .B2(n9176), .A(n6240), .ZN(P1_U3583) );
  INV_X1 U7964 ( .A(n6261), .ZN(n6337) );
  XNOR2_X1 U7965 ( .A(n6289), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n6274) );
  INV_X1 U7966 ( .A(n6342), .ZN(n6242) );
  AOI21_X1 U7967 ( .B1(n6260), .B2(n6243), .A(n6340), .ZN(n6250) );
  INV_X1 U7968 ( .A(n6244), .ZN(n6278) );
  XNOR2_X1 U7969 ( .A(n6289), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n6279) );
  AOI21_X1 U7970 ( .B1(n6280), .B2(n6278), .A(n6279), .ZN(n6282) );
  AOI21_X1 U7971 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n6289), .A(n6282), .ZN(
        n6245) );
  OAI21_X1 U7972 ( .B1(n6246), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6350), .ZN(
        n6247) );
  AOI22_X1 U7973 ( .A1(n6247), .A2(n9877), .B1(n9957), .B2(
        P2_ADDR_REG_5__SCAN_IN), .ZN(n6249) );
  INV_X1 U7974 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10404) );
  NOR2_X1 U7975 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10404), .ZN(n6309) );
  INV_X1 U7976 ( .A(n6309), .ZN(n6248) );
  OAI211_X1 U7977 ( .C1(n6250), .C2(n9963), .A(n6249), .B(n6248), .ZN(n6251)
         );
  AOI21_X1 U7978 ( .B1(n6337), .B2(n8492), .A(n6251), .ZN(n6265) );
  INV_X1 U7979 ( .A(n6289), .ZN(n6258) );
  MUX2_X1 U7980 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8561), .Z(n6256) );
  INV_X1 U7981 ( .A(n6256), .ZN(n6257) );
  INV_X1 U7982 ( .A(n6252), .ZN(n6254) );
  XOR2_X1 U7983 ( .A(n6289), .B(n6256), .Z(n6272) );
  NAND2_X1 U7984 ( .A1(n6273), .A2(n6272), .ZN(n6271) );
  OAI21_X1 U7985 ( .B1(n6258), .B2(n6257), .A(n6271), .ZN(n6263) );
  MUX2_X1 U7986 ( .A(n6260), .B(n6259), .S(n8561), .Z(n6336) );
  XNOR2_X1 U7987 ( .A(n6336), .B(n6261), .ZN(n6262) );
  NAND2_X1 U7988 ( .A1(n6263), .A2(n6262), .ZN(n6335) );
  OAI211_X1 U7989 ( .C1(n6263), .C2(n6262), .A(n6335), .B(n9967), .ZN(n6264)
         );
  NAND2_X1 U7990 ( .A1(n6265), .A2(n6264), .ZN(P2_U3187) );
  NAND2_X1 U7991 ( .A1(n6267), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6373) );
  XNOR2_X1 U7992 ( .A(n6373), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9187) );
  INV_X1 U7993 ( .A(n9187), .ZN(n6268) );
  INV_X1 U7994 ( .A(n7509), .ZN(n6269) );
  INV_X1 U7995 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10234) );
  OAI222_X1 U7996 ( .A1(n6268), .A2(P1_U3086), .B1(n7300), .B2(n6269), .C1(
        n10234), .C2(n6832), .ZN(P1_U3341) );
  INV_X1 U7997 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6270) );
  OAI222_X1 U7998 ( .A1(n8991), .A2(n6270), .B1(n8990), .B2(n6269), .C1(
        P2_U3151), .C2(n9940), .ZN(P2_U3281) );
  OAI211_X1 U7999 ( .C1(n6273), .C2(n6272), .A(n6271), .B(n9967), .ZN(n6288)
         );
  AND3_X1 U8000 ( .A1(n6275), .A2(n6274), .A3(n4530), .ZN(n6276) );
  OAI21_X1 U8001 ( .B1(n6277), .B2(n6276), .A(n8462), .ZN(n6285) );
  AND3_X1 U8002 ( .A1(n6280), .A2(n6279), .A3(n6278), .ZN(n6281) );
  OAI21_X1 U8003 ( .B1(n6282), .B2(n6281), .A(n9877), .ZN(n6283) );
  NAND3_X1 U8004 ( .A1(n6285), .A2(n6284), .A3(n6283), .ZN(n6286) );
  AOI21_X1 U8005 ( .B1(n9957), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6286), .ZN(
        n6287) );
  OAI211_X1 U8006 ( .C1(n9977), .C2(n6289), .A(n6288), .B(n6287), .ZN(P2_U3186) );
  INV_X1 U8007 ( .A(n6290), .ZN(n6291) );
  AOI211_X1 U8008 ( .C1(n6293), .C2(n6292), .A(n8421), .B(n6291), .ZN(n6298)
         );
  INV_X1 U8009 ( .A(n8419), .ZN(n8434) );
  INV_X1 U8010 ( .A(n10001), .ZN(n8442) );
  AOI22_X1 U8011 ( .A1(n8431), .A2(n9998), .B1(n8406), .B2(n8442), .ZN(n6295)
         );
  MUX2_X1 U8012 ( .A(n8428), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n6294) );
  OAI211_X1 U8013 ( .C1(n6296), .C2(n8434), .A(n6295), .B(n6294), .ZN(n6297)
         );
  OR2_X1 U8014 ( .A1(n6298), .A2(n6297), .ZN(P2_U3158) );
  INV_X1 U8015 ( .A(n7512), .ZN(n6376) );
  AOI22_X1 U8016 ( .A1(n8536), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n8988), .ZN(n6299) );
  OAI21_X1 U8017 ( .B1(n6376), .B2(n8990), .A(n6299), .ZN(P2_U3280) );
  XOR2_X1 U8018 ( .A(n6301), .B(n6300), .Z(n6305) );
  AOI22_X1 U8019 ( .A1(n8406), .A2(n9998), .B1(n8431), .B2(n8796), .ZN(n6302)
         );
  OAI21_X1 U8020 ( .B1(n8790), .B2(n8434), .A(n6302), .ZN(n6303) );
  AOI21_X1 U8021 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n6319), .A(n6303), .ZN(
        n6304) );
  OAI21_X1 U8022 ( .B1(n8421), .B2(n6305), .A(n6304), .ZN(P2_U3162) );
  NAND2_X1 U8023 ( .A1(n6306), .A2(n10001), .ZN(n6307) );
  XNOR2_X1 U8024 ( .A(n8051), .B(n6427), .ZN(n6363) );
  XNOR2_X1 U8025 ( .A(n6363), .B(n8441), .ZN(n6364) );
  XNOR2_X1 U8026 ( .A(n6365), .B(n6364), .ZN(n6313) );
  AOI22_X1 U8027 ( .A1(n8406), .A2(n8440), .B1(n6427), .B2(n8419), .ZN(n6311)
         );
  AOI21_X1 U8028 ( .B1(n8431), .B2(n8442), .A(n6309), .ZN(n6310) );
  OAI211_X1 U8029 ( .C1(n6424), .C2(n8428), .A(n6311), .B(n6310), .ZN(n6312)
         );
  AOI21_X1 U8030 ( .B1(n6313), .B2(n8423), .A(n6312), .ZN(n6314) );
  INV_X1 U8031 ( .A(n6314), .ZN(P2_U3167) );
  XOR2_X1 U8032 ( .A(n6316), .B(n6315), .Z(n6321) );
  AOI22_X1 U8033 ( .A1(n8431), .A2(n5870), .B1(n8406), .B2(n10008), .ZN(n6317)
         );
  OAI21_X1 U8034 ( .B1(n9989), .B2(n8434), .A(n6317), .ZN(n6318) );
  AOI21_X1 U8035 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n6319), .A(n6318), .ZN(
        n6320) );
  OAI21_X1 U8036 ( .B1(n8421), .B2(n6321), .A(n6320), .ZN(P2_U3177) );
  OAI21_X1 U8037 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n7230), .A(n6322), .ZN(
        n6325) );
  NAND2_X1 U8038 ( .A1(n7253), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6323) );
  OAI21_X1 U8039 ( .B1(n7253), .B2(P1_REG1_REG_10__SCAN_IN), .A(n6323), .ZN(
        n6324) );
  NOR2_X1 U8040 ( .A1(n6324), .A2(n6325), .ZN(n6525) );
  AOI211_X1 U8041 ( .C1(n6325), .C2(n6324), .A(n6525), .B(n9254), .ZN(n6334)
         );
  OAI21_X1 U8042 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n7230), .A(n6326), .ZN(
        n6329) );
  NAND2_X1 U8043 ( .A1(n7253), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6327) );
  OAI21_X1 U8044 ( .B1(n7253), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6327), .ZN(
        n6328) );
  NOR2_X1 U8045 ( .A1(n6328), .A2(n6329), .ZN(n6521) );
  AOI211_X1 U8046 ( .C1(n6329), .C2(n6328), .A(n6521), .B(n9259), .ZN(n6333)
         );
  INV_X1 U8047 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U8048 ( .A1(n9236), .A2(n7253), .ZN(n6330) );
  NAND2_X1 U8049 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n7427) );
  OAI211_X1 U8050 ( .C1(n6331), .C2(n9234), .A(n6330), .B(n7427), .ZN(n6332)
         );
  OR3_X1 U8051 ( .A1(n6334), .A2(n6333), .A3(n6332), .ZN(P1_U3253) );
  MUX2_X1 U8052 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8561), .Z(n6501) );
  XNOR2_X1 U8053 ( .A(n6501), .B(n6505), .ZN(n6339) );
  OAI21_X1 U8054 ( .B1(n6337), .B2(n6336), .A(n6335), .ZN(n6338) );
  NOR2_X1 U8055 ( .A1(n6338), .A2(n6339), .ZN(n6502) );
  AOI21_X1 U8056 ( .B1(n6339), .B2(n6338), .A(n6502), .ZN(n6356) );
  INV_X1 U8057 ( .A(n6505), .ZN(n6509) );
  INV_X1 U8058 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6347) );
  MUX2_X1 U8059 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6508), .S(n6505), .Z(n6341)
         );
  NOR3_X1 U8060 ( .A1(n6342), .A2(n6341), .A3(n6340), .ZN(n6343) );
  OAI21_X1 U8061 ( .B1(n4601), .B2(n6343), .A(n8462), .ZN(n6346) );
  INV_X1 U8062 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6344) );
  NOR2_X1 U8063 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6344), .ZN(n6369) );
  INV_X1 U8064 ( .A(n6369), .ZN(n6345) );
  OAI211_X1 U8065 ( .C1(n9888), .C2(n6347), .A(n6346), .B(n6345), .ZN(n6354)
         );
  INV_X1 U8066 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6348) );
  MUX2_X1 U8067 ( .A(n6348), .B(P2_REG1_REG_6__SCAN_IN), .S(n6505), .Z(n6349)
         );
  INV_X1 U8068 ( .A(n6504), .ZN(n6352) );
  NAND3_X1 U8069 ( .A1(n6350), .A2(n6349), .A3(n4529), .ZN(n6351) );
  AOI21_X1 U8070 ( .B1(n6352), .B2(n6351), .A(n9971), .ZN(n6353) );
  AOI211_X1 U8071 ( .C1(n8492), .C2(n6509), .A(n6354), .B(n6353), .ZN(n6355)
         );
  OAI21_X1 U8072 ( .B1(n6356), .B2(n8566), .A(n6355), .ZN(P2_U3188) );
  INV_X1 U8073 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8012) );
  INV_X1 U8074 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6357) );
  OAI21_X1 U8075 ( .B1(n7987), .B2(n8012), .A(n6357), .ZN(n6358) );
  INV_X1 U8076 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9618) );
  NAND2_X1 U8077 ( .A1(n7989), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6360) );
  NAND2_X1 U8078 ( .A1(n7798), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6359) );
  OAI211_X1 U8079 ( .C1(n7992), .C2(n9618), .A(n6360), .B(n6359), .ZN(n6361)
         );
  NAND2_X1 U8080 ( .A1(n9176), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6362) );
  OAI21_X1 U8081 ( .B1(n9607), .B2(n9176), .A(n6362), .ZN(P1_U3582) );
  XNOR2_X1 U8082 ( .A(n10021), .B(n8051), .ZN(n6582) );
  XNOR2_X1 U8083 ( .A(n6582), .B(n8440), .ZN(n6366) );
  OAI211_X1 U8084 ( .C1(n6367), .C2(n6366), .A(n6585), .B(n8423), .ZN(n6371)
         );
  OAI22_X1 U8085 ( .A1(n8434), .A2(n6766), .B1(n8427), .B2(n6785), .ZN(n6368)
         );
  AOI211_X1 U8086 ( .C1(n8431), .C2(n8441), .A(n6369), .B(n6368), .ZN(n6370)
         );
  OAI211_X1 U8087 ( .C1(n6765), .C2(n8428), .A(n6371), .B(n6370), .ZN(P2_U3179) );
  NAND2_X1 U8088 ( .A1(n6373), .A2(n6372), .ZN(n6374) );
  NAND2_X1 U8089 ( .A1(n6374), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6378) );
  XNOR2_X1 U8090 ( .A(n6378), .B(n10283), .ZN(n9201) );
  INV_X1 U8091 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6375) );
  OAI222_X1 U8092 ( .A1(n9201), .A2(P1_U3086), .B1(n7300), .B2(n6376), .C1(
        n6375), .C2(n6832), .ZN(P1_U3340) );
  INV_X1 U8093 ( .A(n7515), .ZN(n6382) );
  INV_X1 U8094 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6377) );
  OAI222_X1 U8095 ( .A1(n8990), .A2(n6382), .B1(n9956), .B2(P2_U3151), .C1(
        n6377), .C2(n8991), .ZN(P2_U3279) );
  INV_X1 U8096 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10420) );
  NAND2_X1 U8097 ( .A1(n6378), .A2(n10283), .ZN(n6379) );
  NAND2_X1 U8098 ( .A1(n6379), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6380) );
  XNOR2_X1 U8099 ( .A(n6380), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9217) );
  INV_X1 U8100 ( .A(n9217), .ZN(n6381) );
  OAI222_X1 U8101 ( .A1(n6832), .A2(n10420), .B1(n7300), .B2(n6382), .C1(
        P1_U3086), .C2(n6381), .ZN(P1_U3339) );
  OR2_X1 U8102 ( .A1(n6470), .A2(n6469), .ZN(n6904) );
  INV_X1 U8103 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6383) );
  NAND2_X1 U8104 ( .A1(n6395), .A2(n6383), .ZN(n6384) );
  NAND2_X1 U8105 ( .A1(n7558), .A2(n9794), .ZN(n9785) );
  NAND2_X1 U8106 ( .A1(n6384), .A2(n9785), .ZN(n6466) );
  NOR4_X1 U8107 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6393) );
  NOR4_X1 U8108 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6392) );
  INV_X1 U8109 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n9798) );
  INV_X1 U8110 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10429) );
  INV_X1 U8111 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10487) );
  INV_X1 U8112 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10368) );
  NAND4_X1 U8113 ( .A1(n9798), .A2(n10429), .A3(n10487), .A4(n10368), .ZN(
        n6390) );
  NOR4_X1 U8114 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6388) );
  NOR4_X1 U8115 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6387) );
  NOR4_X1 U8116 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6386) );
  NOR4_X1 U8117 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6385) );
  NAND4_X1 U8118 ( .A1(n6388), .A2(n6387), .A3(n6386), .A4(n6385), .ZN(n6389)
         );
  NOR4_X1 U8119 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6390), .A4(n6389), .ZN(n6391) );
  NAND3_X1 U8120 ( .A1(n6393), .A2(n6392), .A3(n6391), .ZN(n6394) );
  NAND2_X1 U8121 ( .A1(n6395), .A2(n6394), .ZN(n6905) );
  NAND2_X1 U8122 ( .A1(n6395), .A2(n10433), .ZN(n6397) );
  INV_X1 U8123 ( .A(n6467), .ZN(n6908) );
  AND2_X1 U8124 ( .A1(n6917), .A2(n9178), .ZN(n8073) );
  AND2_X1 U8125 ( .A1(n5954), .A2(n9343), .ZN(n6399) );
  OR2_X1 U8126 ( .A1(n6470), .A2(n6398), .ZN(n6485) );
  NAND2_X1 U8127 ( .A1(n5954), .A2(n9327), .ZN(n6400) );
  NOR2_X1 U8128 ( .A1(n9834), .A2(n9713), .ZN(n6406) );
  INV_X1 U8129 ( .A(n6470), .ZN(n8259) );
  NAND2_X1 U8130 ( .A1(n4513), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6405) );
  INV_X1 U8131 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7204) );
  OR2_X1 U8132 ( .A1(n6551), .A2(n7204), .ZN(n6404) );
  OR2_X1 U8133 ( .A1(n7981), .A2(n4739), .ZN(n6403) );
  INV_X1 U8134 ( .A(n7933), .ZN(n6401) );
  INV_X1 U8135 ( .A(n9177), .ZN(n6704) );
  OAI222_X1 U8136 ( .A1(n6917), .A2(n6912), .B1(n4528), .B2(n6406), .C1(n9731), 
        .C2(n6704), .ZN(n6410) );
  NAND2_X1 U8137 ( .A1(n6410), .A2(n9838), .ZN(n6407) );
  OAI21_X1 U8138 ( .B1(n9838), .B2(n5931), .A(n6407), .ZN(P1_U3453) );
  NAND2_X1 U8139 ( .A1(n6410), .A2(n9850), .ZN(n6411) );
  OAI21_X1 U8140 ( .B1(n9850), .B2(n6105), .A(n6411), .ZN(P1_U3522) );
  OR2_X1 U8141 ( .A1(n6412), .A2(n7618), .ZN(n6763) );
  INV_X1 U8142 ( .A(n6763), .ZN(n6987) );
  XNOR2_X1 U8143 ( .A(n10011), .B(n6427), .ZN(n7595) );
  XNOR2_X1 U8144 ( .A(n6413), .B(n7595), .ZN(n10015) );
  INV_X1 U8145 ( .A(n10015), .ZN(n6418) );
  XNOR2_X1 U8146 ( .A(n6414), .B(n7595), .ZN(n6416) );
  OAI22_X1 U8147 ( .A1(n10028), .A2(n10025), .B1(n10001), .B2(n10027), .ZN(
        n6415) );
  AOI21_X1 U8148 ( .B1(n6416), .B2(n10005), .A(n6415), .ZN(n6417) );
  OAI21_X1 U8149 ( .B1(n10015), .B2(n9988), .A(n6417), .ZN(n10017) );
  AOI21_X1 U8150 ( .B1(n6987), .B2(n6418), .A(n10017), .ZN(n6429) );
  NAND2_X1 U8151 ( .A1(n6420), .A2(n6419), .ZN(n6421) );
  NOR2_X1 U8152 ( .A1(n8788), .A2(n6424), .ZN(n6426) );
  NOR2_X1 U8153 ( .A1(n8728), .A2(n6260), .ZN(n6425) );
  AOI211_X1 U8154 ( .C1(n8745), .C2(n6427), .A(n6426), .B(n6425), .ZN(n6428)
         );
  OAI21_X1 U8155 ( .B1(n6429), .B2(n8802), .A(n6428), .ZN(P2_U3228) );
  OR2_X1 U8156 ( .A1(n6430), .A2(n7998), .ZN(n6431) );
  NAND2_X1 U8157 ( .A1(n6432), .A2(n6431), .ZN(n6616) );
  NAND2_X1 U8158 ( .A1(n9177), .A2(n6541), .ZN(n6436) );
  NAND2_X1 U8159 ( .A1(n7206), .A2(n4892), .ZN(n6435) );
  NAND2_X1 U8160 ( .A1(n6436), .A2(n6435), .ZN(n6437) );
  XNOR2_X1 U8161 ( .A(n6437), .B(n8292), .ZN(n6441) );
  NAND2_X1 U8162 ( .A1(n9177), .A2(n7959), .ZN(n6439) );
  NAND2_X1 U8163 ( .A1(n7206), .A2(n6541), .ZN(n6438) );
  AND2_X1 U8164 ( .A1(n6439), .A2(n6438), .ZN(n6615) );
  NAND2_X1 U8165 ( .A1(n6441), .A2(n6615), .ZN(n6440) );
  INV_X1 U8166 ( .A(n6441), .ZN(n6617) );
  INV_X1 U8167 ( .A(n6615), .ZN(n6442) );
  OR2_X1 U8168 ( .A1(n6546), .A2(n5196), .ZN(n6447) );
  OR2_X1 U8169 ( .A1(n7229), .A2(n6444), .ZN(n6445) );
  NAND2_X1 U8170 ( .A1(n4513), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6453) );
  INV_X1 U8171 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6484) );
  OR2_X1 U8172 ( .A1(n6551), .A2(n6484), .ZN(n6452) );
  INV_X1 U8173 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6448) );
  OR2_X1 U8174 ( .A1(n7981), .A2(n6448), .ZN(n6451) );
  INV_X1 U8175 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6449) );
  OR2_X1 U8176 ( .A1(n7933), .A2(n6449), .ZN(n6450) );
  NAND2_X1 U8177 ( .A1(n6676), .A2(n6541), .ZN(n6454) );
  OAI21_X1 U8178 ( .B1(n8077), .B2(n7883), .A(n6454), .ZN(n6455) );
  XNOR2_X1 U8179 ( .A(n6455), .B(n8292), .ZN(n6458) );
  OR2_X1 U8180 ( .A1(n8077), .A2(n7307), .ZN(n6457) );
  NAND2_X1 U8181 ( .A1(n9175), .A2(n7959), .ZN(n6456) );
  AND2_X1 U8182 ( .A1(n6457), .A2(n6456), .ZN(n6459) );
  NAND2_X1 U8183 ( .A1(n6458), .A2(n6459), .ZN(n6531) );
  INV_X1 U8184 ( .A(n6458), .ZN(n6461) );
  INV_X1 U8185 ( .A(n6459), .ZN(n6460) );
  NAND2_X1 U8186 ( .A1(n6461), .A2(n6460), .ZN(n6462) );
  NAND2_X1 U8187 ( .A1(n6531), .A2(n6462), .ZN(n6465) );
  INV_X1 U8188 ( .A(n6465), .ZN(n6463) );
  NAND2_X1 U8189 ( .A1(n6465), .A2(n6464), .ZN(n6472) );
  INV_X1 U8190 ( .A(n6466), .ZN(n6907) );
  NAND3_X1 U8191 ( .A1(n6907), .A2(n6467), .A3(n6905), .ZN(n6479) );
  INV_X1 U8192 ( .A(n8271), .ZN(n6468) );
  AND2_X1 U8193 ( .A1(n9831), .A2(n6470), .ZN(n6471) );
  AOI21_X1 U8194 ( .B1(n6532), .B2(n6472), .A(n9164), .ZN(n6495) );
  INV_X1 U8195 ( .A(n6486), .ZN(n6476) );
  NOR2_X1 U8196 ( .A1(n6912), .A2(n6477), .ZN(n6910) );
  INV_X1 U8197 ( .A(n6910), .ZN(n6475) );
  NOR2_X1 U8198 ( .A1(n6477), .A2(P1_U3086), .ZN(n6930) );
  OR2_X1 U8199 ( .A1(n9831), .A2(n6930), .ZN(n6478) );
  NAND2_X1 U8200 ( .A1(n6479), .A2(n6478), .ZN(n6483) );
  INV_X1 U8201 ( .A(n6480), .ZN(n6481) );
  AND3_X1 U8202 ( .A1(n5958), .A2(n6481), .A3(n6904), .ZN(n6482) );
  NAND2_X1 U8203 ( .A1(n6483), .A2(n6482), .ZN(n9088) );
  NOR2_X1 U8204 ( .A1(n9088), .A2(P1_U3086), .ZN(n6619) );
  OAI22_X1 U8205 ( .A1(n9126), .A2(n8077), .B1(n6619), .B2(n6484), .ZN(n6494)
         );
  INV_X1 U8206 ( .A(n6485), .ZN(n8270) );
  NAND2_X1 U8207 ( .A1(n6486), .A2(n8270), .ZN(n6487) );
  INV_X1 U8208 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7122) );
  OR2_X1 U8209 ( .A1(n7981), .A2(n7122), .ZN(n6492) );
  OR2_X1 U8210 ( .A1(n6551), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6491) );
  NAND2_X1 U8211 ( .A1(n7978), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6490) );
  INV_X1 U8212 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6488) );
  OR2_X1 U8213 ( .A1(n7933), .A2(n6488), .ZN(n6489) );
  INV_X1 U8214 ( .A(n9174), .ZN(n8076) );
  OAI22_X1 U8215 ( .A1(n6704), .A2(n9159), .B1(n9158), .B2(n8076), .ZN(n6493)
         );
  OR3_X1 U8216 ( .A1(n6495), .A2(n6494), .A3(n6493), .ZN(P1_U3237) );
  INV_X1 U8217 ( .A(n9158), .ZN(n9072) );
  OAI22_X1 U8218 ( .A1(n9126), .A2(n6917), .B1(n6619), .B2(n6911), .ZN(n6496)
         );
  AOI21_X1 U8219 ( .B1(n9072), .B2(n9177), .A(n6496), .ZN(n6497) );
  OAI21_X1 U8220 ( .B1(n9164), .B2(n6498), .A(n6497), .ZN(P1_U3232) );
  MUX2_X1 U8221 ( .A(n6500), .B(n6499), .S(n8561), .Z(n6815) );
  XNOR2_X1 U8222 ( .A(n6815), .B(n6506), .ZN(n6818) );
  INV_X1 U8223 ( .A(n6501), .ZN(n6503) );
  XOR2_X1 U8224 ( .A(n6818), .B(n6819), .Z(n6518) );
  OAI21_X1 U8225 ( .B1(n6507), .B2(P2_REG1_REG_7__SCAN_IN), .A(n8452), .ZN(
        n6516) );
  OAI21_X1 U8226 ( .B1(n6510), .B2(n6816), .A(n8458), .ZN(n6511) );
  AOI21_X1 U8227 ( .B1(n6500), .B2(n6511), .A(n8461), .ZN(n6514) );
  NOR2_X1 U8228 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5314), .ZN(n6592) );
  NOR2_X1 U8229 ( .A1(n9977), .A2(n6816), .ZN(n6512) );
  AOI211_X1 U8230 ( .C1(n9957), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n6592), .B(
        n6512), .ZN(n6513) );
  OAI21_X1 U8231 ( .B1(n6514), .B2(n9963), .A(n6513), .ZN(n6515) );
  AOI21_X1 U8232 ( .B1(n6516), .B2(n9877), .A(n6515), .ZN(n6517) );
  OAI21_X1 U8233 ( .B1(n6518), .B2(n8566), .A(n6517), .ZN(P2_U3189) );
  INV_X1 U8234 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6520) );
  NAND2_X1 U8235 ( .A1(n9236), .A2(n7340), .ZN(n6519) );
  NAND2_X1 U8236 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n7444) );
  OAI211_X1 U8237 ( .C1(n6520), .C2(n9234), .A(n6519), .B(n7444), .ZN(n6530)
         );
  NAND2_X1 U8238 ( .A1(n7340), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6522) );
  OAI21_X1 U8239 ( .B1(n7340), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6522), .ZN(
        n6523) );
  AOI211_X1 U8240 ( .C1(n6524), .C2(n6523), .A(n6641), .B(n9259), .ZN(n6529)
         );
  INV_X1 U8241 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7264) );
  MUX2_X1 U8242 ( .A(n7264), .B(P1_REG1_REG_11__SCAN_IN), .S(n7340), .Z(n6526)
         );
  AOI211_X1 U8243 ( .C1(n6527), .C2(n6526), .A(n6637), .B(n9254), .ZN(n6528)
         );
  OR3_X1 U8244 ( .A1(n6530), .A2(n6529), .A3(n6528), .ZN(P1_U3254) );
  OR2_X1 U8245 ( .A1(n6546), .A2(n6533), .ZN(n6538) );
  OR2_X1 U8246 ( .A1(n6544), .A2(n6534), .ZN(n6537) );
  OR2_X1 U8247 ( .A1(n7229), .A2(n6535), .ZN(n6536) );
  AND3_X2 U8248 ( .A1(n6538), .A2(n6537), .A3(n6536), .ZN(n6722) );
  NAND2_X1 U8249 ( .A1(n9174), .A2(n6541), .ZN(n6539) );
  OAI21_X1 U8250 ( .B1(n6722), .B2(n7883), .A(n6539), .ZN(n6540) );
  XNOR2_X1 U8251 ( .A(n6540), .B(n8292), .ZN(n6563) );
  OR2_X1 U8252 ( .A1(n6722), .A2(n7307), .ZN(n6543) );
  NAND2_X1 U8253 ( .A1(n9174), .A2(n7959), .ZN(n6542) );
  NAND2_X1 U8254 ( .A1(n6543), .A2(n6542), .ZN(n6561) );
  XNOR2_X1 U8255 ( .A(n6563), .B(n6561), .ZN(n9014) );
  NAND2_X1 U8256 ( .A1(n9013), .A2(n9014), .ZN(n6565) );
  OR2_X1 U8257 ( .A1(n7504), .A2(n6545), .ZN(n6550) );
  OR2_X1 U8258 ( .A1(n7534), .A2(n4707), .ZN(n6549) );
  OR2_X1 U8259 ( .A1(n4512), .A2(n6547), .ZN(n6548) );
  NAND2_X1 U8260 ( .A1(n4513), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6556) );
  OR2_X1 U8261 ( .A1(n7981), .A2(n7016), .ZN(n6555) );
  OAI21_X1 U8262 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n6569), .ZN(n7015) );
  OR2_X1 U8263 ( .A1(n7988), .A2(n7015), .ZN(n6554) );
  INV_X1 U8264 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6552) );
  OR2_X1 U8265 ( .A1(n7933), .A2(n6552), .ZN(n6553) );
  NAND2_X1 U8266 ( .A1(n9173), .A2(n6541), .ZN(n6557) );
  OAI21_X1 U8267 ( .B1(n9801), .B2(n7883), .A(n6557), .ZN(n6558) );
  XNOR2_X1 U8268 ( .A(n6558), .B(n8292), .ZN(n6834) );
  OR2_X1 U8269 ( .A1(n9801), .A2(n7307), .ZN(n6560) );
  NAND2_X1 U8270 ( .A1(n9173), .A2(n7959), .ZN(n6559) );
  NAND2_X1 U8271 ( .A1(n6560), .A2(n6559), .ZN(n6835) );
  XNOR2_X1 U8272 ( .A(n6834), .B(n6835), .ZN(n6566) );
  INV_X1 U8273 ( .A(n6561), .ZN(n6562) );
  NAND2_X1 U8274 ( .A1(n6563), .A2(n6562), .ZN(n6567) );
  AND2_X1 U8275 ( .A1(n6566), .A2(n6567), .ZN(n6564) );
  NAND2_X1 U8276 ( .A1(n6565), .A2(n6564), .ZN(n6838) );
  NAND2_X1 U8277 ( .A1(n6838), .A2(n9143), .ZN(n6581) );
  AOI21_X1 U8278 ( .B1(n6565), .B2(n6567), .A(n6566), .ZN(n6580) );
  NAND2_X1 U8279 ( .A1(n4513), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6575) );
  OR2_X1 U8280 ( .A1(n7981), .A2(n7217), .ZN(n6574) );
  INV_X1 U8281 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6568) );
  NAND2_X1 U8282 ( .A1(n6569), .A2(n6568), .ZN(n6570) );
  NAND2_X1 U8283 ( .A1(n6741), .A2(n6570), .ZN(n9074) );
  OR2_X1 U8284 ( .A1(n7988), .A2(n9074), .ZN(n6573) );
  INV_X1 U8285 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6571) );
  OR2_X1 U8286 ( .A1(n7933), .A2(n6571), .ZN(n6572) );
  INV_X1 U8287 ( .A(n9801), .ZN(n7018) );
  AOI22_X1 U8288 ( .A1(n9072), .A2(n9172), .B1(n7018), .B2(n9162), .ZN(n6579)
         );
  INV_X1 U8289 ( .A(n9159), .ZN(n9077) );
  NOR2_X1 U8290 ( .A1(n9157), .A2(n7015), .ZN(n6576) );
  AOI211_X1 U8291 ( .C1(n9077), .C2(n9174), .A(n6577), .B(n6576), .ZN(n6578)
         );
  OAI211_X1 U8292 ( .C1(n6581), .C2(n6580), .A(n6579), .B(n6578), .ZN(P1_U3230) );
  XNOR2_X1 U8293 ( .A(n10030), .B(n8048), .ZN(n6602) );
  XNOR2_X1 U8294 ( .A(n6602), .B(n8439), .ZN(n6589) );
  INV_X1 U8295 ( .A(n6582), .ZN(n6583) );
  NAND2_X1 U8296 ( .A1(n6583), .A2(n8440), .ZN(n6584) );
  INV_X1 U8297 ( .A(n6589), .ZN(n6586) );
  INV_X1 U8298 ( .A(n6605), .ZN(n6587) );
  AOI21_X1 U8299 ( .B1(n6589), .B2(n6588), .A(n6587), .ZN(n6596) );
  INV_X1 U8300 ( .A(n10030), .ZN(n6590) );
  OAI22_X1 U8301 ( .A1(n8434), .A2(n6590), .B1(n8427), .B2(n10026), .ZN(n6591)
         );
  AOI211_X1 U8302 ( .C1(n8431), .C2(n8440), .A(n6592), .B(n6591), .ZN(n6595)
         );
  INV_X1 U8303 ( .A(n6995), .ZN(n6593) );
  NAND2_X1 U8304 ( .A1(n8415), .A2(n6593), .ZN(n6594) );
  OAI211_X1 U8305 ( .C1(n6596), .C2(n8421), .A(n6595), .B(n6594), .ZN(P2_U3153) );
  NAND2_X1 U8306 ( .A1(n6597), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6598) );
  XNOR2_X1 U8307 ( .A(n6598), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9215) );
  INV_X1 U8308 ( .A(n9215), .ZN(n9238) );
  INV_X1 U8309 ( .A(n7518), .ZN(n6600) );
  OAI222_X1 U8310 ( .A1(n9238), .A2(P1_U3086), .B1(n7300), .B2(n6600), .C1(
        n6599), .C2(n6832), .ZN(P1_U3338) );
  OAI222_X1 U8311 ( .A1(n8991), .A2(n6601), .B1(n8990), .B2(n6600), .C1(
        P2_U3151), .C2(n9976), .ZN(P2_U3278) );
  INV_X1 U8312 ( .A(n6602), .ZN(n6603) );
  NAND2_X1 U8313 ( .A1(n6603), .A2(n6785), .ZN(n6604) );
  XNOR2_X1 U8314 ( .A(n6789), .B(n5869), .ZN(n6606) );
  AND2_X1 U8315 ( .A1(n6606), .A2(n10026), .ZN(n6652) );
  INV_X1 U8316 ( .A(n6652), .ZN(n6608) );
  INV_X1 U8317 ( .A(n6606), .ZN(n6607) );
  NAND2_X1 U8318 ( .A1(n6607), .A2(n10044), .ZN(n6651) );
  NAND2_X1 U8319 ( .A1(n6608), .A2(n6651), .ZN(n6609) );
  XNOR2_X1 U8320 ( .A(n6653), .B(n6609), .ZN(n6614) );
  OR2_X1 U8321 ( .A1(n8427), .A2(n6947), .ZN(n6610) );
  INV_X1 U8322 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10221) );
  OR2_X1 U8323 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10221), .ZN(n8447) );
  OAI211_X1 U8324 ( .C1(n8409), .C2(n6785), .A(n6610), .B(n8447), .ZN(n6612)
         );
  NOR2_X1 U8325 ( .A1(n8428), .A2(n6786), .ZN(n6611) );
  AOI211_X1 U8326 ( .C1(n6789), .C2(n8419), .A(n6612), .B(n6611), .ZN(n6613)
         );
  OAI21_X1 U8327 ( .B1(n6614), .B2(n8421), .A(n6613), .ZN(P2_U3161) );
  XNOR2_X1 U8328 ( .A(n6616), .B(n6615), .ZN(n6618) );
  XNOR2_X1 U8329 ( .A(n6618), .B(n6617), .ZN(n6623) );
  INV_X1 U8330 ( .A(n9175), .ZN(n6677) );
  NOR2_X1 U8331 ( .A1(n9158), .A2(n6677), .ZN(n6621) );
  INV_X1 U8332 ( .A(n7206), .ZN(n8078) );
  OAI22_X1 U8333 ( .A1(n9126), .A2(n8078), .B1(n6619), .B2(n7204), .ZN(n6620)
         );
  AOI211_X1 U8334 ( .C1(n9077), .C2(n9178), .A(n6621), .B(n6620), .ZN(n6622)
         );
  OAI21_X1 U8335 ( .B1(n6623), .B2(n9164), .A(n6622), .ZN(P1_U3222) );
  INV_X1 U8336 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10446) );
  INV_X1 U8337 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n6629) );
  NAND2_X1 U8338 ( .A1(n5182), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6627) );
  INV_X1 U8339 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6624) );
  OR2_X1 U8340 ( .A1(n6625), .A2(n6624), .ZN(n6626) );
  OAI211_X1 U8341 ( .C1(n6629), .C2(n6628), .A(n6627), .B(n6626), .ZN(n6630)
         );
  INV_X1 U8342 ( .A(n6630), .ZN(n6631) );
  INV_X1 U8343 ( .A(n7794), .ZN(n6633) );
  NAND2_X1 U8344 ( .A1(n6633), .A2(P2_U3893), .ZN(n6634) );
  OAI21_X1 U8345 ( .B1(P2_U3893), .B2(n10446), .A(n6634), .ZN(P2_U3522) );
  NAND2_X1 U8346 ( .A1(n6635), .A2(P2_U3893), .ZN(n6636) );
  OAI21_X1 U8347 ( .B1(n7481), .B2(P2_U3893), .A(n6636), .ZN(P2_U3520) );
  INV_X1 U8348 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9848) );
  AOI22_X1 U8349 ( .A1(n7366), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n9848), .B2(
        n6647), .ZN(n6638) );
  OAI21_X1 U8350 ( .B1(n6639), .B2(n6638), .A(n6792), .ZN(n6649) );
  NOR2_X1 U8351 ( .A1(n7366), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6640) );
  AOI21_X1 U8352 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7366), .A(n6640), .ZN(
        n6643) );
  OAI21_X1 U8353 ( .B1(n6643), .B2(n6642), .A(n6796), .ZN(n6644) );
  NAND2_X1 U8354 ( .A1(n6644), .A2(n9230), .ZN(n6646) );
  AND2_X1 U8355 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9048) );
  AOI21_X1 U8356 ( .B1(n9261), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n9048), .ZN(
        n6645) );
  OAI211_X1 U8357 ( .C1(n9258), .C2(n6647), .A(n6646), .B(n6645), .ZN(n6648)
         );
  AOI21_X1 U8358 ( .B1(n9255), .B2(n6649), .A(n6648), .ZN(n6650) );
  INV_X1 U8359 ( .A(n6650), .ZN(P1_U3255) );
  XNOR2_X1 U8360 ( .A(n10045), .B(n8051), .ZN(n6943) );
  XNOR2_X1 U8361 ( .A(n6943), .B(n8438), .ZN(n6654) );
  NAND2_X1 U8362 ( .A1(n6655), .A2(n6654), .ZN(n6946) );
  OAI211_X1 U8363 ( .C1(n6655), .C2(n6654), .A(n6946), .B(n8423), .ZN(n6660)
         );
  OR2_X1 U8364 ( .A1(n8409), .A2(n10026), .ZN(n6656) );
  OR2_X1 U8365 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5348), .ZN(n6811) );
  OAI211_X1 U8366 ( .C1(n8427), .C2(n7186), .A(n6656), .B(n6811), .ZN(n6658)
         );
  NOR2_X1 U8367 ( .A1(n8428), .A2(n6970), .ZN(n6657) );
  AOI211_X1 U8368 ( .C1(n10045), .C2(n8419), .A(n6658), .B(n6657), .ZN(n6659)
         );
  NAND2_X1 U8369 ( .A1(n6660), .A2(n6659), .ZN(P2_U3171) );
  AND2_X1 U8370 ( .A1(n9178), .A2(n6664), .ZN(n6662) );
  INV_X1 U8371 ( .A(n6680), .ZN(n6661) );
  AOI21_X1 U8372 ( .B1(n6662), .B2(n6673), .A(n6661), .ZN(n7210) );
  AOI22_X1 U8373 ( .A1(n9721), .A2(n9178), .B1(n9175), .B2(n9720), .ZN(n6666)
         );
  AOI21_X1 U8374 ( .B1(n7206), .B2(n6664), .A(n9494), .ZN(n6665) );
  NAND2_X1 U8375 ( .A1(n6665), .A2(n6706), .ZN(n7209) );
  OAI211_X1 U8376 ( .C1(n7210), .C2(n9717), .A(n6666), .B(n7209), .ZN(n6668)
         );
  XOR2_X1 U8377 ( .A(n6673), .B(n6672), .Z(n6667) );
  NOR2_X1 U8378 ( .A1(n6667), .A2(n9693), .ZN(n7213) );
  NOR2_X1 U8379 ( .A1(n6668), .A2(n7213), .ZN(n6697) );
  INV_X1 U8380 ( .A(n9831), .ZN(n9712) );
  INV_X1 U8381 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6669) );
  OAI22_X1 U8382 ( .A1(n9783), .A2(n8078), .B1(n9838), .B2(n6669), .ZN(n6670)
         );
  INV_X1 U8383 ( .A(n6670), .ZN(n6671) );
  OAI21_X1 U8384 ( .B1(n6697), .B2(n9836), .A(n6671), .ZN(P1_U3456) );
  NAND2_X1 U8385 ( .A1(n6673), .A2(n6672), .ZN(n6675) );
  NAND2_X1 U8386 ( .A1(n6704), .A2(n7206), .ZN(n6674) );
  XNOR2_X1 U8387 ( .A(n8077), .B(n6676), .ZN(n6702) );
  INV_X1 U8388 ( .A(n6702), .ZN(n8213) );
  NAND2_X1 U8389 ( .A1(n6677), .A2(n6707), .ZN(n6678) );
  INV_X1 U8390 ( .A(n6684), .ZN(n8210) );
  XNOR2_X1 U8391 ( .A(n6735), .B(n8210), .ZN(n7121) );
  OR2_X1 U8392 ( .A1(n7206), .A2(n9177), .ZN(n6679) );
  NAND2_X1 U8393 ( .A1(n6703), .A2(n6702), .ZN(n6701) );
  OR2_X1 U8394 ( .A1(n6707), .A2(n9175), .ZN(n6681) );
  NAND2_X1 U8395 ( .A1(n6701), .A2(n6681), .ZN(n6685) );
  AND2_X1 U8396 ( .A1(n6702), .A2(n6684), .ZN(n6683) );
  NOR2_X1 U8397 ( .A1(n8210), .A2(n6681), .ZN(n6682) );
  OAI21_X1 U8398 ( .B1(n6685), .B2(n6684), .A(n6724), .ZN(n7128) );
  INV_X1 U8399 ( .A(n7128), .ZN(n6687) );
  AOI22_X1 U8400 ( .A1(n9721), .A2(n9175), .B1(n9173), .B2(n9720), .ZN(n6686)
         );
  NAND2_X1 U8401 ( .A1(n6705), .A2(n6722), .ZN(n7012) );
  OAI211_X1 U8402 ( .C1(n6705), .C2(n6722), .A(n7012), .B(n9593), .ZN(n7126)
         );
  OAI211_X1 U8403 ( .C1(n6687), .C2(n9717), .A(n6686), .B(n7126), .ZN(n6688)
         );
  AOI21_X1 U8404 ( .B1(n9713), .B2(n7121), .A(n6688), .ZN(n6694) );
  OAI22_X1 U8405 ( .A1(n9783), .A2(n6722), .B1(n9838), .B2(n6488), .ZN(n6689)
         );
  INV_X1 U8406 ( .A(n6689), .ZN(n6690) );
  OAI21_X1 U8407 ( .B1(n6694), .B2(n9836), .A(n6690), .ZN(P1_U3462) );
  INV_X1 U8408 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6691) );
  OAI22_X1 U8409 ( .A1(n9742), .A2(n6722), .B1(n9850), .B2(n6691), .ZN(n6692)
         );
  INV_X1 U8410 ( .A(n6692), .ZN(n6693) );
  OAI21_X1 U8411 ( .B1(n6694), .B2(n9847), .A(n6693), .ZN(P1_U3525) );
  OAI22_X1 U8412 ( .A1(n9742), .A2(n8078), .B1(n9850), .B2(n4644), .ZN(n6695)
         );
  INV_X1 U8413 ( .A(n6695), .ZN(n6696) );
  OAI21_X1 U8414 ( .B1(n6697), .B2(n9847), .A(n6696), .ZN(P1_U3523) );
  INV_X1 U8415 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10235) );
  INV_X1 U8416 ( .A(n7521), .ZN(n6771) );
  NAND2_X1 U8417 ( .A1(n4598), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6698) );
  XNOR2_X1 U8418 ( .A(n6698), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9241) );
  INV_X1 U8419 ( .A(n9241), .ZN(n6699) );
  OAI222_X1 U8420 ( .A1(n6832), .A2(n10235), .B1(n7300), .B2(n6771), .C1(
        P1_U3086), .C2(n6699), .ZN(P1_U3337) );
  XNOR2_X1 U8421 ( .A(n6700), .B(n6702), .ZN(n7182) );
  OAI21_X1 U8422 ( .B1(n6703), .B2(n6702), .A(n6701), .ZN(n7179) );
  OAI22_X1 U8423 ( .A1(n6704), .A2(n9708), .B1(n8076), .B2(n9731), .ZN(n6708)
         );
  AOI211_X1 U8424 ( .C1(n6707), .C2(n6706), .A(n9494), .B(n6705), .ZN(n7178)
         );
  AOI211_X1 U8425 ( .C1(n9834), .C2(n7179), .A(n6708), .B(n7178), .ZN(n6709)
         );
  OAI21_X1 U8426 ( .B1(n9693), .B2(n7182), .A(n6709), .ZN(n6714) );
  OAI22_X1 U8427 ( .A1(n9783), .A2(n8077), .B1(n9838), .B2(n6449), .ZN(n6710)
         );
  AOI21_X1 U8428 ( .B1(n6714), .B2(n9838), .A(n6710), .ZN(n6711) );
  INV_X1 U8429 ( .A(n6711), .ZN(P1_U3459) );
  INV_X1 U8430 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6712) );
  OAI22_X1 U8431 ( .A1(n9742), .A2(n8077), .B1(n9850), .B2(n6712), .ZN(n6713)
         );
  AOI21_X1 U8432 ( .B1(n6714), .B2(n9850), .A(n6713), .ZN(n6715) );
  INV_X1 U8433 ( .A(n6715), .ZN(P1_U3524) );
  NAND2_X1 U8434 ( .A1(n8745), .A2(n5191), .ZN(n6716) );
  OAI21_X1 U8435 ( .B1(n8788), .B2(n6717), .A(n6716), .ZN(n6720) );
  NOR3_X1 U8436 ( .A1(n8802), .A2(n9978), .A3(n6718), .ZN(n6719) );
  AOI211_X1 U8437 ( .C1(n8802), .C2(P2_REG2_REG_0__SCAN_IN), .A(n6720), .B(
        n6719), .ZN(n6721) );
  OAI21_X1 U8438 ( .B1(n5005), .B2(n8731), .A(n6721), .ZN(P2_U3233) );
  INV_X1 U8439 ( .A(n6722), .ZN(n9016) );
  OR2_X1 U8440 ( .A1(n9016), .A2(n9174), .ZN(n6723) );
  OR2_X1 U8441 ( .A1(n9801), .A2(n9173), .ZN(n6736) );
  NAND2_X1 U8442 ( .A1(n9801), .A2(n9173), .ZN(n8079) );
  NAND2_X1 U8443 ( .A1(n6736), .A2(n8079), .ZN(n8209) );
  NAND2_X1 U8444 ( .A1(n7010), .A2(n8209), .ZN(n7009) );
  OR2_X1 U8445 ( .A1(n7018), .A2(n9173), .ZN(n6725) );
  NAND2_X1 U8446 ( .A1(n7009), .A2(n6725), .ZN(n6732) );
  OR2_X1 U8447 ( .A1(n7534), .A2(n6726), .ZN(n6731) );
  OR2_X1 U8448 ( .A1(n7504), .A2(n6727), .ZN(n6730) );
  OR2_X1 U8449 ( .A1(n7229), .A2(n6728), .ZN(n6729) );
  OR2_X1 U8450 ( .A1(n6844), .A2(n9172), .ZN(n8109) );
  NAND2_X1 U8451 ( .A1(n6844), .A2(n9172), .ZN(n8108) );
  NAND2_X1 U8452 ( .A1(n8109), .A2(n8108), .ZN(n6738) );
  NAND2_X1 U8453 ( .A1(n6732), .A2(n6738), .ZN(n7024) );
  OAI21_X1 U8454 ( .B1(n6732), .B2(n6738), .A(n7024), .ZN(n7224) );
  INV_X1 U8455 ( .A(n9173), .ZN(n7218) );
  OR2_X1 U8456 ( .A1(n7012), .A2(n7018), .ZN(n7013) );
  INV_X1 U8457 ( .A(n7013), .ZN(n6734) );
  INV_X1 U8458 ( .A(n6844), .ZN(n9071) );
  INV_X1 U8459 ( .A(n7078), .ZN(n6733) );
  OAI211_X1 U8460 ( .C1(n6844), .C2(n6734), .A(n6733), .B(n9593), .ZN(n7222)
         );
  OAI21_X1 U8461 ( .B1(n7218), .B2(n9708), .A(n7222), .ZN(n6748) );
  INV_X1 U8462 ( .A(n6736), .ZN(n6737) );
  INV_X1 U8463 ( .A(n6738), .ZN(n8212) );
  XNOR2_X1 U8464 ( .A(n7046), .B(n8212), .ZN(n6747) );
  NAND2_X1 U8465 ( .A1(n4513), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6746) );
  INV_X1 U8466 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6739) );
  OR2_X1 U8467 ( .A1(n4602), .A2(n6739), .ZN(n6745) );
  INV_X1 U8468 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6740) );
  NAND2_X1 U8469 ( .A1(n6741), .A2(n6740), .ZN(n6742) );
  NAND2_X1 U8470 ( .A1(n6864), .A2(n6742), .ZN(n7080) );
  OR2_X1 U8471 ( .A1(n7988), .A2(n7080), .ZN(n6744) );
  OR2_X1 U8472 ( .A1(n7981), .A2(n7081), .ZN(n6743) );
  NAND4_X1 U8473 ( .A1(n6746), .A2(n6745), .A3(n6744), .A4(n6743), .ZN(n9171)
         );
  INV_X1 U8474 ( .A(n9171), .ZN(n7090) );
  OAI22_X1 U8475 ( .A1(n6747), .A2(n9693), .B1(n7090), .B2(n9731), .ZN(n7216)
         );
  AOI211_X1 U8476 ( .C1(n9834), .C2(n7224), .A(n6748), .B(n7216), .ZN(n6754)
         );
  OAI22_X1 U8477 ( .A1(n9783), .A2(n6844), .B1(n9838), .B2(n6571), .ZN(n6749)
         );
  INV_X1 U8478 ( .A(n6749), .ZN(n6750) );
  OAI21_X1 U8479 ( .B1(n6754), .B2(n9836), .A(n6750), .ZN(P1_U3468) );
  INV_X1 U8480 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6751) );
  OAI22_X1 U8481 ( .A1(n9742), .A2(n6844), .B1(n9850), .B2(n6751), .ZN(n6752)
         );
  INV_X1 U8482 ( .A(n6752), .ZN(n6753) );
  OAI21_X1 U8483 ( .B1(n6754), .B2(n9847), .A(n6753), .ZN(P1_U3527) );
  AND2_X1 U8484 ( .A1(n6755), .A2(n6998), .ZN(n7597) );
  INV_X1 U8485 ( .A(n7597), .ZN(n6756) );
  XNOR2_X1 U8486 ( .A(n6757), .B(n6756), .ZN(n6758) );
  NAND2_X1 U8487 ( .A1(n6758), .A2(n10005), .ZN(n6760) );
  AOI22_X1 U8488 ( .A1(n10043), .A2(n8441), .B1(n8439), .B2(n10042), .ZN(n6759) );
  NAND2_X1 U8489 ( .A1(n6760), .A2(n6759), .ZN(n10023) );
  INV_X1 U8490 ( .A(n10023), .ZN(n6770) );
  NAND2_X1 U8491 ( .A1(n6761), .A2(n7660), .ZN(n6762) );
  XNOR2_X1 U8492 ( .A(n6762), .B(n7597), .ZN(n10020) );
  AND2_X1 U8493 ( .A1(n9988), .A2(n6763), .ZN(n6764) );
  NOR2_X1 U8494 ( .A1(n8728), .A2(n6508), .ZN(n6768) );
  INV_X1 U8495 ( .A(n8757), .ZN(n8791) );
  OAI22_X1 U8496 ( .A1(n8791), .A2(n6766), .B1(n6765), .B2(n8788), .ZN(n6767)
         );
  AOI211_X1 U8497 ( .C1(n10020), .C2(n8793), .A(n6768), .B(n6767), .ZN(n6769)
         );
  OAI21_X1 U8498 ( .B1(n6770), .B2(n8802), .A(n6769), .ZN(P2_U3227) );
  INV_X1 U8499 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6772) );
  INV_X1 U8500 ( .A(n8558), .ZN(n8544) );
  OAI222_X1 U8501 ( .A1(n8991), .A2(n6772), .B1(n8544), .B2(P2_U3151), .C1(
        n8990), .C2(n6771), .ZN(P2_U3277) );
  XNOR2_X1 U8502 ( .A(n6773), .B(n7590), .ZN(n9993) );
  XNOR2_X1 U8503 ( .A(n7635), .B(n6774), .ZN(n6775) );
  NOR2_X1 U8504 ( .A1(n6775), .A2(n9979), .ZN(n9990) );
  OAI22_X1 U8505 ( .A1(n9989), .A2(n8778), .B1(n9874), .B2(n8788), .ZN(n6776)
         );
  NOR2_X1 U8506 ( .A1(n9990), .A2(n6776), .ZN(n6777) );
  MUX2_X1 U8507 ( .A(n6778), .B(n6777), .S(n8728), .Z(n6780) );
  NAND2_X1 U8508 ( .A1(n8728), .A2(n10043), .ZN(n8712) );
  INV_X1 U8509 ( .A(n8712), .ZN(n8797) );
  AOI22_X1 U8510 ( .A1(n8797), .A2(n5870), .B1(n8795), .B2(n10008), .ZN(n6779)
         );
  OAI211_X1 U8511 ( .C1(n8784), .C2(n9993), .A(n6780), .B(n6779), .ZN(P2_U3231) );
  NAND2_X1 U8512 ( .A1(n7652), .A2(n7670), .ZN(n7599) );
  NAND2_X1 U8513 ( .A1(n6993), .A2(n6781), .ZN(n6782) );
  XOR2_X1 U8514 ( .A(n7599), .B(n6782), .Z(n10038) );
  XNOR2_X1 U8515 ( .A(n6783), .B(n7599), .ZN(n6784) );
  OAI222_X1 U8516 ( .A1(n10027), .A2(n6785), .B1(n10025), .B2(n6947), .C1(
        n6784), .C2(n9979), .ZN(n10040) );
  NAND2_X1 U8517 ( .A1(n10040), .A2(n8728), .ZN(n6791) );
  OAI22_X1 U8518 ( .A1(n8728), .A2(n6787), .B1(n6786), .B2(n8788), .ZN(n6788)
         );
  AOI21_X1 U8519 ( .B1(n8757), .B2(n6789), .A(n6788), .ZN(n6790) );
  OAI211_X1 U8520 ( .C1(n10038), .C2(n8784), .A(n6791), .B(n6790), .ZN(
        P2_U3225) );
  OAI21_X1 U8521 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n7366), .A(n6792), .ZN(
        n6795) );
  INV_X1 U8522 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6793) );
  MUX2_X1 U8523 ( .A(n6793), .B(P1_REG1_REG_13__SCAN_IN), .S(n7506), .Z(n6794)
         );
  NOR2_X1 U8524 ( .A1(n6794), .A2(n6795), .ZN(n6956) );
  AOI211_X1 U8525 ( .C1(n6795), .C2(n6794), .A(n6956), .B(n9254), .ZN(n6804)
         );
  OAI21_X1 U8526 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7366), .A(n6796), .ZN(
        n6799) );
  NAND2_X1 U8527 ( .A1(n7506), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6797) );
  OAI21_X1 U8528 ( .B1(n7506), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6797), .ZN(
        n6798) );
  NOR2_X1 U8529 ( .A1(n6798), .A2(n6799), .ZN(n6959) );
  AOI211_X1 U8530 ( .C1(n6799), .C2(n6798), .A(n6959), .B(n9259), .ZN(n6803)
         );
  INV_X1 U8531 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6801) );
  NAND2_X1 U8532 ( .A1(n9236), .A2(n7506), .ZN(n6800) );
  NAND2_X1 U8533 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9120) );
  OAI211_X1 U8534 ( .C1(n6801), .C2(n9234), .A(n6800), .B(n9120), .ZN(n6802)
         );
  OR3_X1 U8535 ( .A1(n6804), .A2(n6803), .A3(n6802), .ZN(P1_U3256) );
  INV_X1 U8536 ( .A(n8461), .ZN(n6806) );
  MUX2_X1 U8537 ( .A(n6787), .B(P2_REG2_REG_8__SCAN_IN), .S(n8450), .Z(n8460)
         );
  INV_X1 U8538 ( .A(n8460), .ZN(n6805) );
  AOI21_X1 U8539 ( .B1(n6806), .B2(n8458), .A(n6805), .ZN(n8463) );
  AOI21_X1 U8540 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n6814), .A(n8463), .ZN(
        n6891) );
  AOI21_X1 U8541 ( .B1(n6807), .B2(n6971), .A(n6893), .ZN(n6830) );
  INV_X1 U8542 ( .A(n8455), .ZN(n6809) );
  INV_X1 U8543 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6808) );
  MUX2_X1 U8544 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6808), .S(n8450), .Z(n8451)
         );
  AOI21_X2 U8545 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n6814), .A(n8457), .ZN(
        n6877) );
  XOR2_X1 U8546 ( .A(n6877), .B(n6882), .Z(n6810) );
  AOI21_X1 U8547 ( .B1(n5352), .B2(n6810), .A(n6878), .ZN(n6827) );
  INV_X1 U8548 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n6812) );
  OAI21_X1 U8549 ( .B1(n9888), .B2(n6812), .A(n6811), .ZN(n6813) );
  AOI21_X1 U8550 ( .B1(n8492), .B2(n6892), .A(n6813), .ZN(n6826) );
  MUX2_X1 U8551 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8561), .Z(n6883) );
  XNOR2_X1 U8552 ( .A(n6883), .B(n6892), .ZN(n6823) );
  MUX2_X1 U8553 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8561), .Z(n6820) );
  OR2_X1 U8554 ( .A1(n6820), .A2(n6814), .ZN(n6821) );
  INV_X1 U8555 ( .A(n6815), .ZN(n6817) );
  OAI22_X1 U8556 ( .A1(n6819), .A2(n6818), .B1(n6817), .B2(n6816), .ZN(n8445)
         );
  XNOR2_X1 U8557 ( .A(n6820), .B(n8450), .ZN(n8444) );
  NAND2_X1 U8558 ( .A1(n8445), .A2(n8444), .ZN(n8443) );
  NAND2_X1 U8559 ( .A1(n6821), .A2(n8443), .ZN(n6822) );
  NAND2_X1 U8560 ( .A1(n6823), .A2(n6822), .ZN(n6884) );
  OAI21_X1 U8561 ( .B1(n6823), .B2(n6822), .A(n6884), .ZN(n6824) );
  NAND2_X1 U8562 ( .A1(n6824), .A2(n9967), .ZN(n6825) );
  OAI211_X1 U8563 ( .C1(n6827), .C2(n9971), .A(n6826), .B(n6825), .ZN(n6828)
         );
  INV_X1 U8564 ( .A(n6828), .ZN(n6829) );
  OAI21_X1 U8565 ( .B1(n6830), .B2(n9963), .A(n6829), .ZN(P2_U3191) );
  INV_X1 U8566 ( .A(n7524), .ZN(n6833) );
  OAI222_X1 U8567 ( .A1(n8991), .A2(n6831), .B1(n8990), .B2(n6833), .C1(n5139), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  OAI222_X1 U8568 ( .A1(n9343), .A2(P1_U3086), .B1(n7300), .B2(n6833), .C1(
        n10247), .C2(n6832), .ZN(P1_U3336) );
  INV_X1 U8569 ( .A(n6834), .ZN(n6836) );
  NAND2_X1 U8570 ( .A1(n6836), .A2(n6835), .ZN(n6837) );
  NAND2_X1 U8571 ( .A1(n6838), .A2(n6837), .ZN(n6842) );
  NAND2_X1 U8572 ( .A1(n9172), .A2(n6541), .ZN(n6839) );
  OAI21_X1 U8573 ( .B1(n6844), .B2(n7883), .A(n6839), .ZN(n6840) );
  XNOR2_X1 U8574 ( .A(n6840), .B(n7998), .ZN(n6841) );
  NAND2_X1 U8575 ( .A1(n6842), .A2(n6841), .ZN(n6843) );
  OR2_X1 U8576 ( .A1(n6844), .A2(n7307), .ZN(n6846) );
  NAND2_X1 U8577 ( .A1(n9172), .A2(n7959), .ZN(n6845) );
  AND2_X1 U8578 ( .A1(n6846), .A2(n6845), .ZN(n9069) );
  OR2_X1 U8579 ( .A1(n7504), .A2(n6848), .ZN(n6853) );
  OR2_X1 U8580 ( .A1(n7534), .A2(n6849), .ZN(n6852) );
  OR2_X1 U8581 ( .A1(n4512), .A2(n6850), .ZN(n6851) );
  NAND2_X1 U8582 ( .A1(n9171), .A2(n6541), .ZN(n6854) );
  OAI21_X1 U8583 ( .B1(n9806), .B2(n7883), .A(n6854), .ZN(n6855) );
  XNOR2_X1 U8584 ( .A(n6855), .B(n7998), .ZN(n6858) );
  OR2_X1 U8585 ( .A1(n9806), .A2(n7307), .ZN(n6857) );
  NAND2_X1 U8586 ( .A1(n9171), .A2(n7959), .ZN(n6856) );
  NAND2_X1 U8587 ( .A1(n6857), .A2(n6856), .ZN(n6859) );
  NAND2_X1 U8588 ( .A1(n6858), .A2(n6859), .ZN(n7105) );
  INV_X1 U8589 ( .A(n6858), .ZN(n6861) );
  INV_X1 U8590 ( .A(n6859), .ZN(n6860) );
  NAND2_X1 U8591 ( .A1(n6861), .A2(n6860), .ZN(n7107) );
  NAND2_X1 U8592 ( .A1(n7105), .A2(n7107), .ZN(n6862) );
  XNOR2_X1 U8593 ( .A(n7106), .B(n6862), .ZN(n6876) );
  NAND2_X1 U8594 ( .A1(n4513), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6870) );
  INV_X1 U8595 ( .A(n7981), .ZN(n7798) );
  OR2_X1 U8596 ( .A1(n7907), .A2(n7099), .ZN(n6869) );
  INV_X1 U8597 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6863) );
  NAND2_X1 U8598 ( .A1(n6864), .A2(n6863), .ZN(n6865) );
  NAND2_X1 U8599 ( .A1(n7040), .A2(n6865), .ZN(n7115) );
  OR2_X1 U8600 ( .A1(n7988), .A2(n7115), .ZN(n6868) );
  INV_X1 U8601 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6866) );
  OR2_X1 U8602 ( .A1(n4602), .A2(n6866), .ZN(n6867) );
  NAND4_X1 U8603 ( .A1(n6870), .A2(n6869), .A3(n6868), .A4(n6867), .ZN(n9170)
         );
  INV_X1 U8604 ( .A(n9806), .ZN(n7083) );
  AOI22_X1 U8605 ( .A1(n9072), .A2(n9170), .B1(n7083), .B2(n9162), .ZN(n6875)
         );
  INV_X1 U8606 ( .A(n6871), .ZN(n6873) );
  NOR2_X1 U8607 ( .A1(n9157), .A2(n7080), .ZN(n6872) );
  AOI211_X1 U8608 ( .C1(n9077), .C2(n9172), .A(n6873), .B(n6872), .ZN(n6874)
         );
  OAI211_X1 U8609 ( .C1(n6876), .C2(n9164), .A(n6875), .B(n6874), .ZN(P1_U3239) );
  NOR2_X1 U8610 ( .A1(n6892), .A2(n6877), .ZN(n6879) );
  AOI22_X1 U8611 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n6895), .B1(n7140), .B2(
        n5373), .ZN(n6880) );
  AOI21_X1 U8612 ( .B1(n6881), .B2(n6880), .A(n7131), .ZN(n6903) );
  MUX2_X1 U8613 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8561), .Z(n7141) );
  XNOR2_X1 U8614 ( .A(n7141), .B(n6895), .ZN(n6887) );
  OR2_X1 U8615 ( .A1(n6883), .A2(n6882), .ZN(n6885) );
  NAND2_X1 U8616 ( .A1(n6885), .A2(n6884), .ZN(n6886) );
  NAND2_X1 U8617 ( .A1(n6887), .A2(n6886), .ZN(n7142) );
  OAI21_X1 U8618 ( .B1(n6887), .B2(n6886), .A(n7142), .ZN(n6901) );
  INV_X1 U8619 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n6890) );
  NAND2_X1 U8620 ( .A1(n8492), .A2(n6895), .ZN(n6889) );
  INV_X1 U8621 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10397) );
  NOR2_X1 U8622 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10397), .ZN(n6949) );
  INV_X1 U8623 ( .A(n6949), .ZN(n6888) );
  OAI211_X1 U8624 ( .C1(n6890), .C2(n9888), .A(n6889), .B(n6888), .ZN(n6900)
         );
  NOR2_X1 U8625 ( .A1(n6892), .A2(n6891), .ZN(n6894) );
  MUX2_X1 U8626 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n6896), .S(n6895), .Z(n6897)
         );
  AOI21_X1 U8627 ( .B1(n4597), .B2(n6897), .A(n7134), .ZN(n6898) );
  NOR2_X1 U8628 ( .A1(n6898), .A2(n9963), .ZN(n6899) );
  AOI211_X1 U8629 ( .C1(n9967), .C2(n6901), .A(n6900), .B(n6899), .ZN(n6902)
         );
  OAI21_X1 U8630 ( .B1(n6903), .B2(n9971), .A(n6902), .ZN(P2_U3192) );
  AND2_X1 U8631 ( .A1(n6905), .A2(n6904), .ZN(n6906) );
  NAND4_X1 U8632 ( .A1(n6908), .A2(n6907), .A3(n8271), .A4(n6906), .ZN(n6909)
         );
  AOI21_X1 U8633 ( .B1(n9593), .B2(n9538), .A(n9569), .ZN(n6918) );
  OAI22_X1 U8634 ( .A1(n9598), .A2(n5930), .B1(n6911), .B2(n9557), .ZN(n6915)
         );
  INV_X1 U8635 ( .A(n6912), .ZN(n6913) );
  NOR4_X1 U8636 ( .A1(n4528), .A2(n9585), .A3(n8270), .A4(n6913), .ZN(n6914)
         );
  AOI211_X1 U8637 ( .C1(n9587), .C2(n9177), .A(n6915), .B(n6914), .ZN(n6916)
         );
  OAI21_X1 U8638 ( .B1(n6918), .B2(n6917), .A(n6916), .ZN(P1_U3293) );
  XNOR2_X1 U8639 ( .A(n6920), .B(n6919), .ZN(n10003) );
  INV_X1 U8640 ( .A(n10003), .ZN(n6929) );
  INV_X1 U8641 ( .A(n8684), .ZN(n8720) );
  OAI21_X1 U8642 ( .B1(n6922), .B2(n7592), .A(n6921), .ZN(n9996) );
  AOI22_X1 U8643 ( .A1(n8797), .A2(n9998), .B1(n8795), .B2(n8442), .ZN(n6925)
         );
  NOR2_X1 U8644 ( .A1(n8788), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6923) );
  AOI21_X1 U8645 ( .B1(n8745), .B2(n9997), .A(n6923), .ZN(n6924) );
  OAI211_X1 U8646 ( .C1(n6926), .C2(n8728), .A(n6925), .B(n6924), .ZN(n6927)
         );
  AOI21_X1 U8647 ( .B1(n8793), .B2(n9996), .A(n6927), .ZN(n6928) );
  OAI21_X1 U8648 ( .B1(n6929), .B2(n8720), .A(n6928), .ZN(P2_U3230) );
  INV_X1 U8649 ( .A(n7529), .ZN(n6967) );
  AOI21_X1 U8650 ( .B1(P2_DATAO_REG_20__SCAN_IN), .B2(n6931), .A(n6930), .ZN(
        n6932) );
  OAI21_X1 U8651 ( .B1(n6967), .B2(n7300), .A(n6932), .ZN(P1_U3335) );
  XNOR2_X1 U8652 ( .A(n4511), .B(n7642), .ZN(n10013) );
  INV_X1 U8653 ( .A(n10013), .ZN(n6942) );
  OAI22_X1 U8654 ( .A1(n8791), .A2(n6935), .B1(n6934), .B2(n8788), .ZN(n6938)
         );
  OAI22_X1 U8655 ( .A1(n8731), .A2(n10011), .B1(n6936), .B2(n8712), .ZN(n6937)
         );
  AOI211_X1 U8656 ( .C1(P2_REG2_REG_4__SCAN_IN), .C2(n8802), .A(n6938), .B(
        n6937), .ZN(n6941) );
  XNOR2_X1 U8657 ( .A(n6939), .B(n7591), .ZN(n10006) );
  NAND2_X1 U8658 ( .A1(n10006), .A2(n8684), .ZN(n6940) );
  OAI211_X1 U8659 ( .C1(n6942), .C2(n8784), .A(n6941), .B(n6940), .ZN(P2_U3229) );
  XNOR2_X1 U8660 ( .A(n10059), .B(n5869), .ZN(n7164) );
  INV_X1 U8661 ( .A(n6943), .ZN(n6944) );
  NAND2_X1 U8662 ( .A1(n6944), .A2(n8438), .ZN(n6945) );
  XOR2_X1 U8663 ( .A(n7164), .B(n7165), .Z(n6953) );
  NOR2_X1 U8664 ( .A1(n8409), .A2(n6947), .ZN(n6948) );
  AOI211_X1 U8665 ( .C1(n8406), .C2(n8437), .A(n6949), .B(n6948), .ZN(n6950)
         );
  OAI21_X1 U8666 ( .B1(n6988), .B2(n8428), .A(n6950), .ZN(n6951) );
  AOI21_X1 U8667 ( .B1(n10059), .B2(n8419), .A(n6951), .ZN(n6952) );
  OAI21_X1 U8668 ( .B1(n6953), .B2(n8421), .A(n6952), .ZN(P2_U3157) );
  INV_X1 U8669 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n6955) );
  NAND2_X1 U8670 ( .A1(n9236), .A2(n9187), .ZN(n6954) );
  NAND2_X1 U8671 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9001) );
  OAI211_X1 U8672 ( .C1(n6955), .C2(n9234), .A(n6954), .B(n9001), .ZN(n6966)
         );
  XNOR2_X1 U8673 ( .A(n9187), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n6957) );
  AOI211_X1 U8674 ( .C1(n6958), .C2(n6957), .A(n9179), .B(n9254), .ZN(n6965)
         );
  INV_X1 U8675 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6960) );
  MUX2_X1 U8676 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n6960), .S(n9187), .Z(n6961)
         );
  INV_X1 U8677 ( .A(n6961), .ZN(n6962) );
  AOI211_X1 U8678 ( .C1(n6963), .C2(n6962), .A(n9186), .B(n9259), .ZN(n6964)
         );
  OR3_X1 U8679 ( .A1(n6966), .A2(n6965), .A3(n6964), .ZN(P1_U3257) );
  OAI222_X1 U8680 ( .A1(n8990), .A2(n6967), .B1(n8991), .B2(n5551), .C1(n7782), 
        .C2(P2_U3151), .ZN(P2_U3275) );
  XNOR2_X1 U8681 ( .A(n6968), .B(n7601), .ZN(n6969) );
  NAND2_X1 U8682 ( .A1(n6969), .A2(n10005), .ZN(n10049) );
  OAI22_X1 U8683 ( .A1(n8728), .A2(n6971), .B1(n6970), .B2(n8788), .ZN(n6972)
         );
  AOI21_X1 U8684 ( .B1(n8797), .B2(n10044), .A(n6972), .ZN(n6973) );
  OAI21_X1 U8685 ( .B1(n7186), .B2(n8731), .A(n6973), .ZN(n6978) );
  NAND2_X1 U8686 ( .A1(n6975), .A2(n7601), .ZN(n6976) );
  NAND2_X1 U8687 ( .A1(n6974), .A2(n6976), .ZN(n10048) );
  NOR2_X1 U8688 ( .A1(n10048), .A2(n8784), .ZN(n6977) );
  AOI211_X1 U8689 ( .C1(n8757), .C2(n10045), .A(n6978), .B(n6977), .ZN(n6979)
         );
  OAI21_X1 U8690 ( .B1(n8802), .B2(n10049), .A(n6979), .ZN(P2_U3224) );
  NAND2_X1 U8691 ( .A1(n7679), .A2(n7678), .ZN(n7600) );
  INV_X1 U8692 ( .A(n7600), .ZN(n6980) );
  XNOR2_X1 U8693 ( .A(n6981), .B(n6980), .ZN(n10056) );
  INV_X1 U8694 ( .A(n10056), .ZN(n6986) );
  XOR2_X1 U8695 ( .A(n7600), .B(n6982), .Z(n6983) );
  NAND2_X1 U8696 ( .A1(n6983), .A2(n10005), .ZN(n6985) );
  AOI22_X1 U8697 ( .A1(n10043), .A2(n8438), .B1(n8437), .B2(n10042), .ZN(n6984) );
  OAI211_X1 U8698 ( .C1(n10056), .C2(n9988), .A(n6985), .B(n6984), .ZN(n10057)
         );
  AOI21_X1 U8699 ( .B1(n6987), .B2(n6986), .A(n10057), .ZN(n6991) );
  OAI22_X1 U8700 ( .A1(n8728), .A2(n6896), .B1(n6988), .B2(n8788), .ZN(n6989)
         );
  AOI21_X1 U8701 ( .B1(n10059), .B2(n8745), .A(n6989), .ZN(n6990) );
  OAI21_X1 U8702 ( .B1(n6991), .B2(n8802), .A(n6990), .ZN(P2_U3223) );
  INV_X1 U8703 ( .A(n6993), .ZN(n6994) );
  AOI21_X1 U8704 ( .B1(n7596), .B2(n6992), .A(n6994), .ZN(n10035) );
  INV_X1 U8705 ( .A(n10035), .ZN(n10032) );
  OAI22_X1 U8706 ( .A1(n8728), .A2(n6500), .B1(n6995), .B2(n8788), .ZN(n6997)
         );
  OAI22_X1 U8707 ( .A1(n8731), .A2(n10026), .B1(n10028), .B2(n8712), .ZN(n6996) );
  AOI211_X1 U8708 ( .C1(n8745), .C2(n10030), .A(n6997), .B(n6996), .ZN(n7003)
         );
  NAND2_X1 U8709 ( .A1(n6999), .A2(n6998), .ZN(n7000) );
  XNOR2_X1 U8710 ( .A(n7000), .B(n7596), .ZN(n7001) );
  NOR2_X1 U8711 ( .A1(n7001), .A2(n9979), .ZN(n10033) );
  NAND2_X1 U8712 ( .A1(n10033), .A2(n8728), .ZN(n7002) );
  OAI211_X1 U8713 ( .C1(n10032), .C2(n8784), .A(n7003), .B(n7002), .ZN(
        P2_U3226) );
  INV_X1 U8714 ( .A(n8209), .ZN(n7004) );
  XNOR2_X1 U8715 ( .A(n7005), .B(n7004), .ZN(n7006) );
  NAND2_X1 U8716 ( .A1(n7006), .A2(n9713), .ZN(n7008) );
  AOI22_X1 U8717 ( .A1(n9721), .A2(n9174), .B1(n9172), .B2(n9720), .ZN(n7007)
         );
  NAND2_X1 U8718 ( .A1(n7008), .A2(n7007), .ZN(n9802) );
  INV_X1 U8719 ( .A(n9802), .ZN(n7022) );
  OAI21_X1 U8720 ( .B1(n7010), .B2(n8209), .A(n7009), .ZN(n9804) );
  NAND2_X1 U8721 ( .A1(n7355), .A2(n7063), .ZN(n7011) );
  INV_X1 U8722 ( .A(n7012), .ZN(n7014) );
  OAI211_X1 U8723 ( .C1(n7014), .C2(n9801), .A(n9593), .B(n7013), .ZN(n9800)
         );
  OAI22_X1 U8724 ( .A1(n9598), .A2(n7016), .B1(n7015), .B2(n9557), .ZN(n7017)
         );
  AOI21_X1 U8725 ( .B1(n9569), .B2(n7018), .A(n7017), .ZN(n7019) );
  OAI21_X1 U8726 ( .B1(n9800), .B2(n9595), .A(n7019), .ZN(n7020) );
  AOI21_X1 U8727 ( .B1(n9804), .B2(n9556), .A(n7020), .ZN(n7021) );
  OAI21_X1 U8728 ( .B1(n7022), .B2(n9585), .A(n7021), .ZN(P1_U3289) );
  OR2_X1 U8729 ( .A1(n9071), .A2(n9172), .ZN(n7023) );
  NAND2_X1 U8730 ( .A1(n7024), .A2(n7023), .ZN(n7077) );
  OR2_X1 U8731 ( .A1(n9806), .A2(n9171), .ZN(n8207) );
  NAND2_X1 U8732 ( .A1(n9806), .A2(n9171), .ZN(n8112) );
  NAND2_X1 U8733 ( .A1(n8207), .A2(n8112), .ZN(n7076) );
  NAND2_X1 U8734 ( .A1(n7077), .A2(n7076), .ZN(n7075) );
  OR2_X1 U8735 ( .A1(n7083), .A2(n9171), .ZN(n7025) );
  NAND2_X1 U8736 ( .A1(n7075), .A2(n7025), .ZN(n7089) );
  OR2_X1 U8737 ( .A1(n7504), .A2(n7026), .ZN(n7031) );
  OR2_X1 U8738 ( .A1(n7534), .A2(n7027), .ZN(n7030) );
  OR2_X1 U8739 ( .A1(n7229), .A2(n7028), .ZN(n7029) );
  XNOR2_X1 U8740 ( .A(n7260), .B(n9170), .ZN(n8115) );
  NAND2_X1 U8741 ( .A1(n7089), .A2(n8115), .ZN(n7088) );
  INV_X1 U8742 ( .A(n7260), .ZN(n7113) );
  OR2_X1 U8743 ( .A1(n7113), .A2(n9170), .ZN(n7032) );
  NAND2_X1 U8744 ( .A1(n7033), .A2(n4514), .ZN(n7037) );
  OR2_X1 U8745 ( .A1(n4512), .A2(n7034), .ZN(n7036) );
  OR2_X1 U8746 ( .A1(n7534), .A2(n10478), .ZN(n7035) );
  NAND2_X1 U8747 ( .A1(n4513), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7045) );
  INV_X1 U8748 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7038) );
  OR2_X1 U8749 ( .A1(n4602), .A2(n7038), .ZN(n7044) );
  NAND2_X1 U8750 ( .A1(n7040), .A2(n7039), .ZN(n7041) );
  NAND2_X1 U8751 ( .A1(n7054), .A2(n7041), .ZN(n7314) );
  OR2_X1 U8752 ( .A1(n7988), .A2(n7314), .ZN(n7043) );
  OR2_X1 U8753 ( .A1(n7907), .A2(n7066), .ZN(n7042) );
  NAND4_X1 U8754 ( .A1(n7045), .A2(n7044), .A3(n7043), .A4(n7042), .ZN(n9169)
         );
  NAND2_X1 U8755 ( .A1(n9811), .A2(n9169), .ZN(n8123) );
  INV_X1 U8756 ( .A(n9169), .ZN(n7399) );
  NAND2_X1 U8757 ( .A1(n7399), .A2(n7318), .ZN(n8121) );
  XNOR2_X1 U8758 ( .A(n7236), .B(n7235), .ZN(n9814) );
  INV_X1 U8759 ( .A(n7355), .ZN(n7096) );
  NAND2_X1 U8760 ( .A1(n7046), .A2(n8212), .ZN(n7047) );
  NAND2_X1 U8761 ( .A1(n7071), .A2(n8207), .ZN(n8086) );
  NAND2_X1 U8762 ( .A1(n8086), .A2(n8112), .ZN(n7091) );
  OR2_X1 U8763 ( .A1(n7091), .A2(n8115), .ZN(n7093) );
  OR2_X1 U8764 ( .A1(n7260), .A2(n9170), .ZN(n7256) );
  NAND2_X1 U8765 ( .A1(n7093), .A2(n7256), .ZN(n7049) );
  INV_X1 U8766 ( .A(n7235), .ZN(n7048) );
  NAND2_X1 U8767 ( .A1(n7049), .A2(n7048), .ZN(n7051) );
  AND2_X1 U8768 ( .A1(n7235), .A2(n7256), .ZN(n7050) );
  NAND2_X1 U8769 ( .A1(n7093), .A2(n7050), .ZN(n7227) );
  NAND3_X1 U8770 ( .A1(n7051), .A2(n9713), .A3(n7227), .ZN(n7061) );
  NAND2_X1 U8771 ( .A1(n7989), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7059) );
  OR2_X1 U8772 ( .A1(n7992), .A2(n7052), .ZN(n7058) );
  INV_X1 U8773 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7053) );
  NAND2_X1 U8774 ( .A1(n7054), .A2(n7053), .ZN(n7055) );
  NAND2_X1 U8775 ( .A1(n7241), .A2(n7055), .ZN(n7398) );
  OR2_X1 U8776 ( .A1(n7988), .A2(n7398), .ZN(n7057) );
  OR2_X1 U8777 ( .A1(n7981), .A2(n6203), .ZN(n7056) );
  INV_X1 U8778 ( .A(n7428), .ZN(n9168) );
  AOI22_X1 U8779 ( .A1(n9168), .A2(n9720), .B1(n9721), .B2(n9170), .ZN(n7060)
         );
  NAND2_X1 U8780 ( .A1(n7061), .A2(n7060), .ZN(n7062) );
  AOI21_X1 U8781 ( .B1(n9814), .B2(n7096), .A(n7062), .ZN(n9816) );
  INV_X1 U8782 ( .A(n7063), .ZN(n7064) );
  NAND2_X1 U8783 ( .A1(n9598), .A2(n7064), .ZN(n7361) );
  INV_X1 U8784 ( .A(n7361), .ZN(n7103) );
  AND2_X1 U8785 ( .A1(n7078), .A2(n9806), .ZN(n7098) );
  AOI21_X1 U8786 ( .B1(n7097), .B2(n7318), .A(n9494), .ZN(n7065) );
  NAND2_X1 U8787 ( .A1(n7065), .A2(n7279), .ZN(n9810) );
  OAI22_X1 U8788 ( .A1(n9598), .A2(n7066), .B1(n7314), .B2(n9557), .ZN(n7067)
         );
  AOI21_X1 U8789 ( .B1(n9569), .B2(n7318), .A(n7067), .ZN(n7068) );
  OAI21_X1 U8790 ( .B1(n9810), .B2(n9595), .A(n7068), .ZN(n7069) );
  AOI21_X1 U8791 ( .B1(n9814), .B2(n7103), .A(n7069), .ZN(n7070) );
  OAI21_X1 U8792 ( .B1(n9816), .B2(n9585), .A(n7070), .ZN(P1_U3285) );
  XNOR2_X1 U8793 ( .A(n7071), .B(n7076), .ZN(n7072) );
  NAND2_X1 U8794 ( .A1(n7072), .A2(n9713), .ZN(n7074) );
  AOI22_X1 U8795 ( .A1(n9720), .A2(n9170), .B1(n9172), .B2(n9721), .ZN(n7073)
         );
  NAND2_X1 U8796 ( .A1(n7074), .A2(n7073), .ZN(n9807) );
  INV_X1 U8797 ( .A(n9807), .ZN(n7087) );
  OAI21_X1 U8798 ( .B1(n7077), .B2(n7076), .A(n7075), .ZN(n9809) );
  OAI21_X1 U8799 ( .B1(n7078), .B2(n9806), .A(n9593), .ZN(n7079) );
  OR2_X1 U8800 ( .A1(n7098), .A2(n7079), .ZN(n9805) );
  OAI22_X1 U8801 ( .A1(n9598), .A2(n7081), .B1(n7080), .B2(n9557), .ZN(n7082)
         );
  AOI21_X1 U8802 ( .B1(n9569), .B2(n7083), .A(n7082), .ZN(n7084) );
  OAI21_X1 U8803 ( .B1(n9805), .B2(n9595), .A(n7084), .ZN(n7085) );
  AOI21_X1 U8804 ( .B1(n9809), .B2(n9556), .A(n7085), .ZN(n7086) );
  OAI21_X1 U8805 ( .B1(n7087), .B2(n9585), .A(n7086), .ZN(P1_U3287) );
  OAI21_X1 U8806 ( .B1(n7089), .B2(n8115), .A(n7088), .ZN(n7193) );
  OAI22_X1 U8807 ( .A1(n7399), .A2(n9731), .B1(n7090), .B2(n9708), .ZN(n7095)
         );
  NAND2_X1 U8808 ( .A1(n7091), .A2(n8115), .ZN(n7092) );
  AOI21_X1 U8809 ( .B1(n7093), .B2(n7092), .A(n9693), .ZN(n7094) );
  AOI211_X1 U8810 ( .C1(n7096), .C2(n7193), .A(n7095), .B(n7094), .ZN(n7195)
         );
  OAI211_X1 U8811 ( .C1(n7260), .C2(n7098), .A(n7097), .B(n9593), .ZN(n7194)
         );
  OAI22_X1 U8812 ( .A1(n9598), .A2(n7099), .B1(n7115), .B2(n9557), .ZN(n7100)
         );
  AOI21_X1 U8813 ( .B1(n9569), .B2(n7113), .A(n7100), .ZN(n7101) );
  OAI21_X1 U8814 ( .B1(n7194), .B2(n9595), .A(n7101), .ZN(n7102) );
  AOI21_X1 U8815 ( .B1(n7193), .B2(n7103), .A(n7102), .ZN(n7104) );
  OAI21_X1 U8816 ( .B1(n7195), .B2(n9585), .A(n7104), .ZN(P1_U3286) );
  NAND2_X1 U8817 ( .A1(n7108), .A2(n7107), .ZN(n7302) );
  NAND2_X1 U8818 ( .A1(n9170), .A2(n6541), .ZN(n7109) );
  OAI21_X1 U8819 ( .B1(n7260), .B2(n7883), .A(n7109), .ZN(n7110) );
  XNOR2_X1 U8820 ( .A(n7110), .B(n8292), .ZN(n7305) );
  OR2_X1 U8821 ( .A1(n7260), .A2(n7307), .ZN(n7112) );
  NAND2_X1 U8822 ( .A1(n9170), .A2(n7959), .ZN(n7111) );
  NAND2_X1 U8823 ( .A1(n7112), .A2(n7111), .ZN(n7303) );
  XNOR2_X1 U8824 ( .A(n7305), .B(n7303), .ZN(n7301) );
  XOR2_X1 U8825 ( .A(n7302), .B(n7301), .Z(n7120) );
  AOI22_X1 U8826 ( .A1(n9072), .A2(n9169), .B1(n7113), .B2(n9162), .ZN(n7119)
         );
  INV_X1 U8827 ( .A(n7114), .ZN(n7117) );
  NOR2_X1 U8828 ( .A1(n9157), .A2(n7115), .ZN(n7116) );
  AOI211_X1 U8829 ( .C1(n9077), .C2(n9171), .A(n7117), .B(n7116), .ZN(n7118)
         );
  OAI211_X1 U8830 ( .C1(n7120), .C2(n9164), .A(n7119), .B(n7118), .ZN(P1_U3213) );
  INV_X1 U8831 ( .A(n7121), .ZN(n7130) );
  INV_X1 U8832 ( .A(n9548), .ZN(n9492) );
  NAND2_X1 U8833 ( .A1(n9598), .A2(n9721), .ZN(n9561) );
  INV_X1 U8834 ( .A(n9561), .ZN(n7203) );
  AOI22_X1 U8835 ( .A1(n7203), .A2(n9175), .B1(n9587), .B2(n9173), .ZN(n7125)
         );
  OAI22_X1 U8836 ( .A1(n9598), .A2(n7122), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9557), .ZN(n7123) );
  AOI21_X1 U8837 ( .B1(n9569), .B2(n9016), .A(n7123), .ZN(n7124) );
  OAI211_X1 U8838 ( .C1(n9595), .C2(n7126), .A(n7125), .B(n7124), .ZN(n7127)
         );
  AOI21_X1 U8839 ( .B1(n7128), .B2(n9556), .A(n7127), .ZN(n7129) );
  OAI21_X1 U8840 ( .B1(n7130), .B2(n9492), .A(n7129), .ZN(P1_U3290) );
  XNOR2_X1 U8841 ( .A(n8496), .B(n4547), .ZN(n7132) );
  AOI21_X1 U8842 ( .B1(n5387), .B2(n7132), .A(n8497), .ZN(n7151) );
  INV_X1 U8843 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7133) );
  NOR2_X1 U8844 ( .A1(n9888), .A2(n7133), .ZN(n7139) );
  XNOR2_X1 U8845 ( .A(n8496), .B(n8469), .ZN(n7135) );
  AOI21_X1 U8846 ( .B1(n7135), .B2(n7188), .A(n8470), .ZN(n7137) );
  INV_X1 U8847 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10340) );
  NOR2_X1 U8848 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10340), .ZN(n7169) );
  INV_X1 U8849 ( .A(n7169), .ZN(n7136) );
  OAI21_X1 U8850 ( .B1(n9963), .B2(n7137), .A(n7136), .ZN(n7138) );
  NOR2_X1 U8851 ( .A1(n7139), .A2(n7138), .ZN(n7148) );
  MUX2_X1 U8852 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8561), .Z(n8484) );
  XNOR2_X1 U8853 ( .A(n8484), .B(n8496), .ZN(n7145) );
  OR2_X1 U8854 ( .A1(n7141), .A2(n7140), .ZN(n7143) );
  NAND2_X1 U8855 ( .A1(n7143), .A2(n7142), .ZN(n7144) );
  NAND2_X1 U8856 ( .A1(n7145), .A2(n7144), .ZN(n8485) );
  OAI21_X1 U8857 ( .B1(n7145), .B2(n7144), .A(n8485), .ZN(n7146) );
  NAND2_X1 U8858 ( .A1(n7146), .A2(n9967), .ZN(n7147) );
  OAI211_X1 U8859 ( .C1(n9977), .C2(n8483), .A(n7148), .B(n7147), .ZN(n7149)
         );
  INV_X1 U8860 ( .A(n7149), .ZN(n7150) );
  OAI21_X1 U8861 ( .B1(n7151), .B2(n9971), .A(n7150), .ZN(P2_U3193) );
  XOR2_X1 U8862 ( .A(n7684), .B(n7152), .Z(n7322) );
  INV_X1 U8863 ( .A(n7153), .ZN(n7155) );
  INV_X1 U8864 ( .A(n7684), .ZN(n7154) );
  NAND2_X1 U8865 ( .A1(n7155), .A2(n7154), .ZN(n7156) );
  AND2_X1 U8866 ( .A1(n7157), .A2(n7156), .ZN(n7330) );
  NAND2_X1 U8867 ( .A1(n7688), .A2(n8745), .ZN(n7161) );
  OAI22_X1 U8868 ( .A1(n8728), .A2(n7158), .B1(n7292), .B2(n8788), .ZN(n7159)
         );
  AOI21_X1 U8869 ( .B1(n8795), .B2(n8763), .A(n7159), .ZN(n7160) );
  OAI211_X1 U8870 ( .C1(n7321), .C2(n8712), .A(n7161), .B(n7160), .ZN(n7162)
         );
  AOI21_X1 U8871 ( .B1(n7330), .B2(n8793), .A(n7162), .ZN(n7163) );
  OAI21_X1 U8872 ( .B1(n7322), .B2(n8720), .A(n7163), .ZN(P2_U3221) );
  INV_X1 U8873 ( .A(n7190), .ZN(n10063) );
  NAND2_X1 U8874 ( .A1(n7167), .A2(n7166), .ZN(n7603) );
  XNOR2_X1 U8875 ( .A(n7603), .B(n8051), .ZN(n7287) );
  OAI211_X1 U8876 ( .C1(n7168), .C2(n7287), .A(n7286), .B(n8423), .ZN(n7174)
         );
  INV_X1 U8877 ( .A(n7187), .ZN(n7172) );
  AOI21_X1 U8878 ( .B1(n8431), .B2(n10041), .A(n7169), .ZN(n7170) );
  OAI21_X1 U8879 ( .B1(n8392), .B2(n8427), .A(n7170), .ZN(n7171) );
  AOI21_X1 U8880 ( .B1(n7172), .B2(n8415), .A(n7171), .ZN(n7173) );
  OAI211_X1 U8881 ( .C1(n10063), .C2(n8434), .A(n7174), .B(n7173), .ZN(
        P2_U3176) );
  AOI22_X1 U8882 ( .A1(n7203), .A2(n9177), .B1(n9587), .B2(n9174), .ZN(n7176)
         );
  INV_X1 U8883 ( .A(n9557), .ZN(n9583) );
  AOI22_X1 U8884 ( .A1(n9585), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9583), .ZN(n7175) );
  OAI211_X1 U8885 ( .C1(n8077), .C2(n9590), .A(n7176), .B(n7175), .ZN(n7177)
         );
  AOI21_X1 U8886 ( .B1(n9538), .B2(n7178), .A(n7177), .ZN(n7181) );
  NAND2_X1 U8887 ( .A1(n7179), .A2(n9556), .ZN(n7180) );
  OAI211_X1 U8888 ( .C1(n7182), .C2(n9492), .A(n7181), .B(n7180), .ZN(P1_U3291) );
  XOR2_X1 U8889 ( .A(n7603), .B(n7183), .Z(n10065) );
  XNOR2_X1 U8890 ( .A(n7184), .B(n7603), .ZN(n7185) );
  OAI222_X1 U8891 ( .A1(n10025), .A2(n8392), .B1(n10027), .B2(n7186), .C1(
        n7185), .C2(n9979), .ZN(n10067) );
  NAND2_X1 U8892 ( .A1(n10067), .A2(n8728), .ZN(n7192) );
  OAI22_X1 U8893 ( .A1(n8728), .A2(n7188), .B1(n7187), .B2(n8788), .ZN(n7189)
         );
  AOI21_X1 U8894 ( .B1(n7190), .B2(n8745), .A(n7189), .ZN(n7191) );
  OAI211_X1 U8895 ( .C1(n10065), .C2(n8784), .A(n7192), .B(n7191), .ZN(
        P2_U3222) );
  INV_X1 U8896 ( .A(n7193), .ZN(n7196) );
  OAI211_X1 U8897 ( .C1(n7196), .C2(n9737), .A(n7195), .B(n7194), .ZN(n7201)
         );
  INV_X1 U8898 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7197) );
  OAI22_X1 U8899 ( .A1(n9742), .A2(n7260), .B1(n9850), .B2(n7197), .ZN(n7198)
         );
  AOI21_X1 U8900 ( .B1(n7201), .B2(n9850), .A(n7198), .ZN(n7199) );
  INV_X1 U8901 ( .A(n7199), .ZN(P1_U3529) );
  OAI22_X1 U8902 ( .A1(n9783), .A2(n7260), .B1(n9838), .B2(n6866), .ZN(n7200)
         );
  AOI21_X1 U8903 ( .B1(n7201), .B2(n9838), .A(n7200), .ZN(n7202) );
  INV_X1 U8904 ( .A(n7202), .ZN(P1_U3474) );
  AOI22_X1 U8905 ( .A1(n7203), .A2(n9178), .B1(n9587), .B2(n9175), .ZN(n7208)
         );
  OAI22_X1 U8906 ( .A1(n9598), .A2(n4739), .B1(n7204), .B2(n9557), .ZN(n7205)
         );
  AOI21_X1 U8907 ( .B1(n9569), .B2(n7206), .A(n7205), .ZN(n7207) );
  OAI211_X1 U8908 ( .C1(n9595), .C2(n7209), .A(n7208), .B(n7207), .ZN(n7212)
         );
  NOR2_X1 U8909 ( .A1(n7210), .A2(n9600), .ZN(n7211) );
  AOI211_X1 U8910 ( .C1(n7213), .C2(n9598), .A(n7212), .B(n7211), .ZN(n7214)
         );
  INV_X1 U8911 ( .A(n7214), .ZN(P1_U3292) );
  INV_X1 U8912 ( .A(n7501), .ZN(n7285) );
  OAI222_X1 U8913 ( .A1(n8990), .A2(n7285), .B1(P2_U3151), .B2(n7618), .C1(
        n7215), .C2(n8991), .ZN(P2_U3274) );
  INV_X1 U8914 ( .A(n7216), .ZN(n7226) );
  OAI22_X1 U8915 ( .A1(n9598), .A2(n7217), .B1(n9074), .B2(n9557), .ZN(n7220)
         );
  NOR2_X1 U8916 ( .A1(n9561), .A2(n7218), .ZN(n7219) );
  AOI211_X1 U8917 ( .C1(n9569), .C2(n9071), .A(n7220), .B(n7219), .ZN(n7221)
         );
  OAI21_X1 U8918 ( .B1(n7222), .B2(n9595), .A(n7221), .ZN(n7223) );
  AOI21_X1 U8919 ( .B1(n7224), .B2(n9556), .A(n7223), .ZN(n7225) );
  OAI21_X1 U8920 ( .B1(n7226), .B2(n9585), .A(n7225), .ZN(P1_U3288) );
  NAND2_X1 U8921 ( .A1(n7227), .A2(n8123), .ZN(n7233) );
  NAND2_X1 U8922 ( .A1(n7228), .A2(n7533), .ZN(n7232) );
  AOI22_X1 U8923 ( .A1(n7526), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7525), .B2(
        n7230), .ZN(n7231) );
  NAND2_X1 U8924 ( .A1(n7232), .A2(n7231), .ZN(n9817) );
  OR2_X1 U8925 ( .A1(n9817), .A2(n7428), .ZN(n8140) );
  NAND2_X1 U8926 ( .A1(n9817), .A2(n7428), .ZN(n8218) );
  NAND2_X1 U8927 ( .A1(n8140), .A2(n8218), .ZN(n7237) );
  XNOR2_X1 U8928 ( .A(n7233), .B(n7237), .ZN(n7234) );
  AOI22_X1 U8929 ( .A1(n7234), .A2(n9713), .B1(n9721), .B2(n9169), .ZN(n9819)
         );
  OAI21_X1 U8930 ( .B1(n7238), .B2(n7237), .A(n7275), .ZN(n9821) );
  XOR2_X1 U8931 ( .A(n9817), .B(n7279), .Z(n7247) );
  NAND2_X1 U8932 ( .A1(n7989), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7246) );
  INV_X1 U8933 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7239) );
  OR2_X1 U8934 ( .A1(n7992), .A2(n7239), .ZN(n7245) );
  NAND2_X1 U8935 ( .A1(n7241), .A2(n7240), .ZN(n7242) );
  NAND2_X1 U8936 ( .A1(n7266), .A2(n7242), .ZN(n7426) );
  OR2_X1 U8937 ( .A1(n7988), .A2(n7426), .ZN(n7244) );
  INV_X1 U8938 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7278) );
  OR2_X1 U8939 ( .A1(n7907), .A2(n7278), .ZN(n7243) );
  INV_X1 U8940 ( .A(n7446), .ZN(n9167) );
  AOI22_X1 U8941 ( .A1(n7247), .A2(n9593), .B1(n9720), .B2(n9167), .ZN(n9818)
         );
  OAI22_X1 U8942 ( .A1(n9598), .A2(n6203), .B1(n7398), .B2(n9557), .ZN(n7248)
         );
  AOI21_X1 U8943 ( .B1(n9569), .B2(n9817), .A(n7248), .ZN(n7249) );
  OAI21_X1 U8944 ( .B1(n9818), .B2(n9595), .A(n7249), .ZN(n7250) );
  AOI21_X1 U8945 ( .B1(n9821), .B2(n9556), .A(n7250), .ZN(n7251) );
  OAI21_X1 U8946 ( .B1(n9585), .B2(n9819), .A(n7251), .ZN(P1_U3284) );
  OR2_X1 U8947 ( .A1(n7252), .A2(n7504), .ZN(n7255) );
  AOI22_X1 U8948 ( .A1(n7526), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7525), .B2(
        n7253), .ZN(n7254) );
  OR2_X1 U8949 ( .A1(n7422), .A2(n7446), .ZN(n8139) );
  NAND2_X1 U8950 ( .A1(n7422), .A2(n7446), .ZN(n8087) );
  NAND2_X1 U8951 ( .A1(n8139), .A2(n8087), .ZN(n7276) );
  INV_X1 U8952 ( .A(n7276), .ZN(n8219) );
  INV_X1 U8953 ( .A(n8218), .ZN(n7257) );
  NAND2_X1 U8954 ( .A1(n8121), .A2(n7256), .ZN(n8214) );
  OR3_X1 U8955 ( .A1(n8086), .A2(n7257), .A3(n8214), .ZN(n7262) );
  NAND2_X1 U8956 ( .A1(n8214), .A2(n8123), .ZN(n7258) );
  NAND2_X1 U8957 ( .A1(n7258), .A2(n8218), .ZN(n7259) );
  NAND2_X1 U8958 ( .A1(n7259), .A2(n8140), .ZN(n8081) );
  NAND2_X1 U8959 ( .A1(n7260), .A2(n9170), .ZN(n7261) );
  AND2_X1 U8960 ( .A1(n8123), .A2(n7261), .ZN(n8118) );
  NAND3_X1 U8961 ( .A1(n8118), .A2(n8140), .A3(n8112), .ZN(n8217) );
  NAND2_X1 U8962 ( .A1(n8081), .A2(n8217), .ZN(n8084) );
  OAI21_X1 U8963 ( .B1(n8219), .B2(n7263), .A(n7364), .ZN(n7273) );
  NAND2_X1 U8964 ( .A1(n7989), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7271) );
  OR2_X1 U8965 ( .A1(n7992), .A2(n7264), .ZN(n7270) );
  INV_X1 U8966 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7356) );
  OR2_X1 U8967 ( .A1(n7907), .A2(n7356), .ZN(n7269) );
  INV_X1 U8968 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7265) );
  NAND2_X1 U8969 ( .A1(n7266), .A2(n7265), .ZN(n7267) );
  NAND2_X1 U8970 ( .A1(n7346), .A2(n7267), .ZN(n7445) );
  OR2_X1 U8971 ( .A1(n7988), .A2(n7445), .ZN(n7268) );
  OAI22_X1 U8972 ( .A1(n7428), .A2(n9708), .B1(n9046), .B2(n9731), .ZN(n7272)
         );
  AOI21_X1 U8973 ( .B1(n7273), .B2(n9713), .A(n7272), .ZN(n9824) );
  NAND2_X1 U8974 ( .A1(n7277), .A2(n7276), .ZN(n7338) );
  OAI21_X1 U8975 ( .B1(n7277), .B2(n7276), .A(n7338), .ZN(n9827) );
  NAND2_X1 U8976 ( .A1(n9827), .A2(n9556), .ZN(n7284) );
  OAI22_X1 U8977 ( .A1(n9598), .A2(n7278), .B1(n7426), .B2(n9557), .ZN(n7282)
         );
  OAI21_X1 U8978 ( .B1(n7279), .B2(n9817), .A(n7422), .ZN(n7280) );
  NAND3_X1 U8979 ( .A1(n4709), .A2(n9593), .A3(n7280), .ZN(n9823) );
  NOR2_X1 U8980 ( .A1(n9823), .A2(n9595), .ZN(n7281) );
  AOI211_X1 U8981 ( .C1(n9569), .C2(n7422), .A(n7282), .B(n7281), .ZN(n7283)
         );
  OAI211_X1 U8982 ( .C1(n9585), .C2(n9824), .A(n7284), .B(n7283), .ZN(P1_U3283) );
  OAI222_X1 U8983 ( .A1(n6832), .A2(n10416), .B1(n7300), .B2(n7285), .C1(
        P1_U3086), .C2(n8267), .ZN(P1_U3334) );
  XNOR2_X1 U8984 ( .A(n7688), .B(n8051), .ZN(n8018) );
  XOR2_X1 U8985 ( .A(n8775), .B(n8018), .Z(n7289) );
  AOI21_X1 U8986 ( .B1(n7289), .B2(n7288), .A(n4585), .ZN(n7295) );
  OAI22_X1 U8987 ( .A1(n8409), .A2(n7321), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10476), .ZN(n7290) );
  AOI21_X1 U8988 ( .B1(n8406), .B2(n8763), .A(n7290), .ZN(n7291) );
  OAI21_X1 U8989 ( .B1(n7292), .B2(n8428), .A(n7291), .ZN(n7293) );
  AOI21_X1 U8990 ( .B1(n7688), .B2(n8419), .A(n7293), .ZN(n7294) );
  OAI21_X1 U8991 ( .B1(n7295), .B2(n8421), .A(n7294), .ZN(P2_U3164) );
  INV_X1 U8992 ( .A(n7497), .ZN(n7299) );
  OAI222_X1 U8993 ( .A1(n8991), .A2(n7297), .B1(n8990), .B2(n7299), .C1(n7296), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U8994 ( .A1(n6832), .A2(n7498), .B1(n7300), .B2(n7299), .C1(n7298), 
        .C2(P1_U3086), .ZN(P1_U3333) );
  INV_X1 U8995 ( .A(n7303), .ZN(n7304) );
  NAND2_X1 U8996 ( .A1(n7305), .A2(n7304), .ZN(n7306) );
  NAND2_X1 U8997 ( .A1(n9169), .A2(n6541), .ZN(n7308) );
  OAI21_X1 U8998 ( .B1(n9811), .B2(n7883), .A(n7308), .ZN(n7309) );
  XNOR2_X1 U8999 ( .A(n7309), .B(n7998), .ZN(n7412) );
  INV_X1 U9000 ( .A(n7412), .ZN(n7409) );
  XNOR2_X1 U9001 ( .A(n7404), .B(n7409), .ZN(n7312) );
  OR2_X1 U9002 ( .A1(n9811), .A2(n7307), .ZN(n7311) );
  NAND2_X1 U9003 ( .A1(n9169), .A2(n7959), .ZN(n7310) );
  NAND2_X1 U9004 ( .A1(n7311), .A2(n7310), .ZN(n7410) );
  NOR2_X1 U9005 ( .A1(n7312), .A2(n7410), .ZN(n7389) );
  AOI21_X1 U9006 ( .B1(n7312), .B2(n7410), .A(n7389), .ZN(n7320) );
  OAI21_X1 U9007 ( .B1(n9157), .B2(n7314), .A(n7313), .ZN(n7317) );
  INV_X1 U9008 ( .A(n9170), .ZN(n7315) );
  OAI22_X1 U9009 ( .A1(n7315), .A2(n9159), .B1(n9158), .B2(n7428), .ZN(n7316)
         );
  AOI211_X1 U9010 ( .C1(n7318), .C2(n9162), .A(n7317), .B(n7316), .ZN(n7319)
         );
  OAI21_X1 U9011 ( .B1(n7320), .B2(n9164), .A(n7319), .ZN(P1_U3221) );
  OAI22_X1 U9012 ( .A1(n7321), .A2(n10027), .B1(n8021), .B2(n10025), .ZN(n7324) );
  NOR2_X1 U9013 ( .A1(n7322), .A2(n9979), .ZN(n7323) );
  AOI211_X1 U9014 ( .C1(n10060), .C2(n7688), .A(n7324), .B(n7323), .ZN(n7332)
         );
  INV_X1 U9015 ( .A(n8893), .ZN(n7327) );
  NOR2_X1 U9016 ( .A1(n10087), .A2(n7325), .ZN(n7326) );
  AOI21_X1 U9017 ( .B1(n7330), .B2(n7327), .A(n7326), .ZN(n7328) );
  OAI21_X1 U9018 ( .B1(n7332), .B2(n10085), .A(n7328), .ZN(P2_U3471) );
  INV_X1 U9019 ( .A(n8974), .ZN(n7329) );
  AOI22_X1 U9020 ( .A1(n7330), .A2(n7329), .B1(P2_REG0_REG_12__SCAN_IN), .B2(
        n10070), .ZN(n7331) );
  OAI21_X1 U9021 ( .B1(n7332), .B2(n10070), .A(n7331), .ZN(P2_U3426) );
  NAND2_X1 U9022 ( .A1(n7493), .A2(n8981), .ZN(n7334) );
  NAND2_X1 U9023 ( .A1(n7333), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7791) );
  OAI211_X1 U9024 ( .C1(n7335), .C2(n8991), .A(n7334), .B(n7791), .ZN(P2_U3272) );
  NAND2_X1 U9025 ( .A1(n7493), .A2(n9790), .ZN(n7336) );
  OAI211_X1 U9026 ( .C1(n7494), .C2(n6832), .A(n7336), .B(n8285), .ZN(P1_U3332) );
  NAND2_X1 U9027 ( .A1(n7338), .A2(n7337), .ZN(n7343) );
  NAND2_X1 U9028 ( .A1(n7339), .A2(n7533), .ZN(n7342) );
  AOI22_X1 U9029 ( .A1(n7526), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7525), .B2(
        n7340), .ZN(n7341) );
  OR2_X1 U9030 ( .A1(n7449), .A2(n9046), .ZN(n8127) );
  NAND2_X1 U9031 ( .A1(n7449), .A2(n9046), .ZN(n8128) );
  NAND2_X1 U9032 ( .A1(n8127), .A2(n8128), .ZN(n8223) );
  OAI21_X1 U9033 ( .B1(n7343), .B2(n8223), .A(n7381), .ZN(n9740) );
  INV_X1 U9034 ( .A(n9740), .ZN(n7362) );
  NAND2_X1 U9035 ( .A1(n7364), .A2(n8087), .ZN(n7344) );
  XOR2_X1 U9036 ( .A(n8223), .B(n7344), .Z(n7353) );
  NAND2_X1 U9037 ( .A1(n7989), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7351) );
  OR2_X1 U9038 ( .A1(n7992), .A2(n9848), .ZN(n7350) );
  NAND2_X1 U9039 ( .A1(n7346), .A2(n7345), .ZN(n7347) );
  NAND2_X1 U9040 ( .A1(n7371), .A2(n7347), .ZN(n9045) );
  OR2_X1 U9041 ( .A1(n7988), .A2(n9045), .ZN(n7349) );
  INV_X1 U9042 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7383) );
  OR2_X1 U9043 ( .A1(n7981), .A2(n7383), .ZN(n7348) );
  OAI22_X1 U9044 ( .A1(n7446), .A2(n9708), .B1(n9580), .B2(n9731), .ZN(n7352)
         );
  AOI21_X1 U9045 ( .B1(n7353), .B2(n9713), .A(n7352), .ZN(n7354) );
  OAI21_X1 U9046 ( .B1(n7362), .B2(n7355), .A(n7354), .ZN(n9738) );
  NAND2_X1 U9047 ( .A1(n9738), .A2(n9598), .ZN(n7360) );
  AOI211_X1 U9048 ( .C1(n7449), .C2(n4709), .A(n9494), .B(n7384), .ZN(n9739)
         );
  NOR2_X1 U9049 ( .A1(n9784), .A2(n9590), .ZN(n7358) );
  OAI22_X1 U9050 ( .A1(n9598), .A2(n7356), .B1(n7445), .B2(n9557), .ZN(n7357)
         );
  AOI211_X1 U9051 ( .C1(n9739), .C2(n9538), .A(n7358), .B(n7357), .ZN(n7359)
         );
  OAI211_X1 U9052 ( .C1(n7362), .C2(n7361), .A(n7360), .B(n7359), .ZN(P1_U3282) );
  INV_X1 U9053 ( .A(n8087), .ZN(n8126) );
  NOR2_X1 U9054 ( .A1(n8223), .A2(n8126), .ZN(n7363) );
  OR2_X1 U9055 ( .A1(n7365), .A2(n7504), .ZN(n7368) );
  AOI22_X1 U9056 ( .A1(n7526), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7525), .B2(
        n7366), .ZN(n7367) );
  NAND2_X1 U9057 ( .A1(n7368), .A2(n7367), .ZN(n9270) );
  OR2_X1 U9058 ( .A1(n9270), .A2(n9580), .ZN(n8132) );
  NAND2_X1 U9059 ( .A1(n9270), .A2(n9580), .ZN(n9574) );
  NAND2_X1 U9060 ( .A1(n8132), .A2(n9574), .ZN(n8236) );
  XNOR2_X1 U9061 ( .A(n8237), .B(n8236), .ZN(n7379) );
  NAND2_X1 U9062 ( .A1(n4513), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7377) );
  INV_X1 U9063 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7369) );
  OR2_X1 U9064 ( .A1(n7907), .A2(n7369), .ZN(n7376) );
  NAND2_X1 U9065 ( .A1(n7371), .A2(n7370), .ZN(n7372) );
  NAND2_X1 U9066 ( .A1(n7834), .A2(n7372), .ZN(n9119) );
  OR2_X1 U9067 ( .A1(n7988), .A2(n9119), .ZN(n7375) );
  INV_X1 U9068 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7373) );
  OR2_X1 U9069 ( .A1(n4602), .A2(n7373), .ZN(n7374) );
  OAI22_X1 U9070 ( .A1(n9046), .A2(n9708), .B1(n9562), .B2(n9731), .ZN(n7378)
         );
  AOI21_X1 U9071 ( .B1(n7379), .B2(n9713), .A(n7378), .ZN(n9830) );
  INV_X1 U9072 ( .A(n9046), .ZN(n9166) );
  OAI21_X1 U9073 ( .B1(n7382), .B2(n8236), .A(n9271), .ZN(n9835) );
  NAND2_X1 U9074 ( .A1(n9835), .A2(n9556), .ZN(n7388) );
  OAI22_X1 U9075 ( .A1(n9598), .A2(n7383), .B1(n9045), .B2(n9557), .ZN(n7386)
         );
  INV_X1 U9076 ( .A(n9270), .ZN(n9832) );
  NAND2_X1 U9077 ( .A1(n7384), .A2(n9832), .ZN(n9591) );
  OAI211_X1 U9078 ( .C1(n7384), .C2(n9832), .A(n9593), .B(n9591), .ZN(n9829)
         );
  NOR2_X1 U9079 ( .A1(n9829), .A2(n9595), .ZN(n7385) );
  AOI211_X1 U9080 ( .C1(n9569), .C2(n9270), .A(n7386), .B(n7385), .ZN(n7387)
         );
  OAI211_X1 U9081 ( .C1(n9585), .C2(n9830), .A(n7388), .B(n7387), .ZN(P1_U3281) );
  AOI21_X1 U9082 ( .B1(n7409), .B2(n7404), .A(n7389), .ZN(n7396) );
  NAND2_X1 U9083 ( .A1(n9817), .A2(n8289), .ZN(n7391) );
  OR2_X1 U9084 ( .A1(n7428), .A2(n7307), .ZN(n7390) );
  NAND2_X1 U9085 ( .A1(n7391), .A2(n7390), .ZN(n7392) );
  XNOR2_X1 U9086 ( .A(n7392), .B(n7998), .ZN(n7414) );
  NAND2_X1 U9087 ( .A1(n9817), .A2(n6541), .ZN(n7394) );
  OR2_X1 U9088 ( .A1(n7428), .A2(n8295), .ZN(n7393) );
  NAND2_X1 U9089 ( .A1(n7394), .A2(n7393), .ZN(n7411) );
  INV_X1 U9090 ( .A(n7411), .ZN(n7407) );
  XNOR2_X1 U9091 ( .A(n7414), .B(n7407), .ZN(n7395) );
  XNOR2_X1 U9092 ( .A(n7396), .B(n7395), .ZN(n7403) );
  OAI21_X1 U9093 ( .B1(n9157), .B2(n7398), .A(n7397), .ZN(n7401) );
  OAI22_X1 U9094 ( .A1(n7399), .A2(n9159), .B1(n9158), .B2(n7446), .ZN(n7400)
         );
  AOI211_X1 U9095 ( .C1(n9817), .C2(n9162), .A(n7401), .B(n7400), .ZN(n7402)
         );
  OAI21_X1 U9096 ( .B1(n7403), .B2(n9164), .A(n7402), .ZN(P1_U3231) );
  INV_X1 U9097 ( .A(n7422), .ZN(n9825) );
  OAI22_X1 U9098 ( .A1(n7414), .A2(n7411), .B1(n7412), .B2(n7410), .ZN(n7405)
         );
  INV_X1 U9099 ( .A(n7405), .ZN(n7406) );
  INV_X1 U9100 ( .A(n7410), .ZN(n7408) );
  OAI21_X1 U9101 ( .B1(n7409), .B2(n7408), .A(n7407), .ZN(n7415) );
  AND2_X1 U9102 ( .A1(n7411), .A2(n7410), .ZN(n7413) );
  AOI22_X1 U9103 ( .A1(n7415), .A2(n7414), .B1(n7413), .B2(n7412), .ZN(n7416)
         );
  NAND2_X1 U9104 ( .A1(n7422), .A2(n8289), .ZN(n7419) );
  OR2_X1 U9105 ( .A1(n7446), .A2(n7307), .ZN(n7418) );
  NAND2_X1 U9106 ( .A1(n7419), .A2(n7418), .ZN(n7420) );
  XNOR2_X1 U9107 ( .A(n7420), .B(n8292), .ZN(n7435) );
  XNOR2_X1 U9108 ( .A(n7434), .B(n7435), .ZN(n7424) );
  NOR2_X1 U9109 ( .A1(n7446), .A2(n8295), .ZN(n7421) );
  AOI21_X1 U9110 ( .B1(n7422), .B2(n6541), .A(n7421), .ZN(n7423) );
  NAND2_X1 U9111 ( .A1(n7424), .A2(n7423), .ZN(n7438) );
  OAI21_X1 U9112 ( .B1(n7424), .B2(n7423), .A(n7438), .ZN(n7425) );
  NAND2_X1 U9113 ( .A1(n7425), .A2(n9143), .ZN(n7433) );
  INV_X1 U9114 ( .A(n7426), .ZN(n7431) );
  INV_X1 U9115 ( .A(n9157), .ZN(n9123) );
  INV_X1 U9116 ( .A(n7427), .ZN(n7430) );
  OAI22_X1 U9117 ( .A1(n7428), .A2(n9159), .B1(n9158), .B2(n9046), .ZN(n7429)
         );
  AOI211_X1 U9118 ( .C1(n7431), .C2(n9123), .A(n7430), .B(n7429), .ZN(n7432)
         );
  OAI211_X1 U9119 ( .C1(n9825), .C2(n9126), .A(n7433), .B(n7432), .ZN(P1_U3217) );
  INV_X1 U9120 ( .A(n7434), .ZN(n7436) );
  NAND2_X1 U9121 ( .A1(n7436), .A2(n7435), .ZN(n7437) );
  NAND2_X1 U9122 ( .A1(n7449), .A2(n8289), .ZN(n7440) );
  OR2_X1 U9123 ( .A1(n9046), .A2(n7307), .ZN(n7439) );
  NAND2_X1 U9124 ( .A1(n7440), .A2(n7439), .ZN(n7441) );
  XNOR2_X1 U9125 ( .A(n7441), .B(n8292), .ZN(n7811) );
  NOR2_X1 U9126 ( .A1(n9046), .A2(n8295), .ZN(n7442) );
  AOI21_X1 U9127 ( .B1(n7449), .B2(n6541), .A(n7442), .ZN(n7812) );
  XNOR2_X1 U9128 ( .A(n7811), .B(n7812), .ZN(n7443) );
  XNOR2_X1 U9129 ( .A(n7810), .B(n7443), .ZN(n7451) );
  OAI21_X1 U9130 ( .B1(n9157), .B2(n7445), .A(n7444), .ZN(n7448) );
  OAI22_X1 U9131 ( .A1(n7446), .A2(n9159), .B1(n9158), .B2(n9580), .ZN(n7447)
         );
  AOI211_X1 U9132 ( .C1(n7449), .C2(n9162), .A(n7448), .B(n7447), .ZN(n7450)
         );
  OAI21_X1 U9133 ( .B1(n7451), .B2(n9164), .A(n7450), .ZN(P1_U3236) );
  INV_X1 U9134 ( .A(n7490), .ZN(n7561) );
  OAI222_X1 U9135 ( .A1(n6832), .A2(n7491), .B1(n7300), .B2(n7561), .C1(
        P1_U3086), .C2(n7452), .ZN(P1_U3331) );
  INV_X1 U9136 ( .A(n7453), .ZN(n7454) );
  NAND2_X1 U9137 ( .A1(n7454), .A2(SI_29_), .ZN(n7460) );
  INV_X1 U9138 ( .A(n7455), .ZN(n7458) );
  INV_X1 U9139 ( .A(n7456), .ZN(n7457) );
  NAND2_X1 U9140 ( .A1(n7458), .A2(n7457), .ZN(n7459) );
  NAND2_X1 U9141 ( .A1(n7460), .A2(n7459), .ZN(n7476) );
  INV_X1 U9142 ( .A(n7476), .ZN(n7466) );
  INV_X1 U9143 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10448) );
  MUX2_X1 U9144 ( .A(n10448), .B(n7552), .S(n7468), .Z(n7462) );
  INV_X1 U9145 ( .A(SI_30_), .ZN(n7461) );
  NAND2_X1 U9146 ( .A1(n7462), .A2(n7461), .ZN(n7467) );
  INV_X1 U9147 ( .A(n7462), .ZN(n7463) );
  NAND2_X1 U9148 ( .A1(n7463), .A2(SI_30_), .ZN(n7464) );
  NAND2_X1 U9149 ( .A1(n7467), .A2(n7464), .ZN(n7475) );
  INV_X1 U9150 ( .A(n7475), .ZN(n7465) );
  NAND2_X1 U9151 ( .A1(n7466), .A2(n7465), .ZN(n7478) );
  NAND2_X1 U9152 ( .A1(n7478), .A2(n7467), .ZN(n7472) );
  MUX2_X1 U9153 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7468), .Z(n7470) );
  INV_X1 U9154 ( .A(SI_31_), .ZN(n7469) );
  XNOR2_X1 U9155 ( .A(n7470), .B(n7469), .ZN(n7471) );
  NAND2_X1 U9156 ( .A1(n8976), .A2(n4514), .ZN(n7474) );
  OR2_X1 U9157 ( .A1(n7534), .A2(n10446), .ZN(n7473) );
  NAND2_X1 U9158 ( .A1(n7476), .A2(n7475), .ZN(n7477) );
  NAND2_X1 U9159 ( .A1(n7478), .A2(n7477), .ZN(n7580) );
  NAND2_X1 U9160 ( .A1(n7580), .A2(n7533), .ZN(n7480) );
  OR2_X1 U9161 ( .A1(n7534), .A2(n10448), .ZN(n7479) );
  NAND2_X1 U9162 ( .A1(n7549), .A2(n4514), .ZN(n7483) );
  OR2_X1 U9163 ( .A1(n7534), .A2(n7481), .ZN(n7482) );
  NAND2_X1 U9164 ( .A1(n8308), .A2(n4514), .ZN(n7485) );
  INV_X1 U9165 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10285) );
  OR2_X1 U9166 ( .A1(n7534), .A2(n10285), .ZN(n7484) );
  NAND2_X1 U9167 ( .A1(n7557), .A2(n7533), .ZN(n7487) );
  OR2_X1 U9168 ( .A1(n7534), .A2(n7559), .ZN(n7486) );
  NAND2_X1 U9169 ( .A1(n7555), .A2(n4514), .ZN(n7489) );
  OR2_X1 U9170 ( .A1(n7534), .A2(n10489), .ZN(n7488) );
  OR2_X1 U9171 ( .A1(n7534), .A2(n7491), .ZN(n7492) );
  NAND2_X1 U9172 ( .A1(n7493), .A2(n4514), .ZN(n7496) );
  OR2_X1 U9173 ( .A1(n7534), .A2(n7494), .ZN(n7495) );
  NAND2_X1 U9174 ( .A1(n7497), .A2(n7533), .ZN(n7500) );
  OR2_X1 U9175 ( .A1(n7534), .A2(n7498), .ZN(n7499) );
  NAND2_X1 U9176 ( .A1(n7501), .A2(n7533), .ZN(n7503) );
  OR2_X1 U9177 ( .A1(n7534), .A2(n10416), .ZN(n7502) );
  OR2_X1 U9178 ( .A1(n7505), .A2(n7504), .ZN(n7508) );
  AOI22_X1 U9179 ( .A1(n7526), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7525), .B2(
        n7506), .ZN(n7507) );
  OR2_X1 U9180 ( .A1(n9591), .A2(n9272), .ZN(n9592) );
  NAND2_X1 U9181 ( .A1(n7509), .A2(n7533), .ZN(n7511) );
  AOI22_X1 U9182 ( .A1(n7526), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7525), .B2(
        n9187), .ZN(n7510) );
  NAND2_X1 U9183 ( .A1(n7512), .A2(n7533), .ZN(n7514) );
  INV_X1 U9184 ( .A(n9201), .ZN(n9182) );
  AOI22_X1 U9185 ( .A1(n7526), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7525), .B2(
        n9182), .ZN(n7513) );
  INV_X1 U9186 ( .A(n9711), .ZN(n9546) );
  NAND2_X1 U9187 ( .A1(n7515), .A2(n7533), .ZN(n7517) );
  AOI22_X1 U9188 ( .A1(n7526), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7525), .B2(
        n9217), .ZN(n7516) );
  NAND2_X1 U9189 ( .A1(n7518), .A2(n7533), .ZN(n7520) );
  AOI22_X1 U9190 ( .A1(n7526), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7525), .B2(
        n9215), .ZN(n7519) );
  NAND2_X1 U9191 ( .A1(n7521), .A2(n4514), .ZN(n7523) );
  AOI22_X1 U9192 ( .A1(n7526), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7525), .B2(
        n9241), .ZN(n7522) );
  NAND2_X1 U9193 ( .A1(n7524), .A2(n4514), .ZN(n7528) );
  AOI22_X1 U9194 ( .A1(n7526), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9327), .B2(
        n7525), .ZN(n7527) );
  NAND2_X1 U9195 ( .A1(n7529), .A2(n4514), .ZN(n7532) );
  INV_X1 U9196 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7530) );
  OR2_X1 U9197 ( .A1(n7534), .A2(n7530), .ZN(n7531) );
  NAND2_X1 U9198 ( .A1(n9468), .A2(n9448), .ZN(n9445) );
  NAND2_X1 U9199 ( .A1(n9661), .A2(n9434), .ZN(n9417) );
  NOR2_X4 U9200 ( .A1(n9390), .A2(n9401), .ZN(n9389) );
  OR2_X1 U9201 ( .A1(n7534), .A2(n10190), .ZN(n7535) );
  NOR2_X2 U9202 ( .A1(n8101), .A2(n9326), .ZN(n9293) );
  NAND2_X1 U9203 ( .A1(n9746), .A2(n9293), .ZN(n9262) );
  XNOR2_X1 U9204 ( .A(n8105), .B(n9262), .ZN(n7537) );
  INV_X1 U9205 ( .A(n9793), .ZN(n7538) );
  AND2_X1 U9206 ( .A1(n7538), .A2(P1_B_REG_SCAN_IN), .ZN(n7539) );
  NOR2_X1 U9207 ( .A1(n8252), .A2(n9310), .ZN(n9602) );
  NOR2_X1 U9208 ( .A1(n7545), .A2(n9602), .ZN(n7542) );
  MUX2_X1 U9209 ( .A(n7540), .B(n7542), .S(n9838), .Z(n7541) );
  OAI21_X1 U9210 ( .B1(n8188), .B2(n9783), .A(n7541), .ZN(P1_U3521) );
  INV_X1 U9211 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n7543) );
  MUX2_X1 U9212 ( .A(n7543), .B(n7542), .S(n9850), .Z(n7544) );
  OAI21_X1 U9213 ( .B1(n8188), .B2(n9742), .A(n7544), .ZN(P1_U3553) );
  NAND2_X1 U9214 ( .A1(n7545), .A2(n9538), .ZN(n7548) );
  INV_X1 U9215 ( .A(n9602), .ZN(n7546) );
  NOR2_X1 U9216 ( .A1(n9585), .A2(n7546), .ZN(n9266) );
  AOI21_X1 U9217 ( .B1(n9585), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9266), .ZN(
        n7547) );
  OAI211_X1 U9218 ( .C1(n8188), .C2(n9590), .A(n7548), .B(n7547), .ZN(P1_U3263) );
  INV_X1 U9219 ( .A(n7549), .ZN(n8288) );
  OAI222_X1 U9220 ( .A1(n7300), .A2(n8288), .B1(n6832), .B2(n7481), .C1(
        P1_U3086), .C2(n7550), .ZN(P1_U3326) );
  INV_X1 U9221 ( .A(n7580), .ZN(n7553) );
  OAI222_X1 U9222 ( .A1(n6832), .A2(n10448), .B1(n7300), .B2(n7553), .C1(
        P1_U3086), .C2(n7551), .ZN(P1_U3325) );
  OAI222_X1 U9223 ( .A1(n7554), .A2(P2_U3151), .B1(n8990), .B2(n7553), .C1(
        n8991), .C2(n7552), .ZN(P2_U3265) );
  INV_X1 U9224 ( .A(n7555), .ZN(n9795) );
  OAI222_X1 U9225 ( .A1(n8990), .A2(n9795), .B1(P2_U3151), .B2(n5794), .C1(
        n7556), .C2(n8991), .ZN(P2_U3270) );
  INV_X1 U9226 ( .A(n7557), .ZN(n8994) );
  OAI222_X1 U9227 ( .A1(n6832), .A2(n7559), .B1(n7300), .B2(n8994), .C1(
        P1_U3086), .C2(n7558), .ZN(P1_U3329) );
  OAI222_X1 U9228 ( .A1(n8990), .A2(n7561), .B1(P2_U3151), .B2(n5791), .C1(
        n7560), .C2(n8991), .ZN(P2_U3271) );
  NAND2_X1 U9229 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n7564) );
  AOI211_X1 U9230 ( .C1(n7564), .C2(n7563), .A(n7562), .B(n9254), .ZN(n7569)
         );
  AOI211_X1 U9231 ( .C1(n7567), .C2(n7566), .A(n7565), .B(n9259), .ZN(n7568)
         );
  NOR2_X1 U9232 ( .A1(n7569), .A2(n7568), .ZN(n7571) );
  AOI22_X1 U9233 ( .A1(n9261), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n7570) );
  OAI211_X1 U9234 ( .C1(n7572), .C2(n9258), .A(n7571), .B(n7570), .ZN(P1_U3244) );
  NAND2_X1 U9235 ( .A1(n8976), .A2(n7579), .ZN(n7576) );
  OR2_X1 U9236 ( .A1(n7577), .A2(n6128), .ZN(n7575) );
  NOR2_X1 U9237 ( .A1(n7783), .A2(n7794), .ZN(n7779) );
  NOR2_X1 U9238 ( .A1(n7577), .A2(n7552), .ZN(n7578) );
  NOR2_X1 U9239 ( .A1(n8809), .A2(n8436), .ZN(n7774) );
  NOR2_X1 U9240 ( .A1(n7779), .A2(n7774), .ZN(n7614) );
  NAND3_X1 U9241 ( .A1(n7614), .A2(n7583), .A3(n5717), .ZN(n7584) );
  AND2_X1 U9242 ( .A1(n8809), .A2(n8436), .ZN(n7769) );
  INV_X1 U9243 ( .A(n7769), .ZN(n7611) );
  INV_X1 U9244 ( .A(n8586), .ZN(n8588) );
  NAND2_X1 U9245 ( .A1(n7757), .A2(n7758), .ZN(n8611) );
  INV_X1 U9246 ( .A(n7747), .ZN(n7587) );
  NOR2_X1 U9247 ( .A1(n7587), .A2(n7586), .ZN(n8643) );
  INV_X1 U9248 ( .A(n8708), .ZN(n8715) );
  INV_X1 U9249 ( .A(n8762), .ZN(n7606) );
  INV_X1 U9250 ( .A(n8748), .ZN(n8750) );
  NOR2_X1 U9251 ( .A1(n7591), .A2(n7590), .ZN(n7594) );
  NAND4_X1 U9252 ( .A1(n7594), .A2(n7593), .A3(n7592), .A4(n9978), .ZN(n7598)
         );
  OR4_X1 U9253 ( .A1(n7598), .A2(n7597), .A3(n7596), .A4(n7595), .ZN(n7602) );
  NOR4_X1 U9254 ( .A1(n7602), .A2(n7601), .A3(n7600), .A4(n7599), .ZN(n7604)
         );
  NAND4_X1 U9255 ( .A1(n8773), .A2(n7604), .A3(n7603), .A4(n7684), .ZN(n7605)
         );
  NOR4_X1 U9256 ( .A1(n8737), .A2(n7606), .A3(n8750), .A4(n7605), .ZN(n7607)
         );
  NAND4_X1 U9257 ( .A1(n8700), .A2(n7706), .A3(n8715), .A4(n7607), .ZN(n7608)
         );
  NOR4_X1 U9258 ( .A1(n8659), .A2(n5750), .A3(n8676), .A4(n7608), .ZN(n7609)
         );
  NAND4_X1 U9259 ( .A1(n8622), .A2(n8643), .A3(n8649), .A4(n7609), .ZN(n7610)
         );
  NOR4_X1 U9260 ( .A1(n8588), .A2(n8598), .A3(n8611), .A4(n7610), .ZN(n7612)
         );
  NAND4_X1 U9261 ( .A1(n7614), .A2(n7613), .A3(n7612), .A4(n7611), .ZN(n7615)
         );
  NOR2_X1 U9262 ( .A1(n7619), .A2(n7768), .ZN(n7620) );
  OAI22_X1 U9263 ( .A1(n7620), .A2(n7766), .B1(n8591), .B2(n7768), .ZN(n7763)
         );
  MUX2_X1 U9264 ( .A(n8816), .B(n7621), .S(n7768), .Z(n7764) );
  INV_X1 U9265 ( .A(n7764), .ZN(n7762) );
  MUX2_X1 U9266 ( .A(n8614), .B(n8607), .S(n7768), .Z(n7760) );
  NAND2_X1 U9267 ( .A1(n8681), .A2(n7723), .ZN(n7624) );
  NAND2_X1 U9268 ( .A1(n8668), .A2(n7727), .ZN(n7623) );
  MUX2_X1 U9269 ( .A(n7624), .B(n7623), .S(n7775), .Z(n7732) );
  XNOR2_X1 U9270 ( .A(n7625), .B(n7775), .ZN(n7705) );
  NAND2_X1 U9271 ( .A1(n7627), .A2(n7626), .ZN(n7632) );
  NAND3_X1 U9272 ( .A1(n7632), .A2(n7629), .A3(n8787), .ZN(n7628) );
  NAND2_X1 U9273 ( .A1(n7628), .A2(n7633), .ZN(n7631) );
  INV_X1 U9274 ( .A(n7629), .ZN(n7630) );
  MUX2_X1 U9275 ( .A(n7631), .B(n7630), .S(n7775), .Z(n7641) );
  INV_X1 U9276 ( .A(n7632), .ZN(n7634) );
  NAND3_X1 U9277 ( .A1(n7634), .A2(n7789), .A3(n7633), .ZN(n7636) );
  NAND2_X1 U9278 ( .A1(n7636), .A2(n7635), .ZN(n7640) );
  OAI21_X1 U9279 ( .B1(n7641), .B2(n7640), .A(n7639), .ZN(n7643) );
  NAND2_X1 U9280 ( .A1(n7643), .A2(n7642), .ZN(n7662) );
  INV_X1 U9281 ( .A(n7644), .ZN(n7646) );
  OAI211_X1 U9282 ( .C1(n7662), .C2(n7646), .A(n7664), .B(n7645), .ZN(n7648)
         );
  NAND2_X1 U9283 ( .A1(n7648), .A2(n7647), .ZN(n7649) );
  NAND3_X1 U9284 ( .A1(n7649), .A2(n7667), .A3(n7663), .ZN(n7651) );
  NAND2_X1 U9285 ( .A1(n7651), .A2(n7650), .ZN(n7657) );
  AND2_X1 U9286 ( .A1(n7672), .A2(n7670), .ZN(n7654) );
  AND2_X1 U9287 ( .A1(n7655), .A2(n7652), .ZN(n7653) );
  MUX2_X1 U9288 ( .A(n7654), .B(n7653), .S(n7775), .Z(n7674) );
  NAND2_X1 U9289 ( .A1(n7679), .A2(n7655), .ZN(n7656) );
  AOI21_X1 U9290 ( .B1(n7657), .B2(n7674), .A(n7656), .ZN(n7677) );
  INV_X1 U9291 ( .A(n7658), .ZN(n7661) );
  NAND3_X1 U9292 ( .A1(n7665), .A2(n7664), .A3(n7663), .ZN(n7668) );
  NAND3_X1 U9293 ( .A1(n7668), .A2(n7667), .A3(n7666), .ZN(n7671) );
  NAND3_X1 U9294 ( .A1(n7671), .A2(n7670), .A3(n7669), .ZN(n7675) );
  NAND2_X1 U9295 ( .A1(n7678), .A2(n7672), .ZN(n7673) );
  AOI21_X1 U9296 ( .B1(n7675), .B2(n7674), .A(n7673), .ZN(n7676) );
  MUX2_X1 U9297 ( .A(n7677), .B(n7676), .S(n7775), .Z(n7687) );
  NAND2_X1 U9298 ( .A1(n7683), .A2(n7678), .ZN(n7681) );
  NAND2_X1 U9299 ( .A1(n7682), .A2(n7679), .ZN(n7680) );
  MUX2_X1 U9300 ( .A(n7681), .B(n7680), .S(n7775), .Z(n7686) );
  MUX2_X1 U9301 ( .A(n7683), .B(n7682), .S(n7768), .Z(n7685) );
  OAI211_X1 U9302 ( .C1(n7687), .C2(n7686), .A(n7685), .B(n7684), .ZN(n7693)
         );
  NAND2_X1 U9303 ( .A1(n7688), .A2(n8392), .ZN(n7689) );
  MUX2_X1 U9304 ( .A(n7690), .B(n7689), .S(n7768), .Z(n7692) );
  AOI21_X1 U9305 ( .B1(n7693), .B2(n7692), .A(n7691), .ZN(n7697) );
  MUX2_X1 U9306 ( .A(n7695), .B(n7694), .S(n7775), .Z(n7696) );
  OAI21_X1 U9307 ( .B1(n7697), .B2(n7696), .A(n8762), .ZN(n7701) );
  MUX2_X1 U9308 ( .A(n7699), .B(n7698), .S(n7775), .Z(n7700) );
  NAND2_X1 U9309 ( .A1(n7701), .A2(n7700), .ZN(n7702) );
  NAND2_X1 U9310 ( .A1(n7707), .A2(n7706), .ZN(n7711) );
  NAND2_X1 U9311 ( .A1(n7725), .A2(n7708), .ZN(n7709) );
  INV_X1 U9312 ( .A(n7724), .ZN(n7717) );
  INV_X1 U9313 ( .A(n7712), .ZN(n7714) );
  INV_X1 U9314 ( .A(n5740), .ZN(n7713) );
  AOI211_X1 U9315 ( .C1(n7715), .C2(n7714), .A(n7775), .B(n7713), .ZN(n7716)
         );
  NOR2_X1 U9316 ( .A1(n7717), .A2(n7716), .ZN(n7721) );
  INV_X1 U9317 ( .A(n7718), .ZN(n7720) );
  NOR3_X1 U9318 ( .A1(n7721), .A2(n7720), .A3(n7719), .ZN(n7729) );
  INV_X1 U9319 ( .A(n7725), .ZN(n7726) );
  INV_X1 U9320 ( .A(n7727), .ZN(n7728) );
  OAI22_X1 U9321 ( .A1(n7732), .A2(n7731), .B1(n7775), .B2(n7730), .ZN(n7741)
         );
  INV_X1 U9322 ( .A(n7741), .ZN(n7737) );
  INV_X1 U9323 ( .A(n7740), .ZN(n7735) );
  OAI211_X1 U9324 ( .C1(n7735), .C2(n7734), .A(n7775), .B(n7733), .ZN(n7736)
         );
  OAI21_X1 U9325 ( .B1(n7737), .B2(n8676), .A(n7736), .ZN(n7739) );
  NAND3_X1 U9326 ( .A1(n7741), .A2(n8656), .A3(n7740), .ZN(n7743) );
  NAND2_X1 U9327 ( .A1(n7749), .A2(n7746), .ZN(n7748) );
  OAI21_X1 U9328 ( .B1(n7751), .B2(n7750), .A(n7749), .ZN(n7752) );
  MUX2_X1 U9329 ( .A(n7755), .B(n7754), .S(n7775), .Z(n7756) );
  MUX2_X1 U9330 ( .A(n7758), .B(n7757), .S(n7775), .Z(n7759) );
  INV_X1 U9331 ( .A(n7765), .ZN(n7761) );
  AOI21_X1 U9332 ( .B1(n7763), .B2(n7762), .A(n7761), .ZN(n7778) );
  NOR3_X1 U9333 ( .A1(n7776), .A2(n7769), .A3(n7766), .ZN(n7767) );
  OAI21_X1 U9334 ( .B1(n7778), .B2(n8898), .A(n7767), .ZN(n7772) );
  NOR2_X1 U9335 ( .A1(n7774), .A2(n7768), .ZN(n7770) );
  OAI21_X1 U9336 ( .B1(n7778), .B2(n8602), .A(n7777), .ZN(n7780) );
  XNOR2_X1 U9337 ( .A(n7785), .B(n7784), .ZN(n7792) );
  NAND3_X1 U9338 ( .A1(n7787), .A2(n7786), .A3(n8561), .ZN(n7788) );
  OAI211_X1 U9339 ( .C1(n7789), .C2(n7791), .A(n7788), .B(P2_B_REG_SCAN_IN), 
        .ZN(n7790) );
  OAI21_X1 U9340 ( .B1(n7792), .B2(n7791), .A(n7790), .ZN(P2_U3296) );
  NOR2_X1 U9341 ( .A1(n8807), .A2(n10070), .ZN(n8894) );
  AOI21_X1 U9342 ( .B1(n10070), .B2(P2_REG0_REG_30__SCAN_IN), .A(n8894), .ZN(
        n7795) );
  OAI21_X1 U9343 ( .B1(n8809), .B2(n8933), .A(n7795), .ZN(P2_U3457) );
  NAND2_X1 U9344 ( .A1(n7796), .A2(n8756), .ZN(n8579) );
  OAI21_X1 U9345 ( .B1(n8802), .B2(n8807), .A(n8579), .ZN(n8575) );
  AOI21_X1 U9346 ( .B1(n8802), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8575), .ZN(
        n7797) );
  OAI21_X1 U9347 ( .B1(n8809), .B2(n8791), .A(n7797), .ZN(P2_U3203) );
  NAND2_X1 U9348 ( .A1(n9620), .A2(n8289), .ZN(n7805) );
  XNOR2_X1 U9349 ( .A(n7987), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9336) );
  NAND2_X1 U9350 ( .A1(n9336), .A2(n7962), .ZN(n7803) );
  INV_X1 U9351 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9624) );
  NAND2_X1 U9352 ( .A1(n7798), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n7800) );
  NAND2_X1 U9353 ( .A1(n7989), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n7799) );
  OAI211_X1 U9354 ( .C1(n7992), .C2(n9624), .A(n7800), .B(n7799), .ZN(n7801)
         );
  INV_X1 U9355 ( .A(n7801), .ZN(n7802) );
  OR2_X1 U9356 ( .A1(n9627), .A2(n7307), .ZN(n7804) );
  NAND2_X1 U9357 ( .A1(n7805), .A2(n7804), .ZN(n7806) );
  XNOR2_X1 U9358 ( .A(n7806), .B(n8292), .ZN(n7809) );
  NOR2_X1 U9359 ( .A1(n9627), .A2(n8295), .ZN(n7807) );
  AOI21_X1 U9360 ( .B1(n9620), .B2(n6541), .A(n7807), .ZN(n7808) );
  NAND2_X1 U9361 ( .A1(n7809), .A2(n7808), .ZN(n8301) );
  OAI21_X1 U9362 ( .B1(n7809), .B2(n7808), .A(n8301), .ZN(n8011) );
  INV_X1 U9363 ( .A(n7811), .ZN(n7814) );
  INV_X1 U9364 ( .A(n7812), .ZN(n7813) );
  NAND2_X1 U9365 ( .A1(n7814), .A2(n7813), .ZN(n7815) );
  NAND2_X1 U9366 ( .A1(n9270), .A2(n8289), .ZN(n7818) );
  OR2_X1 U9367 ( .A1(n9580), .A2(n7307), .ZN(n7817) );
  NAND2_X1 U9368 ( .A1(n7818), .A2(n7817), .ZN(n7819) );
  XNOR2_X1 U9369 ( .A(n7819), .B(n8292), .ZN(n7822) );
  NOR2_X1 U9370 ( .A1(n9580), .A2(n8295), .ZN(n7820) );
  AOI21_X1 U9371 ( .B1(n9270), .B2(n6541), .A(n7820), .ZN(n7821) );
  NAND2_X1 U9372 ( .A1(n7822), .A2(n7821), .ZN(n7824) );
  OR2_X1 U9373 ( .A1(n7822), .A2(n7821), .ZN(n7823) );
  AND2_X1 U9374 ( .A1(n7824), .A2(n7823), .ZN(n9043) );
  NAND2_X1 U9375 ( .A1(n9042), .A2(n7824), .ZN(n9116) );
  NAND2_X1 U9376 ( .A1(n9272), .A2(n8289), .ZN(n7826) );
  OR2_X1 U9377 ( .A1(n9562), .A2(n7307), .ZN(n7825) );
  NAND2_X1 U9378 ( .A1(n7826), .A2(n7825), .ZN(n7827) );
  XNOR2_X1 U9379 ( .A(n7827), .B(n7998), .ZN(n7829) );
  NOR2_X1 U9380 ( .A1(n9562), .A2(n8295), .ZN(n7828) );
  AOI21_X1 U9381 ( .B1(n9272), .B2(n6541), .A(n7828), .ZN(n7830) );
  XNOR2_X1 U9382 ( .A(n7829), .B(n7830), .ZN(n9117) );
  INV_X1 U9383 ( .A(n7829), .ZN(n7831) );
  NAND2_X1 U9384 ( .A1(n7831), .A2(n7830), .ZN(n7832) );
  NAND2_X1 U9385 ( .A1(n7989), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7839) );
  INV_X1 U9386 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9728) );
  OR2_X1 U9387 ( .A1(n7992), .A2(n9728), .ZN(n7838) );
  INV_X1 U9388 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7833) );
  NAND2_X1 U9389 ( .A1(n7834), .A2(n7833), .ZN(n7835) );
  NAND2_X1 U9390 ( .A1(n7847), .A2(n7835), .ZN(n9558) );
  OR2_X1 U9391 ( .A1(n7988), .A2(n9558), .ZN(n7837) );
  OR2_X1 U9392 ( .A1(n7907), .A2(n6960), .ZN(n7836) );
  OAI22_X1 U9393 ( .A1(n9776), .A2(n7883), .B1(n9732), .B2(n7307), .ZN(n7840)
         );
  XNOR2_X1 U9394 ( .A(n7840), .B(n8292), .ZN(n7843) );
  OR2_X1 U9395 ( .A1(n9776), .A2(n7307), .ZN(n7842) );
  OR2_X1 U9396 ( .A1(n9732), .A2(n8295), .ZN(n7841) );
  AND2_X1 U9397 ( .A1(n7842), .A2(n7841), .ZN(n8999) );
  NAND2_X1 U9398 ( .A1(n8998), .A2(n8999), .ZN(n7845) );
  NAND2_X1 U9399 ( .A1(n7844), .A2(n7843), .ZN(n8997) );
  NAND2_X1 U9400 ( .A1(n7845), .A2(n8997), .ZN(n7858) );
  NAND2_X1 U9401 ( .A1(n9711), .A2(n8289), .ZN(n7854) );
  NAND2_X1 U9402 ( .A1(n7989), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7852) );
  INV_X1 U9403 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9180) );
  OR2_X1 U9404 ( .A1(n7992), .A2(n9180), .ZN(n7851) );
  INV_X1 U9405 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7846) );
  NAND2_X1 U9406 ( .A1(n7847), .A2(n7846), .ZN(n7848) );
  NAND2_X1 U9407 ( .A1(n7864), .A2(n7848), .ZN(n9539) );
  OR2_X1 U9408 ( .A1(n7988), .A2(n9539), .ZN(n7850) );
  INV_X1 U9409 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9540) );
  OR2_X1 U9410 ( .A1(n7907), .A2(n9540), .ZN(n7849) );
  NAND4_X1 U9411 ( .A1(n7852), .A2(n7851), .A3(n7850), .A4(n7849), .ZN(n9719)
         );
  NAND2_X1 U9412 ( .A1(n9719), .A2(n6541), .ZN(n7853) );
  NAND2_X1 U9413 ( .A1(n7854), .A2(n7853), .ZN(n7855) );
  XNOR2_X1 U9414 ( .A(n7855), .B(n8292), .ZN(n7859) );
  NAND2_X1 U9415 ( .A1(n7858), .A2(n7859), .ZN(n9152) );
  NAND2_X1 U9416 ( .A1(n9711), .A2(n6541), .ZN(n7857) );
  NAND2_X1 U9417 ( .A1(n9719), .A2(n7959), .ZN(n7856) );
  NAND2_X1 U9418 ( .A1(n7857), .A2(n7856), .ZN(n9155) );
  NAND2_X1 U9419 ( .A1(n9152), .A2(n9155), .ZN(n7862) );
  INV_X1 U9420 ( .A(n7858), .ZN(n7861) );
  INV_X1 U9421 ( .A(n7859), .ZN(n7860) );
  NAND2_X1 U9422 ( .A1(n7861), .A2(n7860), .ZN(n9153) );
  NAND2_X1 U9423 ( .A1(n7862), .A2(n9153), .ZN(n9063) );
  NAND2_X1 U9424 ( .A1(n9528), .A2(n8289), .ZN(n7871) );
  NAND2_X1 U9425 ( .A1(n7989), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n7869) );
  INV_X1 U9426 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9195) );
  OR2_X1 U9427 ( .A1(n7992), .A2(n9195), .ZN(n7868) );
  NAND2_X1 U9428 ( .A1(n7864), .A2(n7863), .ZN(n7865) );
  NAND2_X1 U9429 ( .A1(n9087), .A2(n7865), .ZN(n9523) );
  OR2_X1 U9430 ( .A1(n7988), .A2(n9523), .ZN(n7867) );
  INV_X1 U9431 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9524) );
  OR2_X1 U9432 ( .A1(n7981), .A2(n9524), .ZN(n7866) );
  OR2_X1 U9433 ( .A1(n9707), .A2(n7307), .ZN(n7870) );
  NAND2_X1 U9434 ( .A1(n7871), .A2(n7870), .ZN(n7872) );
  XNOR2_X1 U9435 ( .A(n7872), .B(n7998), .ZN(n7875) );
  NAND2_X1 U9436 ( .A1(n9528), .A2(n6541), .ZN(n7874) );
  OR2_X1 U9437 ( .A1(n9707), .A2(n8295), .ZN(n7873) );
  NAND2_X1 U9438 ( .A1(n7874), .A2(n7873), .ZN(n7876) );
  AND2_X1 U9439 ( .A1(n7875), .A2(n7876), .ZN(n9061) );
  INV_X1 U9440 ( .A(n7875), .ZN(n7878) );
  INV_X1 U9441 ( .A(n7876), .ZN(n7877) );
  NAND2_X1 U9442 ( .A1(n7878), .A2(n7877), .ZN(n9060) );
  NAND2_X1 U9443 ( .A1(n7989), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n7882) );
  INV_X1 U9444 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9237) );
  OR2_X1 U9445 ( .A1(n7992), .A2(n9237), .ZN(n7881) );
  INV_X1 U9446 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9497) );
  OR2_X1 U9447 ( .A1(n7907), .A2(n9497), .ZN(n7880) );
  INV_X1 U9448 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9089) );
  XNOR2_X1 U9449 ( .A(n9087), .B(n9089), .ZN(n9496) );
  OR2_X1 U9450 ( .A1(n7988), .A2(n9496), .ZN(n7879) );
  OAI22_X1 U9451 ( .A1(n9495), .A2(n7883), .B1(n9685), .B2(n7307), .ZN(n7884)
         );
  XNOR2_X1 U9452 ( .A(n7884), .B(n8292), .ZN(n9083) );
  OR2_X1 U9453 ( .A1(n9495), .A2(n7307), .ZN(n7886) );
  OR2_X1 U9454 ( .A1(n9685), .A2(n8295), .ZN(n7885) );
  AND2_X1 U9455 ( .A1(n9083), .A2(n9082), .ZN(n7890) );
  INV_X1 U9456 ( .A(n9083), .ZN(n7888) );
  INV_X1 U9457 ( .A(n9082), .ZN(n7887) );
  NAND2_X1 U9458 ( .A1(n7888), .A2(n7887), .ZN(n7889) );
  NAND2_X1 U9459 ( .A1(n9681), .A2(n8289), .ZN(n7900) );
  NAND2_X1 U9460 ( .A1(n7989), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n7898) );
  INV_X1 U9461 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n7891) );
  OR2_X1 U9462 ( .A1(n7992), .A2(n7891), .ZN(n7897) );
  NAND2_X1 U9463 ( .A1(n7906), .A2(n7892), .ZN(n7893) );
  NAND2_X1 U9464 ( .A1(n7934), .A2(n7893), .ZN(n9031) );
  OR2_X1 U9465 ( .A1(n7988), .A2(n9031), .ZN(n7896) );
  INV_X1 U9466 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n7894) );
  OR2_X1 U9467 ( .A1(n7981), .A2(n7894), .ZN(n7895) );
  NAND4_X1 U9468 ( .A1(n7898), .A2(n7897), .A3(n7896), .A4(n7895), .ZN(n9485)
         );
  NAND2_X1 U9469 ( .A1(n9485), .A2(n6541), .ZN(n7899) );
  NAND2_X1 U9470 ( .A1(n7900), .A2(n7899), .ZN(n7901) );
  XNOR2_X1 U9471 ( .A(n7901), .B(n8292), .ZN(n9026) );
  AND2_X1 U9472 ( .A1(n9485), .A2(n7959), .ZN(n7902) );
  AOI21_X1 U9473 ( .B1(n9681), .B2(n6541), .A(n7902), .ZN(n9025) );
  NOR2_X1 U9474 ( .A1(n9026), .A2(n9025), .ZN(n9106) );
  INV_X1 U9475 ( .A(n9106), .ZN(n7918) );
  NAND2_X1 U9476 ( .A1(n9689), .A2(n8289), .ZN(n7913) );
  NAND2_X1 U9477 ( .A1(n7989), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n7911) );
  INV_X1 U9478 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n7903) );
  OR2_X1 U9479 ( .A1(n7992), .A2(n7903), .ZN(n7910) );
  INV_X1 U9480 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n7904) );
  OAI21_X1 U9481 ( .B1(n9087), .B2(n9089), .A(n7904), .ZN(n7905) );
  NAND2_X1 U9482 ( .A1(n7906), .A2(n7905), .ZN(n9481) );
  OR2_X1 U9483 ( .A1(n7988), .A2(n9481), .ZN(n7909) );
  INV_X1 U9484 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9482) );
  OR2_X1 U9485 ( .A1(n7907), .A2(n9482), .ZN(n7908) );
  NAND4_X1 U9486 ( .A1(n7911), .A2(n7910), .A3(n7909), .A4(n7908), .ZN(n9505)
         );
  NAND2_X1 U9487 ( .A1(n9505), .A2(n6541), .ZN(n7912) );
  NAND2_X1 U9488 ( .A1(n7913), .A2(n7912), .ZN(n7914) );
  XNOR2_X1 U9489 ( .A(n7914), .B(n7998), .ZN(n9023) );
  NAND2_X1 U9490 ( .A1(n9689), .A2(n6541), .ZN(n7916) );
  NAND2_X1 U9491 ( .A1(n9505), .A2(n7959), .ZN(n7915) );
  NAND2_X1 U9492 ( .A1(n7916), .A2(n7915), .ZN(n9138) );
  INV_X1 U9493 ( .A(n9023), .ZN(n7922) );
  INV_X1 U9494 ( .A(n9138), .ZN(n7923) );
  AOI21_X1 U9495 ( .B1(n7922), .B2(n7923), .A(n9025), .ZN(n7926) );
  INV_X1 U9496 ( .A(n9026), .ZN(n7925) );
  OAI22_X1 U9497 ( .A1(n9448), .A2(n7307), .B1(n9437), .B2(n8295), .ZN(n7930)
         );
  NAND2_X1 U9498 ( .A1(n9676), .A2(n8289), .ZN(n7920) );
  NAND2_X1 U9499 ( .A1(n9666), .A2(n6541), .ZN(n7919) );
  NAND2_X1 U9500 ( .A1(n7920), .A2(n7919), .ZN(n7921) );
  XNOR2_X1 U9501 ( .A(n7921), .B(n7998), .ZN(n7929) );
  XOR2_X1 U9502 ( .A(n7930), .B(n7929), .Z(n9109) );
  NAND3_X1 U9503 ( .A1(n9025), .A2(n7923), .A3(n7922), .ZN(n7924) );
  OAI211_X1 U9504 ( .C1(n7926), .C2(n7925), .A(n9109), .B(n7924), .ZN(n7927)
         );
  INV_X1 U9505 ( .A(n7927), .ZN(n7928) );
  NAND2_X1 U9506 ( .A1(n4513), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n7939) );
  INV_X1 U9507 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n7932) );
  OR2_X1 U9508 ( .A1(n4602), .A2(n7932), .ZN(n7938) );
  INV_X1 U9509 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9037) );
  OAI21_X1 U9510 ( .B1(n7934), .B2(n9110), .A(n9037), .ZN(n7935) );
  NAND2_X1 U9511 ( .A1(n7935), .A2(n7945), .ZN(n9435) );
  OR2_X1 U9512 ( .A1(n7988), .A2(n9435), .ZN(n7937) );
  INV_X1 U9513 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9436) );
  OR2_X1 U9514 ( .A1(n7981), .A2(n9436), .ZN(n7936) );
  NAND4_X1 U9515 ( .A1(n7939), .A2(n7938), .A3(n7937), .A4(n7936), .ZN(n9657)
         );
  OAI22_X1 U9516 ( .A1(n9281), .A2(n7307), .B1(n9280), .B2(n8295), .ZN(n7943)
         );
  AOI22_X1 U9517 ( .A1(n9431), .A2(n8289), .B1(n6541), .B2(n9657), .ZN(n7940)
         );
  XNOR2_X1 U9518 ( .A(n7940), .B(n7998), .ZN(n7941) );
  XOR2_X1 U9519 ( .A(n7943), .B(n7941), .Z(n9036) );
  INV_X1 U9520 ( .A(n7941), .ZN(n7942) );
  NAND2_X1 U9521 ( .A1(n7989), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n7951) );
  INV_X1 U9522 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n7944) );
  OR2_X1 U9523 ( .A1(n7992), .A2(n7944), .ZN(n7950) );
  NAND2_X1 U9524 ( .A1(n7945), .A2(n9131), .ZN(n7946) );
  NAND2_X1 U9525 ( .A1(n7947), .A2(n7946), .ZN(n9418) );
  OR2_X1 U9526 ( .A1(n7988), .A2(n9418), .ZN(n7949) );
  INV_X1 U9527 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9419) );
  OR2_X1 U9528 ( .A1(n7981), .A2(n9419), .ZN(n7948) );
  AOI22_X1 U9529 ( .A1(n9422), .A2(n8289), .B1(n6541), .B2(n9667), .ZN(n7952)
         );
  XNOR2_X1 U9530 ( .A(n7952), .B(n7998), .ZN(n7957) );
  NAND2_X1 U9531 ( .A1(n9408), .A2(n8289), .ZN(n7954) );
  NAND2_X1 U9532 ( .A1(n9658), .A2(n6541), .ZN(n7953) );
  NAND2_X1 U9533 ( .A1(n7954), .A2(n7953), .ZN(n7955) );
  XNOR2_X1 U9534 ( .A(n7955), .B(n7998), .ZN(n7971) );
  AND2_X1 U9535 ( .A1(n9658), .A2(n7959), .ZN(n7956) );
  AOI21_X1 U9536 ( .B1(n9408), .B2(n6541), .A(n7956), .ZN(n7969) );
  XNOR2_X1 U9537 ( .A(n7971), .B(n7969), .ZN(n9007) );
  AOI22_X1 U9538 ( .A1(n9422), .A2(n6541), .B1(n7959), .B2(n9667), .ZN(n9129)
         );
  NAND2_X1 U9539 ( .A1(n7960), .A2(n9101), .ZN(n7961) );
  AND2_X1 U9540 ( .A1(n7976), .A2(n7961), .ZN(n9391) );
  NAND2_X1 U9541 ( .A1(n9391), .A2(n7962), .ZN(n7965) );
  AOI22_X1 U9542 ( .A1(n4513), .A2(P1_REG1_REG_24__SCAN_IN), .B1(n7989), .B2(
        P1_REG0_REG_24__SCAN_IN), .ZN(n7964) );
  NAND2_X1 U9543 ( .A1(n7798), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n7963) );
  AOI22_X1 U9544 ( .A1(n9390), .A2(n8289), .B1(n6541), .B2(n9649), .ZN(n7966)
         );
  XOR2_X1 U9545 ( .A(n7998), .B(n7966), .Z(n7968) );
  OAI22_X1 U9546 ( .A1(n9763), .A2(n7307), .B1(n9374), .B2(n8295), .ZN(n7967)
         );
  NOR2_X1 U9547 ( .A1(n7968), .A2(n7967), .ZN(n7973) );
  AOI21_X1 U9548 ( .B1(n7968), .B2(n7967), .A(n7973), .ZN(n9096) );
  INV_X1 U9549 ( .A(n7969), .ZN(n7970) );
  NAND2_X1 U9550 ( .A1(n7971), .A2(n7970), .ZN(n9097) );
  INV_X1 U9551 ( .A(n7973), .ZN(n7974) );
  NAND2_X1 U9552 ( .A1(n9095), .A2(n7974), .ZN(n9053) );
  INV_X1 U9553 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9371) );
  INV_X1 U9554 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n7975) );
  NAND2_X1 U9555 ( .A1(n7976), .A2(n7975), .ZN(n7977) );
  NAND2_X1 U9556 ( .A1(n7985), .A2(n7977), .ZN(n9370) );
  OR2_X1 U9557 ( .A1(n9370), .A2(n7988), .ZN(n7980) );
  AOI22_X1 U9558 ( .A1(n4513), .A2(P1_REG1_REG_25__SCAN_IN), .B1(n7989), .B2(
        P1_REG0_REG_25__SCAN_IN), .ZN(n7979) );
  OAI211_X1 U9559 ( .C1(n7981), .C2(n9371), .A(n7980), .B(n7979), .ZN(n9386)
         );
  OAI22_X1 U9560 ( .A1(n9639), .A2(n7307), .B1(n9626), .B2(n8295), .ZN(n8002)
         );
  NAND2_X1 U9561 ( .A1(n9376), .A2(n8289), .ZN(n7983) );
  NAND2_X1 U9562 ( .A1(n9386), .A2(n6541), .ZN(n7982) );
  NAND2_X1 U9563 ( .A1(n7983), .A2(n7982), .ZN(n7984) );
  XNOR2_X1 U9564 ( .A(n7984), .B(n7998), .ZN(n8001) );
  XOR2_X1 U9565 ( .A(n8002), .B(n8001), .Z(n9054) );
  NAND2_X1 U9566 ( .A1(n9053), .A2(n9054), .ZN(n9052) );
  NAND2_X1 U9567 ( .A1(n9355), .A2(n8289), .ZN(n7997) );
  NAND2_X1 U9568 ( .A1(n7985), .A2(n9146), .ZN(n7986) );
  NAND2_X1 U9569 ( .A1(n7987), .A2(n7986), .ZN(n9356) );
  INV_X1 U9570 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9634) );
  NAND2_X1 U9571 ( .A1(n7989), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n7991) );
  NAND2_X1 U9572 ( .A1(n7798), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n7990) );
  OAI211_X1 U9573 ( .C1(n7992), .C2(n9634), .A(n7991), .B(n7990), .ZN(n7993)
         );
  INV_X1 U9574 ( .A(n7993), .ZN(n7994) );
  NAND2_X1 U9575 ( .A1(n9636), .A2(n6541), .ZN(n7996) );
  NAND2_X1 U9576 ( .A1(n7997), .A2(n7996), .ZN(n7999) );
  XNOR2_X1 U9577 ( .A(n7999), .B(n7998), .ZN(n8007) );
  NOR2_X1 U9578 ( .A1(n9341), .A2(n8295), .ZN(n8000) );
  AOI21_X1 U9579 ( .B1(n9355), .B2(n6541), .A(n8000), .ZN(n8005) );
  XNOR2_X1 U9580 ( .A(n8007), .B(n8005), .ZN(n9144) );
  INV_X1 U9581 ( .A(n8001), .ZN(n8004) );
  INV_X1 U9582 ( .A(n8002), .ZN(n8003) );
  NAND2_X1 U9583 ( .A1(n8004), .A2(n8003), .ZN(n9145) );
  INV_X1 U9584 ( .A(n8005), .ZN(n8006) );
  INV_X1 U9585 ( .A(n8009), .ZN(n8008) );
  NAND2_X1 U9586 ( .A1(n4872), .A2(n8008), .ZN(n8010) );
  AOI21_X1 U9587 ( .B1(n8011), .B2(n8010), .A(n8307), .ZN(n8017) );
  INV_X1 U9588 ( .A(n9336), .ZN(n8013) );
  OAI22_X1 U9589 ( .A1(n9157), .A2(n8013), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8012), .ZN(n8015) );
  OAI22_X1 U9590 ( .A1(n9607), .A2(n9158), .B1(n9341), .B2(n9159), .ZN(n8014)
         );
  AOI211_X1 U9591 ( .C1(n9620), .C2(n9162), .A(n8015), .B(n8014), .ZN(n8016)
         );
  OAI21_X1 U9592 ( .B1(n8017), .B2(n9164), .A(n8016), .ZN(P1_U3214) );
  XNOR2_X1 U9593 ( .A(n8733), .B(n5869), .ZN(n8029) );
  INV_X1 U9594 ( .A(n8029), .ZN(n8030) );
  INV_X1 U9595 ( .A(n8018), .ZN(n8019) );
  NOR2_X1 U9596 ( .A1(n8019), .A2(n8775), .ZN(n8388) );
  XNOR2_X1 U9597 ( .A(n8971), .B(n8051), .ZN(n8020) );
  XNOR2_X1 U9598 ( .A(n8020), .B(n8763), .ZN(n8387) );
  NAND2_X1 U9599 ( .A1(n8020), .A2(n8021), .ZN(n8022) );
  NAND2_X1 U9600 ( .A1(n8386), .A2(n8022), .ZN(n8318) );
  XNOR2_X1 U9601 ( .A(n8964), .B(n5869), .ZN(n8024) );
  XNOR2_X1 U9602 ( .A(n8024), .B(n8774), .ZN(n8319) );
  XNOR2_X1 U9603 ( .A(n8958), .B(n8051), .ZN(n8025) );
  XNOR2_X1 U9604 ( .A(n8025), .B(n8764), .ZN(n8425) );
  NAND2_X1 U9605 ( .A1(n8426), .A2(n8425), .ZN(n8424) );
  XNOR2_X1 U9606 ( .A(n5741), .B(n8051), .ZN(n8027) );
  XOR2_X1 U9607 ( .A(n8752), .B(n8027), .Z(n8354) );
  INV_X1 U9608 ( .A(n8027), .ZN(n8028) );
  NOR2_X1 U9609 ( .A1(n8028), .A2(n8752), .ZN(n8363) );
  XNOR2_X1 U9610 ( .A(n8029), .B(n8740), .ZN(n8362) );
  XNOR2_X1 U9611 ( .A(n8873), .B(n8051), .ZN(n8031) );
  XNOR2_X1 U9612 ( .A(n8031), .B(n8694), .ZN(n8405) );
  XNOR2_X1 U9613 ( .A(n8863), .B(n8051), .ZN(n8032) );
  XNOR2_X1 U9614 ( .A(n8032), .B(n8855), .ZN(n8332) );
  XNOR2_X1 U9615 ( .A(n8937), .B(n8051), .ZN(n8034) );
  XOR2_X1 U9616 ( .A(n8862), .B(n8034), .Z(n8380) );
  INV_X1 U9617 ( .A(n8034), .ZN(n8035) );
  XNOR2_X1 U9618 ( .A(n8845), .B(n5869), .ZN(n8036) );
  XNOR2_X1 U9619 ( .A(n8036), .B(n8856), .ZN(n8339) );
  AND2_X1 U9620 ( .A1(n8036), .A2(n8663), .ZN(n8037) );
  XNOR2_X1 U9621 ( .A(n8665), .B(n8051), .ZN(n8038) );
  XNOR2_X1 U9622 ( .A(n8038), .B(n8846), .ZN(n8398) );
  INV_X1 U9623 ( .A(n8038), .ZN(n8040) );
  XNOR2_X1 U9624 ( .A(n8922), .B(n8048), .ZN(n8042) );
  XNOR2_X1 U9625 ( .A(n8376), .B(n8051), .ZN(n8043) );
  XNOR2_X1 U9626 ( .A(n8043), .B(n8650), .ZN(n8372) );
  XNOR2_X1 U9627 ( .A(n8830), .B(n8051), .ZN(n8044) );
  XOR2_X1 U9628 ( .A(n8613), .B(n8044), .Z(n8347) );
  INV_X1 U9629 ( .A(n8044), .ZN(n8045) );
  XNOR2_X1 U9630 ( .A(n8907), .B(n8051), .ZN(n8046) );
  XNOR2_X1 U9631 ( .A(n8046), .B(n8631), .ZN(n8414) );
  NAND2_X1 U9632 ( .A1(n8046), .A2(n8827), .ZN(n8047) );
  XNOR2_X1 U9633 ( .A(n8607), .B(n8048), .ZN(n8049) );
  NAND2_X1 U9634 ( .A1(n8049), .A2(n8614), .ZN(n8050) );
  OAI21_X1 U9635 ( .B1(n8049), .B2(n8614), .A(n8050), .ZN(n8310) );
  NAND2_X1 U9636 ( .A1(n8311), .A2(n8050), .ZN(n8053) );
  XNOR2_X1 U9637 ( .A(n8586), .B(n8051), .ZN(n8052) );
  XNOR2_X1 U9638 ( .A(n8053), .B(n8052), .ZN(n8059) );
  INV_X1 U9639 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8054) );
  OAI22_X1 U9640 ( .A1(n8590), .A2(n8409), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8054), .ZN(n8057) );
  INV_X1 U9641 ( .A(n8595), .ZN(n8055) );
  OAI22_X1 U9642 ( .A1(n8591), .A2(n8427), .B1(n8055), .B2(n8428), .ZN(n8056)
         );
  AOI211_X1 U9643 ( .C1(n8898), .C2(n8419), .A(n8057), .B(n8056), .ZN(n8058)
         );
  OAI21_X1 U9644 ( .B1(n8059), .B2(n8421), .A(n8058), .ZN(P2_U3160) );
  NAND2_X1 U9645 ( .A1(n9620), .A2(n9627), .ZN(n9306) );
  OR2_X1 U9646 ( .A1(n9620), .A2(n9627), .ZN(n8196) );
  OR2_X1 U9647 ( .A1(n9355), .A2(n9341), .ZN(n8197) );
  OR2_X1 U9648 ( .A1(n9408), .A2(n9285), .ZN(n8199) );
  NAND2_X1 U9649 ( .A1(n9661), .A2(n9667), .ZN(n8060) );
  NAND2_X1 U9650 ( .A1(n8199), .A2(n8060), .ZN(n8162) );
  NAND2_X1 U9651 ( .A1(n8162), .A2(n9381), .ZN(n8061) );
  NAND2_X1 U9652 ( .A1(n9302), .A2(n8061), .ZN(n8062) );
  NAND2_X1 U9653 ( .A1(n9390), .A2(n9374), .ZN(n8169) );
  NAND2_X1 U9654 ( .A1(n8062), .A2(n8169), .ZN(n8067) );
  NOR2_X1 U9655 ( .A1(n9431), .A2(n9280), .ZN(n8155) );
  NAND2_X1 U9656 ( .A1(n9431), .A2(n9280), .ZN(n9297) );
  NAND2_X1 U9657 ( .A1(n9676), .A2(n9437), .ZN(n8200) );
  AND2_X1 U9658 ( .A1(n9297), .A2(n8200), .ZN(n8158) );
  NAND2_X1 U9659 ( .A1(n9422), .A2(n9405), .ZN(n9298) );
  NAND2_X1 U9660 ( .A1(n9381), .A2(n9298), .ZN(n8160) );
  INV_X1 U9661 ( .A(n8160), .ZN(n8063) );
  OAI211_X1 U9662 ( .C1(n8155), .C2(n8158), .A(n8169), .B(n8063), .ZN(n8064)
         );
  NAND2_X1 U9663 ( .A1(n9376), .A2(n9626), .ZN(n9303) );
  NAND2_X1 U9664 ( .A1(n9355), .A2(n9341), .ZN(n9305) );
  INV_X1 U9665 ( .A(n9305), .ZN(n8178) );
  INV_X1 U9666 ( .A(n8155), .ZN(n8065) );
  NAND2_X1 U9667 ( .A1(n8065), .A2(n9296), .ZN(n8152) );
  INV_X1 U9668 ( .A(n8152), .ZN(n8066) );
  NAND3_X1 U9669 ( .A1(n8067), .A2(n8198), .A3(n8066), .ZN(n8071) );
  OR2_X1 U9670 ( .A1(n8068), .A2(n9607), .ZN(n8195) );
  OAI21_X1 U9671 ( .B1(n8069), .B2(n4702), .A(n8195), .ZN(n8070) );
  OR2_X1 U9672 ( .A1(n8101), .A2(n9319), .ZN(n8184) );
  INV_X1 U9673 ( .A(n8254), .ZN(n8103) );
  NAND2_X1 U9674 ( .A1(n9528), .A2(n9707), .ZN(n8244) );
  NAND2_X1 U9675 ( .A1(n9711), .A2(n9525), .ZN(n8242) );
  NAND2_X1 U9676 ( .A1(n9568), .A2(n9732), .ZN(n8241) );
  AND2_X1 U9677 ( .A1(n8242), .A2(n8241), .ZN(n8072) );
  AND2_X1 U9678 ( .A1(n8244), .A2(n8072), .ZN(n8134) );
  INV_X1 U9679 ( .A(n8073), .ZN(n8074) );
  OAI211_X1 U9680 ( .C1(n9016), .C2(n8076), .A(n8075), .B(n8074), .ZN(n8083)
         );
  AOI22_X1 U9681 ( .A1(n8078), .A2(n9177), .B1(n8077), .B2(n9175), .ZN(n8080)
         );
  NAND3_X1 U9682 ( .A1(n8080), .A2(n8108), .A3(n8079), .ZN(n8082) );
  OAI21_X1 U9683 ( .B1(n8083), .B2(n8082), .A(n8081), .ZN(n8085) );
  OAI211_X1 U9684 ( .C1(n8086), .C2(n8085), .A(n8139), .B(n8084), .ZN(n8088)
         );
  AND2_X1 U9685 ( .A1(n8128), .A2(n8087), .ZN(n8143) );
  NAND2_X1 U9686 ( .A1(n8132), .A2(n8127), .ZN(n8142) );
  AOI21_X1 U9687 ( .B1(n8088), .B2(n8143), .A(n8142), .ZN(n8090) );
  NAND2_X1 U9688 ( .A1(n9272), .A2(n9562), .ZN(n8206) );
  NAND2_X1 U9689 ( .A1(n8206), .A2(n9574), .ZN(n8089) );
  OR2_X1 U9690 ( .A1(n9568), .A2(n9732), .ZN(n8145) );
  OAI21_X1 U9691 ( .B1(n8090), .B2(n8089), .A(n8145), .ZN(n8092) );
  OR2_X1 U9692 ( .A1(n9528), .A2(n9707), .ZN(n8204) );
  INV_X1 U9693 ( .A(n8204), .ZN(n8091) );
  AOI211_X1 U9694 ( .C1(n8134), .C2(n8092), .A(n8091), .B(n4761), .ZN(n8098)
         );
  INV_X1 U9695 ( .A(n8134), .ZN(n8093) );
  OR2_X1 U9696 ( .A1(n9272), .A2(n9562), .ZN(n8240) );
  OR2_X1 U9697 ( .A1(n8093), .A2(n8240), .ZN(n8096) );
  OR2_X1 U9698 ( .A1(n9711), .A2(n9525), .ZN(n8205) );
  INV_X1 U9699 ( .A(n8205), .ZN(n8094) );
  NAND2_X1 U9700 ( .A1(n8244), .A2(n8094), .ZN(n8095) );
  AND2_X1 U9701 ( .A1(n8096), .A2(n8095), .ZN(n8136) );
  NAND2_X1 U9702 ( .A1(n9689), .A2(n9277), .ZN(n9464) );
  NAND2_X1 U9703 ( .A1(n9696), .A2(n9685), .ZN(n8203) );
  AND2_X1 U9704 ( .A1(n9464), .A2(n8203), .ZN(n8149) );
  INV_X1 U9705 ( .A(n8149), .ZN(n8097) );
  AOI21_X1 U9706 ( .B1(n8098), .B2(n8136), .A(n8097), .ZN(n8100) );
  OR2_X1 U9707 ( .A1(n9681), .A2(n9686), .ZN(n8250) );
  OR2_X1 U9708 ( .A1(n9689), .A2(n9277), .ZN(n8202) );
  AND2_X1 U9709 ( .A1(n8250), .A2(n8202), .ZN(n8150) );
  INV_X1 U9710 ( .A(n8150), .ZN(n8099) );
  NAND2_X1 U9711 ( .A1(n9681), .A2(n9686), .ZN(n8201) );
  OAI211_X1 U9712 ( .C1(n8100), .C2(n8099), .A(n8251), .B(n8201), .ZN(n8102)
         );
  NAND2_X1 U9713 ( .A1(n9265), .A2(n9311), .ZN(n8233) );
  NAND2_X1 U9714 ( .A1(n8101), .A2(n9319), .ZN(n8185) );
  NAND2_X1 U9715 ( .A1(n8233), .A2(n8185), .ZN(n8255) );
  AOI21_X1 U9716 ( .B1(n8103), .B2(n8102), .A(n8255), .ZN(n8104) );
  NOR2_X1 U9717 ( .A1(n9265), .A2(n9311), .ZN(n8258) );
  NOR2_X1 U9718 ( .A1(n8104), .A2(n8258), .ZN(n8106) );
  NAND2_X1 U9719 ( .A1(n8105), .A2(n8252), .ZN(n8276) );
  OAI21_X1 U9720 ( .B1(n8106), .B2(n8273), .A(n8276), .ZN(n8107) );
  XNOR2_X1 U9721 ( .A(n8107), .B(n9343), .ZN(n8269) );
  INV_X1 U9722 ( .A(n8195), .ZN(n8183) );
  INV_X1 U9723 ( .A(n8277), .ZN(n8194) );
  NAND2_X1 U9724 ( .A1(n8175), .A2(n8194), .ZN(n8177) );
  INV_X1 U9725 ( .A(n8177), .ZN(n8182) );
  INV_X1 U9726 ( .A(n8108), .ZN(n8110) );
  OAI211_X1 U9727 ( .C1(n7046), .C2(n8110), .A(n8207), .B(n8109), .ZN(n8111)
         );
  NAND2_X1 U9728 ( .A1(n8111), .A2(n8112), .ZN(n8114) );
  INV_X1 U9729 ( .A(n8112), .ZN(n8113) );
  INV_X1 U9730 ( .A(n8115), .ZN(n8116) );
  INV_X1 U9731 ( .A(n8214), .ZN(n8117) );
  MUX2_X1 U9732 ( .A(n8118), .B(n8117), .S(n8277), .Z(n8119) );
  NAND2_X1 U9733 ( .A1(n8120), .A2(n8119), .ZN(n8125) );
  AND2_X1 U9734 ( .A1(n8218), .A2(n8121), .ZN(n8122) );
  MUX2_X1 U9735 ( .A(n8123), .B(n8122), .S(n8194), .Z(n8124) );
  NAND2_X1 U9736 ( .A1(n8125), .A2(n8124), .ZN(n8138) );
  AOI21_X1 U9737 ( .B1(n8138), .B2(n8140), .A(n8126), .ZN(n8130) );
  NAND2_X1 U9738 ( .A1(n8127), .A2(n8139), .ZN(n8129) );
  OAI211_X1 U9739 ( .C1(n8130), .C2(n8129), .A(n8128), .B(n9574), .ZN(n8133)
         );
  INV_X1 U9740 ( .A(n8206), .ZN(n8131) );
  AOI21_X1 U9741 ( .B1(n8133), .B2(n8132), .A(n8131), .ZN(n8135) );
  INV_X1 U9742 ( .A(n9552), .ZN(n9554) );
  OAI21_X1 U9743 ( .B1(n8135), .B2(n9554), .A(n8134), .ZN(n8137) );
  NAND3_X1 U9744 ( .A1(n8137), .A2(n8136), .A3(n8204), .ZN(n8148) );
  NAND2_X1 U9745 ( .A1(n8138), .A2(n8218), .ZN(n8141) );
  NAND3_X1 U9746 ( .A1(n8141), .A2(n8140), .A3(n8139), .ZN(n8144) );
  INV_X1 U9747 ( .A(n9574), .ZN(n8238) );
  NAND2_X1 U9748 ( .A1(n8146), .A2(n8242), .ZN(n8147) );
  OAI21_X1 U9749 ( .B1(n4531), .B2(n4761), .A(n8149), .ZN(n8151) );
  NAND2_X1 U9750 ( .A1(n8151), .A2(n8150), .ZN(n8154) );
  AND2_X1 U9751 ( .A1(n8200), .A2(n8201), .ZN(n8153) );
  AOI21_X1 U9752 ( .B1(n8154), .B2(n8153), .A(n8152), .ZN(n8168) );
  NAND3_X1 U9753 ( .A1(n4531), .A2(n8202), .A3(n8246), .ZN(n8156) );
  NAND3_X1 U9754 ( .A1(n8156), .A2(n8201), .A3(n9464), .ZN(n8157) );
  NAND3_X1 U9755 ( .A1(n8157), .A2(n8250), .A3(n9296), .ZN(n8159) );
  XNOR2_X1 U9756 ( .A(n9422), .B(n9667), .ZN(n9415) );
  NOR3_X1 U9757 ( .A1(n8160), .A2(n8194), .A3(n9415), .ZN(n8161) );
  NOR2_X1 U9758 ( .A1(n8162), .A2(n8277), .ZN(n8165) );
  INV_X1 U9759 ( .A(n9415), .ZN(n9413) );
  NAND2_X1 U9760 ( .A1(n9658), .A2(n8277), .ZN(n8163) );
  OAI22_X1 U9761 ( .A1(n9381), .A2(n8277), .B1(n9408), .B2(n8163), .ZN(n8164)
         );
  AOI21_X1 U9762 ( .B1(n8165), .B2(n9413), .A(n8164), .ZN(n8166) );
  MUX2_X1 U9763 ( .A(n9302), .B(n8169), .S(n8277), .Z(n8170) );
  INV_X1 U9764 ( .A(n8176), .ZN(n8172) );
  INV_X1 U9765 ( .A(n8198), .ZN(n8171) );
  OAI211_X1 U9766 ( .C1(n8172), .C2(n8171), .A(n9305), .B(n9303), .ZN(n8173)
         );
  NAND4_X1 U9767 ( .A1(n8173), .A2(n8196), .A3(n8197), .A4(n8277), .ZN(n8174)
         );
  NAND2_X1 U9768 ( .A1(n8176), .A2(n9303), .ZN(n8179) );
  AOI211_X1 U9769 ( .C1(n8198), .C2(n8179), .A(n8178), .B(n8177), .ZN(n8180)
         );
  NAND2_X1 U9770 ( .A1(n8186), .A2(n8276), .ZN(n8193) );
  AOI21_X1 U9771 ( .B1(n8257), .B2(n8187), .A(n8273), .ZN(n8192) );
  NOR2_X1 U9772 ( .A1(n8188), .A2(n9311), .ZN(n8191) );
  AOI22_X1 U9773 ( .A1(n8193), .A2(n8192), .B1(n8191), .B2(n8190), .ZN(n8274)
         );
  NAND2_X1 U9774 ( .A1(n8197), .A2(n9305), .ZN(n9304) );
  NAND2_X1 U9775 ( .A1(n8198), .A2(n9303), .ZN(n9367) );
  NAND2_X1 U9776 ( .A1(n8250), .A2(n8201), .ZN(n9460) );
  INV_X1 U9777 ( .A(n9460), .ZN(n9463) );
  NAND2_X1 U9778 ( .A1(n8202), .A2(n9464), .ZN(n9476) );
  NAND2_X1 U9779 ( .A1(n8246), .A2(n8203), .ZN(n9500) );
  NAND2_X1 U9780 ( .A1(n8204), .A2(n8244), .ZN(n9517) );
  NAND2_X1 U9781 ( .A1(n8240), .A2(n8206), .ZN(n9576) );
  INV_X1 U9782 ( .A(n9576), .ZN(n8225) );
  NAND2_X1 U9783 ( .A1(n8207), .A2(n8267), .ZN(n8208) );
  NOR2_X1 U9784 ( .A1(n8209), .A2(n8208), .ZN(n8211) );
  NAND4_X1 U9785 ( .A1(n4528), .A2(n8212), .A3(n8211), .A4(n8210), .ZN(n8216)
         );
  NAND2_X1 U9786 ( .A1(n8213), .A2(n6673), .ZN(n8215) );
  NOR3_X1 U9787 ( .A1(n8216), .A2(n8215), .A3(n8214), .ZN(n8221) );
  INV_X1 U9788 ( .A(n8217), .ZN(n8220) );
  NAND4_X1 U9789 ( .A1(n8221), .A2(n8220), .A3(n8219), .A4(n8218), .ZN(n8222)
         );
  NOR3_X1 U9790 ( .A1(n8236), .A2(n8223), .A3(n8222), .ZN(n8224) );
  NAND4_X1 U9791 ( .A1(n9534), .A2(n9552), .A3(n8225), .A4(n8224), .ZN(n8226)
         );
  OR3_X1 U9792 ( .A1(n9500), .A2(n9517), .A3(n8226), .ZN(n8227) );
  NOR2_X1 U9793 ( .A1(n9476), .A2(n8227), .ZN(n8228) );
  AND3_X1 U9794 ( .A1(n9454), .A2(n9463), .A3(n8228), .ZN(n8229) );
  XNOR2_X1 U9795 ( .A(n9431), .B(n9280), .ZN(n9427) );
  INV_X1 U9796 ( .A(n9427), .ZN(n9430) );
  NAND4_X1 U9797 ( .A1(n9399), .A2(n8229), .A3(n9415), .A4(n9430), .ZN(n8230)
         );
  OR3_X1 U9798 ( .A1(n9367), .A2(n8230), .A3(n9382), .ZN(n8231) );
  NOR2_X1 U9799 ( .A1(n9304), .A2(n8231), .ZN(n8232) );
  NAND4_X1 U9800 ( .A1(n8233), .A2(n9322), .A3(n9344), .A4(n8232), .ZN(n8234)
         );
  NOR4_X1 U9801 ( .A1(n8273), .A2(n9308), .A3(n8258), .A4(n8234), .ZN(n8235)
         );
  NAND2_X1 U9802 ( .A1(n8235), .A2(n8276), .ZN(n8265) );
  OR2_X2 U9803 ( .A1(n8237), .A2(n8236), .ZN(n9575) );
  NOR2_X1 U9804 ( .A1(n9576), .A2(n8238), .ZN(n8239) );
  NAND2_X1 U9805 ( .A1(n8243), .A2(n8242), .ZN(n9521) );
  INV_X1 U9806 ( .A(n9517), .ZN(n9520) );
  NAND2_X1 U9807 ( .A1(n9521), .A2(n9520), .ZN(n9519) );
  INV_X1 U9808 ( .A(n8244), .ZN(n9501) );
  NOR2_X1 U9809 ( .A1(n9500), .A2(n9501), .ZN(n8245) );
  INV_X1 U9810 ( .A(n9464), .ZN(n8248) );
  NOR2_X1 U9811 ( .A1(n9460), .A2(n8248), .ZN(n8249) );
  NAND2_X1 U9812 ( .A1(n9474), .A2(n8249), .ZN(n9462) );
  NAND2_X1 U9813 ( .A1(n9462), .A2(n8250), .ZN(n9455) );
  AND2_X1 U9814 ( .A1(n8251), .A2(n9455), .ZN(n8253) );
  AOI21_X1 U9815 ( .B1(n8258), .B2(n8257), .A(n8256), .ZN(n8262) );
  NAND2_X1 U9816 ( .A1(n8265), .A2(n8263), .ZN(n8264) );
  MUX2_X1 U9817 ( .A(n8265), .B(n8264), .S(n9343), .Z(n8266) );
  NAND3_X1 U9818 ( .A1(n8271), .A2(n8270), .A3(n5110), .ZN(n8272) );
  OR2_X1 U9819 ( .A1(n8285), .A2(n5954), .ZN(n8279) );
  NAND3_X1 U9820 ( .A1(n8272), .A2(P1_B_REG_SCAN_IN), .A3(n8279), .ZN(n8284)
         );
  INV_X1 U9821 ( .A(n8273), .ZN(n8282) );
  INV_X1 U9822 ( .A(n8274), .ZN(n8275) );
  OAI21_X1 U9823 ( .B1(n8277), .B2(n8276), .A(n8275), .ZN(n8281) );
  NOR2_X1 U9824 ( .A1(n8279), .A2(n8278), .ZN(n8280) );
  OAI211_X1 U9825 ( .C1(n8282), .C2(n9343), .A(n8281), .B(n8280), .ZN(n8283)
         );
  OAI222_X1 U9826 ( .A1(n8990), .A2(n8288), .B1(P2_U3151), .B2(n8287), .C1(
        n8286), .C2(n8991), .ZN(P2_U3266) );
  NAND2_X1 U9827 ( .A1(n8068), .A2(n8289), .ZN(n8291) );
  OR2_X1 U9828 ( .A1(n9607), .A2(n7307), .ZN(n8290) );
  NAND2_X1 U9829 ( .A1(n8291), .A2(n8290), .ZN(n8293) );
  XNOR2_X1 U9830 ( .A(n8293), .B(n8292), .ZN(n8297) );
  NAND2_X1 U9831 ( .A1(n8068), .A2(n6541), .ZN(n8294) );
  OAI21_X1 U9832 ( .B1(n9607), .B2(n8295), .A(n8294), .ZN(n8296) );
  XNOR2_X1 U9833 ( .A(n8297), .B(n8296), .ZN(n8298) );
  INV_X1 U9834 ( .A(n8298), .ZN(n8302) );
  NAND3_X1 U9835 ( .A1(n8302), .A2(n9143), .A3(n8301), .ZN(n8306) );
  INV_X1 U9836 ( .A(n9627), .ZN(n9360) );
  NAND2_X1 U9837 ( .A1(n9360), .A2(n9077), .ZN(n8300) );
  AOI22_X1 U9838 ( .A1(n9123), .A2(n9328), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n8299) );
  OAI211_X1 U9839 ( .C1(n9319), .C2(n9158), .A(n8300), .B(n8299), .ZN(n8304)
         );
  NOR3_X1 U9840 ( .A1(n8302), .A2(n9164), .A3(n8301), .ZN(n8303) );
  AOI211_X1 U9841 ( .C1(n8068), .C2(n9162), .A(n8304), .B(n8303), .ZN(n8305)
         );
  INV_X1 U9842 ( .A(n8308), .ZN(n8985) );
  OAI222_X1 U9843 ( .A1(n6832), .A2(n10285), .B1(P1_U3086), .B2(n5968), .C1(
        n8985), .C2(n7300), .ZN(P1_U3327) );
  AOI21_X1 U9844 ( .B1(n8309), .B2(n8310), .A(n8421), .ZN(n8312) );
  NAND2_X1 U9845 ( .A1(n8312), .A2(n8311), .ZN(n8317) );
  INV_X1 U9846 ( .A(n8603), .ZN(n8314) );
  AOI22_X1 U9847 ( .A1(n8631), .A2(n8431), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8313) );
  OAI21_X1 U9848 ( .B1(n8314), .B2(n8428), .A(n8313), .ZN(n8315) );
  AOI21_X1 U9849 ( .B1(n8406), .B2(n8602), .A(n8315), .ZN(n8316) );
  OAI211_X1 U9850 ( .C1(n4801), .C2(n8434), .A(n8317), .B(n8316), .ZN(P2_U3154) );
  XOR2_X1 U9851 ( .A(n8319), .B(n8318), .Z(n8324) );
  INV_X1 U9852 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10396) );
  OAI22_X1 U9853 ( .A1(n8427), .A2(n8357), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10396), .ZN(n8320) );
  AOI21_X1 U9854 ( .B1(n8431), .B2(n8763), .A(n8320), .ZN(n8321) );
  OAI21_X1 U9855 ( .B1(n8766), .B2(n8428), .A(n8321), .ZN(n8322) );
  AOI21_X1 U9856 ( .B1(n8964), .B2(n8419), .A(n8322), .ZN(n8323) );
  OAI21_X1 U9857 ( .B1(n8324), .B2(n8421), .A(n8323), .ZN(P2_U3155) );
  XNOR2_X1 U9858 ( .A(n8325), .B(n8637), .ZN(n8330) );
  AOI22_X1 U9859 ( .A1(n8846), .A2(n8431), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8327) );
  NAND2_X1 U9860 ( .A1(n8415), .A2(n8653), .ZN(n8326) );
  OAI211_X1 U9861 ( .C1(n8826), .C2(n8427), .A(n8327), .B(n8326), .ZN(n8328)
         );
  AOI21_X1 U9862 ( .B1(n8922), .B2(n8419), .A(n8328), .ZN(n8329) );
  OAI21_X1 U9863 ( .B1(n8330), .B2(n8421), .A(n8329), .ZN(P2_U3156) );
  INV_X1 U9864 ( .A(n8863), .ZN(n8338) );
  OAI211_X1 U9865 ( .C1(n8333), .C2(n8332), .A(n8331), .B(n8423), .ZN(n8337)
         );
  NAND2_X1 U9866 ( .A1(n8431), .A2(n8694), .ZN(n8334) );
  NAND2_X1 U9867 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8568) );
  OAI211_X1 U9868 ( .C1(n8699), .C2(n8427), .A(n8334), .B(n8568), .ZN(n8335)
         );
  AOI21_X1 U9869 ( .B1(n8697), .B2(n8415), .A(n8335), .ZN(n8336) );
  OAI211_X1 U9870 ( .C1(n8338), .C2(n8434), .A(n8337), .B(n8336), .ZN(P2_U3159) );
  XOR2_X1 U9871 ( .A(n8340), .B(n8339), .Z(n8345) );
  AOI22_X1 U9872 ( .A1(n8846), .A2(n8406), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8342) );
  NAND2_X1 U9873 ( .A1(n8415), .A2(n8671), .ZN(n8341) );
  OAI211_X1 U9874 ( .C1(n8699), .C2(n8409), .A(n8342), .B(n8341), .ZN(n8343)
         );
  AOI21_X1 U9875 ( .B1(n8845), .B2(n8419), .A(n8343), .ZN(n8344) );
  OAI21_X1 U9876 ( .B1(n8345), .B2(n8421), .A(n8344), .ZN(P2_U3163) );
  XOR2_X1 U9877 ( .A(n8347), .B(n8346), .Z(n8352) );
  AOI22_X1 U9878 ( .A1(n8650), .A2(n8431), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8349) );
  NAND2_X1 U9879 ( .A1(n8625), .A2(n8415), .ZN(n8348) );
  OAI211_X1 U9880 ( .C1(n8827), .C2(n8427), .A(n8349), .B(n8348), .ZN(n8350)
         );
  AOI21_X1 U9881 ( .B1(n8830), .B2(n8419), .A(n8350), .ZN(n8351) );
  OAI21_X1 U9882 ( .B1(n8352), .B2(n8421), .A(n8351), .ZN(P2_U3165) );
  AOI21_X1 U9883 ( .B1(n8354), .B2(n8353), .A(n8364), .ZN(n8360) );
  AOI22_X1 U9884 ( .A1(n8406), .A2(n8740), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3151), .ZN(n8356) );
  NAND2_X1 U9885 ( .A1(n8415), .A2(n8744), .ZN(n8355) );
  OAI211_X1 U9886 ( .C1(n8357), .C2(n8409), .A(n8356), .B(n8355), .ZN(n8358)
         );
  AOI21_X1 U9887 ( .B1(n5741), .B2(n8419), .A(n8358), .ZN(n8359) );
  OAI21_X1 U9888 ( .B1(n8360), .B2(n8421), .A(n8359), .ZN(P2_U3166) );
  INV_X1 U9889 ( .A(n8733), .ZN(n8877) );
  INV_X1 U9890 ( .A(n8361), .ZN(n8366) );
  NOR3_X1 U9891 ( .A1(n8364), .A2(n8363), .A3(n8362), .ZN(n8365) );
  OAI21_X1 U9892 ( .B1(n8366), .B2(n8365), .A(n8423), .ZN(n8370) );
  AOI22_X1 U9893 ( .A1(n8406), .A2(n8694), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3151), .ZN(n8367) );
  OAI21_X1 U9894 ( .B1(n8726), .B2(n8409), .A(n8367), .ZN(n8368) );
  AOI21_X1 U9895 ( .B1(n8729), .B2(n8415), .A(n8368), .ZN(n8369) );
  OAI211_X1 U9896 ( .C1(n8877), .C2(n8434), .A(n8370), .B(n8369), .ZN(P2_U3168) );
  XOR2_X1 U9897 ( .A(n8372), .B(n8371), .Z(n8378) );
  AOI22_X1 U9898 ( .A1(n8613), .A2(n8406), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8374) );
  NAND2_X1 U9899 ( .A1(n8639), .A2(n8415), .ZN(n8373) );
  OAI211_X1 U9900 ( .C1(n8637), .C2(n8409), .A(n8374), .B(n8373), .ZN(n8375)
         );
  AOI21_X1 U9901 ( .B1(n8376), .B2(n8419), .A(n8375), .ZN(n8377) );
  OAI21_X1 U9902 ( .B1(n8378), .B2(n8421), .A(n8377), .ZN(P2_U3169) );
  AOI21_X1 U9903 ( .B1(n8380), .B2(n8379), .A(n4563), .ZN(n8385) );
  AOI22_X1 U9904 ( .A1(n8406), .A2(n8856), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8382) );
  NAND2_X1 U9905 ( .A1(n8415), .A2(n8685), .ZN(n8381) );
  OAI211_X1 U9906 ( .C1(n8869), .C2(n8409), .A(n8382), .B(n8381), .ZN(n8383)
         );
  AOI21_X1 U9907 ( .B1(n8937), .B2(n8419), .A(n8383), .ZN(n8384) );
  OAI21_X1 U9908 ( .B1(n8385), .B2(n8421), .A(n8384), .ZN(P2_U3173) );
  INV_X1 U9909 ( .A(n8971), .ZN(n8779) );
  INV_X1 U9910 ( .A(n8386), .ZN(n8390) );
  NOR3_X1 U9911 ( .A1(n4585), .A2(n8388), .A3(n8387), .ZN(n8389) );
  OAI21_X1 U9912 ( .B1(n8390), .B2(n8389), .A(n8423), .ZN(n8396) );
  INV_X1 U9913 ( .A(n8777), .ZN(n8394) );
  AOI22_X1 U9914 ( .A1(n8406), .A2(n8774), .B1(P2_REG3_REG_13__SCAN_IN), .B2(
        P2_U3151), .ZN(n8391) );
  OAI21_X1 U9915 ( .B1(n8392), .B2(n8409), .A(n8391), .ZN(n8393) );
  AOI21_X1 U9916 ( .B1(n8394), .B2(n8415), .A(n8393), .ZN(n8395) );
  OAI211_X1 U9917 ( .C1(n8779), .C2(n8434), .A(n8396), .B(n8395), .ZN(P2_U3174) );
  OAI211_X1 U9918 ( .C1(n8399), .C2(n8398), .A(n8397), .B(n8423), .ZN(n8403)
         );
  AOI22_X1 U9919 ( .A1(n8431), .A2(n8856), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8400) );
  OAI21_X1 U9920 ( .B1(n8637), .B2(n8427), .A(n8400), .ZN(n8401) );
  AOI21_X1 U9921 ( .B1(n8660), .B2(n8415), .A(n8401), .ZN(n8402) );
  OAI211_X1 U9922 ( .C1(n8929), .C2(n8434), .A(n8403), .B(n8402), .ZN(P2_U3175) );
  XOR2_X1 U9923 ( .A(n8405), .B(n8404), .Z(n8412) );
  AOI22_X1 U9924 ( .A1(n8406), .A2(n8855), .B1(P2_REG3_REG_18__SCAN_IN), .B2(
        P2_U3151), .ZN(n8408) );
  NAND2_X1 U9925 ( .A1(n8415), .A2(n8709), .ZN(n8407) );
  OAI211_X1 U9926 ( .C1(n8868), .C2(n8409), .A(n8408), .B(n8407), .ZN(n8410)
         );
  AOI21_X1 U9927 ( .B1(n8873), .B2(n8419), .A(n8410), .ZN(n8411) );
  OAI21_X1 U9928 ( .B1(n8412), .B2(n8421), .A(n8411), .ZN(P2_U3178) );
  XOR2_X1 U9929 ( .A(n8414), .B(n8413), .Z(n8422) );
  AOI22_X1 U9930 ( .A1(n8613), .A2(n8431), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8417) );
  NAND2_X1 U9931 ( .A1(n8617), .A2(n8415), .ZN(n8416) );
  OAI211_X1 U9932 ( .C1(n8590), .C2(n8427), .A(n8417), .B(n8416), .ZN(n8418)
         );
  AOI21_X1 U9933 ( .B1(n8907), .B2(n8419), .A(n8418), .ZN(n8420) );
  OAI21_X1 U9934 ( .B1(n8422), .B2(n8421), .A(n8420), .ZN(P2_U3180) );
  INV_X1 U9935 ( .A(n8958), .ZN(n8435) );
  OAI211_X1 U9936 ( .C1(n8426), .C2(n8425), .A(n8424), .B(n8423), .ZN(n8433)
         );
  NAND2_X1 U9937 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8493) );
  OAI21_X1 U9938 ( .B1(n8427), .B2(n8726), .A(n8493), .ZN(n8430) );
  NOR2_X1 U9939 ( .A1(n8428), .A2(n8754), .ZN(n8429) );
  AOI211_X1 U9940 ( .C1(n8431), .C2(n8774), .A(n8430), .B(n8429), .ZN(n8432)
         );
  OAI211_X1 U9941 ( .C1(n8435), .C2(n8434), .A(n8433), .B(n8432), .ZN(P2_U3181) );
  MUX2_X1 U9942 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8436), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9943 ( .A(n8602), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8531), .Z(
        P2_U3519) );
  MUX2_X1 U9944 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8614), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9945 ( .A(n8631), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8531), .Z(
        P2_U3517) );
  MUX2_X1 U9946 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8613), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9947 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8650), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9948 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8846), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9949 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8856), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9950 ( .A(n8862), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8531), .Z(
        P2_U3511) );
  MUX2_X1 U9951 ( .A(n8855), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8531), .Z(
        P2_U3510) );
  MUX2_X1 U9952 ( .A(n8694), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8531), .Z(
        P2_U3509) );
  MUX2_X1 U9953 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8740), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9954 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8752), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9955 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8764), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9956 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8774), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9957 ( .A(n8775), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8531), .Z(
        P2_U3503) );
  MUX2_X1 U9958 ( .A(n8437), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8531), .Z(
        P2_U3502) );
  MUX2_X1 U9959 ( .A(n10041), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8531), .Z(
        P2_U3501) );
  MUX2_X1 U9960 ( .A(n8438), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8531), .Z(
        P2_U3500) );
  MUX2_X1 U9961 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n10044), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U9962 ( .A(n8439), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8531), .Z(
        P2_U3498) );
  MUX2_X1 U9963 ( .A(n8440), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8531), .Z(
        P2_U3497) );
  MUX2_X1 U9964 ( .A(n8441), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8531), .Z(
        P2_U3496) );
  MUX2_X1 U9965 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8442), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U9966 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n10008), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U9967 ( .A(n9998), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8531), .Z(
        P2_U3493) );
  MUX2_X1 U9968 ( .A(n5870), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8531), .Z(
        P2_U3492) );
  MUX2_X1 U9969 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8796), .S(P2_U3893), .Z(
        P2_U3491) );
  OAI21_X1 U9970 ( .B1(n8445), .B2(n8444), .A(n8443), .ZN(n8446) );
  NAND2_X1 U9971 ( .A1(n8446), .A2(n9967), .ZN(n8468) );
  INV_X1 U9972 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n8448) );
  OAI21_X1 U9973 ( .B1(n9888), .B2(n8448), .A(n8447), .ZN(n8449) );
  AOI21_X1 U9974 ( .B1(n8492), .B2(n8450), .A(n8449), .ZN(n8467) );
  INV_X1 U9975 ( .A(n8451), .ZN(n8454) );
  INV_X1 U9976 ( .A(n8452), .ZN(n8453) );
  NOR3_X1 U9977 ( .A1(n8455), .A2(n8454), .A3(n8453), .ZN(n8456) );
  OAI21_X1 U9978 ( .B1(n8457), .B2(n8456), .A(n9877), .ZN(n8466) );
  INV_X1 U9979 ( .A(n8458), .ZN(n8459) );
  NOR3_X1 U9980 ( .A1(n8461), .A2(n8460), .A3(n8459), .ZN(n8464) );
  OAI21_X1 U9981 ( .B1(n8464), .B2(n8463), .A(n8462), .ZN(n8465) );
  NAND4_X1 U9982 ( .A1(n8468), .A2(n8467), .A3(n8466), .A4(n8465), .ZN(
        P2_U3190) );
  NOR2_X1 U9983 ( .A1(n8496), .A2(n8469), .ZN(n8471) );
  NAND2_X1 U9984 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n9905), .ZN(n8472) );
  OAI21_X1 U9985 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n9905), .A(n8472), .ZN(
        n9893) );
  NOR2_X1 U9986 ( .A1(n8500), .A2(n8473), .ZN(n8474) );
  XOR2_X1 U9987 ( .A(n8473), .B(n9923), .Z(n9914) );
  NOR2_X1 U9988 ( .A1(n9915), .A2(n9914), .ZN(n9913) );
  NAND2_X1 U9989 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n9940), .ZN(n8475) );
  OAI21_X1 U9990 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n9940), .A(n8475), .ZN(
        n9931) );
  NOR2_X1 U9991 ( .A1(n9932), .A2(n9931), .ZN(n9930) );
  INV_X1 U9992 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8476) );
  AOI21_X1 U9993 ( .B1(n8477), .B2(n8476), .A(n8512), .ZN(n8510) );
  MUX2_X1 U9994 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8561), .Z(n8521) );
  XNOR2_X1 U9995 ( .A(n8521), .B(n8536), .ZN(n8491) );
  MUX2_X1 U9996 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8561), .Z(n8479) );
  OR2_X1 U9997 ( .A1(n8479), .A2(n9940), .ZN(n8489) );
  XNOR2_X1 U9998 ( .A(n8479), .B(n8478), .ZN(n9928) );
  MUX2_X1 U9999 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8561), .Z(n8480) );
  OR2_X1 U10000 ( .A1(n8480), .A2(n9923), .ZN(n8488) );
  XNOR2_X1 U10001 ( .A(n8480), .B(n8500), .ZN(n9911) );
  MUX2_X1 U10002 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8561), .Z(n8482) );
  OR2_X1 U10003 ( .A1(n8482), .A2(n9905), .ZN(n8487) );
  XNOR2_X1 U10004 ( .A(n8482), .B(n8481), .ZN(n9897) );
  OR2_X1 U10005 ( .A1(n8484), .A2(n8483), .ZN(n8486) );
  NAND2_X1 U10006 ( .A1(n8486), .A2(n8485), .ZN(n9896) );
  NAND2_X1 U10007 ( .A1(n9897), .A2(n9896), .ZN(n9895) );
  NAND2_X1 U10008 ( .A1(n8487), .A2(n9895), .ZN(n9910) );
  NAND2_X1 U10009 ( .A1(n9911), .A2(n9910), .ZN(n9909) );
  NAND2_X1 U10010 ( .A1(n8488), .A2(n9909), .ZN(n9927) );
  NAND2_X1 U10011 ( .A1(n9928), .A2(n9927), .ZN(n9926) );
  NAND2_X1 U10012 ( .A1(n8489), .A2(n9926), .ZN(n8490) );
  OAI21_X1 U10013 ( .B1(n8491), .B2(n8490), .A(n8523), .ZN(n8508) );
  INV_X1 U10014 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8495) );
  NAND2_X1 U10015 ( .A1(n8492), .A2(n8536), .ZN(n8494) );
  OAI211_X1 U10016 ( .C1(n8495), .C2(n9888), .A(n8494), .B(n8493), .ZN(n8507)
         );
  NOR2_X1 U10017 ( .A1(n8496), .A2(n4547), .ZN(n8498) );
  NAND2_X1 U10018 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n9905), .ZN(n8499) );
  OAI21_X1 U10019 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n9905), .A(n8499), .ZN(
        n9891) );
  NAND2_X1 U10020 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n9940), .ZN(n8502) );
  OAI21_X1 U10021 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n9940), .A(n8502), .ZN(
        n9924) );
  AOI21_X1 U10022 ( .B1(n8884), .B2(n8504), .A(n8538), .ZN(n8505) );
  NOR2_X1 U10023 ( .A1(n8505), .A2(n9971), .ZN(n8506) );
  AOI211_X1 U10024 ( .C1(n9967), .C2(n8508), .A(n8507), .B(n8506), .ZN(n8509)
         );
  OAI21_X1 U10025 ( .B1(n8510), .B2(n9963), .A(n8509), .ZN(P2_U3197) );
  NOR2_X1 U10026 ( .A1(n8536), .A2(n8511), .ZN(n8513) );
  NAND2_X1 U10027 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n9956), .ZN(n8514) );
  OAI21_X1 U10028 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n9956), .A(n8514), .ZN(
        n9944) );
  NOR2_X1 U10029 ( .A1(n8541), .A2(n8515), .ZN(n8516) );
  XOR2_X1 U10030 ( .A(n8515), .B(n9976), .Z(n9962) );
  NOR2_X1 U10031 ( .A1(n8519), .A2(n9962), .ZN(n9961) );
  NAND2_X1 U10032 ( .A1(n8544), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8550) );
  OAI21_X1 U10033 ( .B1(n8544), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8550), .ZN(
        n8517) );
  AOI21_X1 U10034 ( .B1(n8518), .B2(n8517), .A(n8552), .ZN(n8549) );
  MUX2_X1 U10035 ( .A(n8519), .B(n9960), .S(n8561), .Z(n8527) );
  XNOR2_X1 U10036 ( .A(n8527), .B(n9976), .ZN(n9966) );
  MUX2_X1 U10037 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8561), .Z(n8520) );
  OR2_X1 U10038 ( .A1(n8520), .A2(n9956), .ZN(n8525) );
  XNOR2_X1 U10039 ( .A(n8520), .B(n8539), .ZN(n9948) );
  INV_X1 U10040 ( .A(n8521), .ZN(n8522) );
  NAND2_X1 U10041 ( .A1(n8536), .A2(n8522), .ZN(n8524) );
  NAND2_X1 U10042 ( .A1(n8524), .A2(n8523), .ZN(n9947) );
  NAND2_X1 U10043 ( .A1(n9948), .A2(n9947), .ZN(n9946) );
  NAND2_X1 U10044 ( .A1(n8525), .A2(n9946), .ZN(n9965) );
  NAND2_X1 U10045 ( .A1(n9966), .A2(n9965), .ZN(n9964) );
  INV_X1 U10046 ( .A(n9964), .ZN(n8526) );
  MUX2_X1 U10047 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8561), .Z(n8528) );
  NOR2_X1 U10048 ( .A1(n8529), .A2(n8528), .ZN(n8559) );
  INV_X1 U10049 ( .A(n8559), .ZN(n8530) );
  NAND2_X1 U10050 ( .A1(n8529), .A2(n8528), .ZN(n8557) );
  NAND2_X1 U10051 ( .A1(n8530), .A2(n8557), .ZN(n8532) );
  OAI21_X1 U10052 ( .B1(n8532), .B2(n8531), .A(n9977), .ZN(n8547) );
  INV_X1 U10053 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10114) );
  NAND3_X1 U10054 ( .A1(n8532), .A2(n9967), .A3(n8544), .ZN(n8534) );
  INV_X1 U10055 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10475) );
  OR2_X1 U10056 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10475), .ZN(n8533) );
  OAI211_X1 U10057 ( .C1(n10114), .C2(n9888), .A(n8534), .B(n8533), .ZN(n8546)
         );
  NOR2_X1 U10058 ( .A1(n8536), .A2(n8535), .ZN(n8537) );
  AOI22_X1 U10059 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8539), .B1(n9956), .B2(
        n8881), .ZN(n9942) );
  NOR2_X1 U10060 ( .A1(n8541), .A2(n8542), .ZN(n8543) );
  NAND2_X1 U10061 ( .A1(n8544), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8553) );
  OAI21_X1 U10062 ( .B1(n8544), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8553), .ZN(
        n8545) );
  OAI21_X1 U10063 ( .B1(n8549), .B2(n9963), .A(n8548), .ZN(P2_U3200) );
  INV_X1 U10064 ( .A(n8550), .ZN(n8551) );
  MUX2_X1 U10065 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n5546), .S(n5139), .Z(n8563) );
  INV_X1 U10066 ( .A(n8553), .ZN(n8554) );
  XNOR2_X1 U10067 ( .A(n5139), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8560) );
  XNOR2_X1 U10068 ( .A(n8556), .B(n8560), .ZN(n8572) );
  INV_X1 U10069 ( .A(n8560), .ZN(n8562) );
  MUX2_X1 U10070 ( .A(n8563), .B(n8562), .S(n8561), .Z(n8564) );
  XNOR2_X1 U10071 ( .A(n8565), .B(n8564), .ZN(n8567) );
  NOR2_X1 U10072 ( .A1(n8567), .A2(n8566), .ZN(n8571) );
  NAND2_X1 U10073 ( .A1(n9957), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8569) );
  OAI211_X1 U10074 ( .C1(n9977), .C2(n5139), .A(n8569), .B(n8568), .ZN(n8570)
         );
  OAI21_X1 U10075 ( .B1(n9963), .B2(n8574), .A(n8573), .ZN(P2_U3201) );
  AOI21_X1 U10076 ( .B1(n8802), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8575), .ZN(
        n8576) );
  OAI21_X1 U10077 ( .B1(n7582), .B2(n8791), .A(n8576), .ZN(P2_U3202) );
  INV_X1 U10078 ( .A(n8577), .ZN(n8585) );
  NAND2_X1 U10079 ( .A1(n8802), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8578) );
  OAI211_X1 U10080 ( .C1(n8816), .C2(n8712), .A(n8579), .B(n8578), .ZN(n8580)
         );
  AOI21_X1 U10081 ( .B1(n8581), .B2(n8757), .A(n8580), .ZN(n8584) );
  NAND2_X1 U10082 ( .A1(n8582), .A2(n8793), .ZN(n8583) );
  OAI211_X1 U10083 ( .C1(n8585), .C2(n8802), .A(n8584), .B(n8583), .ZN(
        P2_U3204) );
  XNOR2_X1 U10084 ( .A(n8587), .B(n8586), .ZN(n8901) );
  XNOR2_X1 U10085 ( .A(n8589), .B(n8588), .ZN(n8593) );
  OAI22_X1 U10086 ( .A1(n8591), .A2(n10025), .B1(n8590), .B2(n10027), .ZN(
        n8592) );
  AOI21_X1 U10087 ( .B1(n8593), .B2(n10005), .A(n8592), .ZN(n8897) );
  MUX2_X1 U10088 ( .A(n8897), .B(n8594), .S(n8802), .Z(n8597) );
  AOI22_X1 U10089 ( .A1(n8898), .A2(n8757), .B1(n8756), .B2(n8595), .ZN(n8596)
         );
  OAI211_X1 U10090 ( .C1(n8901), .C2(n8784), .A(n8597), .B(n8596), .ZN(
        P2_U3205) );
  XNOR2_X1 U10091 ( .A(n8599), .B(n8598), .ZN(n8817) );
  XNOR2_X1 U10092 ( .A(n8601), .B(n8600), .ZN(n8820) );
  NAND2_X1 U10093 ( .A1(n8820), .A2(n8684), .ZN(n8609) );
  NAND2_X1 U10094 ( .A1(n8602), .A2(n8795), .ZN(n8605) );
  AOI22_X1 U10095 ( .A1(n8603), .A2(n8756), .B1(n8802), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8604) );
  OAI211_X1 U10096 ( .C1(n8827), .C2(n8712), .A(n8605), .B(n8604), .ZN(n8606)
         );
  AOI21_X1 U10097 ( .B1(n8607), .B2(n8745), .A(n8606), .ZN(n8608) );
  OAI211_X1 U10098 ( .C1(n8817), .C2(n8784), .A(n8609), .B(n8608), .ZN(
        P2_U3206) );
  XOR2_X1 U10099 ( .A(n8611), .B(n8610), .Z(n8910) );
  XNOR2_X1 U10100 ( .A(n8612), .B(n8611), .ZN(n8615) );
  AOI222_X1 U10101 ( .A1(n10005), .A2(n8615), .B1(n8614), .B2(n10042), .C1(
        n8613), .C2(n10043), .ZN(n8905) );
  MUX2_X1 U10102 ( .A(n8616), .B(n8905), .S(n8728), .Z(n8619) );
  AOI22_X1 U10103 ( .A1(n8907), .A2(n8745), .B1(n8756), .B2(n8617), .ZN(n8618)
         );
  OAI211_X1 U10104 ( .C1(n8910), .C2(n8784), .A(n8619), .B(n8618), .ZN(
        P2_U3207) );
  XNOR2_X1 U10105 ( .A(n8621), .B(n8620), .ZN(n8914) );
  XNOR2_X1 U10106 ( .A(n8623), .B(n8622), .ZN(n8624) );
  NOR2_X1 U10107 ( .A1(n8624), .A2(n9979), .ZN(n8828) );
  INV_X1 U10108 ( .A(n8830), .ZN(n8627) );
  INV_X1 U10109 ( .A(n8625), .ZN(n8626) );
  OAI22_X1 U10110 ( .A1(n8627), .A2(n8778), .B1(n8626), .B2(n8788), .ZN(n8628)
         );
  OAI21_X1 U10111 ( .B1(n8828), .B2(n8628), .A(n8728), .ZN(n8633) );
  OAI22_X1 U10112 ( .A1(n8826), .A2(n8712), .B1(n8728), .B2(n8629), .ZN(n8630)
         );
  AOI21_X1 U10113 ( .B1(n8795), .B2(n8631), .A(n8630), .ZN(n8632) );
  OAI211_X1 U10114 ( .C1(n8914), .C2(n8784), .A(n8633), .B(n8632), .ZN(
        P2_U3208) );
  NOR2_X1 U10115 ( .A1(n8916), .A2(n8778), .ZN(n8638) );
  XOR2_X1 U10116 ( .A(n8643), .B(n8634), .Z(n8635) );
  OAI222_X1 U10117 ( .A1(n10027), .A2(n8637), .B1(n10025), .B2(n8636), .C1(
        n8635), .C2(n9979), .ZN(n8915) );
  AOI211_X1 U10118 ( .C1(n8756), .C2(n8639), .A(n8638), .B(n8915), .ZN(n8646)
         );
  NAND2_X1 U10119 ( .A1(n8641), .A2(n8640), .ZN(n8642) );
  XOR2_X1 U10120 ( .A(n8643), .B(n8642), .Z(n8917) );
  INV_X1 U10121 ( .A(n8917), .ZN(n8644) );
  AOI22_X1 U10122 ( .A1(n8644), .A2(n8793), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n8802), .ZN(n8645) );
  OAI21_X1 U10123 ( .B1(n8646), .B2(n8802), .A(n8645), .ZN(P2_U3209) );
  XOR2_X1 U10124 ( .A(n8647), .B(n8649), .Z(n8925) );
  XOR2_X1 U10125 ( .A(n8649), .B(n8648), .Z(n8651) );
  AOI222_X1 U10126 ( .A1(n10005), .A2(n8651), .B1(n8846), .B2(n10043), .C1(
        n8650), .C2(n10042), .ZN(n8920) );
  MUX2_X1 U10127 ( .A(n8652), .B(n8920), .S(n8728), .Z(n8655) );
  AOI22_X1 U10128 ( .A1(n8922), .A2(n8757), .B1(n8756), .B2(n8653), .ZN(n8654)
         );
  OAI211_X1 U10129 ( .C1(n8925), .C2(n8784), .A(n8655), .B(n8654), .ZN(
        P2_U3210) );
  XNOR2_X1 U10130 ( .A(n8657), .B(n8656), .ZN(n8840) );
  XNOR2_X1 U10131 ( .A(n8658), .B(n8659), .ZN(n8842) );
  NAND2_X1 U10132 ( .A1(n8842), .A2(n8684), .ZN(n8667) );
  NAND2_X1 U10133 ( .A1(n8838), .A2(n8795), .ZN(n8662) );
  AOI22_X1 U10134 ( .A1(n8756), .A2(n8660), .B1(n8802), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n8661) );
  OAI211_X1 U10135 ( .C1(n8663), .C2(n8712), .A(n8662), .B(n8661), .ZN(n8664)
         );
  AOI21_X1 U10136 ( .B1(n8665), .B2(n8757), .A(n8664), .ZN(n8666) );
  OAI211_X1 U10137 ( .C1(n8840), .C2(n8784), .A(n8667), .B(n8666), .ZN(
        P2_U3211) );
  INV_X1 U10138 ( .A(n8668), .ZN(n8669) );
  NOR2_X1 U10139 ( .A1(n4552), .A2(n8669), .ZN(n8670) );
  XOR2_X1 U10140 ( .A(n8676), .B(n8670), .Z(n8848) );
  NAND2_X1 U10141 ( .A1(n8795), .A2(n8846), .ZN(n8673) );
  AOI22_X1 U10142 ( .A1(n8802), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8756), .B2(
        n8671), .ZN(n8672) );
  OAI211_X1 U10143 ( .C1(n8712), .C2(n8699), .A(n8673), .B(n8672), .ZN(n8674)
         );
  AOI21_X1 U10144 ( .B1(n8845), .B2(n8745), .A(n8674), .ZN(n8678) );
  XNOR2_X1 U10145 ( .A(n8675), .B(n8676), .ZN(n8850) );
  NAND2_X1 U10146 ( .A1(n8850), .A2(n8684), .ZN(n8677) );
  OAI211_X1 U10147 ( .C1(n8848), .C2(n8784), .A(n8678), .B(n8677), .ZN(
        P2_U3212) );
  XNOR2_X1 U10148 ( .A(n8679), .B(n8681), .ZN(n8859) );
  NAND2_X1 U10149 ( .A1(n8682), .A2(n8681), .ZN(n8683) );
  NAND2_X1 U10150 ( .A1(n8680), .A2(n8683), .ZN(n8854) );
  NAND2_X1 U10151 ( .A1(n8854), .A2(n8684), .ZN(n8690) );
  NAND2_X1 U10152 ( .A1(n8795), .A2(n8856), .ZN(n8687) );
  AOI22_X1 U10153 ( .A1(n8802), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8756), .B2(
        n8685), .ZN(n8686) );
  OAI211_X1 U10154 ( .C1(n8712), .C2(n8869), .A(n8687), .B(n8686), .ZN(n8688)
         );
  AOI21_X1 U10155 ( .B1(n8937), .B2(n8745), .A(n8688), .ZN(n8689) );
  OAI211_X1 U10156 ( .C1(n8859), .C2(n8784), .A(n8690), .B(n8689), .ZN(
        P2_U3213) );
  NAND2_X1 U10157 ( .A1(n8691), .A2(n8700), .ZN(n8692) );
  NAND3_X1 U10158 ( .A1(n8693), .A2(n10005), .A3(n8692), .ZN(n8696) );
  NAND2_X1 U10159 ( .A1(n8694), .A2(n10043), .ZN(n8695) );
  AND2_X1 U10160 ( .A1(n8696), .A2(n8695), .ZN(n8865) );
  AOI22_X1 U10161 ( .A1(n8802), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8756), .B2(
        n8697), .ZN(n8698) );
  OAI21_X1 U10162 ( .B1(n8731), .B2(n8699), .A(n8698), .ZN(n8705) );
  OR2_X1 U10163 ( .A1(n8701), .A2(n8700), .ZN(n8702) );
  NAND2_X1 U10164 ( .A1(n8703), .A2(n8702), .ZN(n8942) );
  NOR2_X1 U10165 ( .A1(n8942), .A2(n8784), .ZN(n8704) );
  AOI211_X1 U10166 ( .C1(n8757), .C2(n8863), .A(n8705), .B(n8704), .ZN(n8706)
         );
  OAI21_X1 U10167 ( .B1(n8802), .B2(n8865), .A(n8706), .ZN(P2_U3214) );
  XNOR2_X1 U10168 ( .A(n8707), .B(n8708), .ZN(n8870) );
  NAND2_X1 U10169 ( .A1(n8795), .A2(n8855), .ZN(n8711) );
  AOI22_X1 U10170 ( .A1(n8802), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8756), .B2(
        n8709), .ZN(n8710) );
  OAI211_X1 U10171 ( .C1(n8712), .C2(n8868), .A(n8711), .B(n8710), .ZN(n8718)
         );
  INV_X1 U10172 ( .A(n8713), .ZN(n8716) );
  OAI21_X1 U10173 ( .B1(n8716), .B2(n8715), .A(n8714), .ZN(n8946) );
  NOR2_X1 U10174 ( .A1(n8946), .A2(n8784), .ZN(n8717) );
  AOI211_X1 U10175 ( .C1(n8757), .C2(n8873), .A(n8718), .B(n8717), .ZN(n8719)
         );
  OAI21_X1 U10176 ( .B1(n8720), .B2(n8870), .A(n8719), .ZN(P2_U3215) );
  INV_X1 U10177 ( .A(n8721), .ZN(n8722) );
  AOI21_X1 U10178 ( .B1(n8725), .B2(n8723), .A(n8722), .ZN(n8950) );
  XNOR2_X1 U10179 ( .A(n8724), .B(n8725), .ZN(n8727) );
  OAI22_X1 U10180 ( .A1(n8727), .A2(n9979), .B1(n8726), .B2(n10027), .ZN(n8879) );
  NAND2_X1 U10181 ( .A1(n8879), .A2(n8728), .ZN(n8735) );
  AOI22_X1 U10182 ( .A1(n8802), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8756), .B2(
        n8729), .ZN(n8730) );
  OAI21_X1 U10183 ( .B1(n8731), .B2(n8876), .A(n8730), .ZN(n8732) );
  AOI21_X1 U10184 ( .B1(n8733), .B2(n8745), .A(n8732), .ZN(n8734) );
  OAI211_X1 U10185 ( .C1(n8950), .C2(n8784), .A(n8735), .B(n8734), .ZN(
        P2_U3216) );
  XOR2_X1 U10186 ( .A(n8736), .B(n8737), .Z(n8955) );
  XNOR2_X1 U10187 ( .A(n8738), .B(n7704), .ZN(n8739) );
  NAND2_X1 U10188 ( .A1(n8739), .A2(n10005), .ZN(n8742) );
  AOI22_X1 U10189 ( .A1(n10043), .A2(n8764), .B1(n8740), .B2(n10042), .ZN(
        n8741) );
  MUX2_X1 U10190 ( .A(n8743), .B(n8951), .S(n8728), .Z(n8747) );
  AOI22_X1 U10191 ( .A1(n5741), .A2(n8745), .B1(n8756), .B2(n8744), .ZN(n8746)
         );
  OAI211_X1 U10192 ( .C1(n8955), .C2(n8784), .A(n8747), .B(n8746), .ZN(
        P2_U3217) );
  XNOR2_X1 U10193 ( .A(n8749), .B(n8748), .ZN(n8961) );
  XNOR2_X1 U10194 ( .A(n8751), .B(n8750), .ZN(n8753) );
  AOI222_X1 U10195 ( .A1(n10005), .A2(n8753), .B1(n8752), .B2(n10042), .C1(
        n8774), .C2(n10043), .ZN(n8956) );
  MUX2_X1 U10196 ( .A(n8476), .B(n8956), .S(n8728), .Z(n8759) );
  INV_X1 U10197 ( .A(n8754), .ZN(n8755) );
  AOI22_X1 U10198 ( .A1(n8958), .A2(n8757), .B1(n8756), .B2(n8755), .ZN(n8758)
         );
  OAI211_X1 U10199 ( .C1(n8961), .C2(n8784), .A(n8759), .B(n8758), .ZN(
        P2_U3218) );
  XNOR2_X1 U10200 ( .A(n4510), .B(n8762), .ZN(n8967) );
  XNOR2_X1 U10201 ( .A(n8761), .B(n8762), .ZN(n8765) );
  AOI222_X1 U10202 ( .A1(n10005), .A2(n8765), .B1(n8764), .B2(n10042), .C1(
        n8763), .C2(n10043), .ZN(n8962) );
  INV_X1 U10203 ( .A(n8962), .ZN(n8768) );
  OAI22_X1 U10204 ( .A1(n5021), .A2(n8778), .B1(n8766), .B2(n8788), .ZN(n8767)
         );
  OAI21_X1 U10205 ( .B1(n8768), .B2(n8767), .A(n8728), .ZN(n8770) );
  NAND2_X1 U10206 ( .A1(n8802), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8769) );
  OAI211_X1 U10207 ( .C1(n8967), .C2(n8784), .A(n8770), .B(n8769), .ZN(
        P2_U3219) );
  XNOR2_X1 U10208 ( .A(n8771), .B(n8773), .ZN(n8975) );
  XNOR2_X1 U10209 ( .A(n8772), .B(n8773), .ZN(n8776) );
  AOI222_X1 U10210 ( .A1(n10005), .A2(n8776), .B1(n8775), .B2(n10043), .C1(
        n8774), .C2(n10042), .ZN(n8968) );
  INV_X1 U10211 ( .A(n8968), .ZN(n8781) );
  OAI22_X1 U10212 ( .A1(n8779), .A2(n8778), .B1(n8777), .B2(n8788), .ZN(n8780)
         );
  OAI21_X1 U10213 ( .B1(n8781), .B2(n8780), .A(n8728), .ZN(n8783) );
  NAND2_X1 U10214 ( .A1(n8802), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8782) );
  OAI211_X1 U10215 ( .C1(n8975), .C2(n8784), .A(n8783), .B(n8782), .ZN(
        P2_U3220) );
  INV_X1 U10216 ( .A(n8785), .ZN(n8786) );
  AOI21_X1 U10217 ( .B1(n8787), .B2(n8799), .A(n8786), .ZN(n9983) );
  INV_X1 U10218 ( .A(n9983), .ZN(n8794) );
  OAI22_X1 U10219 ( .A1(n8791), .A2(n8790), .B1(n8789), .B2(n8788), .ZN(n8792)
         );
  AOI21_X1 U10220 ( .B1(n8794), .B2(n8793), .A(n8792), .ZN(n8806) );
  AOI22_X1 U10221 ( .A1(n8797), .A2(n8796), .B1(n8795), .B2(n9998), .ZN(n8805)
         );
  OAI21_X1 U10222 ( .B1(n8800), .B2(n8799), .A(n8798), .ZN(n8801) );
  NAND2_X1 U10223 ( .A1(n8801), .A2(n10005), .ZN(n9985) );
  MUX2_X1 U10224 ( .A(n9985), .B(n8803), .S(n8802), .Z(n8804) );
  NAND3_X1 U10225 ( .A1(n8806), .A2(n8805), .A3(n8804), .ZN(P2_U3232) );
  NOR2_X1 U10226 ( .A1(n8807), .A2(n10085), .ZN(n8810) );
  AOI21_X1 U10227 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n10085), .A(n8810), .ZN(
        n8808) );
  OAI21_X1 U10228 ( .B1(n7582), .B2(n8853), .A(n8808), .ZN(P2_U3490) );
  NAND2_X1 U10229 ( .A1(n7581), .A2(n8890), .ZN(n8812) );
  INV_X1 U10230 ( .A(n8810), .ZN(n8811) );
  OAI211_X1 U10231 ( .C1(n10087), .C2(n5769), .A(n8812), .B(n8811), .ZN(
        P2_U3489) );
  INV_X1 U10232 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8813) );
  MUX2_X1 U10233 ( .A(n8897), .B(n8813), .S(n10085), .Z(n8815) );
  NAND2_X1 U10234 ( .A1(n8898), .A2(n8890), .ZN(n8814) );
  OAI211_X1 U10235 ( .C1(n8901), .C2(n8893), .A(n8815), .B(n8814), .ZN(
        P2_U3487) );
  INV_X1 U10236 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8821) );
  OAI22_X1 U10237 ( .A1(n8816), .A2(n10025), .B1(n8827), .B2(n10027), .ZN(
        n8819) );
  NOR2_X1 U10238 ( .A1(n8817), .A2(n10064), .ZN(n8818) );
  AOI211_X1 U10239 ( .C1(n10005), .C2(n8820), .A(n8819), .B(n8818), .ZN(n8902)
         );
  MUX2_X1 U10240 ( .A(n8821), .B(n8902), .S(n10087), .Z(n8822) );
  OAI21_X1 U10241 ( .B1(n4801), .B2(n8853), .A(n8822), .ZN(P2_U3486) );
  INV_X1 U10242 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8823) );
  MUX2_X1 U10243 ( .A(n8823), .B(n8905), .S(n10087), .Z(n8825) );
  NAND2_X1 U10244 ( .A1(n8907), .A2(n8890), .ZN(n8824) );
  OAI211_X1 U10245 ( .C1(n8910), .C2(n8893), .A(n8825), .B(n8824), .ZN(
        P2_U3485) );
  INV_X1 U10246 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8831) );
  OAI22_X1 U10247 ( .A1(n8827), .A2(n10025), .B1(n8826), .B2(n10027), .ZN(
        n8829) );
  AOI211_X1 U10248 ( .C1(n10060), .C2(n8830), .A(n8829), .B(n8828), .ZN(n8911)
         );
  MUX2_X1 U10249 ( .A(n8831), .B(n8911), .S(n10087), .Z(n8832) );
  OAI21_X1 U10250 ( .B1(n8914), .B2(n8893), .A(n8832), .ZN(P2_U3484) );
  MUX2_X1 U10251 ( .A(n8915), .B(P2_REG1_REG_24__SCAN_IN), .S(n10085), .Z(
        n8834) );
  OAI22_X1 U10252 ( .A1(n8917), .A2(n8893), .B1(n8916), .B2(n8853), .ZN(n8833)
         );
  OR2_X1 U10253 ( .A1(n8834), .A2(n8833), .ZN(P2_U3483) );
  INV_X1 U10254 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8835) );
  MUX2_X1 U10255 ( .A(n8835), .B(n8920), .S(n10087), .Z(n8837) );
  NAND2_X1 U10256 ( .A1(n8922), .A2(n8890), .ZN(n8836) );
  OAI211_X1 U10257 ( .C1(n8925), .C2(n8893), .A(n8837), .B(n8836), .ZN(
        P2_U3482) );
  INV_X1 U10258 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8843) );
  AOI22_X1 U10259 ( .A1(n8838), .A2(n10042), .B1(n10043), .B2(n8856), .ZN(
        n8839) );
  OAI21_X1 U10260 ( .B1(n8840), .B2(n10064), .A(n8839), .ZN(n8841) );
  AOI21_X1 U10261 ( .B1(n10005), .B2(n8842), .A(n8841), .ZN(n8926) );
  MUX2_X1 U10262 ( .A(n8843), .B(n8926), .S(n10087), .Z(n8844) );
  OAI21_X1 U10263 ( .B1(n8929), .B2(n8853), .A(n8844), .ZN(P2_U3481) );
  INV_X1 U10264 ( .A(n8845), .ZN(n8934) );
  INV_X1 U10265 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8851) );
  AOI22_X1 U10266 ( .A1(n8846), .A2(n10042), .B1(n10043), .B2(n8862), .ZN(
        n8847) );
  OAI21_X1 U10267 ( .B1(n8848), .B2(n10064), .A(n8847), .ZN(n8849) );
  AOI21_X1 U10268 ( .B1(n10005), .B2(n8850), .A(n8849), .ZN(n8930) );
  MUX2_X1 U10269 ( .A(n8851), .B(n8930), .S(n10087), .Z(n8852) );
  OAI21_X1 U10270 ( .B1(n8934), .B2(n8853), .A(n8852), .ZN(P2_U3480) );
  NAND2_X1 U10271 ( .A1(n8854), .A2(n10005), .ZN(n8858) );
  AOI22_X1 U10272 ( .A1(n8856), .A2(n10042), .B1(n10043), .B2(n8855), .ZN(
        n8857) );
  OAI211_X1 U10273 ( .C1(n10064), .C2(n8859), .A(n8858), .B(n8857), .ZN(n8935)
         );
  MUX2_X1 U10274 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8935), .S(n10087), .Z(
        n8860) );
  AOI21_X1 U10275 ( .B1(n8890), .B2(n8937), .A(n8860), .ZN(n8861) );
  INV_X1 U10276 ( .A(n8861), .ZN(P2_U3479) );
  AOI22_X1 U10277 ( .A1(n8863), .A2(n10060), .B1(n10042), .B2(n8862), .ZN(
        n8864) );
  NAND2_X1 U10278 ( .A1(n8865), .A2(n8864), .ZN(n8939) );
  MUX2_X1 U10279 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8939), .S(n10087), .Z(
        n8866) );
  INV_X1 U10280 ( .A(n8866), .ZN(n8867) );
  OAI21_X1 U10281 ( .B1(n8893), .B2(n8942), .A(n8867), .ZN(P2_U3478) );
  INV_X1 U10282 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8874) );
  OAI22_X1 U10283 ( .A1(n8869), .A2(n10025), .B1(n8868), .B2(n10027), .ZN(
        n8872) );
  NOR2_X1 U10284 ( .A1(n8870), .A2(n9979), .ZN(n8871) );
  AOI211_X1 U10285 ( .C1(n10060), .C2(n8873), .A(n8872), .B(n8871), .ZN(n8943)
         );
  MUX2_X1 U10286 ( .A(n8874), .B(n8943), .S(n10087), .Z(n8875) );
  OAI21_X1 U10287 ( .B1(n8893), .B2(n8946), .A(n8875), .ZN(P2_U3477) );
  OAI22_X1 U10288 ( .A1(n8877), .A2(n10062), .B1(n8876), .B2(n10025), .ZN(
        n8878) );
  NOR2_X1 U10289 ( .A1(n8879), .A2(n8878), .ZN(n8947) );
  MUX2_X1 U10290 ( .A(n9960), .B(n8947), .S(n10087), .Z(n8880) );
  OAI21_X1 U10291 ( .B1(n8950), .B2(n8893), .A(n8880), .ZN(P2_U3476) );
  MUX2_X1 U10292 ( .A(n8881), .B(n8951), .S(n10087), .Z(n8883) );
  NAND2_X1 U10293 ( .A1(n5741), .A2(n8890), .ZN(n8882) );
  OAI211_X1 U10294 ( .C1(n8955), .C2(n8893), .A(n8883), .B(n8882), .ZN(
        P2_U3475) );
  MUX2_X1 U10295 ( .A(n8884), .B(n8956), .S(n10087), .Z(n8886) );
  NAND2_X1 U10296 ( .A1(n8958), .A2(n8890), .ZN(n8885) );
  OAI211_X1 U10297 ( .C1(n8961), .C2(n8893), .A(n8886), .B(n8885), .ZN(
        P2_U3474) );
  MUX2_X1 U10298 ( .A(n8887), .B(n8962), .S(n10087), .Z(n8889) );
  NAND2_X1 U10299 ( .A1(n8964), .A2(n8890), .ZN(n8888) );
  OAI211_X1 U10300 ( .C1(n8967), .C2(n8893), .A(n8889), .B(n8888), .ZN(
        P2_U3473) );
  MUX2_X1 U10301 ( .A(n9908), .B(n8968), .S(n10087), .Z(n8892) );
  NAND2_X1 U10302 ( .A1(n8971), .A2(n8890), .ZN(n8891) );
  OAI211_X1 U10303 ( .C1(n8893), .C2(n8975), .A(n8892), .B(n8891), .ZN(
        P2_U3472) );
  AOI21_X1 U10304 ( .B1(n10070), .B2(P2_REG0_REG_31__SCAN_IN), .A(n8894), .ZN(
        n8895) );
  OAI21_X1 U10305 ( .B1(n7582), .B2(n8933), .A(n8895), .ZN(P2_U3458) );
  INV_X1 U10306 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8896) );
  MUX2_X1 U10307 ( .A(n8897), .B(n8896), .S(n10070), .Z(n8900) );
  NAND2_X1 U10308 ( .A1(n8898), .A2(n8970), .ZN(n8899) );
  OAI211_X1 U10309 ( .C1(n8901), .C2(n8974), .A(n8900), .B(n8899), .ZN(
        P2_U3455) );
  INV_X1 U10310 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8903) );
  MUX2_X1 U10311 ( .A(n8903), .B(n8902), .S(n10068), .Z(n8904) );
  OAI21_X1 U10312 ( .B1(n4801), .B2(n8933), .A(n8904), .ZN(P2_U3454) );
  INV_X1 U10313 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8906) );
  MUX2_X1 U10314 ( .A(n8906), .B(n8905), .S(n10068), .Z(n8909) );
  NAND2_X1 U10315 ( .A1(n8907), .A2(n8970), .ZN(n8908) );
  OAI211_X1 U10316 ( .C1(n8910), .C2(n8974), .A(n8909), .B(n8908), .ZN(
        P2_U3453) );
  INV_X1 U10317 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8912) );
  MUX2_X1 U10318 ( .A(n8912), .B(n8911), .S(n10068), .Z(n8913) );
  OAI21_X1 U10319 ( .B1(n8914), .B2(n8974), .A(n8913), .ZN(P2_U3452) );
  MUX2_X1 U10320 ( .A(n8915), .B(P2_REG0_REG_24__SCAN_IN), .S(n10070), .Z(
        n8919) );
  OAI22_X1 U10321 ( .A1(n8917), .A2(n8974), .B1(n8916), .B2(n8933), .ZN(n8918)
         );
  OR2_X1 U10322 ( .A1(n8919), .A2(n8918), .ZN(P2_U3451) );
  INV_X1 U10323 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8921) );
  MUX2_X1 U10324 ( .A(n8921), .B(n8920), .S(n10068), .Z(n8924) );
  NAND2_X1 U10325 ( .A1(n8922), .A2(n8970), .ZN(n8923) );
  OAI211_X1 U10326 ( .C1(n8925), .C2(n8974), .A(n8924), .B(n8923), .ZN(
        P2_U3450) );
  INV_X1 U10327 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8927) );
  MUX2_X1 U10328 ( .A(n8927), .B(n8926), .S(n10068), .Z(n8928) );
  OAI21_X1 U10329 ( .B1(n8929), .B2(n8933), .A(n8928), .ZN(P2_U3449) );
  INV_X1 U10330 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8931) );
  MUX2_X1 U10331 ( .A(n8931), .B(n8930), .S(n10068), .Z(n8932) );
  OAI21_X1 U10332 ( .B1(n8934), .B2(n8933), .A(n8932), .ZN(P2_U3448) );
  MUX2_X1 U10333 ( .A(n8935), .B(P2_REG0_REG_20__SCAN_IN), .S(n10070), .Z(
        n8936) );
  AOI21_X1 U10334 ( .B1(n8970), .B2(n8937), .A(n8936), .ZN(n8938) );
  INV_X1 U10335 ( .A(n8938), .ZN(P2_U3447) );
  MUX2_X1 U10336 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8939), .S(n10068), .Z(
        n8940) );
  INV_X1 U10337 ( .A(n8940), .ZN(n8941) );
  OAI21_X1 U10338 ( .B1(n8942), .B2(n8974), .A(n8941), .ZN(P2_U3446) );
  INV_X1 U10339 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8944) );
  MUX2_X1 U10340 ( .A(n8944), .B(n8943), .S(n10068), .Z(n8945) );
  OAI21_X1 U10341 ( .B1(n8946), .B2(n8974), .A(n8945), .ZN(P2_U3444) );
  MUX2_X1 U10342 ( .A(n8948), .B(n8947), .S(n10068), .Z(n8949) );
  OAI21_X1 U10343 ( .B1(n8950), .B2(n8974), .A(n8949), .ZN(P2_U3441) );
  MUX2_X1 U10344 ( .A(n8952), .B(n8951), .S(n10068), .Z(n8954) );
  NAND2_X1 U10345 ( .A1(n5741), .A2(n8970), .ZN(n8953) );
  OAI211_X1 U10346 ( .C1(n8955), .C2(n8974), .A(n8954), .B(n8953), .ZN(
        P2_U3438) );
  INV_X1 U10347 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8957) );
  MUX2_X1 U10348 ( .A(n8957), .B(n8956), .S(n10068), .Z(n8960) );
  NAND2_X1 U10349 ( .A1(n8958), .A2(n8970), .ZN(n8959) );
  OAI211_X1 U10350 ( .C1(n8961), .C2(n8974), .A(n8960), .B(n8959), .ZN(
        P2_U3435) );
  INV_X1 U10351 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8963) );
  MUX2_X1 U10352 ( .A(n8963), .B(n8962), .S(n10068), .Z(n8966) );
  NAND2_X1 U10353 ( .A1(n8964), .A2(n8970), .ZN(n8965) );
  OAI211_X1 U10354 ( .C1(n8967), .C2(n8974), .A(n8966), .B(n8965), .ZN(
        P2_U3432) );
  INV_X1 U10355 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8969) );
  MUX2_X1 U10356 ( .A(n8969), .B(n8968), .S(n10068), .Z(n8973) );
  NAND2_X1 U10357 ( .A1(n8971), .A2(n8970), .ZN(n8972) );
  OAI211_X1 U10358 ( .C1(n8975), .C2(n8974), .A(n8973), .B(n8972), .ZN(
        P2_U3429) );
  NAND3_X1 U10359 ( .A1(n8977), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n8978) );
  OAI22_X1 U10360 ( .A1(n8979), .A2(n8978), .B1(n6128), .B2(n8991), .ZN(n8980)
         );
  AOI21_X1 U10361 ( .B1(n8976), .B2(n8981), .A(n8980), .ZN(n8982) );
  INV_X1 U10362 ( .A(n8982), .ZN(P2_U3264) );
  AOI21_X1 U10363 ( .B1(n8988), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8983), .ZN(
        n8984) );
  OAI21_X1 U10364 ( .B1(n8985), .B2(n8990), .A(n8984), .ZN(P2_U3267) );
  INV_X1 U10365 ( .A(n8986), .ZN(n9792) );
  AOI21_X1 U10366 ( .B1(n8988), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n8987), .ZN(
        n8989) );
  OAI21_X1 U10367 ( .B1(n9792), .B2(n8990), .A(n8989), .ZN(P2_U3268) );
  OAI222_X1 U10368 ( .A1(n8990), .A2(n8994), .B1(P2_U3151), .B2(n8993), .C1(
        n8992), .C2(n8991), .ZN(P2_U3269) );
  INV_X1 U10369 ( .A(n8995), .ZN(n8996) );
  MUX2_X1 U10370 ( .A(n8996), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  NAND2_X1 U10371 ( .A1(n8998), .A2(n8997), .ZN(n9000) );
  XNOR2_X1 U10372 ( .A(n9000), .B(n8999), .ZN(n9005) );
  OAI21_X1 U10373 ( .B1(n9157), .B2(n9558), .A(n9001), .ZN(n9003) );
  OAI22_X1 U10374 ( .A1(n9562), .A2(n9159), .B1(n9158), .B2(n9525), .ZN(n9002)
         );
  AOI211_X1 U10375 ( .C1(n9568), .C2(n9162), .A(n9003), .B(n9002), .ZN(n9004)
         );
  OAI21_X1 U10376 ( .B1(n9005), .B2(n9164), .A(n9004), .ZN(P1_U3215) );
  AND2_X1 U10377 ( .A1(n9128), .A2(n9006), .ZN(n9008) );
  OAI211_X1 U10378 ( .C1(n9008), .C2(n9007), .A(n9143), .B(n9098), .ZN(n9012)
         );
  NOR2_X1 U10379 ( .A1(n9157), .A2(n9403), .ZN(n9010) );
  OAI22_X1 U10380 ( .A1(n9405), .A2(n9159), .B1(n9158), .B2(n9374), .ZN(n9009)
         );
  AOI211_X1 U10381 ( .C1(P1_REG3_REG_23__SCAN_IN), .C2(P1_U3086), .A(n9010), 
        .B(n9009), .ZN(n9011) );
  OAI211_X1 U10382 ( .C1(n9652), .C2(n9126), .A(n9012), .B(n9011), .ZN(
        P1_U3216) );
  OAI21_X1 U10383 ( .B1(n9014), .B2(n9013), .A(n6565), .ZN(n9015) );
  NAND2_X1 U10384 ( .A1(n9015), .A2(n9143), .ZN(n9022) );
  AOI22_X1 U10385 ( .A1(n9072), .A2(n9173), .B1(n9016), .B2(n9162), .ZN(n9021)
         );
  INV_X1 U10386 ( .A(n9017), .ZN(n9019) );
  NOR2_X1 U10387 ( .A1(n9157), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9018) );
  AOI211_X1 U10388 ( .C1(n9077), .C2(n9175), .A(n9019), .B(n9018), .ZN(n9020)
         );
  NAND3_X1 U10389 ( .A1(n9022), .A2(n9021), .A3(n9020), .ZN(P1_U3218) );
  XNOR2_X1 U10390 ( .A(n9024), .B(n9023), .ZN(n9137) );
  NOR2_X1 U10391 ( .A1(n9137), .A2(n9138), .ZN(n9136) );
  NOR2_X1 U10392 ( .A1(n9024), .A2(n9023), .ZN(n9028) );
  XNOR2_X1 U10393 ( .A(n9026), .B(n9025), .ZN(n9027) );
  NOR3_X1 U10394 ( .A1(n9136), .A2(n9028), .A3(n9027), .ZN(n9107) );
  INV_X1 U10395 ( .A(n9107), .ZN(n9030) );
  OAI21_X1 U10396 ( .B1(n9136), .B2(n9028), .A(n9027), .ZN(n9029) );
  NAND3_X1 U10397 ( .A1(n9030), .A2(n9143), .A3(n9029), .ZN(n9034) );
  INV_X1 U10398 ( .A(n9031), .ZN(n9469) );
  AND2_X1 U10399 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9260) );
  OAI22_X1 U10400 ( .A1(n9277), .A2(n9159), .B1(n9158), .B2(n9437), .ZN(n9032)
         );
  AOI211_X1 U10401 ( .C1(n9123), .C2(n9469), .A(n9260), .B(n9032), .ZN(n9033)
         );
  OAI211_X1 U10402 ( .C1(n4711), .C2(n9126), .A(n9034), .B(n9033), .ZN(
        P1_U3219) );
  XOR2_X1 U10403 ( .A(n9036), .B(n9035), .Z(n9041) );
  OAI22_X1 U10404 ( .A1(n9157), .A2(n9435), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9037), .ZN(n9039) );
  OAI22_X1 U10405 ( .A1(n9437), .A2(n9159), .B1(n9158), .B2(n9405), .ZN(n9038)
         );
  AOI211_X1 U10406 ( .C1(n9431), .C2(n9162), .A(n9039), .B(n9038), .ZN(n9040)
         );
  OAI21_X1 U10407 ( .B1(n9041), .B2(n9164), .A(n9040), .ZN(P1_U3223) );
  OAI21_X1 U10408 ( .B1(n9043), .B2(n4527), .A(n9042), .ZN(n9044) );
  NAND2_X1 U10409 ( .A1(n9044), .A2(n9143), .ZN(n9051) );
  INV_X1 U10410 ( .A(n9045), .ZN(n9049) );
  OAI22_X1 U10411 ( .A1(n9046), .A2(n9159), .B1(n9158), .B2(n9562), .ZN(n9047)
         );
  AOI211_X1 U10412 ( .C1(n9123), .C2(n9049), .A(n9048), .B(n9047), .ZN(n9050)
         );
  OAI211_X1 U10413 ( .C1(n9832), .C2(n9126), .A(n9051), .B(n9050), .ZN(
        P1_U3224) );
  OAI21_X1 U10414 ( .B1(n9054), .B2(n9053), .A(n9052), .ZN(n9055) );
  NAND2_X1 U10415 ( .A1(n9055), .A2(n9143), .ZN(n9059) );
  NOR2_X1 U10416 ( .A1(n9157), .A2(n9370), .ZN(n9057) );
  OAI22_X1 U10417 ( .A1(n9374), .A2(n9159), .B1(n9158), .B2(n9341), .ZN(n9056)
         );
  AOI211_X1 U10418 ( .C1(P1_REG3_REG_25__SCAN_IN), .C2(P1_U3086), .A(n9057), 
        .B(n9056), .ZN(n9058) );
  OAI211_X1 U10419 ( .C1(n9639), .C2(n9126), .A(n9059), .B(n9058), .ZN(
        P1_U3225) );
  NOR2_X1 U10420 ( .A1(n4868), .A2(n9061), .ZN(n9062) );
  XNOR2_X1 U10421 ( .A(n9063), .B(n9062), .ZN(n9067) );
  NAND2_X1 U10422 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9198) );
  OAI21_X1 U10423 ( .B1(n9157), .B2(n9523), .A(n9198), .ZN(n9065) );
  OAI22_X1 U10424 ( .A1(n9525), .A2(n9159), .B1(n9158), .B2(n9685), .ZN(n9064)
         );
  AOI211_X1 U10425 ( .C1(n9528), .C2(n9162), .A(n9065), .B(n9064), .ZN(n9066)
         );
  OAI21_X1 U10426 ( .B1(n9067), .B2(n9164), .A(n9066), .ZN(P1_U3226) );
  OAI21_X1 U10427 ( .B1(n9069), .B2(n4600), .A(n9068), .ZN(n9070) );
  NAND2_X1 U10428 ( .A1(n9070), .A2(n9143), .ZN(n9080) );
  AOI22_X1 U10429 ( .A1(n9072), .A2(n9171), .B1(n9071), .B2(n9162), .ZN(n9079)
         );
  INV_X1 U10430 ( .A(n9073), .ZN(n9076) );
  NOR2_X1 U10431 ( .A1(n9157), .A2(n9074), .ZN(n9075) );
  AOI211_X1 U10432 ( .C1(n9077), .C2(n9173), .A(n9076), .B(n9075), .ZN(n9078)
         );
  NAND3_X1 U10433 ( .A1(n9080), .A2(n9079), .A3(n9078), .ZN(P1_U3227) );
  XNOR2_X1 U10434 ( .A(n9083), .B(n9082), .ZN(n9084) );
  XNOR2_X1 U10435 ( .A(n9081), .B(n9084), .ZN(n9094) );
  NAND3_X1 U10436 ( .A1(n9123), .A2(n9085), .A3(n9089), .ZN(n9086) );
  OAI21_X1 U10437 ( .B1(n9159), .B2(n9707), .A(n9086), .ZN(n9092) );
  AOI21_X1 U10438 ( .B1(n9088), .B2(n9087), .A(P1_U3086), .ZN(n9090) );
  OAI22_X1 U10439 ( .A1(n9158), .A2(n9277), .B1(n9090), .B2(n9089), .ZN(n9091)
         );
  AOI211_X1 U10440 ( .C1(n9696), .C2(n9162), .A(n9092), .B(n9091), .ZN(n9093)
         );
  OAI21_X1 U10441 ( .B1(n9094), .B2(n9164), .A(n9093), .ZN(P1_U3228) );
  INV_X1 U10442 ( .A(n9095), .ZN(n9100) );
  AOI21_X1 U10443 ( .B1(n9098), .B2(n9097), .A(n9096), .ZN(n9099) );
  OAI21_X1 U10444 ( .B1(n9100), .B2(n9099), .A(n9143), .ZN(n9105) );
  NOR2_X1 U10445 ( .A1(n9101), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9103) );
  OAI22_X1 U10446 ( .A1(n9285), .A2(n9159), .B1(n9158), .B2(n9626), .ZN(n9102)
         );
  AOI211_X1 U10447 ( .C1(n9123), .C2(n9391), .A(n9103), .B(n9102), .ZN(n9104)
         );
  OAI211_X1 U10448 ( .C1(n9763), .C2(n9126), .A(n9105), .B(n9104), .ZN(
        P1_U3229) );
  NOR2_X1 U10449 ( .A1(n9107), .A2(n9106), .ZN(n9108) );
  XOR2_X1 U10450 ( .A(n9109), .B(n9108), .Z(n9114) );
  OAI22_X1 U10451 ( .A1(n9157), .A2(n9449), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9110), .ZN(n9112) );
  OAI22_X1 U10452 ( .A1(n9686), .A2(n9159), .B1(n9158), .B2(n9280), .ZN(n9111)
         );
  AOI211_X1 U10453 ( .C1(n9676), .C2(n9162), .A(n9112), .B(n9111), .ZN(n9113)
         );
  OAI21_X1 U10454 ( .B1(n9114), .B2(n9164), .A(n9113), .ZN(P1_U3233) );
  OAI21_X1 U10455 ( .B1(n9117), .B2(n9116), .A(n9115), .ZN(n9118) );
  NAND2_X1 U10456 ( .A1(n9118), .A2(n9143), .ZN(n9125) );
  INV_X1 U10457 ( .A(n9119), .ZN(n9584) );
  INV_X1 U10458 ( .A(n9120), .ZN(n9122) );
  OAI22_X1 U10459 ( .A1(n9580), .A2(n9159), .B1(n9158), .B2(n9732), .ZN(n9121)
         );
  AOI211_X1 U10460 ( .C1(n9123), .C2(n9584), .A(n9122), .B(n9121), .ZN(n9124)
         );
  OAI211_X1 U10461 ( .C1(n9779), .C2(n9126), .A(n9125), .B(n9124), .ZN(
        P1_U3234) );
  NAND2_X1 U10462 ( .A1(n9128), .A2(n9127), .ZN(n9130) );
  XNOR2_X1 U10463 ( .A(n9130), .B(n9129), .ZN(n9135) );
  OAI22_X1 U10464 ( .A1(n9157), .A2(n9418), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9131), .ZN(n9133) );
  OAI22_X1 U10465 ( .A1(n9280), .A2(n9159), .B1(n9158), .B2(n9285), .ZN(n9132)
         );
  AOI211_X1 U10466 ( .C1(n9422), .C2(n9162), .A(n9133), .B(n9132), .ZN(n9134)
         );
  OAI21_X1 U10467 ( .B1(n9135), .B2(n9164), .A(n9134), .ZN(P1_U3235) );
  AOI21_X1 U10468 ( .B1(n9138), .B2(n9137), .A(n9136), .ZN(n9142) );
  NAND2_X1 U10469 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9233) );
  OAI21_X1 U10470 ( .B1(n9157), .B2(n9481), .A(n9233), .ZN(n9140) );
  OAI22_X1 U10471 ( .A1(n9685), .A2(n9159), .B1(n9158), .B2(n9686), .ZN(n9139)
         );
  AOI211_X1 U10472 ( .C1(n9689), .C2(n9162), .A(n9140), .B(n9139), .ZN(n9141)
         );
  OAI21_X1 U10473 ( .B1(n9142), .B2(n9164), .A(n9141), .ZN(P1_U3238) );
  NAND2_X1 U10474 ( .A1(n4872), .A2(n9143), .ZN(n9151) );
  AOI21_X1 U10475 ( .B1(n9052), .B2(n9145), .A(n9144), .ZN(n9150) );
  OAI22_X1 U10476 ( .A1(n9157), .A2(n9356), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9146), .ZN(n9148) );
  OAI22_X1 U10477 ( .A1(n9627), .A2(n9158), .B1(n9159), .B2(n9626), .ZN(n9147)
         );
  AOI211_X1 U10478 ( .C1(n9355), .C2(n9162), .A(n9148), .B(n9147), .ZN(n9149)
         );
  OAI21_X1 U10479 ( .B1(n9151), .B2(n9150), .A(n9149), .ZN(P1_U3240) );
  NAND2_X1 U10480 ( .A1(n9153), .A2(n9152), .ZN(n9154) );
  XOR2_X1 U10481 ( .A(n9155), .B(n9154), .Z(n9165) );
  NAND2_X1 U10482 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9183) );
  OAI21_X1 U10483 ( .B1(n9157), .B2(n9539), .A(n9183), .ZN(n9161) );
  OAI22_X1 U10484 ( .A1(n9732), .A2(n9159), .B1(n9158), .B2(n9707), .ZN(n9160)
         );
  AOI211_X1 U10485 ( .C1(n9711), .C2(n9162), .A(n9161), .B(n9160), .ZN(n9163)
         );
  OAI21_X1 U10486 ( .B1(n9165), .B2(n9164), .A(n9163), .ZN(P1_U3241) );
  MUX2_X1 U10487 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9360), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10488 ( .A(n9636), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9176), .Z(
        P1_U3580) );
  MUX2_X1 U10489 ( .A(n9386), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9176), .Z(
        P1_U3579) );
  MUX2_X1 U10490 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9649), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10491 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9667), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10492 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9657), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10493 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9485), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10494 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9505), .S(P1_U3973), .Z(
        P1_U3572) );
  INV_X1 U10495 ( .A(n9685), .ZN(n9699) );
  MUX2_X1 U10496 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9699), .S(P1_U3973), .Z(
        P1_U3571) );
  INV_X1 U10497 ( .A(n9707), .ZN(n9543) );
  MUX2_X1 U10498 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9543), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10499 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9719), .S(P1_U3973), .Z(
        P1_U3569) );
  INV_X1 U10500 ( .A(n9732), .ZN(n9586) );
  MUX2_X1 U10501 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9586), .S(P1_U3973), .Z(
        P1_U3568) );
  INV_X1 U10502 ( .A(n9562), .ZN(n9722) );
  MUX2_X1 U10503 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9722), .S(P1_U3973), .Z(
        P1_U3567) );
  INV_X1 U10504 ( .A(n9580), .ZN(n9269) );
  MUX2_X1 U10505 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9269), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10506 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9166), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10507 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9167), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10508 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9168), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10509 ( .A(n9169), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9176), .Z(
        P1_U3562) );
  MUX2_X1 U10510 ( .A(n9170), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9176), .Z(
        P1_U3561) );
  MUX2_X1 U10511 ( .A(n9171), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9176), .Z(
        P1_U3560) );
  MUX2_X1 U10512 ( .A(n9172), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9176), .Z(
        P1_U3559) );
  MUX2_X1 U10513 ( .A(n9173), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9176), .Z(
        P1_U3558) );
  MUX2_X1 U10514 ( .A(n9174), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9176), .Z(
        P1_U3557) );
  MUX2_X1 U10515 ( .A(n9175), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9176), .Z(
        P1_U3556) );
  MUX2_X1 U10516 ( .A(n9177), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9176), .Z(
        P1_U3555) );
  MUX2_X1 U10517 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9178), .S(P1_U3973), .Z(
        P1_U3554) );
  NOR2_X1 U10518 ( .A1(n9180), .A2(n9181), .ZN(n9193) );
  AOI211_X1 U10519 ( .C1(n9181), .C2(n9180), .A(n9193), .B(n9254), .ZN(n9191)
         );
  INV_X1 U10520 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9185) );
  NAND2_X1 U10521 ( .A1(n9236), .A2(n9182), .ZN(n9184) );
  OAI211_X1 U10522 ( .C1(n9185), .C2(n9234), .A(n9184), .B(n9183), .ZN(n9190)
         );
  NOR2_X1 U10523 ( .A1(n9540), .A2(n9188), .ZN(n9203) );
  AOI211_X1 U10524 ( .C1(n9188), .C2(n9540), .A(n9203), .B(n9259), .ZN(n9189)
         );
  OR3_X1 U10525 ( .A1(n9191), .A2(n9190), .A3(n9189), .ZN(P1_U3258) );
  NOR2_X1 U10526 ( .A1(n9192), .A2(n9201), .ZN(n9194) );
  XNOR2_X1 U10527 ( .A(n9217), .B(n9195), .ZN(n9196) );
  OAI21_X1 U10528 ( .B1(n9197), .B2(n9196), .A(n9216), .ZN(n9210) );
  INV_X1 U10529 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9200) );
  NAND2_X1 U10530 ( .A1(n9236), .A2(n9217), .ZN(n9199) );
  OAI211_X1 U10531 ( .C1(n9200), .C2(n9234), .A(n9199), .B(n9198), .ZN(n9209)
         );
  NOR2_X1 U10532 ( .A1(n9202), .A2(n9201), .ZN(n9204) );
  NOR2_X1 U10533 ( .A1(n9204), .A2(n9203), .ZN(n9207) );
  NAND2_X1 U10534 ( .A1(n9217), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9205) );
  OAI21_X1 U10535 ( .B1(n9217), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9205), .ZN(
        n9206) );
  NOR2_X1 U10536 ( .A1(n9207), .A2(n9206), .ZN(n9212) );
  AOI211_X1 U10537 ( .C1(n9207), .C2(n9206), .A(n9212), .B(n9259), .ZN(n9208)
         );
  AOI211_X1 U10538 ( .C1(n9255), .C2(n9210), .A(n9209), .B(n9208), .ZN(n9211)
         );
  INV_X1 U10539 ( .A(n9211), .ZN(P1_U3259) );
  NOR2_X1 U10540 ( .A1(n9215), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9226) );
  AOI21_X1 U10541 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n9215), .A(n9226), .ZN(
        n9214) );
  OAI21_X1 U10542 ( .B1(n9214), .B2(n9213), .A(n9228), .ZN(n9224) );
  AOI22_X1 U10543 ( .A1(n9215), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n9237), .B2(
        n9238), .ZN(n9219) );
  OAI21_X1 U10544 ( .B1(n9219), .B2(n9218), .A(n9240), .ZN(n9220) );
  NAND2_X1 U10545 ( .A1(n9220), .A2(n9255), .ZN(n9222) );
  AOI22_X1 U10546 ( .A1(n9261), .A2(P1_ADDR_REG_17__SCAN_IN), .B1(
        P1_REG3_REG_17__SCAN_IN), .B2(P1_U3086), .ZN(n9221) );
  OAI211_X1 U10547 ( .C1(n9258), .C2(n9238), .A(n9222), .B(n9221), .ZN(n9223)
         );
  AOI21_X1 U10548 ( .B1(n9230), .B2(n9224), .A(n9223), .ZN(n9225) );
  INV_X1 U10549 ( .A(n9225), .ZN(P1_U3260) );
  INV_X1 U10550 ( .A(n9226), .ZN(n9227) );
  OR2_X1 U10551 ( .A1(n9241), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9229) );
  NAND2_X1 U10552 ( .A1(n9241), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9248) );
  AND2_X1 U10553 ( .A1(n9229), .A2(n9248), .ZN(n9231) );
  OAI211_X1 U10554 ( .C1(n9232), .C2(n9231), .A(n9249), .B(n9230), .ZN(n9247)
         );
  INV_X1 U10555 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10111) );
  OAI21_X1 U10556 ( .B1(n9234), .B2(n10111), .A(n9233), .ZN(n9235) );
  AOI21_X1 U10557 ( .B1(n9236), .B2(n9241), .A(n9235), .ZN(n9246) );
  NAND2_X1 U10558 ( .A1(n9238), .A2(n9237), .ZN(n9239) );
  AND2_X1 U10559 ( .A1(n9240), .A2(n9239), .ZN(n9244) );
  OR2_X1 U10560 ( .A1(n9241), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9242) );
  NAND2_X1 U10561 ( .A1(n9241), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9251) );
  AND2_X1 U10562 ( .A1(n9242), .A2(n9251), .ZN(n9243) );
  NAND2_X1 U10563 ( .A1(n9244), .A2(n9243), .ZN(n9252) );
  OAI211_X1 U10564 ( .C1(n9244), .C2(n9243), .A(n9252), .B(n9255), .ZN(n9245)
         );
  NAND3_X1 U10565 ( .A1(n9247), .A2(n9246), .A3(n9245), .ZN(P1_U3261) );
  NAND2_X1 U10566 ( .A1(n9249), .A2(n9248), .ZN(n9250) );
  NAND2_X1 U10567 ( .A1(n9252), .A2(n9251), .ZN(n9253) );
  XNOR2_X1 U10568 ( .A(n9253), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9256) );
  NAND2_X1 U10569 ( .A1(n9256), .A2(n9255), .ZN(n9257) );
  INV_X1 U10570 ( .A(n9293), .ZN(n9264) );
  INV_X1 U10571 ( .A(n9262), .ZN(n9263) );
  AOI211_X1 U10572 ( .C1(n9265), .C2(n9264), .A(n9494), .B(n9263), .ZN(n9603)
         );
  NAND2_X1 U10573 ( .A1(n9603), .A2(n9538), .ZN(n9268) );
  AOI21_X1 U10574 ( .B1(n9585), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9266), .ZN(
        n9267) );
  OAI211_X1 U10575 ( .C1(n9746), .C2(n9590), .A(n9268), .B(n9267), .ZN(
        P1_U3264) );
  NAND2_X1 U10576 ( .A1(n9573), .A2(n9576), .ZN(n9572) );
  AOI21_X1 U10577 ( .B1(n9732), .B2(n9776), .A(n9555), .ZN(n9512) );
  NAND2_X1 U10578 ( .A1(n9711), .A2(n9719), .ZN(n9515) );
  NAND2_X1 U10579 ( .A1(n9568), .A2(n9586), .ZN(n9510) );
  NAND2_X1 U10580 ( .A1(n9515), .A2(n9510), .ZN(n9274) );
  OR2_X1 U10581 ( .A1(n9711), .A2(n9719), .ZN(n9513) );
  OAI211_X1 U10582 ( .C1(n9512), .C2(n9274), .A(n9517), .B(n9513), .ZN(n9516)
         );
  OAI21_X1 U10583 ( .B1(n9707), .B2(n9702), .A(n9516), .ZN(n9493) );
  NAND2_X1 U10584 ( .A1(n9495), .A2(n9685), .ZN(n9276) );
  INV_X1 U10585 ( .A(n9689), .ZN(n9487) );
  OAI21_X1 U10586 ( .B1(n9444), .B2(n5105), .A(n4586), .ZN(n9279) );
  INV_X1 U10587 ( .A(n9279), .ZN(n9428) );
  NAND2_X1 U10588 ( .A1(n9281), .A2(n9280), .ZN(n9282) );
  NAND2_X1 U10589 ( .A1(n9661), .A2(n9405), .ZN(n9283) );
  NOR2_X1 U10590 ( .A1(n9763), .A2(n9374), .ZN(n9286) );
  NAND2_X1 U10591 ( .A1(n9355), .A2(n9636), .ZN(n9287) );
  NAND2_X1 U10592 ( .A1(n9288), .A2(n9287), .ZN(n9345) );
  OAI22_X1 U10593 ( .A1(n9345), .A2(n9344), .B1(n9360), .B2(n9620), .ZN(n9323)
         );
  NAND2_X1 U10594 ( .A1(n9325), .A2(n5108), .ZN(n9290) );
  XNOR2_X1 U10595 ( .A(n9290), .B(n9289), .ZN(n9606) );
  INV_X1 U10596 ( .A(n9606), .ZN(n9316) );
  INV_X1 U10597 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9291) );
  OAI22_X1 U10598 ( .A1(n9607), .A2(n9561), .B1(n9598), .B2(n9291), .ZN(n9292)
         );
  AOI21_X1 U10599 ( .B1(n8101), .B2(n9569), .A(n9292), .ZN(n9315) );
  AOI211_X1 U10600 ( .C1(n8101), .C2(n9326), .A(n9494), .B(n9293), .ZN(n9610)
         );
  INV_X1 U10601 ( .A(n9610), .ZN(n9295) );
  OAI22_X1 U10602 ( .A1(n9295), .A2(n9327), .B1(n9557), .B2(n9294), .ZN(n9313)
         );
  NAND2_X1 U10603 ( .A1(n9455), .A2(n9454), .ZN(n9453) );
  NAND2_X1 U10604 ( .A1(n9299), .A2(n9298), .ZN(n9400) );
  NAND2_X1 U10605 ( .A1(n9400), .A2(n9399), .ZN(n9398) );
  INV_X1 U10606 ( .A(n9381), .ZN(n9300) );
  NOR2_X1 U10607 ( .A1(n9382), .A2(n9300), .ZN(n9301) );
  NAND2_X1 U10608 ( .A1(n9398), .A2(n9301), .ZN(n9384) );
  NAND2_X1 U10609 ( .A1(n9350), .A2(n9305), .ZN(n9338) );
  NAND2_X1 U10610 ( .A1(n9338), .A2(n9344), .ZN(n9337) );
  AND2_X1 U10611 ( .A1(n9337), .A2(n9306), .ZN(n9318) );
  INV_X1 U10612 ( .A(n9322), .ZN(n9317) );
  XNOR2_X1 U10613 ( .A(n9309), .B(n9308), .ZN(n9312) );
  OAI21_X1 U10614 ( .B1(n9313), .B2(n9612), .A(n9598), .ZN(n9314) );
  OAI211_X1 U10615 ( .C1(n9316), .C2(n9600), .A(n9315), .B(n9314), .ZN(
        P1_U3356) );
  XNOR2_X1 U10616 ( .A(n9318), .B(n9317), .ZN(n9321) );
  OAI22_X1 U10617 ( .A1(n9627), .A2(n9708), .B1(n9319), .B2(n9731), .ZN(n9320)
         );
  AOI21_X1 U10618 ( .B1(n9321), .B2(n9713), .A(n9320), .ZN(n9615) );
  NAND2_X1 U10619 ( .A1(n9323), .A2(n9322), .ZN(n9324) );
  NAND2_X1 U10620 ( .A1(n9617), .A2(n9556), .ZN(n9333) );
  OAI211_X1 U10621 ( .C1(n9751), .C2(n9334), .A(n9593), .B(n9326), .ZN(n9614)
         );
  INV_X1 U10622 ( .A(n9614), .ZN(n9331) );
  NOR2_X1 U10623 ( .A1(n9585), .A2(n9327), .ZN(n9489) );
  AOI22_X1 U10624 ( .A1(n9328), .A2(n9583), .B1(n9585), .B2(
        P1_REG2_REG_28__SCAN_IN), .ZN(n9329) );
  OAI21_X1 U10625 ( .B1(n9751), .B2(n9590), .A(n9329), .ZN(n9330) );
  AOI21_X1 U10626 ( .B1(n9331), .B2(n9489), .A(n9330), .ZN(n9332) );
  OAI211_X1 U10627 ( .C1(n9615), .C2(n9585), .A(n9333), .B(n9332), .ZN(
        P1_U3265) );
  AOI21_X1 U10628 ( .B1(n9620), .B2(n9353), .A(n9494), .ZN(n9335) );
  AND2_X1 U10629 ( .A1(n9336), .A2(n9583), .ZN(n9342) );
  OAI21_X1 U10630 ( .B1(n9344), .B2(n9338), .A(n9337), .ZN(n9339) );
  INV_X1 U10631 ( .A(n9339), .ZN(n9340) );
  OAI222_X1 U10632 ( .A1(n9708), .A2(n9341), .B1(n9731), .B2(n9607), .C1(n9693), .C2(n9340), .ZN(n9621) );
  AOI211_X1 U10633 ( .C1(n9622), .C2(n9343), .A(n9342), .B(n9621), .ZN(n9348)
         );
  XNOR2_X1 U10634 ( .A(n9345), .B(n9344), .ZN(n9623) );
  NAND2_X1 U10635 ( .A1(n9623), .A2(n9556), .ZN(n9347) );
  AOI22_X1 U10636 ( .A1(n9620), .A2(n9569), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9585), .ZN(n9346) );
  OAI211_X1 U10637 ( .C1(n9585), .C2(n9348), .A(n9347), .B(n9346), .ZN(
        P1_U3266) );
  XNOR2_X1 U10638 ( .A(n9349), .B(n9351), .ZN(n9633) );
  INV_X1 U10639 ( .A(n9633), .ZN(n9365) );
  OAI21_X1 U10640 ( .B1(n9352), .B2(n9351), .A(n9350), .ZN(n9630) );
  INV_X1 U10641 ( .A(n9355), .ZN(n9758) );
  INV_X1 U10642 ( .A(n9353), .ZN(n9354) );
  AOI211_X1 U10643 ( .C1(n9355), .C2(n9369), .A(n9494), .B(n9354), .ZN(n9628)
         );
  NAND2_X1 U10644 ( .A1(n9628), .A2(n9538), .ZN(n9362) );
  INV_X1 U10645 ( .A(n9356), .ZN(n9357) );
  AOI22_X1 U10646 ( .A1(n9585), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9357), .B2(
        n9583), .ZN(n9358) );
  OAI21_X1 U10647 ( .B1(n9626), .B2(n9561), .A(n9358), .ZN(n9359) );
  AOI21_X1 U10648 ( .B1(n9587), .B2(n9360), .A(n9359), .ZN(n9361) );
  OAI211_X1 U10649 ( .C1(n9758), .C2(n9590), .A(n9362), .B(n9361), .ZN(n9363)
         );
  AOI21_X1 U10650 ( .B1(n9548), .B2(n9630), .A(n9363), .ZN(n9364) );
  OAI21_X1 U10651 ( .B1(n9365), .B2(n9600), .A(n9364), .ZN(P1_U3267) );
  XOR2_X1 U10652 ( .A(n9366), .B(n9367), .Z(n9643) );
  OAI21_X1 U10653 ( .B1(n4554), .B2(n4747), .A(n9368), .ZN(n9641) );
  OAI211_X1 U10654 ( .C1(n9639), .C2(n9389), .A(n9593), .B(n9369), .ZN(n9638)
         );
  OAI22_X1 U10655 ( .A1(n9598), .A2(n9371), .B1(n9370), .B2(n9557), .ZN(n9372)
         );
  AOI21_X1 U10656 ( .B1(n9636), .B2(n9587), .A(n9372), .ZN(n9373) );
  OAI21_X1 U10657 ( .B1(n9374), .B2(n9561), .A(n9373), .ZN(n9375) );
  AOI21_X1 U10658 ( .B1(n9376), .B2(n9569), .A(n9375), .ZN(n9377) );
  OAI21_X1 U10659 ( .B1(n9638), .B2(n9595), .A(n9377), .ZN(n9378) );
  AOI21_X1 U10660 ( .B1(n9641), .B2(n9548), .A(n9378), .ZN(n9379) );
  OAI21_X1 U10661 ( .B1(n9643), .B2(n9600), .A(n9379), .ZN(P1_U3268) );
  XOR2_X1 U10662 ( .A(n9382), .B(n9380), .Z(n9646) );
  INV_X1 U10663 ( .A(n9646), .ZN(n9396) );
  NAND2_X1 U10664 ( .A1(n9398), .A2(n9381), .ZN(n9383) );
  NAND2_X1 U10665 ( .A1(n9383), .A2(n9382), .ZN(n9385) );
  NAND3_X1 U10666 ( .A1(n9385), .A2(n9713), .A3(n9384), .ZN(n9388) );
  AOI22_X1 U10667 ( .A1(n9386), .A2(n9720), .B1(n9721), .B2(n9658), .ZN(n9387)
         );
  NAND2_X1 U10668 ( .A1(n9388), .A2(n9387), .ZN(n9644) );
  AOI211_X1 U10669 ( .C1(n9390), .C2(n9401), .A(n9494), .B(n9389), .ZN(n9645)
         );
  NAND2_X1 U10670 ( .A1(n9645), .A2(n9489), .ZN(n9393) );
  AOI22_X1 U10671 ( .A1(n9585), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9391), .B2(
        n9583), .ZN(n9392) );
  OAI211_X1 U10672 ( .C1(n9763), .C2(n9590), .A(n9393), .B(n9392), .ZN(n9394)
         );
  AOI21_X1 U10673 ( .B1(n9598), .B2(n9644), .A(n9394), .ZN(n9395) );
  OAI21_X1 U10674 ( .B1(n9396), .B2(n9600), .A(n9395), .ZN(P1_U3269) );
  XNOR2_X1 U10675 ( .A(n9397), .B(n9399), .ZN(n9656) );
  OAI21_X1 U10676 ( .B1(n9400), .B2(n9399), .A(n9398), .ZN(n9654) );
  AOI21_X1 U10677 ( .B1(n9408), .B2(n9417), .A(n9494), .ZN(n9402) );
  NAND2_X1 U10678 ( .A1(n9402), .A2(n9401), .ZN(n9651) );
  OAI22_X1 U10679 ( .A1(n9598), .A2(n9404), .B1(n9403), .B2(n9557), .ZN(n9407)
         );
  NOR2_X1 U10680 ( .A1(n9561), .A2(n9405), .ZN(n9406) );
  AOI211_X1 U10681 ( .C1(n9587), .C2(n9649), .A(n9407), .B(n9406), .ZN(n9410)
         );
  NAND2_X1 U10682 ( .A1(n9408), .A2(n9569), .ZN(n9409) );
  OAI211_X1 U10683 ( .C1(n9651), .C2(n9595), .A(n9410), .B(n9409), .ZN(n9411)
         );
  AOI21_X1 U10684 ( .B1(n9654), .B2(n9548), .A(n9411), .ZN(n9412) );
  OAI21_X1 U10685 ( .B1(n9656), .B2(n9600), .A(n9412), .ZN(P1_U3270) );
  XNOR2_X1 U10686 ( .A(n9414), .B(n9413), .ZN(n9665) );
  XNOR2_X1 U10687 ( .A(n9416), .B(n9415), .ZN(n9663) );
  OAI211_X1 U10688 ( .C1(n9661), .C2(n9434), .A(n9593), .B(n9417), .ZN(n9660)
         );
  OAI22_X1 U10689 ( .A1(n9598), .A2(n9419), .B1(n9418), .B2(n9557), .ZN(n9421)
         );
  NOR2_X1 U10690 ( .A1(n9561), .A2(n9280), .ZN(n9420) );
  AOI211_X1 U10691 ( .C1(n9587), .C2(n9658), .A(n9421), .B(n9420), .ZN(n9424)
         );
  NAND2_X1 U10692 ( .A1(n9422), .A2(n9569), .ZN(n9423) );
  OAI211_X1 U10693 ( .C1(n9660), .C2(n9595), .A(n9424), .B(n9423), .ZN(n9425)
         );
  AOI21_X1 U10694 ( .B1(n9663), .B2(n9548), .A(n9425), .ZN(n9426) );
  OAI21_X1 U10695 ( .B1(n9665), .B2(n9600), .A(n9426), .ZN(P1_U3271) );
  XNOR2_X1 U10696 ( .A(n9428), .B(n9427), .ZN(n9673) );
  OAI21_X1 U10697 ( .B1(n5106), .B2(n9430), .A(n9429), .ZN(n9671) );
  NAND2_X1 U10698 ( .A1(n9431), .A2(n9445), .ZN(n9432) );
  NAND2_X1 U10699 ( .A1(n9432), .A2(n9593), .ZN(n9433) );
  NOR2_X1 U10700 ( .A1(n9434), .A2(n9433), .ZN(n9670) );
  NAND2_X1 U10701 ( .A1(n9670), .A2(n9538), .ZN(n9441) );
  OAI22_X1 U10702 ( .A1(n9598), .A2(n9436), .B1(n9435), .B2(n9557), .ZN(n9439)
         );
  NOR2_X1 U10703 ( .A1(n9561), .A2(n9437), .ZN(n9438) );
  AOI211_X1 U10704 ( .C1(n9587), .C2(n9667), .A(n9439), .B(n9438), .ZN(n9440)
         );
  OAI211_X1 U10705 ( .C1(n9281), .C2(n9590), .A(n9441), .B(n9440), .ZN(n9442)
         );
  AOI21_X1 U10706 ( .B1(n9671), .B2(n9548), .A(n9442), .ZN(n9443) );
  OAI21_X1 U10707 ( .B1(n9673), .B2(n9600), .A(n9443), .ZN(P1_U3272) );
  XOR2_X1 U10708 ( .A(n9444), .B(n9454), .Z(n9678) );
  INV_X1 U10709 ( .A(n9468), .ZN(n9447) );
  INV_X1 U10710 ( .A(n9445), .ZN(n9446) );
  AOI211_X1 U10711 ( .C1(n9676), .C2(n9447), .A(n9494), .B(n9446), .ZN(n9675)
         );
  NOR2_X1 U10712 ( .A1(n9448), .A2(n9590), .ZN(n9452) );
  OAI22_X1 U10713 ( .A1(n9598), .A2(n9450), .B1(n9449), .B2(n9557), .ZN(n9451)
         );
  AOI211_X1 U10714 ( .C1(n9675), .C2(n9538), .A(n9452), .B(n9451), .ZN(n9459)
         );
  OAI211_X1 U10715 ( .C1(n9455), .C2(n9454), .A(n9453), .B(n9713), .ZN(n9457)
         );
  AOI22_X1 U10716 ( .A1(n9721), .A2(n9485), .B1(n9657), .B2(n9720), .ZN(n9456)
         );
  NAND2_X1 U10717 ( .A1(n9457), .A2(n9456), .ZN(n9674) );
  NAND2_X1 U10718 ( .A1(n9674), .A2(n9598), .ZN(n9458) );
  OAI211_X1 U10719 ( .C1(n9678), .C2(n9600), .A(n9459), .B(n9458), .ZN(
        P1_U3273) );
  XNOR2_X1 U10720 ( .A(n9461), .B(n9460), .ZN(n9683) );
  NAND2_X1 U10721 ( .A1(n9462), .A2(n9713), .ZN(n9467) );
  AOI21_X1 U10722 ( .B1(n9474), .B2(n9464), .A(n9463), .ZN(n9466) );
  AOI22_X1 U10723 ( .A1(n9721), .A2(n9505), .B1(n9666), .B2(n9720), .ZN(n9465)
         );
  OAI21_X1 U10724 ( .B1(n9467), .B2(n9466), .A(n9465), .ZN(n9679) );
  AOI211_X1 U10725 ( .C1(n9681), .C2(n9479), .A(n9494), .B(n9468), .ZN(n9680)
         );
  NAND2_X1 U10726 ( .A1(n9680), .A2(n9538), .ZN(n9471) );
  AOI22_X1 U10727 ( .A1(n9585), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9469), .B2(
        n9583), .ZN(n9470) );
  OAI211_X1 U10728 ( .C1(n4711), .C2(n9590), .A(n9471), .B(n9470), .ZN(n9472)
         );
  AOI21_X1 U10729 ( .B1(n9598), .B2(n9679), .A(n9472), .ZN(n9473) );
  OAI21_X1 U10730 ( .B1(n9683), .B2(n9600), .A(n9473), .ZN(P1_U3274) );
  AOI21_X1 U10731 ( .B1(n9476), .B2(n9475), .A(n8247), .ZN(n9692) );
  XNOR2_X1 U10732 ( .A(n9477), .B(n9476), .ZN(n9684) );
  NAND2_X1 U10733 ( .A1(n9684), .A2(n9556), .ZN(n9491) );
  INV_X1 U10734 ( .A(n9479), .ZN(n9480) );
  AOI211_X1 U10735 ( .C1(n9689), .C2(n4715), .A(n9494), .B(n9480), .ZN(n9687)
         );
  OAI22_X1 U10736 ( .A1(n9598), .A2(n9482), .B1(n9481), .B2(n9557), .ZN(n9484)
         );
  NOR2_X1 U10737 ( .A1(n9561), .A2(n9685), .ZN(n9483) );
  AOI211_X1 U10738 ( .C1(n9587), .C2(n9485), .A(n9484), .B(n9483), .ZN(n9486)
         );
  OAI21_X1 U10739 ( .B1(n9487), .B2(n9590), .A(n9486), .ZN(n9488) );
  AOI21_X1 U10740 ( .B1(n9687), .B2(n9489), .A(n9488), .ZN(n9490) );
  OAI211_X1 U10741 ( .C1(n9692), .C2(n9492), .A(n9491), .B(n9490), .ZN(
        P1_U3275) );
  XNOR2_X1 U10742 ( .A(n9493), .B(n9500), .ZN(n9698) );
  AOI211_X1 U10743 ( .C1(n9696), .C2(n9522), .A(n9494), .B(n9478), .ZN(n9695)
         );
  NOR2_X1 U10744 ( .A1(n9495), .A2(n9590), .ZN(n9499) );
  OAI22_X1 U10745 ( .A1(n9598), .A2(n9497), .B1(n9496), .B2(n9557), .ZN(n9498)
         );
  AOI211_X1 U10746 ( .C1(n9695), .C2(n9538), .A(n9499), .B(n9498), .ZN(n9509)
         );
  INV_X1 U10747 ( .A(n9519), .ZN(n9502) );
  OAI21_X1 U10748 ( .B1(n9502), .B2(n9501), .A(n9500), .ZN(n9504) );
  NAND3_X1 U10749 ( .A1(n9504), .A2(n9503), .A3(n9713), .ZN(n9507) );
  NAND2_X1 U10750 ( .A1(n9505), .A2(n9720), .ZN(n9506) );
  OAI211_X1 U10751 ( .C1(n9707), .C2(n9708), .A(n9507), .B(n9506), .ZN(n9694)
         );
  NAND2_X1 U10752 ( .A1(n9694), .A2(n9598), .ZN(n9508) );
  OAI211_X1 U10753 ( .C1(n9698), .C2(n9600), .A(n9509), .B(n9508), .ZN(
        P1_U3276) );
  INV_X1 U10754 ( .A(n9510), .ZN(n9511) );
  NOR2_X1 U10755 ( .A1(n9512), .A2(n9511), .ZN(n9533) );
  INV_X1 U10756 ( .A(n9513), .ZN(n9514) );
  AOI21_X1 U10757 ( .B1(n9533), .B2(n9515), .A(n9514), .ZN(n9518) );
  OAI21_X1 U10758 ( .B1(n9518), .B2(n9517), .A(n9516), .ZN(n9706) );
  OAI21_X1 U10759 ( .B1(n9521), .B2(n9520), .A(n9519), .ZN(n9704) );
  OAI211_X1 U10760 ( .C1(n9536), .C2(n9702), .A(n9593), .B(n9522), .ZN(n9701)
         );
  OAI22_X1 U10761 ( .A1(n9598), .A2(n9524), .B1(n9523), .B2(n9557), .ZN(n9527)
         );
  NOR2_X1 U10762 ( .A1(n9561), .A2(n9525), .ZN(n9526) );
  AOI211_X1 U10763 ( .C1(n9587), .C2(n9699), .A(n9527), .B(n9526), .ZN(n9530)
         );
  NAND2_X1 U10764 ( .A1(n9528), .A2(n9569), .ZN(n9529) );
  OAI211_X1 U10765 ( .C1(n9701), .C2(n9595), .A(n9530), .B(n9529), .ZN(n9531)
         );
  AOI21_X1 U10766 ( .B1(n9704), .B2(n9548), .A(n9531), .ZN(n9532) );
  OAI21_X1 U10767 ( .B1(n9706), .B2(n9600), .A(n9532), .ZN(P1_U3277) );
  XNOR2_X1 U10768 ( .A(n9533), .B(n9534), .ZN(n9718) );
  XNOR2_X1 U10769 ( .A(n9535), .B(n9534), .ZN(n9714) );
  OAI21_X1 U10770 ( .B1(n9565), .B2(n9546), .A(n9593), .ZN(n9537) );
  NOR2_X1 U10771 ( .A1(n9537), .A2(n9536), .ZN(n9709) );
  NAND2_X1 U10772 ( .A1(n9709), .A2(n9538), .ZN(n9545) );
  OAI22_X1 U10773 ( .A1(n9598), .A2(n9540), .B1(n9539), .B2(n9557), .ZN(n9542)
         );
  NOR2_X1 U10774 ( .A1(n9561), .A2(n9732), .ZN(n9541) );
  AOI211_X1 U10775 ( .C1(n9587), .C2(n9543), .A(n9542), .B(n9541), .ZN(n9544)
         );
  OAI211_X1 U10776 ( .C1(n9546), .C2(n9590), .A(n9545), .B(n9544), .ZN(n9547)
         );
  AOI21_X1 U10777 ( .B1(n9714), .B2(n9548), .A(n9547), .ZN(n9549) );
  OAI21_X1 U10778 ( .B1(n9718), .B2(n9600), .A(n9549), .ZN(P1_U3278) );
  OAI21_X1 U10779 ( .B1(n9552), .B2(n9551), .A(n9550), .ZN(n9553) );
  NAND2_X1 U10780 ( .A1(n9553), .A2(n9713), .ZN(n9725) );
  XNOR2_X1 U10781 ( .A(n9555), .B(n9554), .ZN(n9727) );
  NAND2_X1 U10782 ( .A1(n9727), .A2(n9556), .ZN(n9571) );
  OAI22_X1 U10783 ( .A1(n9598), .A2(n6960), .B1(n9558), .B2(n9557), .ZN(n9559)
         );
  AOI21_X1 U10784 ( .B1(n9587), .B2(n9719), .A(n9559), .ZN(n9560) );
  OAI21_X1 U10785 ( .B1(n9562), .B2(n9561), .A(n9560), .ZN(n9567) );
  NAND2_X1 U10786 ( .A1(n9592), .A2(n9568), .ZN(n9563) );
  NAND2_X1 U10787 ( .A1(n9563), .A2(n9593), .ZN(n9564) );
  OR2_X1 U10788 ( .A1(n9565), .A2(n9564), .ZN(n9723) );
  NOR2_X1 U10789 ( .A1(n9723), .A2(n9595), .ZN(n9566) );
  AOI211_X1 U10790 ( .C1(n9569), .C2(n9568), .A(n9567), .B(n9566), .ZN(n9570)
         );
  OAI211_X1 U10791 ( .C1(n9585), .C2(n9725), .A(n9571), .B(n9570), .ZN(
        P1_U3279) );
  OAI21_X1 U10792 ( .B1(n9573), .B2(n9576), .A(n9572), .ZN(n9735) );
  INV_X1 U10793 ( .A(n9735), .ZN(n9601) );
  NAND2_X1 U10794 ( .A1(n9575), .A2(n9574), .ZN(n9577) );
  NAND2_X1 U10795 ( .A1(n9577), .A2(n9576), .ZN(n9579) );
  NAND3_X1 U10796 ( .A1(n9579), .A2(n9578), .A3(n9713), .ZN(n9582) );
  OR2_X1 U10797 ( .A1(n9580), .A2(n9708), .ZN(n9581) );
  NAND2_X1 U10798 ( .A1(n9582), .A2(n9581), .ZN(n9734) );
  AOI22_X1 U10799 ( .A1(n9585), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9584), .B2(
        n9583), .ZN(n9589) );
  NAND2_X1 U10800 ( .A1(n9587), .A2(n9586), .ZN(n9588) );
  OAI211_X1 U10801 ( .C1(n9779), .C2(n9590), .A(n9589), .B(n9588), .ZN(n9597)
         );
  INV_X1 U10802 ( .A(n9591), .ZN(n9594) );
  OAI211_X1 U10803 ( .C1(n9594), .C2(n9779), .A(n9593), .B(n9592), .ZN(n9730)
         );
  NOR2_X1 U10804 ( .A1(n9730), .A2(n9595), .ZN(n9596) );
  AOI211_X1 U10805 ( .C1(n9734), .C2(n9598), .A(n9597), .B(n9596), .ZN(n9599)
         );
  OAI21_X1 U10806 ( .B1(n9601), .B2(n9600), .A(n9599), .ZN(P1_U3280) );
  NOR2_X1 U10807 ( .A1(n9603), .A2(n9602), .ZN(n9743) );
  MUX2_X1 U10808 ( .A(n9604), .B(n9743), .S(n9850), .Z(n9605) );
  OAI21_X1 U10809 ( .B1(n9746), .B2(n9742), .A(n9605), .ZN(P1_U3552) );
  NAND2_X1 U10810 ( .A1(n9606), .A2(n9834), .ZN(n9613) );
  INV_X1 U10811 ( .A(n8101), .ZN(n9608) );
  OAI22_X1 U10812 ( .A1(n9608), .A2(n9831), .B1(n9607), .B2(n9708), .ZN(n9609)
         );
  NAND2_X1 U10813 ( .A1(n9615), .A2(n9614), .ZN(n9616) );
  AOI21_X1 U10814 ( .B1(n9617), .B2(n9834), .A(n9616), .ZN(n9748) );
  MUX2_X1 U10815 ( .A(n9618), .B(n9748), .S(n9850), .Z(n9619) );
  OAI21_X1 U10816 ( .B1(n9751), .B2(n9742), .A(n9619), .ZN(P1_U3550) );
  AOI211_X1 U10817 ( .C1(n9623), .C2(n9834), .A(n9622), .B(n9621), .ZN(n9752)
         );
  MUX2_X1 U10818 ( .A(n9624), .B(n9752), .S(n9850), .Z(n9625) );
  OAI21_X1 U10819 ( .B1(n4717), .B2(n9742), .A(n9625), .ZN(P1_U3549) );
  OAI22_X1 U10820 ( .A1(n9627), .A2(n9731), .B1(n9626), .B2(n9708), .ZN(n9629)
         );
  AOI211_X1 U10821 ( .C1(n9713), .C2(n9630), .A(n9629), .B(n9628), .ZN(n9631)
         );
  INV_X1 U10822 ( .A(n9631), .ZN(n9632) );
  AOI21_X1 U10823 ( .B1(n9633), .B2(n9834), .A(n9632), .ZN(n9755) );
  MUX2_X1 U10824 ( .A(n9634), .B(n9755), .S(n9850), .Z(n9635) );
  OAI21_X1 U10825 ( .B1(n9758), .B2(n9742), .A(n9635), .ZN(P1_U3548) );
  AOI22_X1 U10826 ( .A1(n9636), .A2(n9720), .B1(n9721), .B2(n9649), .ZN(n9637)
         );
  OAI211_X1 U10827 ( .C1(n9639), .C2(n9831), .A(n9638), .B(n9637), .ZN(n9640)
         );
  AOI21_X1 U10828 ( .B1(n9641), .B2(n9713), .A(n9640), .ZN(n9642) );
  OAI21_X1 U10829 ( .B1(n9643), .B2(n9717), .A(n9642), .ZN(n9759) );
  MUX2_X1 U10830 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9759), .S(n9850), .Z(
        P1_U3547) );
  INV_X1 U10831 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9647) );
  AOI211_X1 U10832 ( .C1(n9646), .C2(n9834), .A(n9645), .B(n9644), .ZN(n9760)
         );
  MUX2_X1 U10833 ( .A(n9647), .B(n9760), .S(n9850), .Z(n9648) );
  OAI21_X1 U10834 ( .B1(n9763), .B2(n9742), .A(n9648), .ZN(P1_U3546) );
  AOI22_X1 U10835 ( .A1(n9649), .A2(n9720), .B1(n9721), .B2(n9667), .ZN(n9650)
         );
  OAI211_X1 U10836 ( .C1(n9652), .C2(n9831), .A(n9651), .B(n9650), .ZN(n9653)
         );
  AOI21_X1 U10837 ( .B1(n9654), .B2(n9713), .A(n9653), .ZN(n9655) );
  OAI21_X1 U10838 ( .B1(n9656), .B2(n9717), .A(n9655), .ZN(n9764) );
  MUX2_X1 U10839 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9764), .S(n9850), .Z(
        P1_U3545) );
  AOI22_X1 U10840 ( .A1(n9658), .A2(n9720), .B1(n9657), .B2(n9721), .ZN(n9659)
         );
  OAI211_X1 U10841 ( .C1(n9661), .C2(n9831), .A(n9660), .B(n9659), .ZN(n9662)
         );
  AOI21_X1 U10842 ( .B1(n9663), .B2(n9713), .A(n9662), .ZN(n9664) );
  OAI21_X1 U10843 ( .B1(n9665), .B2(n9717), .A(n9664), .ZN(n9765) );
  MUX2_X1 U10844 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9765), .S(n9850), .Z(
        P1_U3544) );
  AOI22_X1 U10845 ( .A1(n9667), .A2(n9720), .B1(n9721), .B2(n9666), .ZN(n9668)
         );
  OAI21_X1 U10846 ( .B1(n9281), .B2(n9831), .A(n9668), .ZN(n9669) );
  AOI211_X1 U10847 ( .C1(n9671), .C2(n9713), .A(n9670), .B(n9669), .ZN(n9672)
         );
  OAI21_X1 U10848 ( .B1(n9673), .B2(n9717), .A(n9672), .ZN(n9766) );
  MUX2_X1 U10849 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9766), .S(n9850), .Z(
        P1_U3543) );
  AOI211_X1 U10850 ( .C1(n9712), .C2(n9676), .A(n9675), .B(n9674), .ZN(n9677)
         );
  OAI21_X1 U10851 ( .B1(n9678), .B2(n9717), .A(n9677), .ZN(n9767) );
  MUX2_X1 U10852 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9767), .S(n9850), .Z(
        P1_U3542) );
  AOI211_X1 U10853 ( .C1(n9712), .C2(n9681), .A(n9680), .B(n9679), .ZN(n9682)
         );
  OAI21_X1 U10854 ( .B1(n9683), .B2(n9717), .A(n9682), .ZN(n9768) );
  MUX2_X1 U10855 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9768), .S(n9850), .Z(
        P1_U3541) );
  NAND2_X1 U10856 ( .A1(n9684), .A2(n9834), .ZN(n9691) );
  OAI22_X1 U10857 ( .A1(n9686), .A2(n9731), .B1(n9685), .B2(n9708), .ZN(n9688)
         );
  AOI211_X1 U10858 ( .C1(n9712), .C2(n9689), .A(n9688), .B(n9687), .ZN(n9690)
         );
  OAI211_X1 U10859 ( .C1(n9693), .C2(n9692), .A(n9691), .B(n9690), .ZN(n9769)
         );
  MUX2_X1 U10860 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9769), .S(n9850), .Z(
        P1_U3540) );
  AOI211_X1 U10861 ( .C1(n9712), .C2(n9696), .A(n9695), .B(n9694), .ZN(n9697)
         );
  OAI21_X1 U10862 ( .B1(n9698), .B2(n9717), .A(n9697), .ZN(n9770) );
  MUX2_X1 U10863 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9770), .S(n9850), .Z(
        P1_U3539) );
  AOI22_X1 U10864 ( .A1(n9699), .A2(n9720), .B1(n9721), .B2(n9719), .ZN(n9700)
         );
  OAI211_X1 U10865 ( .C1(n9702), .C2(n9831), .A(n9701), .B(n9700), .ZN(n9703)
         );
  AOI21_X1 U10866 ( .B1(n9704), .B2(n9713), .A(n9703), .ZN(n9705) );
  OAI21_X1 U10867 ( .B1(n9706), .B2(n9717), .A(n9705), .ZN(n9771) );
  MUX2_X1 U10868 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9771), .S(n9850), .Z(
        P1_U3538) );
  OAI22_X1 U10869 ( .A1(n9732), .A2(n9708), .B1(n9707), .B2(n9731), .ZN(n9710)
         );
  AOI211_X1 U10870 ( .C1(n9712), .C2(n9711), .A(n9710), .B(n9709), .ZN(n9716)
         );
  NAND2_X1 U10871 ( .A1(n9714), .A2(n9713), .ZN(n9715) );
  OAI211_X1 U10872 ( .C1(n9718), .C2(n9717), .A(n9716), .B(n9715), .ZN(n9772)
         );
  MUX2_X1 U10873 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9772), .S(n9850), .Z(
        P1_U3537) );
  AOI22_X1 U10874 ( .A1(n9722), .A2(n9721), .B1(n9720), .B2(n9719), .ZN(n9724)
         );
  NAND3_X1 U10875 ( .A1(n9725), .A2(n9724), .A3(n9723), .ZN(n9726) );
  AOI21_X1 U10876 ( .B1(n9727), .B2(n9834), .A(n9726), .ZN(n9773) );
  MUX2_X1 U10877 ( .A(n9728), .B(n9773), .S(n9850), .Z(n9729) );
  OAI21_X1 U10878 ( .B1(n9776), .B2(n9742), .A(n9729), .ZN(P1_U3536) );
  OAI21_X1 U10879 ( .B1(n9732), .B2(n9731), .A(n9730), .ZN(n9733) );
  AOI211_X1 U10880 ( .C1(n9735), .C2(n9834), .A(n9734), .B(n9733), .ZN(n9777)
         );
  MUX2_X1 U10881 ( .A(n6793), .B(n9777), .S(n9850), .Z(n9736) );
  OAI21_X1 U10882 ( .B1(n9779), .B2(n9742), .A(n9736), .ZN(P1_U3535) );
  INV_X1 U10883 ( .A(n9737), .ZN(n9813) );
  AOI211_X1 U10884 ( .C1(n9813), .C2(n9740), .A(n9739), .B(n9738), .ZN(n9780)
         );
  MUX2_X1 U10885 ( .A(n7264), .B(n9780), .S(n9850), .Z(n9741) );
  OAI21_X1 U10886 ( .B1(n9784), .B2(n9742), .A(n9741), .ZN(P1_U3533) );
  MUX2_X1 U10887 ( .A(n9744), .B(n9743), .S(n9838), .Z(n9745) );
  OAI21_X1 U10888 ( .B1(n9746), .B2(n9783), .A(n9745), .ZN(P1_U3520) );
  MUX2_X1 U10889 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9747), .S(n9838), .Z(
        P1_U3519) );
  INV_X1 U10890 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9749) );
  MUX2_X1 U10891 ( .A(n9749), .B(n9748), .S(n9838), .Z(n9750) );
  OAI21_X1 U10892 ( .B1(n9751), .B2(n9783), .A(n9750), .ZN(P1_U3518) );
  INV_X1 U10893 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9753) );
  MUX2_X1 U10894 ( .A(n9753), .B(n9752), .S(n9838), .Z(n9754) );
  OAI21_X1 U10895 ( .B1(n4717), .B2(n9783), .A(n9754), .ZN(P1_U3517) );
  INV_X1 U10896 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9756) );
  MUX2_X1 U10897 ( .A(n9756), .B(n9755), .S(n9838), .Z(n9757) );
  OAI21_X1 U10898 ( .B1(n9758), .B2(n9783), .A(n9757), .ZN(P1_U3516) );
  MUX2_X1 U10899 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9759), .S(n9838), .Z(
        P1_U3515) );
  INV_X1 U10900 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9761) );
  MUX2_X1 U10901 ( .A(n9761), .B(n9760), .S(n9838), .Z(n9762) );
  OAI21_X1 U10902 ( .B1(n9763), .B2(n9783), .A(n9762), .ZN(P1_U3514) );
  MUX2_X1 U10903 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9764), .S(n9838), .Z(
        P1_U3513) );
  MUX2_X1 U10904 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9765), .S(n9838), .Z(
        P1_U3512) );
  MUX2_X1 U10905 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9766), .S(n9838), .Z(
        P1_U3511) );
  MUX2_X1 U10906 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9767), .S(n9838), .Z(
        P1_U3510) );
  MUX2_X1 U10907 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9768), .S(n9838), .Z(
        P1_U3509) );
  MUX2_X1 U10908 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9769), .S(n9838), .Z(
        P1_U3507) );
  MUX2_X1 U10909 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9770), .S(n9838), .Z(
        P1_U3504) );
  MUX2_X1 U10910 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9771), .S(n9838), .Z(
        P1_U3501) );
  MUX2_X1 U10911 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9772), .S(n9838), .Z(
        P1_U3498) );
  INV_X1 U10912 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9774) );
  MUX2_X1 U10913 ( .A(n9774), .B(n9773), .S(n9838), .Z(n9775) );
  OAI21_X1 U10914 ( .B1(n9776), .B2(n9783), .A(n9775), .ZN(P1_U3495) );
  MUX2_X1 U10915 ( .A(n7373), .B(n9777), .S(n9838), .Z(n9778) );
  OAI21_X1 U10916 ( .B1(n9779), .B2(n9783), .A(n9778), .ZN(P1_U3492) );
  INV_X1 U10917 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9781) );
  MUX2_X1 U10918 ( .A(n9781), .B(n9780), .S(n9838), .Z(n9782) );
  OAI21_X1 U10919 ( .B1(n9784), .B2(n9783), .A(n9782), .ZN(P1_U3486) );
  MUX2_X1 U10920 ( .A(n9785), .B(P1_D_REG_1__SCAN_IN), .S(n9797), .Z(P1_U3440)
         );
  NAND3_X1 U10921 ( .A1(n9786), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n9787) );
  OAI22_X1 U10922 ( .A1(n9788), .A2(n9787), .B1(n10446), .B2(n6832), .ZN(n9789) );
  AOI21_X1 U10923 ( .B1(n8976), .B2(n9790), .A(n9789), .ZN(n9791) );
  INV_X1 U10924 ( .A(n9791), .ZN(P1_U3324) );
  OAI222_X1 U10925 ( .A1(n6832), .A2(n10190), .B1(P1_U3086), .B2(n9793), .C1(
        n9792), .C2(n7300), .ZN(P1_U3328) );
  OAI222_X1 U10926 ( .A1(n6832), .A2(n10489), .B1(n7300), .B2(n9795), .C1(
        P1_U3086), .C2(n9794), .ZN(P1_U3330) );
  MUX2_X1 U10927 ( .A(n9796), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U10928 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10929 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  AND2_X1 U10930 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9797), .ZN(P1_U3294) );
  AND2_X1 U10931 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9797), .ZN(P1_U3295) );
  AND2_X1 U10932 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9797), .ZN(P1_U3296) );
  AND2_X1 U10933 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9797), .ZN(P1_U3297) );
  AND2_X1 U10934 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9797), .ZN(P1_U3298) );
  AND2_X1 U10935 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9797), .ZN(P1_U3299) );
  AND2_X1 U10936 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9797), .ZN(P1_U3300) );
  AND2_X1 U10937 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9797), .ZN(P1_U3301) );
  AND2_X1 U10938 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9797), .ZN(P1_U3302) );
  AND2_X1 U10939 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9797), .ZN(P1_U3303) );
  AND2_X1 U10940 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9797), .ZN(P1_U3304) );
  AND2_X1 U10941 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9797), .ZN(P1_U3305) );
  AND2_X1 U10942 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9797), .ZN(P1_U3306) );
  AND2_X1 U10943 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9797), .ZN(P1_U3307) );
  AND2_X1 U10944 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9797), .ZN(P1_U3308) );
  AND2_X1 U10945 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9797), .ZN(P1_U3309) );
  AND2_X1 U10946 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9797), .ZN(P1_U3310) );
  AND2_X1 U10947 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9797), .ZN(P1_U3311) );
  AND2_X1 U10948 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9797), .ZN(P1_U3312) );
  AND2_X1 U10949 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9797), .ZN(P1_U3313) );
  AND2_X1 U10950 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9797), .ZN(P1_U3314) );
  AND2_X1 U10951 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9797), .ZN(P1_U3315) );
  AND2_X1 U10952 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9797), .ZN(P1_U3316) );
  AND2_X1 U10953 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9797), .ZN(P1_U3317) );
  AND2_X1 U10954 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9797), .ZN(P1_U3318) );
  AND2_X1 U10955 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9797), .ZN(P1_U3319) );
  NOR2_X1 U10956 ( .A1(n9799), .A2(n10429), .ZN(P1_U3320) );
  NOR2_X1 U10957 ( .A1(n9799), .A2(n10487), .ZN(P1_U3321) );
  NOR2_X1 U10958 ( .A1(n9799), .A2(n10368), .ZN(P1_U3322) );
  NOR2_X1 U10959 ( .A1(n9799), .A2(n9798), .ZN(P1_U3323) );
  OAI21_X1 U10960 ( .B1(n9801), .B2(n9831), .A(n9800), .ZN(n9803) );
  AOI211_X1 U10961 ( .C1(n9834), .C2(n9804), .A(n9803), .B(n9802), .ZN(n9840)
         );
  AOI22_X1 U10962 ( .A1(n9838), .A2(n9840), .B1(n6552), .B2(n9836), .ZN(
        P1_U3465) );
  OAI21_X1 U10963 ( .B1(n9806), .B2(n9831), .A(n9805), .ZN(n9808) );
  AOI211_X1 U10964 ( .C1(n9834), .C2(n9809), .A(n9808), .B(n9807), .ZN(n9842)
         );
  AOI22_X1 U10965 ( .A1(n9838), .A2(n9842), .B1(n6739), .B2(n9836), .ZN(
        P1_U3471) );
  OAI21_X1 U10966 ( .B1(n9811), .B2(n9831), .A(n9810), .ZN(n9812) );
  AOI21_X1 U10967 ( .B1(n9814), .B2(n9813), .A(n9812), .ZN(n9815) );
  AND2_X1 U10968 ( .A1(n9816), .A2(n9815), .ZN(n9844) );
  AOI22_X1 U10969 ( .A1(n9838), .A2(n9844), .B1(n7038), .B2(n9836), .ZN(
        P1_U3477) );
  OAI211_X1 U10970 ( .C1(n7274), .C2(n9831), .A(n9819), .B(n9818), .ZN(n9820)
         );
  AOI21_X1 U10971 ( .B1(n9834), .B2(n9821), .A(n9820), .ZN(n9845) );
  INV_X1 U10972 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9822) );
  AOI22_X1 U10973 ( .A1(n9838), .A2(n9845), .B1(n9822), .B2(n9836), .ZN(
        P1_U3480) );
  OAI211_X1 U10974 ( .C1(n9825), .C2(n9831), .A(n9824), .B(n9823), .ZN(n9826)
         );
  AOI21_X1 U10975 ( .B1(n9827), .B2(n9834), .A(n9826), .ZN(n9846) );
  INV_X1 U10976 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9828) );
  AOI22_X1 U10977 ( .A1(n9838), .A2(n9846), .B1(n9828), .B2(n9836), .ZN(
        P1_U3483) );
  OAI211_X1 U10978 ( .C1(n9832), .C2(n9831), .A(n9830), .B(n9829), .ZN(n9833)
         );
  AOI21_X1 U10979 ( .B1(n9835), .B2(n9834), .A(n9833), .ZN(n9849) );
  INV_X1 U10980 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9837) );
  AOI22_X1 U10981 ( .A1(n9838), .A2(n9849), .B1(n9837), .B2(n9836), .ZN(
        P1_U3489) );
  INV_X1 U10982 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9839) );
  AOI22_X1 U10983 ( .A1(n9850), .A2(n9840), .B1(n9839), .B2(n9847), .ZN(
        P1_U3526) );
  INV_X1 U10984 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9841) );
  AOI22_X1 U10985 ( .A1(n9850), .A2(n9842), .B1(n9841), .B2(n9847), .ZN(
        P1_U3528) );
  INV_X1 U10986 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9843) );
  AOI22_X1 U10987 ( .A1(n9850), .A2(n9844), .B1(n9843), .B2(n9847), .ZN(
        P1_U3530) );
  AOI22_X1 U10988 ( .A1(n9850), .A2(n9845), .B1(n7052), .B2(n9847), .ZN(
        P1_U3531) );
  AOI22_X1 U10989 ( .A1(n9850), .A2(n9846), .B1(n7239), .B2(n9847), .ZN(
        P1_U3532) );
  AOI22_X1 U10990 ( .A1(n9850), .A2(n9849), .B1(n9848), .B2(n9847), .ZN(
        P1_U3534) );
  INV_X1 U10991 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10091) );
  NAND2_X1 U10992 ( .A1(n9851), .A2(n6155), .ZN(n9852) );
  NAND2_X1 U10993 ( .A1(n9853), .A2(n9852), .ZN(n9854) );
  AOI22_X1 U10994 ( .A1(n9877), .A2(n9854), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        P2_U3151), .ZN(n9859) );
  OAI211_X1 U10995 ( .C1(n9857), .C2(n9856), .A(n9855), .B(n9967), .ZN(n9858)
         );
  OAI211_X1 U10996 ( .C1(n9977), .C2(n9860), .A(n9859), .B(n9858), .ZN(n9861)
         );
  INV_X1 U10997 ( .A(n9861), .ZN(n9866) );
  AOI21_X1 U10998 ( .B1(n8803), .B2(n9863), .A(n9862), .ZN(n9864) );
  OR2_X1 U10999 ( .A1(n9963), .A2(n9864), .ZN(n9865) );
  OAI211_X1 U11000 ( .C1(n10091), .C2(n9888), .A(n9866), .B(n9865), .ZN(
        P2_U3183) );
  INV_X1 U11001 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n9889) );
  OAI211_X1 U11002 ( .C1(n9869), .C2(n9868), .A(n9867), .B(n9967), .ZN(n9879)
         );
  INV_X1 U11003 ( .A(n9870), .ZN(n9871) );
  OAI21_X1 U11004 ( .B1(n9873), .B2(n9872), .A(n9871), .ZN(n9876) );
  NOR2_X1 U11005 ( .A1(n9874), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9875) );
  AOI21_X1 U11006 ( .B1(n9877), .B2(n9876), .A(n9875), .ZN(n9878) );
  OAI211_X1 U11007 ( .C1(n9977), .C2(n9880), .A(n9879), .B(n9878), .ZN(n9881)
         );
  INV_X1 U11008 ( .A(n9881), .ZN(n9887) );
  AOI21_X1 U11009 ( .B1(n9884), .B2(n9883), .A(n9882), .ZN(n9885) );
  OR2_X1 U11010 ( .A1(n9963), .A2(n9885), .ZN(n9886) );
  OAI211_X1 U11011 ( .C1(n9889), .C2(n9888), .A(n9887), .B(n9886), .ZN(
        P2_U3184) );
  AOI22_X1 U11012 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3151), .B1(n9957), 
        .B2(P2_ADDR_REG_12__SCAN_IN), .ZN(n9904) );
  AOI21_X1 U11013 ( .B1(n4594), .B2(n9891), .A(n9890), .ZN(n9901) );
  AOI21_X1 U11014 ( .B1(n4595), .B2(n9893), .A(n9892), .ZN(n9894) );
  OR2_X1 U11015 ( .A1(n9894), .A2(n9963), .ZN(n9900) );
  OAI21_X1 U11016 ( .B1(n9897), .B2(n9896), .A(n9895), .ZN(n9898) );
  NAND2_X1 U11017 ( .A1(n9898), .A2(n9967), .ZN(n9899) );
  OAI211_X1 U11018 ( .C1(n9901), .C2(n9971), .A(n9900), .B(n9899), .ZN(n9902)
         );
  INV_X1 U11019 ( .A(n9902), .ZN(n9903) );
  OAI211_X1 U11020 ( .C1(n9977), .C2(n9905), .A(n9904), .B(n9903), .ZN(
        P2_U3194) );
  AOI22_X1 U11021 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3151), .B1(n9957), 
        .B2(P2_ADDR_REG_13__SCAN_IN), .ZN(n9922) );
  AOI21_X1 U11022 ( .B1(n9908), .B2(n9907), .A(n9906), .ZN(n9919) );
  OAI21_X1 U11023 ( .B1(n9911), .B2(n9910), .A(n9909), .ZN(n9912) );
  NAND2_X1 U11024 ( .A1(n9912), .A2(n9967), .ZN(n9918) );
  AOI21_X1 U11025 ( .B1(n9915), .B2(n9914), .A(n9913), .ZN(n9916) );
  OR2_X1 U11026 ( .A1(n9916), .A2(n9963), .ZN(n9917) );
  OAI211_X1 U11027 ( .C1(n9919), .C2(n9971), .A(n9918), .B(n9917), .ZN(n9920)
         );
  INV_X1 U11028 ( .A(n9920), .ZN(n9921) );
  OAI211_X1 U11029 ( .C1(n9977), .C2(n9923), .A(n9922), .B(n9921), .ZN(
        P2_U3195) );
  AOI22_X1 U11030 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3151), .B1(n9957), 
        .B2(P2_ADDR_REG_14__SCAN_IN), .ZN(n9939) );
  AOI21_X1 U11031 ( .B1(n9925), .B2(n9924), .A(n4544), .ZN(n9936) );
  OAI21_X1 U11032 ( .B1(n9928), .B2(n9927), .A(n9926), .ZN(n9929) );
  NAND2_X1 U11033 ( .A1(n9929), .A2(n9967), .ZN(n9935) );
  AOI21_X1 U11034 ( .B1(n9932), .B2(n9931), .A(n9930), .ZN(n9933) );
  OR2_X1 U11035 ( .A1(n9933), .A2(n9963), .ZN(n9934) );
  OAI211_X1 U11036 ( .C1(n9936), .C2(n9971), .A(n9935), .B(n9934), .ZN(n9937)
         );
  INV_X1 U11037 ( .A(n9937), .ZN(n9938) );
  OAI211_X1 U11038 ( .C1(n9977), .C2(n9940), .A(n9939), .B(n9938), .ZN(
        P2_U3196) );
  AOI22_X1 U11039 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3151), .B1(n9957), 
        .B2(P2_ADDR_REG_16__SCAN_IN), .ZN(n9955) );
  AOI21_X1 U11040 ( .B1(n4559), .B2(n9942), .A(n9941), .ZN(n9952) );
  AOI21_X1 U11041 ( .B1(n4560), .B2(n9944), .A(n9943), .ZN(n9945) );
  OR2_X1 U11042 ( .A1(n9945), .A2(n9963), .ZN(n9951) );
  OAI21_X1 U11043 ( .B1(n9948), .B2(n9947), .A(n9946), .ZN(n9949) );
  NAND2_X1 U11044 ( .A1(n9949), .A2(n9967), .ZN(n9950) );
  OAI211_X1 U11045 ( .C1(n9952), .C2(n9971), .A(n9951), .B(n9950), .ZN(n9953)
         );
  INV_X1 U11046 ( .A(n9953), .ZN(n9954) );
  OAI211_X1 U11047 ( .C1(n9977), .C2(n9956), .A(n9955), .B(n9954), .ZN(
        P2_U3198) );
  AOI22_X1 U11048 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3151), .B1(n9957), 
        .B2(P2_ADDR_REG_17__SCAN_IN), .ZN(n9975) );
  AOI21_X1 U11049 ( .B1(n9960), .B2(n9959), .A(n9958), .ZN(n9972) );
  OAI21_X1 U11050 ( .B1(n9966), .B2(n9965), .A(n9964), .ZN(n9968) );
  NAND2_X1 U11051 ( .A1(n9968), .A2(n9967), .ZN(n9969) );
  OAI211_X1 U11052 ( .C1(n9972), .C2(n9971), .A(n9970), .B(n9969), .ZN(n9973)
         );
  INV_X1 U11053 ( .A(n9973), .ZN(n9974) );
  OAI211_X1 U11054 ( .C1(n9977), .C2(n9976), .A(n9975), .B(n9974), .ZN(
        P2_U3199) );
  INV_X1 U11055 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9982) );
  INV_X1 U11056 ( .A(n9978), .ZN(n9981) );
  NAND2_X1 U11057 ( .A1(n10064), .A2(n9979), .ZN(n9980) );
  AOI222_X1 U11058 ( .A1(n9981), .A2(n9980), .B1(n5191), .B2(n10060), .C1(
        n5870), .C2(n10042), .ZN(n10071) );
  AOI22_X1 U11059 ( .A1(n10070), .A2(n9982), .B1(n10071), .B2(n10068), .ZN(
        P2_U3390) );
  AOI21_X1 U11060 ( .B1(n10055), .B2(n9988), .A(n9983), .ZN(n9987) );
  AOI22_X1 U11061 ( .A1(n9998), .A2(n10042), .B1(n5868), .B2(n10060), .ZN(
        n9984) );
  OAI211_X1 U11062 ( .C1(n5721), .C2(n10027), .A(n9985), .B(n9984), .ZN(n9986)
         );
  NOR2_X1 U11063 ( .A1(n9987), .A2(n9986), .ZN(n10072) );
  AOI22_X1 U11064 ( .A1(n10070), .A2(n5176), .B1(n10072), .B2(n10068), .ZN(
        P2_U3393) );
  INV_X1 U11065 ( .A(n9988), .ZN(n10053) );
  INV_X1 U11066 ( .A(n9993), .ZN(n9995) );
  OAI22_X1 U11067 ( .A1(n5005), .A2(n10027), .B1(n9989), .B2(n10062), .ZN(
        n9991) );
  AOI211_X1 U11068 ( .C1(n10042), .C2(n10008), .A(n9991), .B(n9990), .ZN(n9992) );
  OAI21_X1 U11069 ( .B1(n10055), .B2(n9993), .A(n9992), .ZN(n9994) );
  AOI21_X1 U11070 ( .B1(n10053), .B2(n9995), .A(n9994), .ZN(n10074) );
  AOI22_X1 U11071 ( .A1(n10070), .A2(n5205), .B1(n10074), .B2(n10068), .ZN(
        P2_U3396) );
  INV_X1 U11072 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10004) );
  NAND2_X1 U11073 ( .A1(n9996), .A2(n10019), .ZN(n10000) );
  AOI22_X1 U11074 ( .A1(n9998), .A2(n10043), .B1(n9997), .B2(n10060), .ZN(
        n9999) );
  OAI211_X1 U11075 ( .C1(n10001), .C2(n10025), .A(n10000), .B(n9999), .ZN(
        n10002) );
  AOI21_X1 U11076 ( .B1(n10005), .B2(n10003), .A(n10002), .ZN(n10076) );
  AOI22_X1 U11077 ( .A1(n10070), .A2(n10004), .B1(n10076), .B2(n10068), .ZN(
        P2_U3399) );
  NAND2_X1 U11078 ( .A1(n10006), .A2(n10005), .ZN(n10010) );
  AOI22_X1 U11079 ( .A1(n10008), .A2(n10043), .B1(n10060), .B2(n10007), .ZN(
        n10009) );
  OAI211_X1 U11080 ( .C1(n10011), .C2(n10025), .A(n10010), .B(n10009), .ZN(
        n10012) );
  AOI21_X1 U11081 ( .B1(n10013), .B2(n10019), .A(n10012), .ZN(n10078) );
  AOI22_X1 U11082 ( .A1(n10070), .A2(n5234), .B1(n10078), .B2(n10068), .ZN(
        P2_U3402) );
  INV_X1 U11083 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10018) );
  OAI22_X1 U11084 ( .A1(n10015), .A2(n10055), .B1(n10014), .B2(n10062), .ZN(
        n10016) );
  NOR2_X1 U11085 ( .A1(n10017), .A2(n10016), .ZN(n10079) );
  AOI22_X1 U11086 ( .A1(n10070), .A2(n10018), .B1(n10079), .B2(n10068), .ZN(
        P2_U3405) );
  AND2_X1 U11087 ( .A1(n10020), .A2(n10019), .ZN(n10024) );
  AND2_X1 U11088 ( .A1(n10021), .A2(n10060), .ZN(n10022) );
  NOR3_X1 U11089 ( .A1(n10024), .A2(n10023), .A3(n10022), .ZN(n10080) );
  AOI22_X1 U11090 ( .A1(n10070), .A2(n5294), .B1(n10080), .B2(n10068), .ZN(
        P2_U3408) );
  INV_X1 U11091 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10036) );
  OAI22_X1 U11092 ( .A1(n10028), .A2(n10027), .B1(n10026), .B2(n10025), .ZN(
        n10029) );
  AOI21_X1 U11093 ( .B1(n10060), .B2(n10030), .A(n10029), .ZN(n10031) );
  OAI21_X1 U11094 ( .B1(n10032), .B2(n10055), .A(n10031), .ZN(n10034) );
  AOI211_X1 U11095 ( .C1(n10053), .C2(n10035), .A(n10034), .B(n10033), .ZN(
        n10081) );
  AOI22_X1 U11096 ( .A1(n10070), .A2(n10036), .B1(n10081), .B2(n10068), .ZN(
        P2_U3411) );
  OAI22_X1 U11097 ( .A1(n10038), .A2(n10064), .B1(n10037), .B2(n10062), .ZN(
        n10039) );
  NOR2_X1 U11098 ( .A1(n10040), .A2(n10039), .ZN(n10082) );
  AOI22_X1 U11099 ( .A1(n10070), .A2(n5329), .B1(n10082), .B2(n10068), .ZN(
        P2_U3414) );
  INV_X1 U11100 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10054) );
  INV_X1 U11101 ( .A(n10048), .ZN(n10052) );
  AOI22_X1 U11102 ( .A1(n10044), .A2(n10043), .B1(n10042), .B2(n10041), .ZN(
        n10047) );
  NAND2_X1 U11103 ( .A1(n10045), .A2(n10060), .ZN(n10046) );
  OAI211_X1 U11104 ( .C1(n10048), .C2(n10055), .A(n10047), .B(n10046), .ZN(
        n10051) );
  INV_X1 U11105 ( .A(n10049), .ZN(n10050) );
  AOI211_X1 U11106 ( .C1(n10053), .C2(n10052), .A(n10051), .B(n10050), .ZN(
        n10083) );
  AOI22_X1 U11107 ( .A1(n10070), .A2(n10054), .B1(n10083), .B2(n10068), .ZN(
        P2_U3417) );
  INV_X1 U11108 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10061) );
  NOR2_X1 U11109 ( .A1(n10056), .A2(n10055), .ZN(n10058) );
  AOI211_X1 U11110 ( .C1(n10060), .C2(n10059), .A(n10058), .B(n10057), .ZN(
        n10084) );
  AOI22_X1 U11111 ( .A1(n10070), .A2(n10061), .B1(n10084), .B2(n10068), .ZN(
        P2_U3420) );
  INV_X1 U11112 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10069) );
  OAI22_X1 U11113 ( .A1(n10065), .A2(n10064), .B1(n10063), .B2(n10062), .ZN(
        n10066) );
  NOR2_X1 U11114 ( .A1(n10067), .A2(n10066), .ZN(n10086) );
  AOI22_X1 U11115 ( .A1(n10070), .A2(n10069), .B1(n10086), .B2(n10068), .ZN(
        P2_U3423) );
  AOI22_X1 U11116 ( .A1(n10087), .A2(n10071), .B1(n5183), .B2(n10085), .ZN(
        P2_U3459) );
  AOI22_X1 U11117 ( .A1(n10087), .A2(n10072), .B1(n6155), .B2(n10085), .ZN(
        P2_U3460) );
  INV_X1 U11118 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10073) );
  AOI22_X1 U11119 ( .A1(n10087), .A2(n10074), .B1(n10073), .B2(n10085), .ZN(
        P2_U3461) );
  INV_X1 U11120 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10075) );
  AOI22_X1 U11121 ( .A1(n10087), .A2(n10076), .B1(n10075), .B2(n10085), .ZN(
        P2_U3462) );
  INV_X1 U11122 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10077) );
  AOI22_X1 U11123 ( .A1(n10087), .A2(n10078), .B1(n10077), .B2(n10085), .ZN(
        P2_U3463) );
  AOI22_X1 U11124 ( .A1(n10087), .A2(n10079), .B1(n6259), .B2(n10085), .ZN(
        P2_U3464) );
  AOI22_X1 U11125 ( .A1(n10087), .A2(n10080), .B1(n6348), .B2(n10085), .ZN(
        P2_U3465) );
  AOI22_X1 U11126 ( .A1(n10087), .A2(n10081), .B1(n6499), .B2(n10085), .ZN(
        P2_U3466) );
  AOI22_X1 U11127 ( .A1(n10087), .A2(n10082), .B1(n6808), .B2(n10085), .ZN(
        P2_U3467) );
  AOI22_X1 U11128 ( .A1(n10087), .A2(n10083), .B1(n5352), .B2(n10085), .ZN(
        P2_U3468) );
  AOI22_X1 U11129 ( .A1(n10087), .A2(n10084), .B1(n5373), .B2(n10085), .ZN(
        P2_U3469) );
  AOI22_X1 U11130 ( .A1(n10087), .A2(n10086), .B1(n5387), .B2(n10085), .ZN(
        P2_U3470) );
  NAND3_X1 U11131 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10090) );
  AND2_X1 U11132 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n10088) );
  NOR2_X1 U11133 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n10088), .ZN(n10089) );
  INV_X1 U11134 ( .A(n10089), .ZN(n10106) );
  NAND2_X1 U11135 ( .A1(n10091), .A2(n10090), .ZN(n10105) );
  OAI222_X1 U11136 ( .A1(n10091), .A2(n10090), .B1(n10091), .B2(n10106), .C1(
        n10089), .C2(n10105), .ZN(ADD_1068_U5) );
  XOR2_X1 U11137 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11138 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10092) );
  AOI21_X1 U11139 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10092), .ZN(n10117) );
  NOR2_X1 U11140 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10093) );
  AOI21_X1 U11141 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10093), .ZN(n10120) );
  NOR2_X1 U11142 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10094) );
  AOI21_X1 U11143 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10094), .ZN(n10123) );
  NOR2_X1 U11144 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10095) );
  AOI21_X1 U11145 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10095), .ZN(n10126) );
  NOR2_X1 U11146 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10096) );
  AOI21_X1 U11147 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10096), .ZN(n10129) );
  NOR2_X1 U11148 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10097) );
  AOI21_X1 U11149 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10097), .ZN(n10132) );
  NOR2_X1 U11150 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10098) );
  AOI21_X1 U11151 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10098), .ZN(n10135) );
  NOR2_X1 U11152 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10099) );
  AOI21_X1 U11153 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10099), .ZN(n10138) );
  NOR2_X1 U11154 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10100) );
  AOI21_X1 U11155 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n10100), .ZN(n10520) );
  NOR2_X1 U11156 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10101) );
  AOI21_X1 U11157 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n10101), .ZN(n10532) );
  NOR2_X1 U11158 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10102) );
  AOI21_X1 U11159 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n10102), .ZN(n10529) );
  NOR2_X1 U11160 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n10103) );
  AOI21_X1 U11161 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10103), .ZN(n10535) );
  NOR2_X1 U11162 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10104) );
  AOI21_X1 U11163 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10104), .ZN(n10526) );
  NAND2_X1 U11164 ( .A1(n10106), .A2(n10105), .ZN(n10523) );
  NAND2_X1 U11165 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10107) );
  OAI21_X1 U11166 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10107), .ZN(n10522) );
  NOR2_X1 U11167 ( .A1(n10523), .A2(n10522), .ZN(n10521) );
  AOI21_X1 U11168 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10521), .ZN(n10538) );
  NAND2_X1 U11169 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10108) );
  OAI21_X1 U11170 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10108), .ZN(n10537) );
  NOR2_X1 U11171 ( .A1(n10538), .A2(n10537), .ZN(n10536) );
  AOI21_X1 U11172 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10536), .ZN(n10541) );
  NOR2_X1 U11173 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10109) );
  AOI21_X1 U11174 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n10109), .ZN(n10540) );
  NAND2_X1 U11175 ( .A1(n10541), .A2(n10540), .ZN(n10539) );
  OAI21_X1 U11176 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10539), .ZN(n10525) );
  NAND2_X1 U11177 ( .A1(n10526), .A2(n10525), .ZN(n10524) );
  OAI21_X1 U11178 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10524), .ZN(n10534) );
  NAND2_X1 U11179 ( .A1(n10535), .A2(n10534), .ZN(n10533) );
  OAI21_X1 U11180 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n10533), .ZN(n10528) );
  NAND2_X1 U11181 ( .A1(n10529), .A2(n10528), .ZN(n10527) );
  OAI21_X1 U11182 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10527), .ZN(n10531) );
  NAND2_X1 U11183 ( .A1(n10532), .A2(n10531), .ZN(n10530) );
  OAI21_X1 U11184 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10530), .ZN(n10519) );
  NAND2_X1 U11185 ( .A1(n10520), .A2(n10519), .ZN(n10518) );
  OAI21_X1 U11186 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10518), .ZN(n10137) );
  NAND2_X1 U11187 ( .A1(n10138), .A2(n10137), .ZN(n10136) );
  OAI21_X1 U11188 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10136), .ZN(n10134) );
  NAND2_X1 U11189 ( .A1(n10135), .A2(n10134), .ZN(n10133) );
  OAI21_X1 U11190 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10133), .ZN(n10131) );
  NAND2_X1 U11191 ( .A1(n10132), .A2(n10131), .ZN(n10130) );
  OAI21_X1 U11192 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10130), .ZN(n10128) );
  NAND2_X1 U11193 ( .A1(n10129), .A2(n10128), .ZN(n10127) );
  OAI21_X1 U11194 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10127), .ZN(n10125) );
  NAND2_X1 U11195 ( .A1(n10126), .A2(n10125), .ZN(n10124) );
  OAI21_X1 U11196 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10124), .ZN(n10122) );
  NAND2_X1 U11197 ( .A1(n10123), .A2(n10122), .ZN(n10121) );
  OAI21_X1 U11198 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10121), .ZN(n10119) );
  NAND2_X1 U11199 ( .A1(n10120), .A2(n10119), .ZN(n10118) );
  OAI21_X1 U11200 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10118), .ZN(n10116) );
  NAND2_X1 U11201 ( .A1(n10117), .A2(n10116), .ZN(n10115) );
  OAI21_X1 U11202 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10115), .ZN(n10110) );
  OR2_X1 U11203 ( .A1(n10111), .A2(n10110), .ZN(n10113) );
  NAND2_X1 U11204 ( .A1(n10111), .A2(n10110), .ZN(n10511) );
  INV_X1 U11205 ( .A(n10511), .ZN(n10112) );
  NAND2_X1 U11206 ( .A1(n10114), .A2(n10113), .ZN(n10512) );
  OAI222_X1 U11207 ( .A1(n10114), .A2(n10113), .B1(n10114), .B2(n10511), .C1(
        n10112), .C2(n10512), .ZN(ADD_1068_U55) );
  OAI21_X1 U11208 ( .B1(n10117), .B2(n10116), .A(n10115), .ZN(ADD_1068_U56) );
  OAI21_X1 U11209 ( .B1(n10120), .B2(n10119), .A(n10118), .ZN(ADD_1068_U57) );
  OAI21_X1 U11210 ( .B1(n10123), .B2(n10122), .A(n10121), .ZN(ADD_1068_U58) );
  OAI21_X1 U11211 ( .B1(n10126), .B2(n10125), .A(n10124), .ZN(ADD_1068_U59) );
  OAI21_X1 U11212 ( .B1(n10129), .B2(n10128), .A(n10127), .ZN(ADD_1068_U60) );
  OAI21_X1 U11213 ( .B1(n10132), .B2(n10131), .A(n10130), .ZN(ADD_1068_U61) );
  OAI21_X1 U11214 ( .B1(n10135), .B2(n10134), .A(n10133), .ZN(ADD_1068_U62) );
  OAI21_X1 U11215 ( .B1(n10138), .B2(n10137), .A(n10136), .ZN(ADD_1068_U63) );
  OAI22_X1 U11216 ( .A1(SI_16_), .A2(keyinput_g16), .B1(keyinput_g50), .B2(
        P2_REG3_REG_17__SCAN_IN), .ZN(n10139) );
  AOI221_X1 U11217 ( .B1(SI_16_), .B2(keyinput_g16), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput_g50), .A(n10139), .ZN(n10147)
         );
  OAI22_X1 U11218 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(keyinput_g86), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .ZN(n10140) );
  AOI221_X1 U11219 ( .B1(P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_g86), .C1(
        keyinput_g36), .C2(P2_REG3_REG_27__SCAN_IN), .A(n10140), .ZN(n10146)
         );
  OAI22_X1 U11220 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput_g91), .B1(
        keyinput_g14), .B2(SI_18_), .ZN(n10142) );
  AOI221_X1 U11221 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput_g91), .C1(SI_18_), 
        .C2(keyinput_g14), .A(n10142), .ZN(n10145) );
  OAI22_X1 U11222 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(keyinput_g106), .B1(
        keyinput_g123), .B2(P1_D_REG_1__SCAN_IN), .ZN(n10143) );
  AOI221_X1 U11223 ( .B1(P1_IR_REG_16__SCAN_IN), .B2(keyinput_g106), .C1(
        P1_D_REG_1__SCAN_IN), .C2(keyinput_g123), .A(n10143), .ZN(n10144) );
  NAND4_X1 U11224 ( .A1(n10147), .A2(n10146), .A3(n10145), .A4(n10144), .ZN(
        n10175) );
  OAI22_X1 U11225 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(keyinput_g101), .B1(
        P1_IR_REG_4__SCAN_IN), .B2(keyinput_g94), .ZN(n10148) );
  AOI221_X1 U11226 ( .B1(P1_IR_REG_11__SCAN_IN), .B2(keyinput_g101), .C1(
        keyinput_g94), .C2(P1_IR_REG_4__SCAN_IN), .A(n10148), .ZN(n10155) );
  OAI22_X1 U11227 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput_g99), .B1(
        keyinput_g63), .B2(P2_REG3_REG_15__SCAN_IN), .ZN(n10149) );
  AOI221_X1 U11228 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput_g99), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput_g63), .A(n10149), .ZN(n10154)
         );
  OAI22_X1 U11229 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(keyinput_g100), .B1(
        P1_IR_REG_3__SCAN_IN), .B2(keyinput_g93), .ZN(n10150) );
  AOI221_X1 U11230 ( .B1(P1_IR_REG_10__SCAN_IN), .B2(keyinput_g100), .C1(
        keyinput_g93), .C2(P1_IR_REG_3__SCAN_IN), .A(n10150), .ZN(n10153) );
  OAI22_X1 U11231 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(keyinput_g85), .B1(
        keyinput_g61), .B2(P2_REG3_REG_6__SCAN_IN), .ZN(n10151) );
  AOI221_X1 U11232 ( .B1(P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_g85), .C1(
        P2_REG3_REG_6__SCAN_IN), .C2(keyinput_g61), .A(n10151), .ZN(n10152) );
  NAND4_X1 U11233 ( .A1(n10155), .A2(n10154), .A3(n10153), .A4(n10152), .ZN(
        n10174) );
  OAI22_X1 U11234 ( .A1(P1_D_REG_0__SCAN_IN), .A2(keyinput_g122), .B1(SI_12_), 
        .B2(keyinput_g20), .ZN(n10156) );
  AOI221_X1 U11235 ( .B1(P1_D_REG_0__SCAN_IN), .B2(keyinput_g122), .C1(
        keyinput_g20), .C2(SI_12_), .A(n10156), .ZN(n10163) );
  OAI22_X1 U11236 ( .A1(SI_21_), .A2(keyinput_g11), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .ZN(n10157) );
  AOI221_X1 U11237 ( .B1(SI_21_), .B2(keyinput_g11), .C1(keyinput_g57), .C2(
        P2_REG3_REG_22__SCAN_IN), .A(n10157), .ZN(n10162) );
  OAI22_X1 U11238 ( .A1(SI_2_), .A2(keyinput_g30), .B1(keyinput_g56), .B2(
        P2_REG3_REG_13__SCAN_IN), .ZN(n10158) );
  AOI221_X1 U11239 ( .B1(SI_2_), .B2(keyinput_g30), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput_g56), .A(n10158), .ZN(n10161)
         );
  OAI22_X1 U11240 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(keyinput_g71), .B1(
        keyinput_g65), .B2(P2_DATAO_REG_31__SCAN_IN), .ZN(n10159) );
  AOI221_X1 U11241 ( .B1(P2_DATAO_REG_25__SCAN_IN), .B2(keyinput_g71), .C1(
        P2_DATAO_REG_31__SCAN_IN), .C2(keyinput_g65), .A(n10159), .ZN(n10160)
         );
  NAND4_X1 U11242 ( .A1(n10163), .A2(n10162), .A3(n10161), .A4(n10160), .ZN(
        n10173) );
  OAI22_X1 U11243 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(keyinput_g111), .B1(
        keyinput_g48), .B2(P2_REG3_REG_16__SCAN_IN), .ZN(n10164) );
  AOI221_X1 U11244 ( .B1(P1_IR_REG_21__SCAN_IN), .B2(keyinput_g111), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput_g48), .A(n10164), .ZN(n10171)
         );
  OAI22_X1 U11245 ( .A1(P1_D_REG_4__SCAN_IN), .A2(keyinput_g126), .B1(SI_3_), 
        .B2(keyinput_g29), .ZN(n10165) );
  AOI221_X1 U11246 ( .B1(P1_D_REG_4__SCAN_IN), .B2(keyinput_g126), .C1(
        keyinput_g29), .C2(SI_3_), .A(n10165), .ZN(n10170) );
  OAI22_X1 U11247 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(keyinput_g116), .B1(
        keyinput_g37), .B2(P2_REG3_REG_14__SCAN_IN), .ZN(n10166) );
  AOI221_X1 U11248 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(keyinput_g116), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput_g37), .A(n10166), .ZN(n10169)
         );
  OAI22_X1 U11249 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(keyinput_g114), .B1(
        keyinput_g13), .B2(SI_19_), .ZN(n10167) );
  AOI221_X1 U11250 ( .B1(P1_IR_REG_24__SCAN_IN), .B2(keyinput_g114), .C1(
        SI_19_), .C2(keyinput_g13), .A(n10167), .ZN(n10168) );
  NAND4_X1 U11251 ( .A1(n10171), .A2(n10170), .A3(n10169), .A4(n10168), .ZN(
        n10172) );
  NOR4_X1 U11252 ( .A1(n10175), .A2(n10174), .A3(n10173), .A4(n10172), .ZN(
        n10312) );
  OAI22_X1 U11253 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(keyinput_g81), .B1(
        P2_REG3_REG_23__SCAN_IN), .B2(keyinput_g38), .ZN(n10176) );
  AOI221_X1 U11254 ( .B1(P2_DATAO_REG_15__SCAN_IN), .B2(keyinput_g81), .C1(
        keyinput_g38), .C2(P2_REG3_REG_23__SCAN_IN), .A(n10176), .ZN(n10183)
         );
  OAI22_X1 U11255 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(keyinput_g70), .B1(
        keyinput_g74), .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n10177) );
  AOI221_X1 U11256 ( .B1(P2_DATAO_REG_26__SCAN_IN), .B2(keyinput_g70), .C1(
        P2_DATAO_REG_22__SCAN_IN), .C2(keyinput_g74), .A(n10177), .ZN(n10182)
         );
  OAI22_X1 U11257 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(keyinput_g92), .B1(
        keyinput_g2), .B2(SI_30_), .ZN(n10178) );
  AOI221_X1 U11258 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(keyinput_g92), .C1(SI_30_), 
        .C2(keyinput_g2), .A(n10178), .ZN(n10181) );
  OAI22_X1 U11259 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(keyinput_g121), .B1(SI_10_), .B2(keyinput_g22), .ZN(n10179) );
  AOI221_X1 U11260 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(keyinput_g121), .C1(
        keyinput_g22), .C2(SI_10_), .A(n10179), .ZN(n10180) );
  NAND4_X1 U11261 ( .A1(n10183), .A2(n10182), .A3(n10181), .A4(n10180), .ZN(
        n10310) );
  OAI22_X1 U11262 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(keyinput_g118), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_g75), .ZN(n10184) );
  AOI221_X1 U11263 ( .B1(P1_IR_REG_28__SCAN_IN), .B2(keyinput_g118), .C1(
        keyinput_g75), .C2(P2_DATAO_REG_21__SCAN_IN), .A(n10184), .ZN(n10210)
         );
  OAI22_X1 U11264 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_g60), .B1(
        keyinput_g49), .B2(P2_REG3_REG_5__SCAN_IN), .ZN(n10185) );
  AOI221_X1 U11265 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .C1(
        P2_REG3_REG_5__SCAN_IN), .C2(keyinput_g49), .A(n10185), .ZN(n10188) );
  OAI22_X1 U11266 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(keyinput_g76), .B1(
        SI_17_), .B2(keyinput_g15), .ZN(n10186) );
  AOI221_X1 U11267 ( .B1(P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_g76), .C1(
        keyinput_g15), .C2(SI_17_), .A(n10186), .ZN(n10187) );
  OAI211_X1 U11268 ( .C1(n10190), .C2(keyinput_g69), .A(n10188), .B(n10187), 
        .ZN(n10189) );
  AOI21_X1 U11269 ( .B1(n10190), .B2(keyinput_g69), .A(n10189), .ZN(n10209) );
  AOI22_X1 U11270 ( .A1(SI_7_), .A2(keyinput_g25), .B1(P1_IR_REG_14__SCAN_IN), 
        .B2(keyinput_g104), .ZN(n10191) );
  OAI221_X1 U11271 ( .B1(SI_7_), .B2(keyinput_g25), .C1(P1_IR_REG_14__SCAN_IN), 
        .C2(keyinput_g104), .A(n10191), .ZN(n10198) );
  AOI22_X1 U11272 ( .A1(SI_29_), .A2(keyinput_g3), .B1(P1_IR_REG_27__SCAN_IN), 
        .B2(keyinput_g117), .ZN(n10192) );
  OAI221_X1 U11273 ( .B1(SI_29_), .B2(keyinput_g3), .C1(P1_IR_REG_27__SCAN_IN), 
        .C2(keyinput_g117), .A(n10192), .ZN(n10197) );
  AOI22_X1 U11274 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_g44), .B1(SI_4_), 
        .B2(keyinput_g28), .ZN(n10193) );
  OAI221_X1 U11275 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .C1(SI_4_), .C2(keyinput_g28), .A(n10193), .ZN(n10196) );
  AOI22_X1 U11276 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_g58), .B1(
        P2_RD_REG_SCAN_IN), .B2(keyinput_g33), .ZN(n10194) );
  OAI221_X1 U11277 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .C1(
        P2_RD_REG_SCAN_IN), .C2(keyinput_g33), .A(n10194), .ZN(n10195) );
  NOR4_X1 U11278 ( .A1(n10198), .A2(n10197), .A3(n10196), .A4(n10195), .ZN(
        n10208) );
  AOI22_X1 U11279 ( .A1(SI_20_), .A2(keyinput_g12), .B1(P1_IR_REG_6__SCAN_IN), 
        .B2(keyinput_g96), .ZN(n10199) );
  OAI221_X1 U11280 ( .B1(SI_20_), .B2(keyinput_g12), .C1(P1_IR_REG_6__SCAN_IN), 
        .C2(keyinput_g96), .A(n10199), .ZN(n10206) );
  AOI22_X1 U11281 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(keyinput_g67), .B1(
        SI_0_), .B2(keyinput_g32), .ZN(n10200) );
  OAI221_X1 U11282 ( .B1(P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_g67), .C1(
        SI_0_), .C2(keyinput_g32), .A(n10200), .ZN(n10205) );
  AOI22_X1 U11283 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_g40), .B1(
        P2_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .ZN(n10201) );
  OAI221_X1 U11284 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_g40), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_g46), .A(n10201), .ZN(n10204)
         );
  AOI22_X1 U11285 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_g53), .B1(SI_23_), .B2(keyinput_g9), .ZN(n10202) );
  OAI221_X1 U11286 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_g53), .C1(
        SI_23_), .C2(keyinput_g9), .A(n10202), .ZN(n10203) );
  NOR4_X1 U11287 ( .A1(n10206), .A2(n10205), .A3(n10204), .A4(n10203), .ZN(
        n10207) );
  NAND4_X1 U11288 ( .A1(n10210), .A2(n10209), .A3(n10208), .A4(n10207), .ZN(
        n10309) );
  AOI22_X1 U11289 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_g0), .B1(
        P1_D_REG_2__SCAN_IN), .B2(keyinput_g124), .ZN(n10211) );
  OAI221_X1 U11290 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_g0), .C1(
        P1_D_REG_2__SCAN_IN), .C2(keyinput_g124), .A(n10211), .ZN(n10219) );
  AOI22_X1 U11291 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_g55), .B1(
        P1_IR_REG_23__SCAN_IN), .B2(keyinput_g113), .ZN(n10212) );
  OAI221_X1 U11292 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .C1(
        P1_IR_REG_23__SCAN_IN), .C2(keyinput_g113), .A(n10212), .ZN(n10218) );
  AOI22_X1 U11293 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(keyinput_g79), .B1(
        P1_IR_REG_13__SCAN_IN), .B2(keyinput_g103), .ZN(n10213) );
  OAI221_X1 U11294 ( .B1(P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_g79), .C1(
        P1_IR_REG_13__SCAN_IN), .C2(keyinput_g103), .A(n10213), .ZN(n10217) );
  XNOR2_X1 U11295 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_g95), .ZN(n10215) );
  XNOR2_X1 U11296 ( .A(SI_6_), .B(keyinput_g26), .ZN(n10214) );
  NAND2_X1 U11297 ( .A1(n10215), .A2(n10214), .ZN(n10216) );
  NOR4_X1 U11298 ( .A1(n10219), .A2(n10218), .A3(n10217), .A4(n10216), .ZN(
        n10257) );
  AOI22_X1 U11299 ( .A1(n10221), .A2(keyinput_g43), .B1(n10368), .B2(
        keyinput_g125), .ZN(n10220) );
  OAI221_X1 U11300 ( .B1(n10221), .B2(keyinput_g43), .C1(n10368), .C2(
        keyinput_g125), .A(n10220), .ZN(n10229) );
  INV_X1 U11301 ( .A(SI_9_), .ZN(n10391) );
  AOI22_X1 U11302 ( .A1(n7469), .A2(keyinput_g1), .B1(n10391), .B2(
        keyinput_g23), .ZN(n10222) );
  OAI221_X1 U11303 ( .B1(n7469), .B2(keyinput_g1), .C1(n10391), .C2(
        keyinput_g23), .A(n10222), .ZN(n10228) );
  XNOR2_X1 U11304 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_g89), .ZN(n10226)
         );
  XNOR2_X1 U11305 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_g98), .ZN(n10225) );
  XNOR2_X1 U11306 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_g108), .ZN(n10224)
         );
  XNOR2_X1 U11307 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_g88), .ZN(n10223)
         );
  NAND4_X1 U11308 ( .A1(n10226), .A2(n10225), .A3(n10224), .A4(n10223), .ZN(
        n10227) );
  NOR3_X1 U11309 ( .A1(n10229), .A2(n10228), .A3(n10227), .ZN(n10256) );
  AOI22_X1 U11310 ( .A1(n5069), .A2(keyinput_g107), .B1(keyinput_g97), .B2(
        n6041), .ZN(n10230) );
  OAI221_X1 U11311 ( .B1(n5069), .B2(keyinput_g107), .C1(n6041), .C2(
        keyinput_g97), .A(n10230), .ZN(n10241) );
  INV_X1 U11312 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n10232) );
  AOI22_X1 U11313 ( .A1(n10232), .A2(keyinput_g112), .B1(keyinput_g80), .B2(
        n10420), .ZN(n10231) );
  OAI221_X1 U11314 ( .B1(n10232), .B2(keyinput_g112), .C1(n10420), .C2(
        keyinput_g80), .A(n10231), .ZN(n10240) );
  AOI22_X1 U11315 ( .A1(n10235), .A2(keyinput_g78), .B1(keyinput_g82), .B2(
        n10234), .ZN(n10233) );
  OAI221_X1 U11316 ( .B1(n10235), .B2(keyinput_g78), .C1(n10234), .C2(
        keyinput_g82), .A(n10233), .ZN(n10239) );
  XNOR2_X1 U11317 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_g102), .ZN(n10237)
         );
  XNOR2_X1 U11318 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput_g41), .ZN(n10236)
         );
  NAND2_X1 U11319 ( .A1(n10237), .A2(n10236), .ZN(n10238) );
  NOR4_X1 U11320 ( .A1(n10241), .A2(n10240), .A3(n10239), .A4(n10238), .ZN(
        n10255) );
  AOI22_X1 U11321 ( .A1(n10243), .A2(keyinput_g7), .B1(keyinput_g35), .B2(
        n5314), .ZN(n10242) );
  OAI221_X1 U11322 ( .B1(n10243), .B2(keyinput_g7), .C1(n5314), .C2(
        keyinput_g35), .A(n10242), .ZN(n10253) );
  INV_X1 U11323 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10407) );
  AOI22_X1 U11324 ( .A1(n10452), .A2(keyinput_g83), .B1(keyinput_g62), .B2(
        n10407), .ZN(n10244) );
  OAI221_X1 U11325 ( .B1(n10452), .B2(keyinput_g83), .C1(n10407), .C2(
        keyinput_g62), .A(n10244), .ZN(n10252) );
  AOI22_X1 U11326 ( .A1(n10247), .A2(keyinput_g77), .B1(keyinput_g19), .B2(
        n10246), .ZN(n10245) );
  OAI221_X1 U11327 ( .B1(n10247), .B2(keyinput_g77), .C1(n10246), .C2(
        keyinput_g19), .A(n10245), .ZN(n10251) );
  XNOR2_X1 U11328 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_g72), .ZN(n10249) );
  XNOR2_X1 U11329 ( .A(SI_1_), .B(keyinput_g31), .ZN(n10248) );
  NAND2_X1 U11330 ( .A1(n10249), .A2(n10248), .ZN(n10250) );
  NOR4_X1 U11331 ( .A1(n10253), .A2(n10252), .A3(n10251), .A4(n10250), .ZN(
        n10254) );
  NAND4_X1 U11332 ( .A1(n10257), .A2(n10256), .A3(n10255), .A4(n10254), .ZN(
        n10308) );
  AOI22_X1 U11333 ( .A1(n10260), .A2(keyinput_g10), .B1(keyinput_g84), .B2(
        n10259), .ZN(n10258) );
  OAI221_X1 U11334 ( .B1(n10260), .B2(keyinput_g10), .C1(n10259), .C2(
        keyinput_g84), .A(n10258), .ZN(n10269) );
  XNOR2_X1 U11335 ( .A(n10261), .B(keyinput_g109), .ZN(n10268) );
  XNOR2_X1 U11336 ( .A(SI_5_), .B(keyinput_g27), .ZN(n10265) );
  XNOR2_X1 U11337 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_g52), .ZN(n10264)
         );
  XNOR2_X1 U11338 ( .A(SI_8_), .B(keyinput_g24), .ZN(n10263) );
  XNOR2_X1 U11339 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_g90), .ZN(n10262) );
  NAND4_X1 U11340 ( .A1(n10265), .A2(n10264), .A3(n10263), .A4(n10262), .ZN(
        n10267) );
  XNOR2_X1 U11341 ( .A(keyinput_g120), .B(n9786), .ZN(n10266) );
  NOR4_X1 U11342 ( .A1(n10269), .A2(n10268), .A3(n10267), .A4(n10266), .ZN(
        n10306) );
  AOI22_X1 U11343 ( .A1(n5642), .A2(keyinput_g47), .B1(keyinput_g51), .B2(
        n10479), .ZN(n10270) );
  OAI221_X1 U11344 ( .B1(n5642), .B2(keyinput_g47), .C1(n10479), .C2(
        keyinput_g51), .A(n10270), .ZN(n10279) );
  AOI22_X1 U11345 ( .A1(n7494), .A2(keyinput_g73), .B1(keyinput_g66), .B2(
        n10448), .ZN(n10271) );
  OAI221_X1 U11346 ( .B1(n7494), .B2(keyinput_g73), .C1(n10448), .C2(
        keyinput_g66), .A(n10271), .ZN(n10278) );
  INV_X1 U11347 ( .A(P2_B_REG_SCAN_IN), .ZN(n10273) );
  AOI22_X1 U11348 ( .A1(n10273), .A2(keyinput_g64), .B1(n10419), .B2(
        keyinput_g6), .ZN(n10272) );
  OAI221_X1 U11349 ( .B1(n10273), .B2(keyinput_g64), .C1(n10419), .C2(
        keyinput_g6), .A(n10272), .ZN(n10277) );
  XNOR2_X1 U11350 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_g87), .ZN(n10275)
         );
  XNOR2_X1 U11351 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_g59), .ZN(n10274)
         );
  NAND2_X1 U11352 ( .A1(n10275), .A2(n10274), .ZN(n10276) );
  NOR4_X1 U11353 ( .A1(n10279), .A2(n10278), .A3(n10277), .A4(n10276), .ZN(
        n10305) );
  INV_X1 U11354 ( .A(SI_14_), .ZN(n10281) );
  AOI22_X1 U11355 ( .A1(n10281), .A2(keyinput_g18), .B1(n10429), .B2(
        keyinput_g127), .ZN(n10280) );
  OAI221_X1 U11356 ( .B1(n10281), .B2(keyinput_g18), .C1(n10429), .C2(
        keyinput_g127), .A(n10280), .ZN(n10291) );
  INV_X1 U11357 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n10283) );
  AOI22_X1 U11358 ( .A1(n10406), .A2(keyinput_g5), .B1(n10283), .B2(
        keyinput_g105), .ZN(n10282) );
  OAI221_X1 U11359 ( .B1(n10406), .B2(keyinput_g5), .C1(n10283), .C2(
        keyinput_g105), .A(n10282), .ZN(n10290) );
  AOI22_X1 U11360 ( .A1(n5474), .A2(keyinput_g17), .B1(keyinput_g68), .B2(
        n10285), .ZN(n10284) );
  OAI221_X1 U11361 ( .B1(n5474), .B2(keyinput_g17), .C1(n10285), .C2(
        keyinput_g68), .A(n10284), .ZN(n10289) );
  XOR2_X1 U11362 ( .A(n6717), .B(keyinput_g54), .Z(n10287) );
  XNOR2_X1 U11363 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_g115), .ZN(n10286)
         );
  NAND2_X1 U11364 ( .A1(n10287), .A2(n10286), .ZN(n10288) );
  NOR4_X1 U11365 ( .A1(n10291), .A2(n10290), .A3(n10289), .A4(n10288), .ZN(
        n10304) );
  AOI22_X1 U11366 ( .A1(n10293), .A2(keyinput_g8), .B1(keyinput_g45), .B2(
        n5566), .ZN(n10292) );
  OAI221_X1 U11367 ( .B1(n10293), .B2(keyinput_g8), .C1(n5566), .C2(
        keyinput_g45), .A(n10292), .ZN(n10302) );
  INV_X1 U11368 ( .A(SI_11_), .ZN(n10430) );
  AOI22_X1 U11369 ( .A1(P2_U3151), .A2(keyinput_g34), .B1(n10430), .B2(
        keyinput_g21), .ZN(n10294) );
  OAI221_X1 U11370 ( .B1(P2_U3151), .B2(keyinput_g34), .C1(n10430), .C2(
        keyinput_g21), .A(n10294), .ZN(n10301) );
  XNOR2_X1 U11371 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_g39), .ZN(n10299)
         );
  XNOR2_X1 U11372 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_g119), .ZN(n10298)
         );
  XNOR2_X1 U11373 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_g110), .ZN(n10297)
         );
  XNOR2_X1 U11374 ( .A(SI_28_), .B(keyinput_g4), .ZN(n10296) );
  NAND4_X1 U11375 ( .A1(n10299), .A2(n10298), .A3(n10297), .A4(n10296), .ZN(
        n10300) );
  NOR3_X1 U11376 ( .A1(n10302), .A2(n10301), .A3(n10300), .ZN(n10303) );
  NAND4_X1 U11377 ( .A1(n10306), .A2(n10305), .A3(n10304), .A4(n10303), .ZN(
        n10307) );
  NOR4_X1 U11378 ( .A1(n10310), .A2(n10309), .A3(n10308), .A4(n10307), .ZN(
        n10311) );
  AOI22_X1 U11379 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_g42), .B1(
        n10312), .B2(n10311), .ZN(n10510) );
  OAI22_X1 U11380 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput_f91), .B1(
        keyinput_f106), .B2(P1_IR_REG_16__SCAN_IN), .ZN(n10313) );
  AOI221_X1 U11381 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput_f91), .C1(
        P1_IR_REG_16__SCAN_IN), .C2(keyinput_f106), .A(n10313), .ZN(n10320) );
  OAI22_X1 U11382 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(keyinput_f72), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_f67), .ZN(n10314) );
  AOI221_X1 U11383 ( .B1(P2_DATAO_REG_24__SCAN_IN), .B2(keyinput_f72), .C1(
        keyinput_f67), .C2(P2_DATAO_REG_29__SCAN_IN), .A(n10314), .ZN(n10319)
         );
  OAI22_X1 U11384 ( .A1(SI_2_), .A2(keyinput_f30), .B1(keyinput_f4), .B2(
        SI_28_), .ZN(n10315) );
  AOI221_X1 U11385 ( .B1(SI_2_), .B2(keyinput_f30), .C1(SI_28_), .C2(
        keyinput_f4), .A(n10315), .ZN(n10318) );
  OAI22_X1 U11386 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput_f93), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(keyinput_f54), .ZN(n10316) );
  AOI221_X1 U11387 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput_f93), .C1(
        keyinput_f54), .C2(P2_REG3_REG_0__SCAN_IN), .A(n10316), .ZN(n10317) );
  NAND4_X1 U11388 ( .A1(n10320), .A2(n10319), .A3(n10318), .A4(n10317), .ZN(
        n10353) );
  OAI22_X1 U11389 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(keyinput_f117), .B1(SI_31_), .B2(keyinput_f1), .ZN(n10321) );
  AOI221_X1 U11390 ( .B1(P1_IR_REG_27__SCAN_IN), .B2(keyinput_f117), .C1(
        keyinput_f1), .C2(SI_31_), .A(n10321), .ZN(n10328) );
  OAI22_X1 U11391 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(keyinput_f115), .B1(
        keyinput_f68), .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n10322) );
  AOI221_X1 U11392 ( .B1(P1_IR_REG_25__SCAN_IN), .B2(keyinput_f115), .C1(
        P2_DATAO_REG_28__SCAN_IN), .C2(keyinput_f68), .A(n10322), .ZN(n10327)
         );
  OAI22_X1 U11393 ( .A1(P1_D_REG_2__SCAN_IN), .A2(keyinput_f124), .B1(
        keyinput_f10), .B2(SI_22_), .ZN(n10323) );
  AOI221_X1 U11394 ( .B1(P1_D_REG_2__SCAN_IN), .B2(keyinput_f124), .C1(SI_22_), 
        .C2(keyinput_f10), .A(n10323), .ZN(n10326) );
  OAI22_X1 U11395 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(keyinput_f120), .B1(
        keyinput_f48), .B2(P2_REG3_REG_16__SCAN_IN), .ZN(n10324) );
  AOI221_X1 U11396 ( .B1(P1_IR_REG_30__SCAN_IN), .B2(keyinput_f120), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput_f48), .A(n10324), .ZN(n10325)
         );
  NAND4_X1 U11397 ( .A1(n10328), .A2(n10327), .A3(n10326), .A4(n10325), .ZN(
        n10352) );
  OAI22_X1 U11398 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(keyinput_f96), .B1(
        keyinput_f89), .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n10329) );
  AOI221_X1 U11399 ( .B1(P1_IR_REG_6__SCAN_IN), .B2(keyinput_f96), .C1(
        P2_DATAO_REG_7__SCAN_IN), .C2(keyinput_f89), .A(n10329), .ZN(n10336)
         );
  OAI22_X1 U11400 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(keyinput_f108), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_f79), .ZN(n10330) );
  AOI221_X1 U11401 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(keyinput_f108), .C1(
        keyinput_f79), .C2(P2_DATAO_REG_17__SCAN_IN), .A(n10330), .ZN(n10335)
         );
  OAI22_X1 U11402 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(keyinput_f105), .B1(
        keyinput_f29), .B2(SI_3_), .ZN(n10331) );
  AOI221_X1 U11403 ( .B1(P1_IR_REG_15__SCAN_IN), .B2(keyinput_f105), .C1(SI_3_), .C2(keyinput_f29), .A(n10331), .ZN(n10334) );
  OAI22_X1 U11404 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(keyinput_f113), .B1(
        keyinput_f19), .B2(SI_13_), .ZN(n10332) );
  AOI221_X1 U11405 ( .B1(P1_IR_REG_23__SCAN_IN), .B2(keyinput_f113), .C1(
        SI_13_), .C2(keyinput_f19), .A(n10332), .ZN(n10333) );
  NAND4_X1 U11406 ( .A1(n10336), .A2(n10335), .A3(n10334), .A4(n10333), .ZN(
        n10351) );
  OAI22_X1 U11407 ( .A1(n10338), .A2(keyinput_f26), .B1(n5566), .B2(
        keyinput_f45), .ZN(n10337) );
  AOI221_X1 U11408 ( .B1(n10338), .B2(keyinput_f26), .C1(keyinput_f45), .C2(
        n5566), .A(n10337), .ZN(n10349) );
  OAI22_X1 U11409 ( .A1(n10340), .A2(keyinput_f58), .B1(keyinput_f33), .B2(
        P2_RD_REG_SCAN_IN), .ZN(n10339) );
  AOI221_X1 U11410 ( .B1(n10340), .B2(keyinput_f58), .C1(P2_RD_REG_SCAN_IN), 
        .C2(keyinput_f33), .A(n10339), .ZN(n10348) );
  OAI22_X1 U11411 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(keyinput_f104), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(keyinput_f74), .ZN(n10341) );
  AOI221_X1 U11412 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput_f104), .C1(
        keyinput_f74), .C2(P2_DATAO_REG_22__SCAN_IN), .A(n10341), .ZN(n10347)
         );
  XNOR2_X1 U11413 ( .A(n10342), .B(keyinput_f114), .ZN(n10345) );
  XNOR2_X1 U11414 ( .A(n10343), .B(keyinput_f31), .ZN(n10344) );
  NOR2_X1 U11415 ( .A1(n10345), .A2(n10344), .ZN(n10346) );
  NAND4_X1 U11416 ( .A1(n10349), .A2(n10348), .A3(n10347), .A4(n10346), .ZN(
        n10350) );
  NOR4_X1 U11417 ( .A1(n10353), .A2(n10352), .A3(n10351), .A4(n10350), .ZN(
        n10507) );
  OAI22_X1 U11418 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput_f87), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .ZN(n10354) );
  AOI221_X1 U11419 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_f87), .C1(
        keyinput_f63), .C2(P2_REG3_REG_15__SCAN_IN), .A(n10354), .ZN(n10361)
         );
  OAI22_X1 U11420 ( .A1(SI_20_), .A2(keyinput_f12), .B1(P2_B_REG_SCAN_IN), 
        .B2(keyinput_f64), .ZN(n10355) );
  AOI221_X1 U11421 ( .B1(SI_20_), .B2(keyinput_f12), .C1(keyinput_f64), .C2(
        P2_B_REG_SCAN_IN), .A(n10355), .ZN(n10360) );
  OAI22_X1 U11422 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput_f109), .B1(
        keyinput_f18), .B2(SI_14_), .ZN(n10356) );
  AOI221_X1 U11423 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(keyinput_f109), .C1(
        SI_14_), .C2(keyinput_f18), .A(n10356), .ZN(n10359) );
  OAI22_X1 U11424 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_f50), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .ZN(n10357) );
  AOI221_X1 U11425 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_f50), .C1(
        keyinput_f44), .C2(P2_REG3_REG_1__SCAN_IN), .A(n10357), .ZN(n10358) );
  NAND4_X1 U11426 ( .A1(n10361), .A2(n10360), .A3(n10359), .A4(n10358), .ZN(
        n10505) );
  OAI22_X1 U11427 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(keyinput_f86), .B1(
        keyinput_f119), .B2(P1_IR_REG_29__SCAN_IN), .ZN(n10362) );
  AOI221_X1 U11428 ( .B1(P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_f86), .C1(
        P1_IR_REG_29__SCAN_IN), .C2(keyinput_f119), .A(n10362), .ZN(n10388) );
  OAI22_X1 U11429 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_f36), .B1(
        P2_REG3_REG_20__SCAN_IN), .B2(keyinput_f55), .ZN(n10363) );
  AOI221_X1 U11430 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .C1(
        keyinput_f55), .C2(P2_REG3_REG_20__SCAN_IN), .A(n10363), .ZN(n10366)
         );
  OAI22_X1 U11431 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(keyinput_f84), .B1(
        keyinput_f85), .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n10364) );
  AOI221_X1 U11432 ( .B1(P2_DATAO_REG_12__SCAN_IN), .B2(keyinput_f84), .C1(
        P2_DATAO_REG_11__SCAN_IN), .C2(keyinput_f85), .A(n10364), .ZN(n10365)
         );
  OAI211_X1 U11433 ( .C1(n10368), .C2(keyinput_f125), .A(n10366), .B(n10365), 
        .ZN(n10367) );
  AOI21_X1 U11434 ( .B1(n10368), .B2(keyinput_f125), .A(n10367), .ZN(n10387)
         );
  AOI22_X1 U11435 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(keyinput_f70), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_f69), .ZN(n10369) );
  OAI221_X1 U11436 ( .B1(P2_DATAO_REG_26__SCAN_IN), .B2(keyinput_f70), .C1(
        P2_DATAO_REG_27__SCAN_IN), .C2(keyinput_f69), .A(n10369), .ZN(n10376)
         );
  AOI22_X1 U11437 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_f43), .B1(
        P1_D_REG_1__SCAN_IN), .B2(keyinput_f123), .ZN(n10370) );
  OAI221_X1 U11438 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .C1(
        P1_D_REG_1__SCAN_IN), .C2(keyinput_f123), .A(n10370), .ZN(n10375) );
  AOI22_X1 U11439 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(keyinput_f82), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(keyinput_f81), .ZN(n10371) );
  OAI221_X1 U11440 ( .B1(P2_DATAO_REG_14__SCAN_IN), .B2(keyinput_f82), .C1(
        P2_DATAO_REG_15__SCAN_IN), .C2(keyinput_f81), .A(n10371), .ZN(n10374)
         );
  AOI22_X1 U11441 ( .A1(SI_7_), .A2(keyinput_f25), .B1(P1_IR_REG_20__SCAN_IN), 
        .B2(keyinput_f110), .ZN(n10372) );
  OAI221_X1 U11442 ( .B1(SI_7_), .B2(keyinput_f25), .C1(P1_IR_REG_20__SCAN_IN), 
        .C2(keyinput_f110), .A(n10372), .ZN(n10373) );
  NOR4_X1 U11443 ( .A1(n10376), .A2(n10375), .A3(n10374), .A4(n10373), .ZN(
        n10386) );
  AOI22_X1 U11444 ( .A1(SI_12_), .A2(keyinput_f20), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_f76), .ZN(n10377) );
  OAI221_X1 U11445 ( .B1(SI_12_), .B2(keyinput_f20), .C1(
        P2_DATAO_REG_20__SCAN_IN), .C2(keyinput_f76), .A(n10377), .ZN(n10384)
         );
  AOI22_X1 U11446 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_f34), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(keyinput_f73), .ZN(n10378) );
  OAI221_X1 U11447 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_f34), .C1(
        P2_DATAO_REG_23__SCAN_IN), .C2(keyinput_f73), .A(n10378), .ZN(n10383)
         );
  AOI22_X1 U11448 ( .A1(SI_29_), .A2(keyinput_f3), .B1(P1_IR_REG_22__SCAN_IN), 
        .B2(keyinput_f112), .ZN(n10379) );
  OAI221_X1 U11449 ( .B1(SI_29_), .B2(keyinput_f3), .C1(P1_IR_REG_22__SCAN_IN), 
        .C2(keyinput_f112), .A(n10379), .ZN(n10382) );
  AOI22_X1 U11450 ( .A1(SI_25_), .A2(keyinput_f7), .B1(P1_IR_REG_4__SCAN_IN), 
        .B2(keyinput_f94), .ZN(n10380) );
  OAI221_X1 U11451 ( .B1(SI_25_), .B2(keyinput_f7), .C1(P1_IR_REG_4__SCAN_IN), 
        .C2(keyinput_f94), .A(n10380), .ZN(n10381) );
  NOR4_X1 U11452 ( .A1(n10384), .A2(n10383), .A3(n10382), .A4(n10381), .ZN(
        n10385) );
  NAND4_X1 U11453 ( .A1(n10388), .A2(n10387), .A3(n10386), .A4(n10385), .ZN(
        n10504) );
  INV_X1 U11454 ( .A(SI_21_), .ZN(n10390) );
  AOI22_X1 U11455 ( .A1(n10391), .A2(keyinput_f23), .B1(n10390), .B2(
        keyinput_f11), .ZN(n10389) );
  OAI221_X1 U11456 ( .B1(n10391), .B2(keyinput_f23), .C1(n10390), .C2(
        keyinput_f11), .A(n10389), .ZN(n10402) );
  INV_X1 U11457 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10393) );
  AOI22_X1 U11458 ( .A1(n10394), .A2(keyinput_f13), .B1(keyinput_f56), .B2(
        n10393), .ZN(n10392) );
  OAI221_X1 U11459 ( .B1(n10394), .B2(keyinput_f13), .C1(n10393), .C2(
        keyinput_f56), .A(n10392), .ZN(n10401) );
  AOI22_X1 U11460 ( .A1(n10397), .A2(keyinput_f39), .B1(n10396), .B2(
        keyinput_f37), .ZN(n10395) );
  OAI221_X1 U11461 ( .B1(n10397), .B2(keyinput_f39), .C1(n10396), .C2(
        keyinput_f37), .A(n10395), .ZN(n10400) );
  AOI22_X1 U11462 ( .A1(n5837), .A2(keyinput_f92), .B1(keyinput_f53), .B2(
        n5348), .ZN(n10398) );
  OAI221_X1 U11463 ( .B1(n5837), .B2(keyinput_f92), .C1(n5348), .C2(
        keyinput_f53), .A(n10398), .ZN(n10399) );
  NOR4_X1 U11464 ( .A1(n10402), .A2(n10401), .A3(n10400), .A4(n10399), .ZN(
        n10444) );
  AOI22_X1 U11465 ( .A1(n10404), .A2(keyinput_f49), .B1(n5314), .B2(
        keyinput_f35), .ZN(n10403) );
  OAI221_X1 U11466 ( .B1(n10404), .B2(keyinput_f49), .C1(n5314), .C2(
        keyinput_f35), .A(n10403), .ZN(n10414) );
  AOI22_X1 U11467 ( .A1(n10407), .A2(keyinput_f62), .B1(n10406), .B2(
        keyinput_f5), .ZN(n10405) );
  OAI221_X1 U11468 ( .B1(n10407), .B2(keyinput_f62), .C1(n10406), .C2(
        keyinput_f5), .A(n10405), .ZN(n10413) );
  XOR2_X1 U11469 ( .A(n5642), .B(keyinput_f47), .Z(n10411) );
  XNOR2_X1 U11470 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_f59), .ZN(n10410)
         );
  XNOR2_X1 U11471 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_f98), .ZN(n10409) );
  XNOR2_X1 U11472 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_f102), .ZN(n10408)
         );
  NAND4_X1 U11473 ( .A1(n10411), .A2(n10410), .A3(n10409), .A4(n10408), .ZN(
        n10412) );
  NOR3_X1 U11474 ( .A1(n10414), .A2(n10413), .A3(n10412), .ZN(n10443) );
  AOI22_X1 U11475 ( .A1(n10417), .A2(keyinput_f24), .B1(n10416), .B2(
        keyinput_f75), .ZN(n10415) );
  OAI221_X1 U11476 ( .B1(n10417), .B2(keyinput_f24), .C1(n10416), .C2(
        keyinput_f75), .A(n10415), .ZN(n10427) );
  AOI22_X1 U11477 ( .A1(n10420), .A2(keyinput_f80), .B1(n10419), .B2(
        keyinput_f6), .ZN(n10418) );
  OAI221_X1 U11478 ( .B1(n10420), .B2(keyinput_f80), .C1(n10419), .C2(
        keyinput_f6), .A(n10418), .ZN(n10426) );
  XOR2_X1 U11479 ( .A(n5514), .B(keyinput_f14), .Z(n10424) );
  XNOR2_X1 U11480 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_f52), .ZN(n10423)
         );
  XNOR2_X1 U11481 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_f77), .ZN(n10422) );
  XNOR2_X1 U11482 ( .A(SI_5_), .B(keyinput_f27), .ZN(n10421) );
  NAND4_X1 U11483 ( .A1(n10424), .A2(n10423), .A3(n10422), .A4(n10421), .ZN(
        n10425) );
  NOR3_X1 U11484 ( .A1(n10427), .A2(n10426), .A3(n10425), .ZN(n10442) );
  AOI22_X1 U11485 ( .A1(n10430), .A2(keyinput_f21), .B1(n10429), .B2(
        keyinput_f127), .ZN(n10428) );
  OAI221_X1 U11486 ( .B1(n10430), .B2(keyinput_f21), .C1(n10429), .C2(
        keyinput_f127), .A(n10428), .ZN(n10440) );
  AOI22_X1 U11487 ( .A1(n5948), .A2(keyinput_f118), .B1(n6041), .B2(
        keyinput_f97), .ZN(n10431) );
  OAI221_X1 U11488 ( .B1(n5948), .B2(keyinput_f118), .C1(n6041), .C2(
        keyinput_f97), .A(n10431), .ZN(n10439) );
  AOI22_X1 U11489 ( .A1(n10434), .A2(keyinput_f15), .B1(n10433), .B2(
        keyinput_f122), .ZN(n10432) );
  OAI221_X1 U11490 ( .B1(n10434), .B2(keyinput_f15), .C1(n10433), .C2(
        keyinput_f122), .A(n10432), .ZN(n10438) );
  XOR2_X1 U11491 ( .A(n5848), .B(keyinput_f116), .Z(n10436) );
  XNOR2_X1 U11492 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_f121), .ZN(n10435)
         );
  NAND2_X1 U11493 ( .A1(n10436), .A2(n10435), .ZN(n10437) );
  NOR4_X1 U11494 ( .A1(n10440), .A2(n10439), .A3(n10438), .A4(n10437), .ZN(
        n10441) );
  NAND4_X1 U11495 ( .A1(n10444), .A2(n10443), .A3(n10442), .A4(n10441), .ZN(
        n10503) );
  AOI22_X1 U11496 ( .A1(n5474), .A2(keyinput_f17), .B1(keyinput_f65), .B2(
        n10446), .ZN(n10445) );
  OAI221_X1 U11497 ( .B1(n5474), .B2(keyinput_f17), .C1(n10446), .C2(
        keyinput_f65), .A(n10445), .ZN(n10458) );
  AOI22_X1 U11498 ( .A1(n10448), .A2(keyinput_f66), .B1(n5069), .B2(
        keyinput_f107), .ZN(n10447) );
  OAI221_X1 U11499 ( .B1(n10448), .B2(keyinput_f66), .C1(n5069), .C2(
        keyinput_f107), .A(n10447), .ZN(n10457) );
  INV_X1 U11500 ( .A(SI_0_), .ZN(n10450) );
  AOI22_X1 U11501 ( .A1(n10451), .A2(keyinput_f22), .B1(keyinput_f32), .B2(
        n10450), .ZN(n10449) );
  OAI221_X1 U11502 ( .B1(n10451), .B2(keyinput_f22), .C1(n10450), .C2(
        keyinput_f32), .A(n10449), .ZN(n10456) );
  XOR2_X1 U11503 ( .A(n10452), .B(keyinput_f83), .Z(n10454) );
  XNOR2_X1 U11504 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_f95), .ZN(n10453) );
  NAND2_X1 U11505 ( .A1(n10454), .A2(n10453), .ZN(n10455) );
  NOR4_X1 U11506 ( .A1(n10458), .A2(n10457), .A3(n10456), .A4(n10455), .ZN(
        n10501) );
  INV_X1 U11507 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10460) );
  AOI22_X1 U11508 ( .A1(n10460), .A2(keyinput_f38), .B1(n5840), .B2(
        keyinput_f101), .ZN(n10459) );
  OAI221_X1 U11509 ( .B1(n10460), .B2(keyinput_f38), .C1(n5840), .C2(
        keyinput_f101), .A(n10459), .ZN(n10470) );
  INV_X1 U11510 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10462) );
  AOI22_X1 U11511 ( .A1(n10463), .A2(keyinput_f41), .B1(n10462), .B2(
        keyinput_f57), .ZN(n10461) );
  OAI221_X1 U11512 ( .B1(n10463), .B2(keyinput_f41), .C1(n10462), .C2(
        keyinput_f57), .A(n10461), .ZN(n10469) );
  XNOR2_X1 U11513 ( .A(SI_24_), .B(keyinput_f8), .ZN(n10467) );
  XNOR2_X1 U11514 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_f40), .ZN(n10466)
         );
  XNOR2_X1 U11515 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_f99), .ZN(n10465) );
  XNOR2_X1 U11516 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_f78), .ZN(n10464) );
  NAND4_X1 U11517 ( .A1(n10467), .A2(n10466), .A3(n10465), .A4(n10464), .ZN(
        n10468) );
  NOR3_X1 U11518 ( .A1(n10470), .A2(n10469), .A3(n10468), .ZN(n10500) );
  INV_X1 U11519 ( .A(keyinput_f0), .ZN(n10472) );
  AOI22_X1 U11520 ( .A1(n10473), .A2(keyinput_f9), .B1(P2_WR_REG_SCAN_IN), 
        .B2(n10472), .ZN(n10471) );
  OAI221_X1 U11521 ( .B1(n10473), .B2(keyinput_f9), .C1(n10472), .C2(
        P2_WR_REG_SCAN_IN), .A(n10471), .ZN(n10485) );
  AOI22_X1 U11522 ( .A1(n10476), .A2(keyinput_f46), .B1(n10475), .B2(
        keyinput_f60), .ZN(n10474) );
  OAI221_X1 U11523 ( .B1(n10476), .B2(keyinput_f46), .C1(n10475), .C2(
        keyinput_f60), .A(n10474), .ZN(n10484) );
  AOI22_X1 U11524 ( .A1(n10479), .A2(keyinput_f51), .B1(n10478), .B2(
        keyinput_f88), .ZN(n10477) );
  OAI221_X1 U11525 ( .B1(n10479), .B2(keyinput_f51), .C1(n10478), .C2(
        keyinput_f88), .A(n10477), .ZN(n10483) );
  XNOR2_X1 U11526 ( .A(SI_4_), .B(keyinput_f28), .ZN(n10481) );
  XNOR2_X1 U11527 ( .A(SI_16_), .B(keyinput_f16), .ZN(n10480) );
  NAND2_X1 U11528 ( .A1(n10481), .A2(n10480), .ZN(n10482) );
  NOR4_X1 U11529 ( .A1(n10485), .A2(n10484), .A3(n10483), .A4(n10482), .ZN(
        n10499) );
  AOI22_X1 U11530 ( .A1(n5855), .A2(keyinput_f111), .B1(keyinput_f126), .B2(
        n10487), .ZN(n10486) );
  OAI221_X1 U11531 ( .B1(n5855), .B2(keyinput_f111), .C1(n10487), .C2(
        keyinput_f126), .A(n10486), .ZN(n10497) );
  INV_X1 U11532 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n10490) );
  AOI22_X1 U11533 ( .A1(n10490), .A2(keyinput_f100), .B1(keyinput_f71), .B2(
        n10489), .ZN(n10488) );
  OAI221_X1 U11534 ( .B1(n10490), .B2(keyinput_f100), .C1(n10489), .C2(
        keyinput_f71), .A(n10488), .ZN(n10496) );
  XNOR2_X1 U11535 ( .A(SI_30_), .B(keyinput_f2), .ZN(n10494) );
  XNOR2_X1 U11536 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_f103), .ZN(n10493)
         );
  XNOR2_X1 U11537 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_f90), .ZN(n10492) );
  XNOR2_X1 U11538 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_f61), .ZN(n10491)
         );
  NAND4_X1 U11539 ( .A1(n10494), .A2(n10493), .A3(n10492), .A4(n10491), .ZN(
        n10495) );
  NOR3_X1 U11540 ( .A1(n10497), .A2(n10496), .A3(n10495), .ZN(n10498) );
  NAND4_X1 U11541 ( .A1(n10501), .A2(n10500), .A3(n10499), .A4(n10498), .ZN(
        n10502) );
  NOR4_X1 U11542 ( .A1(n10505), .A2(n10504), .A3(n10503), .A4(n10502), .ZN(
        n10506) );
  AOI22_X1 U11543 ( .A1(n10507), .A2(n10506), .B1(keyinput_f42), .B2(
        P2_REG3_REG_28__SCAN_IN), .ZN(n10508) );
  OAI21_X1 U11544 ( .B1(keyinput_f42), .B2(P2_REG3_REG_28__SCAN_IN), .A(n10508), .ZN(n10509) );
  OAI211_X1 U11545 ( .C1(P2_REG3_REG_28__SCAN_IN), .C2(keyinput_g42), .A(
        n10510), .B(n10509), .ZN(n10517) );
  NAND2_X1 U11546 ( .A1(n10512), .A2(n10511), .ZN(n10515) );
  XNOR2_X1 U11547 ( .A(n10513), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n10514) );
  XNOR2_X1 U11548 ( .A(n10515), .B(n10514), .ZN(n10516) );
  XNOR2_X1 U11549 ( .A(n10517), .B(n10516), .ZN(ADD_1068_U4) );
  OAI21_X1 U11550 ( .B1(n10520), .B2(n10519), .A(n10518), .ZN(ADD_1068_U47) );
  AOI21_X1 U11551 ( .B1(n10523), .B2(n10522), .A(n10521), .ZN(ADD_1068_U54) );
  OAI21_X1 U11552 ( .B1(n10526), .B2(n10525), .A(n10524), .ZN(ADD_1068_U51) );
  OAI21_X1 U11553 ( .B1(n10529), .B2(n10528), .A(n10527), .ZN(ADD_1068_U49) );
  OAI21_X1 U11554 ( .B1(n10532), .B2(n10531), .A(n10530), .ZN(ADD_1068_U48) );
  OAI21_X1 U11555 ( .B1(n10535), .B2(n10534), .A(n10533), .ZN(ADD_1068_U50) );
  AOI21_X1 U11556 ( .B1(n10538), .B2(n10537), .A(n10536), .ZN(ADD_1068_U53) );
  OAI21_X1 U11557 ( .B1(n10541), .B2(n10540), .A(n10539), .ZN(ADD_1068_U52) );
  BUF_X1 U5076 ( .A(n5212), .Z(n6625) );
  OR2_X1 U5055 ( .A1(n7183), .A2(n5394), .ZN(n5395) );
  CLKBUF_X1 U5074 ( .A(n7933), .Z(n4602) );
  CLKBUF_X2 U5246 ( .A(n5214), .Z(n6628) );
endmodule

