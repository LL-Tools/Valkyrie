

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput63, keyinput62, keyinput61, 
        keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, 
        keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, 
        keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, 
        keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, 
        keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, 
        keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, 
        keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, 
        keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, 
        keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, 
        keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, 
        keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput63, keyinput62,
         keyinput61, keyinput60, keyinput59, keyinput58, keyinput57,
         keyinput56, keyinput55, keyinput54, keyinput53, keyinput52,
         keyinput51, keyinput50, keyinput49, keyinput48, keyinput47,
         keyinput46, keyinput45, keyinput44, keyinput43, keyinput42,
         keyinput41, keyinput40, keyinput39, keyinput38, keyinput37,
         keyinput36, keyinput35, keyinput34, keyinput33, keyinput32,
         keyinput31, keyinput30, keyinput29, keyinput28, keyinput27,
         keyinput26, keyinput25, keyinput24, keyinput23, keyinput22,
         keyinput21, keyinput20, keyinput19, keyinput18, keyinput17,
         keyinput16, keyinput15, keyinput14, keyinput13, keyinput12,
         keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6,
         keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740;

  CLKBUF_X1 U3410 ( .A(n4011), .Z(n4025) );
  CLKBUF_X2 U3411 ( .A(n3262), .Z(n4141) );
  CLKBUF_X2 U3412 ( .A(n3161), .Z(n4214) );
  CLKBUF_X2 U3413 ( .A(n3228), .Z(n4664) );
  CLKBUF_X2 U3414 ( .A(n3166), .Z(n4224) );
  CLKBUF_X2 U3415 ( .A(n3646), .Z(n4225) );
  CLKBUF_X2 U3416 ( .A(n3953), .Z(n4628) );
  NOR2_X1 U3417 ( .A1(n3205), .A2(n3282), .ZN(n3285) );
  NAND2_X1 U3418 ( .A1(n2967), .A2(n3183), .ZN(n3205) );
  AND4_X1 U3419 ( .A1(n3077), .A2(n3076), .A3(n3075), .A4(n3074), .ZN(n3194)
         );
  AND4_X1 U3420 ( .A1(n3046), .A2(n3045), .A3(n3044), .A4(n3043), .ZN(n3176)
         );
  AND4_X1 U3421 ( .A1(n3049), .A2(n3050), .A3(n3048), .A4(n3047), .ZN(n3174)
         );
  NOR2_X2 U3423 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4667) );
  AND4_X1 U3424 ( .A1(n3177), .A2(n3176), .A3(n3175), .A4(n3174), .ZN(n3178)
         );
  OAI21_X1 U3425 ( .B1(n3284), .B2(n3186), .A(n5171), .ZN(n3207) );
  AND2_X2 U3426 ( .A1(n3010), .A2(n4662), .ZN(n3247) );
  AND4_X1 U3427 ( .A1(n3042), .A2(n3041), .A3(n3040), .A4(n3039), .ZN(n3175)
         );
  NAND2_X1 U3429 ( .A1(n4813), .A2(n3192), .ZN(n5174) );
  BUF_X1 U3430 ( .A(n3560), .Z(n4726) );
  AND2_X1 U3431 ( .A1(n3132), .A2(n3131), .ZN(n4606) );
  AND2_X1 U3432 ( .A1(n5556), .A2(n6616), .ZN(n6160) );
  NAND2_X1 U3433 ( .A1(n2991), .A2(n5494), .ZN(n5525) );
  INV_X1 U3434 ( .A(n6160), .ZN(n6146) );
  NAND2_X1 U3435 ( .A1(n5668), .A2(n4756), .ZN(n5935) );
  NOR2_X1 U3437 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n2995) );
  AND2_X2 U3438 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4670) );
  OR2_X2 U3440 ( .A1(n4878), .A2(n4959), .ZN(n5039) );
  NAND2_X2 U3441 ( .A1(n2971), .A2(n2972), .ZN(n3195) );
  NAND2_X2 U3442 ( .A1(n3305), .A2(n3304), .ZN(n2970) );
  NAND2_X2 U3443 ( .A1(n3485), .A2(n3484), .ZN(n5193) );
  XNOR2_X1 U34460 ( .A(n3408), .B(n3409), .ZN(n3390) );
  AND2_X2 U34470 ( .A1(n3924), .A2(n4628), .ZN(n4518) );
  INV_X2 U34480 ( .A(n4557), .ZN(n2962) );
  CLKBUF_X2 U3449 ( .A(n3188), .Z(n4802) );
  INV_X1 U3450 ( .A(n3194), .ZN(n3956) );
  INV_X1 U34510 ( .A(n2973), .ZN(n3204) );
  INV_X1 U34520 ( .A(n3179), .ZN(n2963) );
  NAND4_X2 U34530 ( .A1(n3018), .A2(n3017), .A3(n3016), .A4(n3015), .ZN(n3189)
         );
  CLKBUF_X2 U3454 ( .A(n3263), .Z(n4215) );
  CLKBUF_X2 U34550 ( .A(n4218), .Z(n3661) );
  BUF_X1 U34560 ( .A(n4439), .Z(n5698) );
  OR2_X1 U3457 ( .A1(n4289), .A2(n4288), .ZN(n4290) );
  CLKBUF_X1 U3458 ( .A(n3920), .Z(n4289) );
  CLKBUF_X1 U34590 ( .A(n3526), .Z(n5701) );
  OAI22_X1 U34600 ( .A1(n5931), .A2(n5935), .B1(n5930), .B2(n5929), .ZN(n5932)
         );
  OAI21_X1 U34610 ( .B1(n4438), .B2(n4437), .A(n5627), .ZN(n5635) );
  AND2_X1 U34620 ( .A1(n4480), .A2(n4479), .ZN(n5579) );
  CLKBUF_X2 U34630 ( .A(n4477), .Z(n4480) );
  AND2_X1 U34640 ( .A1(n2975), .A2(n2976), .ZN(n4477) );
  AND2_X1 U34650 ( .A1(n5598), .A2(n3868), .ZN(n4455) );
  NOR2_X1 U3466 ( .A1(n5597), .A2(n5601), .ZN(n5598) );
  CLKBUF_X1 U3467 ( .A(n5650), .Z(n5651) );
  NAND2_X1 U34680 ( .A1(n3767), .A2(n3766), .ZN(n5512) );
  AOI211_X1 U34690 ( .C1(n4294), .C2(n6330), .A(n5554), .B(n4293), .ZN(n4298)
         );
  CLKBUF_X1 U34700 ( .A(n5036), .Z(n5160) );
  INV_X1 U34710 ( .A(n4874), .ZN(n3640) );
  INV_X4 U34720 ( .A(n4451), .ZN(n5848) );
  NOR2_X1 U34730 ( .A1(n5637), .A2(n5638), .ZN(n4069) );
  OR2_X1 U34740 ( .A1(n3508), .A2(n3458), .ZN(n3519) );
  XNOR2_X1 U3475 ( .A(n3468), .B(n3467), .ZN(n3528) );
  XNOR2_X1 U3476 ( .A(n3452), .B(n4845), .ZN(n4838) );
  NAND2_X1 U3477 ( .A1(n3387), .A2(n3455), .ZN(n3468) );
  OAI21_X2 U3478 ( .B1(n3566), .B2(n3458), .A(n3439), .ZN(n3440) );
  OR2_X1 U3479 ( .A1(n3566), .A2(n3711), .ZN(n3576) );
  INV_X1 U3480 ( .A(n3457), .ZN(n3387) );
  OAI21_X1 U3481 ( .B1(n4726), .B2(n3711), .A(n3565), .ZN(n4548) );
  BUF_X1 U3482 ( .A(n3405), .Z(n3425) );
  INV_X1 U3483 ( .A(n4704), .ZN(n3350) );
  NAND2_X1 U3484 ( .A1(n4594), .A2(n3550), .ZN(n4554) );
  AND2_X1 U3485 ( .A1(n3349), .A2(n3348), .ZN(n4704) );
  XNOR2_X1 U3486 ( .A(n3390), .B(n3389), .ZN(n4701) );
  AND2_X1 U3487 ( .A1(n3301), .A2(n3389), .ZN(n3407) );
  AND2_X1 U3488 ( .A1(n4760), .A2(n4759), .ZN(n4880) );
  NAND2_X1 U3489 ( .A1(n3300), .A2(n3299), .ZN(n3389) );
  CLKBUF_X1 U3490 ( .A(n4595), .Z(n6163) );
  NAND2_X1 U3491 ( .A1(n3227), .A2(n6615), .ZN(n3401) );
  CLKBUF_X1 U3492 ( .A(n3544), .Z(n5540) );
  NAND2_X1 U3493 ( .A1(n3296), .A2(n3226), .ZN(n3544) );
  BUF_X1 U3494 ( .A(n3303), .Z(n3296) );
  NAND2_X1 U3495 ( .A1(n3333), .A2(n3332), .ZN(n6391) );
  INV_X1 U3496 ( .A(n2965), .ZN(n3328) );
  CLKBUF_X1 U3497 ( .A(n3951), .Z(n4748) );
  CLKBUF_X1 U3498 ( .A(n3924), .Z(n4599) );
  AND2_X1 U3499 ( .A1(n3279), .A2(n3278), .ZN(n3924) );
  AND2_X1 U3500 ( .A1(n3191), .A2(n4596), .ZN(n3210) );
  NOR2_X1 U3501 ( .A1(n3257), .A2(n6615), .ZN(n3388) );
  NAND2_X1 U3502 ( .A1(n4305), .A2(n3502), .ZN(n3465) );
  INV_X2 U3503 ( .A(n3978), .ZN(n4557) );
  AND2_X2 U3504 ( .A1(n3081), .A2(n3956), .ZN(n3374) );
  AND2_X1 U3505 ( .A1(n4628), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3081) );
  OR2_X1 U3506 ( .A1(n3256), .A2(n3255), .ZN(n3392) );
  NAND2_X1 U3507 ( .A1(n3241), .A2(n2983), .ZN(n3479) );
  NOR2_X1 U3508 ( .A1(n3213), .A2(n3204), .ZN(n3280) );
  NAND2_X1 U3509 ( .A1(n2963), .A2(n3183), .ZN(n3198) );
  CLKBUF_X1 U3510 ( .A(n3195), .Z(n5533) );
  INV_X1 U3511 ( .A(n3189), .ZN(n3188) );
  NOR2_X2 U3512 ( .A1(n3189), .A2(n3953), .ZN(n5171) );
  INV_X1 U3513 ( .A(n3953), .ZN(n4813) );
  AND2_X2 U3514 ( .A1(n3160), .A2(n2978), .ZN(n2973) );
  NAND4_X2 U3515 ( .A1(n3038), .A2(n3037), .A3(n3036), .A4(n3035), .ZN(n3953)
         );
  AND4_X1 U3516 ( .A1(n3009), .A2(n3008), .A3(n3007), .A4(n3006), .ZN(n3016)
         );
  AND4_X1 U3517 ( .A1(n3069), .A2(n3068), .A3(n3067), .A4(n3066), .ZN(n3075)
         );
  AND4_X1 U3518 ( .A1(n3022), .A2(n3021), .A3(n3020), .A4(n3019), .ZN(n3038)
         );
  AND4_X1 U3519 ( .A1(n3026), .A2(n3025), .A3(n3024), .A4(n3023), .ZN(n3037)
         );
  AND4_X1 U3520 ( .A1(n3155), .A2(n3154), .A3(n3153), .A4(n3152), .ZN(n3160)
         );
  AND4_X1 U3521 ( .A1(n3073), .A2(n3072), .A3(n3071), .A4(n3070), .ZN(n3074)
         );
  AND4_X1 U3522 ( .A1(n3004), .A2(n3003), .A3(n3002), .A4(n3001), .ZN(n3017)
         );
  AND4_X1 U3523 ( .A1(n3151), .A2(n3150), .A3(n3149), .A4(n3148), .ZN(n2972)
         );
  AND4_X1 U3524 ( .A1(n3034), .A2(n3033), .A3(n3032), .A4(n3031), .ZN(n3035)
         );
  AND4_X1 U3525 ( .A1(n3030), .A2(n3029), .A3(n3028), .A4(n3027), .ZN(n3036)
         );
  AND4_X1 U3526 ( .A1(n3061), .A2(n3060), .A3(n3059), .A4(n3058), .ZN(n3077)
         );
  AND4_X1 U3527 ( .A1(n3147), .A2(n3146), .A3(n3145), .A4(n3144), .ZN(n2971)
         );
  AND4_X1 U3528 ( .A1(n2999), .A2(n2998), .A3(n2997), .A4(n2996), .ZN(n3018)
         );
  AND4_X1 U3529 ( .A1(n3065), .A2(n3064), .A3(n3063), .A4(n3062), .ZN(n3076)
         );
  AND4_X1 U3530 ( .A1(n3137), .A2(n3136), .A3(n3135), .A4(n3134), .ZN(n3143)
         );
  AND4_X1 U3531 ( .A1(n3014), .A2(n3013), .A3(n3012), .A4(n3011), .ZN(n3015)
         );
  CLKBUF_X1 U3532 ( .A(n4127), .Z(n4216) );
  CLKBUF_X1 U3533 ( .A(n3334), .Z(n3235) );
  AND2_X1 U3534 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4603) );
  INV_X2 U3535 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6615) );
  AND2_X1 U3536 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        STATE2_REG_0__SCAN_IN), .ZN(n2964) );
  NAND2_X1 U3537 ( .A1(n3201), .A2(STATE2_REG_0__SCAN_IN), .ZN(n2965) );
  AND2_X1 U3538 ( .A1(n3929), .A2(n3199), .ZN(n3208) );
  AND2_X1 U3539 ( .A1(n3197), .A2(n3196), .ZN(n3929) );
  NAND2_X1 U3540 ( .A1(n3541), .A2(n3540), .ZN(n4552) );
  AND2_X2 U3541 ( .A1(n3010), .A2(n4660), .ZN(n3341) );
  AND2_X2 U3542 ( .A1(n3005), .A2(n4603), .ZN(n3228) );
  AOI22_X1 U3543 ( .A1(n3262), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3161), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3136) );
  AND2_X2 U3544 ( .A1(n4610), .A2(n4667), .ZN(n4223) );
  NAND2_X1 U3545 ( .A1(n3968), .A2(n3221), .ZN(n3223) );
  AND2_X1 U3546 ( .A1(n3220), .A2(n3219), .ZN(n3221) );
  CLKBUF_X1 U3547 ( .A(n4719), .Z(n2966) );
  AND4_X1 U3548 ( .A1(n3077), .A2(n3076), .A3(n3075), .A4(n3074), .ZN(n2967)
         );
  AND4_X1 U3549 ( .A1(n3077), .A2(n3076), .A3(n3075), .A4(n3074), .ZN(n2968)
         );
  NAND2_X1 U3550 ( .A1(n3433), .A2(n3432), .ZN(n4719) );
  NOR2_X4 U3551 ( .A1(n5039), .A2(n5038), .ZN(n5326) );
  NOR2_X2 U3552 ( .A1(n4654), .A2(n4010), .ZN(n4760) );
  INV_X1 U3553 ( .A(n3198), .ZN(n2969) );
  NAND2_X1 U3555 ( .A1(n4303), .A2(n3187), .ZN(n3932) );
  CLKBUF_X1 U3556 ( .A(n4133), .Z(n4195) );
  NAND2_X1 U3557 ( .A1(n3442), .A2(n3441), .ZN(n4839) );
  NAND2_X1 U3558 ( .A1(n4439), .A2(n4441), .ZN(n5709) );
  NOR2_X1 U3559 ( .A1(n5597), .A2(n5601), .ZN(n2975) );
  AND2_X1 U3560 ( .A1(n4456), .A2(n3868), .ZN(n2976) );
  NAND2_X1 U3561 ( .A1(n4477), .A2(n4210), .ZN(n4300) );
  XNOR2_X1 U3562 ( .A(n4571), .B(n6391), .ZN(n4661) );
  AND2_X2 U3563 ( .A1(n4547), .A2(n4548), .ZN(n4546) );
  NAND2_X2 U3564 ( .A1(n2979), .A2(n3559), .ZN(n4547) );
  AND2_X2 U3565 ( .A1(n4576), .A2(n4649), .ZN(n4651) );
  AND2_X2 U3566 ( .A1(n4546), .A2(n4577), .ZN(n4576) );
  AND2_X2 U3567 ( .A1(n4651), .A2(n5043), .ZN(n4708) );
  NAND2_X1 U3568 ( .A1(n3682), .A2(n3681), .ZN(n5285) );
  OR2_X2 U3570 ( .A1(n4553), .A2(n3556), .ZN(n2979) );
  AND2_X2 U3571 ( .A1(n5337), .A2(n3713), .ZN(n5437) );
  AND2_X2 U3572 ( .A1(n5437), .A2(n5479), .ZN(n5478) );
  AOI21_X1 U3573 ( .B1(n4302), .B2(n4300), .A(n4301), .ZN(n5687) );
  NAND2_X1 U3574 ( .A1(n3222), .A2(n3223), .ZN(n3303) );
  INV_X1 U3575 ( .A(n4248), .ZN(n4236) );
  OR2_X1 U3576 ( .A1(n5533), .A2(n6514), .ZN(n4304) );
  INV_X1 U3577 ( .A(n4304), .ZN(n4243) );
  OR2_X1 U3578 ( .A1(n3384), .A2(n3383), .ZN(n3470) );
  NAND2_X1 U3579 ( .A1(n3457), .A2(n3445), .ZN(n3577) );
  OR2_X1 U3580 ( .A1(n3319), .A2(n3318), .ZN(n3416) );
  CLKBUF_X1 U3581 ( .A(n3339), .Z(n3340) );
  OR2_X1 U3582 ( .A1(n4628), .A2(n6615), .ZN(n3502) );
  INV_X1 U3583 ( .A(n3130), .ZN(n3120) );
  NAND2_X1 U3584 ( .A1(n3503), .A2(n3938), .ZN(n3113) );
  NAND2_X1 U3585 ( .A1(n3118), .A2(n3117), .ZN(n3125) );
  OR2_X1 U3586 ( .A1(n3116), .A2(n3115), .ZN(n3118) );
  AND2_X2 U3587 ( .A1(n4660), .A2(n4603), .ZN(n3339) );
  OR2_X1 U3588 ( .A1(n3956), .A2(n6615), .ZN(n4305) );
  AND2_X1 U3589 ( .A1(n4189), .A2(n4476), .ZN(n4479) );
  NAND2_X1 U3590 ( .A1(n3784), .A2(n3783), .ZN(n5519) );
  INV_X1 U3591 ( .A(n5521), .ZN(n3783) );
  INV_X1 U3592 ( .A(n5512), .ZN(n3784) );
  INV_X1 U3593 ( .A(n4207), .ZN(n4239) );
  NAND2_X1 U3594 ( .A1(n5848), .A2(n5967), .ZN(n3919) );
  NAND2_X1 U3595 ( .A1(n2963), .A2(n3195), .ZN(n3212) );
  NAND2_X1 U3596 ( .A1(n3203), .A2(n3202), .ZN(n3222) );
  NAND2_X1 U3597 ( .A1(n2964), .A2(n3201), .ZN(n3203) );
  AND2_X1 U3598 ( .A1(n3374), .A2(n3509), .ZN(n3130) );
  NOR2_X1 U3599 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4725), .ZN(n4768) );
  INV_X1 U3600 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6575) );
  AND2_X1 U3601 ( .A1(n4687), .A2(n4686), .ZN(n6581) );
  AND3_X1 U3602 ( .A1(n4039), .A2(n4063), .A3(n4038), .ZN(n5482) );
  NAND2_X1 U3603 ( .A1(n4752), .A2(n6273), .ZN(n5531) );
  AOI21_X1 U3604 ( .B1(n3680), .B2(n3679), .A(n3678), .ZN(n5286) );
  NOR2_X2 U3605 ( .A1(n5640), .A2(n4504), .ZN(n5590) );
  INV_X1 U3606 ( .A(n4054), .ZN(n4055) );
  OR2_X1 U3607 ( .A1(n5848), .A2(n5987), .ZN(n5501) );
  OAI21_X1 U3608 ( .B1(n4750), .B2(n3950), .A(n3949), .ZN(n4097) );
  NAND2_X1 U3609 ( .A1(n3948), .A2(n6612), .ZN(n3949) );
  OR2_X1 U3610 ( .A1(n3954), .A2(n4513), .ZN(n4749) );
  OR2_X1 U3611 ( .A1(n4980), .A2(n4702), .ZN(n4890) );
  AND2_X1 U3612 ( .A1(n6467), .A2(n4892), .ZN(n6349) );
  OR2_X1 U3613 ( .A1(n3330), .A2(n6615), .ZN(n6598) );
  NOR2_X1 U3614 ( .A1(n6693), .A2(n5587), .ZN(n5876) );
  AND2_X1 U3615 ( .A1(n4485), .A2(n6727), .ZN(n6161) );
  INV_X1 U3616 ( .A(n6158), .ZN(n6144) );
  AND2_X1 U3617 ( .A1(n6170), .A2(n4557), .ZN(n6140) );
  INV_X1 U3618 ( .A(n6140), .ZN(n6157) );
  XNOR2_X1 U3619 ( .A(n4255), .B(n4254), .ZN(n5621) );
  OAI21_X1 U3620 ( .B1(n4253), .B2(n4252), .A(n4251), .ZN(n4255) );
  INV_X1 U3621 ( .A(n4435), .ZN(n4438) );
  AND2_X1 U3622 ( .A1(n4627), .A2(n6638), .ZN(n6210) );
  INV_X1 U3623 ( .A(n5955), .ZN(n5961) );
  INV_X1 U3624 ( .A(n6016), .ZN(n6296) );
  INV_X1 U3625 ( .A(n5977), .ZN(n5030) );
  NAND2_X2 U3626 ( .A1(n3401), .A2(n3400), .ZN(n5387) );
  CLKBUF_X1 U3627 ( .A(n6389), .Z(n6513) );
  INV_X1 U3628 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6501) );
  NOR2_X1 U3629 ( .A1(n5171), .A2(n3057), .ZN(n3102) );
  AOI22_X1 U3630 ( .A1(n4133), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3228), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3151) );
  AOI22_X1 U3631 ( .A1(n4218), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3166), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3147) );
  CLKBUF_X1 U3632 ( .A(n3341), .Z(n3230) );
  OAI21_X1 U3633 ( .B1(n3503), .B2(n3386), .A(n3385), .ZN(n3455) );
  XNOR2_X1 U3634 ( .A(n3325), .B(n3324), .ZN(n3406) );
  NAND2_X1 U3635 ( .A1(n3322), .A2(n3321), .ZN(n3325) );
  AND3_X1 U3636 ( .A1(n4303), .A2(n3212), .A3(n2968), .ZN(n3185) );
  OR2_X1 U3637 ( .A1(n3347), .A2(n3346), .ZN(n3428) );
  AND2_X1 U3638 ( .A1(n4188), .A2(n4436), .ZN(n4476) );
  AND2_X1 U3639 ( .A1(n5541), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4207) );
  NAND2_X1 U3640 ( .A1(n3619), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3624)
         );
  AND2_X1 U3641 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3561), .ZN(n3572)
         );
  NAND2_X1 U3642 ( .A1(n2969), .A2(n2967), .ZN(n3197) );
  NAND2_X1 U3643 ( .A1(n3519), .A2(n3482), .ZN(n3483) );
  NAND2_X1 U3644 ( .A1(n4002), .A2(n4001), .ZN(n4654) );
  INV_X1 U3645 ( .A(n4656), .ZN(n4001) );
  INV_X1 U3646 ( .A(n4655), .ZN(n4002) );
  AND2_X2 U3647 ( .A1(n3401), .A2(n3259), .ZN(n3408) );
  AND3_X1 U3648 ( .A1(n3277), .A2(n3276), .A3(n3275), .ZN(n3409) );
  OR2_X1 U3649 ( .A1(n3969), .A2(n3715), .ZN(n3930) );
  XNOR2_X1 U3650 ( .A(n3298), .B(n3297), .ZN(n4595) );
  INV_X1 U3651 ( .A(n3296), .ZN(n3297) );
  AOI21_X1 U3652 ( .B1(n3114), .B2(n3113), .A(n3112), .ZN(n3122) );
  AND2_X1 U3653 ( .A1(n3127), .A2(n3126), .ZN(n3937) );
  AND2_X1 U3654 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6586), .ZN(n3124)
         );
  NAND2_X1 U3655 ( .A1(n3935), .A2(n4802), .ZN(n3951) );
  AND2_X1 U3656 ( .A1(n3329), .A2(n5151), .ZN(n5065) );
  AOI21_X1 U3657 ( .B1(n6603), .B2(n6619), .A(n5562), .ZN(n4725) );
  NAND2_X1 U3658 ( .A1(n4518), .A2(n4625), .ZN(n4527) );
  NAND2_X1 U3659 ( .A1(n5892), .A2(n2986), .ZN(n4266) );
  AND2_X1 U3660 ( .A1(n3881), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3883)
         );
  NAND2_X1 U3661 ( .A1(n3883), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4157)
         );
  AND2_X1 U3662 ( .A1(n4018), .A2(n4017), .ZN(n4879) );
  AND2_X1 U3663 ( .A1(n4004), .A2(n4003), .ZN(n4712) );
  NAND2_X1 U3664 ( .A1(n3536), .A2(n3535), .ZN(n4711) );
  NAND2_X1 U3665 ( .A1(n3558), .A2(n3885), .ZN(n4588) );
  NOR2_X2 U3666 ( .A1(n4300), .A2(n4302), .ZN(n4301) );
  NAND2_X1 U3667 ( .A1(n4158), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4211)
         );
  AND2_X1 U3668 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n4179), .ZN(n4178)
         );
  NAND2_X1 U3669 ( .A1(n4480), .A2(n4187), .ZN(n4435) );
  AND2_X1 U3670 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n3835), .ZN(n3836)
         );
  AND2_X1 U3671 ( .A1(n3836), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3881)
         );
  OR2_X1 U3672 ( .A1(n5728), .A2(n4248), .ZN(n3841) );
  NOR2_X1 U3673 ( .A1(n3800), .A2(n5745), .ZN(n3801) );
  NOR2_X1 U3674 ( .A1(n3762), .A2(n5490), .ZN(n3763) );
  NAND2_X1 U3675 ( .A1(n3763), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3800)
         );
  INV_X1 U3676 ( .A(n5513), .ZN(n3766) );
  INV_X1 U3677 ( .A(n5485), .ZN(n3767) );
  NAND2_X1 U3678 ( .A1(n3731), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3762)
         );
  AND2_X1 U3679 ( .A1(n3714), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3731)
         );
  NOR2_X1 U3680 ( .A1(n3697), .A2(n6058), .ZN(n3714) );
  CLKBUF_X1 U3681 ( .A(n5337), .Z(n5338) );
  NOR2_X1 U3682 ( .A1(n3674), .A2(n6081), .ZN(n3675) );
  INV_X1 U3683 ( .A(n5286), .ZN(n3681) );
  INV_X1 U3684 ( .A(n5157), .ZN(n3682) );
  OR2_X1 U3685 ( .A1(n3657), .A2(n5273), .ZN(n3674) );
  AND3_X1 U3686 ( .A1(n3607), .A2(n3606), .A3(n3605), .ZN(n4745) );
  CLKBUF_X1 U3687 ( .A(n4743), .Z(n4744) );
  INV_X1 U3688 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U3689 ( .A1(n3588), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3590)
         );
  CLKBUF_X1 U3690 ( .A(n4708), .Z(n5044) );
  NAND2_X1 U3691 ( .A1(n3572), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3579)
         );
  NAND2_X1 U3692 ( .A1(n3578), .A2(n3679), .ZN(n3584) );
  NOR2_X1 U3693 ( .A1(n6145), .A2(n3551), .ZN(n3561) );
  NAND2_X1 U3694 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4111) );
  INV_X1 U3695 ( .A(n4439), .ZN(n3921) );
  NOR2_X2 U3696 ( .A1(n5709), .A2(n4111), .ZN(n4463) );
  OR2_X1 U3697 ( .A1(n5848), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5699)
         );
  BUF_X1 U3698 ( .A(n5637), .Z(n5645) );
  AND2_X1 U3699 ( .A1(n4046), .A2(n4045), .ZN(n5523) );
  CLKBUF_X1 U3700 ( .A(n5750), .Z(n5751) );
  INV_X1 U3701 ( .A(n5482), .ZN(n4040) );
  AND2_X1 U3702 ( .A1(n4043), .A2(n4042), .ZN(n5494) );
  CLKBUF_X1 U3703 ( .A(n5754), .Z(n5755) );
  NAND3_X1 U3704 ( .A1(n5171), .A2(n3281), .A3(n3280), .ZN(n4597) );
  AND2_X1 U3705 ( .A1(n5327), .A2(n5289), .ZN(n4031) );
  NAND2_X1 U3706 ( .A1(n5848), .A2(n5320), .ZN(n3491) );
  NAND2_X1 U3707 ( .A1(n5848), .A2(n5322), .ZN(n5265) );
  AND3_X1 U3708 ( .A1(n4020), .A2(n4063), .A3(n4019), .ZN(n4959) );
  NAND2_X1 U3709 ( .A1(n3992), .A2(n3991), .ZN(n4586) );
  INV_X1 U3710 ( .A(n4584), .ZN(n3992) );
  NOR2_X2 U3711 ( .A1(n4586), .A2(n4550), .ZN(n4580) );
  AND2_X1 U3712 ( .A1(n5464), .A2(n5995), .ZN(n4867) );
  OR2_X1 U3713 ( .A1(n4867), .A2(n4618), .ZN(n6338) );
  OR2_X1 U3714 ( .A1(n4726), .A2(n3557), .ZN(n6506) );
  INV_X1 U3715 ( .A(n3935), .ZN(n4256) );
  NOR2_X1 U3716 ( .A1(n3930), .A2(n3204), .ZN(n5541) );
  CLKBUF_X1 U3717 ( .A(n4675), .Z(n5862) );
  INV_X1 U3718 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3000) );
  AND4_X1 U3719 ( .A1(n4568), .A2(n4567), .A3(n4566), .A4(n4565), .ZN(n6579)
         );
  INV_X1 U3720 ( .A(n5202), .ZN(n5210) );
  NOR2_X1 U3721 ( .A1(n6506), .A2(n4702), .ZN(n5202) );
  CLKBUF_X1 U3722 ( .A(n2963), .Z(n3529) );
  INV_X1 U3723 ( .A(n6506), .ZN(n5070) );
  OR2_X1 U3724 ( .A1(n6714), .A2(n4725), .ZN(n4951) );
  INV_X1 U3725 ( .A(n5387), .ZN(n5209) );
  NOR2_X1 U3726 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6389) );
  NOR2_X1 U3727 ( .A1(n6345), .A2(n4727), .ZN(n5119) );
  AOI21_X1 U3728 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5385), .A(n5123), .ZN(
        n6510) );
  NAND2_X1 U3729 ( .A1(n6514), .A2(n6015), .ZN(n4248) );
  AND2_X1 U3730 ( .A1(n6513), .A2(n6614), .ZN(n6007) );
  AND2_X1 U3731 ( .A1(n5874), .A2(n4278), .ZN(n5582) );
  INV_X1 U3732 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6111) );
  NOR2_X1 U3733 ( .A1(n5184), .A2(n5183), .ZN(n6126) );
  NAND2_X1 U3734 ( .A1(n4316), .A2(n4315), .ZN(n4317) );
  AND2_X1 U3735 ( .A1(n6182), .A2(n5533), .ZN(n6179) );
  AND2_X1 U3736 ( .A1(n6182), .A2(n5669), .ZN(n6178) );
  INV_X1 U3737 ( .A(n6182), .ZN(n5641) );
  NAND2_X2 U3738 ( .A1(n4310), .A2(n4309), .ZN(n6182) );
  OR2_X1 U3739 ( .A1(n4568), .A2(n6598), .ZN(n4310) );
  INV_X1 U3740 ( .A(n6179), .ZN(n5667) );
  INV_X1 U3741 ( .A(n5935), .ZN(n6191) );
  AND2_X1 U3742 ( .A1(n5668), .A2(n5534), .ZN(n6190) );
  INV_X1 U3743 ( .A(n5668), .ZN(n6193) );
  NAND2_X1 U3744 ( .A1(n5531), .A2(n4757), .ZN(n5452) );
  INV_X2 U3745 ( .A(n6199), .ZN(n6226) );
  INV_X1 U3746 ( .A(n6280), .ZN(n4658) );
  NAND2_X1 U3747 ( .A1(n4625), .A2(n4533), .ZN(n6282) );
  INV_X2 U3748 ( .A(n4658), .ZN(n6276) );
  OR2_X1 U3749 ( .A1(n4246), .A2(n4245), .ZN(n4247) );
  CLKBUF_X1 U3750 ( .A(n5471), .Z(n5472) );
  OR2_X1 U3751 ( .A1(n5824), .A2(n3977), .ZN(n5965) );
  INV_X1 U3752 ( .A(n5965), .ZN(n5782) );
  NAND2_X1 U3753 ( .A1(n5853), .A2(n4105), .ZN(n5824) );
  CLKBUF_X1 U3754 ( .A(n5821), .Z(n5822) );
  AND2_X1 U3755 ( .A1(n4102), .A2(n6306), .ZN(n5853) );
  CLKBUF_X1 U3756 ( .A(n5499), .Z(n5500) );
  NAND2_X1 U3757 ( .A1(n5817), .A2(n5994), .ZN(n6306) );
  INV_X1 U3758 ( .A(n5997), .ZN(n6336) );
  INV_X1 U3759 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5385) );
  CLKBUF_X1 U3760 ( .A(n4701), .Z(n4702) );
  CLKBUF_X1 U3761 ( .A(n4700), .Z(n6345) );
  INV_X1 U3762 ( .A(n2977), .ZN(n6467) );
  INV_X1 U3763 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6586) );
  OAI21_X1 U3764 ( .B1(n4695), .B2(n6713), .A(n5123), .ZN(n6344) );
  INV_X1 U3765 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6614) );
  AND2_X2 U3766 ( .A1(n3292), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4608)
         );
  NOR2_X1 U3767 ( .A1(n6716), .A2(n4606), .ZN(n5562) );
  INV_X1 U3768 ( .A(n5343), .ZN(n5384) );
  OAI21_X1 U3769 ( .B1(n4968), .B2(n4896), .A(n4895), .ZN(n4964) );
  INV_X1 U3770 ( .A(n5000), .ZN(n5426) );
  INV_X1 U3771 ( .A(n5211), .ZN(n5259) );
  NOR2_X1 U3772 ( .A1(n4951), .A2(n4813), .ZN(n6504) );
  NOR2_X1 U3773 ( .A1(n4951), .A2(n2973), .ZN(n6529) );
  NOR2_X1 U3774 ( .A1(n4951), .A2(n4822), .ZN(n6535) );
  NOR2_X1 U3775 ( .A1(n4951), .A2(n2967), .ZN(n6541) );
  NAND2_X1 U3776 ( .A1(n5070), .A2(n6423), .ZN(n6569) );
  NOR2_X1 U3777 ( .A1(n6253), .A2(n5123), .ZN(n6524) );
  NOR2_X1 U3778 ( .A1(n6255), .A2(n5123), .ZN(n6530) );
  NOR2_X1 U3779 ( .A1(n6257), .A2(n5123), .ZN(n6536) );
  NOR2_X1 U3780 ( .A1(n6261), .A2(n5123), .ZN(n6548) );
  NOR2_X1 U3781 ( .A1(n5047), .A2(n5123), .ZN(n6555) );
  INV_X1 U3782 ( .A(n6523), .ZN(n5431) );
  INV_X1 U3783 ( .A(n6530), .ZN(n5363) );
  INV_X1 U3784 ( .A(n6529), .ZN(n5415) );
  INV_X1 U3785 ( .A(n6536), .ZN(n5352) );
  INV_X1 U3786 ( .A(n6535), .ZN(n5403) );
  INV_X1 U3787 ( .A(n6542), .ZN(n5383) );
  INV_X1 U3788 ( .A(n6541), .ZN(n5419) );
  INV_X1 U3789 ( .A(n6548), .ZN(n5367) );
  INV_X1 U3790 ( .A(n6547), .ZN(n5423) );
  NAND2_X1 U3791 ( .A1(n5119), .A2(n5209), .ZN(n5149) );
  NAND2_X1 U3792 ( .A1(n5119), .A2(n5387), .ZN(n5150) );
  INV_X1 U3793 ( .A(n6563), .ZN(n5407) );
  AND2_X1 U3794 ( .A1(n6602), .A2(n6601), .ZN(n6621) );
  INV_X1 U3795 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6716) );
  INV_X1 U3796 ( .A(n6708), .ZN(n6740) );
  AOI21_X1 U3797 ( .B1(n5881), .B2(n5880), .A(n5879), .ZN(n5882) );
  NAND2_X1 U3798 ( .A1(n5878), .A2(n5877), .ZN(n5879) );
  NAND2_X1 U3799 ( .A1(n5876), .A2(n6695), .ZN(n5877) );
  NOR2_X1 U3800 ( .A1(n4508), .A2(n4507), .ZN(n4509) );
  INV_X1 U3801 ( .A(n4498), .ZN(n4510) );
  OAI21_X1 U3802 ( .B1(n5780), .B2(n6157), .A(n4506), .ZN(n4507) );
  OAI21_X1 U3803 ( .B1(n5955), .B2(n5588), .A(n4443), .ZN(n4444) );
  NOR2_X1 U3804 ( .A1(n4461), .A2(n4460), .ZN(n4462) );
  INV_X1 U3805 ( .A(n4459), .ZN(n4460) );
  AND2_X1 U3806 ( .A1(n4298), .A2(n4297), .ZN(n4299) );
  AND2_X1 U3807 ( .A1(n4474), .A2(n4473), .ZN(n4475) );
  AND2_X1 U3808 ( .A1(n4113), .A2(n4112), .ZN(n4114) );
  NAND2_X1 U3809 ( .A1(n3640), .A2(n3639), .ZN(n4962) );
  AND4_X1 U3810 ( .A1(n3159), .A2(n3158), .A3(n3157), .A4(n3156), .ZN(n2978)
         );
  OAI21_X1 U3811 ( .B1(n3577), .B2(n3458), .A(n3451), .ZN(n3452) );
  NAND2_X1 U3812 ( .A1(n5478), .A2(n5486), .ZN(n5485) );
  AND2_X1 U3813 ( .A1(n4284), .A2(n4283), .ZN(n2980) );
  OR2_X1 U3814 ( .A1(n6298), .A2(n3912), .ZN(n5955) );
  INV_X1 U3815 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3292) );
  INV_X1 U3816 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n2993) );
  NAND2_X1 U3817 ( .A1(n3529), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3711) );
  INV_X1 U3818 ( .A(n3711), .ZN(n3679) );
  OAI21_X1 U3819 ( .B1(n5193), .B2(n3487), .A(n3486), .ZN(n5026) );
  INV_X1 U3820 ( .A(n3212), .ZN(n3542) );
  AND2_X2 U3821 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4660) );
  INV_X1 U3822 ( .A(n4961), .ZN(n3639) );
  INV_X1 U3823 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3570) );
  NAND2_X1 U3824 ( .A1(n5936), .A2(n6288), .ZN(n4446) );
  AND2_X1 U3825 ( .A1(n5939), .A2(n6288), .ZN(n4461) );
  AND2_X1 U3826 ( .A1(n3285), .A2(n4813), .ZN(n2981) );
  INV_X1 U3827 ( .A(n4702), .ZN(n4983) );
  AND3_X1 U3828 ( .A1(n5851), .A2(n3518), .A3(n5820), .ZN(n2982) );
  NOR2_X1 U3829 ( .A1(n3240), .A2(n3239), .ZN(n2983) );
  AND4_X1 U3830 ( .A1(REIP_REG_30__SCAN_IN), .A2(REIP_REG_29__SCAN_IN), .A3(
        n5585), .A4(n6705), .ZN(n2984) );
  AND3_X1 U3831 ( .A1(n4495), .A2(n4494), .A3(n2989), .ZN(n2985) );
  AND3_X1 U3832 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .A3(
        REIP_REG_22__SCAN_IN), .ZN(n2986) );
  AND2_X1 U3833 ( .A1(n4451), .A2(n3524), .ZN(n2987) );
  INV_X1 U3834 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3551) );
  NAND2_X1 U3835 ( .A1(n5848), .A2(n5032), .ZN(n2988) );
  OR2_X1 U3836 ( .A1(n4493), .A2(REIP_REG_28__SCAN_IN), .ZN(n2989) );
  INV_X1 U3837 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6081) );
  INV_X1 U3838 ( .A(n6039), .ZN(n5880) );
  NAND2_X1 U3839 ( .A1(n3983), .A2(n3982), .ZN(n3986) );
  AND2_X1 U3840 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n2990) );
  INV_X1 U3841 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3078) );
  AND2_X1 U3842 ( .A1(n5440), .A2(n4040), .ZN(n2991) );
  INV_X1 U3843 ( .A(n6726), .ZN(n6708) );
  AND2_X1 U3844 ( .A1(n6007), .A2(n6615), .ZN(n6328) );
  INV_X1 U3846 ( .A(n5338), .ZN(n5438) );
  NAND2_X1 U3847 ( .A1(n4527), .A2(n4528), .ZN(n6727) );
  INV_X1 U3848 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3099) );
  INV_X1 U3849 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3110) );
  AND2_X2 U3850 ( .A1(n4667), .A2(n4603), .ZN(n3334) );
  AND2_X2 U3851 ( .A1(n3189), .A2(n3213), .ZN(n5515) );
  OR2_X1 U3852 ( .A1(n6727), .A2(n4263), .ZN(n4264) );
  OR2_X1 U3853 ( .A1(n3293), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n2992)
         );
  AND2_X2 U3854 ( .A1(n6016), .A2(n3909), .ZN(n6298) );
  AOI21_X1 U3855 ( .B1(n3082), .B2(n3465), .A(n3130), .ZN(n3083) );
  OR2_X1 U3856 ( .A1(n3087), .A2(n3086), .ZN(n3090) );
  OR2_X1 U3857 ( .A1(n3361), .A2(n3360), .ZN(n3446) );
  OAI22_X1 U3858 ( .A1(n3109), .A2(n3108), .B1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n6582), .ZN(n3116) );
  NAND2_X1 U3859 ( .A1(n3262), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3052)
         );
  AOI22_X1 U3860 ( .A1(n3247), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3341), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3138) );
  NAND2_X1 U3861 ( .A1(n3098), .A2(n3097), .ZN(n3109) );
  AND2_X1 U3862 ( .A1(n5385), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3096)
         );
  OAI21_X1 U3863 ( .B1(n3503), .B2(n4932), .A(n3362), .ZN(n3434) );
  OR2_X1 U3864 ( .A1(n5848), .A2(n6002), .ZN(n3514) );
  OR2_X1 U3865 ( .A1(n3373), .A2(n3372), .ZN(n3449) );
  NAND2_X1 U3866 ( .A1(n4595), .A2(n6615), .ZN(n3300) );
  INV_X1 U3867 ( .A(n3374), .ZN(n3503) );
  OAI21_X1 U3868 ( .B1(n3503), .B2(n4861), .A(n3466), .ZN(n3467) );
  NOR2_X1 U3869 ( .A1(n4157), .A2(n4503), .ZN(n4179) );
  INV_X1 U3870 ( .A(n5439), .ZN(n3713) );
  CLKBUF_X2 U3871 ( .A(n3261), .Z(n4213) );
  AND2_X1 U3872 ( .A1(n3585), .A2(n3679), .ZN(n3586) );
  INV_X1 U3873 ( .A(n5458), .ZN(n3510) );
  OR2_X1 U3874 ( .A1(n3274), .A2(n3273), .ZN(n3391) );
  OR2_X1 U3875 ( .A1(n3125), .A2(n3124), .ZN(n3127) );
  INV_X1 U3876 ( .A(n3834), .ZN(n3835) );
  OR2_X1 U3877 ( .A1(n3978), .A2(n5662), .ZN(n3987) );
  AND2_X1 U3878 ( .A1(n4178), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4158)
         );
  NOR2_X1 U3879 ( .A1(n3624), .A2(n5196), .ZN(n3641) );
  NAND2_X1 U3880 ( .A1(n3468), .A2(n3388), .ZN(n3508) );
  AOI21_X1 U3881 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6615), .A(n3123), 
        .ZN(n3129) );
  OAI21_X1 U3882 ( .B1(n2965), .B2(n3099), .A(n3309), .ZN(n3326) );
  AND2_X1 U3883 ( .A1(n4280), .A2(REIP_REG_31__SCAN_IN), .ZN(n4281) );
  OR2_X1 U3884 ( .A1(n5886), .A2(n5898), .ZN(n4496) );
  INV_X1 U3885 ( .A(n4270), .ZN(n4261) );
  BUF_X1 U3886 ( .A(n3987), .Z(n4076) );
  NAND2_X1 U3887 ( .A1(n4557), .A2(n5662), .ZN(n4082) );
  AND2_X1 U3888 ( .A1(n4479), .A2(n5578), .ZN(n4210) );
  INV_X1 U3889 ( .A(n3885), .ZN(n4242) );
  AND2_X1 U3890 ( .A1(n3818), .A2(n3817), .ZN(n5652) );
  INV_X1 U3891 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5273) );
  NOR2_X1 U3892 ( .A1(n4451), .A2(n5974), .ZN(n4441) );
  AND2_X1 U3893 ( .A1(n5848), .A2(n5987), .ZN(n5502) );
  INV_X1 U3894 ( .A(n6338), .ZN(n4716) );
  AND2_X1 U3895 ( .A1(n3192), .A2(n3183), .ZN(n3509) );
  NAND2_X1 U3896 ( .A1(n3425), .A2(n3415), .ZN(n4700) );
  XNOR2_X1 U3897 ( .A(n3399), .B(n3398), .ZN(n3400) );
  OR2_X1 U3898 ( .A1(n5621), .A2(n6157), .ZN(n4284) );
  NAND2_X1 U3899 ( .A1(n6161), .A2(EBX_REG_25__SCAN_IN), .ZN(n4506) );
  NAND2_X1 U3900 ( .A1(n6045), .A2(n4261), .ZN(n5488) );
  INV_X1 U3901 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6058) );
  NOR2_X1 U3902 ( .A1(n6095), .A2(n3590), .ZN(n3619) );
  INV_X1 U3903 ( .A(n4264), .ZN(n4267) );
  AND2_X1 U3904 ( .A1(n4311), .A2(n4250), .ZN(n4251) );
  NAND2_X1 U3905 ( .A1(n5575), .A2(n6178), .ZN(n4316) );
  INV_X1 U3906 ( .A(n5522), .ZN(n5661) );
  INV_X1 U3907 ( .A(n5440), .ZN(n5481) );
  INV_X1 U3908 ( .A(n4583), .ZN(n3991) );
  OR2_X1 U3909 ( .A1(n4480), .A2(n4187), .ZN(n3906) );
  AND2_X1 U3910 ( .A1(n3914), .A2(n3913), .ZN(n3915) );
  AND2_X1 U3911 ( .A1(n3549), .A2(n3548), .ZN(n4591) );
  INV_X1 U3912 ( .A(n6330), .ZN(n5996) );
  NAND2_X1 U3913 ( .A1(n3422), .A2(n3421), .ZN(n6286) );
  NAND2_X1 U3914 ( .A1(n4097), .A2(n4516), .ZN(n5816) );
  NAND2_X1 U3915 ( .A1(n4733), .A2(n5387), .ZN(n5379) );
  OR2_X1 U3916 ( .A1(n4980), .A2(n4891), .ZN(n4965) );
  INV_X1 U3917 ( .A(n5087), .ZN(n5113) );
  INV_X1 U3918 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6582) );
  INV_X1 U3919 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6631) );
  NOR2_X1 U3920 ( .A1(n6697), .A2(n4493), .ZN(n5585) );
  AND2_X1 U3921 ( .A1(n3884), .A2(n4157), .ZN(n5884) );
  NOR2_X1 U3922 ( .A1(n5488), .A2(n5489), .ZN(n6034) );
  NAND2_X1 U3923 ( .A1(n3675), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3697)
         );
  INV_X1 U3924 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5196) );
  NOR2_X1 U3925 ( .A1(n3579), .A2(n6111), .ZN(n3588) );
  NOR2_X1 U3926 ( .A1(n4262), .A2(n4265), .ZN(n6170) );
  NAND2_X1 U3927 ( .A1(n4025), .A2(n5662), .ZN(n4542) );
  NAND2_X1 U3928 ( .A1(n4435), .A2(n3906), .ZN(n5548) );
  CLKBUF_X1 U3929 ( .A(n4576), .Z(n4650) );
  INV_X1 U3930 ( .A(n6597), .ZN(n6730) );
  OAI21_X1 U3931 ( .B1(n6731), .B2(n6729), .A(n4532), .ZN(n6280) );
  NAND2_X1 U3932 ( .A1(n3801), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3834)
         );
  INV_X1 U3933 ( .A(n5758), .ZN(n6192) );
  NOR2_X1 U3934 ( .A1(n4606), .A2(n6598), .ZN(n4625) );
  OR2_X1 U3935 ( .A1(n4592), .A2(n4591), .ZN(n4594) );
  AOI22_X1 U3936 ( .A1(n5702), .A2(n5710), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5974), .ZN(n5703) );
  AND2_X1 U3937 ( .A1(n5799), .A2(n5809), .ZN(n5791) );
  INV_X1 U3938 ( .A(n6309), .ZN(n6284) );
  OR2_X1 U3939 ( .A1(n5462), .A2(n4093), .ZN(n5977) );
  CLKBUF_X1 U3940 ( .A(n5454), .Z(n5457) );
  CLKBUF_X1 U3941 ( .A(n5026), .Z(n5029) );
  CLKBUF_X1 U3942 ( .A(n4862), .Z(n4863) );
  INV_X1 U3943 ( .A(n5816), .ZN(n6332) );
  AND2_X1 U3944 ( .A1(n4097), .A2(n4091), .ZN(n6330) );
  INV_X1 U3945 ( .A(n4768), .ZN(n5123) );
  NOR2_X1 U3946 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6611) );
  INV_X1 U3947 ( .A(n4965), .ZN(n6377) );
  AND2_X1 U3948 ( .A1(n5862), .A2(n5860), .ZN(n5217) );
  AND2_X1 U3949 ( .A1(n6424), .A2(n5388), .ZN(n6418) );
  OR3_X1 U3950 ( .A1(n6397), .A2(n6396), .A3(n6395), .ZN(n6419) );
  INV_X1 U3951 ( .A(n6499), .ZN(n6464) );
  NOR2_X1 U3952 ( .A1(n6345), .A2(n3350), .ZN(n6424) );
  AND2_X1 U3953 ( .A1(n4702), .A2(n5387), .ZN(n6385) );
  INV_X1 U3954 ( .A(n5069), .ZN(n6423) );
  NOR2_X1 U3955 ( .A1(n6251), .A2(n5123), .ZN(n6518) );
  NOR2_X1 U3956 ( .A1(n6259), .A2(n5123), .ZN(n6542) );
  NOR2_X1 U3957 ( .A1(n6264), .A2(n5123), .ZN(n6565) );
  NOR2_X1 U3958 ( .A1(n4951), .A2(n4802), .ZN(n6523) );
  NOR2_X1 U3959 ( .A1(n4951), .A2(n3281), .ZN(n6547) );
  NOR2_X1 U3960 ( .A1(n4951), .A2(n5669), .ZN(n6563) );
  INV_X1 U3961 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6015) );
  OR2_X1 U3962 ( .A1(n5556), .A2(n4486), .ZN(n6039) );
  INV_X1 U3963 ( .A(n6161), .ZN(n6129) );
  AOI21_X1 U3964 ( .B1(n5687), .B2(n6179), .A(n4317), .ZN(n4434) );
  INV_X1 U3965 ( .A(n6178), .ZN(n5666) );
  OR2_X1 U3966 ( .A1(n5531), .A2(n4754), .ZN(n5668) );
  OR2_X1 U3967 ( .A1(n6210), .A2(n6730), .ZN(n6199) );
  INV_X1 U3968 ( .A(n6210), .ZN(n6228) );
  NAND2_X2 U3969 ( .A1(n4625), .A2(n4535), .ZN(n6273) );
  AOI21_X1 U3970 ( .B1(n5971), .B2(n6296), .A(n4444), .ZN(n4445) );
  NAND2_X2 U3971 ( .A1(n4625), .A2(n3952), .ZN(n6016) );
  AND2_X1 U3972 ( .A1(n5791), .A2(n4110), .ZN(n5975) );
  INV_X1 U3973 ( .A(n6328), .ZN(n6309) );
  NAND2_X1 U3974 ( .A1(n4097), .A2(n3959), .ZN(n5997) );
  AND2_X1 U3975 ( .A1(n4737), .A2(n4736), .ZN(n4958) );
  INV_X1 U3976 ( .A(n4950), .ZN(n4937) );
  AOI21_X1 U3977 ( .B1(n6352), .B2(n6353), .A(n6351), .ZN(n6384) );
  NAND2_X1 U3978 ( .A1(n6424), .A2(n6385), .ZN(n6459) );
  NAND2_X1 U3979 ( .A1(n6424), .A2(n6423), .ZN(n6499) );
  INV_X1 U3980 ( .A(n6518), .ZN(n5375) );
  INV_X1 U3981 ( .A(n6524), .ZN(n5371) );
  INV_X1 U3982 ( .A(n6565), .ZN(n5356) );
  NAND2_X1 U3983 ( .A1(n5070), .A2(n6385), .ZN(n6558) );
  AND2_X1 U3984 ( .A1(n5068), .A2(n5067), .ZN(n5115) );
  INV_X1 U3985 ( .A(n6504), .ZN(n5411) );
  INV_X1 U3986 ( .A(n6555), .ZN(n5398) );
  INV_X1 U3987 ( .A(n6621), .ZN(n6715) );
  INV_X1 U3988 ( .A(n6712), .ZN(n6630) );
  INV_X1 U3989 ( .A(n6700), .ZN(n6702) );
  OAI21_X1 U3990 ( .B1(n5931), .B2(n6039), .A(n2985), .ZN(U2799) );
  NAND2_X1 U3991 ( .A1(n4446), .A2(n4445), .ZN(U2960) );
  NOR2_X2 U3992 ( .A1(n2993), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4610)
         );
  AND2_X2 U3993 ( .A1(n4610), .A2(n4660), .ZN(n3262) );
  NAND2_X1 U3994 ( .A1(n3262), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n2999)
         );
  INV_X1 U3995 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n2994) );
  AND2_X2 U3996 ( .A1(n2994), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3005)
         );
  AND2_X4 U3997 ( .A1(n4608), .A2(n3005), .ZN(n4218) );
  NAND2_X1 U3998 ( .A1(n4218), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n2998) );
  AND2_X2 U3999 ( .A1(n4608), .A2(n4667), .ZN(n3166) );
  NAND2_X1 U4000 ( .A1(n3166), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n2997) );
  AND2_X4 U4001 ( .A1(n4670), .A2(n2995), .ZN(n4127) );
  NAND2_X1 U4002 ( .A1(n4127), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n2996) );
  AND2_X2 U4003 ( .A1(n3000), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4662)
         );
  AND2_X2 U4004 ( .A1(n4608), .A2(n4662), .ZN(n3263) );
  NAND2_X1 U4005 ( .A1(n3263), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3004) );
  NOR2_X4 U4006 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3010) );
  AND2_X4 U4007 ( .A1(n3005), .A2(n3010), .ZN(n4133) );
  NAND2_X1 U4008 ( .A1(n4133), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3003) );
  AND2_X2 U4009 ( .A1(n4662), .A2(n4603), .ZN(n3161) );
  NAND2_X1 U4010 ( .A1(n3161), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3002)
         );
  NAND2_X1 U4011 ( .A1(n3339), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3001)
         );
  AND2_X2 U4012 ( .A1(n4608), .A2(n4660), .ZN(n3646) );
  NAND2_X1 U4013 ( .A1(n3646), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3009)
         );
  NAND2_X1 U4014 ( .A1(n3228), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3008) );
  NAND2_X1 U4015 ( .A1(n3247), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3007) );
  NAND2_X1 U4016 ( .A1(n3341), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3006)
         );
  AND2_X2 U4017 ( .A1(n4610), .A2(n4662), .ZN(n3261) );
  NAND2_X1 U4018 ( .A1(n3261), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3014)
         );
  NAND2_X1 U4019 ( .A1(n4223), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3013) );
  AND2_X2 U4020 ( .A1(n3010), .A2(n4667), .ZN(n3133) );
  NAND2_X1 U4021 ( .A1(n3133), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3012) );
  NAND2_X1 U4022 ( .A1(n3334), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3011) );
  NAND2_X1 U4023 ( .A1(n3166), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3022) );
  NAND2_X1 U4024 ( .A1(n4218), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3021) );
  NAND2_X1 U4025 ( .A1(n3262), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3020)
         );
  NAND2_X1 U4026 ( .A1(n3161), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3019)
         );
  NAND2_X1 U4027 ( .A1(n4223), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3026) );
  NAND2_X1 U4028 ( .A1(n3263), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3025) );
  NAND2_X1 U4029 ( .A1(n3646), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3024)
         );
  NAND2_X1 U4030 ( .A1(n3339), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3023)
         );
  NAND2_X1 U4031 ( .A1(n3228), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3030) );
  NAND2_X1 U4032 ( .A1(n4133), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3029) );
  NAND2_X1 U4033 ( .A1(n3247), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3028) );
  NAND2_X1 U4034 ( .A1(n3341), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3027)
         );
  NAND2_X1 U4035 ( .A1(n3261), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3034)
         );
  NAND2_X1 U4036 ( .A1(n3133), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3033) );
  NAND2_X1 U4037 ( .A1(n3334), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3032) );
  NAND2_X1 U4038 ( .A1(n4127), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3031) );
  NAND2_X1 U4039 ( .A1(n3263), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3042) );
  NAND2_X1 U4040 ( .A1(n3228), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3041) );
  NAND2_X1 U4041 ( .A1(n3247), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3040) );
  NAND2_X1 U4042 ( .A1(n3341), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3039)
         );
  NAND2_X1 U4043 ( .A1(n4218), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3046) );
  NAND2_X1 U4044 ( .A1(n3261), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3045)
         );
  NAND2_X1 U4045 ( .A1(n3161), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3044)
         );
  NAND2_X1 U4046 ( .A1(n3133), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3043) );
  NAND2_X1 U4047 ( .A1(n4223), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3050) );
  NAND2_X1 U4048 ( .A1(n4133), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3049) );
  NAND2_X1 U4049 ( .A1(n3646), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3048)
         );
  NAND2_X1 U4050 ( .A1(n3339), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3047)
         );
  NAND2_X1 U4051 ( .A1(n3166), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3051) );
  NAND2_X1 U4052 ( .A1(n3052), .A2(n3051), .ZN(n3056) );
  NAND2_X1 U4053 ( .A1(n4127), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3054) );
  NAND2_X1 U4054 ( .A1(n3334), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3053) );
  NAND2_X1 U4055 ( .A1(n3054), .A2(n3053), .ZN(n3055) );
  NOR2_X2 U4056 ( .A1(n3056), .A2(n3055), .ZN(n3177) );
  NAND4_X4 U4057 ( .A1(n3177), .A2(n3176), .A3(n3174), .A4(n3175), .ZN(n3183)
         );
  AND2_X1 U4058 ( .A1(n4802), .A2(n3183), .ZN(n3057) );
  NAND2_X1 U4059 ( .A1(n3261), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3061)
         );
  NAND2_X1 U4060 ( .A1(n3133), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3060) );
  NAND2_X1 U4061 ( .A1(n3334), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3059) );
  NAND2_X1 U4062 ( .A1(n4127), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3058) );
  NAND2_X1 U4063 ( .A1(n3166), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3065) );
  NAND2_X1 U4064 ( .A1(n4218), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3064) );
  NAND2_X1 U4065 ( .A1(n3262), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3063)
         );
  NAND2_X1 U4066 ( .A1(n3161), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3062)
         );
  NAND2_X1 U4067 ( .A1(n3228), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3069) );
  NAND2_X1 U4068 ( .A1(n4133), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3068) );
  NAND2_X1 U4069 ( .A1(n3247), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3067) );
  NAND2_X1 U4070 ( .A1(n3341), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3066)
         );
  NAND2_X1 U4071 ( .A1(n4223), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3073) );
  NAND2_X1 U4072 ( .A1(n3263), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3072) );
  NAND2_X1 U4073 ( .A1(n3646), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3071)
         );
  NAND2_X1 U4074 ( .A1(n3339), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3070)
         );
  INV_X1 U4075 ( .A(n3205), .ZN(n3190) );
  AND2_X1 U4076 ( .A1(n3078), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3079)
         );
  NOR2_X1 U4077 ( .A1(n3096), .A2(n3079), .ZN(n3082) );
  INV_X1 U4078 ( .A(n3082), .ZN(n3080) );
  OAI21_X1 U4079 ( .B1(n3190), .B2(n3080), .A(n3081), .ZN(n3084) );
  AOI21_X1 U4080 ( .B1(n3102), .B2(n3084), .A(n3083), .ZN(n3087) );
  XNOR2_X1 U4081 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3095) );
  INV_X1 U4082 ( .A(n3095), .ZN(n3085) );
  XNOR2_X1 U4083 ( .A(n3085), .B(n3096), .ZN(n3942) );
  INV_X1 U4084 ( .A(n3942), .ZN(n3088) );
  AND2_X1 U4085 ( .A1(n3130), .A2(n3088), .ZN(n3086) );
  INV_X1 U4086 ( .A(n3090), .ZN(n3094) );
  OAI21_X1 U4087 ( .B1(n3088), .B2(n6615), .A(n3120), .ZN(n3089) );
  INV_X1 U4088 ( .A(n3089), .ZN(n3093) );
  INV_X1 U4089 ( .A(n3183), .ZN(n3281) );
  AOI21_X1 U4090 ( .B1(n3465), .B2(n3192), .A(n3281), .ZN(n3092) );
  NOR2_X1 U4091 ( .A1(n3090), .A2(n3089), .ZN(n3091) );
  OAI22_X1 U4092 ( .A1(n3094), .A2(n3093), .B1(n3092), .B2(n3091), .ZN(n3106)
         );
  NAND2_X1 U4093 ( .A1(n3096), .A2(n3095), .ZN(n3098) );
  NAND2_X1 U4094 ( .A1(n6575), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3097) );
  XNOR2_X1 U4095 ( .A(n3099), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3100)
         );
  XNOR2_X1 U4096 ( .A(n3109), .B(n3100), .ZN(n3939) );
  NAND2_X1 U4097 ( .A1(n3465), .A2(n3939), .ZN(n3101) );
  OAI211_X1 U4098 ( .C1(n3503), .C2(n3939), .A(n3102), .B(n3101), .ZN(n3105)
         );
  INV_X1 U4099 ( .A(n3101), .ZN(n3104) );
  INV_X1 U4100 ( .A(n3102), .ZN(n3103) );
  AOI22_X1 U4101 ( .A1(n3106), .A2(n3105), .B1(n3104), .B2(n3103), .ZN(n3107)
         );
  INV_X1 U4102 ( .A(n3107), .ZN(n3114) );
  NOR2_X1 U4103 ( .A1(n3099), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3108)
         );
  XNOR2_X1 U4104 ( .A(n3110), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3111)
         );
  XNOR2_X1 U4105 ( .A(n3116), .B(n3111), .ZN(n3938) );
  AND2_X1 U4106 ( .A1(n3130), .A2(n3938), .ZN(n3112) );
  NOR2_X1 U4107 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n6501), .ZN(n3115)
         );
  NAND2_X1 U4108 ( .A1(n6501), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3117) );
  INV_X1 U4109 ( .A(n3125), .ZN(n3119) );
  NAND3_X1 U4110 ( .A1(n3119), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(n3570), .ZN(n3941) );
  NOR2_X1 U4111 ( .A1(n3374), .A2(n3941), .ZN(n3121) );
  OAI22_X1 U4112 ( .A1(n3122), .A2(n3121), .B1(n3120), .B2(n3941), .ZN(n3123)
         );
  NAND2_X1 U4113 ( .A1(n3570), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3126) );
  NAND2_X1 U4114 ( .A1(n3465), .A2(n3937), .ZN(n3128) );
  NAND2_X1 U4115 ( .A1(n3129), .A2(n3128), .ZN(n3132) );
  NAND2_X1 U4116 ( .A1(n3130), .A2(n3937), .ZN(n3131) );
  NAND2_X1 U4117 ( .A1(n6614), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3330) );
  AOI22_X1 U4118 ( .A1(n4218), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3166), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3137) );
  AOI22_X1 U4119 ( .A1(n3133), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3135) );
  AOI22_X1 U4120 ( .A1(n3261), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3334), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3134) );
  AOI22_X1 U4121 ( .A1(n3263), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3141) );
  AOI22_X1 U4122 ( .A1(n4133), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3228), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3140) );
  AOI22_X1 U4123 ( .A1(n3646), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3339), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3139) );
  AND4_X2 U4124 ( .A1(n3141), .A2(n3140), .A3(n3139), .A4(n3138), .ZN(n3142)
         );
  NAND2_X2 U4125 ( .A1(n3143), .A2(n3142), .ZN(n3179) );
  AOI22_X1 U4126 ( .A1(n3262), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3161), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3146) );
  AOI22_X1 U4127 ( .A1(n3133), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3145) );
  AOI22_X1 U4128 ( .A1(n3261), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3334), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3144) );
  AOI22_X1 U4129 ( .A1(n3263), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3150) );
  AOI22_X1 U4130 ( .A1(n3646), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3339), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3149) );
  AOI22_X1 U4131 ( .A1(n3247), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3341), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3148) );
  NAND2_X1 U4132 ( .A1(n3179), .A2(n3195), .ZN(n3282) );
  AOI22_X1 U4133 ( .A1(n3262), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3161), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3155) );
  AOI22_X1 U4134 ( .A1(n3261), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3334), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3154) );
  AOI22_X1 U4135 ( .A1(n3133), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3153) );
  AOI22_X1 U4136 ( .A1(n4218), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3166), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3152) );
  AOI22_X1 U4137 ( .A1(n4133), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3228), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3159) );
  AOI22_X1 U4138 ( .A1(n3263), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4223), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3158) );
  AOI22_X1 U4139 ( .A1(n3646), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3339), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3157) );
  AOI22_X1 U4140 ( .A1(n3247), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3341), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3156) );
  AOI22_X1 U4141 ( .A1(n3161), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3646), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3165) );
  AOI22_X1 U4142 ( .A1(n3228), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3164) );
  AOI22_X1 U4143 ( .A1(n3261), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3163) );
  AOI22_X1 U4144 ( .A1(n4218), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3262), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3162) );
  NAND4_X1 U4145 ( .A1(n3165), .A2(n3164), .A3(n3163), .A4(n3162), .ZN(n3172)
         );
  AOI22_X1 U4146 ( .A1(n3263), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3166), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3170) );
  AOI22_X1 U4147 ( .A1(n4133), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3341), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3169) );
  AOI22_X1 U4148 ( .A1(n3334), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3168) );
  AOI22_X1 U4149 ( .A1(n4223), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3339), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3167) );
  NAND4_X1 U4150 ( .A1(n3170), .A2(n3169), .A3(n3168), .A4(n3167), .ZN(n3171)
         );
  OR2_X2 U4151 ( .A1(n3172), .A2(n3171), .ZN(n3213) );
  NAND2_X2 U4152 ( .A1(n2973), .A2(n3213), .ZN(n3974) );
  NOR2_X1 U4153 ( .A1(n3974), .A2(n4813), .ZN(n3173) );
  AND2_X1 U4154 ( .A1(n3285), .A2(n3173), .ZN(n3952) );
  NAND2_X1 U4155 ( .A1(n3542), .A2(n3956), .ZN(n3182) );
  NAND2_X2 U4156 ( .A1(n3179), .A2(n3178), .ZN(n4303) );
  NAND2_X1 U4157 ( .A1(n4303), .A2(n2973), .ZN(n3180) );
  NAND2_X1 U4158 ( .A1(n3180), .A2(n3195), .ZN(n3181) );
  NAND2_X1 U4159 ( .A1(n3182), .A2(n3181), .ZN(n3184) );
  NAND2_X1 U4160 ( .A1(n3198), .A2(n3213), .ZN(n3211) );
  NAND2_X1 U4161 ( .A1(n3184), .A2(n3211), .ZN(n3284) );
  NOR2_X1 U4162 ( .A1(n3185), .A2(n2973), .ZN(n3186) );
  AND2_X1 U4163 ( .A1(n3194), .A2(n3195), .ZN(n3187) );
  AND2_X4 U4164 ( .A1(n3953), .A2(n3188), .ZN(n6731) );
  NAND2_X1 U4165 ( .A1(n3932), .A2(n6731), .ZN(n3191) );
  NAND2_X1 U4166 ( .A1(n3190), .A2(n5515), .ZN(n4596) );
  NAND2_X1 U4167 ( .A1(n5174), .A2(n3183), .ZN(n3193) );
  XNOR2_X1 U4168 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .ZN(
        n3925) );
  NAND2_X1 U4169 ( .A1(n4802), .A2(n3925), .ZN(n3283) );
  AOI21_X1 U4170 ( .B1(n3193), .B2(n3283), .A(n3974), .ZN(n3200) );
  AND2_X1 U4171 ( .A1(n4303), .A2(n3195), .ZN(n3196) );
  NAND2_X1 U4172 ( .A1(n4755), .A2(n3956), .ZN(n3199) );
  NAND4_X1 U4173 ( .A1(n3207), .A2(n3210), .A3(n3200), .A4(n3208), .ZN(n3201)
         );
  INV_X1 U4174 ( .A(n3330), .ZN(n6607) );
  NAND2_X1 U4175 ( .A1(n6611), .A2(n6615), .ZN(n3908) );
  MUX2_X1 U4176 ( .A(n6607), .B(n3908), .S(n5385), .Z(n3202) );
  INV_X1 U4177 ( .A(n5174), .ZN(n4514) );
  AOI22_X1 U4178 ( .A1(n4514), .A2(n3205), .B1(n4628), .B2(n3204), .ZN(n3206)
         );
  AND2_X1 U4179 ( .A1(n3207), .A2(n3206), .ZN(n3968) );
  INV_X1 U4180 ( .A(n3208), .ZN(n3209) );
  NAND2_X1 U4181 ( .A1(n3209), .A2(n3192), .ZN(n3220) );
  INV_X1 U4182 ( .A(n3210), .ZN(n3218) );
  NAND2_X1 U4183 ( .A1(n3211), .A2(n6731), .ZN(n3216) );
  NAND2_X1 U4184 ( .A1(n3969), .A2(n4802), .ZN(n3214) );
  INV_X1 U4185 ( .A(n3213), .ZN(n4822) );
  NAND2_X1 U4186 ( .A1(n3214), .A2(n4822), .ZN(n3215) );
  NAND4_X1 U4187 ( .A1(n3216), .A2(n6611), .A3(n3215), .A4(
        STATE2_REG_0__SCAN_IN), .ZN(n3217) );
  NOR2_X1 U4188 ( .A1(n3218), .A2(n3217), .ZN(n3219) );
  INV_X1 U4189 ( .A(n3222), .ZN(n3225) );
  INV_X1 U4190 ( .A(n3223), .ZN(n3224) );
  NAND2_X1 U4191 ( .A1(n3225), .A2(n3224), .ZN(n3226) );
  INV_X1 U4192 ( .A(n3544), .ZN(n3227) );
  AOI22_X1 U4193 ( .A1(n4141), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3241) );
  AOI22_X1 U4194 ( .A1(n4133), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4664), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3234) );
  AOI22_X1 U4196 ( .A1(n3263), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3233) );
  AOI22_X1 U4198 ( .A1(n4225), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3232) );
  BUF_X1 U4199 ( .A(n3247), .Z(n3264) );
  AOI22_X1 U4200 ( .A1(n3264), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3230), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3231) );
  NAND4_X1 U4201 ( .A1(n3234), .A2(n3233), .A3(n3232), .A4(n3231), .ZN(n3240)
         );
  AOI22_X1 U4202 ( .A1(n4218), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3238) );
  AOI22_X1 U4203 ( .A1(n4213), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3235), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3237) );
  AOI22_X1 U4204 ( .A1(n3823), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3236) );
  NAND3_X1 U4205 ( .A1(n3238), .A2(n3237), .A3(n3236), .ZN(n3239) );
  NOR2_X1 U4206 ( .A1(n4305), .A2(n3479), .ZN(n3260) );
  NAND2_X1 U4207 ( .A1(n2968), .A2(n3479), .ZN(n3257) );
  AOI22_X1 U4208 ( .A1(n4213), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3246) );
  AOI22_X1 U4209 ( .A1(n4664), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3263), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3245) );
  AOI22_X1 U4211 ( .A1(n3661), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3244) );
  BUF_X1 U4212 ( .A(n3823), .Z(n4190) );
  AOI22_X1 U4213 ( .A1(n3823), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3243) );
  NAND4_X1 U4214 ( .A1(n3246), .A2(n3245), .A3(n3244), .A4(n3243), .ZN(n3256)
         );
  AOI22_X1 U4215 ( .A1(n4141), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3254) );
  AOI22_X1 U4218 ( .A1(n4132), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3248), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3253) );
  BUF_X1 U4219 ( .A(n3341), .Z(n3249) );
  AOI22_X1 U4220 ( .A1(n4133), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3252) );
  AOI22_X1 U4221 ( .A1(n4225), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3251) );
  NAND4_X1 U4222 ( .A1(n3254), .A2(n3253), .A3(n3252), .A4(n3251), .ZN(n3255)
         );
  INV_X1 U4223 ( .A(n3392), .ZN(n3402) );
  MUX2_X1 U4224 ( .A(n3260), .B(n3388), .S(n3402), .Z(n3399) );
  INV_X1 U4225 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4889) );
  AOI21_X1 U4226 ( .B1(n4813), .B2(n3392), .A(n6615), .ZN(n3258) );
  OAI211_X1 U4227 ( .C1(n3503), .C2(n4889), .A(n3258), .B(n3257), .ZN(n3397)
         );
  AOI21_X1 U4228 ( .B1(n3399), .B2(n3397), .A(n3388), .ZN(n3259) );
  NAND2_X1 U4229 ( .A1(n3374), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3277) );
  INV_X1 U4230 ( .A(n3260), .ZN(n3276) );
  INV_X1 U4231 ( .A(n3502), .ZN(n3323) );
  AOI22_X1 U4232 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n4213), .B1(n4141), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3268) );
  AOI22_X1 U4233 ( .A1(n4215), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3267) );
  AOI22_X1 U4234 ( .A1(n4224), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3266) );
  AOI22_X1 U4235 ( .A1(n4132), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3265) );
  NAND4_X1 U4236 ( .A1(n3268), .A2(n3267), .A3(n3266), .A4(n3265), .ZN(n3274)
         );
  AOI22_X1 U4237 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n4195), .B1(n4664), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3272) );
  AOI22_X1 U4238 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n3661), .B1(n3242), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3271) );
  AOI22_X1 U4239 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4190), .B1(n3248), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3270) );
  AOI22_X1 U4240 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n4225), .B1(n3249), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3269) );
  NAND4_X1 U4241 ( .A1(n3272), .A2(n3271), .A3(n3270), .A4(n3269), .ZN(n3273)
         );
  NAND2_X1 U4242 ( .A1(n3323), .A2(n3391), .ZN(n3275) );
  NAND2_X1 U4243 ( .A1(n3408), .A2(n3409), .ZN(n3301) );
  NOR2_X1 U4244 ( .A1(n3974), .A2(n3183), .ZN(n3279) );
  INV_X1 U4245 ( .A(n3932), .ZN(n3278) );
  INV_X1 U4246 ( .A(n3282), .ZN(n3537) );
  NOR2_X2 U4247 ( .A1(n4597), .A2(n3282), .ZN(n3955) );
  AOI21_X1 U4248 ( .B1(n4518), .B2(n3283), .A(n3955), .ZN(n3287) );
  INV_X1 U4249 ( .A(n3284), .ZN(n3286) );
  AND2_X2 U4250 ( .A1(n3286), .A2(n2981), .ZN(n3935) );
  NAND2_X1 U4251 ( .A1(n3287), .A2(n3951), .ZN(n3288) );
  NAND2_X1 U4252 ( .A1(n3288), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3295) );
  INV_X1 U4253 ( .A(n3295), .ZN(n3291) );
  XNOR2_X1 U4254 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5064) );
  OR2_X1 U4255 ( .A1(n5064), .A2(n3908), .ZN(n3290) );
  NAND2_X1 U4256 ( .A1(n3330), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3289) );
  NAND2_X1 U4257 ( .A1(n3290), .A2(n3289), .ZN(n3293) );
  NAND2_X1 U4258 ( .A1(n3291), .A2(n2992), .ZN(n3302) );
  INV_X1 U4259 ( .A(n3293), .ZN(n3294) );
  OAI211_X1 U4260 ( .C1(n2965), .C2(n2993), .A(n3295), .B(n3294), .ZN(n3304)
         );
  NAND2_X1 U4261 ( .A1(n3302), .A2(n3304), .ZN(n3298) );
  INV_X1 U4262 ( .A(n4305), .ZN(n3320) );
  NAND2_X1 U4263 ( .A1(n3320), .A2(n3391), .ZN(n3299) );
  NAND2_X1 U4264 ( .A1(n3303), .A2(n3302), .ZN(n3305) );
  INV_X1 U4265 ( .A(n3908), .ZN(n3331) );
  AND2_X1 U4266 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3306) );
  NAND2_X1 U4267 ( .A1(n3306), .A2(n6582), .ZN(n6502) );
  INV_X1 U4268 ( .A(n3306), .ZN(n3307) );
  NAND2_X1 U4269 ( .A1(n3307), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3308) );
  NAND2_X1 U4270 ( .A1(n6502), .A2(n3308), .ZN(n4735) );
  AOI22_X1 U4271 ( .A1(n3331), .A2(n4735), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3330), .ZN(n3309) );
  XNOR2_X1 U4272 ( .A(n2970), .B(n3326), .ZN(n4675) );
  NAND2_X1 U4273 ( .A1(n4675), .A2(n6615), .ZN(n3322) );
  AOI22_X1 U4274 ( .A1(n4218), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4275 ( .A1(n4141), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3312) );
  AOI22_X1 U4276 ( .A1(n4190), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3311) );
  AOI22_X1 U4277 ( .A1(n4213), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3248), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3310) );
  NAND4_X1 U4278 ( .A1(n3313), .A2(n3312), .A3(n3311), .A4(n3310), .ZN(n3319)
         );
  AOI22_X1 U4279 ( .A1(n4133), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4664), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3317) );
  AOI22_X1 U4280 ( .A1(n4215), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4281 ( .A1(n4225), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3315) );
  AOI22_X1 U4282 ( .A1(n4132), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3314) );
  NAND4_X1 U4283 ( .A1(n3317), .A2(n3316), .A3(n3315), .A4(n3314), .ZN(n3318)
         );
  NAND2_X1 U4284 ( .A1(n3320), .A2(n3416), .ZN(n3321) );
  AOI22_X1 U4285 ( .A1(n3374), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3323), 
        .B2(n3416), .ZN(n3324) );
  NAND2_X1 U4286 ( .A1(n3407), .A2(n3406), .ZN(n3405) );
  INV_X1 U4287 ( .A(n3405), .ZN(n3351) );
  INV_X1 U4288 ( .A(n2970), .ZN(n3327) );
  NAND2_X1 U4289 ( .A1(n3327), .A2(n3326), .ZN(n4571) );
  NAND2_X1 U4290 ( .A1(n3328), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3333) );
  NAND3_X1 U4291 ( .A1(n6501), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6430) );
  INV_X1 U4292 ( .A(n6430), .ZN(n6429) );
  NAND2_X1 U4293 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6429), .ZN(n6422) );
  NAND2_X1 U4294 ( .A1(n6501), .A2(n6422), .ZN(n3329) );
  NOR3_X1 U4295 ( .A1(n6501), .A2(n6582), .A3(n6575), .ZN(n5126) );
  NAND2_X1 U4296 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5126), .ZN(n5151) );
  AOI22_X1 U4297 ( .A1(n3331), .A2(n5065), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3330), .ZN(n3332) );
  NAND2_X1 U4298 ( .A1(n4661), .A2(n6615), .ZN(n3349) );
  AOI22_X1 U4299 ( .A1(n3661), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3338) );
  AOI22_X1 U4300 ( .A1(n4141), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3337) );
  INV_X1 U4301 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4374) );
  AOI22_X1 U4302 ( .A1(n4190), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3336) );
  AOI22_X1 U4303 ( .A1(n4213), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3248), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3335) );
  NAND4_X1 U4304 ( .A1(n3338), .A2(n3337), .A3(n3336), .A4(n3335), .ZN(n3347)
         );
  AOI22_X1 U4305 ( .A1(n4195), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4664), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3345) );
  AOI22_X1 U4306 ( .A1(n4215), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3344) );
  AOI22_X1 U4307 ( .A1(n4225), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3343) );
  AOI22_X1 U4308 ( .A1(n4132), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3342) );
  NAND4_X1 U4309 ( .A1(n3345), .A2(n3344), .A3(n3343), .A4(n3342), .ZN(n3346)
         );
  AOI22_X1 U4310 ( .A1(n3374), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3465), 
        .B2(n3428), .ZN(n3348) );
  NAND2_X1 U4311 ( .A1(n3351), .A2(n3350), .ZN(n3436) );
  INV_X1 U4312 ( .A(n3436), .ZN(n3363) );
  INV_X1 U4313 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4932) );
  AOI22_X1 U4314 ( .A1(n4141), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3355) );
  AOI22_X1 U4315 ( .A1(n4215), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3354) );
  AOI22_X1 U4316 ( .A1(n3661), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4317 ( .A1(n4195), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3352) );
  NAND4_X1 U4318 ( .A1(n3355), .A2(n3354), .A3(n3353), .A4(n3352), .ZN(n3361)
         );
  AOI22_X1 U4319 ( .A1(n4224), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4320 ( .A1(n4664), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4132), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4321 ( .A1(n4190), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3357) );
  AOI22_X1 U4322 ( .A1(n4213), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3248), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3356) );
  NAND4_X1 U4323 ( .A1(n3359), .A2(n3358), .A3(n3357), .A4(n3356), .ZN(n3360)
         );
  NAND2_X1 U4324 ( .A1(n3465), .A2(n3446), .ZN(n3362) );
  NAND2_X1 U4325 ( .A1(n3363), .A2(n3434), .ZN(n3444) );
  AOI22_X1 U4326 ( .A1(n3661), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4327 ( .A1(n4141), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4328 ( .A1(n4190), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3365) );
  AOI22_X1 U4329 ( .A1(n4213), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3248), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3364) );
  NAND4_X1 U4330 ( .A1(n3367), .A2(n3366), .A3(n3365), .A4(n3364), .ZN(n3373)
         );
  AOI22_X1 U4331 ( .A1(n4195), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4664), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3371) );
  AOI22_X1 U4332 ( .A1(n4215), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3370) );
  AOI22_X1 U4333 ( .A1(n4225), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4334 ( .A1(n4132), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3368) );
  NAND4_X1 U4335 ( .A1(n3371), .A2(n3370), .A3(n3369), .A4(n3368), .ZN(n3372)
         );
  AOI22_X1 U4336 ( .A1(n3374), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3465), 
        .B2(n3449), .ZN(n3443) );
  OR2_X2 U4337 ( .A1(n3444), .A2(n3443), .ZN(n3457) );
  INV_X1 U4338 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3386) );
  AOI22_X1 U4339 ( .A1(n3661), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4664), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4340 ( .A1(n4213), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3377) );
  AOI22_X1 U4341 ( .A1(n4190), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3376) );
  AOI22_X1 U4342 ( .A1(n4224), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3375) );
  NAND4_X1 U4343 ( .A1(n3378), .A2(n3377), .A3(n3376), .A4(n3375), .ZN(n3384)
         );
  AOI22_X1 U4344 ( .A1(n4215), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4345 ( .A1(n4225), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4132), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3381) );
  AOI22_X1 U4346 ( .A1(n4195), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3248), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3380) );
  AOI22_X1 U4347 ( .A1(n3242), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3379) );
  NAND4_X1 U4348 ( .A1(n3382), .A2(n3381), .A3(n3380), .A4(n3379), .ZN(n3383)
         );
  NAND2_X1 U4349 ( .A1(n3465), .A2(n3470), .ZN(n3385) );
  INV_X1 U4350 ( .A(n3509), .ZN(n3458) );
  XNOR2_X1 U4351 ( .A(n5848), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3527)
         );
  NAND2_X1 U4352 ( .A1(n4701), .A2(n3509), .ZN(n3396) );
  NAND2_X1 U4353 ( .A1(n3392), .A2(n3391), .ZN(n3417) );
  OAI211_X1 U4354 ( .C1(n3392), .C2(n3391), .A(n6731), .B(n3417), .ZN(n3394)
         );
  NOR2_X1 U4355 ( .A1(n3974), .A2(n3281), .ZN(n3393) );
  AND2_X1 U4356 ( .A1(n3394), .A2(n3393), .ZN(n3395) );
  NAND2_X1 U4357 ( .A1(n3396), .A2(n3395), .ZN(n4615) );
  INV_X1 U4358 ( .A(n3397), .ZN(n3398) );
  AND2_X1 U4359 ( .A1(n4813), .A2(n3213), .ZN(n3419) );
  AOI21_X1 U4360 ( .B1(n3402), .B2(n6731), .A(n3419), .ZN(n3403) );
  OAI21_X1 U4361 ( .B1(n5387), .B2(n3458), .A(n3403), .ZN(n4538) );
  NAND2_X1 U4362 ( .A1(n4538), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4537)
         );
  XNOR2_X1 U4363 ( .A(n4537), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4614)
         );
  NAND2_X1 U4364 ( .A1(n4615), .A2(n4614), .ZN(n4617) );
  INV_X1 U4365 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6339) );
  OR2_X1 U4366 ( .A1(n4537), .A2(n6339), .ZN(n3404) );
  NAND2_X1 U4367 ( .A1(n4617), .A2(n3404), .ZN(n6285) );
  INV_X1 U4368 ( .A(n3406), .ZN(n3414) );
  INV_X1 U4369 ( .A(n3407), .ZN(n3413) );
  INV_X1 U4370 ( .A(n3408), .ZN(n3411) );
  INV_X1 U4371 ( .A(n3409), .ZN(n3410) );
  NAND2_X1 U4372 ( .A1(n3411), .A2(n3410), .ZN(n3412) );
  NAND3_X1 U4373 ( .A1(n3414), .A2(n3413), .A3(n3412), .ZN(n3415) );
  OR2_X1 U4374 ( .A1(n4700), .A2(n3458), .ZN(n3422) );
  INV_X1 U4375 ( .A(n3416), .ZN(n3418) );
  NAND2_X1 U4376 ( .A1(n3417), .A2(n3418), .ZN(n3427) );
  OAI21_X1 U4377 ( .B1(n3418), .B2(n3417), .A(n3427), .ZN(n3420) );
  AOI21_X1 U4378 ( .B1(n3420), .B2(n6731), .A(n3419), .ZN(n3421) );
  OAI21_X1 U4379 ( .B1(n6285), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .A(n6286), 
        .ZN(n3424) );
  NAND2_X1 U4380 ( .A1(n6285), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3423)
         );
  NAND2_X1 U4381 ( .A1(n3424), .A2(n3423), .ZN(n4784) );
  NAND2_X1 U4382 ( .A1(n3425), .A2(n4704), .ZN(n3426) );
  NAND2_X1 U4383 ( .A1(n3426), .A2(n3436), .ZN(n3560) );
  NAND2_X1 U4384 ( .A1(n3427), .A2(n3428), .ZN(n3448) );
  OAI211_X1 U4385 ( .C1(n3428), .C2(n3427), .A(n3448), .B(n6731), .ZN(n3429)
         );
  OAI21_X2 U4386 ( .B1(n3560), .B2(n3458), .A(n3429), .ZN(n3431) );
  INV_X1 U4387 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3430) );
  XNOR2_X1 U4388 ( .A(n3431), .B(n3430), .ZN(n4782) );
  NAND2_X1 U4389 ( .A1(n4784), .A2(n4782), .ZN(n3433) );
  NAND2_X1 U4390 ( .A1(n3431), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3432)
         );
  INV_X1 U4391 ( .A(n3434), .ZN(n3435) );
  NAND2_X1 U4392 ( .A1(n3436), .A2(n3435), .ZN(n3437) );
  NAND2_X1 U4393 ( .A1(n3444), .A2(n3437), .ZN(n3566) );
  XNOR2_X1 U4394 ( .A(n3448), .B(n3446), .ZN(n3438) );
  NAND2_X1 U4395 ( .A1(n3438), .A2(n6731), .ZN(n3439) );
  INV_X1 U4396 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3995) );
  XNOR2_X1 U4397 ( .A(n3440), .B(n3995), .ZN(n4718) );
  NAND2_X1 U4398 ( .A1(n4719), .A2(n4718), .ZN(n3442) );
  NAND2_X1 U4399 ( .A1(n3440), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3441)
         );
  NAND2_X1 U4400 ( .A1(n3444), .A2(n3443), .ZN(n3445) );
  INV_X1 U4401 ( .A(n3446), .ZN(n3447) );
  NOR2_X1 U4402 ( .A1(n3448), .A2(n3447), .ZN(n3450) );
  NAND2_X1 U4403 ( .A1(n3450), .A2(n3449), .ZN(n3469) );
  OAI211_X1 U4404 ( .C1(n3450), .C2(n3449), .A(n3469), .B(n6731), .ZN(n3451)
         );
  NAND2_X1 U4405 ( .A1(n4839), .A2(n4838), .ZN(n3454) );
  NAND2_X1 U4406 ( .A1(n3452), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3453)
         );
  NAND2_X1 U4407 ( .A1(n3454), .A2(n3453), .ZN(n4938) );
  INV_X1 U4408 ( .A(n3455), .ZN(n3456) );
  NAND2_X1 U4409 ( .A1(n3457), .A2(n3456), .ZN(n3585) );
  NAND3_X1 U4410 ( .A1(n3468), .A2(n3585), .A3(n3509), .ZN(n3461) );
  XNOR2_X1 U4411 ( .A(n3469), .B(n3470), .ZN(n3459) );
  NAND2_X1 U4412 ( .A1(n3459), .A2(n6731), .ZN(n3460) );
  NAND2_X1 U4413 ( .A1(n3461), .A2(n3460), .ZN(n3462) );
  INV_X1 U4414 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4005) );
  XNOR2_X1 U4415 ( .A(n3462), .B(n4005), .ZN(n4940) );
  NAND2_X1 U4416 ( .A1(n4938), .A2(n4940), .ZN(n3464) );
  NAND2_X1 U4417 ( .A1(n3462), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3463)
         );
  NAND2_X1 U4418 ( .A1(n3464), .A2(n3463), .ZN(n5163) );
  INV_X1 U4419 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4861) );
  NAND2_X1 U4420 ( .A1(n3465), .A2(n3479), .ZN(n3466) );
  NAND2_X1 U4421 ( .A1(n3528), .A2(n3509), .ZN(n3474) );
  INV_X1 U4422 ( .A(n3469), .ZN(n3471) );
  NAND2_X1 U4423 ( .A1(n3471), .A2(n3470), .ZN(n3481) );
  XNOR2_X1 U4424 ( .A(n3481), .B(n3479), .ZN(n3472) );
  NAND2_X1 U4425 ( .A1(n3472), .A2(n6731), .ZN(n3473) );
  NAND2_X1 U4426 ( .A1(n3474), .A2(n3473), .ZN(n3476) );
  INV_X1 U4427 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3475) );
  XNOR2_X1 U4428 ( .A(n3476), .B(n3475), .ZN(n5162) );
  NAND2_X1 U4429 ( .A1(n5163), .A2(n5162), .ZN(n3478) );
  NAND2_X1 U4430 ( .A1(n3476), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3477)
         );
  NAND2_X1 U4431 ( .A1(n3478), .A2(n3477), .ZN(n4862) );
  NAND2_X1 U4432 ( .A1(n6731), .A2(n3479), .ZN(n3480) );
  OR2_X1 U4433 ( .A1(n3481), .A2(n3480), .ZN(n3482) );
  INV_X1 U4434 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4012) );
  XNOR2_X1 U4435 ( .A(n3483), .B(n4012), .ZN(n4864) );
  NAND2_X1 U4436 ( .A1(n4862), .A2(n4864), .ZN(n3485) );
  NAND2_X1 U4437 ( .A1(n3483), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3484)
         );
  INV_X1 U4438 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5194) );
  NOR2_X1 U4439 ( .A1(n3519), .A2(n5194), .ZN(n3487) );
  NAND2_X1 U4440 ( .A1(n5848), .A2(n5194), .ZN(n3486) );
  INV_X1 U4441 ( .A(n5026), .ZN(n3488) );
  INV_X1 U4442 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5032) );
  NAND2_X1 U4443 ( .A1(n3488), .A2(n2988), .ZN(n3489) );
  OR2_X1 U4444 ( .A1(n5848), .A2(n5032), .ZN(n5027) );
  NAND2_X1 U4445 ( .A1(n3489), .A2(n5027), .ZN(n5263) );
  INV_X1 U4446 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U4447 ( .A1(n5263), .A2(n5265), .ZN(n3490) );
  OR2_X1 U4448 ( .A1(n5848), .A2(n5322), .ZN(n5266) );
  NAND2_X1 U4449 ( .A1(n3490), .A2(n5266), .ZN(n5318) );
  INV_X1 U4450 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5320) );
  NAND2_X1 U4451 ( .A1(n5318), .A2(n3491), .ZN(n3493) );
  OR2_X1 U4452 ( .A1(n5848), .A2(n5320), .ZN(n3492) );
  NAND2_X1 U4453 ( .A1(n3493), .A2(n3492), .ZN(n5454) );
  INV_X1 U4454 ( .A(n5454), .ZN(n3511) );
  AOI22_X1 U4455 ( .A1(n3661), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3497) );
  AOI22_X1 U4456 ( .A1(n4195), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3496) );
  AOI22_X1 U4457 ( .A1(n4225), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3248), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3495) );
  AOI22_X1 U4458 ( .A1(n4132), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3494) );
  NAND4_X1 U4459 ( .A1(n3497), .A2(n3496), .A3(n3495), .A4(n3494), .ZN(n3506)
         );
  AOI22_X1 U4460 ( .A1(n4664), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3501) );
  AOI22_X1 U4461 ( .A1(n4215), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4190), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3500) );
  AOI22_X1 U4462 ( .A1(n4141), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3499) );
  AOI22_X1 U4463 ( .A1(n4214), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3498) );
  NAND4_X1 U4464 ( .A1(n3501), .A2(n3500), .A3(n3499), .A4(n3498), .ZN(n3505)
         );
  NAND2_X1 U4465 ( .A1(n3503), .A2(n3502), .ZN(n3504) );
  OAI21_X1 U4466 ( .B1(n3506), .B2(n3505), .A(n3504), .ZN(n3507) );
  NAND2_X1 U4467 ( .A1(n3508), .A2(n3507), .ZN(n3680) );
  NAND2_X1 U4468 ( .A1(n3680), .A2(n3509), .ZN(n3512) );
  XNOR2_X1 U4469 ( .A(n3512), .B(n4343), .ZN(n5458) );
  NAND2_X1 U4470 ( .A1(n3511), .A2(n3510), .ZN(n5455) );
  NAND2_X1 U4471 ( .A1(n3512), .A2(n4343), .ZN(n3513) );
  NAND2_X1 U4472 ( .A1(n5455), .A2(n3513), .ZN(n5471) );
  INV_X1 U4473 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U4474 ( .A1(n5471), .A2(n3514), .ZN(n3516) );
  NAND2_X1 U4475 ( .A1(n5848), .A2(n6002), .ZN(n3515) );
  NAND2_X1 U4476 ( .A1(n3516), .A2(n3515), .ZN(n5499) );
  INV_X1 U4477 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5987) );
  OAI21_X2 U4478 ( .B1(n5499), .B2(n5502), .A(n5501), .ZN(n5754) );
  INV_X1 U4479 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3518) );
  NAND2_X1 U4480 ( .A1(n5848), .A2(n3518), .ZN(n5752) );
  NAND2_X1 U4481 ( .A1(n5754), .A2(n5752), .ZN(n5750) );
  INV_X1 U4482 ( .A(n5750), .ZN(n3517) );
  AND2_X1 U4483 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4105) );
  NAND2_X1 U4484 ( .A1(n3517), .A2(n4105), .ZN(n5716) );
  INV_X1 U4485 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5851) );
  INV_X1 U4486 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5820) );
  NAND2_X1 U4487 ( .A1(n5750), .A2(n2982), .ZN(n3520) );
  NAND2_X1 U4488 ( .A1(n3520), .A2(n4451), .ZN(n3521) );
  NAND2_X1 U4489 ( .A1(n5716), .A2(n3521), .ZN(n4447) );
  NOR2_X1 U4490 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5825) );
  NOR2_X1 U4491 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3523) );
  INV_X1 U4492 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3522) );
  INV_X1 U4493 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5812) );
  NAND4_X1 U4494 ( .A1(n5825), .A2(n3523), .A3(n3522), .A4(n5812), .ZN(n3524)
         );
  AND2_X1 U4495 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5826) );
  AND2_X1 U4496 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4095) );
  AND2_X1 U4497 ( .A1(n5826), .A2(n4095), .ZN(n5793) );
  AND2_X1 U4498 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4108) );
  NAND2_X1 U4499 ( .A1(n5793), .A2(n4108), .ZN(n3977) );
  NAND2_X1 U4500 ( .A1(n5848), .A2(n3977), .ZN(n3525) );
  OAI21_X1 U4501 ( .B1(n4447), .B2(n2987), .A(n3525), .ZN(n3526) );
  NAND2_X1 U4502 ( .A1(n3526), .A2(n3527), .ZN(n3920) );
  OAI21_X1 U4503 ( .B1(n3527), .B2(n5701), .A(n4289), .ZN(n5778) );
  INV_X1 U4504 ( .A(n5778), .ZN(n3918) );
  NAND2_X1 U4505 ( .A1(n3528), .A2(n3679), .ZN(n3536) );
  INV_X2 U4506 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6514) );
  INV_X1 U4507 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3533) );
  INV_X1 U4508 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U4509 ( .A1(n3590), .A2(n6095), .ZN(n3531) );
  INV_X1 U4510 ( .A(n3619), .ZN(n3530) );
  NAND2_X1 U4511 ( .A1(n3531), .A2(n3530), .ZN(n6100) );
  NAND2_X1 U4512 ( .A1(n6514), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4513 ( .A1(n6100), .A2(n4236), .B1(n4242), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3532) );
  OAI21_X1 U4514 ( .B1(n4304), .B2(n3533), .A(n3532), .ZN(n3534) );
  INV_X1 U4515 ( .A(n3534), .ZN(n3535) );
  NAND2_X1 U4516 ( .A1(n4701), .A2(n3679), .ZN(n3541) );
  AND2_X1 U4517 ( .A1(n3537), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3567) );
  INV_X1 U4518 ( .A(EAX_REG_1__SCAN_IN), .ZN(n3538) );
  OAI22_X1 U4519 ( .A1(n4304), .A2(n3538), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3551), .ZN(n3539) );
  AOI21_X1 U4520 ( .B1(n3567), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3539), 
        .ZN(n3540) );
  NAND2_X1 U4521 ( .A1(n5387), .A2(n3542), .ZN(n3543) );
  NAND2_X1 U4522 ( .A1(n3543), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4592) );
  OR2_X1 U4523 ( .A1(n5540), .A2(n3711), .ZN(n3549) );
  INV_X1 U4524 ( .A(EAX_REG_0__SCAN_IN), .ZN(n3546) );
  INV_X1 U4525 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3545) );
  OAI22_X1 U4526 ( .A1(n4304), .A2(n3546), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3545), .ZN(n3547) );
  AOI21_X1 U4527 ( .B1(n3567), .B2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(n3547), 
        .ZN(n3548) );
  NAND2_X1 U4528 ( .A1(n4591), .A2(n4236), .ZN(n3550) );
  NAND2_X1 U4529 ( .A1(n4552), .A2(n4554), .ZN(n4553) );
  INV_X1 U4530 ( .A(EAX_REG_2__SCAN_IN), .ZN(n3554) );
  AOI21_X1 U4531 ( .B1(n6145), .B2(n3551), .A(n3561), .ZN(n3552) );
  INV_X1 U4532 ( .A(n3552), .ZN(n6292) );
  AOI22_X1 U4533 ( .A1(n6292), .A2(n4236), .B1(n4242), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3553) );
  OAI21_X1 U4534 ( .B1(n4304), .B2(n3554), .A(n3553), .ZN(n3555) );
  AOI21_X1 U4535 ( .B1(n3567), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3555), 
        .ZN(n3556) );
  NAND2_X1 U4536 ( .A1(n4553), .A2(n3556), .ZN(n4587) );
  INV_X1 U4537 ( .A(n4700), .ZN(n3557) );
  NAND2_X1 U4538 ( .A1(n3557), .A2(n3679), .ZN(n3558) );
  NAND2_X1 U4539 ( .A1(n4587), .A2(n4588), .ZN(n3559) );
  INV_X1 U4540 ( .A(EAX_REG_3__SCAN_IN), .ZN(n3563) );
  XNOR2_X1 U4541 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .B(n3561), .ZN(n6133) );
  AOI22_X1 U4542 ( .A1(n4236), .A2(n6133), .B1(n4242), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3562) );
  OAI21_X1 U4543 ( .B1(n4304), .B2(n3563), .A(n3562), .ZN(n3564) );
  AOI21_X1 U4544 ( .B1(n3567), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n3564), 
        .ZN(n3565) );
  INV_X1 U4545 ( .A(n3567), .ZN(n3571) );
  NAND2_X1 U4546 ( .A1(n6514), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3569)
         );
  NAND2_X1 U4547 ( .A1(n4243), .A2(EAX_REG_4__SCAN_IN), .ZN(n3568) );
  OAI211_X1 U4548 ( .C1(n3571), .C2(n3570), .A(n3569), .B(n3568), .ZN(n3574)
         );
  OAI21_X1 U4549 ( .B1(n3572), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3579), 
        .ZN(n6122) );
  AND2_X1 U4550 ( .A1(n6122), .A2(n4236), .ZN(n3573) );
  AOI21_X1 U4551 ( .B1(n3574), .B2(n4248), .A(n3573), .ZN(n3575) );
  NAND2_X1 U4552 ( .A1(n3576), .A2(n3575), .ZN(n4577) );
  INV_X1 U4553 ( .A(n3577), .ZN(n3578) );
  AND2_X1 U4554 ( .A1(n3579), .A2(n6111), .ZN(n3580) );
  OR2_X1 U4555 ( .A1(n3580), .A2(n3588), .ZN(n6117) );
  NAND2_X1 U4556 ( .A1(n6117), .A2(n4236), .ZN(n3581) );
  OAI21_X1 U4557 ( .B1(n6111), .B2(n3885), .A(n3581), .ZN(n3582) );
  AOI21_X1 U4558 ( .B1(n4243), .B2(EAX_REG_5__SCAN_IN), .A(n3582), .ZN(n3583)
         );
  NAND2_X1 U4559 ( .A1(n3584), .A2(n3583), .ZN(n4649) );
  NAND2_X1 U4560 ( .A1(n3468), .A2(n3586), .ZN(n3594) );
  INV_X1 U4561 ( .A(EAX_REG_6__SCAN_IN), .ZN(n5048) );
  INV_X1 U4562 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3587) );
  OAI22_X1 U4563 ( .A1(n4304), .A2(n5048), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3587), .ZN(n3592) );
  OR2_X1 U4564 ( .A1(n3588), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3589) );
  NAND2_X1 U4565 ( .A1(n3590), .A2(n3589), .ZN(n6105) );
  AND2_X1 U4566 ( .A1(n6105), .A2(n4236), .ZN(n3591) );
  AOI21_X1 U4567 ( .B1(n3592), .B2(n4248), .A(n3591), .ZN(n3593) );
  NAND2_X1 U4568 ( .A1(n3594), .A2(n3593), .ZN(n5043) );
  NAND2_X1 U4569 ( .A1(n4711), .A2(n4708), .ZN(n4709) );
  AOI22_X1 U4570 ( .A1(n4215), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4132), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4571 ( .A1(n4664), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4572 ( .A1(n4141), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4573 ( .A1(n4224), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3595) );
  NAND4_X1 U4574 ( .A1(n3598), .A2(n3597), .A3(n3596), .A4(n3595), .ZN(n3604)
         );
  AOI22_X1 U4575 ( .A1(n3661), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3602) );
  AOI22_X1 U4576 ( .A1(n4195), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4190), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3601) );
  AOI22_X1 U4577 ( .A1(n4214), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3248), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3600) );
  AOI22_X1 U4578 ( .A1(n3242), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3599) );
  NAND4_X1 U4579 ( .A1(n3602), .A2(n3601), .A3(n3600), .A4(n3599), .ZN(n3603)
         );
  OAI21_X1 U4580 ( .B1(n3604), .B2(n3603), .A(n3679), .ZN(n3607) );
  XOR2_X1 U4581 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3619), .Z(n5613) );
  INV_X1 U4582 ( .A(n5613), .ZN(n5314) );
  AOI22_X1 U4583 ( .A1(n4236), .A2(n5314), .B1(n4242), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3606) );
  NAND2_X1 U4584 ( .A1(n4243), .A2(EAX_REG_8__SCAN_IN), .ZN(n3605) );
  NOR2_X2 U4585 ( .A1(n4709), .A2(n4745), .ZN(n4743) );
  INV_X1 U4586 ( .A(EAX_REG_9__SCAN_IN), .ZN(n3623) );
  AOI22_X1 U4587 ( .A1(n4215), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U4588 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4664), .B1(n3242), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3610) );
  AOI22_X1 U4589 ( .A1(n4190), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3609) );
  AOI22_X1 U4590 ( .A1(n4213), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3248), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3608) );
  NAND4_X1 U4591 ( .A1(n3611), .A2(n3610), .A3(n3609), .A4(n3608), .ZN(n3617)
         );
  AOI22_X1 U4592 ( .A1(n3661), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4593 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n4195), .B1(n4132), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4594 ( .A1(n4214), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3613) );
  AOI22_X1 U4595 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n4225), .B1(n3249), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3612) );
  NAND4_X1 U4596 ( .A1(n3615), .A2(n3614), .A3(n3613), .A4(n3612), .ZN(n3616)
         );
  OR2_X1 U4597 ( .A1(n3617), .A2(n3616), .ZN(n3618) );
  NAND2_X1 U4598 ( .A1(n3679), .A2(n3618), .ZN(n3622) );
  INV_X1 U4599 ( .A(n3624), .ZN(n3620) );
  XNOR2_X1 U4600 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3620), .ZN(n5189) );
  AOI22_X1 U4601 ( .A1(n4236), .A2(n5189), .B1(n4242), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3621) );
  OAI211_X1 U4602 ( .C1(n4304), .C2(n3623), .A(n3622), .B(n3621), .ZN(n4876)
         );
  NAND2_X1 U4603 ( .A1(n4743), .A2(n4876), .ZN(n4874) );
  XOR2_X1 U4604 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3641), .Z(n5296) );
  INV_X1 U4605 ( .A(n5296), .ZN(n5082) );
  AOI22_X1 U4606 ( .A1(n3661), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3628) );
  AOI22_X1 U4607 ( .A1(n4664), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3627) );
  AOI22_X1 U4608 ( .A1(n4224), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4609 ( .A1(n4215), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3248), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3625) );
  NAND4_X1 U4610 ( .A1(n3628), .A2(n3627), .A3(n3626), .A4(n3625), .ZN(n3634)
         );
  AOI22_X1 U4611 ( .A1(n4141), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3632) );
  AOI22_X1 U4612 ( .A1(n4195), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4132), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3631) );
  AOI22_X1 U4613 ( .A1(n4190), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4614 ( .A1(n4225), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3629) );
  NAND4_X1 U4615 ( .A1(n3632), .A2(n3631), .A3(n3630), .A4(n3629), .ZN(n3633)
         );
  NOR2_X1 U4616 ( .A1(n3634), .A2(n3633), .ZN(n3637) );
  NAND2_X1 U4617 ( .A1(n4243), .A2(EAX_REG_10__SCAN_IN), .ZN(n3636) );
  NAND2_X1 U4618 ( .A1(n4242), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3635)
         );
  OAI211_X1 U4619 ( .C1(n3711), .C2(n3637), .A(n3636), .B(n3635), .ZN(n3638)
         );
  AOI21_X1 U4620 ( .B1(n5082), .B2(n4236), .A(n3638), .ZN(n4961) );
  NAND2_X1 U4621 ( .A1(n3641), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3657)
         );
  XNOR2_X1 U4622 ( .A(n3657), .B(n5273), .ZN(n5277) );
  AOI22_X1 U4623 ( .A1(n4214), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4624 ( .A1(n4195), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4132), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4625 ( .A1(n4213), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4626 ( .A1(n3249), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3642) );
  NAND4_X1 U4627 ( .A1(n3645), .A2(n3644), .A3(n3643), .A4(n3642), .ZN(n3652)
         );
  AOI22_X1 U4628 ( .A1(n3661), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4215), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3650) );
  AOI22_X1 U4629 ( .A1(n4664), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3649) );
  AOI22_X1 U4630 ( .A1(n4224), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4190), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3648) );
  AOI22_X1 U4631 ( .A1(n4141), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3248), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3647) );
  NAND4_X1 U4632 ( .A1(n3650), .A2(n3649), .A3(n3648), .A4(n3647), .ZN(n3651)
         );
  NOR2_X1 U4633 ( .A1(n3652), .A2(n3651), .ZN(n3655) );
  NAND2_X1 U4634 ( .A1(n4243), .A2(EAX_REG_11__SCAN_IN), .ZN(n3654) );
  NAND2_X1 U4635 ( .A1(n4242), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3653)
         );
  OAI211_X1 U4636 ( .C1(n3711), .C2(n3655), .A(n3654), .B(n3653), .ZN(n3656)
         );
  AOI21_X1 U4637 ( .B1(n5277), .B2(n4236), .A(n3656), .ZN(n5037) );
  NOR2_X2 U4638 ( .A1(n4962), .A2(n5037), .ZN(n5036) );
  XOR2_X1 U4639 ( .A(n6081), .B(n3674), .Z(n6078) );
  NAND2_X1 U4640 ( .A1(n6078), .A2(n4236), .ZN(n3660) );
  INV_X1 U4641 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5161) );
  OAI21_X1 U4642 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6015), .A(n6514), 
        .ZN(n3658) );
  OAI21_X1 U4643 ( .B1(n4304), .B2(n5161), .A(n3658), .ZN(n3659) );
  NAND2_X1 U4644 ( .A1(n3660), .A2(n3659), .ZN(n3673) );
  AOI22_X1 U4645 ( .A1(n3661), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3665) );
  AOI22_X1 U4646 ( .A1(n4664), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3664) );
  AOI22_X1 U4647 ( .A1(n4214), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4648 ( .A1(n3264), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3662) );
  NAND4_X1 U4649 ( .A1(n3665), .A2(n3664), .A3(n3663), .A4(n3662), .ZN(n3671)
         );
  AOI22_X1 U4650 ( .A1(n4141), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4651 ( .A1(n4215), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4652 ( .A1(n4195), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4190), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4653 ( .A1(n4213), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3248), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3666) );
  NAND4_X1 U4654 ( .A1(n3669), .A2(n3668), .A3(n3667), .A4(n3666), .ZN(n3670)
         );
  OAI21_X1 U4655 ( .B1(n3671), .B2(n3670), .A(n3679), .ZN(n3672) );
  NAND2_X1 U4656 ( .A1(n3673), .A2(n3672), .ZN(n5159) );
  NAND2_X1 U4657 ( .A1(n5036), .A2(n5159), .ZN(n5157) );
  OAI21_X1 U4658 ( .B1(n3675), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n3697), 
        .ZN(n6076) );
  NAND2_X1 U4659 ( .A1(n6076), .A2(n4236), .ZN(n3677) );
  AOI22_X1 U4660 ( .A1(n4243), .A2(EAX_REG_13__SCAN_IN), .B1(n4242), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3676) );
  NAND2_X1 U4661 ( .A1(n3677), .A2(n3676), .ZN(n3678) );
  XOR2_X1 U4662 ( .A(n6058), .B(n3697), .Z(n6061) );
  INV_X1 U4663 ( .A(n6061), .ZN(n5475) );
  AOI22_X1 U4664 ( .A1(n3661), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4665 ( .A1(n4664), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4132), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4666 ( .A1(n4141), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3684) );
  AOI22_X1 U4667 ( .A1(n4225), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3683) );
  NAND4_X1 U4668 ( .A1(n3686), .A2(n3685), .A3(n3684), .A4(n3683), .ZN(n3692)
         );
  AOI22_X1 U4669 ( .A1(n4195), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4215), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4670 ( .A1(n4214), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4190), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4671 ( .A1(n3242), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3248), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4672 ( .A1(n4224), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3687) );
  NAND4_X1 U4673 ( .A1(n3690), .A2(n3689), .A3(n3688), .A4(n3687), .ZN(n3691)
         );
  NOR2_X1 U4674 ( .A1(n3692), .A2(n3691), .ZN(n3695) );
  NAND2_X1 U4675 ( .A1(n4243), .A2(EAX_REG_14__SCAN_IN), .ZN(n3694) );
  NAND2_X1 U4676 ( .A1(n4242), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3693)
         );
  OAI211_X1 U4677 ( .C1(n3711), .C2(n3695), .A(n3694), .B(n3693), .ZN(n3696)
         );
  AOI21_X1 U4678 ( .B1(n5475), .B2(n4236), .A(n3696), .ZN(n5339) );
  NOR2_X2 U4679 ( .A1(n5285), .A2(n5339), .ZN(n5337) );
  XNOR2_X1 U4680 ( .A(n3714), .B(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5506)
         );
  AOI22_X1 U4681 ( .A1(n3661), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3701) );
  AOI22_X1 U4682 ( .A1(n4215), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3700) );
  AOI22_X1 U4683 ( .A1(n4195), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4190), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U4684 ( .A1(n4214), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3248), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3698) );
  NAND4_X1 U4685 ( .A1(n3701), .A2(n3700), .A3(n3699), .A4(n3698), .ZN(n3707)
         );
  AOI22_X1 U4686 ( .A1(n4224), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4687 ( .A1(n4664), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4688 ( .A1(n4141), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4689 ( .A1(n3264), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3702) );
  NAND4_X1 U4690 ( .A1(n3705), .A2(n3704), .A3(n3703), .A4(n3702), .ZN(n3706)
         );
  NOR2_X1 U4691 ( .A1(n3707), .A2(n3706), .ZN(n3710) );
  NAND2_X1 U4692 ( .A1(n4243), .A2(EAX_REG_15__SCAN_IN), .ZN(n3709) );
  NAND2_X1 U4693 ( .A1(n4242), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3708)
         );
  OAI211_X1 U4694 ( .C1(n3711), .C2(n3710), .A(n3709), .B(n3708), .ZN(n3712)
         );
  AOI21_X1 U4695 ( .B1(n5506), .B2(n4236), .A(n3712), .ZN(n5439) );
  XOR2_X1 U4696 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3731), .Z(n6050) );
  NAND2_X1 U4697 ( .A1(n3183), .A2(n3956), .ZN(n3715) );
  AOI22_X1 U4698 ( .A1(n3661), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4699 ( .A1(n4215), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4700 ( .A1(n4141), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4701 ( .A1(n3230), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3716) );
  NAND4_X1 U4702 ( .A1(n3719), .A2(n3718), .A3(n3717), .A4(n3716), .ZN(n3725)
         );
  AOI22_X1 U4703 ( .A1(n4195), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4664), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4704 ( .A1(n4225), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3264), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4705 ( .A1(n4213), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4706 ( .A1(n4214), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3248), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3720) );
  NAND4_X1 U4707 ( .A1(n3723), .A2(n3722), .A3(n3721), .A4(n3720), .ZN(n3724)
         );
  OR2_X1 U4708 ( .A1(n3725), .A2(n3724), .ZN(n3729) );
  INV_X1 U4709 ( .A(EAX_REG_16__SCAN_IN), .ZN(n3727) );
  INV_X1 U4710 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3726) );
  OAI22_X1 U4711 ( .A1(n4304), .A2(n3727), .B1(n3885), .B2(n3726), .ZN(n3728)
         );
  AOI21_X1 U4712 ( .B1(n4207), .B2(n3729), .A(n3728), .ZN(n3730) );
  OAI21_X1 U4713 ( .B1(n6050), .B2(n4248), .A(n3730), .ZN(n5479) );
  XNOR2_X1 U4714 ( .A(n3762), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5960)
         );
  AOI22_X1 U4715 ( .A1(n3661), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4716 ( .A1(n4141), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3734) );
  AOI22_X1 U4717 ( .A1(n3823), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3733) );
  AOI22_X1 U4718 ( .A1(n4213), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3235), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3732) );
  NAND4_X1 U4719 ( .A1(n3735), .A2(n3734), .A3(n3733), .A4(n3732), .ZN(n3741)
         );
  INV_X1 U4720 ( .A(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4422) );
  AOI22_X1 U4721 ( .A1(n4195), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4664), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4722 ( .A1(n4215), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4723 ( .A1(n4225), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4724 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n4132), .B1(n3230), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3736) );
  NAND4_X1 U4725 ( .A1(n3739), .A2(n3738), .A3(n3737), .A4(n3736), .ZN(n3740)
         );
  OR2_X1 U4726 ( .A1(n3741), .A2(n3740), .ZN(n3745) );
  INV_X1 U4727 ( .A(EAX_REG_17__SCAN_IN), .ZN(n3743) );
  OAI21_X1 U4728 ( .B1(n6015), .B2(PHYADDRPOINTER_REG_17__SCAN_IN), .A(n6514), 
        .ZN(n3742) );
  OAI21_X1 U4729 ( .B1(n4304), .B2(n3743), .A(n3742), .ZN(n3744) );
  AOI21_X1 U4730 ( .B1(n4207), .B2(n3745), .A(n3744), .ZN(n3746) );
  AOI21_X1 U4731 ( .B1(n5960), .B2(n4236), .A(n3746), .ZN(n5486) );
  AOI22_X1 U4732 ( .A1(n4213), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3750) );
  AOI22_X1 U4733 ( .A1(n4214), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3749) );
  AOI22_X1 U4734 ( .A1(n3823), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4735 ( .A1(n4664), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3747) );
  NAND4_X1 U4736 ( .A1(n3750), .A2(n3749), .A3(n3748), .A4(n3747), .ZN(n3756)
         );
  AOI22_X1 U4737 ( .A1(n3661), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3754) );
  AOI22_X1 U4738 ( .A1(n4215), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4739 ( .A1(n3264), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3235), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4740 ( .A1(n4195), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3230), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3751) );
  NAND4_X1 U4741 ( .A1(n3754), .A2(n3753), .A3(n3752), .A4(n3751), .ZN(n3755)
         );
  NOR2_X1 U4742 ( .A1(n3756), .A2(n3755), .ZN(n3761) );
  INV_X1 U4743 ( .A(EAX_REG_18__SCAN_IN), .ZN(n3758) );
  NAND2_X1 U4744 ( .A1(n6514), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3757)
         );
  OAI211_X1 U4745 ( .C1(n4304), .C2(n3758), .A(n4248), .B(n3757), .ZN(n3759)
         );
  INV_X1 U4746 ( .A(n3759), .ZN(n3760) );
  OAI21_X1 U4747 ( .B1(n4239), .B2(n3761), .A(n3760), .ZN(n3765) );
  INV_X1 U4748 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5490) );
  OAI21_X1 U4749 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n3763), .A(n3800), 
        .ZN(n6044) );
  OR2_X1 U4750 ( .A1(n4248), .A2(n6044), .ZN(n3764) );
  NAND2_X1 U4751 ( .A1(n3765), .A2(n3764), .ZN(n5513) );
  AOI22_X1 U4752 ( .A1(n3661), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4753 ( .A1(n4141), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4754 ( .A1(n3823), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3769) );
  AOI22_X1 U4755 ( .A1(n4213), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3235), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3768) );
  NAND4_X1 U4756 ( .A1(n3771), .A2(n3770), .A3(n3769), .A4(n3768), .ZN(n3777)
         );
  AOI22_X1 U4757 ( .A1(n4195), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4664), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4758 ( .A1(n4215), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4759 ( .A1(n4225), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4760 ( .A1(n3264), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3772) );
  NAND4_X1 U4761 ( .A1(n3775), .A2(n3774), .A3(n3773), .A4(n3772), .ZN(n3776)
         );
  NOR2_X1 U4762 ( .A1(n3777), .A2(n3776), .ZN(n3780) );
  NAND2_X1 U4763 ( .A1(n4243), .A2(EAX_REG_19__SCAN_IN), .ZN(n3779) );
  OAI21_X1 U4764 ( .B1(n6015), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6514), 
        .ZN(n3778) );
  OAI211_X1 U4765 ( .C1(n4239), .C2(n3780), .A(n3779), .B(n3778), .ZN(n3782)
         );
  XNOR2_X1 U4766 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n3800), .ZN(n5923)
         );
  NAND2_X1 U4767 ( .A1(n4236), .A2(n5923), .ZN(n3781) );
  NAND2_X1 U4768 ( .A1(n3782), .A2(n3781), .ZN(n5521) );
  AOI22_X1 U4769 ( .A1(n4195), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4664), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4770 ( .A1(n4215), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4771 ( .A1(n4141), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4772 ( .A1(n3264), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3785) );
  NAND4_X1 U4773 ( .A1(n3788), .A2(n3787), .A3(n3786), .A4(n3785), .ZN(n3794)
         );
  AOI22_X1 U4774 ( .A1(n4218), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4775 ( .A1(n3229), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3248), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4776 ( .A1(n4225), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3230), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4777 ( .A1(n4224), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3789) );
  NAND4_X1 U4778 ( .A1(n3792), .A2(n3791), .A3(n3790), .A4(n3789), .ZN(n3793)
         );
  NOR2_X1 U4779 ( .A1(n3794), .A2(n3793), .ZN(n3799) );
  INV_X1 U4780 ( .A(EAX_REG_20__SCAN_IN), .ZN(n3796) );
  NAND2_X1 U4781 ( .A1(n6514), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3795)
         );
  OAI211_X1 U4782 ( .C1(n4304), .C2(n3796), .A(n4248), .B(n3795), .ZN(n3797)
         );
  INV_X1 U4783 ( .A(n3797), .ZN(n3798) );
  OAI21_X1 U4784 ( .B1(n4239), .B2(n3799), .A(n3798), .ZN(n3803) );
  INV_X1 U4785 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5745) );
  OAI21_X1 U4786 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n3801), .A(n3834), 
        .ZN(n5954) );
  OR2_X1 U4787 ( .A1(n4248), .A2(n5954), .ZN(n3802) );
  NAND2_X1 U4788 ( .A1(n3803), .A2(n3802), .ZN(n5659) );
  NOR2_X2 U4789 ( .A1(n5519), .A2(n5659), .ZN(n5650) );
  AOI22_X1 U4790 ( .A1(n4218), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4215), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4791 ( .A1(n4195), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4664), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4792 ( .A1(n4225), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4132), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4793 ( .A1(n3823), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3248), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3804) );
  NAND4_X1 U4794 ( .A1(n3807), .A2(n3806), .A3(n3805), .A4(n3804), .ZN(n3813)
         );
  AOI22_X1 U4795 ( .A1(n4213), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4796 ( .A1(n4214), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4797 ( .A1(n4224), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4798 ( .A1(n3249), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3808) );
  NAND4_X1 U4799 ( .A1(n3811), .A2(n3810), .A3(n3809), .A4(n3808), .ZN(n3812)
         );
  NOR2_X1 U4800 ( .A1(n3813), .A2(n3812), .ZN(n3816) );
  INV_X1 U4801 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5902) );
  OAI21_X1 U4802 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5902), .A(n4248), .ZN(
        n3814) );
  AOI21_X1 U4803 ( .B1(n4243), .B2(EAX_REG_21__SCAN_IN), .A(n3814), .ZN(n3815)
         );
  OAI21_X1 U4804 ( .B1(n4239), .B2(n3816), .A(n3815), .ZN(n3818) );
  XNOR2_X1 U4805 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n3834), .ZN(n5905)
         );
  NAND2_X1 U4806 ( .A1(n4236), .A2(n5905), .ZN(n3817) );
  NAND2_X1 U4807 ( .A1(n5650), .A2(n5652), .ZN(n5597) );
  AOI22_X1 U4808 ( .A1(n4224), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4132), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4809 ( .A1(n4218), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4810 ( .A1(n4215), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4811 ( .A1(n4664), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3819) );
  NAND4_X1 U4812 ( .A1(n3822), .A2(n3821), .A3(n3820), .A4(n3819), .ZN(n3829)
         );
  AOI22_X1 U4813 ( .A1(n3242), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4814 ( .A1(n4141), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4815 ( .A1(n3248), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4816 ( .A1(n4133), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3824) );
  NAND4_X1 U4817 ( .A1(n3827), .A2(n3826), .A3(n3825), .A4(n3824), .ZN(n3828)
         );
  NOR2_X1 U4818 ( .A1(n3829), .A2(n3828), .ZN(n3833) );
  INV_X1 U4819 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4638) );
  OAI21_X1 U4820 ( .B1(PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6015), .A(n6514), 
        .ZN(n3830) );
  OAI21_X1 U4821 ( .B1(n4304), .B2(n4638), .A(n3830), .ZN(n3831) );
  INV_X1 U4822 ( .A(n3831), .ZN(n3832) );
  OAI21_X1 U4823 ( .B1(n4239), .B2(n3833), .A(n3832), .ZN(n3842) );
  INV_X1 U4824 ( .A(n3881), .ZN(n3840) );
  INV_X1 U4825 ( .A(n3836), .ZN(n3838) );
  INV_X1 U4826 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3837) );
  NAND2_X1 U4827 ( .A1(n3838), .A2(n3837), .ZN(n3839) );
  NAND2_X1 U4828 ( .A1(n3840), .A2(n3839), .ZN(n5728) );
  NAND2_X1 U4829 ( .A1(n3842), .A2(n3841), .ZN(n5601) );
  AOI22_X1 U4830 ( .A1(n3661), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4831 ( .A1(n4664), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4132), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4832 ( .A1(n4190), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4833 ( .A1(n4224), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3843) );
  NAND4_X1 U4834 ( .A1(n3846), .A2(n3845), .A3(n3844), .A4(n3843), .ZN(n3852)
         );
  AOI22_X1 U4835 ( .A1(n4215), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4836 ( .A1(n3242), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4837 ( .A1(n4141), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3235), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4838 ( .A1(n4133), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3847) );
  NAND4_X1 U4839 ( .A1(n3850), .A2(n3849), .A3(n3848), .A4(n3847), .ZN(n3851)
         );
  NOR2_X1 U4840 ( .A1(n3852), .A2(n3851), .ZN(n3869) );
  AOI22_X1 U4841 ( .A1(n3661), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4842 ( .A1(n4215), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4843 ( .A1(n4213), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3248), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4844 ( .A1(n4132), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3230), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3853) );
  NAND4_X1 U4845 ( .A1(n3856), .A2(n3855), .A3(n3854), .A4(n3853), .ZN(n3862)
         );
  AOI22_X1 U4846 ( .A1(n4133), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4664), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4847 ( .A1(n4214), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4190), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4848 ( .A1(n4224), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4849 ( .A1(n3242), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3857) );
  NAND4_X1 U4850 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(n3861)
         );
  NOR2_X1 U4851 ( .A1(n3862), .A2(n3861), .ZN(n3870) );
  XNOR2_X1 U4852 ( .A(n3869), .B(n3870), .ZN(n3865) );
  INV_X1 U4853 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5901) );
  OAI21_X1 U4854 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5901), .A(n4248), .ZN(
        n3863) );
  AOI21_X1 U4855 ( .B1(n4243), .B2(EAX_REG_23__SCAN_IN), .A(n3863), .ZN(n3864)
         );
  OAI21_X1 U4856 ( .B1(n4239), .B2(n3865), .A(n3864), .ZN(n3867) );
  XNOR2_X1 U4857 ( .A(n3881), .B(n5901), .ZN(n5891) );
  NAND2_X1 U4858 ( .A1(n5891), .A2(n4236), .ZN(n3866) );
  NAND2_X1 U4859 ( .A1(n3867), .A2(n3866), .ZN(n5644) );
  INV_X1 U4860 ( .A(n5644), .ZN(n3868) );
  OR2_X1 U4861 ( .A1(n3870), .A2(n3869), .ZN(n3900) );
  AOI22_X1 U4862 ( .A1(n4224), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3264), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4863 ( .A1(n4215), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4864 ( .A1(n4133), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4865 ( .A1(n4213), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3871) );
  NAND4_X1 U4866 ( .A1(n3874), .A2(n3873), .A3(n3872), .A4(n3871), .ZN(n3880)
         );
  AOI22_X1 U4867 ( .A1(n4141), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4868 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n3229), .B1(n3249), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4869 ( .A1(n3661), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4870 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n4664), .B1(n3235), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3875) );
  NAND4_X1 U4871 ( .A1(n3878), .A2(n3877), .A3(n3876), .A4(n3875), .ZN(n3879)
         );
  NOR2_X1 U4872 ( .A1(n3880), .A2(n3879), .ZN(n3899) );
  XNOR2_X1 U4873 ( .A(n3900), .B(n3899), .ZN(n3888) );
  INV_X1 U4874 ( .A(n3883), .ZN(n3882) );
  INV_X1 U4875 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4457) );
  NAND2_X1 U4876 ( .A1(n3882), .A2(n4457), .ZN(n3884) );
  OAI22_X1 U4877 ( .A1(n5884), .A2(n4248), .B1(n4457), .B2(n3885), .ZN(n3886)
         );
  AOI21_X1 U4878 ( .B1(n4243), .B2(EAX_REG_24__SCAN_IN), .A(n3886), .ZN(n3887)
         );
  OAI21_X1 U4879 ( .B1(n4239), .B2(n3888), .A(n3887), .ZN(n4456) );
  AOI22_X1 U4880 ( .A1(n4133), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4664), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4881 ( .A1(n3661), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4215), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4882 ( .A1(n4141), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3235), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4883 ( .A1(n3242), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3230), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3889) );
  NAND4_X1 U4884 ( .A1(n3892), .A2(n3891), .A3(n3890), .A4(n3889), .ZN(n3898)
         );
  AOI22_X1 U4885 ( .A1(n4213), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4886 ( .A1(n4225), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4132), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4887 ( .A1(n3823), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4888 ( .A1(n4214), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3893) );
  NAND4_X1 U4889 ( .A1(n3896), .A2(n3895), .A3(n3894), .A4(n3893), .ZN(n3897)
         );
  OR2_X1 U4890 ( .A1(n3898), .A2(n3897), .ZN(n4126) );
  NOR2_X1 U4891 ( .A1(n3900), .A2(n3899), .ZN(n4125) );
  XOR2_X1 U4892 ( .A(n4126), .B(n4125), .Z(n3901) );
  NAND2_X1 U4893 ( .A1(n3901), .A2(n4207), .ZN(n3905) );
  INV_X1 U4894 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4503) );
  OAI21_X1 U4895 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4503), .A(n4248), .ZN(
        n3902) );
  AOI21_X1 U4896 ( .B1(n4243), .B2(EAX_REG_25__SCAN_IN), .A(n3902), .ZN(n3904)
         );
  XNOR2_X1 U4897 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .B(n4157), .ZN(n4501)
         );
  AND2_X1 U4898 ( .A1(n4236), .A2(n4501), .ZN(n3903) );
  AOI21_X1 U4899 ( .B1(n3905), .B2(n3904), .A(n3903), .ZN(n4187) );
  NAND3_X1 U4900 ( .A1(n6615), .A2(STATE2_REG_1__SCAN_IN), .A3(
        STATEBS16_REG_SCAN_IN), .ZN(n6623) );
  INV_X1 U4901 ( .A(n6623), .ZN(n3907) );
  NAND2_X1 U4902 ( .A1(n3907), .A2(n6389), .ZN(n6301) );
  INV_X1 U4903 ( .A(n6389), .ZN(n6352) );
  NAND2_X1 U4904 ( .A1(n6352), .A2(n3908), .ZN(n6728) );
  NAND2_X1 U4905 ( .A1(n6728), .A2(n6615), .ZN(n3909) );
  NAND2_X1 U4906 ( .A1(n6615), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3911) );
  NAND2_X1 U4907 ( .A1(n6015), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3910) );
  NAND2_X1 U4908 ( .A1(n3911), .A2(n3910), .ZN(n6297) );
  INV_X1 U4909 ( .A(n6297), .ZN(n3912) );
  NAND2_X1 U4910 ( .A1(n5961), .A2(n4501), .ZN(n3914) );
  AOI22_X1 U4911 ( .A1(n6298), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .B1(n6284), 
        .B2(REIP_REG_25__SCAN_IN), .ZN(n3913) );
  OAI21_X1 U4912 ( .B1(n5548), .B2(n6301), .A(n3915), .ZN(n3916) );
  INV_X1 U4913 ( .A(n3916), .ZN(n3917) );
  OAI21_X1 U4914 ( .B1(n6016), .B2(n3918), .A(n3917), .ZN(U2961) );
  INV_X1 U4915 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5967) );
  AND2_X2 U4916 ( .A1(n3920), .A2(n3919), .ZN(n4439) );
  INV_X1 U4917 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5974) );
  INV_X1 U4918 ( .A(n4463), .ZN(n3922) );
  NOR3_X1 U4919 ( .A1(n5699), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4287) );
  NAND2_X1 U4920 ( .A1(n3921), .A2(n4287), .ZN(n4464) );
  NAND2_X1 U4921 ( .A1(n3922), .A2(n4464), .ZN(n3923) );
  XNOR2_X1 U4922 ( .A(n3923), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5697)
         );
  INV_X1 U4923 ( .A(n4625), .ZN(n4750) );
  INV_X1 U4924 ( .A(n3925), .ZN(n3926) );
  AND2_X1 U4925 ( .A1(n3926), .A2(n6631), .ZN(n6638) );
  INV_X1 U4926 ( .A(n6638), .ZN(n4559) );
  NAND2_X1 U4927 ( .A1(n4802), .A2(n4559), .ZN(n4259) );
  NAND3_X1 U4928 ( .A1(n4599), .A2(n4259), .A3(n6729), .ZN(n3927) );
  NAND3_X1 U4929 ( .A1(n3927), .A2(n4628), .A3(n3282), .ZN(n3928) );
  NAND2_X1 U4930 ( .A1(n3928), .A2(n2973), .ZN(n3950) );
  NAND3_X1 U4931 ( .A1(n4606), .A2(n5541), .A3(n3189), .ZN(n3947) );
  AOI21_X1 U4932 ( .B1(n3930), .B2(n4813), .A(n3974), .ZN(n3931) );
  NAND2_X1 U4933 ( .A1(n3929), .A2(n3931), .ZN(n3954) );
  NAND3_X1 U4934 ( .A1(n3932), .A2(n4628), .A3(n4755), .ZN(n3934) );
  NAND2_X1 U4935 ( .A1(n2969), .A2(n6731), .ZN(n3933) );
  NAND2_X1 U4936 ( .A1(n3934), .A2(n3933), .ZN(n3961) );
  OR2_X1 U4937 ( .A1(n3954), .A2(n3961), .ZN(n3936) );
  NAND2_X1 U4938 ( .A1(n3936), .A2(n4256), .ZN(n4562) );
  NAND2_X1 U4939 ( .A1(n3192), .A2(n4559), .ZN(n3945) );
  INV_X1 U4940 ( .A(n3937), .ZN(n3944) );
  INV_X1 U4941 ( .A(n3938), .ZN(n3940) );
  NAND4_X1 U4942 ( .A1(n3942), .A2(n3941), .A3(n3940), .A4(n3939), .ZN(n3943)
         );
  NAND2_X1 U4943 ( .A1(n3944), .A2(n3943), .ZN(n4517) );
  NOR2_X1 U4944 ( .A1(READY_N), .A2(n4517), .ZN(n4746) );
  NAND3_X1 U4945 ( .A1(n3945), .A2(n4746), .A3(n3204), .ZN(n3946) );
  NAND3_X1 U4946 ( .A1(n3947), .A2(n4562), .A3(n3946), .ZN(n3948) );
  INV_X1 U4947 ( .A(n6598), .ZN(n6612) );
  INV_X1 U4948 ( .A(n3952), .ZN(n6590) );
  NAND2_X1 U4949 ( .A1(n3192), .A2(n3953), .ZN(n3978) );
  NAND2_X1 U4950 ( .A1(n4599), .A2(n4557), .ZN(n4534) );
  AND2_X1 U4951 ( .A1(n6590), .A2(n4534), .ZN(n3958) );
  INV_X1 U4952 ( .A(n5171), .ZN(n4513) );
  NAND2_X1 U4953 ( .A1(n3955), .A2(n3956), .ZN(n3957) );
  NAND4_X1 U4954 ( .A1(n4748), .A2(n3958), .A3(n4749), .A4(n3957), .ZN(n3959)
         );
  INV_X1 U4955 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4343) );
  NAND2_X1 U4956 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5465) );
  NOR2_X1 U4957 ( .A1(n4343), .A2(n5465), .ZN(n6003) );
  NAND2_X1 U4958 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6003), .ZN(n5985) );
  NAND2_X1 U4959 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5980) );
  NOR2_X1 U4960 ( .A1(n5985), .A2(n5980), .ZN(n4102) );
  NOR2_X1 U4961 ( .A1(n4012), .A2(n3475), .ZN(n5031) );
  NAND3_X1 U4962 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n5031), .ZN(n3976) );
  INV_X1 U4963 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4845) );
  NAND2_X1 U4964 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4840) );
  NAND2_X1 U4965 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4841) );
  NOR4_X1 U4966 ( .A1(n4005), .A2(n4845), .A3(n4840), .A4(n4841), .ZN(n4866)
         );
  INV_X1 U4967 ( .A(n4866), .ZN(n3960) );
  NOR2_X1 U4968 ( .A1(n3976), .A2(n3960), .ZN(n4099) );
  NOR2_X1 U4969 ( .A1(n4256), .A2(n4802), .ZN(n5537) );
  NAND2_X1 U4970 ( .A1(n4097), .A2(n5537), .ZN(n5464) );
  INV_X4 U4971 ( .A(n5515), .ZN(n5662) );
  INV_X1 U4972 ( .A(n3961), .ZN(n3965) );
  NAND2_X1 U4973 ( .A1(n4822), .A2(n4628), .ZN(n4011) );
  INV_X1 U4974 ( .A(n4542), .ZN(n4086) );
  OAI21_X1 U4975 ( .B1(n2973), .B2(n3282), .A(n4514), .ZN(n3962) );
  NAND2_X1 U4976 ( .A1(n4086), .A2(n3962), .ZN(n3963) );
  NAND2_X1 U4977 ( .A1(n3963), .A2(n3974), .ZN(n3964) );
  OAI211_X1 U4978 ( .C1(n5662), .C2(n3929), .A(n3965), .B(n3964), .ZN(n3966)
         );
  INV_X1 U4979 ( .A(n3966), .ZN(n3967) );
  AND2_X1 U4980 ( .A1(n3968), .A2(n3967), .ZN(n4602) );
  OAI22_X1 U4981 ( .A1(n4597), .A2(n3969), .B1(n4596), .B2(n4628), .ZN(n3970)
         );
  INV_X1 U4982 ( .A(n3970), .ZN(n3972) );
  NOR2_X1 U4983 ( .A1(n3213), .A2(n4628), .ZN(n3971) );
  NAND2_X1 U4984 ( .A1(n5541), .A2(n3971), .ZN(n4681) );
  NAND3_X1 U4985 ( .A1(n4602), .A2(n3972), .A3(n4681), .ZN(n3973) );
  NAND2_X1 U4986 ( .A1(n4097), .A2(n3973), .ZN(n5995) );
  INV_X1 U4987 ( .A(n5464), .ZN(n4093) );
  NOR2_X1 U4988 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n4093), .ZN(n4618)
         );
  NAND2_X1 U4989 ( .A1(n4099), .A2(n4716), .ZN(n5817) );
  NOR2_X1 U4990 ( .A1(n3974), .A2(n2962), .ZN(n3975) );
  AND2_X1 U4991 ( .A1(n5541), .A2(n3975), .ZN(n4516) );
  AOI21_X1 U4992 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6334) );
  NOR2_X1 U4993 ( .A1(n6334), .A2(n4840), .ZN(n4844) );
  NAND3_X1 U4994 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n4844), .ZN(n4869) );
  NOR2_X1 U4995 ( .A1(n4869), .A2(n3976), .ZN(n4101) );
  NAND2_X1 U4996 ( .A1(n6332), .A2(n4101), .ZN(n5994) );
  AND2_X1 U4997 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5966) );
  NAND2_X1 U4998 ( .A1(n5782), .A2(n5966), .ZN(n5771) );
  NOR2_X1 U4999 ( .A1(n5771), .A2(n4111), .ZN(n4470) );
  INV_X1 U5000 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4286) );
  AND2_X1 U5001 ( .A1(n6284), .A2(REIP_REG_29__SCAN_IN), .ZN(n5691) );
  OR2_X1 U5002 ( .A1(n3987), .A2(EBX_REG_1__SCAN_IN), .ZN(n3983) );
  NAND2_X1 U5003 ( .A1(n4011), .A2(n6339), .ZN(n3981) );
  INV_X1 U5004 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3979) );
  NAND2_X1 U5005 ( .A1(n4557), .A2(n3979), .ZN(n3980) );
  NAND3_X1 U5006 ( .A1(n3981), .A2(n3980), .A3(n5662), .ZN(n3982) );
  NAND2_X1 U5007 ( .A1(n4011), .A2(EBX_REG_0__SCAN_IN), .ZN(n3985) );
  INV_X1 U5008 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5176) );
  NAND2_X1 U5009 ( .A1(n5662), .A2(n5176), .ZN(n3984) );
  NAND2_X1 U5010 ( .A1(n3985), .A2(n3984), .ZN(n4541) );
  XNOR2_X1 U5011 ( .A(n3986), .B(n4541), .ZN(n4555) );
  NAND2_X1 U5012 ( .A1(n4555), .A2(n4557), .ZN(n4556) );
  NAND2_X1 U5013 ( .A1(n4556), .A2(n3986), .ZN(n4584) );
  MUX2_X1 U5014 ( .A(n4076), .B(n4011), .S(EBX_REG_2__SCAN_IN), .Z(n3990) );
  INV_X1 U5015 ( .A(n4011), .ZN(n3988) );
  NAND2_X1 U5016 ( .A1(n3988), .A2(n2962), .ZN(n4063) );
  NAND2_X1 U5017 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n2962), .ZN(n3989)
         );
  AND3_X1 U5018 ( .A1(n3990), .A2(n4063), .A3(n3989), .ZN(n4583) );
  MUX2_X1 U5019 ( .A(n4082), .B(n5662), .S(EBX_REG_3__SCAN_IN), .Z(n3994) );
  OR2_X1 U5020 ( .A1(n4542), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3993)
         );
  NAND2_X1 U5021 ( .A1(n3994), .A2(n3993), .ZN(n4550) );
  OR2_X1 U5022 ( .A1(n4076), .A2(EBX_REG_4__SCAN_IN), .ZN(n3999) );
  NAND2_X1 U5023 ( .A1(n4025), .A2(n3995), .ZN(n3997) );
  INV_X1 U5024 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6130) );
  NAND2_X1 U5025 ( .A1(n4557), .A2(n6130), .ZN(n3996) );
  NAND3_X1 U5026 ( .A1(n3997), .A2(n3996), .A3(n5662), .ZN(n3998) );
  NAND2_X1 U5027 ( .A1(n3999), .A2(n3998), .ZN(n4579) );
  NAND2_X1 U5028 ( .A1(n4580), .A2(n4579), .ZN(n4655) );
  MUX2_X1 U5029 ( .A(n4082), .B(n5662), .S(EBX_REG_5__SCAN_IN), .Z(n4000) );
  OAI21_X1 U5030 ( .B1(n4542), .B2(INSTADDRPOINTER_REG_5__SCAN_IN), .A(n4000), 
        .ZN(n4656) );
  NAND2_X1 U5031 ( .A1(n3475), .A2(n4086), .ZN(n4004) );
  MUX2_X1 U5032 ( .A(n4082), .B(n5662), .S(EBX_REG_7__SCAN_IN), .Z(n4003) );
  OR2_X1 U5033 ( .A1(n4076), .A2(EBX_REG_6__SCAN_IN), .ZN(n4009) );
  NAND2_X1 U5034 ( .A1(n4025), .A2(n4005), .ZN(n4007) );
  INV_X1 U5035 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U5036 ( .A1(n4557), .A2(n6183), .ZN(n4006) );
  NAND3_X1 U5037 ( .A1(n4007), .A2(n4006), .A3(n5662), .ZN(n4008) );
  NAND2_X1 U5038 ( .A1(n4009), .A2(n4008), .ZN(n4941) );
  NAND2_X1 U5039 ( .A1(n4712), .A2(n4941), .ZN(n4010) );
  OR2_X1 U5040 ( .A1(n4076), .A2(EBX_REG_8__SCAN_IN), .ZN(n4016) );
  NAND2_X1 U5041 ( .A1(n4025), .A2(n4012), .ZN(n4014) );
  INV_X1 U5042 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U5043 ( .A1(n4557), .A2(n5611), .ZN(n4013) );
  NAND3_X1 U5044 ( .A1(n4014), .A2(n4013), .A3(n5662), .ZN(n4015) );
  NAND2_X1 U5045 ( .A1(n4016), .A2(n4015), .ZN(n4759) );
  NAND2_X1 U5046 ( .A1(n5194), .A2(n4086), .ZN(n4018) );
  MUX2_X1 U5047 ( .A(n4082), .B(n5662), .S(EBX_REG_9__SCAN_IN), .Z(n4017) );
  NAND2_X1 U5048 ( .A1(n4880), .A2(n4879), .ZN(n4878) );
  MUX2_X1 U5049 ( .A(n4076), .B(n4025), .S(EBX_REG_10__SCAN_IN), .Z(n4020) );
  NAND2_X1 U5050 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n2962), .ZN(n4019) );
  OR2_X1 U5051 ( .A1(n4082), .A2(EBX_REG_11__SCAN_IN), .ZN(n4023) );
  NAND2_X1 U5052 ( .A1(n5662), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4021) );
  OAI211_X1 U5053 ( .C1(n2962), .C2(EBX_REG_11__SCAN_IN), .A(n4025), .B(n4021), 
        .ZN(n4022) );
  NAND2_X1 U5054 ( .A1(n4023), .A2(n4022), .ZN(n5038) );
  NAND2_X1 U5055 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n2962), .ZN(n4024) );
  AND2_X1 U5056 ( .A1(n4063), .A2(n4024), .ZN(n4027) );
  MUX2_X1 U5057 ( .A(n4076), .B(n4025), .S(EBX_REG_12__SCAN_IN), .Z(n4026) );
  NAND2_X1 U5058 ( .A1(n4027), .A2(n4026), .ZN(n5327) );
  OR2_X1 U5059 ( .A1(n4082), .A2(EBX_REG_13__SCAN_IN), .ZN(n4030) );
  NAND2_X1 U5060 ( .A1(n5662), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4028) );
  OAI211_X1 U5061 ( .C1(EBX_REG_13__SCAN_IN), .C2(n2962), .A(n4025), .B(n4028), 
        .ZN(n4029) );
  AND2_X1 U5062 ( .A1(n4030), .A2(n4029), .ZN(n5289) );
  AND2_X2 U5063 ( .A1(n5326), .A2(n4031), .ZN(n5433) );
  NAND2_X1 U5064 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n2962), .ZN(n4032) );
  AND2_X1 U5065 ( .A1(n4063), .A2(n4032), .ZN(n4034) );
  MUX2_X1 U5066 ( .A(n4076), .B(n4025), .S(EBX_REG_14__SCAN_IN), .Z(n4033) );
  NAND2_X1 U5067 ( .A1(n4034), .A2(n4033), .ZN(n5432) );
  NAND2_X1 U5068 ( .A1(n5433), .A2(n5432), .ZN(n5442) );
  OR2_X1 U5069 ( .A1(n4082), .A2(EBX_REG_15__SCAN_IN), .ZN(n4037) );
  NAND2_X1 U5070 ( .A1(n5662), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4035) );
  OAI211_X1 U5071 ( .C1(n2962), .C2(EBX_REG_15__SCAN_IN), .A(n4025), .B(n4035), 
        .ZN(n4036) );
  NAND2_X1 U5072 ( .A1(n4037), .A2(n4036), .ZN(n5443) );
  NOR2_X2 U5073 ( .A1(n5442), .A2(n5443), .ZN(n5440) );
  MUX2_X1 U5074 ( .A(n4076), .B(n4025), .S(EBX_REG_16__SCAN_IN), .Z(n4039) );
  NAND2_X1 U5075 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n2962), .ZN(n4038) );
  OR2_X1 U5076 ( .A1(n4082), .A2(EBX_REG_17__SCAN_IN), .ZN(n4043) );
  NAND2_X1 U5077 ( .A1(n5662), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4041) );
  OAI211_X1 U5078 ( .C1(n2962), .C2(EBX_REG_17__SCAN_IN), .A(n4025), .B(n4041), 
        .ZN(n4042) );
  INV_X1 U5079 ( .A(n4076), .ZN(n4070) );
  INV_X1 U5080 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5528) );
  NAND2_X1 U5081 ( .A1(n4070), .A2(n5528), .ZN(n4046) );
  INV_X1 U5082 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5836) );
  NAND2_X1 U5083 ( .A1(n4025), .A2(n5836), .ZN(n4044) );
  OAI211_X1 U5084 ( .C1(n2962), .C2(EBX_REG_19__SCAN_IN), .A(n4044), .B(n5662), 
        .ZN(n4045) );
  NOR2_X2 U5085 ( .A1(n5525), .A2(n5523), .ZN(n5522) );
  NAND2_X1 U5086 ( .A1(n4542), .A2(EBX_REG_18__SCAN_IN), .ZN(n4048) );
  NAND2_X1 U5087 ( .A1(n2962), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4047) );
  NAND2_X1 U5088 ( .A1(n4048), .A2(n4047), .ZN(n5516) );
  INV_X1 U5089 ( .A(n5516), .ZN(n5663) );
  OR2_X1 U5090 ( .A1(n4542), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4050)
         );
  INV_X1 U5091 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5912) );
  NAND2_X1 U5092 ( .A1(n4557), .A2(n5912), .ZN(n4049) );
  AND2_X1 U5093 ( .A1(n4050), .A2(n4049), .ZN(n4051) );
  INV_X1 U5094 ( .A(n4051), .ZN(n5664) );
  NAND2_X1 U5095 ( .A1(n5663), .A2(n5664), .ZN(n4053) );
  NAND2_X1 U5096 ( .A1(n4051), .A2(n5516), .ZN(n4052) );
  MUX2_X1 U5097 ( .A(n4053), .B(n4052), .S(n5662), .Z(n4054) );
  NAND2_X1 U5098 ( .A1(n5522), .A2(n4055), .ZN(n5654) );
  INV_X1 U5099 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U5100 ( .A1(n4070), .A2(n5903), .ZN(n4058) );
  NAND2_X1 U5101 ( .A1(n4025), .A2(n5812), .ZN(n4056) );
  OAI211_X1 U5102 ( .C1(n2962), .C2(EBX_REG_21__SCAN_IN), .A(n4056), .B(n5662), 
        .ZN(n4057) );
  AND2_X1 U5103 ( .A1(n4058), .A2(n4057), .ZN(n5653) );
  NOR2_X2 U5104 ( .A1(n5654), .A2(n5653), .ZN(n5655) );
  OR2_X1 U5105 ( .A1(n4082), .A2(EBX_REG_22__SCAN_IN), .ZN(n4061) );
  NAND2_X1 U5106 ( .A1(n5662), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4059) );
  OAI211_X1 U5107 ( .C1(n2962), .C2(EBX_REG_22__SCAN_IN), .A(n4025), .B(n4059), 
        .ZN(n4060) );
  AND2_X1 U5108 ( .A1(n4061), .A2(n4060), .ZN(n5603) );
  AND2_X2 U5109 ( .A1(n5655), .A2(n5603), .ZN(n5647) );
  NAND2_X1 U5110 ( .A1(n2962), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4062) );
  AND2_X1 U5111 ( .A1(n4063), .A2(n4062), .ZN(n4065) );
  MUX2_X1 U5112 ( .A(n4076), .B(n4025), .S(EBX_REG_23__SCAN_IN), .Z(n4064) );
  NAND2_X1 U5113 ( .A1(n4065), .A2(n4064), .ZN(n5646) );
  NAND2_X1 U5114 ( .A1(n5647), .A2(n5646), .ZN(n5637) );
  OR2_X1 U5115 ( .A1(n4082), .A2(EBX_REG_24__SCAN_IN), .ZN(n4068) );
  NAND2_X1 U5116 ( .A1(n5662), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4066) );
  OAI211_X1 U5117 ( .C1(EBX_REG_24__SCAN_IN), .C2(n2962), .A(n4025), .B(n4066), 
        .ZN(n4067) );
  NAND2_X1 U5118 ( .A1(n4068), .A2(n4067), .ZN(n5638) );
  INV_X1 U5119 ( .A(n4069), .ZN(n5640) );
  INV_X1 U5120 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U5121 ( .A1(n4070), .A2(n5549), .ZN(n4073) );
  NAND2_X1 U5122 ( .A1(n4025), .A2(n5967), .ZN(n4071) );
  OAI211_X1 U5123 ( .C1(n2962), .C2(EBX_REG_25__SCAN_IN), .A(n4071), .B(n5662), 
        .ZN(n4072) );
  AND2_X1 U5124 ( .A1(n4073), .A2(n4072), .ZN(n4504) );
  MUX2_X1 U5125 ( .A(n4082), .B(n5662), .S(EBX_REG_26__SCAN_IN), .Z(n4075) );
  OR2_X1 U5126 ( .A1(n4542), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4074)
         );
  AND2_X1 U5127 ( .A1(n4075), .A2(n4074), .ZN(n5591) );
  AND2_X2 U5128 ( .A1(n5590), .A2(n5591), .ZN(n5630) );
  OR2_X1 U5129 ( .A1(n4076), .A2(EBX_REG_27__SCAN_IN), .ZN(n4081) );
  INV_X1 U5130 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4077) );
  NAND2_X1 U5131 ( .A1(n4025), .A2(n4077), .ZN(n4079) );
  INV_X1 U5132 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U5133 ( .A1(n4557), .A2(n5632), .ZN(n4078) );
  NAND3_X1 U5134 ( .A1(n4079), .A2(n4078), .A3(n5662), .ZN(n4080) );
  NAND2_X1 U5135 ( .A1(n4081), .A2(n4080), .ZN(n5629) );
  NAND2_X1 U5136 ( .A1(n5630), .A2(n5629), .ZN(n4489) );
  MUX2_X1 U5137 ( .A(n4082), .B(n5662), .S(EBX_REG_28__SCAN_IN), .Z(n4084) );
  OR2_X1 U5138 ( .A1(n4542), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4083)
         );
  NAND2_X1 U5139 ( .A1(n4084), .A2(n4083), .ZN(n4490) );
  OR2_X2 U5140 ( .A1(n4489), .A2(n4490), .ZN(n4492) );
  NOR2_X1 U5141 ( .A1(n2962), .A2(EBX_REG_29__SCAN_IN), .ZN(n4085) );
  AOI21_X1 U5142 ( .B1(n4086), .B2(n4286), .A(n4085), .ZN(n4312) );
  OR2_X1 U5143 ( .A1(n4312), .A2(n5515), .ZN(n4250) );
  NAND2_X1 U5144 ( .A1(n5515), .A2(EBX_REG_29__SCAN_IN), .ZN(n4087) );
  NAND2_X1 U5145 ( .A1(n4250), .A2(n4087), .ZN(n4088) );
  OR2_X2 U5146 ( .A1(n4492), .A2(n4088), .ZN(n4253) );
  NAND2_X1 U5147 ( .A1(n4492), .A2(n4088), .ZN(n4089) );
  NAND2_X1 U5148 ( .A1(n4253), .A2(n4089), .ZN(n5622) );
  NAND2_X1 U5149 ( .A1(n3955), .A2(n2968), .ZN(n4090) );
  NAND2_X1 U5150 ( .A1(n4599), .A2(n6731), .ZN(n6600) );
  NAND2_X1 U5151 ( .A1(n4090), .A2(n6600), .ZN(n4091) );
  NOR2_X1 U5152 ( .A1(n5622), .A2(n5996), .ZN(n4092) );
  AOI211_X1 U5153 ( .C1(n4470), .C2(n4286), .A(n5691), .B(n4092), .ZN(n4113)
         );
  NAND2_X1 U5154 ( .A1(n5816), .A2(n5995), .ZN(n5462) );
  INV_X1 U5155 ( .A(n5826), .ZN(n4094) );
  NOR2_X1 U5156 ( .A1(n5824), .A2(n4094), .ZN(n5813) );
  INV_X1 U5157 ( .A(n4095), .ZN(n4096) );
  NAND2_X1 U5158 ( .A1(n5813), .A2(n4096), .ZN(n5799) );
  INV_X1 U5159 ( .A(n5995), .ZN(n4098) );
  INV_X1 U5160 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6331) );
  OR2_X1 U5161 ( .A1(n4097), .A2(n6284), .ZN(n4539) );
  INV_X1 U5162 ( .A(n4539), .ZN(n4619) );
  AOI21_X1 U5163 ( .B1(n4098), .B2(n6331), .A(n4619), .ZN(n4865) );
  OAI21_X1 U5164 ( .B1(n4867), .B2(n4099), .A(n4865), .ZN(n5325) );
  INV_X1 U5165 ( .A(n5325), .ZN(n4100) );
  OAI21_X1 U5166 ( .B1(n5816), .B2(n4101), .A(n4100), .ZN(n5976) );
  INV_X1 U5167 ( .A(n4102), .ZN(n4103) );
  AND2_X1 U5168 ( .A1(n5977), .A2(n4103), .ZN(n4104) );
  OR2_X1 U5169 ( .A1(n5976), .A2(n4104), .ZN(n5857) );
  NAND2_X1 U5170 ( .A1(n5826), .A2(n4105), .ZN(n4106) );
  AND2_X1 U5171 ( .A1(n5977), .A2(n4106), .ZN(n4107) );
  NOR2_X1 U5172 ( .A1(n5857), .A2(n4107), .ZN(n5809) );
  NAND2_X1 U5173 ( .A1(n6338), .A2(n5816), .ZN(n5324) );
  INV_X1 U5174 ( .A(n4108), .ZN(n4109) );
  NAND2_X1 U5175 ( .A1(n5324), .A2(n4109), .ZN(n4110) );
  OAI21_X1 U5176 ( .B1(n5030), .B2(n5966), .A(n5975), .ZN(n5775) );
  AOI21_X1 U5177 ( .B1(n4111), .B2(n5977), .A(n5775), .ZN(n4295) );
  OR2_X1 U5178 ( .A1(n4295), .A2(n4286), .ZN(n4112) );
  OAI21_X1 U5179 ( .B1(n5697), .B2(n5997), .A(n4114), .ZN(U2989) );
  AOI22_X1 U5180 ( .A1(n4133), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4664), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4118) );
  AOI22_X1 U5181 ( .A1(n4213), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4117) );
  AOI22_X1 U5182 ( .A1(n4224), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3235), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4116) );
  AOI22_X1 U5183 ( .A1(n4225), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4115) );
  NAND4_X1 U5184 ( .A1(n4118), .A2(n4117), .A3(n4116), .A4(n4115), .ZN(n4124)
         );
  AOI22_X1 U5185 ( .A1(n4141), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4122) );
  AOI22_X1 U5186 ( .A1(n4215), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4121) );
  AOI22_X1 U5187 ( .A1(n3661), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4120) );
  AOI22_X1 U5188 ( .A1(n4132), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4119) );
  NAND4_X1 U5189 ( .A1(n4122), .A2(n4121), .A3(n4120), .A4(n4119), .ZN(n4123)
         );
  OR2_X1 U5190 ( .A1(n4124), .A2(n4123), .ZN(n4165) );
  NAND2_X1 U5191 ( .A1(n4126), .A2(n4125), .ZN(n4173) );
  AOI22_X1 U5192 ( .A1(n4215), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4213), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U5193 ( .A1(n3661), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4130) );
  AOI22_X1 U5194 ( .A1(n3250), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4129) );
  AOI22_X1 U5195 ( .A1(n4214), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3248), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4128) );
  NAND4_X1 U5196 ( .A1(n4131), .A2(n4130), .A3(n4129), .A4(n4128), .ZN(n4139)
         );
  AOI22_X1 U5197 ( .A1(n4141), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4225), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4137) );
  AOI22_X1 U5198 ( .A1(n4664), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4132), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4136) );
  AOI22_X1 U5199 ( .A1(n4133), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4135) );
  AOI22_X1 U5200 ( .A1(n3229), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3230), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4134) );
  NAND4_X1 U5201 ( .A1(n4137), .A2(n4136), .A3(n4135), .A4(n4134), .ZN(n4138)
         );
  OR2_X1 U5202 ( .A1(n4139), .A2(n4138), .ZN(n4172) );
  INV_X1 U5203 ( .A(n4172), .ZN(n4140) );
  NOR2_X1 U5204 ( .A1(n4173), .A2(n4140), .ZN(n4164) );
  AND2_X1 U5205 ( .A1(n4165), .A2(n4164), .ZN(n4203) );
  AOI22_X1 U5206 ( .A1(n4218), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4145) );
  AOI22_X1 U5207 ( .A1(n4141), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4144) );
  AOI22_X1 U5208 ( .A1(n3823), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4143) );
  AOI22_X1 U5209 ( .A1(n4213), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3248), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4142) );
  NAND4_X1 U5210 ( .A1(n4145), .A2(n4144), .A3(n4143), .A4(n4142), .ZN(n4151)
         );
  AOI22_X1 U5211 ( .A1(n4133), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4664), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U5212 ( .A1(n4215), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U5213 ( .A1(n4225), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4147) );
  AOI22_X1 U5214 ( .A1(n4132), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4146) );
  NAND4_X1 U5215 ( .A1(n4149), .A2(n4148), .A3(n4147), .A4(n4146), .ZN(n4150)
         );
  OR2_X1 U5216 ( .A1(n4151), .A2(n4150), .ZN(n4202) );
  XNOR2_X1 U5217 ( .A(n4203), .B(n4202), .ZN(n4156) );
  INV_X1 U5218 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4153) );
  NAND2_X1 U5219 ( .A1(n6514), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4152)
         );
  OAI211_X1 U5220 ( .C1(n4304), .C2(n4153), .A(n4248), .B(n4152), .ZN(n4154)
         );
  INV_X1 U5221 ( .A(n4154), .ZN(n4155) );
  OAI21_X1 U5222 ( .B1(n4156), .B2(n4239), .A(n4155), .ZN(n4163) );
  INV_X1 U5223 ( .A(n4158), .ZN(n4160) );
  INV_X1 U5224 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4159) );
  NAND2_X1 U5225 ( .A1(n4160), .A2(n4159), .ZN(n4161) );
  NAND2_X1 U5226 ( .A1(n4211), .A2(n4161), .ZN(n5705) );
  OR2_X1 U5227 ( .A1(n5705), .A2(n4248), .ZN(n4162) );
  NAND2_X1 U5228 ( .A1(n4163), .A2(n4162), .ZN(n4478) );
  INV_X1 U5229 ( .A(n4478), .ZN(n4189) );
  XOR2_X1 U5230 ( .A(n4165), .B(n4164), .Z(n4168) );
  NAND2_X1 U5231 ( .A1(n6514), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4166)
         );
  OAI211_X1 U5232 ( .C1(n4304), .C2(n4647), .A(n4248), .B(n4166), .ZN(n4167)
         );
  AOI21_X1 U5233 ( .B1(n4168), .B2(n4207), .A(n4167), .ZN(n4169) );
  INV_X1 U5234 ( .A(n4169), .ZN(n4171) );
  INV_X1 U5235 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5713) );
  XNOR2_X1 U5236 ( .A(n4178), .B(n5713), .ZN(n5871) );
  NAND2_X1 U5237 ( .A1(n5871), .A2(n4236), .ZN(n4170) );
  NAND2_X1 U5238 ( .A1(n4171), .A2(n4170), .ZN(n5628) );
  INV_X1 U5239 ( .A(n5628), .ZN(n4188) );
  XNOR2_X1 U5240 ( .A(n4173), .B(n4172), .ZN(n4174) );
  NAND2_X1 U5241 ( .A1(n4174), .A2(n4207), .ZN(n4186) );
  INV_X1 U5242 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4176) );
  NAND2_X1 U5243 ( .A1(n6514), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4175)
         );
  OAI211_X1 U5244 ( .C1(n4304), .C2(n4176), .A(n4248), .B(n4175), .ZN(n4177)
         );
  INV_X1 U5245 ( .A(n4177), .ZN(n4185) );
  INV_X1 U5246 ( .A(n4178), .ZN(n4183) );
  INV_X1 U5247 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4181) );
  INV_X1 U5248 ( .A(n4179), .ZN(n4180) );
  NAND2_X1 U5249 ( .A1(n4181), .A2(n4180), .ZN(n4182) );
  NAND2_X1 U5250 ( .A1(n4183), .A2(n4182), .ZN(n5588) );
  NOR2_X1 U5251 ( .A1(n5588), .A2(n4248), .ZN(n4184) );
  AOI21_X1 U5252 ( .B1(n4186), .B2(n4185), .A(n4184), .ZN(n4437) );
  AND2_X1 U5253 ( .A1(n4437), .A2(n4187), .ZN(n4436) );
  XNOR2_X1 U5254 ( .A(n4211), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5580)
         );
  AOI22_X1 U5255 ( .A1(n4218), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4224), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4194) );
  AOI22_X1 U5256 ( .A1(n4141), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4193) );
  AOI22_X1 U5257 ( .A1(n3823), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4192) );
  AOI22_X1 U5258 ( .A1(n4213), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3248), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4191) );
  NAND4_X1 U5259 ( .A1(n4194), .A2(n4193), .A3(n4192), .A4(n4191), .ZN(n4201)
         );
  AOI22_X1 U5260 ( .A1(n4195), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4664), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4199) );
  AOI22_X1 U5261 ( .A1(n4215), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4198) );
  AOI22_X1 U5262 ( .A1(n4225), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4197) );
  AOI22_X1 U5263 ( .A1(n3264), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4196) );
  NAND4_X1 U5264 ( .A1(n4199), .A2(n4198), .A3(n4197), .A4(n4196), .ZN(n4200)
         );
  NOR2_X1 U5265 ( .A1(n4201), .A2(n4200), .ZN(n4233) );
  NAND2_X1 U5266 ( .A1(n4203), .A2(n4202), .ZN(n4232) );
  XOR2_X1 U5267 ( .A(n4233), .B(n4232), .Z(n4208) );
  INV_X1 U5268 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4205) );
  NAND2_X1 U5269 ( .A1(n4243), .A2(EAX_REG_29__SCAN_IN), .ZN(n4204) );
  OAI211_X1 U5270 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n4205), .A(n4204), .B(
        n4248), .ZN(n4206) );
  AOI21_X1 U5271 ( .B1(n4208), .B2(n4207), .A(n4206), .ZN(n4209) );
  AOI21_X1 U5272 ( .B1(n4236), .B2(n5580), .A(n4209), .ZN(n5578) );
  INV_X1 U5273 ( .A(n4211), .ZN(n4212) );
  NAND2_X1 U5274 ( .A1(n4212), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4246)
         );
  INV_X1 U5275 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4245) );
  XNOR2_X1 U5276 ( .A(n4246), .B(n4245), .ZN(n5685) );
  AOI22_X1 U5277 ( .A1(n4213), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4141), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4222) );
  AOI22_X1 U5278 ( .A1(n4215), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4221) );
  AOI22_X1 U5279 ( .A1(n3823), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4220) );
  AOI22_X1 U5280 ( .A1(n4218), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3248), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4219) );
  NAND4_X1 U5281 ( .A1(n4222), .A2(n4221), .A3(n4220), .A4(n4219), .ZN(n4231)
         );
  AOI22_X1 U5282 ( .A1(n4133), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4664), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4229) );
  AOI22_X1 U5283 ( .A1(n4224), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4228) );
  AOI22_X1 U5284 ( .A1(n4225), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3340), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4227) );
  AOI22_X1 U5285 ( .A1(n3264), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3230), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4226) );
  NAND4_X1 U5286 ( .A1(n4229), .A2(n4228), .A3(n4227), .A4(n4226), .ZN(n4230)
         );
  NOR2_X1 U5287 ( .A1(n4231), .A2(n4230), .ZN(n4235) );
  NOR2_X1 U5288 ( .A1(n4233), .A2(n4232), .ZN(n4234) );
  XOR2_X1 U5289 ( .A(n4235), .B(n4234), .Z(n4240) );
  AOI21_X1 U5290 ( .B1(PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6514), .A(n4236), 
        .ZN(n4238) );
  NAND2_X1 U5291 ( .A1(n4243), .A2(EAX_REG_30__SCAN_IN), .ZN(n4237) );
  OAI211_X1 U5292 ( .C1(n4240), .C2(n4239), .A(n4238), .B(n4237), .ZN(n4241)
         );
  OAI21_X1 U5293 ( .B1(n4248), .B2(n5685), .A(n4241), .ZN(n4302) );
  AOI22_X1 U5294 ( .A1(n4243), .A2(EAX_REG_31__SCAN_IN), .B1(n4242), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4244) );
  XNOR2_X1 U5295 ( .A(n4301), .B(n4244), .ZN(n5670) );
  INV_X1 U5296 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4356) );
  XNOR2_X1 U5297 ( .A(n4247), .B(n4356), .ZN(n5556) );
  NOR3_X1 U5298 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6614), .A3(n4248), .ZN(
        n6616) );
  INV_X1 U5299 ( .A(n6616), .ZN(n4486) );
  NAND2_X1 U5300 ( .A1(n5670), .A2(n5880), .ZN(n4285) );
  AND2_X1 U5301 ( .A1(n2962), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4249)
         );
  AOI21_X1 U5302 ( .B1(n4542), .B2(EBX_REG_30__SCAN_IN), .A(n4249), .ZN(n4314)
         );
  INV_X1 U5303 ( .A(n4314), .ZN(n4252) );
  NAND2_X1 U5304 ( .A1(n4492), .A2(n5662), .ZN(n4311) );
  OAI22_X1 U5305 ( .A1(n4542), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n2962), .ZN(n4254) );
  INV_X1 U5306 ( .A(READY_N), .ZN(n6729) );
  NAND2_X1 U5307 ( .A1(n6729), .A2(n6015), .ZN(n4482) );
  INV_X1 U5308 ( .A(n4482), .ZN(n4262) );
  NOR2_X1 U5309 ( .A1(n4256), .A2(n4517), .ZN(n4511) );
  NAND2_X1 U5310 ( .A1(n4511), .A2(n6612), .ZN(n4528) );
  INV_X1 U5311 ( .A(n6727), .ZN(n5173) );
  NAND2_X1 U5312 ( .A1(EBX_REG_31__SCAN_IN), .A2(n6727), .ZN(n4265) );
  INV_X1 U5313 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6697) );
  INV_X1 U5314 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6693) );
  INV_X1 U5315 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6691) );
  NOR2_X1 U5316 ( .A1(n4482), .A2(n5173), .ZN(n4257) );
  AND2_X1 U5317 ( .A1(n4628), .A2(n4257), .ZN(n4258) );
  NAND2_X2 U5318 ( .A1(n4259), .A2(n4258), .ZN(n6131) );
  INV_X1 U5319 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6670) );
  NAND3_X1 U5320 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6086) );
  INV_X1 U5321 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6654) );
  INV_X1 U5322 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6655) );
  NOR2_X1 U5323 ( .A1(n6654), .A2(n6655), .ZN(n6089) );
  INV_X1 U5324 ( .A(n6089), .ZN(n4260) );
  NAND3_X1 U5325 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_6__SCAN_IN), .ZN(n5279) );
  NOR3_X1 U5326 ( .A1(n6086), .A2(n4260), .A3(n5279), .ZN(n5186) );
  AND4_X1 U5327 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .A4(n5186), .ZN(n5280) );
  NAND2_X1 U5328 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5280), .ZN(n6069) );
  NOR2_X1 U5329 ( .A1(n6670), .A2(n6069), .ZN(n6056) );
  NAND2_X1 U5330 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6056), .ZN(n4268) );
  NOR2_X2 U5331 ( .A1(n6131), .A2(n4268), .ZN(n6045) );
  NAND2_X1 U5332 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .ZN(
        n4270) );
  INV_X1 U5333 ( .A(REIP_REG_17__SCAN_IN), .ZN(n5489) );
  NAND3_X1 U5334 ( .A1(n6034), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n5918) );
  INV_X1 U5335 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6683) );
  NOR2_X2 U5336 ( .A1(n5918), .A2(n6683), .ZN(n5892) );
  NOR2_X1 U5337 ( .A1(n6691), .A2(n4266), .ZN(n4500) );
  NAND2_X1 U5338 ( .A1(REIP_REG_25__SCAN_IN), .A2(n4500), .ZN(n5587) );
  NAND2_X1 U5339 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5876), .ZN(n4493) );
  INV_X1 U5340 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6705) );
  NAND2_X1 U5341 ( .A1(n6638), .A2(n4262), .ZN(n6599) );
  NAND2_X1 U5342 ( .A1(n6731), .A2(n6599), .ZN(n4484) );
  NOR2_X1 U5343 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6735) );
  NAND3_X1 U5344 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), 
        .A3(n6735), .ZN(n6608) );
  NAND3_X1 U5345 ( .A1(n6309), .A2(n6608), .A3(n4486), .ZN(n4263) );
  NOR2_X2 U5346 ( .A1(n6716), .A2(n4267), .ZN(n6158) );
  OAI22_X1 U5347 ( .A1(n4484), .A2(n4265), .B1(n4356), .B2(n6144), .ZN(n4282)
         );
  NAND2_X1 U5348 ( .A1(REIP_REG_30__SCAN_IN), .A2(REIP_REG_29__SCAN_IN), .ZN(
        n5569) );
  INV_X1 U5349 ( .A(n5569), .ZN(n4279) );
  NOR2_X1 U5350 ( .A1(REIP_REG_24__SCAN_IN), .A2(n4266), .ZN(n5886) );
  NOR2_X1 U5351 ( .A1(n4268), .A2(n4267), .ZN(n6054) );
  INV_X1 U5352 ( .A(n6054), .ZN(n4269) );
  NOR2_X1 U5353 ( .A1(n4270), .A2(n4269), .ZN(n4271) );
  AND2_X1 U5354 ( .A1(n4264), .A2(n6131), .ZN(n6055) );
  AOI21_X1 U5355 ( .B1(REIP_REG_17__SCAN_IN), .B2(n4271), .A(n6055), .ZN(n6035) );
  NAND2_X1 U5356 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5924) );
  NOR2_X1 U5357 ( .A1(n5924), .A2(n6683), .ZN(n4272) );
  NOR2_X1 U5358 ( .A1(n6055), .A2(n4272), .ZN(n4273) );
  NOR2_X1 U5359 ( .A1(n6035), .A2(n4273), .ZN(n5919) );
  OR2_X1 U5360 ( .A1(n6131), .A2(n2986), .ZN(n4274) );
  NAND2_X1 U5361 ( .A1(n5919), .A2(n4274), .ZN(n5898) );
  AND2_X1 U5362 ( .A1(REIP_REG_25__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .ZN(
        n4275) );
  NOR2_X1 U5363 ( .A1(n6131), .A2(n4275), .ZN(n4276) );
  NOR2_X1 U5364 ( .A1(n4496), .A2(n4276), .ZN(n5874) );
  INV_X1 U5365 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6695) );
  NOR2_X1 U5366 ( .A1(n6697), .A2(n6695), .ZN(n4277) );
  OR2_X1 U5367 ( .A1(n6131), .A2(n4277), .ZN(n4278) );
  OAI21_X1 U5368 ( .B1(n4279), .B2(n6131), .A(n5582), .ZN(n4280) );
  NOR3_X1 U5369 ( .A1(n2984), .A2(n4282), .A3(n4281), .ZN(n4283) );
  NAND2_X1 U5370 ( .A1(n4285), .A2(n2980), .ZN(U2796) );
  NAND2_X1 U5371 ( .A1(n4463), .A2(n2990), .ZN(n4291) );
  INV_X1 U5372 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4469) );
  NAND3_X1 U5373 ( .A1(n4287), .A2(n4469), .A3(n4286), .ZN(n4288) );
  NAND2_X1 U5374 ( .A1(n4291), .A2(n4290), .ZN(n4292) );
  XNOR2_X1 U5375 ( .A(n4292), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5559)
         );
  INV_X1 U5376 ( .A(n5621), .ZN(n4294) );
  AND2_X1 U5377 ( .A1(n6284), .A2(REIP_REG_31__SCAN_IN), .ZN(n5554) );
  INV_X1 U5378 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4607) );
  AND4_X1 U5379 ( .A1(n4470), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n4607), .ZN(n4293) );
  OAI21_X1 U5380 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5030), .A(n4295), 
        .ZN(n4472) );
  NOR2_X1 U5381 ( .A1(n5030), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4296)
         );
  OAI21_X1 U5382 ( .B1(n4472), .B2(n4296), .A(INSTADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n4297) );
  OAI21_X1 U5383 ( .B1(n5559), .B2(n5997), .A(n4299), .ZN(U2987) );
  NAND2_X1 U5384 ( .A1(n4606), .A2(n4516), .ZN(n4568) );
  AND3_X1 U5385 ( .A1(n4822), .A2(n2973), .A3(n6614), .ZN(n4308) );
  INV_X1 U5386 ( .A(n4303), .ZN(n4307) );
  NOR2_X1 U5387 ( .A1(n4305), .A2(n4304), .ZN(n4306) );
  AND3_X1 U5388 ( .A1(n4308), .A2(n4307), .A3(n4306), .ZN(n4753) );
  NAND2_X1 U5389 ( .A1(n4753), .A2(n4557), .ZN(n4309) );
  OAI21_X1 U5390 ( .B1(n4312), .B2(n4492), .A(n4311), .ZN(n4313) );
  XOR2_X1 U5391 ( .A(n4314), .B(n4313), .Z(n5575) );
  INV_X1 U5392 ( .A(n5533), .ZN(n5669) );
  NAND2_X1 U5393 ( .A1(n5641), .A2(EBX_REG_30__SCAN_IN), .ZN(n4315) );
  INV_X1 U5394 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6246) );
  NOR4_X1 U5395 ( .A1(EAX_REG_30__SCAN_IN), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .A3(n3837), .A4(n6246), .ZN(n4321) );
  NOR4_X1 U5396 ( .A1(EAX_REG_21__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n5974), .A4(n3623), .ZN(n4320)
         );
  NOR4_X1 U5397 ( .A1(EBX_REG_12__SCAN_IN), .A2(EBX_REG_10__SCAN_IN), .A3(
        n4343), .A4(n5836), .ZN(n4319) );
  NOR4_X1 U5398 ( .A1(ADDRESS_REG_13__SCAN_IN), .A2(ADDRESS_REG_4__SCAN_IN), 
        .A3(BE_N_REG_0__SCAN_IN), .A4(n3430), .ZN(n4318) );
  NAND4_X1 U5399 ( .A1(n4321), .A2(n4320), .A3(n4319), .A4(n4318), .ZN(n4326)
         );
  INV_X1 U5400 ( .A(EAX_REG_31__SCAN_IN), .ZN(n4390) );
  NAND4_X1 U5401 ( .A1(ADDRESS_REG_29__SCAN_IN), .A2(ADDRESS_REG_10__SCAN_IN), 
        .A3(ADDRESS_REG_8__SCAN_IN), .A4(n4390), .ZN(n4325) );
  NAND4_X1 U5402 ( .A1(UWORD_REG_1__SCAN_IN), .A2(ADDRESS_REG_2__SCAN_IN), 
        .A3(LWORD_REG_12__SCAN_IN), .A4(ADS_N_REG_SCAN_IN), .ZN(n4324) );
  NOR2_X1 U5403 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(DATAWIDTH_REG_28__SCAN_IN), .ZN(n6020) );
  NOR4_X1 U5404 ( .A1(PHYADDRPOINTER_REG_31__SCAN_IN), .A2(DATAI_21_), .A3(
        DATAI_10_), .A4(DATAI_11_), .ZN(n4322) );
  INV_X1 U5405 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6032) );
  INV_X1 U5406 ( .A(DATAI_3_), .ZN(n6257) );
  NAND4_X1 U5407 ( .A1(n6020), .A2(n4322), .A3(n6032), .A4(n6257), .ZN(n4323)
         );
  NOR4_X1 U5408 ( .A1(n4326), .A2(n4325), .A3(n4324), .A4(n4323), .ZN(n4338)
         );
  NAND4_X1 U5409 ( .A1(DATAO_REG_24__SCAN_IN), .A2(DATAWIDTH_REG_3__SCAN_IN), 
        .A3(ADDRESS_REG_14__SCAN_IN), .A4(DATAWIDTH_REG_5__SCAN_IN), .ZN(n4330) );
  NAND4_X1 U5410 ( .A1(DATAI_15_), .A2(REIP_REG_8__SCAN_IN), .A3(
        DATAO_REG_11__SCAN_IN), .A4(LWORD_REG_5__SCAN_IN), .ZN(n4329) );
  NAND4_X1 U5411 ( .A1(REIP_REG_4__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .A3(
        DATAI_25_), .A4(DATAI_6_), .ZN(n4328) );
  NAND4_X1 U5412 ( .A1(REIP_REG_28__SCAN_IN), .A2(DATAI_28_), .A3(DATAI_26_), 
        .A4(DATAI_30_), .ZN(n4327) );
  NOR4_X1 U5413 ( .A1(n4330), .A2(n4329), .A3(n4328), .A4(n4327), .ZN(n4337)
         );
  INV_X1 U5414 ( .A(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n6358) );
  NOR4_X1 U5415 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(
        INSTQUEUE_REG_14__0__SCAN_IN), .A3(INSTQUEUE_REG_13__0__SCAN_IN), .A4(
        n6358), .ZN(n4336) );
  NAND4_X1 U5416 ( .A1(INSTQUEUE_REG_15__3__SCAN_IN), .A2(
        INSTQUEUE_REG_7__1__SCAN_IN), .A3(INSTQUEUE_REG_15__7__SCAN_IN), .A4(
        n4374), .ZN(n4332) );
  INV_X1 U5417 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n6370) );
  INV_X1 U5418 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4402) );
  NAND3_X1 U5419 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n6370), .A3(n4402), 
        .ZN(n4331) );
  NOR3_X1 U5420 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4332), .A3(n4331), 
        .ZN(n4334) );
  NOR2_X1 U5421 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4333) );
  AND4_X1 U5422 ( .A1(n4334), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .A3(
        INSTQUEUE_REG_15__2__SCAN_IN), .A4(n4333), .ZN(n4335) );
  NAND4_X1 U5423 ( .A1(n4338), .A2(n4337), .A3(n4336), .A4(n4335), .ZN(n4432)
         );
  INV_X1 U5424 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4340) );
  AOI22_X1 U5425 ( .A1(n4340), .A2(keyinput22), .B1(keyinput52), .B2(n6032), 
        .ZN(n4339) );
  OAI221_X1 U5426 ( .B1(n4340), .B2(keyinput22), .C1(n6032), .C2(keyinput52), 
        .A(n4339), .ZN(n4350) );
  INV_X1 U5427 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4342) );
  AOI22_X1 U5428 ( .A1(n4343), .A2(keyinput47), .B1(n4342), .B2(keyinput58), 
        .ZN(n4341) );
  OAI221_X1 U5429 ( .B1(n4343), .B2(keyinput47), .C1(n4342), .C2(keyinput58), 
        .A(n4341), .ZN(n4349) );
  INV_X1 U5430 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6661) );
  AOI22_X1 U5431 ( .A1(n6661), .A2(keyinput2), .B1(n3430), .B2(keyinput16), 
        .ZN(n4344) );
  OAI221_X1 U5432 ( .B1(n6661), .B2(keyinput2), .C1(n3430), .C2(keyinput16), 
        .A(n4344), .ZN(n4348) );
  INV_X1 U5433 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6176) );
  INV_X1 U5434 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n4346) );
  AOI22_X1 U5435 ( .A1(n6176), .A2(keyinput4), .B1(keyinput31), .B2(n4346), 
        .ZN(n4345) );
  OAI221_X1 U5436 ( .B1(n6176), .B2(keyinput4), .C1(n4346), .C2(keyinput31), 
        .A(n4345), .ZN(n4347) );
  NOR4_X1 U5437 ( .A1(n4350), .A2(n4349), .A3(n4348), .A4(n4347), .ZN(n4384)
         );
  INV_X1 U5438 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4352) );
  INV_X1 U5439 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6717) );
  AOI22_X1 U5440 ( .A1(n4352), .A2(keyinput25), .B1(keyinput10), .B2(n6717), 
        .ZN(n4351) );
  OAI221_X1 U5441 ( .B1(n4352), .B2(keyinput25), .C1(n6717), .C2(keyinput10), 
        .A(n4351), .ZN(n4361) );
  INV_X1 U5442 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n4354) );
  AOI22_X1 U5443 ( .A1(n4354), .A2(keyinput51), .B1(n3837), .B2(keyinput0), 
        .ZN(n4353) );
  OAI221_X1 U5444 ( .B1(n4354), .B2(keyinput51), .C1(n3837), .C2(keyinput0), 
        .A(n4353), .ZN(n4360) );
  INV_X1 U5445 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n6200) );
  AOI22_X1 U5446 ( .A1(n4356), .A2(keyinput23), .B1(keyinput26), .B2(n6200), 
        .ZN(n4355) );
  OAI221_X1 U5447 ( .B1(n4356), .B2(keyinput23), .C1(n6200), .C2(keyinput26), 
        .A(n4355), .ZN(n4359) );
  AOI22_X1 U5448 ( .A1(n6246), .A2(keyinput54), .B1(n5974), .B2(keyinput13), 
        .ZN(n4357) );
  OAI221_X1 U5449 ( .B1(n6246), .B2(keyinput54), .C1(n5974), .C2(keyinput13), 
        .A(n4357), .ZN(n4358) );
  NOR4_X1 U5450 ( .A1(n4361), .A2(n4360), .A3(n4359), .A4(n4358), .ZN(n4383)
         );
  INV_X1 U5451 ( .A(DATAI_30_), .ZN(n4953) );
  INV_X1 U5452 ( .A(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6629) );
  AOI22_X1 U5453 ( .A1(n4953), .A2(keyinput60), .B1(n6629), .B2(keyinput8), 
        .ZN(n4362) );
  OAI221_X1 U5454 ( .B1(n4953), .B2(keyinput60), .C1(n6629), .C2(keyinput8), 
        .A(n4362), .ZN(n4370) );
  INV_X1 U5455 ( .A(DATAI_15_), .ZN(n5451) );
  INV_X1 U5456 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6249) );
  AOI22_X1 U5457 ( .A1(n5451), .A2(keyinput33), .B1(n6249), .B2(keyinput30), 
        .ZN(n4363) );
  OAI221_X1 U5458 ( .B1(n5451), .B2(keyinput33), .C1(n6249), .C2(keyinput30), 
        .A(n4363), .ZN(n4369) );
  INV_X1 U5459 ( .A(DATAI_11_), .ZN(n6274) );
  AOI22_X1 U5460 ( .A1(n6274), .A2(keyinput34), .B1(keyinput11), .B2(n6654), 
        .ZN(n4364) );
  OAI221_X1 U5461 ( .B1(n6274), .B2(keyinput34), .C1(n6654), .C2(keyinput11), 
        .A(n4364), .ZN(n4368) );
  INV_X1 U5462 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4366) );
  INV_X1 U5463 ( .A(DATAI_28_), .ZN(n4797) );
  AOI22_X1 U5464 ( .A1(n4366), .A2(keyinput56), .B1(keyinput18), .B2(n4797), 
        .ZN(n4365) );
  OAI221_X1 U5465 ( .B1(n4366), .B2(keyinput56), .C1(n4797), .C2(keyinput18), 
        .A(n4365), .ZN(n4367) );
  NOR4_X1 U5466 ( .A1(n4370), .A2(n4369), .A3(n4368), .A4(n4367), .ZN(n4382)
         );
  INV_X1 U5467 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6006) );
  INV_X1 U5468 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4372) );
  AOI22_X1 U5469 ( .A1(n6006), .A2(keyinput14), .B1(n4372), .B2(keyinput15), 
        .ZN(n4371) );
  OAI221_X1 U5470 ( .B1(n6006), .B2(keyinput14), .C1(n4372), .C2(keyinput15), 
        .A(n4371), .ZN(n4380) );
  AOI22_X1 U5471 ( .A1(n5836), .A2(keyinput53), .B1(n4374), .B2(keyinput41), 
        .ZN(n4373) );
  OAI221_X1 U5472 ( .B1(n5836), .B2(keyinput53), .C1(n4374), .C2(keyinput41), 
        .A(n4373), .ZN(n4379) );
  INV_X1 U5473 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n6651) );
  AOI22_X1 U5474 ( .A1(n3623), .A2(keyinput7), .B1(keyinput39), .B2(n6651), 
        .ZN(n4375) );
  OAI221_X1 U5475 ( .B1(n3623), .B2(keyinput7), .C1(n6651), .C2(keyinput39), 
        .A(n4375), .ZN(n4378) );
  INV_X1 U5476 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n6203) );
  INV_X1 U5477 ( .A(LWORD_REG_12__SCAN_IN), .ZN(n6209) );
  AOI22_X1 U5478 ( .A1(n6203), .A2(keyinput24), .B1(keyinput40), .B2(n6209), 
        .ZN(n4376) );
  OAI221_X1 U5479 ( .B1(n6203), .B2(keyinput24), .C1(n6209), .C2(keyinput40), 
        .A(n4376), .ZN(n4377) );
  NOR4_X1 U5480 ( .A1(n4380), .A2(n4379), .A3(n4378), .A4(n4377), .ZN(n4381)
         );
  NAND4_X1 U5481 ( .A1(n4384), .A2(n4383), .A3(n4382), .A4(n4381), .ZN(n4398)
         );
  INV_X1 U5482 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4386) );
  AOI22_X1 U5483 ( .A1(n4386), .A2(keyinput37), .B1(keyinput45), .B2(n5047), 
        .ZN(n4385) );
  OAI221_X1 U5484 ( .B1(n4386), .B2(keyinput37), .C1(n5047), .C2(keyinput45), 
        .A(n4385), .ZN(n4397) );
  INV_X1 U5485 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n6656) );
  INV_X1 U5486 ( .A(DATAI_21_), .ZN(n4388) );
  AOI22_X1 U5487 ( .A1(n6656), .A2(keyinput17), .B1(keyinput62), .B2(n4388), 
        .ZN(n4387) );
  OAI221_X1 U5488 ( .B1(n6656), .B2(keyinput17), .C1(n4388), .C2(keyinput62), 
        .A(n4387), .ZN(n4396) );
  AOI22_X1 U5489 ( .A1(n4390), .A2(keyinput50), .B1(n4457), .B2(keyinput1), 
        .ZN(n4389) );
  OAI221_X1 U5490 ( .B1(n4390), .B2(keyinput50), .C1(n4457), .C2(keyinput1), 
        .A(n4389), .ZN(n4394) );
  XNOR2_X1 U5491 ( .A(n3099), .B(keyinput3), .ZN(n4393) );
  INV_X1 U5492 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4391) );
  XNOR2_X1 U5493 ( .A(keyinput12), .B(n4391), .ZN(n4392) );
  OR3_X1 U5494 ( .A1(n4394), .A2(n4393), .A3(n4392), .ZN(n4395) );
  NOR4_X1 U5495 ( .A1(n4398), .A2(n4397), .A3(n4396), .A4(n4395), .ZN(n4430)
         );
  INV_X1 U5496 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n6667) );
  INV_X1 U5497 ( .A(DATAI_26_), .ZN(n4808) );
  AOI22_X1 U5498 ( .A1(n6667), .A2(keyinput46), .B1(keyinput48), .B2(n4808), 
        .ZN(n4399) );
  OAI221_X1 U5499 ( .B1(n6667), .B2(keyinput46), .C1(n4808), .C2(keyinput48), 
        .A(n4399), .ZN(n4407) );
  INV_X1 U5500 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n6673) );
  AOI22_X1 U5501 ( .A1(n6673), .A2(keyinput29), .B1(n6358), .B2(keyinput36), 
        .ZN(n4400) );
  OAI221_X1 U5502 ( .B1(n6673), .B2(keyinput29), .C1(n6358), .C2(keyinput36), 
        .A(n4400), .ZN(n4406) );
  INV_X1 U5503 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4963) );
  AOI22_X1 U5504 ( .A1(n4402), .A2(keyinput27), .B1(n4963), .B2(keyinput55), 
        .ZN(n4401) );
  OAI221_X1 U5505 ( .B1(n4402), .B2(keyinput27), .C1(n4963), .C2(keyinput55), 
        .A(n4401), .ZN(n4405) );
  INV_X1 U5506 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6627) );
  INV_X1 U5507 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6707) );
  AOI22_X1 U5508 ( .A1(n6627), .A2(keyinput5), .B1(n6707), .B2(keyinput44), 
        .ZN(n4403) );
  OAI221_X1 U5509 ( .B1(n6627), .B2(keyinput5), .C1(n6707), .C2(keyinput44), 
        .A(n4403), .ZN(n4404) );
  NOR4_X1 U5510 ( .A1(n4407), .A2(n4406), .A3(n4405), .A4(n4404), .ZN(n4429)
         );
  INV_X1 U5511 ( .A(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n6364) );
  INV_X1 U5512 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n6704) );
  AOI22_X1 U5513 ( .A1(n6364), .A2(keyinput32), .B1(keyinput43), .B2(n6704), 
        .ZN(n4408) );
  OAI221_X1 U5514 ( .B1(n6364), .B2(keyinput32), .C1(n6704), .C2(keyinput43), 
        .A(n4408), .ZN(n4415) );
  INV_X1 U5515 ( .A(DATAI_10_), .ZN(n6270) );
  INV_X1 U5516 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6674) );
  AOI22_X1 U5517 ( .A1(n6270), .A2(keyinput38), .B1(keyinput57), .B2(n6674), 
        .ZN(n4409) );
  OAI221_X1 U5518 ( .B1(n6270), .B2(keyinput38), .C1(n6674), .C2(keyinput57), 
        .A(n4409), .ZN(n4414) );
  INV_X1 U5519 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n6663) );
  AOI22_X1 U5520 ( .A1(n6663), .A2(keyinput35), .B1(n6501), .B2(keyinput49), 
        .ZN(n4410) );
  OAI221_X1 U5521 ( .B1(n6663), .B2(keyinput35), .C1(n6501), .C2(keyinput49), 
        .A(n4410), .ZN(n4413) );
  AOI22_X1 U5522 ( .A1(n6257), .A2(keyinput6), .B1(n6697), .B2(keyinput63), 
        .ZN(n4411) );
  OAI221_X1 U5523 ( .B1(n6257), .B2(keyinput6), .C1(n6697), .C2(keyinput63), 
        .A(n4411), .ZN(n4412) );
  NOR4_X1 U5524 ( .A1(n4415), .A2(n4414), .A3(n4413), .A4(n4412), .ZN(n4428)
         );
  INV_X1 U5525 ( .A(DATAWIDTH_REG_28__SCAN_IN), .ZN(n6626) );
  INV_X1 U5526 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4636) );
  AOI22_X1 U5527 ( .A1(n6626), .A2(keyinput9), .B1(n4636), .B2(keyinput20), 
        .ZN(n4416) );
  OAI221_X1 U5528 ( .B1(n6626), .B2(keyinput9), .C1(n4636), .C2(keyinput20), 
        .A(n4416), .ZN(n4426) );
  INV_X1 U5529 ( .A(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4418) );
  AOI22_X1 U5530 ( .A1(n4418), .A2(keyinput19), .B1(n6370), .B2(keyinput61), 
        .ZN(n4417) );
  OAI221_X1 U5531 ( .B1(n4418), .B2(keyinput19), .C1(n6370), .C2(keyinput61), 
        .A(n4417), .ZN(n4425) );
  INV_X1 U5532 ( .A(DATAI_25_), .ZN(n4803) );
  INV_X1 U5533 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4420) );
  AOI22_X1 U5534 ( .A1(n4803), .A2(keyinput21), .B1(n4420), .B2(keyinput42), 
        .ZN(n4419) );
  OAI221_X1 U5535 ( .B1(n4803), .B2(keyinput21), .C1(n4420), .C2(keyinput42), 
        .A(n4419), .ZN(n4424) );
  INV_X1 U5536 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6628) );
  AOI22_X1 U5537 ( .A1(n6628), .A2(keyinput28), .B1(n4422), .B2(keyinput59), 
        .ZN(n4421) );
  OAI221_X1 U5538 ( .B1(n6628), .B2(keyinput28), .C1(n4422), .C2(keyinput59), 
        .A(n4421), .ZN(n4423) );
  NOR4_X1 U5539 ( .A1(n4426), .A2(n4425), .A3(n4424), .A4(n4423), .ZN(n4427)
         );
  NAND4_X1 U5540 ( .A1(n4430), .A2(n4429), .A3(n4428), .A4(n4427), .ZN(n4431)
         );
  XOR2_X1 U5541 ( .A(n4432), .B(n4431), .Z(n4433) );
  XNOR2_X1 U5542 ( .A(n4434), .B(n4433), .ZN(U2829) );
  NAND2_X1 U5543 ( .A1(n4480), .A2(n4436), .ZN(n5627) );
  INV_X1 U5544 ( .A(n5635), .ZN(n5936) );
  INV_X1 U5545 ( .A(n6301), .ZN(n6288) );
  INV_X1 U5546 ( .A(n5699), .ZN(n4440) );
  NOR2_X1 U5547 ( .A1(n4441), .A2(n4440), .ZN(n4442) );
  XNOR2_X1 U5548 ( .A(n5698), .B(n4442), .ZN(n5971) );
  AOI22_X1 U5549 ( .A1(n6328), .A2(REIP_REG_26__SCAN_IN), .B1(n6298), .B2(
        PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4443) );
  INV_X1 U5550 ( .A(n4447), .ZN(n5739) );
  OR2_X1 U5551 ( .A1(n5848), .A2(n5836), .ZN(n5741) );
  AND2_X1 U5552 ( .A1(n5848), .A2(n5836), .ZN(n5740) );
  AOI21_X2 U5553 ( .B1(n5739), .B2(n5741), .A(n5740), .ZN(n5821) );
  INV_X1 U5554 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5831) );
  NAND2_X1 U5555 ( .A1(n5848), .A2(n5831), .ZN(n4449) );
  NOR2_X1 U5556 ( .A1(n5848), .A2(n5831), .ZN(n4448) );
  AOI21_X2 U5557 ( .B1(n5821), .B2(n4449), .A(n4448), .ZN(n5731) );
  XNOR2_X1 U5558 ( .A(n5848), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5733)
         );
  NAND2_X2 U5559 ( .A1(n5731), .A2(n5733), .ZN(n5732) );
  INV_X1 U5560 ( .A(n5732), .ZN(n4450) );
  NOR2_X1 U5561 ( .A1(n5848), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5724)
         );
  NAND2_X1 U5562 ( .A1(n4450), .A2(n5724), .ZN(n5717) );
  OR2_X1 U5563 ( .A1(n4451), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4452)
         );
  NAND2_X1 U5564 ( .A1(n5732), .A2(n4452), .ZN(n5726) );
  NAND3_X1 U5565 ( .A1(n5848), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4453) );
  OAI22_X2 U5566 ( .A1(n5717), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5726), .B2(n4453), .ZN(n4454) );
  XNOR2_X1 U5567 ( .A(n4454), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5790)
         );
  XOR2_X1 U5568 ( .A(n4456), .B(n4455), .Z(n5939) );
  AND2_X1 U5569 ( .A1(n6284), .A2(REIP_REG_24__SCAN_IN), .ZN(n5788) );
  INV_X1 U5570 ( .A(n6298), .ZN(n5746) );
  NOR2_X1 U5571 ( .A1(n5746), .A2(n4457), .ZN(n4458) );
  AOI211_X1 U5572 ( .C1(n5961), .C2(n5884), .A(n5788), .B(n4458), .ZN(n4459)
         );
  OAI21_X1 U5573 ( .B1(n5790), .B2(n6016), .A(n4462), .ZN(U2962) );
  NAND2_X1 U5574 ( .A1(n4463), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4467) );
  INV_X1 U5575 ( .A(n4464), .ZN(n4465) );
  NAND2_X1 U5576 ( .A1(n4465), .A2(n4286), .ZN(n4466) );
  NAND2_X1 U5577 ( .A1(n4467), .A2(n4466), .ZN(n4468) );
  XNOR2_X1 U5578 ( .A(n4468), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5689)
         );
  AND3_X1 U5579 ( .A1(n4470), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n4469), 
        .ZN(n4471) );
  AND2_X1 U5580 ( .A1(n6284), .A2(REIP_REG_30__SCAN_IN), .ZN(n5683) );
  AOI211_X1 U5581 ( .C1(n5575), .C2(n6330), .A(n4471), .B(n5683), .ZN(n4474)
         );
  NAND2_X1 U5582 ( .A1(n4472), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4473) );
  OAI21_X1 U5583 ( .B1(n5689), .B2(n5997), .A(n4475), .ZN(U2988) );
  NAND2_X1 U5584 ( .A1(n4477), .A2(n4476), .ZN(n5625) );
  AND2_X1 U5585 ( .A1(n5625), .A2(n4478), .ZN(n4481) );
  OR2_X2 U5586 ( .A1(n4481), .A2(n5579), .ZN(n5931) );
  INV_X1 U5587 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5620) );
  NAND3_X1 U5588 ( .A1(n4628), .A2(n4482), .A3(n5620), .ZN(n4483) );
  NAND2_X1 U5589 ( .A1(n4484), .A2(n4483), .ZN(n4485) );
  NOR2_X1 U5590 ( .A1(n5705), .A2(n6146), .ZN(n4488) );
  OAI22_X1 U5591 ( .A1(n5582), .A2(n6697), .B1(n4159), .B2(n6144), .ZN(n4487)
         );
  AOI211_X1 U5592 ( .C1(n6161), .C2(EBX_REG_28__SCAN_IN), .A(n4488), .B(n4487), 
        .ZN(n4495) );
  NAND2_X1 U5593 ( .A1(n4489), .A2(n4490), .ZN(n4491) );
  NAND2_X1 U5594 ( .A1(n4492), .A2(n4491), .ZN(n5763) );
  OR2_X1 U5595 ( .A1(n5763), .A2(n6157), .ZN(n4494) );
  INV_X1 U5596 ( .A(n4496), .ZN(n4497) );
  INV_X1 U5597 ( .A(REIP_REG_25__SCAN_IN), .ZN(n4499) );
  OAI22_X1 U5598 ( .A1(n5548), .A2(n6039), .B1(n4497), .B2(n4499), .ZN(n4498)
         );
  AOI22_X1 U5599 ( .A1(n4501), .A2(n6160), .B1(n4500), .B2(n4499), .ZN(n4502)
         );
  OAI21_X1 U5600 ( .B1(n4503), .B2(n6144), .A(n4502), .ZN(n4508) );
  AND2_X1 U5601 ( .A1(n5640), .A2(n4504), .ZN(n4505) );
  OR2_X1 U5602 ( .A1(n4505), .A2(n5590), .ZN(n5780) );
  NAND2_X1 U5603 ( .A1(n4510), .A2(n4509), .ZN(U2802) );
  NOR2_X1 U5604 ( .A1(n4511), .A2(n4518), .ZN(n4512) );
  AOI21_X1 U5605 ( .B1(n4606), .B2(n4513), .A(n4512), .ZN(n6008) );
  OR2_X1 U5606 ( .A1(n6731), .A2(n4514), .ZN(n4531) );
  NAND2_X1 U5607 ( .A1(n4531), .A2(n4559), .ZN(n4515) );
  NAND2_X1 U5608 ( .A1(n4515), .A2(n6729), .ZN(n6732) );
  AND2_X1 U5609 ( .A1(n6008), .A2(n6732), .ZN(n6588) );
  NOR2_X1 U5610 ( .A1(n6588), .A2(n6598), .ZN(n6018) );
  INV_X1 U5611 ( .A(MORE_REG_SCAN_IN), .ZN(n4526) );
  INV_X1 U5612 ( .A(n4516), .ZN(n4666) );
  OR2_X1 U5613 ( .A1(n4606), .A2(n4666), .ZN(n4523) );
  NAND2_X1 U5614 ( .A1(n3935), .A2(n4517), .ZN(n4522) );
  INV_X1 U5615 ( .A(n4518), .ZN(n4519) );
  NAND3_X1 U5616 ( .A1(n4519), .A2(n4749), .A3(n6590), .ZN(n4520) );
  NAND2_X1 U5617 ( .A1(n4606), .A2(n4520), .ZN(n4521) );
  AND3_X1 U5618 ( .A1(n4523), .A2(n4522), .A3(n4521), .ZN(n6591) );
  INV_X1 U5619 ( .A(n6591), .ZN(n4524) );
  NAND2_X1 U5620 ( .A1(n6018), .A2(n4524), .ZN(n4525) );
  OAI21_X1 U5621 ( .B1(n6018), .B2(n4526), .A(n4525), .ZN(U3471) );
  INV_X1 U5622 ( .A(n4527), .ZN(n4532) );
  AOI211_X1 U5623 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4528), .A(n6007), .B(
        n4532), .ZN(n4529) );
  INV_X1 U5624 ( .A(n4529), .ZN(U2788) );
  OAI21_X1 U5625 ( .B1(n6007), .B2(READREQUEST_REG_SCAN_IN), .A(n5173), .ZN(
        n4530) );
  OAI21_X1 U5626 ( .B1(n5173), .B2(n4531), .A(n4530), .ZN(U3474) );
  INV_X1 U5627 ( .A(n6600), .ZN(n4533) );
  INV_X2 U5628 ( .A(n6282), .ZN(n6271) );
  NOR2_X1 U5629 ( .A1(n4534), .A2(READY_N), .ZN(n4535) );
  INV_X1 U5630 ( .A(DATAI_12_), .ZN(n5929) );
  NOR2_X1 U5631 ( .A1(n6273), .A2(n5929), .ZN(n6242) );
  AOI21_X1 U5632 ( .B1(n6271), .B2(EAX_REG_12__SCAN_IN), .A(n6242), .ZN(n4536)
         );
  OAI21_X1 U5633 ( .B1(n4658), .B2(n6209), .A(n4536), .ZN(U2951) );
  OAI21_X1 U5634 ( .B1(n4538), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4537), 
        .ZN(n6293) );
  AOI21_X1 U5635 ( .B1(n5464), .B2(n4539), .A(n6331), .ZN(n4540) );
  AOI21_X1 U5636 ( .B1(n6331), .B2(n5462), .A(n4540), .ZN(n4545) );
  OAI21_X1 U5637 ( .B1(n4542), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4541), 
        .ZN(n5182) );
  INV_X1 U5638 ( .A(n5182), .ZN(n4543) );
  AND2_X1 U5639 ( .A1(n6284), .A2(REIP_REG_0__SCAN_IN), .ZN(n6294) );
  AOI21_X1 U5640 ( .B1(n6330), .B2(n4543), .A(n6294), .ZN(n4544) );
  OAI211_X1 U5641 ( .C1(n5997), .C2(n6293), .A(n4545), .B(n4544), .ZN(U3018)
         );
  NOR2_X1 U5642 ( .A1(n4547), .A2(n4548), .ZN(n4549) );
  OR2_X1 U5643 ( .A1(n4546), .A2(n4549), .ZN(n6137) );
  AOI21_X1 U5644 ( .B1(n4586), .B2(n4550), .A(n4580), .ZN(n6139) );
  AOI22_X1 U5645 ( .A1(n6178), .A2(n6139), .B1(n5641), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4551) );
  OAI21_X1 U5646 ( .B1(n5667), .B2(n6137), .A(n4551), .ZN(U2856) );
  OAI21_X1 U5647 ( .B1(n4552), .B2(n4554), .A(n4553), .ZN(n6167) );
  OAI21_X1 U5648 ( .B1(n4555), .B2(n4557), .A(n4556), .ZN(n4622) );
  AOI22_X1 U5649 ( .A1(n6178), .A2(n4622), .B1(n5641), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4558) );
  OAI21_X1 U5650 ( .B1(n5667), .B2(n6167), .A(n4558), .ZN(U2858) );
  NAND2_X1 U5651 ( .A1(n6615), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6714) );
  INV_X1 U5652 ( .A(n6714), .ZN(n4569) );
  AOI21_X1 U5653 ( .B1(n2962), .B2(n4559), .A(READY_N), .ZN(n4560) );
  OAI21_X1 U5654 ( .B1(n5537), .B2(n4599), .A(n4560), .ZN(n4561) );
  OR2_X1 U5655 ( .A1(n4606), .A2(n4561), .ZN(n4567) );
  OR2_X1 U5656 ( .A1(n4606), .A2(n4749), .ZN(n4566) );
  INV_X1 U5657 ( .A(n4748), .ZN(n4564) );
  OAI21_X1 U5658 ( .B1(n5174), .B2(n3204), .A(n4562), .ZN(n4563) );
  AOI21_X1 U5659 ( .B1(n4564), .B2(n4746), .A(n4563), .ZN(n4565) );
  INV_X1 U5660 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6017) );
  NAND2_X1 U5661 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .ZN(n6619) );
  NOR2_X1 U5662 ( .A1(n6615), .A2(n6619), .ZN(n6625) );
  INV_X1 U5663 ( .A(n6625), .ZN(n6713) );
  OAI22_X1 U5664 ( .A1(n6579), .A2(n6598), .B1(n6017), .B2(n6713), .ZN(n4570)
         );
  NOR2_X1 U5665 ( .A1(n4569), .A2(n4570), .ZN(n5869) );
  INV_X1 U5666 ( .A(n5869), .ZN(n4613) );
  NAND2_X1 U5667 ( .A1(n6716), .A2(n4570), .ZN(n4575) );
  INV_X1 U5668 ( .A(n6391), .ZN(n4982) );
  NOR2_X1 U5669 ( .A1(n4571), .A2(n4982), .ZN(n4572) );
  XNOR2_X1 U5670 ( .A(n4572), .B(n3570), .ZN(n6118) );
  NOR2_X1 U5671 ( .A1(n4748), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4573) );
  AND2_X1 U5672 ( .A1(n6118), .A2(n4573), .ZN(n4693) );
  INV_X1 U5673 ( .A(n4693), .ZN(n4574) );
  OAI22_X1 U5674 ( .A1(n4613), .A2(n3570), .B1(n4575), .B2(n4574), .ZN(U3455)
         );
  NOR2_X1 U5675 ( .A1(n4546), .A2(n4577), .ZN(n4578) );
  OR2_X1 U5676 ( .A1(n4650), .A2(n4578), .ZN(n6123) );
  OR2_X1 U5677 ( .A1(n4580), .A2(n4579), .ZN(n4581) );
  AND2_X1 U5678 ( .A1(n4655), .A2(n4581), .ZN(n6119) );
  AOI22_X1 U5679 ( .A1(n6178), .A2(n6119), .B1(n5641), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4582) );
  OAI21_X1 U5680 ( .B1(n6123), .B2(n5667), .A(n4582), .ZN(U2855) );
  NAND2_X1 U5681 ( .A1(n4584), .A2(n4583), .ZN(n4585) );
  NAND2_X1 U5682 ( .A1(n4586), .A2(n4585), .ZN(n6327) );
  INV_X1 U5683 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4590) );
  NOR2_X1 U5684 ( .A1(n4588), .A2(n4587), .ZN(n4589) );
  OR2_X1 U5685 ( .A1(n4547), .A2(n4589), .ZN(n6143) );
  OAI222_X1 U5686 ( .A1(n6327), .A2(n5666), .B1(n4590), .B2(n6182), .C1(n5667), 
        .C2(n6143), .ZN(U2857) );
  NAND2_X1 U5687 ( .A1(n4592), .A2(n4591), .ZN(n4593) );
  NAND2_X1 U5688 ( .A1(n4594), .A2(n4593), .ZN(n6302) );
  OAI222_X1 U5689 ( .A1(n6302), .A2(n5667), .B1(n6182), .B2(n5176), .C1(n5182), 
        .C2(n5666), .ZN(U2859) );
  NAND2_X1 U5690 ( .A1(n4597), .A2(n4596), .ZN(n4598) );
  NOR2_X1 U5691 ( .A1(n4599), .A2(n4598), .ZN(n4600) );
  AND2_X1 U5692 ( .A1(n4748), .A2(n4600), .ZN(n4601) );
  NAND2_X1 U5693 ( .A1(n4602), .A2(n4601), .ZN(n5538) );
  INV_X1 U5694 ( .A(n5537), .ZN(n6572) );
  CLKBUF_X1 U5695 ( .A(n4603), .Z(n4676) );
  INV_X1 U5696 ( .A(n4676), .ZN(n5563) );
  INV_X1 U5697 ( .A(n3010), .ZN(n4692) );
  NAND3_X1 U5698 ( .A1(n5541), .A2(n5563), .A3(n4692), .ZN(n4604) );
  OAI21_X1 U5699 ( .B1(n6572), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n4604), 
        .ZN(n4605) );
  AOI21_X1 U5700 ( .B1(n6163), .B2(n5538), .A(n4605), .ZN(n6573) );
  INV_X1 U5701 ( .A(n6611), .ZN(n5867) );
  AOI22_X1 U5702 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4607), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6339), .ZN(n5560) );
  NOR2_X1 U5703 ( .A1(n6614), .A2(n6331), .ZN(n5544) );
  AOI22_X1 U5704 ( .A1(n4608), .A2(n5562), .B1(n5560), .B2(n5544), .ZN(n4609)
         );
  OAI21_X1 U5705 ( .B1(n6573), .B2(n5867), .A(n4609), .ZN(n4611) );
  AOI22_X1 U5706 ( .A1(n4613), .A2(n4611), .B1(n4610), .B2(n5562), .ZN(n4612)
         );
  OAI21_X1 U5707 ( .B1(n3292), .B2(n4613), .A(n4612), .ZN(U3460) );
  OR2_X1 U5708 ( .A1(n4615), .A2(n4614), .ZN(n4616) );
  NAND2_X1 U5709 ( .A1(n4617), .A2(n4616), .ZN(n4921) );
  OR3_X1 U5710 ( .A1(n5030), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n4618), 
        .ZN(n4624) );
  AOI21_X1 U5711 ( .B1(n6331), .B2(n5462), .A(n4619), .ZN(n4620) );
  NAND2_X1 U5712 ( .A1(n6284), .A2(REIP_REG_1__SCAN_IN), .ZN(n4920) );
  OAI21_X1 U5713 ( .B1(n4620), .B2(n6339), .A(n4920), .ZN(n4621) );
  AOI21_X1 U5714 ( .B1(n6330), .B2(n4622), .A(n4621), .ZN(n4623) );
  OAI211_X1 U5715 ( .C1(n5997), .C2(n4921), .A(n4624), .B(n4623), .ZN(U3017)
         );
  NAND2_X1 U5716 ( .A1(n4625), .A2(n5537), .ZN(n4626) );
  NAND2_X1 U5717 ( .A1(n6282), .A2(n4626), .ZN(n4627) );
  NAND2_X1 U5718 ( .A1(n6210), .A2(n4628), .ZN(n6197) );
  NOR2_X1 U5719 ( .A1(n6619), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4645) );
  INV_X1 U5720 ( .A(n4645), .ZN(n6597) );
  AOI22_X1 U5721 ( .A1(n4645), .A2(UWORD_REG_0__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4629) );
  OAI21_X1 U5722 ( .B1(n3727), .B2(n6197), .A(n4629), .ZN(U2907) );
  AOI22_X1 U5723 ( .A1(n6730), .A2(UWORD_REG_14__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4630) );
  OAI21_X1 U5724 ( .B1(n6249), .B2(n6197), .A(n4630), .ZN(U2893) );
  AOI22_X1 U5725 ( .A1(n4645), .A2(UWORD_REG_2__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4631) );
  OAI21_X1 U5726 ( .B1(n3758), .B2(n6197), .A(n4631), .ZN(U2905) );
  INV_X1 U5727 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4633) );
  AOI22_X1 U5728 ( .A1(n4645), .A2(UWORD_REG_3__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4632) );
  OAI21_X1 U5729 ( .B1(n4633), .B2(n6197), .A(n4632), .ZN(U2904) );
  AOI22_X1 U5730 ( .A1(n4645), .A2(UWORD_REG_4__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4634) );
  OAI21_X1 U5731 ( .B1(n3796), .B2(n6197), .A(n4634), .ZN(U2903) );
  AOI22_X1 U5732 ( .A1(n4645), .A2(UWORD_REG_5__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4635) );
  OAI21_X1 U5733 ( .B1(n4636), .B2(n6197), .A(n4635), .ZN(U2902) );
  AOI22_X1 U5734 ( .A1(n4645), .A2(UWORD_REG_6__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4637) );
  OAI21_X1 U5735 ( .B1(n4638), .B2(n6197), .A(n4637), .ZN(U2901) );
  AOI22_X1 U5736 ( .A1(n4645), .A2(UWORD_REG_13__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4639) );
  OAI21_X1 U5737 ( .B1(n6246), .B2(n6197), .A(n4639), .ZN(U2894) );
  INV_X1 U5738 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4641) );
  AOI22_X1 U5739 ( .A1(n4645), .A2(UWORD_REG_7__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4640) );
  OAI21_X1 U5740 ( .B1(n4641), .B2(n6197), .A(n4640), .ZN(U2900) );
  INV_X1 U5741 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4643) );
  AOI22_X1 U5742 ( .A1(n4645), .A2(UWORD_REG_9__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4642) );
  OAI21_X1 U5743 ( .B1(n4643), .B2(n6197), .A(n4642), .ZN(U2898) );
  AOI22_X1 U5744 ( .A1(n6730), .A2(UWORD_REG_10__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4644) );
  OAI21_X1 U5745 ( .B1(n4176), .B2(n6197), .A(n4644), .ZN(U2897) );
  INV_X1 U5746 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4647) );
  AOI22_X1 U5747 ( .A1(n4645), .A2(UWORD_REG_11__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4646) );
  OAI21_X1 U5748 ( .B1(n4647), .B2(n6197), .A(n4646), .ZN(U2896) );
  AOI22_X1 U5749 ( .A1(n6730), .A2(UWORD_REG_12__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4648) );
  OAI21_X1 U5750 ( .B1(n4153), .B2(n6197), .A(n4648), .ZN(U2895) );
  INV_X1 U5751 ( .A(n4649), .ZN(n4653) );
  INV_X1 U5752 ( .A(n4650), .ZN(n4652) );
  AOI21_X1 U5753 ( .B1(n4653), .B2(n4652), .A(n4651), .ZN(n6113) );
  INV_X1 U5754 ( .A(n6113), .ZN(n4831) );
  INV_X1 U5755 ( .A(n4654), .ZN(n4713) );
  AOI21_X1 U5756 ( .B1(n4656), .B2(n4655), .A(n4713), .ZN(n6109) );
  AOI22_X1 U5757 ( .A1(n6178), .A2(n6109), .B1(n5641), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n4657) );
  OAI21_X1 U5758 ( .B1(n4831), .B2(n5667), .A(n4657), .ZN(U2854) );
  INV_X1 U5759 ( .A(n6273), .ZN(n6237) );
  AOI222_X1 U5760 ( .A1(n6276), .A2(LWORD_REG_15__SCAN_IN), .B1(n6237), .B2(
        DATAI_15_), .C1(EAX_REG_15__SCAN_IN), .C2(n6271), .ZN(n4659) );
  INV_X1 U5761 ( .A(n4659), .ZN(U2954) );
  NAND2_X1 U5762 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6017), .ZN(n4691) );
  INV_X1 U5763 ( .A(n4660), .ZN(n4690) );
  INV_X1 U5764 ( .A(n4662), .ZN(n4663) );
  OAI21_X1 U5765 ( .B1(n4676), .B2(n3110), .A(n4663), .ZN(n4665) );
  NOR2_X1 U5766 ( .A1(n4665), .A2(n4664), .ZN(n5866) );
  NAND2_X1 U5767 ( .A1(n4666), .A2(n4749), .ZN(n4677) );
  MUX2_X1 U5768 ( .A(n4667), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4676), 
        .Z(n4668) );
  NOR2_X1 U5769 ( .A1(n4668), .A2(n4660), .ZN(n4669) );
  NAND2_X1 U5770 ( .A1(n4677), .A2(n4669), .ZN(n4673) );
  XNOR2_X1 U5771 ( .A(n4670), .B(n3110), .ZN(n4671) );
  NAND2_X1 U5772 ( .A1(n5537), .A2(n4671), .ZN(n4672) );
  OAI211_X1 U5773 ( .C1(n5866), .C2(n4681), .A(n4673), .B(n4672), .ZN(n4674)
         );
  AOI21_X1 U5774 ( .B1(n2977), .B2(n5538), .A(n4674), .ZN(n5868) );
  MUX2_X1 U5775 ( .A(n5868), .B(n3110), .S(n6579), .Z(n6583) );
  INV_X1 U5776 ( .A(n6583), .ZN(n4688) );
  NAND2_X1 U5777 ( .A1(n5862), .A2(n5538), .ZN(n4685) );
  XNOR2_X1 U5778 ( .A(n4676), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4682)
         );
  NAND2_X1 U5779 ( .A1(n4677), .A2(n4682), .ZN(n4680) );
  XNOR2_X1 U5780 ( .A(n3099), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4678)
         );
  NAND2_X1 U5781 ( .A1(n5537), .A2(n4678), .ZN(n4679) );
  OAI211_X1 U5782 ( .C1(n4682), .C2(n4681), .A(n4680), .B(n4679), .ZN(n4683)
         );
  INV_X1 U5783 ( .A(n4683), .ZN(n4684) );
  NAND2_X1 U5784 ( .A1(n4685), .A2(n4684), .ZN(n5566) );
  OR2_X1 U5785 ( .A1(n6579), .A2(n5566), .ZN(n4687) );
  NAND2_X1 U5786 ( .A1(n6579), .A2(n3099), .ZN(n4686) );
  NAND3_X1 U5787 ( .A1(n4688), .A2(n6581), .A3(n6614), .ZN(n4689) );
  OAI21_X1 U5788 ( .B1(n4691), .B2(n4690), .A(n4689), .ZN(n6594) );
  NAND2_X1 U5789 ( .A1(n6594), .A2(n4692), .ZN(n4697) );
  MUX2_X1 U5790 ( .A(n6579), .B(n6017), .S(STATE2_REG_1__SCAN_IN), .Z(n4694)
         );
  AOI21_X1 U5791 ( .B1(n4694), .B2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(n4693), 
        .ZN(n6592) );
  AND3_X1 U5792 ( .A1(n4697), .A2(n6592), .A3(n6017), .ZN(n4695) );
  INV_X1 U5793 ( .A(n6735), .ZN(n6603) );
  INV_X1 U5794 ( .A(n6619), .ZN(n4696) );
  AND3_X1 U5795 ( .A1(n4697), .A2(n6592), .A3(n4696), .ZN(n6605) );
  AND2_X1 U5796 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6716), .ZN(n5863) );
  OAI22_X1 U5797 ( .A1(n5387), .A2(n6352), .B1(n5540), .B2(n5863), .ZN(n4698)
         );
  OAI21_X1 U5798 ( .B1(n6605), .B2(n4698), .A(n6344), .ZN(n4699) );
  OAI21_X1 U5799 ( .B1(n6344), .B2(n5385), .A(n4699), .ZN(U3465) );
  OR3_X1 U5800 ( .A1(n6345), .A2(n4704), .A3(n4702), .ZN(n5071) );
  INV_X1 U5801 ( .A(n5071), .ZN(n4703) );
  NAND2_X1 U5802 ( .A1(n4703), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5219) );
  AND2_X1 U5803 ( .A1(n6506), .A2(n5219), .ZN(n6347) );
  NAND2_X1 U5804 ( .A1(n4702), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6505) );
  INV_X1 U5805 ( .A(n6505), .ZN(n6346) );
  NAND2_X1 U5806 ( .A1(n6424), .A2(n6346), .ZN(n6425) );
  AOI21_X1 U5807 ( .B1(n6347), .B2(n6425), .A(n6352), .ZN(n4706) );
  NAND2_X1 U5808 ( .A1(n6513), .A2(n6015), .ZN(n6393) );
  OAI22_X1 U5809 ( .A1(n4726), .A2(n6393), .B1(n6467), .B2(n5863), .ZN(n4705)
         );
  OAI21_X1 U5810 ( .B1(n4706), .B2(n4705), .A(n6344), .ZN(n4707) );
  OAI21_X1 U5811 ( .B1(n6344), .B2(n6501), .A(n4707), .ZN(U3462) );
  CLKBUF_X1 U5812 ( .A(n4709), .Z(n4710) );
  OAI21_X1 U5813 ( .B1(n5044), .B2(n4711), .A(n4710), .ZN(n5166) );
  INV_X1 U5814 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4715) );
  AOI21_X1 U5815 ( .B1(n4713), .B2(n4941), .A(n4712), .ZN(n4714) );
  OR2_X1 U5816 ( .A1(n4714), .A2(n4760), .ZN(n6093) );
  OAI222_X1 U5817 ( .A1(n5166), .A2(n5667), .B1(n6182), .B2(n4715), .C1(n6093), 
        .C2(n5666), .ZN(U2852) );
  INV_X1 U5818 ( .A(n4841), .ZN(n4717) );
  AOI21_X1 U5819 ( .B1(n4717), .B2(n4716), .A(n6332), .ZN(n4943) );
  AOI211_X1 U5820 ( .C1(n3995), .C2(n3430), .A(n4943), .B(n6334), .ZN(n4723)
         );
  OAI21_X1 U5821 ( .B1(n4867), .B2(n4717), .A(n4865), .ZN(n6337) );
  AOI21_X1 U5822 ( .B1(n6332), .B2(n6334), .A(n6337), .ZN(n4785) );
  AND2_X1 U5823 ( .A1(n6284), .A2(REIP_REG_4__SCAN_IN), .ZN(n5057) );
  AOI21_X1 U5824 ( .B1(n6330), .B2(n6119), .A(n5057), .ZN(n4721) );
  XOR2_X1 U5825 ( .A(n4718), .B(n2966), .Z(n5056) );
  NAND2_X1 U5826 ( .A1(n5056), .A2(n6336), .ZN(n4720) );
  OAI211_X1 U5827 ( .C1(n4785), .C2(n3995), .A(n4721), .B(n4720), .ZN(n4722)
         );
  AOI21_X1 U5828 ( .B1(n4723), .B2(n4840), .A(n4722), .ZN(n4724) );
  INV_X1 U5829 ( .A(n4724), .ZN(U3014) );
  NAND3_X1 U5830 ( .A1(n6501), .A2(n6582), .A3(n6575), .ZN(n5345) );
  NOR2_X1 U5831 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5345), .ZN(n4955)
         );
  INV_X1 U5832 ( .A(n4955), .ZN(n4742) );
  AND2_X1 U5833 ( .A1(n4735), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6468) );
  NAND2_X1 U5834 ( .A1(n4726), .A2(n6345), .ZN(n4980) );
  INV_X1 U5835 ( .A(n6393), .ZN(n4729) );
  AOI21_X1 U5836 ( .B1(n4890), .B2(n6513), .A(n4729), .ZN(n5344) );
  NAND2_X1 U5837 ( .A1(n3350), .A2(n4702), .ZN(n4727) );
  OR2_X1 U5838 ( .A1(n5862), .A2(n6163), .ZN(n6466) );
  NOR2_X1 U5839 ( .A1(n2977), .A2(n6466), .ZN(n5342) );
  INV_X1 U5840 ( .A(n5342), .ZN(n4728) );
  OAI21_X1 U5841 ( .B1(n5149), .B2(n4729), .A(n4728), .ZN(n4730) );
  NOR2_X1 U5842 ( .A1(n5344), .A2(n4730), .ZN(n4731) );
  INV_X1 U5843 ( .A(n5064), .ZN(n6386) );
  NOR2_X1 U5844 ( .A1(n6386), .A2(n5065), .ZN(n4978) );
  OAI21_X1 U5845 ( .B1(n4978), .B2(n6514), .A(n4768), .ZN(n4985) );
  NOR3_X1 U5846 ( .A1(n6468), .A2(n4731), .A3(n4985), .ZN(n4732) );
  OAI21_X1 U5847 ( .B1(n4955), .B2(n6716), .A(n4732), .ZN(n4950) );
  NAND2_X1 U5848 ( .A1(n4950), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4741) );
  INV_X1 U5849 ( .A(n4890), .ZN(n4733) );
  INV_X1 U5850 ( .A(n5379), .ZN(n4739) );
  OR2_X1 U5851 ( .A1(n6301), .A2(n4388), .ZN(n6551) );
  INV_X1 U5852 ( .A(n6551), .ZN(n6486) );
  INV_X1 U5853 ( .A(DATAI_29_), .ZN(n4734) );
  OR2_X1 U5854 ( .A1(n6301), .A2(n4734), .ZN(n6489) );
  NAND2_X1 U5855 ( .A1(n5342), .A2(n6513), .ZN(n4737) );
  NOR2_X1 U5856 ( .A1(n4735), .A2(n6514), .ZN(n5075) );
  NAND2_X1 U5857 ( .A1(n5075), .A2(n4978), .ZN(n4736) );
  INV_X1 U5858 ( .A(DATAI_5_), .ZN(n6261) );
  OAI22_X1 U5859 ( .A1(n5149), .A2(n6489), .B1(n4958), .B2(n5367), .ZN(n4738)
         );
  AOI21_X1 U5860 ( .B1(n4739), .B2(n6486), .A(n4738), .ZN(n4740) );
  OAI211_X1 U5861 ( .C1(n4742), .C2(n5423), .A(n4741), .B(n4740), .ZN(U3025)
         );
  AOI21_X1 U5862 ( .B1(n4745), .B2(n4710), .A(n4744), .ZN(n5614) );
  INV_X1 U5863 ( .A(n5614), .ZN(n4764) );
  NAND2_X1 U5864 ( .A1(n6612), .A2(n4746), .ZN(n4747) );
  OAI22_X1 U5865 ( .A1(n4750), .A2(n4749), .B1(n4748), .B2(n4747), .ZN(n4751)
         );
  INV_X1 U5866 ( .A(n4751), .ZN(n4752) );
  AND2_X1 U5867 ( .A1(n4753), .A2(n5171), .ZN(n4754) );
  NAND2_X1 U5868 ( .A1(n4755), .A2(n5533), .ZN(n4756) );
  INV_X1 U5869 ( .A(n4756), .ZN(n4757) );
  INV_X1 U5870 ( .A(n5452), .ZN(n5340) );
  AOI22_X1 U5871 ( .A1(EAX_REG_8__SCAN_IN), .A2(n6193), .B1(n5340), .B2(
        DATAI_8_), .ZN(n4758) );
  OAI21_X1 U5872 ( .B1(n4764), .B2(n5935), .A(n4758), .ZN(U2883) );
  NOR2_X1 U5873 ( .A1(n4760), .A2(n4759), .ZN(n4761) );
  OR2_X1 U5874 ( .A1(n4880), .A2(n4761), .ZN(n5610) );
  INV_X1 U5875 ( .A(n5610), .ZN(n4762) );
  AOI22_X1 U5876 ( .A1(n6178), .A2(n4762), .B1(n5641), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n4763) );
  OAI21_X1 U5877 ( .B1(n4764), .B2(n5667), .A(n4763), .ZN(U2851) );
  INV_X1 U5878 ( .A(n5126), .ZN(n4765) );
  NOR2_X1 U5879 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4765), .ZN(n4771)
         );
  INV_X1 U5880 ( .A(n4771), .ZN(n4998) );
  NAND2_X1 U5881 ( .A1(n5862), .A2(n6163), .ZN(n6392) );
  INV_X1 U5882 ( .A(n5150), .ZN(n4766) );
  NOR2_X2 U5883 ( .A1(n5071), .A2(n5387), .ZN(n5247) );
  OAI21_X1 U5884 ( .B1(n4766), .B2(n5247), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4767) );
  NAND3_X1 U5885 ( .A1(n6392), .A2(n6513), .A3(n4767), .ZN(n4770) );
  OAI21_X1 U5886 ( .B1(n6386), .B2(n6514), .A(n4768), .ZN(n6397) );
  NOR3_X1 U5887 ( .A1(n6397), .A2(n6501), .A3(n5075), .ZN(n4769) );
  OAI211_X1 U5888 ( .C1(n4771), .C2(n6716), .A(n4770), .B(n4769), .ZN(n4995)
         );
  INV_X1 U5889 ( .A(DATAI_23_), .ZN(n4772) );
  OR2_X1 U5890 ( .A1(n6301), .A2(n4772), .ZN(n6570) );
  INV_X1 U5891 ( .A(DATAI_31_), .ZN(n4773) );
  OR2_X1 U5892 ( .A1(n6301), .A2(n4773), .ZN(n6500) );
  INV_X1 U5893 ( .A(n6500), .ZN(n6560) );
  INV_X1 U5894 ( .A(DATAI_7_), .ZN(n6264) );
  NAND2_X1 U5895 ( .A1(n2977), .A2(n6389), .ZN(n6463) );
  OR2_X1 U5896 ( .A1(n6463), .A2(n6392), .ZN(n4775) );
  NAND3_X1 U5897 ( .A1(n6468), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6386), .ZN(n4774) );
  NAND2_X1 U5898 ( .A1(n4775), .A2(n4774), .ZN(n4992) );
  AOI22_X1 U5899 ( .A1(n5247), .A2(n6560), .B1(n6565), .B2(n4992), .ZN(n4776)
         );
  OAI21_X1 U5900 ( .B1(n6570), .B2(n5150), .A(n4776), .ZN(n4777) );
  AOI21_X1 U5901 ( .B1(n4995), .B2(INSTQUEUE_REG_14__7__SCAN_IN), .A(n4777), 
        .ZN(n4778) );
  OAI21_X1 U5902 ( .B1(n5407), .B2(n4998), .A(n4778), .ZN(U3139) );
  INV_X1 U5903 ( .A(n6489), .ZN(n6546) );
  AOI22_X1 U5904 ( .A1(n5247), .A2(n6546), .B1(n6548), .B2(n4992), .ZN(n4779)
         );
  OAI21_X1 U5905 ( .B1(n6551), .B2(n5150), .A(n4779), .ZN(n4780) );
  AOI21_X1 U5906 ( .B1(n4995), .B2(INSTQUEUE_REG_14__5__SCAN_IN), .A(n4780), 
        .ZN(n4781) );
  OAI21_X1 U5907 ( .B1(n5423), .B2(n4998), .A(n4781), .ZN(U3137) );
  CLKBUF_X1 U5908 ( .A(n4782), .Z(n4783) );
  XNOR2_X1 U5909 ( .A(n4783), .B(n4784), .ZN(n5055) );
  NOR2_X1 U5910 ( .A1(n6334), .A2(n4943), .ZN(n4787) );
  INV_X1 U5911 ( .A(n4785), .ZN(n4786) );
  MUX2_X1 U5912 ( .A(n4787), .B(n4786), .S(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .Z(n4788) );
  INV_X1 U5913 ( .A(n4788), .ZN(n4790) );
  INV_X1 U5914 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6652) );
  NOR2_X1 U5915 ( .A1(n6309), .A2(n6652), .ZN(n5050) );
  AOI21_X1 U5916 ( .B1(n6330), .B2(n6139), .A(n5050), .ZN(n4789) );
  OAI211_X1 U5917 ( .C1(n5997), .C2(n5055), .A(n4790), .B(n4789), .ZN(U3015)
         );
  NAND2_X1 U5918 ( .A1(n5202), .A2(n5209), .ZN(n5211) );
  NAND2_X1 U5919 ( .A1(n5211), .A2(n6558), .ZN(n4791) );
  AOI21_X1 U5920 ( .B1(n4791), .B2(STATEBS16_REG_SCAN_IN), .A(n6352), .ZN(
        n4795) );
  INV_X1 U5921 ( .A(n6163), .ZN(n5860) );
  NOR2_X1 U5922 ( .A1(n5862), .A2(n5860), .ZN(n4892) );
  AND2_X1 U5923 ( .A1(n4892), .A2(n2977), .ZN(n6508) );
  INV_X1 U5924 ( .A(n5075), .ZN(n6462) );
  NOR3_X1 U5925 ( .A1(n6462), .A2(n6501), .A3(n5064), .ZN(n4792) );
  AOI21_X1 U5926 ( .B1(n4795), .B2(n6508), .A(n4792), .ZN(n4977) );
  INV_X1 U5927 ( .A(DATAI_4_), .ZN(n6259) );
  NOR2_X1 U5928 ( .A1(n6468), .A2(n6397), .ZN(n4895) );
  INV_X1 U5929 ( .A(n6508), .ZN(n4794) );
  NAND3_X1 U5930 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6582), .ZN(n6515) );
  NOR2_X1 U5931 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6515), .ZN(n4974)
         );
  INV_X1 U5932 ( .A(n4974), .ZN(n4793) );
  AOI22_X1 U5933 ( .A1(n4795), .A2(n4794), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n4793), .ZN(n4796) );
  OAI211_X1 U5934 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6514), .A(n4895), .B(n4796), .ZN(n4972) );
  NAND2_X1 U5935 ( .A1(n4972), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4801)
         );
  OR2_X1 U5936 ( .A1(n6301), .A2(n4797), .ZN(n6545) );
  INV_X1 U5937 ( .A(DATAI_20_), .ZN(n4798) );
  OR2_X1 U5938 ( .A1(n6301), .A2(n4798), .ZN(n6449) );
  OAI22_X1 U5939 ( .A1(n5211), .A2(n6545), .B1(n6558), .B2(n6449), .ZN(n4799)
         );
  AOI21_X1 U5940 ( .B1(n6541), .B2(n4974), .A(n4799), .ZN(n4800) );
  OAI211_X1 U5941 ( .C1(n4977), .C2(n5383), .A(n4801), .B(n4800), .ZN(U3104)
         );
  INV_X1 U5942 ( .A(DATAI_1_), .ZN(n6253) );
  NAND2_X1 U5943 ( .A1(n4972), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4807)
         );
  OR2_X1 U5944 ( .A1(n6301), .A2(n4803), .ZN(n6527) );
  INV_X1 U5945 ( .A(DATAI_17_), .ZN(n4804) );
  OR2_X1 U5946 ( .A1(n6301), .A2(n4804), .ZN(n6438) );
  OAI22_X1 U5947 ( .A1(n5211), .A2(n6527), .B1(n6558), .B2(n6438), .ZN(n4805)
         );
  AOI21_X1 U5948 ( .B1(n6523), .B2(n4974), .A(n4805), .ZN(n4806) );
  OAI211_X1 U5949 ( .C1(n4977), .C2(n5371), .A(n4807), .B(n4806), .ZN(U3101)
         );
  INV_X1 U5950 ( .A(DATAI_2_), .ZN(n6255) );
  NAND2_X1 U5951 ( .A1(n4972), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4812)
         );
  OR2_X1 U5952 ( .A1(n6301), .A2(n4808), .ZN(n6533) );
  INV_X1 U5953 ( .A(DATAI_18_), .ZN(n4809) );
  OR2_X1 U5954 ( .A1(n6301), .A2(n4809), .ZN(n6442) );
  OAI22_X1 U5955 ( .A1(n5211), .A2(n6533), .B1(n6558), .B2(n6442), .ZN(n4810)
         );
  AOI21_X1 U5956 ( .B1(n6529), .B2(n4974), .A(n4810), .ZN(n4811) );
  OAI211_X1 U5957 ( .C1(n4977), .C2(n5363), .A(n4812), .B(n4811), .ZN(U3102)
         );
  INV_X1 U5958 ( .A(DATAI_0_), .ZN(n6251) );
  NAND2_X1 U5959 ( .A1(n4972), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4818)
         );
  INV_X1 U5960 ( .A(DATAI_24_), .ZN(n4814) );
  OR2_X1 U5961 ( .A1(n6301), .A2(n4814), .ZN(n6477) );
  INV_X1 U5962 ( .A(DATAI_16_), .ZN(n4815) );
  OR2_X1 U5963 ( .A1(n6301), .A2(n4815), .ZN(n6521) );
  OAI22_X1 U5964 ( .A1(n5211), .A2(n6477), .B1(n6558), .B2(n6521), .ZN(n4816)
         );
  AOI21_X1 U5965 ( .B1(n6504), .B2(n4974), .A(n4816), .ZN(n4817) );
  OAI211_X1 U5966 ( .C1(n4977), .C2(n5375), .A(n4818), .B(n4817), .ZN(U3100)
         );
  NAND2_X1 U5967 ( .A1(n4972), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4821)
         );
  OAI22_X1 U5968 ( .A1(n5211), .A2(n6500), .B1(n6558), .B2(n6570), .ZN(n4819)
         );
  AOI21_X1 U5969 ( .B1(n6563), .B2(n4974), .A(n4819), .ZN(n4820) );
  OAI211_X1 U5970 ( .C1(n4977), .C2(n5356), .A(n4821), .B(n4820), .ZN(U3107)
         );
  NAND2_X1 U5971 ( .A1(n4972), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4827)
         );
  INV_X1 U5972 ( .A(DATAI_27_), .ZN(n4823) );
  OR2_X1 U5973 ( .A1(n6301), .A2(n4823), .ZN(n6539) );
  INV_X1 U5974 ( .A(DATAI_19_), .ZN(n4824) );
  OR2_X1 U5975 ( .A1(n6301), .A2(n4824), .ZN(n6407) );
  OAI22_X1 U5976 ( .A1(n5211), .A2(n6539), .B1(n6558), .B2(n6407), .ZN(n4825)
         );
  AOI21_X1 U5977 ( .B1(n6535), .B2(n4974), .A(n4825), .ZN(n4826) );
  OAI211_X1 U5978 ( .C1(n4977), .C2(n5352), .A(n4827), .B(n4826), .ZN(U3103)
         );
  NAND2_X1 U5979 ( .A1(n4972), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4830)
         );
  OAI22_X1 U5980 ( .A1(n5211), .A2(n6489), .B1(n6558), .B2(n6551), .ZN(n4828)
         );
  AOI21_X1 U5981 ( .B1(n6547), .B2(n4974), .A(n4828), .ZN(n4829) );
  OAI211_X1 U5982 ( .C1(n4977), .C2(n5367), .A(n4830), .B(n4829), .ZN(U3105)
         );
  OAI222_X1 U5983 ( .A1(n6302), .A2(n5935), .B1(n5452), .B2(n6251), .C1(n5668), 
        .C2(n3546), .ZN(U2891) );
  INV_X1 U5984 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6222) );
  OAI222_X1 U5985 ( .A1(n6123), .A2(n5935), .B1(n5452), .B2(n6259), .C1(n5668), 
        .C2(n6222), .ZN(U2887) );
  OAI222_X1 U5986 ( .A1(n6143), .A2(n5935), .B1(n5452), .B2(n6255), .C1(n5668), 
        .C2(n3554), .ZN(U2889) );
  INV_X1 U5987 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6220) );
  OAI222_X1 U5988 ( .A1(n4831), .A2(n5935), .B1(n5452), .B2(n6261), .C1(n5668), 
        .C2(n6220), .ZN(U2886) );
  OAI222_X1 U5989 ( .A1(n6137), .A2(n5935), .B1(n5452), .B2(n6257), .C1(n5668), 
        .C2(n3563), .ZN(U2888) );
  INV_X1 U5990 ( .A(n6477), .ZN(n6503) );
  AOI22_X1 U5991 ( .A1(n5247), .A2(n6503), .B1(n6518), .B2(n4992), .ZN(n4832)
         );
  OAI21_X1 U5992 ( .B1(n6521), .B2(n5150), .A(n4832), .ZN(n4833) );
  AOI21_X1 U5993 ( .B1(n4995), .B2(INSTQUEUE_REG_14__0__SCAN_IN), .A(n4833), 
        .ZN(n4834) );
  OAI21_X1 U5994 ( .B1(n5411), .B2(n4998), .A(n4834), .ZN(U3132) );
  INV_X1 U5995 ( .A(n6539), .ZN(n6404) );
  AOI22_X1 U5996 ( .A1(n5247), .A2(n6404), .B1(n6536), .B2(n4992), .ZN(n4835)
         );
  OAI21_X1 U5997 ( .B1(n6407), .B2(n5150), .A(n4835), .ZN(n4836) );
  AOI21_X1 U5998 ( .B1(n4995), .B2(INSTQUEUE_REG_14__3__SCAN_IN), .A(n4836), 
        .ZN(n4837) );
  OAI21_X1 U5999 ( .B1(n5403), .B2(n4998), .A(n4837), .ZN(U3135) );
  XNOR2_X1 U6000 ( .A(n4838), .B(n4839), .ZN(n5307) );
  NOR2_X1 U6001 ( .A1(n6309), .A2(n6655), .ZN(n5303) );
  INV_X1 U6002 ( .A(n4840), .ZN(n4843) );
  NOR2_X1 U6003 ( .A1(n4841), .A2(n6338), .ZN(n4842) );
  AOI22_X1 U6004 ( .A1(n6332), .A2(n4844), .B1(n4843), .B2(n4842), .ZN(n4846)
         );
  NAND2_X1 U6005 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4844), .ZN(n4942)
         );
  AOI21_X1 U6006 ( .B1(n5977), .B2(n4942), .A(n6337), .ZN(n4944) );
  AOI21_X1 U6007 ( .B1(n4846), .B2(n4845), .A(n4944), .ZN(n4847) );
  AOI211_X1 U6008 ( .C1(n6330), .C2(n6109), .A(n5303), .B(n4847), .ZN(n4848)
         );
  OAI21_X1 U6009 ( .B1(n5997), .B2(n5307), .A(n4848), .ZN(U3013) );
  INV_X1 U6010 ( .A(n6545), .ZN(n6446) );
  AOI22_X1 U6011 ( .A1(n5247), .A2(n6446), .B1(n6542), .B2(n4992), .ZN(n4849)
         );
  OAI21_X1 U6012 ( .B1(n6449), .B2(n5150), .A(n4849), .ZN(n4850) );
  AOI21_X1 U6013 ( .B1(n4995), .B2(INSTQUEUE_REG_14__4__SCAN_IN), .A(n4850), 
        .ZN(n4851) );
  OAI21_X1 U6014 ( .B1(n5419), .B2(n4998), .A(n4851), .ZN(U3136) );
  INV_X1 U6015 ( .A(n6533), .ZN(n6439) );
  AOI22_X1 U6016 ( .A1(n5247), .A2(n6439), .B1(n6530), .B2(n4992), .ZN(n4852)
         );
  OAI21_X1 U6017 ( .B1(n6442), .B2(n5150), .A(n4852), .ZN(n4853) );
  AOI21_X1 U6018 ( .B1(n4995), .B2(INSTQUEUE_REG_14__2__SCAN_IN), .A(n4853), 
        .ZN(n4854) );
  OAI21_X1 U6019 ( .B1(n5415), .B2(n4998), .A(n4854), .ZN(U3134) );
  INV_X1 U6020 ( .A(n6527), .ZN(n6435) );
  AOI22_X1 U6021 ( .A1(n5247), .A2(n6435), .B1(n6524), .B2(n4992), .ZN(n4855)
         );
  OAI21_X1 U6022 ( .B1(n6438), .B2(n5150), .A(n4855), .ZN(n4856) );
  AOI21_X1 U6023 ( .B1(n4995), .B2(INSTQUEUE_REG_14__1__SCAN_IN), .A(n4856), 
        .ZN(n4857) );
  OAI21_X1 U6024 ( .B1(n5431), .B2(n4998), .A(n4857), .ZN(U3133) );
  NOR2_X1 U6025 ( .A1(n5379), .A2(n6570), .ZN(n4859) );
  OAI22_X1 U6026 ( .A1(n5149), .A2(n6500), .B1(n4958), .B2(n5356), .ZN(n4858)
         );
  AOI211_X1 U6027 ( .C1(n6563), .C2(n4955), .A(n4859), .B(n4858), .ZN(n4860)
         );
  OAI21_X1 U6028 ( .B1(n4937), .B2(n4861), .A(n4860), .ZN(U3027) );
  XNOR2_X1 U6029 ( .A(n4864), .B(n4863), .ZN(n5317) );
  AOI21_X1 U6030 ( .B1(n4012), .B2(n3475), .A(n5031), .ZN(n4872) );
  NOR2_X1 U6031 ( .A1(n4943), .A2(n4869), .ZN(n6318) );
  OAI21_X1 U6032 ( .B1(n4867), .B2(n4866), .A(n4865), .ZN(n4868) );
  AOI21_X1 U6033 ( .B1(n6332), .B2(n4869), .A(n4868), .ZN(n6326) );
  OR2_X1 U6034 ( .A1(n6326), .A2(n4012), .ZN(n4870) );
  NAND2_X1 U6035 ( .A1(n6284), .A2(REIP_REG_8__SCAN_IN), .ZN(n5313) );
  OAI211_X1 U6036 ( .C1(n5996), .C2(n5610), .A(n4870), .B(n5313), .ZN(n4871)
         );
  AOI21_X1 U6037 ( .B1(n4872), .B2(n6318), .A(n4871), .ZN(n4873) );
  OAI21_X1 U6038 ( .B1(n5997), .B2(n5317), .A(n4873), .ZN(U3010) );
  CLKBUF_X1 U6039 ( .A(n4874), .Z(n4875) );
  OR2_X1 U6040 ( .A1(n4744), .A2(n4876), .ZN(n4877) );
  NAND2_X1 U6041 ( .A1(n4875), .A2(n4877), .ZN(n5201) );
  INV_X1 U6042 ( .A(DATAI_9_), .ZN(n6268) );
  OAI222_X1 U6043 ( .A1(n5201), .A2(n5935), .B1(n5452), .B2(n6268), .C1(n5668), 
        .C2(n3623), .ZN(U2882) );
  OAI21_X1 U6044 ( .B1(n4880), .B2(n4879), .A(n4878), .ZN(n5185) );
  INV_X1 U6045 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4881) );
  OAI222_X1 U6046 ( .A1(n5185), .A2(n5666), .B1(n4881), .B2(n6182), .C1(n5667), 
        .C2(n5201), .ZN(U2850) );
  INV_X1 U6047 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4885) );
  NOR2_X1 U6048 ( .A1(n5379), .A2(n6407), .ZN(n4883) );
  OAI22_X1 U6049 ( .A1(n5149), .A2(n6539), .B1(n4958), .B2(n5352), .ZN(n4882)
         );
  AOI211_X1 U6050 ( .C1(n6535), .C2(n4955), .A(n4883), .B(n4882), .ZN(n4884)
         );
  OAI21_X1 U6051 ( .B1(n4937), .B2(n4885), .A(n4884), .ZN(U3023) );
  NOR2_X1 U6052 ( .A1(n5379), .A2(n6521), .ZN(n4887) );
  OAI22_X1 U6053 ( .A1(n5149), .A2(n6477), .B1(n4958), .B2(n5375), .ZN(n4886)
         );
  AOI211_X1 U6054 ( .C1(n6504), .C2(n4955), .A(n4887), .B(n4886), .ZN(n4888)
         );
  OAI21_X1 U6055 ( .B1(n4937), .B2(n4889), .A(n4888), .ZN(U3020) );
  NAND3_X1 U6056 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6501), .A3(n6582), .ZN(n6353) );
  NOR2_X1 U6057 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6353), .ZN(n4968)
         );
  INV_X1 U6058 ( .A(n4968), .ZN(n4919) );
  NOR2_X2 U6059 ( .A1(n4890), .A2(n5387), .ZN(n5377) );
  INV_X1 U6060 ( .A(n6385), .ZN(n4891) );
  OAI21_X1 U6061 ( .B1(n5377), .B2(n6377), .A(n6393), .ZN(n4894) );
  INV_X1 U6062 ( .A(n6349), .ZN(n4893) );
  AOI21_X1 U6063 ( .B1(n4894), .B2(n4893), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4896) );
  NAND2_X1 U6064 ( .A1(n4964), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4900) );
  NOR3_X1 U6065 ( .A1(n6462), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n5064), 
        .ZN(n4897) );
  AOI21_X1 U6066 ( .B1(n6349), .B2(n6513), .A(n4897), .ZN(n4971) );
  OAI22_X1 U6067 ( .A1(n4965), .A2(n6521), .B1(n4971), .B2(n5375), .ZN(n4898)
         );
  AOI21_X1 U6068 ( .B1(n5377), .B2(n6503), .A(n4898), .ZN(n4899) );
  OAI211_X1 U6069 ( .C1(n5411), .C2(n4919), .A(n4900), .B(n4899), .ZN(U3036)
         );
  NAND2_X1 U6070 ( .A1(n4964), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4903) );
  OAI22_X1 U6071 ( .A1(n4965), .A2(n6407), .B1(n4971), .B2(n5352), .ZN(n4901)
         );
  AOI21_X1 U6072 ( .B1(n5377), .B2(n6404), .A(n4901), .ZN(n4902) );
  OAI211_X1 U6073 ( .C1(n4919), .C2(n5403), .A(n4903), .B(n4902), .ZN(U3039)
         );
  NAND2_X1 U6074 ( .A1(n4964), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4906) );
  OAI22_X1 U6075 ( .A1(n4965), .A2(n6551), .B1(n4971), .B2(n5367), .ZN(n4904)
         );
  AOI21_X1 U6076 ( .B1(n5377), .B2(n6546), .A(n4904), .ZN(n4905) );
  OAI211_X1 U6077 ( .C1(n4919), .C2(n5423), .A(n4906), .B(n4905), .ZN(U3041)
         );
  NAND2_X1 U6078 ( .A1(n4964), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4909) );
  OAI22_X1 U6079 ( .A1(n4965), .A2(n6449), .B1(n4971), .B2(n5383), .ZN(n4907)
         );
  AOI21_X1 U6080 ( .B1(n5377), .B2(n6446), .A(n4907), .ZN(n4908) );
  OAI211_X1 U6081 ( .C1(n4919), .C2(n5419), .A(n4909), .B(n4908), .ZN(U3040)
         );
  NAND2_X1 U6082 ( .A1(n4964), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4912) );
  OAI22_X1 U6083 ( .A1(n4965), .A2(n6438), .B1(n4971), .B2(n5371), .ZN(n4910)
         );
  AOI21_X1 U6084 ( .B1(n5377), .B2(n6435), .A(n4910), .ZN(n4911) );
  OAI211_X1 U6085 ( .C1(n4919), .C2(n5431), .A(n4912), .B(n4911), .ZN(U3037)
         );
  NAND2_X1 U6086 ( .A1(n4964), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4915) );
  OAI22_X1 U6087 ( .A1(n4965), .A2(n6570), .B1(n4971), .B2(n5356), .ZN(n4913)
         );
  AOI21_X1 U6088 ( .B1(n5377), .B2(n6560), .A(n4913), .ZN(n4914) );
  OAI211_X1 U6089 ( .C1(n4919), .C2(n5407), .A(n4915), .B(n4914), .ZN(U3043)
         );
  NAND2_X1 U6090 ( .A1(n4964), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4918) );
  OAI22_X1 U6091 ( .A1(n4965), .A2(n6442), .B1(n4971), .B2(n5363), .ZN(n4916)
         );
  AOI21_X1 U6092 ( .B1(n5377), .B2(n6439), .A(n4916), .ZN(n4917) );
  OAI211_X1 U6093 ( .C1(n4919), .C2(n5415), .A(n4918), .B(n4917), .ZN(U3038)
         );
  OAI21_X1 U6094 ( .B1(n6167), .B2(n6301), .A(n4920), .ZN(n4923) );
  NOR2_X1 U6095 ( .A1(n6016), .A2(n4921), .ZN(n4922) );
  AOI211_X1 U6096 ( .C1(n6298), .C2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4923), 
        .B(n4922), .ZN(n4924) );
  OAI21_X1 U6097 ( .B1(n5955), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4924), 
        .ZN(U2985) );
  INV_X1 U6098 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4928) );
  NOR2_X1 U6099 ( .A1(n5379), .A2(n6438), .ZN(n4926) );
  OAI22_X1 U6100 ( .A1(n5149), .A2(n6527), .B1(n4958), .B2(n5371), .ZN(n4925)
         );
  AOI211_X1 U6101 ( .C1(n6523), .C2(n4955), .A(n4926), .B(n4925), .ZN(n4927)
         );
  OAI21_X1 U6102 ( .B1(n4937), .B2(n4928), .A(n4927), .ZN(U3021) );
  NOR2_X1 U6103 ( .A1(n5379), .A2(n6449), .ZN(n4930) );
  OAI22_X1 U6104 ( .A1(n5149), .A2(n6545), .B1(n4958), .B2(n5383), .ZN(n4929)
         );
  AOI211_X1 U6105 ( .C1(n6541), .C2(n4955), .A(n4930), .B(n4929), .ZN(n4931)
         );
  OAI21_X1 U6106 ( .B1(n4937), .B2(n4932), .A(n4931), .ZN(U3024) );
  INV_X1 U6107 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4936) );
  NOR2_X1 U6108 ( .A1(n5379), .A2(n6442), .ZN(n4934) );
  OAI22_X1 U6109 ( .A1(n5149), .A2(n6533), .B1(n4958), .B2(n5363), .ZN(n4933)
         );
  AOI211_X1 U6110 ( .C1(n6529), .C2(n4955), .A(n4934), .B(n4933), .ZN(n4935)
         );
  OAI21_X1 U6111 ( .B1(n4937), .B2(n4936), .A(n4935), .ZN(U3022) );
  CLKBUF_X1 U6112 ( .A(n4938), .Z(n4939) );
  XNOR2_X1 U6113 ( .A(n4940), .B(n4939), .ZN(n5311) );
  XNOR2_X1 U6114 ( .A(n4654), .B(n4941), .ZN(n6177) );
  INV_X1 U6115 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6658) );
  NOR2_X1 U6116 ( .A1(n6309), .A2(n6658), .ZN(n4948) );
  NOR2_X1 U6117 ( .A1(n4943), .A2(n4942), .ZN(n4946) );
  INV_X1 U6118 ( .A(n4944), .ZN(n4945) );
  MUX2_X1 U6119 ( .A(n4946), .B(n4945), .S(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .Z(n4947) );
  AOI211_X1 U6120 ( .C1(n6330), .C2(n6177), .A(n4948), .B(n4947), .ZN(n4949)
         );
  OAI21_X1 U6121 ( .B1(n5997), .B2(n5311), .A(n4949), .ZN(U3012) );
  NAND2_X1 U6122 ( .A1(n4950), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4957) );
  NOR2_X2 U6123 ( .A1(n4951), .A2(n3529), .ZN(n6554) );
  INV_X1 U6124 ( .A(DATAI_22_), .ZN(n4952) );
  OR2_X1 U6125 ( .A1(n6301), .A2(n4952), .ZN(n6415) );
  OR2_X1 U6126 ( .A1(n6301), .A2(n4953), .ZN(n6559) );
  OAI22_X1 U6127 ( .A1(n5379), .A2(n6415), .B1(n6559), .B2(n5149), .ZN(n4954)
         );
  AOI21_X1 U6128 ( .B1(n6554), .B2(n4955), .A(n4954), .ZN(n4956) );
  OAI211_X1 U6129 ( .C1(n4958), .C2(n5398), .A(n4957), .B(n4956), .ZN(U3026)
         );
  NAND2_X1 U6130 ( .A1(n4878), .A2(n4959), .ZN(n4960) );
  NAND2_X1 U6131 ( .A1(n5039), .A2(n4960), .ZN(n5298) );
  OAI21_X1 U6132 ( .B1(n3640), .B2(n3639), .A(n4962), .ZN(n5302) );
  OAI222_X1 U6133 ( .A1(n5298), .A2(n5666), .B1(n6182), .B2(n4963), .C1(n5667), 
        .C2(n5302), .ZN(U2849) );
  NAND2_X1 U6134 ( .A1(n4964), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4970) );
  INV_X1 U6135 ( .A(n5377), .ZN(n4966) );
  OAI22_X1 U6136 ( .A1(n4966), .A2(n6559), .B1(n6415), .B2(n4965), .ZN(n4967)
         );
  AOI21_X1 U6137 ( .B1(n6554), .B2(n4968), .A(n4967), .ZN(n4969) );
  OAI211_X1 U6138 ( .C1(n4971), .C2(n5398), .A(n4970), .B(n4969), .ZN(U3042)
         );
  NAND2_X1 U6139 ( .A1(n4972), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4976)
         );
  OAI22_X1 U6140 ( .A1(n5211), .A2(n6559), .B1(n6558), .B2(n6415), .ZN(n4973)
         );
  AOI21_X1 U6141 ( .B1(n6554), .B2(n4974), .A(n4973), .ZN(n4975) );
  OAI211_X1 U6142 ( .C1(n4977), .C2(n5398), .A(n4976), .B(n4975), .ZN(U3106)
         );
  NAND2_X1 U6143 ( .A1(n6467), .A2(n6389), .ZN(n6388) );
  INV_X1 U6144 ( .A(n6388), .ZN(n4979) );
  AOI22_X1 U6145 ( .A1(n4979), .A2(n5217), .B1(n4978), .B2(n6468), .ZN(n5001)
         );
  NAND3_X1 U6146 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6501), .A3(n6575), .ZN(n5390) );
  NOR2_X1 U6147 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5390), .ZN(n4999)
         );
  NAND2_X1 U6148 ( .A1(n4702), .A2(n5209), .ZN(n5069) );
  NOR2_X2 U6149 ( .A1(n4980), .A2(n5069), .ZN(n6380) );
  INV_X1 U6150 ( .A(n6380), .ZN(n4989) );
  INV_X1 U6151 ( .A(n6424), .ZN(n4981) );
  NOR3_X1 U6152 ( .A1(n4981), .A2(n5209), .A3(n4702), .ZN(n5000) );
  INV_X1 U6153 ( .A(n6415), .ZN(n6553) );
  AND2_X1 U6154 ( .A1(n5217), .A2(n4982), .ZN(n5386) );
  NAND3_X1 U6155 ( .A1(n6424), .A2(n4983), .A3(STATEBS16_REG_SCAN_IN), .ZN(
        n4984) );
  NAND2_X1 U6156 ( .A1(n4984), .A2(n6389), .ZN(n5389) );
  AOI211_X1 U6157 ( .C1(n6380), .C2(n6393), .A(n5386), .B(n5389), .ZN(n4986)
         );
  NOR3_X1 U6158 ( .A1(n5075), .A2(n4986), .A3(n4985), .ZN(n4987) );
  OAI21_X1 U6159 ( .B1(n4999), .B2(n6716), .A(n4987), .ZN(n5020) );
  AOI22_X1 U6160 ( .A1(n5000), .A2(n6553), .B1(INSTQUEUE_REG_4__6__SCAN_IN), 
        .B2(n5020), .ZN(n4988) );
  OAI21_X1 U6161 ( .B1(n6559), .B2(n4989), .A(n4988), .ZN(n4990) );
  AOI21_X1 U6162 ( .B1(n6554), .B2(n4999), .A(n4990), .ZN(n4991) );
  OAI21_X1 U6163 ( .B1(n5398), .B2(n5001), .A(n4991), .ZN(U3058) );
  INV_X1 U6164 ( .A(n6554), .ZN(n5256) );
  NAND2_X1 U6165 ( .A1(n6555), .A2(n4992), .ZN(n4997) );
  INV_X1 U6166 ( .A(n5247), .ZN(n4993) );
  OAI22_X1 U6167 ( .A1(n4993), .A2(n6559), .B1(n6415), .B2(n5150), .ZN(n4994)
         );
  AOI21_X1 U6168 ( .B1(n4995), .B2(INSTQUEUE_REG_14__6__SCAN_IN), .A(n4994), 
        .ZN(n4996) );
  OAI211_X1 U6169 ( .C1(n5256), .C2(n4998), .A(n4997), .B(n4996), .ZN(U3138)
         );
  INV_X1 U6170 ( .A(n4999), .ZN(n5025) );
  INV_X1 U6171 ( .A(n5001), .ZN(n5021) );
  AOI22_X1 U6172 ( .A1(n5021), .A2(n6542), .B1(INSTQUEUE_REG_4__4__SCAN_IN), 
        .B2(n5020), .ZN(n5002) );
  OAI21_X1 U6173 ( .B1(n5426), .B2(n6449), .A(n5002), .ZN(n5003) );
  AOI21_X1 U6174 ( .B1(n6446), .B2(n6380), .A(n5003), .ZN(n5004) );
  OAI21_X1 U6175 ( .B1(n5419), .B2(n5025), .A(n5004), .ZN(U3056) );
  AOI22_X1 U6176 ( .A1(n5021), .A2(n6524), .B1(INSTQUEUE_REG_4__1__SCAN_IN), 
        .B2(n5020), .ZN(n5005) );
  OAI21_X1 U6177 ( .B1(n5426), .B2(n6438), .A(n5005), .ZN(n5006) );
  AOI21_X1 U6178 ( .B1(n6435), .B2(n6380), .A(n5006), .ZN(n5007) );
  OAI21_X1 U6179 ( .B1(n5431), .B2(n5025), .A(n5007), .ZN(U3053) );
  AOI22_X1 U6180 ( .A1(n5021), .A2(n6530), .B1(INSTQUEUE_REG_4__2__SCAN_IN), 
        .B2(n5020), .ZN(n5008) );
  OAI21_X1 U6181 ( .B1(n5426), .B2(n6442), .A(n5008), .ZN(n5009) );
  AOI21_X1 U6182 ( .B1(n6439), .B2(n6380), .A(n5009), .ZN(n5010) );
  OAI21_X1 U6183 ( .B1(n5415), .B2(n5025), .A(n5010), .ZN(U3054) );
  AOI22_X1 U6184 ( .A1(n5021), .A2(n6518), .B1(INSTQUEUE_REG_4__0__SCAN_IN), 
        .B2(n5020), .ZN(n5011) );
  OAI21_X1 U6185 ( .B1(n5426), .B2(n6521), .A(n5011), .ZN(n5012) );
  AOI21_X1 U6186 ( .B1(n6503), .B2(n6380), .A(n5012), .ZN(n5013) );
  OAI21_X1 U6187 ( .B1(n5411), .B2(n5025), .A(n5013), .ZN(U3052) );
  AOI22_X1 U6188 ( .A1(n5021), .A2(n6536), .B1(INSTQUEUE_REG_4__3__SCAN_IN), 
        .B2(n5020), .ZN(n5014) );
  OAI21_X1 U6189 ( .B1(n5426), .B2(n6407), .A(n5014), .ZN(n5015) );
  AOI21_X1 U6190 ( .B1(n6404), .B2(n6380), .A(n5015), .ZN(n5016) );
  OAI21_X1 U6191 ( .B1(n5403), .B2(n5025), .A(n5016), .ZN(U3055) );
  AOI22_X1 U6192 ( .A1(n5021), .A2(n6565), .B1(INSTQUEUE_REG_4__7__SCAN_IN), 
        .B2(n5020), .ZN(n5017) );
  OAI21_X1 U6193 ( .B1(n5426), .B2(n6570), .A(n5017), .ZN(n5018) );
  AOI21_X1 U6194 ( .B1(n6560), .B2(n6380), .A(n5018), .ZN(n5019) );
  OAI21_X1 U6195 ( .B1(n5407), .B2(n5025), .A(n5019), .ZN(U3059) );
  AOI22_X1 U6196 ( .A1(n5021), .A2(n6548), .B1(INSTQUEUE_REG_4__5__SCAN_IN), 
        .B2(n5020), .ZN(n5022) );
  OAI21_X1 U6197 ( .B1(n5426), .B2(n6551), .A(n5022), .ZN(n5023) );
  AOI21_X1 U6198 ( .B1(n6546), .B2(n6380), .A(n5023), .ZN(n5024) );
  OAI21_X1 U6199 ( .B1(n5423), .B2(n5025), .A(n5024), .ZN(U3057) );
  NAND2_X1 U6200 ( .A1(n2988), .A2(n5027), .ZN(n5028) );
  XNOR2_X1 U6201 ( .A(n5029), .B(n5028), .ZN(n5086) );
  OAI21_X1 U6202 ( .B1(n5030), .B2(n5031), .A(n6326), .ZN(n6313) );
  INV_X1 U6203 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6662) );
  OAI22_X1 U6204 ( .A1(n5996), .A2(n5298), .B1(n6662), .B2(n6309), .ZN(n5034)
         );
  NAND2_X1 U6205 ( .A1(n5031), .A2(n6318), .ZN(n6317) );
  AOI221_X1 U6206 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n5032), .C2(n5194), .A(n6317), 
        .ZN(n5033) );
  AOI211_X1 U6207 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n6313), .A(n5034), .B(n5033), .ZN(n5035) );
  OAI21_X1 U6208 ( .B1(n5997), .B2(n5086), .A(n5035), .ZN(U3008) );
  AOI21_X1 U6209 ( .B1(n5037), .B2(n4962), .A(n5160), .ZN(n5270) );
  INV_X1 U6210 ( .A(n5270), .ZN(n5284) );
  AND2_X1 U6211 ( .A1(n5039), .A2(n5038), .ZN(n5040) );
  NOR2_X1 U6212 ( .A1(n5326), .A2(n5040), .ZN(n6303) );
  AOI22_X1 U6213 ( .A1(n6178), .A2(n6303), .B1(n5641), .B2(EBX_REG_11__SCAN_IN), .ZN(n5041) );
  OAI21_X1 U6214 ( .B1(n5284), .B2(n5667), .A(n5041), .ZN(U2848) );
  OAI222_X1 U6215 ( .A1(n6167), .A2(n5935), .B1(n5452), .B2(n6253), .C1(n5668), 
        .C2(n3538), .ZN(U2890) );
  INV_X1 U6216 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6213) );
  OAI222_X1 U6217 ( .A1(n5302), .A2(n5935), .B1(n5452), .B2(n6270), .C1(n5668), 
        .C2(n6213), .ZN(U2881) );
  INV_X1 U6218 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5042) );
  OAI222_X1 U6219 ( .A1(n5284), .A2(n5935), .B1(n5452), .B2(n6274), .C1(n5668), 
        .C2(n5042), .ZN(U2880) );
  OAI222_X1 U6220 ( .A1(n5166), .A2(n5935), .B1(n5452), .B2(n6264), .C1(n5668), 
        .C2(n3533), .ZN(U2884) );
  INV_X1 U6221 ( .A(n5043), .ZN(n5046) );
  INV_X1 U6222 ( .A(n4651), .ZN(n5045) );
  AOI21_X1 U6223 ( .B1(n5046), .B2(n5045), .A(n5044), .ZN(n6180) );
  INV_X1 U6224 ( .A(n6180), .ZN(n5049) );
  INV_X1 U6225 ( .A(DATAI_6_), .ZN(n5047) );
  OAI222_X1 U6226 ( .A1(n5049), .A2(n5935), .B1(n5668), .B2(n5048), .C1(n5452), 
        .C2(n5047), .ZN(U2885) );
  INV_X1 U6227 ( .A(n6137), .ZN(n5053) );
  AOI21_X1 U6228 ( .B1(n6298), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n5050), 
        .ZN(n5051) );
  OAI21_X1 U6229 ( .B1(n5955), .B2(n6133), .A(n5051), .ZN(n5052) );
  AOI21_X1 U6230 ( .B1(n6288), .B2(n5053), .A(n5052), .ZN(n5054) );
  OAI21_X1 U6231 ( .B1(n6016), .B2(n5055), .A(n5054), .ZN(U2983) );
  INV_X1 U6232 ( .A(n5056), .ZN(n5062) );
  INV_X1 U6233 ( .A(n6123), .ZN(n5060) );
  AOI21_X1 U6234 ( .B1(n6298), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n5057), 
        .ZN(n5058) );
  OAI21_X1 U6235 ( .B1(n5955), .B2(n6122), .A(n5058), .ZN(n5059) );
  AOI21_X1 U6236 ( .B1(n6288), .B2(n5060), .A(n5059), .ZN(n5061) );
  OAI21_X1 U6237 ( .B1(n5062), .B2(n6016), .A(n5061), .ZN(U2982) );
  INV_X1 U6238 ( .A(n5217), .ZN(n5063) );
  OR2_X1 U6239 ( .A1(n6463), .A2(n5063), .ZN(n5068) );
  NAND2_X1 U6240 ( .A1(n5065), .A2(n5064), .ZN(n6461) );
  INV_X1 U6241 ( .A(n6461), .ZN(n5066) );
  NAND2_X1 U6242 ( .A1(n5066), .A2(n6468), .ZN(n5067) );
  NAND3_X1 U6243 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6575), .ZN(n5222) );
  NOR2_X1 U6244 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5222), .ZN(n5112)
         );
  NOR2_X2 U6245 ( .A1(n5071), .A2(n5209), .ZN(n5248) );
  AOI21_X1 U6246 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6461), .A(n5123), .ZN(
        n6472) );
  INV_X1 U6247 ( .A(n5112), .ZN(n5076) );
  INV_X1 U6248 ( .A(n5248), .ZN(n5072) );
  AOI21_X1 U6249 ( .B1(n5072), .B2(n6569), .A(n6015), .ZN(n5073) );
  AOI211_X1 U6250 ( .C1(n5217), .C2(n6391), .A(n5073), .B(n6352), .ZN(n5074)
         );
  AOI211_X1 U6251 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5076), .A(n5075), .B(
        n5074), .ZN(n5077) );
  NAND2_X1 U6252 ( .A1(n6472), .A2(n5077), .ZN(n5087) );
  AOI22_X1 U6253 ( .A1(n5248), .A2(n6553), .B1(INSTQUEUE_REG_12__6__SCAN_IN), 
        .B2(n5087), .ZN(n5078) );
  OAI21_X1 U6254 ( .B1(n6569), .B2(n6559), .A(n5078), .ZN(n5079) );
  AOI21_X1 U6255 ( .B1(n6554), .B2(n5112), .A(n5079), .ZN(n5080) );
  OAI21_X1 U6256 ( .B1(n5398), .B2(n5115), .A(n5080), .ZN(U3122) );
  INV_X1 U6257 ( .A(n5302), .ZN(n5084) );
  AOI22_X1 U6258 ( .A1(n6298), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6284), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5081) );
  OAI21_X1 U6259 ( .B1(n5955), .B2(n5082), .A(n5081), .ZN(n5083) );
  AOI21_X1 U6260 ( .B1(n5084), .B2(n6288), .A(n5083), .ZN(n5085) );
  OAI21_X1 U6261 ( .B1(n5086), .B2(n6016), .A(n5085), .ZN(U2976) );
  NAND2_X1 U6262 ( .A1(n6504), .A2(n5112), .ZN(n5091) );
  INV_X1 U6263 ( .A(n6521), .ZN(n6474) );
  INV_X1 U6264 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5088) );
  OAI22_X1 U6265 ( .A1(n5115), .A2(n5375), .B1(n5088), .B2(n5113), .ZN(n5089)
         );
  AOI21_X1 U6266 ( .B1(n5248), .B2(n6474), .A(n5089), .ZN(n5090) );
  OAI211_X1 U6267 ( .C1(n6569), .C2(n6477), .A(n5091), .B(n5090), .ZN(U3116)
         );
  NAND2_X1 U6268 ( .A1(n6535), .A2(n5112), .ZN(n5095) );
  INV_X1 U6269 ( .A(n6407), .ZN(n6534) );
  INV_X1 U6270 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5092) );
  OAI22_X1 U6271 ( .A1(n5115), .A2(n5352), .B1(n5092), .B2(n5113), .ZN(n5093)
         );
  AOI21_X1 U6272 ( .B1(n5248), .B2(n6534), .A(n5093), .ZN(n5094) );
  OAI211_X1 U6273 ( .C1(n6569), .C2(n6539), .A(n5095), .B(n5094), .ZN(U3119)
         );
  NAND2_X1 U6274 ( .A1(n6523), .A2(n5112), .ZN(n5099) );
  INV_X1 U6275 ( .A(n6438), .ZN(n6522) );
  INV_X1 U6276 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5096) );
  OAI22_X1 U6277 ( .A1(n5115), .A2(n5371), .B1(n5096), .B2(n5113), .ZN(n5097)
         );
  AOI21_X1 U6278 ( .B1(n5248), .B2(n6522), .A(n5097), .ZN(n5098) );
  OAI211_X1 U6279 ( .C1(n6569), .C2(n6527), .A(n5099), .B(n5098), .ZN(U3117)
         );
  NAND2_X1 U6280 ( .A1(n6547), .A2(n5112), .ZN(n5103) );
  INV_X1 U6281 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5100) );
  OAI22_X1 U6282 ( .A1(n5115), .A2(n5367), .B1(n5100), .B2(n5113), .ZN(n5101)
         );
  AOI21_X1 U6283 ( .B1(n5248), .B2(n6486), .A(n5101), .ZN(n5102) );
  OAI211_X1 U6284 ( .C1(n6569), .C2(n6489), .A(n5103), .B(n5102), .ZN(U3121)
         );
  NAND2_X1 U6285 ( .A1(n6529), .A2(n5112), .ZN(n5107) );
  INV_X1 U6286 ( .A(n6442), .ZN(n6528) );
  INV_X1 U6287 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5104) );
  OAI22_X1 U6288 ( .A1(n5115), .A2(n5363), .B1(n5104), .B2(n5113), .ZN(n5105)
         );
  AOI21_X1 U6289 ( .B1(n5248), .B2(n6528), .A(n5105), .ZN(n5106) );
  OAI211_X1 U6290 ( .C1(n6569), .C2(n6533), .A(n5107), .B(n5106), .ZN(U3118)
         );
  NAND2_X1 U6291 ( .A1(n6563), .A2(n5112), .ZN(n5111) );
  INV_X1 U6292 ( .A(n6570), .ZN(n6495) );
  INV_X1 U6293 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5108) );
  OAI22_X1 U6294 ( .A1(n5115), .A2(n5356), .B1(n5108), .B2(n5113), .ZN(n5109)
         );
  AOI21_X1 U6295 ( .B1(n5248), .B2(n6495), .A(n5109), .ZN(n5110) );
  OAI211_X1 U6296 ( .C1(n6569), .C2(n6500), .A(n5111), .B(n5110), .ZN(U3123)
         );
  NAND2_X1 U6297 ( .A1(n6541), .A2(n5112), .ZN(n5118) );
  INV_X1 U6298 ( .A(n6449), .ZN(n6540) );
  INV_X1 U6299 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5114) );
  OAI22_X1 U6300 ( .A1(n5115), .A2(n5383), .B1(n5114), .B2(n5113), .ZN(n5116)
         );
  AOI21_X1 U6301 ( .B1(n5248), .B2(n6540), .A(n5116), .ZN(n5117) );
  OAI211_X1 U6302 ( .C1(n6569), .C2(n6545), .A(n5118), .B(n5117), .ZN(U3120)
         );
  OAI21_X1 U6303 ( .B1(n5119), .B2(n6301), .A(n6393), .ZN(n5122) );
  INV_X1 U6304 ( .A(n5540), .ZN(n6507) );
  AND2_X1 U6305 ( .A1(n2977), .A2(n6507), .ZN(n5218) );
  INV_X1 U6306 ( .A(n6392), .ZN(n5121) );
  INV_X1 U6307 ( .A(n5151), .ZN(n5120) );
  AOI21_X1 U6308 ( .B1(n5218), .B2(n5121), .A(n5120), .ZN(n5125) );
  NAND2_X1 U6309 ( .A1(n5122), .A2(n5125), .ZN(n5124) );
  OAI211_X1 U6310 ( .C1(n5126), .C2(n6513), .A(n5124), .B(n6510), .ZN(n5154)
         );
  NOR2_X1 U6311 ( .A1(n5150), .A2(n6500), .ZN(n5129) );
  INV_X1 U6312 ( .A(n5125), .ZN(n5127) );
  AOI22_X1 U6313 ( .A1(n5127), .A2(n6389), .B1(n5126), .B2(
        STATE2_REG_2__SCAN_IN), .ZN(n5156) );
  OAI22_X1 U6314 ( .A1(n5149), .A2(n6570), .B1(n5156), .B2(n5356), .ZN(n5128)
         );
  AOI211_X1 U6315 ( .C1(INSTQUEUE_REG_15__7__SCAN_IN), .C2(n5154), .A(n5129), 
        .B(n5128), .ZN(n5130) );
  OAI21_X1 U6316 ( .B1(n5407), .B2(n5151), .A(n5130), .ZN(U3147) );
  NOR2_X1 U6317 ( .A1(n5150), .A2(n6533), .ZN(n5132) );
  OAI22_X1 U6318 ( .A1(n5149), .A2(n6442), .B1(n5156), .B2(n5363), .ZN(n5131)
         );
  AOI211_X1 U6319 ( .C1(INSTQUEUE_REG_15__2__SCAN_IN), .C2(n5154), .A(n5132), 
        .B(n5131), .ZN(n5133) );
  OAI21_X1 U6320 ( .B1(n5415), .B2(n5151), .A(n5133), .ZN(U3142) );
  NOR2_X1 U6321 ( .A1(n5150), .A2(n6477), .ZN(n5135) );
  OAI22_X1 U6322 ( .A1(n5149), .A2(n6521), .B1(n5156), .B2(n5375), .ZN(n5134)
         );
  AOI211_X1 U6323 ( .C1(INSTQUEUE_REG_15__0__SCAN_IN), .C2(n5154), .A(n5135), 
        .B(n5134), .ZN(n5136) );
  OAI21_X1 U6324 ( .B1(n5411), .B2(n5151), .A(n5136), .ZN(U3140) );
  NOR2_X1 U6325 ( .A1(n5150), .A2(n6489), .ZN(n5138) );
  OAI22_X1 U6326 ( .A1(n5149), .A2(n6551), .B1(n5156), .B2(n5367), .ZN(n5137)
         );
  AOI211_X1 U6327 ( .C1(INSTQUEUE_REG_15__5__SCAN_IN), .C2(n5154), .A(n5138), 
        .B(n5137), .ZN(n5139) );
  OAI21_X1 U6328 ( .B1(n5423), .B2(n5151), .A(n5139), .ZN(U3145) );
  NOR2_X1 U6329 ( .A1(n5150), .A2(n6527), .ZN(n5141) );
  OAI22_X1 U6330 ( .A1(n5149), .A2(n6438), .B1(n5156), .B2(n5371), .ZN(n5140)
         );
  AOI211_X1 U6331 ( .C1(INSTQUEUE_REG_15__1__SCAN_IN), .C2(n5154), .A(n5141), 
        .B(n5140), .ZN(n5142) );
  OAI21_X1 U6332 ( .B1(n5431), .B2(n5151), .A(n5142), .ZN(U3141) );
  NOR2_X1 U6333 ( .A1(n5150), .A2(n6539), .ZN(n5144) );
  OAI22_X1 U6334 ( .A1(n5149), .A2(n6407), .B1(n5156), .B2(n5352), .ZN(n5143)
         );
  AOI211_X1 U6335 ( .C1(INSTQUEUE_REG_15__3__SCAN_IN), .C2(n5154), .A(n5144), 
        .B(n5143), .ZN(n5145) );
  OAI21_X1 U6336 ( .B1(n5403), .B2(n5151), .A(n5145), .ZN(U3143) );
  NOR2_X1 U6337 ( .A1(n5150), .A2(n6545), .ZN(n5147) );
  OAI22_X1 U6338 ( .A1(n5149), .A2(n6449), .B1(n5156), .B2(n5383), .ZN(n5146)
         );
  AOI211_X1 U6339 ( .C1(INSTQUEUE_REG_15__4__SCAN_IN), .C2(n5154), .A(n5147), 
        .B(n5146), .ZN(n5148) );
  OAI21_X1 U6340 ( .B1(n5419), .B2(n5151), .A(n5148), .ZN(U3144) );
  OAI22_X1 U6341 ( .A1(n6559), .A2(n5150), .B1(n5149), .B2(n6415), .ZN(n5153)
         );
  NOR2_X1 U6342 ( .A1(n5256), .A2(n5151), .ZN(n5152) );
  AOI211_X1 U6343 ( .C1(INSTQUEUE_REG_15__6__SCAN_IN), .C2(n5154), .A(n5153), 
        .B(n5152), .ZN(n5155) );
  OAI21_X1 U6344 ( .B1(n5156), .B2(n5398), .A(n5155), .ZN(U3146) );
  CLKBUF_X1 U6345 ( .A(n5157), .Z(n5158) );
  OAI21_X1 U6346 ( .B1(n5160), .B2(n5159), .A(n5158), .ZN(n6077) );
  OAI222_X1 U6347 ( .A1(n6077), .A2(n5935), .B1(n5668), .B2(n5161), .C1(n5929), 
        .C2(n5452), .ZN(U2879) );
  CLKBUF_X1 U6348 ( .A(n5162), .Z(n5165) );
  CLKBUF_X1 U6349 ( .A(n5163), .Z(n5164) );
  XOR2_X1 U6350 ( .A(n5165), .B(n5164), .Z(n6324) );
  INV_X1 U6351 ( .A(n6324), .ZN(n5170) );
  INV_X1 U6352 ( .A(n5166), .ZN(n6097) );
  NAND2_X1 U6353 ( .A1(n6284), .A2(REIP_REG_7__SCAN_IN), .ZN(n6320) );
  NAND2_X1 U6354 ( .A1(n6298), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5167)
         );
  OAI211_X1 U6355 ( .C1(n5955), .C2(n6100), .A(n6320), .B(n5167), .ZN(n5168)
         );
  AOI21_X1 U6356 ( .B1(n6097), .B2(n6288), .A(n5168), .ZN(n5169) );
  OAI21_X1 U6357 ( .B1(n5170), .B2(n6016), .A(n5169), .ZN(U2979) );
  INV_X1 U6358 ( .A(n6055), .ZN(n5180) );
  NAND2_X1 U6359 ( .A1(n5171), .A2(n6727), .ZN(n5172) );
  NAND2_X1 U6360 ( .A1(n5172), .A2(n6039), .ZN(n6152) );
  INV_X1 U6361 ( .A(n6152), .ZN(n6166) );
  NOR2_X1 U6362 ( .A1(n5174), .A2(n5173), .ZN(n6162) );
  OAI21_X1 U6363 ( .B1(n6160), .B2(n6158), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5175) );
  OAI21_X1 U6364 ( .B1(n6129), .B2(n5176), .A(n5175), .ZN(n5177) );
  AOI21_X1 U6365 ( .B1(n6507), .B2(n6162), .A(n5177), .ZN(n5178) );
  OAI21_X1 U6366 ( .B1(n6302), .B2(n6166), .A(n5178), .ZN(n5179) );
  AOI21_X1 U6367 ( .B1(n5180), .B2(REIP_REG_0__SCAN_IN), .A(n5179), .ZN(n5181)
         );
  OAI21_X1 U6368 ( .B1(n6157), .B2(n5182), .A(n5181), .ZN(U2827) );
  NOR2_X1 U6369 ( .A1(n6131), .A2(n6717), .ZN(n6154) );
  INV_X1 U6370 ( .A(n6154), .ZN(n5184) );
  NAND2_X1 U6371 ( .A1(REIP_REG_3__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .ZN(
        n5183) );
  NAND2_X1 U6372 ( .A1(n6089), .A2(n6126), .ZN(n6101) );
  NOR3_X1 U6373 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5279), .A3(n6101), .ZN(n5293)
         );
  INV_X1 U6374 ( .A(n5185), .ZN(n6312) );
  OR2_X1 U6375 ( .A1(n6131), .A2(n5186), .ZN(n5187) );
  NAND2_X1 U6376 ( .A1(n4264), .A2(n5187), .ZN(n5615) );
  AOI22_X1 U6377 ( .A1(n6140), .A2(n6312), .B1(REIP_REG_9__SCAN_IN), .B2(n5615), .ZN(n5188) );
  OAI211_X1 U6378 ( .C1(n6144), .C2(n5196), .A(n5188), .B(n6309), .ZN(n5192)
         );
  INV_X1 U6379 ( .A(n5189), .ZN(n5198) );
  AOI22_X1 U6380 ( .A1(n6161), .A2(EBX_REG_9__SCAN_IN), .B1(n6160), .B2(n5198), 
        .ZN(n5190) );
  OAI21_X1 U6381 ( .B1(n5201), .B2(n6039), .A(n5190), .ZN(n5191) );
  OR3_X1 U6382 ( .A1(n5293), .A2(n5192), .A3(n5191), .ZN(U2818) );
  XNOR2_X1 U6383 ( .A(n5848), .B(n5194), .ZN(n5195) );
  XNOR2_X1 U6384 ( .A(n5193), .B(n5195), .ZN(n6314) );
  NAND2_X1 U6385 ( .A1(n6314), .A2(n6296), .ZN(n5200) );
  NAND2_X1 U6386 ( .A1(n6284), .A2(REIP_REG_9__SCAN_IN), .ZN(n6310) );
  OAI21_X1 U6387 ( .B1(n5746), .B2(n5196), .A(n6310), .ZN(n5197) );
  AOI21_X1 U6388 ( .B1(n5961), .B2(n5198), .A(n5197), .ZN(n5199) );
  OAI211_X1 U6389 ( .C1(n6301), .C2(n5201), .A(n5200), .B(n5199), .ZN(U2977)
         );
  NAND3_X1 U6390 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6582), .A3(n6575), .ZN(n6460) );
  NOR2_X1 U6391 ( .A1(n5385), .A2(n6460), .ZN(n5203) );
  INV_X1 U6392 ( .A(n5203), .ZN(n5262) );
  OAI21_X1 U6393 ( .B1(n5210), .B2(n6015), .A(n6389), .ZN(n5208) );
  INV_X1 U6394 ( .A(n6466), .ZN(n5204) );
  AOI21_X1 U6395 ( .B1(n5218), .B2(n5204), .A(n5203), .ZN(n5207) );
  INV_X1 U6396 ( .A(n5207), .ZN(n5206) );
  NAND2_X1 U6397 ( .A1(n6352), .A2(n6460), .ZN(n5205) );
  OAI211_X1 U6398 ( .C1(n5208), .C2(n5206), .A(n6510), .B(n5205), .ZN(n5258)
         );
  OAI22_X1 U6399 ( .A1(n5208), .A2(n5207), .B1(n6514), .B2(n6460), .ZN(n5257)
         );
  AOI22_X1 U6400 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5258), .B1(n6565), 
        .B2(n5257), .ZN(n5213) );
  NOR2_X2 U6401 ( .A1(n5210), .A2(n5209), .ZN(n6494) );
  AOI22_X1 U6402 ( .A1(n6494), .A2(n6560), .B1(n5259), .B2(n6495), .ZN(n5212)
         );
  OAI211_X1 U6403 ( .C1(n5407), .C2(n5262), .A(n5213), .B(n5212), .ZN(U3099)
         );
  AOI22_X1 U6404 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5258), .B1(n6548), 
        .B2(n5257), .ZN(n5215) );
  AOI22_X1 U6405 ( .A1(n6494), .A2(n6546), .B1(n5259), .B2(n6486), .ZN(n5214)
         );
  OAI211_X1 U6406 ( .C1(n5423), .C2(n5262), .A(n5215), .B(n5214), .ZN(U3097)
         );
  NOR2_X1 U6407 ( .A1(n5385), .A2(n5222), .ZN(n5216) );
  INV_X1 U6408 ( .A(n5216), .ZN(n5251) );
  AOI21_X1 U6409 ( .B1(n5218), .B2(n5217), .A(n5216), .ZN(n5224) );
  INV_X1 U6410 ( .A(n5224), .ZN(n5221) );
  NAND2_X1 U6411 ( .A1(n6389), .A2(n5219), .ZN(n5223) );
  NAND2_X1 U6412 ( .A1(n6352), .A2(n5222), .ZN(n5220) );
  OAI211_X1 U6413 ( .C1(n5221), .C2(n5223), .A(n6510), .B(n5220), .ZN(n5246)
         );
  OAI22_X1 U6414 ( .A1(n5224), .A2(n5223), .B1(n6514), .B2(n5222), .ZN(n5245)
         );
  AOI22_X1 U6415 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n5246), .B1(n6530), 
        .B2(n5245), .ZN(n5226) );
  AOI22_X1 U6416 ( .A1(n6439), .A2(n5248), .B1(n5247), .B2(n6528), .ZN(n5225)
         );
  OAI211_X1 U6417 ( .C1(n5415), .C2(n5251), .A(n5226), .B(n5225), .ZN(U3126)
         );
  AOI22_X1 U6418 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n5246), .B1(n6536), 
        .B2(n5245), .ZN(n5228) );
  AOI22_X1 U6419 ( .A1(n6404), .A2(n5248), .B1(n5247), .B2(n6534), .ZN(n5227)
         );
  OAI211_X1 U6420 ( .C1(n5403), .C2(n5251), .A(n5228), .B(n5227), .ZN(U3127)
         );
  AOI22_X1 U6421 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n5246), .B1(n6542), 
        .B2(n5245), .ZN(n5230) );
  AOI22_X1 U6422 ( .A1(n6446), .A2(n5248), .B1(n5247), .B2(n6540), .ZN(n5229)
         );
  OAI211_X1 U6423 ( .C1(n5419), .C2(n5251), .A(n5230), .B(n5229), .ZN(U3128)
         );
  AOI22_X1 U6424 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5258), .B1(n6542), 
        .B2(n5257), .ZN(n5232) );
  AOI22_X1 U6425 ( .A1(n6494), .A2(n6446), .B1(n5259), .B2(n6540), .ZN(n5231)
         );
  OAI211_X1 U6426 ( .C1(n5419), .C2(n5262), .A(n5232), .B(n5231), .ZN(U3096)
         );
  AOI22_X1 U6427 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n5246), .B1(n6555), 
        .B2(n5245), .ZN(n5234) );
  INV_X1 U6428 ( .A(n6559), .ZN(n6412) );
  AOI22_X1 U6429 ( .A1(n6412), .A2(n5248), .B1(n5247), .B2(n6553), .ZN(n5233)
         );
  OAI211_X1 U6430 ( .C1(n5256), .C2(n5251), .A(n5234), .B(n5233), .ZN(U3130)
         );
  AOI22_X1 U6431 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n5246), .B1(n6565), 
        .B2(n5245), .ZN(n5236) );
  AOI22_X1 U6432 ( .A1(n6560), .A2(n5248), .B1(n5247), .B2(n6495), .ZN(n5235)
         );
  OAI211_X1 U6433 ( .C1(n5407), .C2(n5251), .A(n5236), .B(n5235), .ZN(U3131)
         );
  AOI22_X1 U6434 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n5258), .B1(n6530), 
        .B2(n5257), .ZN(n5238) );
  AOI22_X1 U6435 ( .A1(n6494), .A2(n6439), .B1(n5259), .B2(n6528), .ZN(n5237)
         );
  OAI211_X1 U6436 ( .C1(n5415), .C2(n5262), .A(n5238), .B(n5237), .ZN(U3094)
         );
  AOI22_X1 U6437 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5258), .B1(n6536), 
        .B2(n5257), .ZN(n5240) );
  AOI22_X1 U6438 ( .A1(n6494), .A2(n6404), .B1(n5259), .B2(n6534), .ZN(n5239)
         );
  OAI211_X1 U6439 ( .C1(n5403), .C2(n5262), .A(n5240), .B(n5239), .ZN(U3095)
         );
  AOI22_X1 U6440 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n5246), .B1(n6548), 
        .B2(n5245), .ZN(n5242) );
  AOI22_X1 U6441 ( .A1(n6546), .A2(n5248), .B1(n5247), .B2(n6486), .ZN(n5241)
         );
  OAI211_X1 U6442 ( .C1(n5423), .C2(n5251), .A(n5242), .B(n5241), .ZN(U3129)
         );
  AOI22_X1 U6443 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n5246), .B1(n6518), 
        .B2(n5245), .ZN(n5244) );
  AOI22_X1 U6444 ( .A1(n6503), .A2(n5248), .B1(n5247), .B2(n6474), .ZN(n5243)
         );
  OAI211_X1 U6445 ( .C1(n5411), .C2(n5251), .A(n5244), .B(n5243), .ZN(U3124)
         );
  AOI22_X1 U6446 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n5246), .B1(n6524), 
        .B2(n5245), .ZN(n5250) );
  AOI22_X1 U6447 ( .A1(n6435), .A2(n5248), .B1(n5247), .B2(n6522), .ZN(n5249)
         );
  OAI211_X1 U6448 ( .C1(n5431), .C2(n5251), .A(n5250), .B(n5249), .ZN(U3125)
         );
  AOI22_X1 U6449 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5258), .B1(n6524), 
        .B2(n5257), .ZN(n5253) );
  AOI22_X1 U6450 ( .A1(n6494), .A2(n6435), .B1(n5259), .B2(n6522), .ZN(n5252)
         );
  OAI211_X1 U6451 ( .C1(n5431), .C2(n5262), .A(n5253), .B(n5252), .ZN(U3093)
         );
  AOI22_X1 U6452 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5258), .B1(n6555), 
        .B2(n5257), .ZN(n5255) );
  AOI22_X1 U6453 ( .A1(n6494), .A2(n6412), .B1(n5259), .B2(n6553), .ZN(n5254)
         );
  OAI211_X1 U6454 ( .C1(n5256), .C2(n5262), .A(n5255), .B(n5254), .ZN(U3098)
         );
  AOI22_X1 U6455 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5258), .B1(n6518), 
        .B2(n5257), .ZN(n5261) );
  AOI22_X1 U6456 ( .A1(n6494), .A2(n6503), .B1(n5259), .B2(n6474), .ZN(n5260)
         );
  OAI211_X1 U6457 ( .C1(n5411), .C2(n5262), .A(n5261), .B(n5260), .ZN(U3092)
         );
  CLKBUF_X1 U6458 ( .A(n5263), .Z(n5264) );
  NAND2_X1 U6459 ( .A1(n5266), .A2(n5265), .ZN(n5267) );
  XNOR2_X1 U6460 ( .A(n5264), .B(n5267), .ZN(n6304) );
  INV_X1 U6461 ( .A(n6304), .ZN(n5272) );
  AOI22_X1 U6462 ( .A1(n6298), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .B1(n6284), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n5268) );
  OAI21_X1 U6463 ( .B1(n5955), .B2(n5277), .A(n5268), .ZN(n5269) );
  AOI21_X1 U6464 ( .B1(n5270), .B2(n6288), .A(n5269), .ZN(n5271) );
  OAI21_X1 U6465 ( .B1(n5272), .B2(n6016), .A(n5271), .ZN(U2975) );
  INV_X1 U6466 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5274) );
  OAI22_X1 U6467 ( .A1(n5274), .A2(n6129), .B1(n5273), .B2(n6144), .ZN(n5275)
         );
  INV_X1 U6468 ( .A(n5275), .ZN(n5276) );
  OAI21_X1 U6469 ( .B1(n5277), .B2(n6146), .A(n5276), .ZN(n5278) );
  AOI211_X1 U6470 ( .C1(n6140), .C2(n6303), .A(n6328), .B(n5278), .ZN(n5283)
         );
  INV_X1 U6471 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6668) );
  INV_X1 U6472 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6664) );
  NOR3_X1 U6473 ( .A1(n6664), .A2(n5279), .A3(n6101), .ZN(n5295) );
  NAND2_X1 U6474 ( .A1(REIP_REG_10__SCAN_IN), .A2(n5295), .ZN(n6073) );
  NAND2_X1 U6475 ( .A1(n6668), .A2(n6073), .ZN(n5281) );
  OAI21_X1 U6476 ( .B1(n5280), .B2(n6131), .A(n4264), .ZN(n6079) );
  NAND2_X1 U6477 ( .A1(n5281), .A2(n6079), .ZN(n5282) );
  OAI211_X1 U6478 ( .C1(n5284), .C2(n6039), .A(n5283), .B(n5282), .ZN(U2816)
         );
  NAND2_X1 U6479 ( .A1(n5158), .A2(n5286), .ZN(n5287) );
  AND2_X1 U6480 ( .A1(n5285), .A2(n5287), .ZN(n6072) );
  INV_X1 U6481 ( .A(n6072), .ZN(n5292) );
  AOI22_X1 U6482 ( .A1(EAX_REG_13__SCAN_IN), .A2(n6193), .B1(n5340), .B2(
        DATAI_13_), .ZN(n5288) );
  OAI21_X1 U6483 ( .B1(n5292), .B2(n5935), .A(n5288), .ZN(U2878) );
  AOI21_X1 U6484 ( .B1(n5326), .B2(n5327), .A(n5289), .ZN(n5290) );
  NOR2_X1 U6485 ( .A1(n5290), .A2(n5433), .ZN(n6066) );
  AOI22_X1 U6486 ( .A1(n6178), .A2(n6066), .B1(n5641), .B2(EBX_REG_13__SCAN_IN), .ZN(n5291) );
  OAI21_X1 U6487 ( .B1(n5292), .B2(n5667), .A(n5291), .ZN(U2846) );
  OR3_X1 U6488 ( .A1(n5293), .A2(n6662), .A3(n5615), .ZN(n5294) );
  OAI21_X1 U6489 ( .B1(n5295), .B2(REIP_REG_10__SCAN_IN), .A(n5294), .ZN(n5301) );
  AOI22_X1 U6490 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6161), .B1(n5296), .B2(n6160), .ZN(n5297) );
  OAI21_X1 U6491 ( .B1(n6157), .B2(n5298), .A(n5297), .ZN(n5299) );
  AOI211_X1 U6492 ( .C1(n6158), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6328), 
        .B(n5299), .ZN(n5300) );
  OAI211_X1 U6493 ( .C1(n5302), .C2(n6039), .A(n5301), .B(n5300), .ZN(U2817)
         );
  AOI21_X1 U6494 ( .B1(n6298), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n5303), 
        .ZN(n5304) );
  OAI21_X1 U6495 ( .B1(n5955), .B2(n6117), .A(n5304), .ZN(n5305) );
  AOI21_X1 U6496 ( .B1(n6113), .B2(n6288), .A(n5305), .ZN(n5306) );
  OAI21_X1 U6497 ( .B1(n6016), .B2(n5307), .A(n5306), .ZN(U2981) );
  AOI22_X1 U6498 ( .A1(n6298), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .B1(n6284), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n5308) );
  OAI21_X1 U6499 ( .B1(n5955), .B2(n6105), .A(n5308), .ZN(n5309) );
  AOI21_X1 U6500 ( .B1(n6180), .B2(n6288), .A(n5309), .ZN(n5310) );
  OAI21_X1 U6501 ( .B1(n6016), .B2(n5311), .A(n5310), .ZN(U2980) );
  NAND2_X1 U6502 ( .A1(n6298), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5312)
         );
  OAI211_X1 U6503 ( .C1(n5955), .C2(n5314), .A(n5313), .B(n5312), .ZN(n5315)
         );
  AOI21_X1 U6504 ( .B1(n5614), .B2(n6288), .A(n5315), .ZN(n5316) );
  OAI21_X1 U6505 ( .B1(n6016), .B2(n5317), .A(n5316), .ZN(U2978) );
  CLKBUF_X1 U6506 ( .A(n5318), .Z(n5319) );
  XNOR2_X1 U6507 ( .A(n5848), .B(n5320), .ZN(n5321) );
  XNOR2_X1 U6508 ( .A(n5319), .B(n5321), .ZN(n5333) );
  INV_X1 U6509 ( .A(n6306), .ZN(n5984) );
  NOR3_X1 U6510 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n5984), .A3(n5322), 
        .ZN(n5331) );
  INV_X1 U6511 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6666) );
  INV_X1 U6512 ( .A(n5976), .ZN(n5323) );
  NAND2_X1 U6513 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n5323), .ZN(n6305) );
  OAI211_X1 U6514 ( .C1(n5325), .C2(n5324), .A(INSTADDRPOINTER_REG_12__SCAN_IN), .B(n6305), .ZN(n5329) );
  XOR2_X1 U6515 ( .A(n5327), .B(n5326), .Z(n6173) );
  NAND2_X1 U6516 ( .A1(n6330), .A2(n6173), .ZN(n5328) );
  OAI211_X1 U6517 ( .C1(n6666), .C2(n6309), .A(n5329), .B(n5328), .ZN(n5330)
         );
  AOI211_X1 U6518 ( .C1(n5333), .C2(n6336), .A(n5331), .B(n5330), .ZN(n5332)
         );
  INV_X1 U6519 ( .A(n5332), .ZN(U3006) );
  NAND2_X1 U6520 ( .A1(n5333), .A2(n6296), .ZN(n5336) );
  OAI22_X1 U6521 ( .A1(n5746), .A2(n6081), .B1(n6309), .B2(n6666), .ZN(n5334)
         );
  AOI21_X1 U6522 ( .B1(n6078), .B2(n5961), .A(n5334), .ZN(n5335) );
  OAI211_X1 U6523 ( .C1(n6301), .C2(n6077), .A(n5336), .B(n5335), .ZN(U2974)
         );
  AOI21_X1 U6524 ( .B1(n5339), .B2(n5285), .A(n5338), .ZN(n6062) );
  INV_X1 U6525 ( .A(n6062), .ZN(n5436) );
  AOI22_X1 U6526 ( .A1(EAX_REG_14__SCAN_IN), .A2(n6193), .B1(n5340), .B2(
        DATAI_14_), .ZN(n5341) );
  OAI21_X1 U6527 ( .B1(n5436), .B2(n5935), .A(n5341), .ZN(U2877) );
  NOR2_X1 U6528 ( .A1(n5385), .A2(n5345), .ZN(n5381) );
  AOI21_X1 U6529 ( .B1(n5342), .B2(n6507), .A(n5381), .ZN(n5347) );
  OAI22_X1 U6530 ( .A1(n5344), .A2(n5347), .B1(n5345), .B2(n6514), .ZN(n5343)
         );
  INV_X1 U6531 ( .A(n5344), .ZN(n5346) );
  AOI22_X1 U6532 ( .A1(n5347), .A2(n5346), .B1(n5345), .B2(n6352), .ZN(n5348)
         );
  NAND2_X1 U6533 ( .A1(n6510), .A2(n5348), .ZN(n5376) );
  AOI22_X1 U6534 ( .A1(n5377), .A2(n6534), .B1(INSTQUEUE_REG_1__3__SCAN_IN), 
        .B2(n5376), .ZN(n5349) );
  OAI21_X1 U6535 ( .B1(n6539), .B2(n5379), .A(n5349), .ZN(n5350) );
  AOI21_X1 U6536 ( .B1(n6535), .B2(n5381), .A(n5350), .ZN(n5351) );
  OAI21_X1 U6537 ( .B1(n5384), .B2(n5352), .A(n5351), .ZN(U3031) );
  AOI22_X1 U6538 ( .A1(n5377), .A2(n6495), .B1(INSTQUEUE_REG_1__7__SCAN_IN), 
        .B2(n5376), .ZN(n5353) );
  OAI21_X1 U6539 ( .B1(n6500), .B2(n5379), .A(n5353), .ZN(n5354) );
  AOI21_X1 U6540 ( .B1(n6563), .B2(n5381), .A(n5354), .ZN(n5355) );
  OAI21_X1 U6541 ( .B1(n5384), .B2(n5356), .A(n5355), .ZN(U3035) );
  AOI22_X1 U6542 ( .A1(n5377), .A2(n6553), .B1(INSTQUEUE_REG_1__6__SCAN_IN), 
        .B2(n5376), .ZN(n5357) );
  OAI21_X1 U6543 ( .B1(n6559), .B2(n5379), .A(n5357), .ZN(n5358) );
  AOI21_X1 U6544 ( .B1(n6554), .B2(n5381), .A(n5358), .ZN(n5359) );
  OAI21_X1 U6545 ( .B1(n5398), .B2(n5384), .A(n5359), .ZN(U3034) );
  AOI22_X1 U6546 ( .A1(n5377), .A2(n6528), .B1(INSTQUEUE_REG_1__2__SCAN_IN), 
        .B2(n5376), .ZN(n5360) );
  OAI21_X1 U6547 ( .B1(n6533), .B2(n5379), .A(n5360), .ZN(n5361) );
  AOI21_X1 U6548 ( .B1(n6529), .B2(n5381), .A(n5361), .ZN(n5362) );
  OAI21_X1 U6549 ( .B1(n5384), .B2(n5363), .A(n5362), .ZN(U3030) );
  AOI22_X1 U6550 ( .A1(n5377), .A2(n6486), .B1(INSTQUEUE_REG_1__5__SCAN_IN), 
        .B2(n5376), .ZN(n5364) );
  OAI21_X1 U6551 ( .B1(n6489), .B2(n5379), .A(n5364), .ZN(n5365) );
  AOI21_X1 U6552 ( .B1(n6547), .B2(n5381), .A(n5365), .ZN(n5366) );
  OAI21_X1 U6553 ( .B1(n5384), .B2(n5367), .A(n5366), .ZN(U3033) );
  AOI22_X1 U6554 ( .A1(n5377), .A2(n6522), .B1(INSTQUEUE_REG_1__1__SCAN_IN), 
        .B2(n5376), .ZN(n5368) );
  OAI21_X1 U6555 ( .B1(n6527), .B2(n5379), .A(n5368), .ZN(n5369) );
  AOI21_X1 U6556 ( .B1(n6523), .B2(n5381), .A(n5369), .ZN(n5370) );
  OAI21_X1 U6557 ( .B1(n5384), .B2(n5371), .A(n5370), .ZN(U3029) );
  AOI22_X1 U6558 ( .A1(n5377), .A2(n6474), .B1(INSTQUEUE_REG_1__0__SCAN_IN), 
        .B2(n5376), .ZN(n5372) );
  OAI21_X1 U6559 ( .B1(n6477), .B2(n5379), .A(n5372), .ZN(n5373) );
  AOI21_X1 U6560 ( .B1(n6504), .B2(n5381), .A(n5373), .ZN(n5374) );
  OAI21_X1 U6561 ( .B1(n5384), .B2(n5375), .A(n5374), .ZN(U3028) );
  AOI22_X1 U6562 ( .A1(n5377), .A2(n6540), .B1(INSTQUEUE_REG_1__4__SCAN_IN), 
        .B2(n5376), .ZN(n5378) );
  OAI21_X1 U6563 ( .B1(n6545), .B2(n5379), .A(n5378), .ZN(n5380) );
  AOI21_X1 U6564 ( .B1(n6541), .B2(n5381), .A(n5380), .ZN(n5382) );
  OAI21_X1 U6565 ( .B1(n5384), .B2(n5383), .A(n5382), .ZN(U3032) );
  NOR2_X1 U6566 ( .A1(n5385), .A2(n5390), .ZN(n5399) );
  AOI21_X1 U6567 ( .B1(n5386), .B2(n6507), .A(n5399), .ZN(n5392) );
  OAI22_X1 U6568 ( .A1(n5389), .A2(n5392), .B1(n5390), .B2(n6514), .ZN(n5428)
         );
  INV_X1 U6569 ( .A(n5428), .ZN(n5397) );
  NOR2_X1 U6570 ( .A1(n4702), .A2(n5387), .ZN(n5388) );
  INV_X1 U6571 ( .A(n5389), .ZN(n5391) );
  AOI22_X1 U6572 ( .A1(n5392), .A2(n5391), .B1(n5390), .B2(n6352), .ZN(n5393)
         );
  NAND2_X1 U6573 ( .A1(n6510), .A2(n5393), .ZN(n5424) );
  AOI22_X1 U6574 ( .A1(n6418), .A2(n6553), .B1(INSTQUEUE_REG_5__6__SCAN_IN), 
        .B2(n5424), .ZN(n5394) );
  OAI21_X1 U6575 ( .B1(n5426), .B2(n6559), .A(n5394), .ZN(n5395) );
  AOI21_X1 U6576 ( .B1(n6554), .B2(n5399), .A(n5395), .ZN(n5396) );
  OAI21_X1 U6577 ( .B1(n5398), .B2(n5397), .A(n5396), .ZN(U3066) );
  INV_X1 U6578 ( .A(n5399), .ZN(n5430) );
  AOI22_X1 U6579 ( .A1(n6418), .A2(n6534), .B1(INSTQUEUE_REG_5__3__SCAN_IN), 
        .B2(n5424), .ZN(n5400) );
  OAI21_X1 U6580 ( .B1(n5426), .B2(n6539), .A(n5400), .ZN(n5401) );
  AOI21_X1 U6581 ( .B1(n6536), .B2(n5428), .A(n5401), .ZN(n5402) );
  OAI21_X1 U6582 ( .B1(n5403), .B2(n5430), .A(n5402), .ZN(U3063) );
  AOI22_X1 U6583 ( .A1(n6418), .A2(n6495), .B1(INSTQUEUE_REG_5__7__SCAN_IN), 
        .B2(n5424), .ZN(n5404) );
  OAI21_X1 U6584 ( .B1(n5426), .B2(n6500), .A(n5404), .ZN(n5405) );
  AOI21_X1 U6585 ( .B1(n6565), .B2(n5428), .A(n5405), .ZN(n5406) );
  OAI21_X1 U6586 ( .B1(n5407), .B2(n5430), .A(n5406), .ZN(U3067) );
  AOI22_X1 U6587 ( .A1(n6418), .A2(n6474), .B1(INSTQUEUE_REG_5__0__SCAN_IN), 
        .B2(n5424), .ZN(n5408) );
  OAI21_X1 U6588 ( .B1(n5426), .B2(n6477), .A(n5408), .ZN(n5409) );
  AOI21_X1 U6589 ( .B1(n6518), .B2(n5428), .A(n5409), .ZN(n5410) );
  OAI21_X1 U6590 ( .B1(n5411), .B2(n5430), .A(n5410), .ZN(U3060) );
  AOI22_X1 U6591 ( .A1(n6418), .A2(n6528), .B1(INSTQUEUE_REG_5__2__SCAN_IN), 
        .B2(n5424), .ZN(n5412) );
  OAI21_X1 U6592 ( .B1(n5426), .B2(n6533), .A(n5412), .ZN(n5413) );
  AOI21_X1 U6593 ( .B1(n6530), .B2(n5428), .A(n5413), .ZN(n5414) );
  OAI21_X1 U6594 ( .B1(n5415), .B2(n5430), .A(n5414), .ZN(U3062) );
  AOI22_X1 U6595 ( .A1(n6418), .A2(n6540), .B1(INSTQUEUE_REG_5__4__SCAN_IN), 
        .B2(n5424), .ZN(n5416) );
  OAI21_X1 U6596 ( .B1(n5426), .B2(n6545), .A(n5416), .ZN(n5417) );
  AOI21_X1 U6597 ( .B1(n6542), .B2(n5428), .A(n5417), .ZN(n5418) );
  OAI21_X1 U6598 ( .B1(n5419), .B2(n5430), .A(n5418), .ZN(U3064) );
  AOI22_X1 U6599 ( .A1(n6418), .A2(n6486), .B1(INSTQUEUE_REG_5__5__SCAN_IN), 
        .B2(n5424), .ZN(n5420) );
  OAI21_X1 U6600 ( .B1(n5426), .B2(n6489), .A(n5420), .ZN(n5421) );
  AOI21_X1 U6601 ( .B1(n6548), .B2(n5428), .A(n5421), .ZN(n5422) );
  OAI21_X1 U6602 ( .B1(n5423), .B2(n5430), .A(n5422), .ZN(U3065) );
  AOI22_X1 U6603 ( .A1(n6418), .A2(n6522), .B1(INSTQUEUE_REG_5__1__SCAN_IN), 
        .B2(n5424), .ZN(n5425) );
  OAI21_X1 U6604 ( .B1(n5426), .B2(n6527), .A(n5425), .ZN(n5427) );
  AOI21_X1 U6605 ( .B1(n6524), .B2(n5428), .A(n5427), .ZN(n5429) );
  OAI21_X1 U6606 ( .B1(n5431), .B2(n5430), .A(n5429), .ZN(U3061) );
  INV_X1 U6607 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5435) );
  OR2_X1 U6608 ( .A1(n5433), .A2(n5432), .ZN(n5434) );
  NAND2_X1 U6609 ( .A1(n5442), .A2(n5434), .ZN(n6065) );
  OAI222_X1 U6610 ( .A1(n5436), .A2(n5667), .B1(n6182), .B2(n5435), .C1(n6065), 
        .C2(n5666), .ZN(U2845) );
  AOI21_X1 U6611 ( .B1(n5439), .B2(n5438), .A(n5437), .ZN(n5508) );
  INV_X1 U6612 ( .A(n5508), .ZN(n5453) );
  INV_X1 U6613 ( .A(n5481), .ZN(n5441) );
  AOI21_X1 U6614 ( .B1(n5443), .B2(n5442), .A(n5441), .ZN(n5989) );
  AOI22_X1 U6615 ( .A1(n5989), .A2(n6178), .B1(n5641), .B2(EBX_REG_15__SCAN_IN), .ZN(n5444) );
  OAI21_X1 U6616 ( .B1(n5453), .B2(n5667), .A(n5444), .ZN(U2844) );
  INV_X1 U6617 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5446) );
  AOI21_X1 U6618 ( .B1(REIP_REG_15__SCAN_IN), .B2(n6054), .A(n6055), .ZN(n6046) );
  OAI21_X1 U6619 ( .B1(n6045), .B2(REIP_REG_15__SCAN_IN), .A(n6046), .ZN(n5445) );
  OAI211_X1 U6620 ( .C1(n6129), .C2(n5446), .A(n6309), .B(n5445), .ZN(n5447)
         );
  AOI21_X1 U6621 ( .B1(PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n6158), .A(n5447), 
        .ZN(n5450) );
  INV_X1 U6622 ( .A(n5506), .ZN(n5448) );
  AOI22_X1 U6623 ( .A1(n6140), .A2(n5989), .B1(n5448), .B2(n6160), .ZN(n5449)
         );
  OAI211_X1 U6624 ( .C1(n5453), .C2(n6039), .A(n5450), .B(n5449), .ZN(U2812)
         );
  INV_X1 U6625 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6205) );
  OAI222_X1 U6626 ( .A1(n5453), .A2(n5935), .B1(n5452), .B2(n5451), .C1(n5668), 
        .C2(n6205), .ZN(U2876) );
  INV_X1 U6627 ( .A(n5455), .ZN(n5456) );
  AOI21_X1 U6628 ( .B1(n5458), .B2(n5457), .A(n5456), .ZN(n5470) );
  NOR2_X1 U6629 ( .A1(n6309), .A2(n6670), .ZN(n5467) );
  AOI21_X1 U6630 ( .B1(n6298), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5467), 
        .ZN(n5459) );
  OAI21_X1 U6631 ( .B1(n5955), .B2(n6076), .A(n5459), .ZN(n5460) );
  AOI21_X1 U6632 ( .B1(n6072), .B2(n6288), .A(n5460), .ZN(n5461) );
  OAI21_X1 U6633 ( .B1(n5470), .B2(n6016), .A(n5461), .ZN(U2973) );
  AOI21_X1 U6634 ( .B1(n5462), .B2(n5465), .A(n5976), .ZN(n5463) );
  OAI21_X1 U6635 ( .B1(n6003), .B2(n5464), .A(n5463), .ZN(n6000) );
  NOR2_X1 U6636 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5465), .ZN(n5466)
         );
  AOI22_X1 U6637 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6000), .B1(n5466), .B2(n6306), .ZN(n5469) );
  AOI21_X1 U6638 ( .B1(n6330), .B2(n6066), .A(n5467), .ZN(n5468) );
  OAI211_X1 U6639 ( .C1(n5470), .C2(n5997), .A(n5469), .B(n5468), .ZN(U3005)
         );
  XNOR2_X1 U6640 ( .A(n5848), .B(n6002), .ZN(n5473) );
  XNOR2_X1 U6641 ( .A(n5472), .B(n5473), .ZN(n5998) );
  AOI22_X1 U6642 ( .A1(n6298), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6284), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5474) );
  OAI21_X1 U6643 ( .B1(n5955), .B2(n5475), .A(n5474), .ZN(n5476) );
  AOI21_X1 U6644 ( .B1(n6062), .B2(n6288), .A(n5476), .ZN(n5477) );
  OAI21_X1 U6645 ( .B1(n5998), .B2(n6016), .A(n5477), .ZN(U2972) );
  NOR2_X1 U6646 ( .A1(n5437), .A2(n5479), .ZN(n5480) );
  OR2_X1 U6647 ( .A1(n5478), .A2(n5480), .ZN(n5758) );
  INV_X1 U6648 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5484) );
  AOI21_X1 U6649 ( .B1(n5482), .B2(n5481), .A(n2991), .ZN(n5483) );
  INV_X1 U6650 ( .A(n5483), .ZN(n6053) );
  OAI222_X1 U6651 ( .A1(n5758), .A2(n5667), .B1(n6182), .B2(n5484), .C1(n6053), 
        .C2(n5666), .ZN(U2843) );
  OR2_X1 U6652 ( .A1(n5478), .A2(n5486), .ZN(n5487) );
  AND2_X1 U6653 ( .A1(n5485), .A2(n5487), .ZN(n6187) );
  INV_X1 U6654 ( .A(n6187), .ZN(n5511) );
  NAND2_X1 U6655 ( .A1(n5489), .A2(n5488), .ZN(n5493) );
  INV_X1 U6656 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5491) );
  OAI22_X1 U6657 ( .A1(n5491), .A2(n6129), .B1(n5490), .B2(n6144), .ZN(n5492)
         );
  AOI211_X1 U6658 ( .C1(n6035), .C2(n5493), .A(n6328), .B(n5492), .ZN(n5498)
         );
  OR2_X1 U6659 ( .A1(n2991), .A2(n5494), .ZN(n5495) );
  NAND2_X1 U6660 ( .A1(n5525), .A2(n5495), .ZN(n5855) );
  INV_X1 U6661 ( .A(n5855), .ZN(n5496) );
  AOI22_X1 U6662 ( .A1(n6140), .A2(n5496), .B1(n6160), .B2(n5960), .ZN(n5497)
         );
  OAI211_X1 U6663 ( .C1(n5511), .C2(n6039), .A(n5498), .B(n5497), .ZN(U2810)
         );
  INV_X1 U6664 ( .A(n5501), .ZN(n5503) );
  NOR2_X1 U6665 ( .A1(n5503), .A2(n5502), .ZN(n5504) );
  XNOR2_X1 U6666 ( .A(n5500), .B(n5504), .ZN(n5990) );
  INV_X1 U6667 ( .A(n5990), .ZN(n5510) );
  AOI22_X1 U6668 ( .A1(n6298), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n6284), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5505) );
  OAI21_X1 U6669 ( .B1(n5955), .B2(n5506), .A(n5505), .ZN(n5507) );
  AOI21_X1 U6670 ( .B1(n5508), .B2(n6288), .A(n5507), .ZN(n5509) );
  OAI21_X1 U6671 ( .B1(n5510), .B2(n6016), .A(n5509), .ZN(U2971) );
  OAI222_X1 U6672 ( .A1(n5855), .A2(n5666), .B1(n5491), .B2(n6182), .C1(n5511), 
        .C2(n5667), .ZN(U2842) );
  NAND2_X1 U6673 ( .A1(n5485), .A2(n5513), .ZN(n5514) );
  AND2_X1 U6674 ( .A1(n5512), .A2(n5514), .ZN(n6184) );
  INV_X1 U6675 ( .A(n6184), .ZN(n6040) );
  INV_X1 U6676 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5518) );
  XNOR2_X1 U6677 ( .A(n5516), .B(n5515), .ZN(n5524) );
  INV_X1 U6678 ( .A(n5524), .ZN(n5517) );
  XNOR2_X1 U6679 ( .A(n5525), .B(n5517), .ZN(n5846) );
  INV_X1 U6680 ( .A(n5846), .ZN(n6038) );
  OAI222_X1 U6681 ( .A1(n5667), .A2(n6040), .B1(n6182), .B2(n5518), .C1(n5666), 
        .C2(n6038), .ZN(U2841) );
  INV_X1 U6682 ( .A(n5519), .ZN(n5520) );
  AOI21_X1 U6683 ( .B1(n5512), .B2(n5521), .A(n5520), .ZN(n5748) );
  OR2_X1 U6684 ( .A1(n5661), .A2(n5524), .ZN(n5527) );
  OAI21_X1 U6685 ( .B1(n5525), .B2(n5524), .A(n5523), .ZN(n5526) );
  NAND2_X1 U6686 ( .A1(n5527), .A2(n5526), .ZN(n5920) );
  OAI22_X1 U6687 ( .A1(n5920), .A2(n5666), .B1(n5528), .B2(n6182), .ZN(n5529)
         );
  AOI21_X1 U6688 ( .B1(n5748), .B2(n6179), .A(n5529), .ZN(n5530) );
  INV_X1 U6689 ( .A(n5530), .ZN(U2840) );
  INV_X1 U6690 ( .A(n5748), .ZN(n5921) );
  INV_X1 U6691 ( .A(n5531), .ZN(n5532) );
  NOR2_X2 U6692 ( .A1(n5532), .A2(n3282), .ZN(n6194) );
  AOI22_X1 U6693 ( .A1(n6194), .A2(DATAI_19_), .B1(n6193), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5536) );
  AND2_X1 U6694 ( .A1(n3281), .A2(n5533), .ZN(n5534) );
  NAND2_X1 U6695 ( .A1(n6190), .A2(DATAI_3_), .ZN(n5535) );
  OAI211_X1 U6696 ( .C1(n5921), .C2(n5935), .A(n5536), .B(n5535), .ZN(U2872)
         );
  AOI21_X1 U6697 ( .B1(n5537), .B2(n6611), .A(n5869), .ZN(n5547) );
  INV_X1 U6698 ( .A(n5538), .ZN(n5539) );
  OR2_X1 U6699 ( .A1(n5540), .A2(n5539), .ZN(n5543) );
  NAND2_X1 U6700 ( .A1(n5541), .A2(n3078), .ZN(n5542) );
  AND2_X1 U6701 ( .A1(n5543), .A2(n5542), .ZN(n6571) );
  OAI21_X1 U6702 ( .B1(n6571), .B2(STATE2_REG_3__SCAN_IN), .A(n6614), .ZN(
        n5545) );
  INV_X1 U6703 ( .A(n5544), .ZN(n5561) );
  AOI22_X1 U6704 ( .A1(n5545), .A2(n5561), .B1(n5562), .B2(n3078), .ZN(n5546)
         );
  OAI22_X1 U6705 ( .A1(n5547), .A2(n3078), .B1(n5869), .B2(n5546), .ZN(U3461)
         );
  OAI22_X1 U6706 ( .A1(n5780), .A2(n5666), .B1(n5549), .B2(n6182), .ZN(n5550)
         );
  INV_X1 U6707 ( .A(n5550), .ZN(n5551) );
  OAI21_X1 U6708 ( .B1(n5548), .B2(n5667), .A(n5551), .ZN(U2834) );
  AOI22_X1 U6709 ( .A1(n6194), .A2(DATAI_25_), .B1(n6193), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5553) );
  NAND2_X1 U6710 ( .A1(n6190), .A2(DATAI_9_), .ZN(n5552) );
  OAI211_X1 U6711 ( .C1(n5548), .C2(n5935), .A(n5553), .B(n5552), .ZN(U2866)
         );
  AOI21_X1 U6712 ( .B1(n6298), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5554), 
        .ZN(n5555) );
  OAI21_X1 U6713 ( .B1(n5955), .B2(n5556), .A(n5555), .ZN(n5557) );
  AOI21_X1 U6714 ( .B1(n5670), .B2(n6288), .A(n5557), .ZN(n5558) );
  OAI21_X1 U6715 ( .B1(n5559), .B2(n6016), .A(n5558), .ZN(U2955) );
  AOI21_X1 U6716 ( .B1(n5562), .B2(n5563), .A(n5869), .ZN(n5568) );
  NOR2_X1 U6717 ( .A1(n5561), .A2(n5560), .ZN(n5565) );
  INV_X1 U6718 ( .A(n5562), .ZN(n6604) );
  NOR3_X1 U6719 ( .A1(n5563), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n6604), 
        .ZN(n5564) );
  AOI211_X1 U6720 ( .C1(n5566), .C2(n6611), .A(n5565), .B(n5564), .ZN(n5567)
         );
  OAI22_X1 U6721 ( .A1(n5568), .A2(n3099), .B1(n5869), .B2(n5567), .ZN(U3459)
         );
  INV_X1 U6722 ( .A(n5687), .ZN(n5675) );
  OAI211_X1 U6723 ( .C1(REIP_REG_30__SCAN_IN), .C2(REIP_REG_29__SCAN_IN), .A(
        n5585), .B(n5569), .ZN(n5577) );
  INV_X1 U6724 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5572) );
  INV_X1 U6725 ( .A(n5685), .ZN(n5570) );
  AOI22_X1 U6726 ( .A1(n6160), .A2(n5570), .B1(PHYADDRPOINTER_REG_30__SCAN_IN), 
        .B2(n6158), .ZN(n5571) );
  OAI21_X1 U6727 ( .B1(n6129), .B2(n5572), .A(n5571), .ZN(n5574) );
  INV_X1 U6728 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6703) );
  NOR2_X1 U6729 ( .A1(n5582), .A2(n6703), .ZN(n5573) );
  AOI211_X1 U6730 ( .C1(n6140), .C2(n5575), .A(n5574), .B(n5573), .ZN(n5576)
         );
  OAI211_X1 U6731 ( .C1(n5675), .C2(n6039), .A(n5577), .B(n5576), .ZN(U2797)
         );
  OAI21_X1 U6732 ( .B1(n5579), .B2(n5578), .A(n4300), .ZN(n5690) );
  INV_X1 U6733 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6699) );
  INV_X1 U6734 ( .A(n5580), .ZN(n5693) );
  OAI22_X1 U6735 ( .A1(n5622), .A2(n6157), .B1(n5693), .B2(n6146), .ZN(n5584)
         );
  AOI22_X1 U6736 ( .A1(EBX_REG_29__SCAN_IN), .A2(n6161), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6158), .ZN(n5581) );
  OAI21_X1 U6737 ( .B1(n5582), .B2(n6699), .A(n5581), .ZN(n5583) );
  AOI211_X1 U6738 ( .C1(n5585), .C2(n6699), .A(n5584), .B(n5583), .ZN(n5586)
         );
  OAI21_X1 U6739 ( .B1(n5690), .B2(n6039), .A(n5586), .ZN(U2798) );
  INV_X1 U6740 ( .A(n5874), .ZN(n5595) );
  NAND2_X1 U6741 ( .A1(n6693), .A2(n5587), .ZN(n5594) );
  OAI22_X1 U6742 ( .A1(n4181), .A2(n6144), .B1(n5588), .B2(n6146), .ZN(n5593)
         );
  INV_X1 U6743 ( .A(n5630), .ZN(n5589) );
  OAI21_X1 U6744 ( .B1(n5591), .B2(n5590), .A(n5589), .ZN(n5969) );
  INV_X1 U6745 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5636) );
  OAI22_X1 U6746 ( .A1(n5969), .A2(n6157), .B1(n6129), .B2(n5636), .ZN(n5592)
         );
  AOI211_X1 U6747 ( .C1(n5595), .C2(n5594), .A(n5593), .B(n5592), .ZN(n5596)
         );
  OAI21_X1 U6748 ( .B1(n5635), .B2(n6039), .A(n5596), .ZN(U2801) );
  INV_X1 U6749 ( .A(n5599), .ZN(n5600) );
  AOI21_X1 U6750 ( .B1(n5601), .B2(n5597), .A(n5599), .ZN(n5942) );
  INV_X1 U6751 ( .A(n5942), .ZN(n5649) );
  NAND2_X1 U6752 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5893) );
  OAI211_X1 U6753 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5892), .B(n5893), .ZN(n5609) );
  INV_X1 U6754 ( .A(n5647), .ZN(n5602) );
  OAI21_X1 U6755 ( .B1(n5603), .B2(n5655), .A(n5602), .ZN(n5800) );
  INV_X1 U6756 ( .A(n5800), .ZN(n5607) );
  INV_X1 U6757 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6685) );
  OAI22_X1 U6758 ( .A1(n5919), .A2(n6685), .B1(n5728), .B2(n6146), .ZN(n5606)
         );
  INV_X1 U6759 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5604) );
  OAI22_X1 U6760 ( .A1(n5604), .A2(n6129), .B1(n3837), .B2(n6144), .ZN(n5605)
         );
  AOI211_X1 U6761 ( .C1(n6140), .C2(n5607), .A(n5606), .B(n5605), .ZN(n5608)
         );
  OAI211_X1 U6762 ( .C1(n5649), .C2(n6039), .A(n5609), .B(n5608), .ZN(U2805)
         );
  OAI22_X1 U6763 ( .A1(n5611), .A2(n6129), .B1(n6157), .B2(n5610), .ZN(n5612)
         );
  AOI211_X1 U6764 ( .C1(n6158), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6328), 
        .B(n5612), .ZN(n5619) );
  AOI22_X1 U6765 ( .A1(n5614), .A2(n5880), .B1(n6160), .B2(n5613), .ZN(n5618)
         );
  NAND2_X1 U6766 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .ZN(
        n6091) );
  OAI21_X1 U6767 ( .B1(n6091), .B2(n6101), .A(n6661), .ZN(n5616) );
  NAND2_X1 U6768 ( .A1(n5616), .A2(n5615), .ZN(n5617) );
  NAND3_X1 U6769 ( .A1(n5619), .A2(n5618), .A3(n5617), .ZN(U2819) );
  OAI22_X1 U6770 ( .A1(n5621), .A2(n5666), .B1(n5620), .B2(n6182), .ZN(U2828)
         );
  INV_X1 U6771 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5623) );
  OAI222_X1 U6772 ( .A1(n5667), .A2(n5690), .B1(n6182), .B2(n5623), .C1(n5622), 
        .C2(n5666), .ZN(U2830) );
  INV_X1 U6773 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5624) );
  OAI222_X1 U6774 ( .A1(n5667), .A2(n5931), .B1(n6182), .B2(n5624), .C1(n5763), 
        .C2(n5666), .ZN(U2831) );
  INV_X1 U6775 ( .A(n5625), .ZN(n5626) );
  AOI21_X2 U6776 ( .B1(n5628), .B2(n5627), .A(n5626), .ZN(n5881) );
  OR2_X1 U6777 ( .A1(n5630), .A2(n5629), .ZN(n5631) );
  NAND2_X1 U6778 ( .A1(n4489), .A2(n5631), .ZN(n5883) );
  OAI22_X1 U6779 ( .A1(n5883), .A2(n5666), .B1(n5632), .B2(n6182), .ZN(n5633)
         );
  AOI21_X1 U6780 ( .B1(n5881), .B2(n6179), .A(n5633), .ZN(n5634) );
  INV_X1 U6781 ( .A(n5634), .ZN(U2832) );
  OAI222_X1 U6782 ( .A1(n5636), .A2(n6182), .B1(n5666), .B2(n5969), .C1(n5635), 
        .C2(n5667), .ZN(U2833) );
  INV_X1 U6783 ( .A(n5939), .ZN(n5643) );
  NAND2_X1 U6784 ( .A1(n5645), .A2(n5638), .ZN(n5639) );
  AND2_X1 U6785 ( .A1(n5640), .A2(n5639), .ZN(n5885) );
  AOI22_X1 U6786 ( .A1(n5885), .A2(n6178), .B1(EBX_REG_24__SCAN_IN), .B2(n5641), .ZN(n5642) );
  OAI21_X1 U6787 ( .B1(n5643), .B2(n5667), .A(n5642), .ZN(U2835) );
  AOI21_X1 U6788 ( .B1(n5644), .B2(n5600), .A(n4455), .ZN(n5722) );
  INV_X1 U6789 ( .A(n5722), .ZN(n5895) );
  INV_X1 U6790 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5648) );
  OAI21_X1 U6791 ( .B1(n5647), .B2(n5646), .A(n5645), .ZN(n5894) );
  OAI222_X1 U6792 ( .A1(n5667), .A2(n5895), .B1(n6182), .B2(n5648), .C1(n5894), 
        .C2(n5666), .ZN(U2836) );
  OAI222_X1 U6793 ( .A1(n5604), .A2(n6182), .B1(n5667), .B2(n5649), .C1(n5666), 
        .C2(n5800), .ZN(U2837) );
  OAI21_X1 U6794 ( .B1(n5651), .B2(n5652), .A(n5597), .ZN(n5735) );
  INV_X1 U6795 ( .A(n5735), .ZN(n5945) );
  AND2_X1 U6796 ( .A1(n5654), .A2(n5653), .ZN(n5656) );
  OR2_X1 U6797 ( .A1(n5656), .A2(n5655), .ZN(n5911) );
  OAI22_X1 U6798 ( .A1(n5911), .A2(n5666), .B1(n5903), .B2(n6182), .ZN(n5657)
         );
  AOI21_X1 U6799 ( .B1(n5945), .B2(n6179), .A(n5657), .ZN(n5658) );
  INV_X1 U6800 ( .A(n5658), .ZN(U2838) );
  AND2_X1 U6801 ( .A1(n5519), .A2(n5659), .ZN(n5660) );
  NOR2_X1 U6802 ( .A1(n5651), .A2(n5660), .ZN(n5950) );
  INV_X1 U6803 ( .A(n5950), .ZN(n5914) );
  MUX2_X1 U6804 ( .A(n5663), .B(n5662), .S(n5661), .Z(n5665) );
  XNOR2_X1 U6805 ( .A(n5665), .B(n5664), .ZN(n5913) );
  OAI222_X1 U6806 ( .A1(n5914), .A2(n5667), .B1(n5666), .B2(n5913), .C1(n6182), 
        .C2(n5912), .ZN(U2839) );
  NAND3_X1 U6807 ( .A1(n5670), .A2(n5669), .A3(n5668), .ZN(n5672) );
  AOI22_X1 U6808 ( .A1(n6194), .A2(DATAI_31_), .B1(n6193), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U6809 ( .A1(n5672), .A2(n5671), .ZN(U2860) );
  AOI22_X1 U6810 ( .A1(n6194), .A2(DATAI_30_), .B1(n6193), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U6811 ( .A1(n6190), .A2(DATAI_14_), .ZN(n5673) );
  OAI211_X1 U6812 ( .C1(n5675), .C2(n5935), .A(n5674), .B(n5673), .ZN(U2861)
         );
  AOI22_X1 U6813 ( .A1(n6194), .A2(DATAI_29_), .B1(n6193), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5677) );
  NAND2_X1 U6814 ( .A1(n6190), .A2(DATAI_13_), .ZN(n5676) );
  OAI211_X1 U6815 ( .C1(n5690), .C2(n5935), .A(n5677), .B(n5676), .ZN(U2862)
         );
  INV_X1 U6816 ( .A(n5881), .ZN(n5680) );
  AOI22_X1 U6817 ( .A1(n6194), .A2(DATAI_27_), .B1(n6193), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U6818 ( .A1(n6190), .A2(DATAI_11_), .ZN(n5678) );
  OAI211_X1 U6819 ( .C1(n5680), .C2(n5935), .A(n5679), .B(n5678), .ZN(U2864)
         );
  AOI22_X1 U6820 ( .A1(n6194), .A2(DATAI_23_), .B1(n6193), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5682) );
  NAND2_X1 U6821 ( .A1(n6190), .A2(DATAI_7_), .ZN(n5681) );
  OAI211_X1 U6822 ( .C1(n5895), .C2(n5935), .A(n5682), .B(n5681), .ZN(U2868)
         );
  AOI21_X1 U6823 ( .B1(n6298), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5683), 
        .ZN(n5684) );
  OAI21_X1 U6824 ( .B1(n5955), .B2(n5685), .A(n5684), .ZN(n5686) );
  AOI21_X1 U6825 ( .B1(n5687), .B2(n6288), .A(n5686), .ZN(n5688) );
  OAI21_X1 U6826 ( .B1(n5689), .B2(n6016), .A(n5688), .ZN(U2956) );
  INV_X1 U6827 ( .A(n5690), .ZN(n5695) );
  AOI21_X1 U6828 ( .B1(n6298), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5691), 
        .ZN(n5692) );
  OAI21_X1 U6829 ( .B1(n5955), .B2(n5693), .A(n5692), .ZN(n5694) );
  AOI21_X1 U6830 ( .B1(n5695), .B2(n6288), .A(n5694), .ZN(n5696) );
  OAI21_X1 U6831 ( .B1(n5697), .B2(n6016), .A(n5696), .ZN(U2957) );
  NAND3_X1 U6832 ( .A1(n5698), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5848), .ZN(n5702) );
  NOR2_X1 U6833 ( .A1(n5699), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5700)
         );
  NAND2_X1 U6834 ( .A1(n5701), .A2(n5700), .ZN(n5710) );
  XNOR2_X1 U6835 ( .A(n5703), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5770)
         );
  INV_X1 U6836 ( .A(n5931), .ZN(n5707) );
  AND2_X1 U6837 ( .A1(n6284), .A2(REIP_REG_28__SCAN_IN), .ZN(n5764) );
  AOI21_X1 U6838 ( .B1(n6298), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5764), 
        .ZN(n5704) );
  OAI21_X1 U6839 ( .B1(n5955), .B2(n5705), .A(n5704), .ZN(n5706) );
  AOI21_X1 U6840 ( .B1(n5707), .B2(n6288), .A(n5706), .ZN(n5708) );
  OAI21_X1 U6841 ( .B1(n5770), .B2(n6016), .A(n5708), .ZN(U2958) );
  NAND2_X1 U6842 ( .A1(n5709), .A2(n5710), .ZN(n5711) );
  XNOR2_X1 U6843 ( .A(n5711), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5777)
         );
  NAND2_X1 U6844 ( .A1(n5961), .A2(n5871), .ZN(n5712) );
  NAND2_X1 U6845 ( .A1(n6284), .A2(REIP_REG_27__SCAN_IN), .ZN(n5772) );
  OAI211_X1 U6846 ( .C1(n5746), .C2(n5713), .A(n5712), .B(n5772), .ZN(n5714)
         );
  AOI21_X1 U6847 ( .B1(n5881), .B2(n6288), .A(n5714), .ZN(n5715) );
  OAI21_X1 U6848 ( .B1(n5777), .B2(n6016), .A(n5715), .ZN(U2959) );
  NAND2_X1 U6849 ( .A1(n5848), .A2(n5793), .ZN(n5718) );
  OAI21_X1 U6850 ( .B1(n5716), .B2(n5718), .A(n5717), .ZN(n5719) );
  XNOR2_X1 U6851 ( .A(n5719), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5798)
         );
  NAND2_X1 U6852 ( .A1(n5961), .A2(n5891), .ZN(n5720) );
  NAND2_X1 U6853 ( .A1(n6284), .A2(REIP_REG_23__SCAN_IN), .ZN(n5794) );
  OAI211_X1 U6854 ( .C1(n5746), .C2(n5901), .A(n5720), .B(n5794), .ZN(n5721)
         );
  AOI21_X1 U6855 ( .B1(n5722), .B2(n6288), .A(n5721), .ZN(n5723) );
  OAI21_X1 U6856 ( .B1(n5798), .B2(n6016), .A(n5723), .ZN(U2963) );
  AOI21_X1 U6857 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5848), .A(n5724), 
        .ZN(n5725) );
  XNOR2_X1 U6858 ( .A(n5726), .B(n5725), .ZN(n5807) );
  NOR2_X1 U6859 ( .A1(n6309), .A2(n6685), .ZN(n5802) );
  AOI21_X1 U6860 ( .B1(n6298), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5802), 
        .ZN(n5727) );
  OAI21_X1 U6861 ( .B1(n5955), .B2(n5728), .A(n5727), .ZN(n5729) );
  AOI21_X1 U6862 ( .B1(n5942), .B2(n6288), .A(n5729), .ZN(n5730) );
  OAI21_X1 U6863 ( .B1(n5807), .B2(n6016), .A(n5730), .ZN(U2964) );
  OAI21_X1 U6864 ( .B1(n5733), .B2(n5731), .A(n5732), .ZN(n5734) );
  INV_X1 U6865 ( .A(n5734), .ZN(n5815) );
  NAND2_X1 U6866 ( .A1(n6284), .A2(REIP_REG_21__SCAN_IN), .ZN(n5808) );
  OAI21_X1 U6867 ( .B1(n5746), .B2(n5902), .A(n5808), .ZN(n5737) );
  NOR2_X1 U6868 ( .A1(n5735), .A2(n6301), .ZN(n5736) );
  AOI211_X1 U6869 ( .C1(n5961), .C2(n5905), .A(n5737), .B(n5736), .ZN(n5738)
         );
  OAI21_X1 U6870 ( .B1(n5815), .B2(n6016), .A(n5738), .ZN(U2965) );
  INV_X1 U6871 ( .A(n5740), .ZN(n5742) );
  NAND2_X1 U6872 ( .A1(n5742), .A2(n5741), .ZN(n5743) );
  XNOR2_X1 U6873 ( .A(n5739), .B(n5743), .ZN(n5839) );
  NAND2_X1 U6874 ( .A1(n5961), .A2(n5923), .ZN(n5744) );
  NAND2_X1 U6875 ( .A1(n6284), .A2(REIP_REG_19__SCAN_IN), .ZN(n5832) );
  OAI211_X1 U6876 ( .C1(n5746), .C2(n5745), .A(n5744), .B(n5832), .ZN(n5747)
         );
  AOI21_X1 U6877 ( .B1(n5748), .B2(n6288), .A(n5747), .ZN(n5749) );
  OAI21_X1 U6878 ( .B1(n5839), .B2(n6016), .A(n5749), .ZN(U2967) );
  NOR2_X1 U6879 ( .A1(n5848), .A2(n3518), .ZN(n5757) );
  INV_X1 U6880 ( .A(n5752), .ZN(n5753) );
  NOR2_X1 U6881 ( .A1(n5757), .A2(n5753), .ZN(n5756) );
  OAI22_X1 U6882 ( .A1(n5751), .A2(n5757), .B1(n5756), .B2(n5755), .ZN(n5978)
         );
  INV_X1 U6883 ( .A(n6050), .ZN(n5760) );
  AOI22_X1 U6884 ( .A1(n6298), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6284), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5759) );
  OAI21_X1 U6885 ( .B1(n5955), .B2(n5760), .A(n5759), .ZN(n5761) );
  AOI21_X1 U6886 ( .B1(n6192), .B2(n6288), .A(n5761), .ZN(n5762) );
  OAI21_X1 U6887 ( .B1(n5978), .B2(n6016), .A(n5762), .ZN(U2970) );
  XNOR2_X1 U6888 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5767) );
  INV_X1 U6889 ( .A(n5763), .ZN(n5765) );
  AOI21_X1 U6890 ( .B1(n5765), .B2(n6330), .A(n5764), .ZN(n5766) );
  OAI21_X1 U6891 ( .B1(n5771), .B2(n5767), .A(n5766), .ZN(n5768) );
  AOI21_X1 U6892 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n5775), .A(n5768), 
        .ZN(n5769) );
  OAI21_X1 U6893 ( .B1(n5770), .B2(n5997), .A(n5769), .ZN(U2990) );
  NOR2_X1 U6894 ( .A1(n5771), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5774)
         );
  OAI21_X1 U6895 ( .B1(n5883), .B2(n5996), .A(n5772), .ZN(n5773) );
  AOI211_X1 U6896 ( .C1(n5775), .C2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5774), .B(n5773), .ZN(n5776) );
  OAI21_X1 U6897 ( .B1(n5777), .B2(n5997), .A(n5776), .ZN(U2991) );
  NAND2_X1 U6898 ( .A1(n5778), .A2(n6336), .ZN(n5784) );
  NAND2_X1 U6899 ( .A1(n6328), .A2(REIP_REG_25__SCAN_IN), .ZN(n5779) );
  OAI21_X1 U6900 ( .B1(n5780), .B2(n5996), .A(n5779), .ZN(n5781) );
  AOI21_X1 U6901 ( .B1(n5782), .B2(n5967), .A(n5781), .ZN(n5783) );
  OAI211_X1 U6902 ( .C1(n5975), .C2(n5967), .A(n5784), .B(n5783), .ZN(U2993)
         );
  INV_X1 U6903 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5786) );
  INV_X1 U6904 ( .A(n5824), .ZN(n5837) );
  NAND3_X1 U6905 ( .A1(n5837), .A2(n5793), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5785) );
  AOI21_X1 U6906 ( .B1(n5786), .B2(n5785), .A(n5975), .ZN(n5787) );
  AOI211_X1 U6907 ( .C1(n6330), .C2(n5885), .A(n5788), .B(n5787), .ZN(n5789)
         );
  OAI21_X1 U6908 ( .B1(n5790), .B2(n5997), .A(n5789), .ZN(U2994) );
  INV_X1 U6909 ( .A(n5791), .ZN(n5804) );
  INV_X1 U6910 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5792) );
  NAND3_X1 U6911 ( .A1(n5837), .A2(n5793), .A3(n5792), .ZN(n5795) );
  OAI211_X1 U6912 ( .C1(n5996), .C2(n5894), .A(n5795), .B(n5794), .ZN(n5796)
         );
  AOI21_X1 U6913 ( .B1(n5804), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n5796), 
        .ZN(n5797) );
  OAI21_X1 U6914 ( .B1(n5798), .B2(n5997), .A(n5797), .ZN(U2995) );
  INV_X1 U6915 ( .A(n5799), .ZN(n5803) );
  NOR2_X1 U6916 ( .A1(n5800), .A2(n5996), .ZN(n5801) );
  AOI211_X1 U6917 ( .C1(n5803), .C2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5802), .B(n5801), .ZN(n5806) );
  NAND2_X1 U6918 ( .A1(n5804), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5805) );
  OAI211_X1 U6919 ( .C1(n5807), .C2(n5997), .A(n5806), .B(n5805), .ZN(U2996)
         );
  OAI21_X1 U6920 ( .B1(n5911), .B2(n5996), .A(n5808), .ZN(n5811) );
  NOR2_X1 U6921 ( .A1(n5809), .A2(n5812), .ZN(n5810) );
  AOI211_X1 U6922 ( .C1(n5813), .C2(n5812), .A(n5811), .B(n5810), .ZN(n5814)
         );
  OAI21_X1 U6923 ( .B1(n5815), .B2(n5997), .A(n5814), .ZN(U2997) );
  AOI21_X1 U6924 ( .B1(n5817), .B2(n5816), .A(INSTADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n5818) );
  NOR2_X1 U6925 ( .A1(n5818), .A2(n5857), .ZN(n5843) );
  INV_X1 U6926 ( .A(n5843), .ZN(n5819) );
  AOI21_X1 U6927 ( .B1(n5820), .B2(n5977), .A(n5819), .ZN(n5833) );
  XNOR2_X1 U6928 ( .A(n5848), .B(n5831), .ZN(n5823) );
  XNOR2_X1 U6929 ( .A(n5822), .B(n5823), .ZN(n5951) );
  NAND2_X1 U6930 ( .A1(n5951), .A2(n6336), .ZN(n5830) );
  NOR3_X1 U6931 ( .A1(n5826), .A2(n5825), .A3(n5824), .ZN(n5828) );
  NOR2_X1 U6932 ( .A1(n5913), .A2(n5996), .ZN(n5827) );
  AOI211_X1 U6933 ( .C1(n6284), .C2(REIP_REG_20__SCAN_IN), .A(n5828), .B(n5827), .ZN(n5829) );
  OAI211_X1 U6934 ( .C1(n5833), .C2(n5831), .A(n5830), .B(n5829), .ZN(U2998)
         );
  OAI21_X1 U6935 ( .B1(n5920), .B2(n5996), .A(n5832), .ZN(n5835) );
  NOR2_X1 U6936 ( .A1(n5833), .A2(n5836), .ZN(n5834) );
  AOI211_X1 U6937 ( .C1(n5837), .C2(n5836), .A(n5835), .B(n5834), .ZN(n5838)
         );
  OAI21_X1 U6938 ( .B1(n5839), .B2(n5997), .A(n5838), .ZN(U2999) );
  NOR3_X1 U6939 ( .A1(n5755), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5848), 
        .ZN(n5850) );
  NOR3_X1 U6940 ( .A1(n5751), .A2(n4451), .A3(n5851), .ZN(n5840) );
  AOI21_X1 U6941 ( .B1(n5850), .B2(n5851), .A(n5840), .ZN(n5841) );
  XNOR2_X1 U6942 ( .A(n5841), .B(n5820), .ZN(n5956) );
  NAND2_X1 U6943 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5853), .ZN(n5844) );
  NAND2_X1 U6944 ( .A1(n6328), .A2(REIP_REG_18__SCAN_IN), .ZN(n5842) );
  OAI221_X1 U6945 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5844), .C1(
        n5820), .C2(n5843), .A(n5842), .ZN(n5845) );
  AOI21_X1 U6946 ( .B1(n6330), .B2(n5846), .A(n5845), .ZN(n5847) );
  OAI21_X1 U6947 ( .B1(n5956), .B2(n5997), .A(n5847), .ZN(U3000) );
  AND3_X1 U6948 ( .A1(n5755), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5848), 
        .ZN(n5849) );
  NOR2_X1 U6949 ( .A1(n5850), .A2(n5849), .ZN(n5852) );
  XNOR2_X1 U6950 ( .A(n5852), .B(n5851), .ZN(n5964) );
  AOI22_X1 U6951 ( .A1(n6284), .A2(REIP_REG_17__SCAN_IN), .B1(n5851), .B2(
        n5853), .ZN(n5854) );
  OAI21_X1 U6952 ( .B1(n5855), .B2(n5996), .A(n5854), .ZN(n5856) );
  AOI21_X1 U6953 ( .B1(n5857), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5856), 
        .ZN(n5858) );
  OAI21_X1 U6954 ( .B1(n5964), .B2(n5997), .A(n5858), .ZN(U3001) );
  OAI211_X1 U6955 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n4702), .A(n6505), .B(
        n6513), .ZN(n5859) );
  OAI21_X1 U6956 ( .B1(n5860), .B2(n5863), .A(n5859), .ZN(n5861) );
  MUX2_X1 U6957 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5861), .S(n6344), 
        .Z(U3464) );
  XNOR2_X1 U6958 ( .A(n6345), .B(n6505), .ZN(n5864) );
  INV_X1 U6959 ( .A(n5862), .ZN(n6150) );
  OAI22_X1 U6960 ( .A1(n5864), .A2(n6352), .B1(n6150), .B2(n5863), .ZN(n5865)
         );
  MUX2_X1 U6961 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5865), .S(n6344), 
        .Z(U3463) );
  OAI22_X1 U6962 ( .A1(n5868), .A2(n5867), .B1(n5866), .B2(n6604), .ZN(n5870)
         );
  MUX2_X1 U6963 ( .A(n5870), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n5869), 
        .Z(U3456) );
  AND2_X1 U6964 ( .A1(n6226), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U6965 ( .A1(n6160), .A2(n5871), .B1(PHYADDRPOINTER_REG_27__SCAN_IN), 
        .B2(n6158), .ZN(n5873) );
  NAND2_X1 U6966 ( .A1(n6161), .A2(EBX_REG_27__SCAN_IN), .ZN(n5872) );
  OAI211_X1 U6967 ( .C1(n5874), .C2(n6695), .A(n5873), .B(n5872), .ZN(n5875)
         );
  INV_X1 U6968 ( .A(n5875), .ZN(n5878) );
  OAI21_X1 U6969 ( .B1(n5883), .B2(n6157), .A(n5882), .ZN(U2800) );
  AOI22_X1 U6970 ( .A1(EBX_REG_24__SCAN_IN), .A2(n6161), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n6158), .ZN(n5890) );
  AOI22_X1 U6971 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5898), .B1(n5884), .B2(
        n6160), .ZN(n5889) );
  AOI22_X1 U6972 ( .A1(n5939), .A2(n5880), .B1(n5885), .B2(n6140), .ZN(n5888)
         );
  INV_X1 U6973 ( .A(n5886), .ZN(n5887) );
  NAND4_X1 U6974 ( .A1(n5890), .A2(n5889), .A3(n5888), .A4(n5887), .ZN(U2803)
         );
  AOI22_X1 U6975 ( .A1(EBX_REG_23__SCAN_IN), .A2(n6161), .B1(n5891), .B2(n6160), .ZN(n5900) );
  INV_X1 U6976 ( .A(n5892), .ZN(n5908) );
  INV_X1 U6977 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6688) );
  OAI21_X1 U6978 ( .B1(n5908), .B2(n5893), .A(n6688), .ZN(n5897) );
  OAI22_X1 U6979 ( .A1(n5895), .A2(n6039), .B1(n5894), .B2(n6157), .ZN(n5896)
         );
  AOI21_X1 U6980 ( .B1(n5898), .B2(n5897), .A(n5896), .ZN(n5899) );
  OAI211_X1 U6981 ( .C1(n5901), .C2(n6144), .A(n5900), .B(n5899), .ZN(U2804)
         );
  INV_X1 U6982 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5907) );
  OAI22_X1 U6983 ( .A1(n5903), .A2(n6129), .B1(n5902), .B2(n6144), .ZN(n5904)
         );
  AOI21_X1 U6984 ( .B1(n5905), .B2(n6160), .A(n5904), .ZN(n5906) );
  OAI221_X1 U6985 ( .B1(REIP_REG_21__SCAN_IN), .B2(n5908), .C1(n5907), .C2(
        n5919), .A(n5906), .ZN(n5909) );
  AOI21_X1 U6986 ( .B1(n5945), .B2(n5880), .A(n5909), .ZN(n5910) );
  OAI21_X1 U6987 ( .B1(n5911), .B2(n6157), .A(n5910), .ZN(U2806) );
  OAI22_X1 U6988 ( .A1(n5912), .A2(n6129), .B1(n5954), .B2(n6146), .ZN(n5916)
         );
  OAI22_X1 U6989 ( .A1(n5914), .A2(n6039), .B1(n5913), .B2(n6157), .ZN(n5915)
         );
  AOI211_X1 U6990 ( .C1(PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n6158), .A(n5916), 
        .B(n5915), .ZN(n5917) );
  OAI221_X1 U6991 ( .B1(n5919), .B2(n6683), .C1(n5919), .C2(n5918), .A(n5917), 
        .ZN(U2807) );
  AOI21_X1 U6992 ( .B1(n6158), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6328), 
        .ZN(n5928) );
  AOI22_X1 U6993 ( .A1(EBX_REG_19__SCAN_IN), .A2(n6161), .B1(
        REIP_REG_19__SCAN_IN), .B2(n6035), .ZN(n5927) );
  OAI22_X1 U6994 ( .A1(n5921), .A2(n6039), .B1(n5920), .B2(n6157), .ZN(n5922)
         );
  AOI21_X1 U6995 ( .B1(n5923), .B2(n6160), .A(n5922), .ZN(n5926) );
  OAI211_X1 U6996 ( .C1(REIP_REG_19__SCAN_IN), .C2(REIP_REG_18__SCAN_IN), .A(
        n6034), .B(n5924), .ZN(n5925) );
  NAND4_X1 U6997 ( .A1(n5928), .A2(n5927), .A3(n5926), .A4(n5925), .ZN(U2808)
         );
  INV_X1 U6998 ( .A(n6190), .ZN(n5930) );
  INV_X1 U6999 ( .A(n5932), .ZN(n5934) );
  AOI22_X1 U7000 ( .A1(n6194), .A2(DATAI_28_), .B1(n6193), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5933) );
  NAND2_X1 U7001 ( .A1(n5934), .A2(n5933), .ZN(U2863) );
  AOI22_X1 U7002 ( .A1(n5936), .A2(n6191), .B1(n6190), .B2(DATAI_10_), .ZN(
        n5938) );
  AOI22_X1 U7003 ( .A1(n6194), .A2(DATAI_26_), .B1(n6193), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5937) );
  NAND2_X1 U7004 ( .A1(n5938), .A2(n5937), .ZN(U2865) );
  AOI22_X1 U7005 ( .A1(n5939), .A2(n6191), .B1(DATAI_8_), .B2(n6190), .ZN(
        n5941) );
  AOI22_X1 U7006 ( .A1(n6194), .A2(DATAI_24_), .B1(n6193), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U7007 ( .A1(n5941), .A2(n5940), .ZN(U2867) );
  AOI22_X1 U7008 ( .A1(n5942), .A2(n6191), .B1(n6190), .B2(DATAI_6_), .ZN(
        n5944) );
  AOI22_X1 U7009 ( .A1(n6194), .A2(DATAI_22_), .B1(n6193), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5943) );
  NAND2_X1 U7010 ( .A1(n5944), .A2(n5943), .ZN(U2869) );
  AOI22_X1 U7011 ( .A1(n5945), .A2(n6191), .B1(n6190), .B2(DATAI_5_), .ZN(
        n5947) );
  AOI22_X1 U7012 ( .A1(n6194), .A2(DATAI_21_), .B1(n6193), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U7013 ( .A1(n5947), .A2(n5946), .ZN(U2870) );
  AOI22_X1 U7014 ( .A1(n5950), .A2(n6191), .B1(n6190), .B2(DATAI_4_), .ZN(
        n5949) );
  AOI22_X1 U7015 ( .A1(n6194), .A2(DATAI_20_), .B1(n6193), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U7016 ( .A1(n5949), .A2(n5948), .ZN(U2871) );
  AOI22_X1 U7017 ( .A1(n6328), .A2(REIP_REG_20__SCAN_IN), .B1(n6298), .B2(
        PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5953) );
  AOI22_X1 U7018 ( .A1(n5951), .A2(n6296), .B1(n6288), .B2(n5950), .ZN(n5952)
         );
  OAI211_X1 U7019 ( .C1(n5955), .C2(n5954), .A(n5953), .B(n5952), .ZN(U2966)
         );
  AOI22_X1 U7020 ( .A1(n6328), .A2(REIP_REG_18__SCAN_IN), .B1(n6298), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5959) );
  INV_X1 U7021 ( .A(n5956), .ZN(n5957) );
  AOI22_X1 U7022 ( .A1(n5957), .A2(n6296), .B1(n6288), .B2(n6184), .ZN(n5958)
         );
  OAI211_X1 U7023 ( .C1(n5955), .C2(n6044), .A(n5959), .B(n5958), .ZN(U2968)
         );
  AOI22_X1 U7024 ( .A1(n6328), .A2(REIP_REG_17__SCAN_IN), .B1(n6298), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5963) );
  AOI22_X1 U7025 ( .A1(n6187), .A2(n6288), .B1(n5961), .B2(n5960), .ZN(n5962)
         );
  OAI211_X1 U7026 ( .C1(n5964), .C2(n6016), .A(n5963), .B(n5962), .ZN(U2969)
         );
  AOI211_X1 U7027 ( .C1(n5974), .C2(n5967), .A(n5966), .B(n5965), .ZN(n5968)
         );
  AOI21_X1 U7028 ( .B1(REIP_REG_26__SCAN_IN), .B2(n6328), .A(n5968), .ZN(n5973) );
  INV_X1 U7029 ( .A(n5969), .ZN(n5970) );
  AOI22_X1 U7030 ( .A1(n5971), .A2(n6336), .B1(n6330), .B2(n5970), .ZN(n5972)
         );
  OAI211_X1 U7031 ( .C1(n5975), .C2(n5974), .A(n5973), .B(n5972), .ZN(U2992)
         );
  AOI21_X1 U7032 ( .B1(n5977), .B2(n5985), .A(n5976), .ZN(n5986) );
  AOI211_X1 U7033 ( .C1(n3518), .C2(n5987), .A(n5984), .B(n5985), .ZN(n5981)
         );
  OAI22_X1 U7034 ( .A1(n5978), .A2(n5997), .B1(n5996), .B2(n6053), .ZN(n5979)
         );
  AOI21_X1 U7035 ( .B1(n5981), .B2(n5980), .A(n5979), .ZN(n5983) );
  NAND2_X1 U7036 ( .A1(n6328), .A2(REIP_REG_16__SCAN_IN), .ZN(n5982) );
  OAI211_X1 U7037 ( .C1(n5986), .C2(n3518), .A(n5983), .B(n5982), .ZN(U3002)
         );
  OR2_X1 U7038 ( .A1(n5985), .A2(n5984), .ZN(n5993) );
  INV_X1 U7039 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6675) );
  OAI22_X1 U7040 ( .A1(n5987), .A2(n5986), .B1(n6309), .B2(n6675), .ZN(n5988)
         );
  INV_X1 U7041 ( .A(n5988), .ZN(n5992) );
  AOI22_X1 U7042 ( .A1(n5990), .A2(n6336), .B1(n6330), .B2(n5989), .ZN(n5991)
         );
  OAI211_X1 U7043 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n5993), .A(n5992), .B(n5991), .ZN(U3003) );
  INV_X1 U7044 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6672) );
  AOI21_X1 U7045 ( .B1(n5995), .B2(n5994), .A(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n6001) );
  OAI22_X1 U7046 ( .A1(n5998), .A2(n5997), .B1(n5996), .B2(n6065), .ZN(n5999)
         );
  AOI221_X1 U7047 ( .B1(n6001), .B2(INSTADDRPOINTER_REG_14__SCAN_IN), .C1(
        n6000), .C2(INSTADDRPOINTER_REG_14__SCAN_IN), .A(n5999), .ZN(n6005) );
  NAND3_X1 U7048 ( .A1(n6003), .A2(n6002), .A3(n6306), .ZN(n6004) );
  OAI211_X1 U7049 ( .C1(n6672), .C2(n6309), .A(n6005), .B(n6004), .ZN(U3004)
         );
  INV_X1 U7050 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6648) );
  AOI21_X1 U7051 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6648), .A(n6631), .ZN(n6013) );
  NAND2_X1 U7052 ( .A1(n6631), .A2(STATE_REG_1__SCAN_IN), .ZN(n6726) );
  AOI21_X1 U7053 ( .B1(n6013), .B2(n6006), .A(n6708), .ZN(U2789) );
  INV_X1 U7054 ( .A(n6007), .ZN(n6011) );
  INV_X1 U7055 ( .A(n6008), .ZN(n6009) );
  OAI21_X1 U7056 ( .B1(n6009), .B2(n6598), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6010) );
  OAI21_X1 U7057 ( .B1(n6011), .B2(n6615), .A(n6010), .ZN(U2790) );
  NOR2_X1 U7058 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n6014) );
  OAI21_X1 U7059 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6014), .A(n6740), .ZN(n6012)
         );
  OAI21_X1 U7060 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6726), .A(n6012), .ZN(
        U2791) );
  NOR2_X1 U7061 ( .A1(n6708), .A2(n6013), .ZN(n6712) );
  OAI21_X1 U7062 ( .B1(n6014), .B2(BS16_N), .A(n6712), .ZN(n6710) );
  OAI21_X1 U7063 ( .B1(n6712), .B2(n6015), .A(n6710), .ZN(U2792) );
  OAI21_X1 U7064 ( .B1(n6018), .B2(n6017), .A(n6016), .ZN(U2793) );
  AOI211_X1 U7065 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_2__SCAN_IN), .B(
        DATAWIDTH_REG_4__SCAN_IN), .ZN(n6019) );
  NAND4_X1 U7066 ( .A1(n6020), .A2(n6019), .A3(n6628), .A4(n6629), .ZN(n6028)
         );
  OR4_X1 U7067 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6027)
         );
  OR4_X1 U7068 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_9__SCAN_IN), .A4(DATAWIDTH_REG_10__SCAN_IN), .ZN(
        n6026) );
  NOR4_X1 U7069 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_21__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n6024) );
  NOR4_X1 U7070 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_17__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n6023) );
  NOR4_X1 U7071 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6022) );
  NOR4_X1 U7072 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n6021) );
  NAND4_X1 U7073 ( .A1(n6024), .A2(n6023), .A3(n6022), .A4(n6021), .ZN(n6025)
         );
  NOR4_X2 U7074 ( .A1(n6028), .A2(n6027), .A3(n6026), .A4(n6025), .ZN(n6724)
         );
  INV_X1 U7075 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6030) );
  NOR3_X1 U7076 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6031) );
  OAI21_X1 U7077 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6031), .A(n6724), .ZN(n6029)
         );
  OAI21_X1 U7078 ( .B1(n6724), .B2(n6030), .A(n6029), .ZN(U2794) );
  INV_X1 U7079 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6711) );
  AOI21_X1 U7080 ( .B1(n6717), .B2(n6711), .A(n6031), .ZN(n6033) );
  INV_X1 U7081 ( .A(n6724), .ZN(n6719) );
  AOI22_X1 U7082 ( .A1(n6724), .A2(n6033), .B1(n6032), .B2(n6719), .ZN(U2795)
         );
  INV_X1 U7083 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6037) );
  INV_X1 U7084 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6680) );
  AOI22_X1 U7085 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6035), .B1(n6034), .B2(
        n6680), .ZN(n6036) );
  OAI211_X1 U7086 ( .C1(n6144), .C2(n6037), .A(n6036), .B(n6309), .ZN(n6042)
         );
  OAI22_X1 U7087 ( .A1(n6040), .A2(n6039), .B1(n6038), .B2(n6157), .ZN(n6041)
         );
  AOI211_X1 U7088 ( .C1(EBX_REG_18__SCAN_IN), .C2(n6161), .A(n6042), .B(n6041), 
        .ZN(n6043) );
  OAI21_X1 U7089 ( .B1(n6044), .B2(n6146), .A(n6043), .ZN(U2809) );
  NAND2_X1 U7090 ( .A1(n6045), .A2(REIP_REG_15__SCAN_IN), .ZN(n6048) );
  AOI22_X1 U7091 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6161), .B1(
        REIP_REG_16__SCAN_IN), .B2(n6046), .ZN(n6047) );
  OAI21_X1 U7092 ( .B1(REIP_REG_16__SCAN_IN), .B2(n6048), .A(n6047), .ZN(n6049) );
  AOI211_X1 U7093 ( .C1(n6158), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6328), 
        .B(n6049), .ZN(n6052) );
  AOI22_X1 U7094 ( .A1(n6192), .A2(n5880), .B1(n6160), .B2(n6050), .ZN(n6051)
         );
  OAI211_X1 U7095 ( .C1(n6157), .C2(n6053), .A(n6052), .B(n6051), .ZN(U2811)
         );
  NOR3_X1 U7096 ( .A1(n6055), .A2(n6054), .A3(n6672), .ZN(n6060) );
  INV_X1 U7097 ( .A(n6131), .ZN(n6159) );
  NAND3_X1 U7098 ( .A1(n6159), .A2(n6672), .A3(n6056), .ZN(n6057) );
  OAI211_X1 U7099 ( .C1(n6144), .C2(n6058), .A(n6309), .B(n6057), .ZN(n6059)
         );
  AOI211_X1 U7100 ( .C1(n6161), .C2(EBX_REG_14__SCAN_IN), .A(n6060), .B(n6059), 
        .ZN(n6064) );
  AOI22_X1 U7101 ( .A1(n6062), .A2(n5880), .B1(n6160), .B2(n6061), .ZN(n6063)
         );
  OAI211_X1 U7102 ( .C1(n6157), .C2(n6065), .A(n6064), .B(n6063), .ZN(U2813)
         );
  INV_X1 U7103 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6068) );
  AOI22_X1 U7104 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6161), .B1(n6140), .B2(n6066), .ZN(n6067) );
  OAI211_X1 U7105 ( .C1(n6144), .C2(n6068), .A(n6067), .B(n6309), .ZN(n6071)
         );
  NOR3_X1 U7106 ( .A1(n6131), .A2(REIP_REG_13__SCAN_IN), .A3(n6069), .ZN(n6070) );
  AOI211_X1 U7107 ( .C1(n6072), .C2(n5880), .A(n6071), .B(n6070), .ZN(n6075)
         );
  NOR3_X1 U7108 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6668), .A3(n6073), .ZN(n6083) );
  OAI21_X1 U7109 ( .B1(n6083), .B2(n6079), .A(REIP_REG_13__SCAN_IN), .ZN(n6074) );
  OAI211_X1 U7110 ( .C1(n6146), .C2(n6076), .A(n6075), .B(n6074), .ZN(U2814)
         );
  INV_X1 U7111 ( .A(n6077), .ZN(n6174) );
  AOI22_X1 U7112 ( .A1(n6174), .A2(n5880), .B1(n6078), .B2(n6160), .ZN(n6085)
         );
  AOI22_X1 U7113 ( .A1(n6140), .A2(n6173), .B1(REIP_REG_12__SCAN_IN), .B2(
        n6079), .ZN(n6080) );
  OAI211_X1 U7114 ( .C1(n6144), .C2(n6081), .A(n6080), .B(n6309), .ZN(n6082)
         );
  AOI211_X1 U7115 ( .C1(n6161), .C2(EBX_REG_12__SCAN_IN), .A(n6083), .B(n6082), 
        .ZN(n6084) );
  NAND2_X1 U7116 ( .A1(n6085), .A2(n6084), .ZN(U2815) );
  INV_X1 U7117 ( .A(n6086), .ZN(n6087) );
  OR2_X1 U7118 ( .A1(n6131), .A2(n6087), .ZN(n6088) );
  AND2_X1 U7119 ( .A1(n4264), .A2(n6088), .ZN(n6142) );
  OAI21_X1 U7120 ( .B1(n6089), .B2(n6131), .A(n6142), .ZN(n6114) );
  INV_X1 U7121 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6090) );
  AOI21_X1 U7122 ( .B1(n6090), .B2(n6658), .A(n6101), .ZN(n6092) );
  AOI22_X1 U7123 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6114), .B1(n6092), .B2(n6091), .ZN(n6099) );
  INV_X1 U7124 ( .A(n6093), .ZN(n6319) );
  AOI22_X1 U7125 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6161), .B1(n6140), .B2(n6319), 
        .ZN(n6094) );
  OAI211_X1 U7126 ( .C1(n6144), .C2(n6095), .A(n6094), .B(n6309), .ZN(n6096)
         );
  AOI21_X1 U7127 ( .B1(n6097), .B2(n5880), .A(n6096), .ZN(n6098) );
  OAI211_X1 U7128 ( .C1(n6100), .C2(n6146), .A(n6099), .B(n6098), .ZN(U2820)
         );
  INV_X1 U7129 ( .A(n6101), .ZN(n6104) );
  AOI22_X1 U7130 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6158), .B1(n6140), 
        .B2(n6177), .ZN(n6102) );
  OAI211_X1 U7131 ( .C1(n6129), .C2(n6183), .A(n6102), .B(n6309), .ZN(n6103)
         );
  AOI221_X1 U7132 ( .B1(n6104), .B2(n6658), .C1(n6114), .C2(
        REIP_REG_6__SCAN_IN), .A(n6103), .ZN(n6108) );
  INV_X1 U7133 ( .A(n6105), .ZN(n6106) );
  AOI22_X1 U7134 ( .A1(n6180), .A2(n5880), .B1(n6106), .B2(n6160), .ZN(n6107)
         );
  NAND2_X1 U7135 ( .A1(n6108), .A2(n6107), .ZN(U2821) );
  AOI22_X1 U7136 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6161), .B1(n6140), .B2(n6109), 
        .ZN(n6110) );
  OAI211_X1 U7137 ( .C1(n6144), .C2(n6111), .A(n6110), .B(n6309), .ZN(n6112)
         );
  AOI21_X1 U7138 ( .B1(n6113), .B2(n6152), .A(n6112), .ZN(n6116) );
  OAI221_X1 U7139 ( .B1(REIP_REG_5__SCAN_IN), .B2(REIP_REG_4__SCAN_IN), .C1(
        REIP_REG_5__SCAN_IN), .C2(n6126), .A(n6114), .ZN(n6115) );
  OAI211_X1 U7140 ( .C1(n6146), .C2(n6117), .A(n6116), .B(n6115), .ZN(U2822)
         );
  AOI22_X1 U7141 ( .A1(n6140), .A2(n6119), .B1(n6162), .B2(n6118), .ZN(n6120)
         );
  INV_X1 U7142 ( .A(n6120), .ZN(n6121) );
  AOI211_X1 U7143 ( .C1(n6158), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6328), 
        .B(n6121), .ZN(n6128) );
  INV_X1 U7144 ( .A(n6142), .ZN(n6125) );
  OAI22_X1 U7145 ( .A1(n6123), .A2(n6166), .B1(n6122), .B2(n6146), .ZN(n6124)
         );
  AOI221_X1 U7146 ( .B1(n6126), .B2(n6654), .C1(n6125), .C2(
        REIP_REG_4__SCAN_IN), .A(n6124), .ZN(n6127) );
  OAI211_X1 U7147 ( .C1(n6130), .C2(n6129), .A(n6128), .B(n6127), .ZN(U2823)
         );
  OAI211_X1 U7148 ( .C1(REIP_REG_1__SCAN_IN), .C2(n6131), .A(n4264), .B(
        REIP_REG_2__SCAN_IN), .ZN(n6153) );
  INV_X1 U7149 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6132) );
  OAI22_X1 U7150 ( .A1(n6146), .A2(n6133), .B1(n6132), .B2(n6144), .ZN(n6134)
         );
  AOI21_X1 U7151 ( .B1(n6161), .B2(EBX_REG_3__SCAN_IN), .A(n6134), .ZN(n6136)
         );
  NAND2_X1 U7152 ( .A1(n2977), .A2(n6162), .ZN(n6135) );
  OAI211_X1 U7153 ( .C1(n6137), .C2(n6166), .A(n6136), .B(n6135), .ZN(n6138)
         );
  AOI21_X1 U7154 ( .B1(n6140), .B2(n6139), .A(n6138), .ZN(n6141) );
  OAI221_X1 U7155 ( .B1(n6142), .B2(n6652), .C1(n6142), .C2(n6153), .A(n6141), 
        .ZN(U2824) );
  INV_X1 U7156 ( .A(n6143), .ZN(n6289) );
  INV_X1 U7157 ( .A(n6162), .ZN(n6149) );
  OAI22_X1 U7158 ( .A1(n6146), .A2(n6292), .B1(n6145), .B2(n6144), .ZN(n6147)
         );
  AOI21_X1 U7159 ( .B1(n6161), .B2(EBX_REG_2__SCAN_IN), .A(n6147), .ZN(n6148)
         );
  OAI21_X1 U7160 ( .B1(n6150), .B2(n6149), .A(n6148), .ZN(n6151) );
  AOI21_X1 U7161 ( .B1(n6289), .B2(n6152), .A(n6151), .ZN(n6156) );
  OAI21_X1 U7162 ( .B1(REIP_REG_2__SCAN_IN), .B2(n6154), .A(n6153), .ZN(n6155)
         );
  OAI211_X1 U7163 ( .C1(n6157), .C2(n6327), .A(n6156), .B(n6155), .ZN(U2825)
         );
  AOI22_X1 U7164 ( .A1(n6159), .A2(n6717), .B1(PHYADDRPOINTER_REG_1__SCAN_IN), 
        .B2(n6158), .ZN(n6172) );
  INV_X1 U7165 ( .A(n4556), .ZN(n6169) );
  AOI22_X1 U7166 ( .A1(n6161), .A2(EBX_REG_1__SCAN_IN), .B1(n6160), .B2(n3551), 
        .ZN(n6165) );
  NAND2_X1 U7167 ( .A1(n6163), .A2(n6162), .ZN(n6164) );
  OAI211_X1 U7168 ( .C1(n6167), .C2(n6166), .A(n6165), .B(n6164), .ZN(n6168)
         );
  AOI21_X1 U7169 ( .B1(n6170), .B2(n6169), .A(n6168), .ZN(n6171) );
  OAI211_X1 U7170 ( .C1(n6717), .C2(n4264), .A(n6172), .B(n6171), .ZN(U2826)
         );
  AOI22_X1 U7171 ( .A1(n6174), .A2(n6179), .B1(n6178), .B2(n6173), .ZN(n6175)
         );
  OAI21_X1 U7172 ( .B1(n6176), .B2(n6182), .A(n6175), .ZN(U2847) );
  AOI22_X1 U7173 ( .A1(n6180), .A2(n6179), .B1(n6178), .B2(n6177), .ZN(n6181)
         );
  OAI21_X1 U7174 ( .B1(n6183), .B2(n6182), .A(n6181), .ZN(U2853) );
  AOI22_X1 U7175 ( .A1(n6184), .A2(n6191), .B1(n6190), .B2(DATAI_2_), .ZN(
        n6186) );
  AOI22_X1 U7176 ( .A1(n6194), .A2(DATAI_18_), .B1(n6193), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6185) );
  NAND2_X1 U7177 ( .A1(n6186), .A2(n6185), .ZN(U2873) );
  AOI22_X1 U7178 ( .A1(n6187), .A2(n6191), .B1(n6190), .B2(DATAI_1_), .ZN(
        n6189) );
  AOI22_X1 U7179 ( .A1(n6194), .A2(DATAI_17_), .B1(n6193), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U7180 ( .A1(n6189), .A2(n6188), .ZN(U2874) );
  AOI22_X1 U7181 ( .A1(n6192), .A2(n6191), .B1(n6190), .B2(DATAI_0_), .ZN(
        n6196) );
  AOI22_X1 U7182 ( .A1(n6194), .A2(DATAI_16_), .B1(n6193), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U7183 ( .A1(n6196), .A2(n6195), .ZN(U2875) );
  INV_X1 U7184 ( .A(n6197), .ZN(n6201) );
  AOI22_X1 U7185 ( .A1(n6201), .A2(EAX_REG_24__SCAN_IN), .B1(
        UWORD_REG_8__SCAN_IN), .B2(n6730), .ZN(n6198) );
  OAI21_X1 U7186 ( .B1(n6200), .B2(n6199), .A(n6198), .ZN(U2899) );
  AOI22_X1 U7187 ( .A1(n6226), .A2(DATAO_REG_17__SCAN_IN), .B1(n6201), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6202) );
  OAI21_X1 U7188 ( .B1(n6203), .B2(n6597), .A(n6202), .ZN(U2906) );
  AOI22_X1 U7189 ( .A1(n6730), .A2(LWORD_REG_15__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6204) );
  OAI21_X1 U7190 ( .B1(n6205), .B2(n6228), .A(n6204), .ZN(U2908) );
  INV_X1 U7191 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6283) );
  AOI22_X1 U7192 ( .A1(n6730), .A2(LWORD_REG_14__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6206) );
  OAI21_X1 U7193 ( .B1(n6283), .B2(n6228), .A(n6206), .ZN(U2909) );
  INV_X1 U7194 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6278) );
  AOI22_X1 U7195 ( .A1(n6730), .A2(LWORD_REG_13__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6207) );
  OAI21_X1 U7196 ( .B1(n6278), .B2(n6228), .A(n6207), .ZN(U2910) );
  AOI22_X1 U7197 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6210), .B1(n6226), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6208) );
  OAI21_X1 U7198 ( .B1(n6209), .B2(n6597), .A(n6208), .ZN(U2911) );
  AOI222_X1 U7199 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n6730), .B1(n6210), .B2(
        EAX_REG_11__SCAN_IN), .C1(n6226), .C2(DATAO_REG_11__SCAN_IN), .ZN(
        n6211) );
  INV_X1 U7200 ( .A(n6211), .ZN(U2912) );
  AOI22_X1 U7201 ( .A1(n6730), .A2(LWORD_REG_10__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6212) );
  OAI21_X1 U7202 ( .B1(n6213), .B2(n6228), .A(n6212), .ZN(U2913) );
  AOI22_X1 U7203 ( .A1(n6730), .A2(LWORD_REG_9__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6214) );
  OAI21_X1 U7204 ( .B1(n3623), .B2(n6228), .A(n6214), .ZN(U2914) );
  INV_X1 U7205 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6216) );
  AOI22_X1 U7206 ( .A1(n6730), .A2(LWORD_REG_8__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6215) );
  OAI21_X1 U7207 ( .B1(n6216), .B2(n6228), .A(n6215), .ZN(U2915) );
  AOI22_X1 U7208 ( .A1(n6730), .A2(LWORD_REG_7__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6217) );
  OAI21_X1 U7209 ( .B1(n3533), .B2(n6228), .A(n6217), .ZN(U2916) );
  AOI22_X1 U7210 ( .A1(n6730), .A2(LWORD_REG_6__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6218) );
  OAI21_X1 U7211 ( .B1(n5048), .B2(n6228), .A(n6218), .ZN(U2917) );
  AOI22_X1 U7212 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n6730), .B1(n6226), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6219) );
  OAI21_X1 U7213 ( .B1(n6220), .B2(n6228), .A(n6219), .ZN(U2918) );
  AOI22_X1 U7214 ( .A1(n6730), .A2(LWORD_REG_4__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6221) );
  OAI21_X1 U7215 ( .B1(n6222), .B2(n6228), .A(n6221), .ZN(U2919) );
  AOI22_X1 U7216 ( .A1(n6730), .A2(LWORD_REG_3__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6223) );
  OAI21_X1 U7217 ( .B1(n3563), .B2(n6228), .A(n6223), .ZN(U2920) );
  AOI22_X1 U7218 ( .A1(n6730), .A2(LWORD_REG_2__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6224) );
  OAI21_X1 U7219 ( .B1(n3554), .B2(n6228), .A(n6224), .ZN(U2921) );
  AOI22_X1 U7220 ( .A1(n6730), .A2(LWORD_REG_1__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6225) );
  OAI21_X1 U7221 ( .B1(n3538), .B2(n6228), .A(n6225), .ZN(U2922) );
  AOI22_X1 U7222 ( .A1(n6730), .A2(LWORD_REG_0__SCAN_IN), .B1(n6226), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6227) );
  OAI21_X1 U7223 ( .B1(n3546), .B2(n6228), .A(n6227), .ZN(U2923) );
  AOI22_X1 U7224 ( .A1(n6276), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n6271), .ZN(n6229) );
  OAI21_X1 U7225 ( .B1(n6273), .B2(n6251), .A(n6229), .ZN(U2924) );
  AOI22_X1 U7226 ( .A1(n6280), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n6271), .ZN(n6230) );
  OAI21_X1 U7227 ( .B1(n6273), .B2(n6253), .A(n6230), .ZN(U2925) );
  AOI22_X1 U7228 ( .A1(n6280), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n6271), .ZN(n6231) );
  OAI21_X1 U7229 ( .B1(n6273), .B2(n6255), .A(n6231), .ZN(U2926) );
  AOI22_X1 U7230 ( .A1(n6276), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n6271), .ZN(n6232) );
  OAI21_X1 U7231 ( .B1(n6257), .B2(n6273), .A(n6232), .ZN(U2927) );
  AOI22_X1 U7232 ( .A1(n6276), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n6271), .ZN(n6233) );
  OAI21_X1 U7233 ( .B1(n6273), .B2(n6259), .A(n6233), .ZN(U2928) );
  AOI22_X1 U7234 ( .A1(n6276), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n6271), .ZN(n6234) );
  OAI21_X1 U7235 ( .B1(n6273), .B2(n6261), .A(n6234), .ZN(U2929) );
  AOI22_X1 U7236 ( .A1(n6276), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n6271), .ZN(n6235) );
  OAI21_X1 U7237 ( .B1(n5047), .B2(n6273), .A(n6235), .ZN(U2930) );
  AOI22_X1 U7238 ( .A1(n6276), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6271), .ZN(n6236) );
  OAI21_X1 U7239 ( .B1(n6273), .B2(n6264), .A(n6236), .ZN(U2931) );
  AOI22_X1 U7240 ( .A1(n6276), .A2(UWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n6271), .ZN(n6238) );
  NAND2_X1 U7241 ( .A1(n6237), .A2(DATAI_8_), .ZN(n6265) );
  NAND2_X1 U7242 ( .A1(n6238), .A2(n6265), .ZN(U2932) );
  AOI22_X1 U7243 ( .A1(n6276), .A2(UWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_25__SCAN_IN), .B2(n6271), .ZN(n6239) );
  OAI21_X1 U7244 ( .B1(n6273), .B2(n6268), .A(n6239), .ZN(U2933) );
  AOI22_X1 U7245 ( .A1(n6276), .A2(UWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_26__SCAN_IN), .B2(n6271), .ZN(n6240) );
  OAI21_X1 U7246 ( .B1(n6270), .B2(n6273), .A(n6240), .ZN(U2934) );
  AOI22_X1 U7247 ( .A1(n6276), .A2(UWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_27__SCAN_IN), .B2(n6271), .ZN(n6241) );
  OAI21_X1 U7248 ( .B1(n6274), .B2(n6273), .A(n6241), .ZN(U2935) );
  AOI21_X1 U7249 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6280), .A(n6242), .ZN(
        n6243) );
  OAI21_X1 U7250 ( .B1(n4153), .B2(n6282), .A(n6243), .ZN(U2936) );
  INV_X1 U7251 ( .A(DATAI_13_), .ZN(n6244) );
  NOR2_X1 U7252 ( .A1(n6273), .A2(n6244), .ZN(n6275) );
  AOI21_X1 U7253 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n6280), .A(n6275), .ZN(
        n6245) );
  OAI21_X1 U7254 ( .B1(n6246), .B2(n6282), .A(n6245), .ZN(U2937) );
  INV_X1 U7255 ( .A(DATAI_14_), .ZN(n6247) );
  NOR2_X1 U7256 ( .A1(n6273), .A2(n6247), .ZN(n6279) );
  AOI21_X1 U7257 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6276), .A(n6279), .ZN(
        n6248) );
  OAI21_X1 U7258 ( .B1(n6249), .B2(n6282), .A(n6248), .ZN(U2938) );
  AOI22_X1 U7259 ( .A1(n6276), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n6271), .ZN(n6250) );
  OAI21_X1 U7260 ( .B1(n6273), .B2(n6251), .A(n6250), .ZN(U2939) );
  AOI22_X1 U7261 ( .A1(n6276), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n6271), .ZN(n6252) );
  OAI21_X1 U7262 ( .B1(n6273), .B2(n6253), .A(n6252), .ZN(U2940) );
  AOI22_X1 U7263 ( .A1(n6276), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6271), .ZN(n6254) );
  OAI21_X1 U7264 ( .B1(n6273), .B2(n6255), .A(n6254), .ZN(U2941) );
  AOI22_X1 U7265 ( .A1(n6276), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6271), .ZN(n6256) );
  OAI21_X1 U7266 ( .B1(n6257), .B2(n6273), .A(n6256), .ZN(U2942) );
  AOI22_X1 U7267 ( .A1(n6276), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6271), .ZN(n6258) );
  OAI21_X1 U7268 ( .B1(n6273), .B2(n6259), .A(n6258), .ZN(U2943) );
  AOI22_X1 U7269 ( .A1(n6276), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6271), .ZN(n6260) );
  OAI21_X1 U7270 ( .B1(n6273), .B2(n6261), .A(n6260), .ZN(U2944) );
  AOI22_X1 U7271 ( .A1(n6276), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n6271), .ZN(n6262) );
  OAI21_X1 U7272 ( .B1(n5047), .B2(n6273), .A(n6262), .ZN(U2945) );
  AOI22_X1 U7273 ( .A1(n6276), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6271), .ZN(n6263) );
  OAI21_X1 U7274 ( .B1(n6273), .B2(n6264), .A(n6263), .ZN(U2946) );
  AOI22_X1 U7275 ( .A1(n6276), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n6271), .ZN(n6266) );
  NAND2_X1 U7276 ( .A1(n6266), .A2(n6265), .ZN(U2947) );
  AOI22_X1 U7277 ( .A1(n6276), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n6271), .ZN(n6267) );
  OAI21_X1 U7278 ( .B1(n6273), .B2(n6268), .A(n6267), .ZN(U2948) );
  AOI22_X1 U7279 ( .A1(n6276), .A2(LWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n6271), .ZN(n6269) );
  OAI21_X1 U7280 ( .B1(n6270), .B2(n6273), .A(n6269), .ZN(U2949) );
  AOI22_X1 U7281 ( .A1(n6276), .A2(LWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_11__SCAN_IN), .B2(n6271), .ZN(n6272) );
  OAI21_X1 U7282 ( .B1(n6274), .B2(n6273), .A(n6272), .ZN(U2950) );
  AOI21_X1 U7283 ( .B1(LWORD_REG_13__SCAN_IN), .B2(n6276), .A(n6275), .ZN(
        n6277) );
  OAI21_X1 U7284 ( .B1(n6278), .B2(n6282), .A(n6277), .ZN(U2952) );
  AOI21_X1 U7285 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n6280), .A(n6279), .ZN(
        n6281) );
  OAI21_X1 U7286 ( .B1(n6283), .B2(n6282), .A(n6281), .ZN(U2953) );
  AOI22_X1 U7287 ( .A1(n6284), .A2(REIP_REG_2__SCAN_IN), .B1(n6298), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6291) );
  XNOR2_X1 U7288 ( .A(n6285), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6287)
         );
  XNOR2_X1 U7289 ( .A(n6287), .B(n6286), .ZN(n6335) );
  AOI22_X1 U7290 ( .A1(n6296), .A2(n6335), .B1(n6289), .B2(n6288), .ZN(n6290)
         );
  OAI211_X1 U7291 ( .C1(n5955), .C2(n6292), .A(n6291), .B(n6290), .ZN(U2984)
         );
  INV_X1 U7292 ( .A(n6293), .ZN(n6295) );
  AOI21_X1 U7293 ( .B1(n6296), .B2(n6295), .A(n6294), .ZN(n6300) );
  OAI21_X1 U7294 ( .B1(n6298), .B2(n6297), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n6299) );
  OAI211_X1 U7295 ( .C1(n6302), .C2(n6301), .A(n6300), .B(n6299), .ZN(U2986)
         );
  AOI22_X1 U7296 ( .A1(n6304), .A2(n6336), .B1(n6330), .B2(n6303), .ZN(n6308)
         );
  OAI21_X1 U7297 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6306), .A(n6305), 
        .ZN(n6307) );
  OAI211_X1 U7298 ( .C1(n6668), .C2(n6309), .A(n6308), .B(n6307), .ZN(U3007)
         );
  INV_X1 U7299 ( .A(n6310), .ZN(n6311) );
  AOI21_X1 U7300 ( .B1(n6330), .B2(n6312), .A(n6311), .ZN(n6316) );
  AOI22_X1 U7301 ( .A1(n6314), .A2(n6336), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6313), .ZN(n6315) );
  OAI211_X1 U7302 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6317), .A(n6316), 
        .B(n6315), .ZN(U3009) );
  INV_X1 U7303 ( .A(n6318), .ZN(n6322) );
  NAND2_X1 U7304 ( .A1(n6330), .A2(n6319), .ZN(n6321) );
  OAI211_X1 U7305 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n6322), .A(n6321), 
        .B(n6320), .ZN(n6323) );
  AOI21_X1 U7306 ( .B1(n6324), .B2(n6336), .A(n6323), .ZN(n6325) );
  OAI21_X1 U7307 ( .B1(n6326), .B2(n3475), .A(n6325), .ZN(U3011) );
  INV_X1 U7308 ( .A(n6327), .ZN(n6329) );
  AOI22_X1 U7309 ( .A1(n6330), .A2(n6329), .B1(n6328), .B2(REIP_REG_2__SCAN_IN), .ZN(n6343) );
  NOR2_X1 U7310 ( .A1(n6331), .A2(n6339), .ZN(n6333) );
  OAI221_X1 U7311 ( .B1(n6334), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .C1(n6334), .C2(n6333), .A(n6332), .ZN(n6342) );
  AOI22_X1 U7312 ( .A1(n6337), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6336), 
        .B2(n6335), .ZN(n6341) );
  OR3_X1 U7313 ( .A1(n6339), .A2(n6338), .A3(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6340) );
  NAND4_X1 U7314 ( .A1(n6343), .A2(n6342), .A3(n6341), .A4(n6340), .ZN(U3016)
         );
  NOR2_X1 U7315 ( .A1(n6586), .A2(n6344), .ZN(U3019) );
  NAND3_X1 U7316 ( .A1(n6347), .A2(n6346), .A3(n6345), .ZN(n6348) );
  NAND2_X1 U7317 ( .A1(n6348), .A2(n6389), .ZN(n6355) );
  NOR2_X1 U7318 ( .A1(n6502), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6378)
         );
  AOI21_X1 U7319 ( .B1(n6349), .B2(n6507), .A(n6378), .ZN(n6354) );
  INV_X1 U7320 ( .A(n6354), .ZN(n6350) );
  OAI21_X1 U7321 ( .B1(n6355), .B2(n6350), .A(n6510), .ZN(n6351) );
  AOI22_X1 U7322 ( .A1(n6504), .A2(n6378), .B1(n6503), .B2(n6377), .ZN(n6357)
         );
  OAI22_X1 U7323 ( .A1(n6355), .A2(n6354), .B1(n6353), .B2(n6514), .ZN(n6379)
         );
  AOI22_X1 U7324 ( .A1(n6474), .A2(n6380), .B1(n6518), .B2(n6379), .ZN(n6356)
         );
  OAI211_X1 U7325 ( .C1(n6384), .C2(n6358), .A(n6357), .B(n6356), .ZN(U3044)
         );
  INV_X1 U7326 ( .A(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n6361) );
  AOI22_X1 U7327 ( .A1(n6523), .A2(n6378), .B1(n6435), .B2(n6377), .ZN(n6360)
         );
  AOI22_X1 U7328 ( .A1(n6522), .A2(n6380), .B1(n6524), .B2(n6379), .ZN(n6359)
         );
  OAI211_X1 U7329 ( .C1(n6384), .C2(n6361), .A(n6360), .B(n6359), .ZN(U3045)
         );
  AOI22_X1 U7330 ( .A1(n6529), .A2(n6378), .B1(n6439), .B2(n6377), .ZN(n6363)
         );
  AOI22_X1 U7331 ( .A1(n6528), .A2(n6380), .B1(n6530), .B2(n6379), .ZN(n6362)
         );
  OAI211_X1 U7332 ( .C1(n6384), .C2(n6364), .A(n6363), .B(n6362), .ZN(U3046)
         );
  INV_X1 U7333 ( .A(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n6367) );
  AOI22_X1 U7334 ( .A1(n6535), .A2(n6378), .B1(n6404), .B2(n6377), .ZN(n6366)
         );
  AOI22_X1 U7335 ( .A1(n6534), .A2(n6380), .B1(n6536), .B2(n6379), .ZN(n6365)
         );
  OAI211_X1 U7336 ( .C1(n6384), .C2(n6367), .A(n6366), .B(n6365), .ZN(U3047)
         );
  AOI22_X1 U7337 ( .A1(n6541), .A2(n6378), .B1(n6446), .B2(n6377), .ZN(n6369)
         );
  AOI22_X1 U7338 ( .A1(n6540), .A2(n6380), .B1(n6542), .B2(n6379), .ZN(n6368)
         );
  OAI211_X1 U7339 ( .C1(n6384), .C2(n6370), .A(n6369), .B(n6368), .ZN(U3048)
         );
  INV_X1 U7340 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n6373) );
  AOI22_X1 U7341 ( .A1(n6547), .A2(n6378), .B1(n6546), .B2(n6377), .ZN(n6372)
         );
  AOI22_X1 U7342 ( .A1(n6486), .A2(n6380), .B1(n6548), .B2(n6379), .ZN(n6371)
         );
  OAI211_X1 U7343 ( .C1(n6384), .C2(n6373), .A(n6372), .B(n6371), .ZN(U3049)
         );
  INV_X1 U7344 ( .A(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n6376) );
  AOI22_X1 U7345 ( .A1(n6554), .A2(n6378), .B1(n6412), .B2(n6377), .ZN(n6375)
         );
  AOI22_X1 U7346 ( .A1(n6553), .A2(n6380), .B1(n6555), .B2(n6379), .ZN(n6374)
         );
  OAI211_X1 U7347 ( .C1(n6384), .C2(n6376), .A(n6375), .B(n6374), .ZN(U3050)
         );
  INV_X1 U7348 ( .A(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n6383) );
  AOI22_X1 U7349 ( .A1(n6563), .A2(n6378), .B1(n6560), .B2(n6377), .ZN(n6382)
         );
  AOI22_X1 U7350 ( .A1(n6495), .A2(n6380), .B1(n6565), .B2(n6379), .ZN(n6381)
         );
  OAI211_X1 U7351 ( .C1(n6384), .C2(n6383), .A(n6382), .B(n6381), .ZN(U3051)
         );
  NOR2_X1 U7352 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6430), .ZN(n6417)
         );
  NAND3_X1 U7353 ( .A1(n6468), .A2(n6386), .A3(n6501), .ZN(n6387) );
  OAI21_X1 U7354 ( .B1(n6388), .B2(n6392), .A(n6387), .ZN(n6416) );
  AOI22_X1 U7355 ( .A1(n6504), .A2(n6417), .B1(n6518), .B2(n6416), .ZN(n6399)
         );
  INV_X1 U7356 ( .A(n6418), .ZN(n6390) );
  NAND3_X1 U7357 ( .A1(n6390), .A2(n6389), .A3(n6459), .ZN(n6394) );
  NOR2_X1 U7358 ( .A1(n6392), .A2(n6391), .ZN(n6426) );
  AOI21_X1 U7359 ( .B1(n6394), .B2(n6393), .A(n6426), .ZN(n6396) );
  OAI211_X1 U7360 ( .C1(n6417), .C2(n6716), .A(n6462), .B(n6501), .ZN(n6395)
         );
  AOI22_X1 U7361 ( .A1(n6419), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6503), 
        .B2(n6418), .ZN(n6398) );
  OAI211_X1 U7362 ( .C1(n6521), .C2(n6459), .A(n6399), .B(n6398), .ZN(U3068)
         );
  AOI22_X1 U7363 ( .A1(n6523), .A2(n6417), .B1(n6524), .B2(n6416), .ZN(n6401)
         );
  AOI22_X1 U7364 ( .A1(n6419), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6435), 
        .B2(n6418), .ZN(n6400) );
  OAI211_X1 U7365 ( .C1(n6438), .C2(n6459), .A(n6401), .B(n6400), .ZN(U3069)
         );
  AOI22_X1 U7366 ( .A1(n6529), .A2(n6417), .B1(n6530), .B2(n6416), .ZN(n6403)
         );
  AOI22_X1 U7367 ( .A1(n6419), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6439), 
        .B2(n6418), .ZN(n6402) );
  OAI211_X1 U7368 ( .C1(n6442), .C2(n6459), .A(n6403), .B(n6402), .ZN(U3070)
         );
  AOI22_X1 U7369 ( .A1(n6535), .A2(n6417), .B1(n6536), .B2(n6416), .ZN(n6406)
         );
  AOI22_X1 U7370 ( .A1(n6419), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6404), 
        .B2(n6418), .ZN(n6405) );
  OAI211_X1 U7371 ( .C1(n6407), .C2(n6459), .A(n6406), .B(n6405), .ZN(U3071)
         );
  AOI22_X1 U7372 ( .A1(n6541), .A2(n6417), .B1(n6542), .B2(n6416), .ZN(n6409)
         );
  AOI22_X1 U7373 ( .A1(n6419), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6446), 
        .B2(n6418), .ZN(n6408) );
  OAI211_X1 U7374 ( .C1(n6449), .C2(n6459), .A(n6409), .B(n6408), .ZN(U3072)
         );
  AOI22_X1 U7375 ( .A1(n6547), .A2(n6417), .B1(n6548), .B2(n6416), .ZN(n6411)
         );
  AOI22_X1 U7376 ( .A1(n6419), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6546), 
        .B2(n6418), .ZN(n6410) );
  OAI211_X1 U7377 ( .C1(n6551), .C2(n6459), .A(n6411), .B(n6410), .ZN(U3073)
         );
  AOI22_X1 U7378 ( .A1(n6555), .A2(n6416), .B1(n6554), .B2(n6417), .ZN(n6414)
         );
  AOI22_X1 U7379 ( .A1(n6419), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6412), 
        .B2(n6418), .ZN(n6413) );
  OAI211_X1 U7380 ( .C1(n6415), .C2(n6459), .A(n6414), .B(n6413), .ZN(U3074)
         );
  AOI22_X1 U7381 ( .A1(n6563), .A2(n6417), .B1(n6565), .B2(n6416), .ZN(n6421)
         );
  AOI22_X1 U7382 ( .A1(n6419), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6560), 
        .B2(n6418), .ZN(n6420) );
  OAI211_X1 U7383 ( .C1(n6570), .C2(n6459), .A(n6421), .B(n6420), .ZN(U3075)
         );
  INV_X1 U7384 ( .A(n6422), .ZN(n6454) );
  AOI22_X1 U7385 ( .A1(n6504), .A2(n6454), .B1(n6474), .B2(n6464), .ZN(n6434)
         );
  NAND2_X1 U7386 ( .A1(n6425), .A2(n6513), .ZN(n6432) );
  INV_X1 U7387 ( .A(n6432), .ZN(n6427) );
  AOI21_X1 U7388 ( .B1(n6426), .B2(n6507), .A(n6454), .ZN(n6431) );
  NAND2_X1 U7389 ( .A1(n6427), .A2(n6431), .ZN(n6428) );
  OAI211_X1 U7390 ( .C1(n6513), .C2(n6429), .A(n6428), .B(n6510), .ZN(n6456)
         );
  OAI22_X1 U7391 ( .A1(n6432), .A2(n6431), .B1(n6430), .B2(n6514), .ZN(n6455)
         );
  AOI22_X1 U7392 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6456), .B1(n6518), 
        .B2(n6455), .ZN(n6433) );
  OAI211_X1 U7393 ( .C1(n6477), .C2(n6459), .A(n6434), .B(n6433), .ZN(U3076)
         );
  INV_X1 U7394 ( .A(n6459), .ZN(n6445) );
  AOI22_X1 U7395 ( .A1(n6523), .A2(n6454), .B1(n6435), .B2(n6445), .ZN(n6437)
         );
  AOI22_X1 U7396 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6456), .B1(n6524), 
        .B2(n6455), .ZN(n6436) );
  OAI211_X1 U7397 ( .C1(n6438), .C2(n6499), .A(n6437), .B(n6436), .ZN(U3077)
         );
  AOI22_X1 U7398 ( .A1(n6529), .A2(n6454), .B1(n6439), .B2(n6445), .ZN(n6441)
         );
  AOI22_X1 U7399 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6456), .B1(n6530), 
        .B2(n6455), .ZN(n6440) );
  OAI211_X1 U7400 ( .C1(n6442), .C2(n6499), .A(n6441), .B(n6440), .ZN(U3078)
         );
  AOI22_X1 U7401 ( .A1(n6535), .A2(n6454), .B1(n6534), .B2(n6464), .ZN(n6444)
         );
  AOI22_X1 U7402 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6456), .B1(n6536), 
        .B2(n6455), .ZN(n6443) );
  OAI211_X1 U7403 ( .C1(n6539), .C2(n6459), .A(n6444), .B(n6443), .ZN(U3079)
         );
  AOI22_X1 U7404 ( .A1(n6541), .A2(n6454), .B1(n6446), .B2(n6445), .ZN(n6448)
         );
  AOI22_X1 U7405 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6456), .B1(n6542), 
        .B2(n6455), .ZN(n6447) );
  OAI211_X1 U7406 ( .C1(n6449), .C2(n6499), .A(n6448), .B(n6447), .ZN(U3080)
         );
  AOI22_X1 U7407 ( .A1(n6547), .A2(n6454), .B1(n6486), .B2(n6464), .ZN(n6451)
         );
  AOI22_X1 U7408 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6456), .B1(n6548), 
        .B2(n6455), .ZN(n6450) );
  OAI211_X1 U7409 ( .C1(n6489), .C2(n6459), .A(n6451), .B(n6450), .ZN(U3081)
         );
  AOI22_X1 U7410 ( .A1(n6554), .A2(n6454), .B1(n6553), .B2(n6464), .ZN(n6453)
         );
  AOI22_X1 U7411 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6456), .B1(n6555), 
        .B2(n6455), .ZN(n6452) );
  OAI211_X1 U7412 ( .C1(n6559), .C2(n6459), .A(n6453), .B(n6452), .ZN(U3082)
         );
  AOI22_X1 U7413 ( .A1(n6563), .A2(n6454), .B1(n6495), .B2(n6464), .ZN(n6458)
         );
  AOI22_X1 U7414 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6456), .B1(n6565), 
        .B2(n6455), .ZN(n6457) );
  OAI211_X1 U7415 ( .C1(n6500), .C2(n6459), .A(n6458), .B(n6457), .ZN(U3083)
         );
  NOR2_X1 U7416 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6460), .ZN(n6493)
         );
  OAI22_X1 U7417 ( .A1(n6463), .A2(n6466), .B1(n6462), .B2(n6461), .ZN(n6492)
         );
  AOI22_X1 U7418 ( .A1(n6504), .A2(n6493), .B1(n6518), .B2(n6492), .ZN(n6476)
         );
  OAI21_X1 U7419 ( .B1(n6494), .B2(n6464), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6465) );
  OAI211_X1 U7420 ( .C1(n6467), .C2(n6466), .A(n6465), .B(n6513), .ZN(n6473)
         );
  INV_X1 U7421 ( .A(n6468), .ZN(n6469) );
  OAI21_X1 U7422 ( .B1(n6716), .B2(n6493), .A(n6469), .ZN(n6470) );
  INV_X1 U7423 ( .A(n6470), .ZN(n6471) );
  NAND3_X1 U7424 ( .A1(n6473), .A2(n6472), .A3(n6471), .ZN(n6496) );
  AOI22_X1 U7425 ( .A1(n6496), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6474), 
        .B2(n6494), .ZN(n6475) );
  OAI211_X1 U7426 ( .C1(n6477), .C2(n6499), .A(n6476), .B(n6475), .ZN(U3084)
         );
  AOI22_X1 U7427 ( .A1(n6523), .A2(n6493), .B1(n6524), .B2(n6492), .ZN(n6479)
         );
  AOI22_X1 U7428 ( .A1(n6496), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6522), 
        .B2(n6494), .ZN(n6478) );
  OAI211_X1 U7429 ( .C1(n6527), .C2(n6499), .A(n6479), .B(n6478), .ZN(U3085)
         );
  AOI22_X1 U7430 ( .A1(n6529), .A2(n6493), .B1(n6530), .B2(n6492), .ZN(n6481)
         );
  AOI22_X1 U7431 ( .A1(n6496), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6528), 
        .B2(n6494), .ZN(n6480) );
  OAI211_X1 U7432 ( .C1(n6533), .C2(n6499), .A(n6481), .B(n6480), .ZN(U3086)
         );
  AOI22_X1 U7433 ( .A1(n6535), .A2(n6493), .B1(n6536), .B2(n6492), .ZN(n6483)
         );
  AOI22_X1 U7434 ( .A1(n6496), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6534), 
        .B2(n6494), .ZN(n6482) );
  OAI211_X1 U7435 ( .C1(n6539), .C2(n6499), .A(n6483), .B(n6482), .ZN(U3087)
         );
  AOI22_X1 U7436 ( .A1(n6541), .A2(n6493), .B1(n6542), .B2(n6492), .ZN(n6485)
         );
  AOI22_X1 U7437 ( .A1(n6496), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6540), 
        .B2(n6494), .ZN(n6484) );
  OAI211_X1 U7438 ( .C1(n6545), .C2(n6499), .A(n6485), .B(n6484), .ZN(U3088)
         );
  AOI22_X1 U7439 ( .A1(n6547), .A2(n6493), .B1(n6548), .B2(n6492), .ZN(n6488)
         );
  AOI22_X1 U7440 ( .A1(n6496), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6486), 
        .B2(n6494), .ZN(n6487) );
  OAI211_X1 U7441 ( .C1(n6489), .C2(n6499), .A(n6488), .B(n6487), .ZN(U3089)
         );
  AOI22_X1 U7442 ( .A1(n6555), .A2(n6492), .B1(n6554), .B2(n6493), .ZN(n6491)
         );
  AOI22_X1 U7443 ( .A1(n6496), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6553), 
        .B2(n6494), .ZN(n6490) );
  OAI211_X1 U7444 ( .C1(n6559), .C2(n6499), .A(n6491), .B(n6490), .ZN(U3090)
         );
  AOI22_X1 U7445 ( .A1(n6563), .A2(n6493), .B1(n6565), .B2(n6492), .ZN(n6498)
         );
  AOI22_X1 U7446 ( .A1(n6496), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6495), 
        .B2(n6494), .ZN(n6497) );
  OAI211_X1 U7447 ( .C1(n6500), .C2(n6499), .A(n6498), .B(n6497), .ZN(U3091)
         );
  NOR2_X1 U7448 ( .A1(n6502), .A2(n6501), .ZN(n6562) );
  INV_X1 U7449 ( .A(n6558), .ZN(n6561) );
  AOI22_X1 U7450 ( .A1(n6504), .A2(n6562), .B1(n6561), .B2(n6503), .ZN(n6520)
         );
  INV_X1 U7451 ( .A(n6515), .ZN(n6512) );
  OAI21_X1 U7452 ( .B1(n6506), .B2(n6505), .A(n6513), .ZN(n6517) );
  INV_X1 U7453 ( .A(n6517), .ZN(n6509) );
  AOI21_X1 U7454 ( .B1(n6508), .B2(n6507), .A(n6562), .ZN(n6516) );
  NAND2_X1 U7455 ( .A1(n6509), .A2(n6516), .ZN(n6511) );
  OAI211_X1 U7456 ( .C1(n6513), .C2(n6512), .A(n6511), .B(n6510), .ZN(n6566)
         );
  OAI22_X1 U7457 ( .A1(n6517), .A2(n6516), .B1(n6515), .B2(n6514), .ZN(n6564)
         );
  AOI22_X1 U7458 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6566), .B1(n6518), 
        .B2(n6564), .ZN(n6519) );
  OAI211_X1 U7459 ( .C1(n6521), .C2(n6569), .A(n6520), .B(n6519), .ZN(U3108)
         );
  INV_X1 U7460 ( .A(n6569), .ZN(n6552) );
  AOI22_X1 U7461 ( .A1(n6523), .A2(n6562), .B1(n6522), .B2(n6552), .ZN(n6526)
         );
  AOI22_X1 U7462 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6566), .B1(n6524), 
        .B2(n6564), .ZN(n6525) );
  OAI211_X1 U7463 ( .C1(n6527), .C2(n6558), .A(n6526), .B(n6525), .ZN(U3109)
         );
  AOI22_X1 U7464 ( .A1(n6529), .A2(n6562), .B1(n6528), .B2(n6552), .ZN(n6532)
         );
  AOI22_X1 U7465 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6566), .B1(n6530), 
        .B2(n6564), .ZN(n6531) );
  OAI211_X1 U7466 ( .C1(n6533), .C2(n6558), .A(n6532), .B(n6531), .ZN(U3110)
         );
  AOI22_X1 U7467 ( .A1(n6535), .A2(n6562), .B1(n6534), .B2(n6552), .ZN(n6538)
         );
  AOI22_X1 U7468 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6566), .B1(n6536), 
        .B2(n6564), .ZN(n6537) );
  OAI211_X1 U7469 ( .C1(n6539), .C2(n6558), .A(n6538), .B(n6537), .ZN(U3111)
         );
  AOI22_X1 U7470 ( .A1(n6541), .A2(n6562), .B1(n6540), .B2(n6552), .ZN(n6544)
         );
  AOI22_X1 U7471 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6566), .B1(n6542), 
        .B2(n6564), .ZN(n6543) );
  OAI211_X1 U7472 ( .C1(n6545), .C2(n6558), .A(n6544), .B(n6543), .ZN(U3112)
         );
  AOI22_X1 U7473 ( .A1(n6547), .A2(n6562), .B1(n6561), .B2(n6546), .ZN(n6550)
         );
  AOI22_X1 U7474 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6566), .B1(n6548), 
        .B2(n6564), .ZN(n6549) );
  OAI211_X1 U7475 ( .C1(n6551), .C2(n6569), .A(n6550), .B(n6549), .ZN(U3113)
         );
  AOI22_X1 U7476 ( .A1(n6554), .A2(n6562), .B1(n6553), .B2(n6552), .ZN(n6557)
         );
  AOI22_X1 U7477 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6566), .B1(n6555), 
        .B2(n6564), .ZN(n6556) );
  OAI211_X1 U7478 ( .C1(n6559), .C2(n6558), .A(n6557), .B(n6556), .ZN(U3114)
         );
  AOI22_X1 U7479 ( .A1(n6563), .A2(n6562), .B1(n6561), .B2(n6560), .ZN(n6568)
         );
  AOI22_X1 U7480 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6566), .B1(n6565), 
        .B2(n6564), .ZN(n6567) );
  OAI211_X1 U7481 ( .C1(n6570), .C2(n6569), .A(n6568), .B(n6567), .ZN(U3115)
         );
  OAI211_X1 U7482 ( .C1(n3078), .C2(n6572), .A(n6571), .B(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6576) );
  INV_X1 U7483 ( .A(n6573), .ZN(n6574) );
  OAI21_X1 U7484 ( .B1(n6576), .B2(n6575), .A(n6574), .ZN(n6578) );
  NAND2_X1 U7485 ( .A1(n6576), .A2(n6575), .ZN(n6577) );
  OAI21_X1 U7486 ( .B1(n6579), .B2(n6578), .A(n6577), .ZN(n6580) );
  AOI222_X1 U7487 ( .A1(n6582), .A2(n6581), .B1(n6582), .B2(n6580), .C1(n6581), 
        .C2(n6580), .ZN(n6584) );
  AND2_X1 U7488 ( .A1(n6584), .A2(n6583), .ZN(n6585) );
  OAI22_X1 U7489 ( .A1(n6585), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(n6584), .B2(n6583), .ZN(n6587) );
  NAND2_X1 U7490 ( .A1(n6587), .A2(n6586), .ZN(n6596) );
  OAI21_X1 U7491 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6588), 
        .ZN(n6589) );
  NAND4_X1 U7492 ( .A1(n6592), .A2(n6591), .A3(n6590), .A4(n6589), .ZN(n6593)
         );
  NOR2_X1 U7493 ( .A1(n6594), .A2(n6593), .ZN(n6595) );
  NAND2_X1 U7494 ( .A1(n6596), .A2(n6595), .ZN(n6606) );
  OAI22_X1 U7495 ( .A1(n6606), .A2(n6598), .B1(n6729), .B2(n6597), .ZN(n6602)
         );
  OR2_X1 U7496 ( .A1(n6600), .A2(n6599), .ZN(n6601) );
  OAI21_X1 U7497 ( .B1(n6604), .B2(n6603), .A(n6715), .ZN(n6610) );
  OAI21_X1 U7498 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6729), .A(n6715), .ZN(
        n6617) );
  AOI211_X1 U7499 ( .C1(n6607), .C2(n6606), .A(n6605), .B(n6617), .ZN(n6609)
         );
  OAI221_X1 U7500 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6610), .C1(n6615), .C2(
        n6609), .A(n6608), .ZN(U3148) );
  AND2_X1 U7501 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6611), .ZN(n6613) );
  AOI21_X1 U7502 ( .B1(n6613), .B2(n6729), .A(n6612), .ZN(n6620) );
  NOR2_X1 U7503 ( .A1(n6615), .A2(n6614), .ZN(n6622) );
  AOI21_X1 U7504 ( .B1(n6622), .B2(n6617), .A(n6616), .ZN(n6618) );
  OAI221_X1 U7505 ( .B1(n6621), .B2(n6620), .C1(n6715), .C2(n6619), .A(n6618), 
        .ZN(U3149) );
  AOI21_X1 U7506 ( .B1(n6622), .B2(n6729), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n6624) );
  OAI21_X1 U7507 ( .B1(n6625), .B2(n6624), .A(n6623), .ZN(U3150) );
  AND2_X1 U7508 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6630), .ZN(U3151) );
  AND2_X1 U7509 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6630), .ZN(U3152) );
  AND2_X1 U7510 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6630), .ZN(U3153) );
  NOR2_X1 U7511 ( .A1(n6712), .A2(n6626), .ZN(U3154) );
  AND2_X1 U7512 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6630), .ZN(U3155) );
  AND2_X1 U7513 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6630), .ZN(U3156) );
  AND2_X1 U7514 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6630), .ZN(U3157) );
  AND2_X1 U7515 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6630), .ZN(U3158) );
  AND2_X1 U7516 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6630), .ZN(U3159) );
  AND2_X1 U7517 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6630), .ZN(U3160) );
  AND2_X1 U7518 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6630), .ZN(U3161) );
  AND2_X1 U7519 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6630), .ZN(U3162) );
  AND2_X1 U7520 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6630), .ZN(U3163) );
  AND2_X1 U7521 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6630), .ZN(U3164) );
  AND2_X1 U7522 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6630), .ZN(U3165) );
  AND2_X1 U7523 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6630), .ZN(U3166) );
  AND2_X1 U7524 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6630), .ZN(U3167) );
  AND2_X1 U7525 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6630), .ZN(U3168) );
  AND2_X1 U7526 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6630), .ZN(U3169) );
  AND2_X1 U7527 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6630), .ZN(U3170) );
  AND2_X1 U7528 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6630), .ZN(U3171) );
  AND2_X1 U7529 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6630), .ZN(U3172) );
  AND2_X1 U7530 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6630), .ZN(U3173) );
  AND2_X1 U7531 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6630), .ZN(U3174) );
  NOR2_X1 U7532 ( .A1(n6712), .A2(n6627), .ZN(U3175) );
  AND2_X1 U7533 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6630), .ZN(U3176) );
  NOR2_X1 U7534 ( .A1(n6712), .A2(n6628), .ZN(U3177) );
  AND2_X1 U7535 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6630), .ZN(U3178) );
  NOR2_X1 U7536 ( .A1(n6712), .A2(n6629), .ZN(U3179) );
  AND2_X1 U7537 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6630), .ZN(U3180) );
  NAND2_X1 U7538 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6640) );
  NAND2_X1 U7539 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6635) );
  INV_X1 U7540 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6632) );
  NAND2_X1 U7541 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6637) );
  OAI21_X1 U7542 ( .B1(n6632), .B2(n6729), .A(n6637), .ZN(n6634) );
  OAI221_X1 U7543 ( .B1(n6632), .B2(n6648), .C1(NA_N), .C2(n6648), .A(n6631), 
        .ZN(n6633) );
  INV_X1 U7544 ( .A(n6633), .ZN(n6647) );
  AOI21_X1 U7545 ( .B1(n6635), .B2(n6634), .A(n6647), .ZN(n6636) );
  OAI221_X1 U7546 ( .B1(n6708), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n6708), 
        .C2(n6640), .A(n6636), .ZN(U3181) );
  INV_X1 U7547 ( .A(n6637), .ZN(n6641) );
  NAND2_X1 U7548 ( .A1(STATE_REG_0__SCAN_IN), .A2(REQUESTPENDING_REG_SCAN_IN), 
        .ZN(n6643) );
  AOI21_X1 U7549 ( .B1(STATE_REG_1__SCAN_IN), .B2(READY_N), .A(n6638), .ZN(
        n6639) );
  OAI221_X1 U7550 ( .B1(n6641), .B2(n6643), .C1(n6641), .C2(n6640), .A(n6639), 
        .ZN(U3182) );
  AOI221_X1 U7551 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6729), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6642) );
  OAI21_X1 U7552 ( .B1(STATE_REG_2__SCAN_IN), .B2(n6642), .A(HOLD), .ZN(n6646)
         );
  OAI21_X1 U7553 ( .B1(NA_N), .B2(n6643), .A(n6648), .ZN(n6644) );
  NAND3_X1 U7554 ( .A1(READY_N), .A2(n6644), .A3(STATE_REG_1__SCAN_IN), .ZN(
        n6645) );
  OAI221_X1 U7555 ( .B1(n6647), .B2(n6646), .C1(n6647), .C2(
        STATE_REG_0__SCAN_IN), .A(n6645), .ZN(U3183) );
  NOR2_X2 U7556 ( .A1(n6648), .A2(n6740), .ZN(n6700) );
  NAND2_X1 U7557 ( .A1(n6648), .A2(n6708), .ZN(n6706) );
  INV_X1 U7558 ( .A(n6706), .ZN(n6689) );
  AOI22_X1 U7559 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6689), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6726), .ZN(n6649) );
  OAI21_X1 U7560 ( .B1(n6717), .B2(n6702), .A(n6649), .ZN(U3184) );
  AOI22_X1 U7561 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6726), .ZN(n6650) );
  OAI21_X1 U7562 ( .B1(n6652), .B2(n6706), .A(n6650), .ZN(U3185) );
  OAI222_X1 U7563 ( .A1(n6702), .A2(n6652), .B1(n6651), .B2(n6708), .C1(n6654), 
        .C2(n6706), .ZN(U3186) );
  AOI22_X1 U7564 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6689), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6726), .ZN(n6653) );
  OAI21_X1 U7565 ( .B1(n6654), .B2(n6702), .A(n6653), .ZN(U3187) );
  OAI222_X1 U7566 ( .A1(n6706), .A2(n6658), .B1(n6656), .B2(n6708), .C1(n6655), 
        .C2(n6702), .ZN(U3188) );
  AOI22_X1 U7567 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6689), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6726), .ZN(n6657) );
  OAI21_X1 U7568 ( .B1(n6658), .B2(n6702), .A(n6657), .ZN(U3189) );
  AOI22_X1 U7569 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6740), .ZN(n6659) );
  OAI21_X1 U7570 ( .B1(n6661), .B2(n6706), .A(n6659), .ZN(U3190) );
  AOI22_X1 U7571 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6689), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6726), .ZN(n6660) );
  OAI21_X1 U7572 ( .B1(n6661), .B2(n6702), .A(n6660), .ZN(U3191) );
  OAI222_X1 U7573 ( .A1(n6702), .A2(n6664), .B1(n6663), .B2(n6708), .C1(n6662), 
        .C2(n6706), .ZN(U3192) );
  AOI22_X1 U7574 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6726), .ZN(n6665) );
  OAI21_X1 U7575 ( .B1(n6668), .B2(n6706), .A(n6665), .ZN(U3193) );
  OAI222_X1 U7576 ( .A1(n6702), .A2(n6668), .B1(n6667), .B2(n6708), .C1(n6666), 
        .C2(n6706), .ZN(U3194) );
  AOI22_X1 U7577 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6726), .ZN(n6669) );
  OAI21_X1 U7578 ( .B1(n6670), .B2(n6706), .A(n6669), .ZN(U3195) );
  AOI22_X1 U7579 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6726), .ZN(n6671) );
  OAI21_X1 U7580 ( .B1(n6672), .B2(n6706), .A(n6671), .ZN(U3196) );
  OAI222_X1 U7581 ( .A1(n6706), .A2(n6675), .B1(n6673), .B2(n6708), .C1(n6672), 
        .C2(n6702), .ZN(U3197) );
  INV_X1 U7582 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6677) );
  OAI222_X1 U7583 ( .A1(n6702), .A2(n6675), .B1(n6674), .B2(n6708), .C1(n6677), 
        .C2(n6706), .ZN(U3198) );
  AOI22_X1 U7584 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6689), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6726), .ZN(n6676) );
  OAI21_X1 U7585 ( .B1(n6677), .B2(n6702), .A(n6676), .ZN(U3199) );
  AOI22_X1 U7586 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6726), .ZN(n6678) );
  OAI21_X1 U7587 ( .B1(n6680), .B2(n6706), .A(n6678), .ZN(U3200) );
  AOI22_X1 U7588 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6689), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6726), .ZN(n6679) );
  OAI21_X1 U7589 ( .B1(n6680), .B2(n6702), .A(n6679), .ZN(U3201) );
  AOI22_X1 U7590 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6726), .ZN(n6681) );
  OAI21_X1 U7591 ( .B1(n6683), .B2(n6706), .A(n6681), .ZN(U3202) );
  AOI22_X1 U7592 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6689), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6726), .ZN(n6682) );
  OAI21_X1 U7593 ( .B1(n6683), .B2(n6702), .A(n6682), .ZN(U3203) );
  AOI22_X1 U7594 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6726), .ZN(n6684) );
  OAI21_X1 U7595 ( .B1(n6685), .B2(n6706), .A(n6684), .ZN(U3204) );
  AOI22_X1 U7596 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6726), .ZN(n6686) );
  OAI21_X1 U7597 ( .B1(n6688), .B2(n6706), .A(n6686), .ZN(U3205) );
  AOI22_X1 U7598 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6689), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6726), .ZN(n6687) );
  OAI21_X1 U7599 ( .B1(n6688), .B2(n6702), .A(n6687), .ZN(U3206) );
  AOI22_X1 U7600 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6689), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6740), .ZN(n6690) );
  OAI21_X1 U7601 ( .B1(n6691), .B2(n6702), .A(n6690), .ZN(U3207) );
  AOI22_X1 U7602 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6740), .ZN(n6692) );
  OAI21_X1 U7603 ( .B1(n6693), .B2(n6706), .A(n6692), .ZN(U3208) );
  AOI22_X1 U7604 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6740), .ZN(n6694) );
  OAI21_X1 U7605 ( .B1(n6695), .B2(n6706), .A(n6694), .ZN(U3209) );
  AOI22_X1 U7606 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6740), .ZN(n6696) );
  OAI21_X1 U7607 ( .B1(n6697), .B2(n6706), .A(n6696), .ZN(U3210) );
  AOI22_X1 U7608 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6740), .ZN(n6698) );
  OAI21_X1 U7609 ( .B1(n6699), .B2(n6706), .A(n6698), .ZN(U3211) );
  AOI22_X1 U7610 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6700), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6740), .ZN(n6701) );
  OAI21_X1 U7611 ( .B1(n6703), .B2(n6706), .A(n6701), .ZN(U3212) );
  OAI222_X1 U7612 ( .A1(n6706), .A2(n6705), .B1(n6704), .B2(n6708), .C1(n6703), 
        .C2(n6702), .ZN(U3213) );
  MUX2_X1 U7613 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6740), .Z(U3445) );
  MUX2_X1 U7614 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6740), .Z(U3446) );
  MUX2_X1 U7615 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6740), .Z(U3447) );
  INV_X1 U7616 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6723) );
  AOI22_X1 U7617 ( .A1(n6708), .A2(n6723), .B1(n6707), .B2(n6740), .ZN(U3448)
         );
  OAI21_X1 U7618 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6712), .A(n6710), .ZN(
        n6709) );
  INV_X1 U7619 ( .A(n6709), .ZN(U3451) );
  OAI21_X1 U7620 ( .B1(n6712), .B2(n6711), .A(n6710), .ZN(U3452) );
  OAI211_X1 U7621 ( .C1(n6716), .C2(n6715), .A(n6714), .B(n6713), .ZN(U3453)
         );
  AOI21_X1 U7622 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6718) );
  AOI22_X1 U7623 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6718), .B2(n6717), .ZN(n6721) );
  INV_X1 U7624 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6720) );
  AOI22_X1 U7625 ( .A1(n6724), .A2(n6721), .B1(n6720), .B2(n6719), .ZN(U3468)
         );
  OAI21_X1 U7626 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6724), .ZN(n6722) );
  OAI21_X1 U7627 ( .B1(n6724), .B2(n6723), .A(n6722), .ZN(U3469) );
  NAND2_X1 U7628 ( .A1(n6726), .A2(W_R_N_REG_SCAN_IN), .ZN(n6725) );
  OAI21_X1 U7629 ( .B1(n6726), .B2(READREQUEST_REG_SCAN_IN), .A(n6725), .ZN(
        U3470) );
  AOI211_X1 U7630 ( .C1(n6730), .C2(n6729), .A(n6728), .B(n6727), .ZN(n6739)
         );
  INV_X1 U7631 ( .A(n6731), .ZN(n6734) );
  INV_X1 U7632 ( .A(n6732), .ZN(n6733) );
  OAI211_X1 U7633 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6734), .A(n6733), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6736) );
  AOI21_X1 U7634 ( .B1(n6736), .B2(STATE2_REG_0__SCAN_IN), .A(n6735), .ZN(
        n6738) );
  NAND2_X1 U7635 ( .A1(n6739), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6737) );
  OAI21_X1 U7636 ( .B1(n6739), .B2(n6738), .A(n6737), .ZN(U3472) );
  MUX2_X1 U7637 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6740), .Z(U3473) );
  CLKBUF_X1 U3422 ( .A(n4223), .Z(n3229) );
  CLKBUF_X1 U3428 ( .A(n3339), .Z(n3250) );
  CLKBUF_X1 U3436 ( .A(n3133), .Z(n3823) );
  CLKBUF_X1 U3439 ( .A(n3247), .Z(n4132) );
  CLKBUF_X1 U3444 ( .A(n3212), .Z(n3969) );
  CLKBUF_X1 U34450 ( .A(n3334), .Z(n3248) );
  CLKBUF_X1 U3554 ( .A(n4223), .Z(n3242) );
  CLKBUF_X1 U3569 ( .A(n3189), .Z(n3192) );
  INV_X1 U3845 ( .A(n3519), .ZN(n4451) );
  CLKBUF_X1 U4195 ( .A(n3198), .Z(n4755) );
  CLKBUF_X1 U4197 ( .A(n5598), .Z(n5599) );
  CLKBUF_X1 U4210 ( .A(n4661), .Z(n2977) );
endmodule

