

module b14_C_SARLock_k_128_8 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943;

  AND2_X1 U2413 ( .A1(n3052), .A2(n3003), .ZN(n2885) );
  CLKBUF_X1 U2414 ( .A(n4943), .Z(U4043) );
  NOR2_X1 U2415 ( .A1(n3052), .A2(n4510), .ZN(n4943) );
  INV_X1 U2416 ( .A(n2885), .ZN(n2872) );
  INV_X1 U2417 ( .A(n2875), .ZN(n2891) );
  INV_X1 U2418 ( .A(n2539), .ZN(n2492) );
  INV_X1 U2419 ( .A(IR_REG_31__SCAN_IN), .ZN(n2768) );
  CLKBUF_X3 U2420 ( .A(n2507), .Z(n2856) );
  AND2_X4 U2421 ( .A1(n2453), .A2(n2452), .ZN(n2506) );
  CLKBUF_X3 U2422 ( .A(n2539), .Z(n2171) );
  NAND2_X1 U2423 ( .A1(n4312), .A2(n2452), .ZN(n2539) );
  CLKBUF_X2 U2424 ( .A(n2533), .Z(n2890) );
  NOR2_X1 U2425 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2247)
         );
  AOI21_X1 U2426 ( .B1(n2373), .B2(n2257), .A(n4584), .ZN(n2256) );
  NAND3_X1 U2427 ( .A1(n2362), .A2(n2361), .A3(n2368), .ZN(n3903) );
  NAND2_X1 U2428 ( .A1(n3002), .A2(n3001), .ZN(n3515) );
  NAND2_X1 U2429 ( .A1(n4480), .A2(n3228), .ZN(n3661) );
  INV_X1 U2430 ( .A(n3213), .ZN(n4480) );
  INV_X1 U2431 ( .A(n3347), .ZN(n3818) );
  AND4_X1 U2432 ( .A1(n2586), .A2(n2585), .A3(n2584), .A4(n2583), .ZN(n3347)
         );
  NAND4_X1 U2433 ( .A1(n2457), .A2(n2456), .A3(n2455), .A4(n2454), .ZN(n3824)
         );
  NAND4_X1 U2434 ( .A1(n2525), .A2(n2524), .A3(n2523), .A4(n2522), .ZN(n3821)
         );
  CLKBUF_X3 U2435 ( .A(n2521), .Z(n3712) );
  INV_X2 U2436 ( .A(n2533), .ZN(n2873) );
  NAND2_X1 U2437 ( .A1(n2450), .A2(n2449), .ZN(n2452) );
  XNOR2_X1 U2438 ( .A(n2447), .B(n2446), .ZN(n2453) );
  NAND2_X1 U2439 ( .A1(n2449), .A2(IR_REG_31__SCAN_IN), .ZN(n2447) );
  NAND3_X2 U2440 ( .A1(n2479), .A2(n2478), .A3(n2477), .ZN(n3716) );
  AND2_X1 U2441 ( .A1(n2430), .A2(n2497), .ZN(n2234) );
  AND2_X1 U2442 ( .A1(n2245), .A2(n2248), .ZN(n2232) );
  INV_X1 U2443 ( .A(n2498), .ZN(n2497) );
  AND3_X1 U2444 ( .A1(n2247), .A2(n2246), .A3(n2433), .ZN(n2245) );
  AND2_X1 U2445 ( .A1(n2435), .A2(n2624), .ZN(n2248) );
  AND4_X1 U2446 ( .A1(n2747), .A2(n2693), .A3(n2436), .A4(n2746), .ZN(n2437)
         );
  NAND2_X1 U2447 ( .A1(n2210), .A2(n2209), .ZN(n2498) );
  NOR2_X1 U2448 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2246)
         );
  NOR2_X1 U2449 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2624)
         );
  NOR2_X1 U2450 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2435)
         );
  INV_X1 U2451 ( .A(IR_REG_3__SCAN_IN), .ZN(n2527) );
  INV_X1 U2452 ( .A(IR_REG_2__SCAN_IN), .ZN(n2433) );
  INV_X1 U2453 ( .A(IR_REG_0__SCAN_IN), .ZN(n2210) );
  INV_X1 U2454 ( .A(IR_REG_1__SCAN_IN), .ZN(n2209) );
  OR2_X1 U2455 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_22__SCAN_IN), .ZN(n2441)
         );
  NOR2_X1 U2456 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2747)
         );
  INV_X1 U2457 ( .A(IR_REG_16__SCAN_IN), .ZN(n2746) );
  OR2_X1 U2458 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2173)
         );
  OAI22_X2 U2459 ( .A1(n3343), .A2(n2972), .B1(n3345), .B2(n3817), .ZN(n3371)
         );
  OAI21_X2 U2460 ( .B1(n3326), .B2(n2971), .A(n2970), .ZN(n3343) );
  INV_X2 U2461 ( .A(n2888), .ZN(n2862) );
  NAND2_X1 U2462 ( .A1(n2232), .A2(n2234), .ZN(n2237) );
  INV_X1 U2463 ( .A(IR_REG_13__SCAN_IN), .ZN(n2693) );
  AND2_X1 U2464 ( .A1(n3003), .A2(n2934), .ZN(n2888) );
  AOI21_X1 U2465 ( .B1(n2382), .B2(n2379), .A(n2378), .ZN(n2377) );
  NAND2_X1 U2466 ( .A1(n2382), .A2(n2381), .ZN(n2380) );
  NOR2_X1 U2467 ( .A1(n3810), .A2(n3592), .ZN(n2378) );
  AND2_X1 U2468 ( .A1(n3735), .A2(n2284), .ZN(n2283) );
  NOR2_X1 U2469 ( .A1(n3730), .A2(n2285), .ZN(n2284) );
  INV_X1 U2470 ( .A(n2286), .ZN(n2285) );
  NAND2_X1 U2471 ( .A1(n4318), .A2(n2927), .ZN(n3003) );
  NAND2_X1 U2472 ( .A1(n3652), .A2(n3655), .ZN(n3005) );
  AND2_X1 U2473 ( .A1(n2427), .A2(n2439), .ZN(n2426) );
  NOR3_X1 U2474 ( .A1(n2173), .A2(IR_REG_25__SCAN_IN), .A3(n2441), .ZN(n2427)
         );
  NAND2_X1 U2475 ( .A1(n2437), .A2(n2438), .ZN(n2235) );
  NOR2_X1 U2476 ( .A1(n2420), .A2(n2242), .ZN(n2241) );
  INV_X1 U2477 ( .A(n2596), .ZN(n2242) );
  INV_X1 U2478 ( .A(n2421), .ZN(n2420) );
  NAND2_X1 U2479 ( .A1(n2193), .A2(n2221), .ZN(n2220) );
  NAND2_X1 U2480 ( .A1(n3628), .A2(n2222), .ZN(n2221) );
  OAI21_X1 U2481 ( .B1(n3607), .B2(n2412), .A(n2402), .ZN(n3584) );
  OAI22_X1 U2482 ( .A1(n3213), .A2(n2873), .B1(n2872), .B2(n3228), .ZN(n2546)
         );
  AOI22_X1 U2483 ( .A1(n2409), .A2(n2403), .B1(n2402), .B2(n2412), .ZN(n2401)
         );
  NAND2_X1 U2484 ( .A1(n3884), .A2(n4855), .ZN(n2298) );
  NOR2_X1 U2485 ( .A1(n4447), .A2(n4448), .ZN(n4446) );
  INV_X1 U2486 ( .A(n2384), .ZN(n2383) );
  OAI21_X1 U2487 ( .B1(n4023), .B2(n2385), .A(n2178), .ZN(n2384) );
  NAND2_X1 U2488 ( .A1(n2357), .A2(n2356), .ZN(n4056) );
  AOI21_X1 U2489 ( .B1(n2358), .B2(n2360), .A(n2180), .ZN(n2356) );
  OR2_X1 U2490 ( .A1(n3516), .A2(n3043), .ZN(n4179) );
  NAND2_X1 U2491 ( .A1(n3924), .A2(n3517), .ZN(n3516) );
  AND2_X1 U2492 ( .A1(n3940), .A2(n3926), .ZN(n3924) );
  OR2_X1 U2493 ( .A1(n4317), .A2(n4502), .ZN(n4253) );
  AND2_X1 U2494 ( .A1(n3256), .A2(n3255), .ZN(n4553) );
  MUX2_X1 U2495 ( .A(IR_REG_31__SCAN_IN), .B(n2448), .S(IR_REG_29__SCAN_IN), 
        .Z(n2450) );
  NAND2_X1 U2496 ( .A1(n2932), .A2(IR_REG_31__SCAN_IN), .ZN(n2448) );
  NAND2_X1 U2497 ( .A1(n2397), .A2(n2396), .ZN(n3307) );
  NAND2_X1 U2498 ( .A1(n2393), .A2(n2392), .ZN(n2396) );
  INV_X1 U2499 ( .A(n2398), .ZN(n2392) );
  NOR2_X1 U2500 ( .A1(n3889), .A2(n3890), .ZN(n4454) );
  NAND2_X1 U2501 ( .A1(n4454), .A2(n4455), .ZN(n4452) );
  NAND2_X1 U2502 ( .A1(n2489), .A2(n2488), .ZN(n3898) );
  NAND2_X1 U2503 ( .A1(n2251), .A2(n4497), .ZN(n2250) );
  INV_X1 U2504 ( .A(n2369), .ZN(n2368) );
  OR2_X1 U2505 ( .A1(n3515), .A2(n2371), .ZN(n2362) );
  INV_X1 U2506 ( .A(n2283), .ZN(n2280) );
  NAND2_X1 U2507 ( .A1(n2283), .A2(n2278), .ZN(n2277) );
  INV_X1 U2508 ( .A(n2281), .ZN(n2278) );
  INV_X1 U2509 ( .A(n3729), .ZN(n2282) );
  NAND2_X1 U2510 ( .A1(n2414), .A2(n2411), .ZN(n2410) );
  INV_X1 U2511 ( .A(n2843), .ZN(n2411) );
  AND2_X1 U2512 ( .A1(n3576), .A2(n2229), .ZN(n2228) );
  NAND2_X1 U2513 ( .A1(n2230), .A2(n3640), .ZN(n2229) );
  NOR2_X1 U2514 ( .A1(n2230), .A2(n3640), .ZN(n2231) );
  NAND2_X1 U2515 ( .A1(n2407), .A2(n2406), .ZN(n2405) );
  INV_X1 U2516 ( .A(n3587), .ZN(n2406) );
  OAI22_X1 U2517 ( .A1(n2701), .A2(n2423), .B1(n2424), .B2(n2196), .ZN(n2734)
         );
  AND2_X1 U2518 ( .A1(n2424), .A2(n2190), .ZN(n2423) );
  INV_X1 U2519 ( .A(n2425), .ZN(n2424) );
  NAND2_X1 U2520 ( .A1(n4577), .A2(n2885), .ZN(n2875) );
  INV_X1 U2521 ( .A(n2992), .ZN(n2360) );
  NAND2_X1 U2522 ( .A1(n2198), .A2(n3696), .ZN(n2286) );
  NAND2_X1 U2523 ( .A1(n3779), .A2(n3671), .ZN(n2289) );
  AND2_X1 U2524 ( .A1(n3696), .A2(n3671), .ZN(n2281) );
  NAND2_X1 U2525 ( .A1(n4460), .A2(n3687), .ZN(n3425) );
  NOR2_X1 U2526 ( .A1(n2975), .A2(n2352), .ZN(n2351) );
  INV_X1 U2527 ( .A(n4459), .ZN(n2352) );
  OAI21_X1 U2528 ( .B1(n3344), .B2(n2261), .A(n2258), .ZN(n3375) );
  AOI21_X1 U2529 ( .B1(n2262), .B2(n2260), .A(n2259), .ZN(n2258) );
  INV_X1 U2530 ( .A(n2262), .ZN(n2261) );
  INV_X1 U2531 ( .A(n3668), .ZN(n2259) );
  NAND2_X1 U2532 ( .A1(n2266), .A2(n3675), .ZN(n2265) );
  NAND2_X1 U2533 ( .A1(n2272), .A2(n3009), .ZN(n2266) );
  NAND2_X1 U2534 ( .A1(n3914), .A2(n3710), .ZN(n3520) );
  INV_X1 U2535 ( .A(n3054), .ZN(n2910) );
  NOR2_X1 U2536 ( .A1(n2174), .A2(IR_REG_26__SCAN_IN), .ZN(n2386) );
  INV_X1 U2537 ( .A(IR_REG_28__SCAN_IN), .ZN(n2445) );
  AND2_X1 U2538 ( .A1(n2245), .A2(n2236), .ZN(n2233) );
  AND2_X1 U2539 ( .A1(n2439), .A2(n2438), .ZN(n2236) );
  INV_X1 U2540 ( .A(n2526), .ZN(n2249) );
  NOR2_X1 U2541 ( .A1(n3237), .A2(n3238), .ZN(n2398) );
  OR2_X1 U2542 ( .A1(n3455), .A2(n3452), .ZN(n2701) );
  NAND2_X1 U2543 ( .A1(n2416), .A2(n2415), .ZN(n2414) );
  INV_X1 U2544 ( .A(n3541), .ZN(n2415) );
  INV_X1 U2545 ( .A(n3542), .ZN(n2416) );
  NOR2_X1 U2546 ( .A1(n3232), .A2(n2215), .ZN(n2214) );
  INV_X1 U2547 ( .A(n2537), .ZN(n2215) );
  NAND2_X1 U2548 ( .A1(n2417), .A2(n2421), .ZN(n3405) );
  NAND2_X1 U2549 ( .A1(n3333), .A2(n3334), .ZN(n2417) );
  XNOR2_X1 U2550 ( .A(n2501), .B(n2888), .ZN(n2502) );
  OAI22_X1 U2551 ( .A1(n2875), .A2(n4501), .B1(n2873), .B2(n3097), .ZN(n2503)
         );
  AND2_X1 U2552 ( .A1(n2861), .A2(n2860), .ZN(n3790) );
  AND4_X1 U2553 ( .A1(n2670), .A2(n2669), .A3(n2668), .A4(n2667), .ZN(n3016)
         );
  AOI22_X1 U2554 ( .A1(n3170), .A2(REG2_REG_3__SCAN_IN), .B1(n4324), .B2(n3169), .ZN(n3284) );
  NAND2_X1 U2555 ( .A1(n4338), .A2(n3286), .ZN(n3287) );
  NAND2_X1 U2556 ( .A1(n2331), .A2(n2330), .ZN(n2329) );
  NAND2_X1 U2557 ( .A1(n3281), .A2(REG1_REG_5__SCAN_IN), .ZN(n2330) );
  INV_X1 U2558 ( .A(n4333), .ZN(n2331) );
  NAND2_X1 U2559 ( .A1(n4396), .A2(n4397), .ZN(n4395) );
  NAND2_X1 U2560 ( .A1(n4395), .A2(n2324), .ZN(n3274) );
  NAND2_X1 U2561 ( .A1(n3278), .A2(REG1_REG_11__SCAN_IN), .ZN(n2324) );
  NAND2_X1 U2562 ( .A1(n2327), .A2(n2202), .ZN(n3862) );
  NAND2_X1 U2563 ( .A1(n3859), .A2(n2328), .ZN(n2327) );
  NAND2_X1 U2564 ( .A1(n4430), .A2(n2332), .ZN(n3864) );
  NAND2_X1 U2565 ( .A1(n3877), .A2(REG1_REG_15__SCAN_IN), .ZN(n2332) );
  INV_X1 U2566 ( .A(IR_REG_19__SCAN_IN), .ZN(n2486) );
  OR2_X1 U2567 ( .A1(n2854), .A2(n4810), .ZN(n2878) );
  AOI21_X1 U2568 ( .B1(n2383), .B2(n2385), .A(n2185), .ZN(n2382) );
  AND2_X1 U2569 ( .A1(n4040), .A2(n2997), .ZN(n2385) );
  NAND2_X1 U2570 ( .A1(n2991), .A2(n2990), .ZN(n4108) );
  NAND2_X1 U2571 ( .A1(n2651), .A2(REG3_REG_11__SCAN_IN), .ZN(n2664) );
  INV_X1 U2572 ( .A(n3099), .ZN(n2343) );
  AND2_X1 U2573 ( .A1(n2244), .A2(n3763), .ZN(n4494) );
  INV_X1 U2574 ( .A(n4317), .ZN(n2244) );
  AND2_X1 U2575 ( .A1(n4028), .A2(n2205), .ZN(n3940) );
  AND2_X1 U2576 ( .A1(n4024), .A2(n4023), .ZN(n4212) );
  NAND2_X1 U2577 ( .A1(n4124), .A2(n2177), .ZN(n4224) );
  NAND2_X1 U2578 ( .A1(n4124), .A2(n2322), .ZN(n4093) );
  NOR2_X1 U2579 ( .A1(n4240), .A2(n3042), .ZN(n4124) );
  NAND2_X1 U2580 ( .A1(n4494), .A2(n2927), .ZN(n4577) );
  AND2_X1 U2581 ( .A1(n2426), .A2(n2443), .ZN(n2300) );
  NAND2_X1 U2582 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_25__SCAN_IN), .ZN(n2459) );
  NAND2_X1 U2583 ( .A1(n2213), .A2(n2212), .ZN(n2482) );
  INV_X1 U2584 ( .A(IR_REG_21__SCAN_IN), .ZN(n2212) );
  INV_X1 U2585 ( .A(n2470), .ZN(n2213) );
  NOR2_X1 U2586 ( .A1(n2557), .A2(IR_REG_5__SCAN_IN), .ZN(n2626) );
  NAND3_X1 U2587 ( .A1(n4315), .A2(n3058), .A3(n4316), .ZN(n3052) );
  OAI21_X1 U2588 ( .B1(n3307), .B2(n2240), .A(n2183), .ZN(n3406) );
  INV_X1 U2589 ( .A(n2241), .ZN(n2240) );
  AOI21_X1 U2590 ( .B1(n2421), .B2(n2419), .A(n2175), .ZN(n2418) );
  INV_X1 U2591 ( .A(n2220), .ZN(n2219) );
  AOI21_X1 U2592 ( .B1(n2224), .B2(n2220), .A(n2218), .ZN(n2217) );
  INV_X1 U2593 ( .A(n3532), .ZN(n2218) );
  INV_X1 U2594 ( .A(n3136), .ZN(n3097) );
  XNOR2_X1 U2595 ( .A(n2502), .B(n2503), .ZN(n3092) );
  AND4_X1 U2596 ( .A1(n2543), .A2(n2542), .A3(n2541), .A4(n2540), .ZN(n3213)
         );
  OAI21_X1 U2597 ( .B1(n3607), .B2(n2409), .A(n2407), .ZN(n3586) );
  OR2_X1 U2598 ( .A1(n2947), .A2(n2946), .ZN(n3620) );
  INV_X1 U2599 ( .A(n3154), .ZN(n2389) );
  INV_X1 U2600 ( .A(n3153), .ZN(n2390) );
  NAND4_X1 U2601 ( .A1(n2779), .A2(n2778), .A3(n2777), .A4(n2776), .ZN(n4102)
         );
  XNOR2_X1 U2602 ( .A(n2329), .B(n4525), .ZN(n4345) );
  XNOR2_X1 U2603 ( .A(n3864), .B(n3878), .ZN(n4440) );
  NOR2_X1 U2604 ( .A1(n4440), .A2(REG1_REG_16__SCAN_IN), .ZN(n4441) );
  AND2_X1 U2605 ( .A1(n3826), .A2(n3164), .ZN(n4453) );
  NAND2_X1 U2606 ( .A1(n4452), .A2(n2207), .ZN(n2326) );
  XNOR2_X1 U2607 ( .A(n2297), .B(n3895), .ZN(n3900) );
  NOR2_X1 U2608 ( .A1(n4446), .A2(n2206), .ZN(n2297) );
  AND2_X1 U2609 ( .A1(n3826), .A2(n3804), .ZN(n4407) );
  NAND2_X1 U2610 ( .A1(n4553), .A2(n2197), .ZN(n4572) );
  OAI21_X1 U2611 ( .B1(n3045), .B2(n3044), .A(n4179), .ZN(n3906) );
  AND2_X1 U2612 ( .A1(n2364), .A2(n2372), .ZN(n2363) );
  OR2_X1 U2613 ( .A1(n3908), .A2(n2365), .ZN(n2364) );
  NAND2_X1 U2614 ( .A1(n4604), .A2(n2366), .ZN(n2365) );
  NAND2_X1 U2615 ( .A1(n3903), .A2(n4561), .ZN(n2257) );
  NOR2_X1 U2616 ( .A1(n3672), .A2(n2263), .ZN(n2262) );
  INV_X1 U2617 ( .A(n3678), .ZN(n2263) );
  INV_X1 U2618 ( .A(n3667), .ZN(n2260) );
  INV_X1 U2619 ( .A(IR_REG_18__SCAN_IN), .ZN(n2438) );
  NOR2_X1 U2620 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2439)
         );
  NAND2_X1 U2621 ( .A1(n2410), .A2(n2842), .ZN(n2404) );
  INV_X1 U2622 ( .A(n2405), .ZN(n2403) );
  INV_X1 U2623 ( .A(n2404), .ZN(n2402) );
  OR2_X1 U2624 ( .A1(n3608), .A2(n2843), .ZN(n2412) );
  NAND2_X1 U2625 ( .A1(n4398), .A2(n3296), .ZN(n3298) );
  INV_X1 U2626 ( .A(n3861), .ZN(n2328) );
  INV_X1 U2627 ( .A(n3299), .ZN(n2294) );
  INV_X1 U2628 ( .A(n2998), .ZN(n2381) );
  NOR2_X1 U2629 ( .A1(n2383), .A2(n2998), .ZN(n2379) );
  AND2_X1 U2630 ( .A1(n2279), .A2(n2176), .ZN(n3971) );
  OR2_X1 U2631 ( .A1(n3505), .A2(n2280), .ZN(n2279) );
  INV_X1 U2632 ( .A(n3733), .ZN(n2276) );
  OR2_X1 U2633 ( .A1(n4038), .A2(n4037), .ZN(n4035) );
  INV_X1 U2634 ( .A(n2359), .ZN(n2358) );
  OAI21_X1 U2635 ( .B1(n2990), .B2(n2360), .A(n2993), .ZN(n2359) );
  INV_X1 U2636 ( .A(n4158), .ZN(n2982) );
  NAND2_X1 U2637 ( .A1(n3156), .A2(n4488), .ZN(n2303) );
  NAND2_X1 U2638 ( .A1(n3650), .A2(n3651), .ZN(n2334) );
  NAND2_X1 U2639 ( .A1(n3913), .A2(n3521), .ZN(n2375) );
  AND2_X1 U2640 ( .A1(n3954), .A2(n2320), .ZN(n2319) );
  AND2_X1 U2641 ( .A1(n4006), .A2(n3980), .ZN(n2320) );
  NOR2_X1 U2642 ( .A1(n4101), .A2(n4091), .ZN(n2322) );
  INV_X1 U2643 ( .A(n4936), .ZN(n3042) );
  NAND2_X1 U2644 ( .A1(n2288), .A2(n3671), .ZN(n4135) );
  OR2_X1 U2645 ( .A1(n3505), .A2(n3779), .ZN(n2288) );
  NAND2_X1 U2646 ( .A1(n2307), .A2(n3644), .ZN(n2306) );
  INV_X1 U2647 ( .A(n2308), .ZN(n2307) );
  NAND2_X1 U2648 ( .A1(n3498), .A2(n3472), .ZN(n2308) );
  NOR2_X1 U2649 ( .A1(n2303), .A2(n3180), .ZN(n2301) );
  INV_X1 U2650 ( .A(n3138), .ZN(n2304) );
  INV_X1 U2651 ( .A(IR_REG_23__SCAN_IN), .ZN(n2912) );
  OR2_X1 U2652 ( .A1(n2749), .A2(IR_REG_14__SCAN_IN), .ZN(n2716) );
  OR2_X1 U2653 ( .A1(n2658), .A2(IR_REG_10__SCAN_IN), .ZN(n2659) );
  INV_X1 U2654 ( .A(IR_REG_11__SCAN_IN), .ZN(n4763) );
  NOR2_X1 U2655 ( .A1(n2395), .A2(n2398), .ZN(n2394) );
  NAND2_X1 U2656 ( .A1(n2399), .A2(n2567), .ZN(n2393) );
  AND2_X1 U2657 ( .A1(n2422), .A2(n3389), .ZN(n2421) );
  NAND2_X1 U2658 ( .A1(n2241), .A2(n2239), .ZN(n2238) );
  INV_X1 U2659 ( .A(n3306), .ZN(n2239) );
  XNOR2_X1 U2660 ( .A(n2532), .B(n2862), .ZN(n2534) );
  AOI21_X1 U2661 ( .B1(n3824), .B2(n2890), .A(n2480), .ZN(n2490) );
  AND2_X1 U2662 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2551) );
  NAND2_X1 U2663 ( .A1(n2408), .A2(n2413), .ZN(n2407) );
  INV_X1 U2664 ( .A(n2410), .ZN(n2408) );
  OR2_X1 U2665 ( .A1(n2412), .A2(n2842), .ZN(n2409) );
  OR2_X1 U2666 ( .A1(n2597), .A2(n3337), .ZN(n2616) );
  OAI21_X1 U2667 ( .B1(n3093), .B2(n2875), .A(n2485), .ZN(n3081) );
  NAND2_X1 U2668 ( .A1(n3082), .A2(n3081), .ZN(n3080) );
  NAND2_X1 U2669 ( .A1(n2785), .A2(REG3_REG_20__SCAN_IN), .ZN(n2801) );
  AND2_X1 U2670 ( .A1(n2774), .A2(REG3_REG_19__SCAN_IN), .ZN(n2785) );
  NAND2_X1 U2671 ( .A1(n2226), .A2(n2225), .ZN(n4925) );
  AOI21_X1 U2672 ( .B1(n2228), .B2(n2231), .A(n2195), .ZN(n2225) );
  NAND2_X1 U2673 ( .A1(n2734), .A2(n2228), .ZN(n2226) );
  NAND2_X1 U2674 ( .A1(n2551), .A2(REG3_REG_5__SCAN_IN), .ZN(n2568) );
  OR2_X1 U2675 ( .A1(n3033), .A2(IR_REG_28__SCAN_IN), .ZN(n2479) );
  NAND2_X1 U2676 ( .A1(n3033), .A2(IR_REG_27__SCAN_IN), .ZN(n2478) );
  NOR2_X1 U2677 ( .A1(n2947), .A2(n3064), .ZN(n2928) );
  NAND2_X1 U2678 ( .A1(n2227), .A2(n2230), .ZN(n3637) );
  INV_X1 U2679 ( .A(n2734), .ZN(n2227) );
  NAND2_X1 U2680 ( .A1(n2734), .A2(n2735), .ZN(n3638) );
  AND2_X1 U2681 ( .A1(n2871), .A2(n2870), .ZN(n3523) );
  AND4_X1 U2682 ( .A1(n2705), .A2(n2704), .A3(n2703), .A4(n2702), .ZN(n3473)
         );
  XNOR2_X1 U2683 ( .A(n3266), .B(n3283), .ZN(n3174) );
  NAND2_X1 U2684 ( .A1(n3174), .A2(REG1_REG_4__SCAN_IN), .ZN(n3265) );
  INV_X1 U2685 ( .A(REG3_REG_8__SCAN_IN), .ZN(n3337) );
  NAND2_X1 U2686 ( .A1(n4360), .A2(n3289), .ZN(n3291) );
  NAND2_X1 U2687 ( .A1(n3293), .A2(n4377), .ZN(n3294) );
  NAND2_X1 U2688 ( .A1(n4385), .A2(n3273), .ZN(n4396) );
  XNOR2_X1 U2689 ( .A(n3298), .B(n4517), .ZN(n4408) );
  NAND2_X1 U2690 ( .A1(n4408), .A2(REG2_REG_12__SCAN_IN), .ZN(n4406) );
  NAND2_X1 U2691 ( .A1(n4412), .A2(n3275), .ZN(n3859) );
  XNOR2_X1 U2692 ( .A(n3873), .B(n2208), .ZN(n4418) );
  NAND2_X1 U2693 ( .A1(n2296), .A2(n2295), .ZN(n3873) );
  OR2_X1 U2694 ( .A1(n4322), .A2(REG2_REG_13__SCAN_IN), .ZN(n2295) );
  NAND2_X1 U2695 ( .A1(n4406), .A2(n2293), .ZN(n2296) );
  NOR2_X1 U2696 ( .A1(n2294), .A2(n3871), .ZN(n2293) );
  AND2_X1 U2697 ( .A1(n2691), .A2(n2437), .ZN(n2751) );
  NAND2_X1 U2698 ( .A1(n4436), .A2(n3880), .ZN(n3881) );
  INV_X1 U2699 ( .A(n4176), .ZN(n2314) );
  NOR2_X1 U2700 ( .A1(n2317), .A2(n3521), .ZN(n2310) );
  NAND2_X1 U2701 ( .A1(n3753), .A2(n2318), .ZN(n2317) );
  NOR2_X1 U2702 ( .A1(n3043), .A2(n4176), .ZN(n2318) );
  AND2_X1 U2703 ( .A1(n2316), .A2(n4176), .ZN(n2315) );
  NOR2_X1 U2704 ( .A1(n2314), .A2(n3517), .ZN(n2313) );
  NAND2_X1 U2705 ( .A1(n3753), .A2(n3044), .ZN(n2316) );
  AND2_X1 U2706 ( .A1(n3716), .A2(DATAI_27_), .ZN(n3920) );
  AND2_X1 U2707 ( .A1(n2850), .A2(n2849), .ZN(n3935) );
  NAND2_X1 U2708 ( .A1(n2287), .A2(n2286), .ZN(n4119) );
  AND4_X1 U2709 ( .A1(n2730), .A2(n2729), .A3(n2728), .A4(n2727), .ZN(n4927)
         );
  OAI21_X1 U2710 ( .B1(n3425), .B2(n3017), .A(n3689), .ZN(n4152) );
  AND2_X1 U2711 ( .A1(n3691), .A2(n3670), .ZN(n4158) );
  OAI21_X1 U2712 ( .B1(n2354), .B2(n2347), .A(n2345), .ZN(n2978) );
  AOI21_X1 U2713 ( .B1(n2346), .B2(n2349), .A(n2179), .ZN(n2345) );
  OR2_X1 U2714 ( .A1(n2664), .A2(n2663), .ZN(n2684) );
  INV_X1 U2715 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3276) );
  AND4_X1 U2716 ( .A1(n2690), .A2(n2689), .A3(n2688), .A4(n2687), .ZN(n4155)
         );
  NAND2_X1 U2717 ( .A1(n3015), .A2(n3681), .ZN(n4460) );
  AND2_X1 U2718 ( .A1(n2191), .A2(n3361), .ZN(n2323) );
  NOR2_X1 U2719 ( .A1(n2616), .A2(n2615), .ZN(n2631) );
  AND2_X1 U2720 ( .A1(n2631), .A2(REG3_REG_10__SCAN_IN), .ZN(n2651) );
  NAND2_X1 U2721 ( .A1(n2264), .A2(n3678), .ZN(n3360) );
  NAND2_X1 U2722 ( .A1(n3344), .A2(n3667), .ZN(n2264) );
  INV_X1 U2723 ( .A(n2268), .ZN(n2267) );
  NAND2_X1 U2724 ( .A1(n2269), .A2(n2270), .ZN(n3247) );
  INV_X1 U2725 ( .A(n2265), .ZN(n2270) );
  NAND2_X1 U2726 ( .A1(n3184), .A2(n2272), .ZN(n2269) );
  NAND2_X1 U2727 ( .A1(n2274), .A2(n3661), .ZN(n3199) );
  NAND2_X1 U2728 ( .A1(n2275), .A2(n3658), .ZN(n2274) );
  INV_X1 U2729 ( .A(n3184), .ZN(n2275) );
  OR2_X1 U2730 ( .A1(n3155), .A2(n4488), .ZN(n2342) );
  NAND2_X1 U2731 ( .A1(n3099), .A2(n2340), .ZN(n2339) );
  INV_X1 U2732 ( .A(n4500), .ZN(n4481) );
  INV_X1 U2733 ( .A(n3007), .ZN(n4488) );
  NOR2_X1 U2734 ( .A1(n3138), .A2(n3117), .ZN(n4489) );
  NAND2_X1 U2735 ( .A1(n2304), .A2(n2302), .ZN(n4487) );
  INV_X1 U2736 ( .A(n2303), .ZN(n2302) );
  NAND2_X1 U2737 ( .A1(n2334), .A2(n3123), .ZN(n3125) );
  INV_X1 U2738 ( .A(n2334), .ZN(n3765) );
  INV_X1 U2739 ( .A(n4159), .ZN(n4498) );
  XNOR2_X1 U2740 ( .A(n2252), .B(n3767), .ZN(n2251) );
  AOI21_X1 U2741 ( .B1(n3520), .B2(n3740), .A(n3030), .ZN(n2252) );
  AND2_X1 U2742 ( .A1(n3762), .A2(n2374), .ZN(n2370) );
  NAND2_X1 U2743 ( .A1(n2375), .A2(n3767), .ZN(n2371) );
  OAI22_X1 U2744 ( .A1(n3762), .A2(n2371), .B1(n2375), .B2(n3767), .ZN(n2369)
         );
  NAND2_X1 U2745 ( .A1(n4494), .A2(n4319), .ZN(n4477) );
  NAND2_X1 U2746 ( .A1(n4028), .A2(n2319), .ZN(n3961) );
  NAND2_X1 U2747 ( .A1(n4028), .A2(n2320), .ZN(n3979) );
  NAND2_X1 U2748 ( .A1(n3716), .A2(DATAI_24_), .ZN(n3980) );
  AND2_X1 U2749 ( .A1(n4028), .A2(n4006), .ZN(n4008) );
  AND2_X1 U2750 ( .A1(n4045), .A2(n4026), .ZN(n4028) );
  AND2_X1 U2751 ( .A1(n4124), .A2(n2321), .ZN(n4045) );
  AND2_X1 U2752 ( .A1(n2177), .A2(n4047), .ZN(n2321) );
  NAND2_X1 U2753 ( .A1(n4124), .A2(n4112), .ZN(n4111) );
  NOR2_X1 U2754 ( .A1(n3479), .A2(n2308), .ZN(n4163) );
  INV_X1 U2755 ( .A(n3446), .ZN(n3430) );
  OR2_X1 U2756 ( .A1(n4572), .A2(n3041), .ZN(n4468) );
  OR2_X1 U2757 ( .A1(n4468), .A2(n3430), .ZN(n3479) );
  AND2_X1 U2758 ( .A1(n4553), .A2(n2323), .ZN(n3383) );
  NAND2_X1 U2759 ( .A1(n4553), .A2(n2191), .ZN(n3365) );
  AND3_X1 U2760 ( .A1(n2304), .A2(n2301), .A3(n3200), .ZN(n3256) );
  NAND2_X1 U2761 ( .A1(n2301), .A2(n2304), .ZN(n3197) );
  INV_X1 U2762 ( .A(n4577), .ZN(n4570) );
  NAND2_X1 U2763 ( .A1(n3097), .A2(n4496), .ZN(n3138) );
  AND3_X1 U2764 ( .A1(n3040), .A2(n3109), .A3(n3039), .ZN(n3049) );
  AND2_X1 U2765 ( .A1(n3052), .A2(n2914), .ZN(n3055) );
  INV_X1 U2766 ( .A(IR_REG_29__SCAN_IN), .ZN(n2253) );
  NAND2_X1 U2767 ( .A1(n2466), .A2(IR_REG_31__SCAN_IN), .ZN(n3033) );
  NAND2_X1 U2768 ( .A1(n2913), .A2(n2912), .ZN(n2911) );
  XNOR2_X1 U2769 ( .A(n2476), .B(n2475), .ZN(n2927) );
  INV_X1 U2770 ( .A(IR_REG_20__SCAN_IN), .ZN(n2475) );
  AND2_X1 U2771 ( .A1(n2560), .A2(n2559), .ZN(n3281) );
  OAI211_X1 U2772 ( .C1(IR_REG_1__SCAN_IN), .C2(IR_REG_31__SCAN_IN), .A(n2299), 
        .B(n2498), .ZN(n3072) );
  NAND2_X1 U2773 ( .A1(IR_REG_31__SCAN_IN), .A2(n2181), .ZN(n2299) );
  INV_X1 U2774 ( .A(n3920), .ZN(n3926) );
  NAND2_X1 U2775 ( .A1(n2216), .A2(n2220), .ZN(n3533) );
  INV_X1 U2776 ( .A(n4164), .ZN(n3498) );
  NAND2_X1 U2777 ( .A1(n2701), .A2(n3451), .ZN(n3495) );
  INV_X1 U2778 ( .A(n4926), .ZN(n3641) );
  NAND2_X1 U2779 ( .A1(n3716), .A2(DATAI_23_), .ZN(n4006) );
  AND4_X1 U2780 ( .A1(n2657), .A2(n2656), .A3(n2655), .A4(n2654), .ZN(n3411)
         );
  INV_X1 U2781 ( .A(n2923), .ZN(n2917) );
  NAND2_X1 U2782 ( .A1(n3307), .A2(n3306), .ZN(n2243) );
  NAND2_X1 U2783 ( .A1(n3229), .A2(n2549), .ZN(n3210) );
  NAND2_X1 U2784 ( .A1(n3210), .A2(n3209), .ZN(n3208) );
  NAND2_X1 U2785 ( .A1(n2538), .A2(n2537), .ZN(n3231) );
  INV_X1 U2786 ( .A(n3135), .ZN(n4496) );
  OAI22_X1 U2787 ( .A1(n3558), .A2(n2814), .B1(n2813), .B2(n2812), .ZN(n3607)
         );
  NOR2_X1 U2788 ( .A1(n3607), .A2(n3608), .ZN(n3606) );
  NAND2_X1 U2789 ( .A1(n3406), .A2(n2650), .ZN(n3437) );
  NAND2_X1 U2790 ( .A1(n3090), .A2(n2505), .ZN(n3153) );
  INV_X1 U2791 ( .A(n3248), .ZN(n3255) );
  AOI21_X1 U2792 ( .B1(n2928), .B2(n4182), .A(n4503), .ZN(n3624) );
  NAND2_X1 U2793 ( .A1(n3208), .A2(n2567), .ZN(n3240) );
  AND2_X1 U2794 ( .A1(n2878), .A2(n2855), .ZN(n3944) );
  INV_X1 U2795 ( .A(n3620), .ZN(n4931) );
  INV_X1 U2796 ( .A(n3019), .ZN(n3644) );
  AND2_X1 U2797 ( .A1(n2890), .A2(n2935), .ZN(n3803) );
  INV_X1 U2798 ( .A(n3523), .ZN(n3937) );
  INV_X1 U2799 ( .A(n3790), .ZN(n3956) );
  INV_X1 U2800 ( .A(n3935), .ZN(n3976) );
  OAI211_X1 U2801 ( .C1(n3982), .C2(n2884), .A(n2838), .B(n2837), .ZN(n3810)
         );
  OAI211_X1 U2802 ( .C1(n4009), .C2(n2884), .A(n2828), .B(n2827), .ZN(n4018)
         );
  NAND4_X1 U2803 ( .A1(n2806), .A2(n2805), .A3(n2804), .A4(n2803), .ZN(n4063)
         );
  NAND4_X1 U2804 ( .A1(n2790), .A2(n2789), .A3(n2788), .A4(n2787), .ZN(n4041)
         );
  INV_X1 U2805 ( .A(n4104), .ZN(n4137) );
  INV_X1 U2806 ( .A(n3473), .ZN(n3812) );
  INV_X1 U2807 ( .A(n4155), .ZN(n3813) );
  INV_X1 U2808 ( .A(n3016), .ZN(n4463) );
  INV_X1 U2809 ( .A(n3411), .ZN(n3814) );
  INV_X1 U2810 ( .A(n2959), .ZN(n3822) );
  NAND2_X1 U2811 ( .A1(n2506), .A2(REG0_REG_1__SCAN_IN), .ZN(n2494) );
  NAND2_X1 U2812 ( .A1(n3837), .A2(n3838), .ZN(n3849) );
  XNOR2_X1 U2813 ( .A(n3284), .B(n4323), .ZN(n3282) );
  NAND2_X1 U2814 ( .A1(n2292), .A2(n2290), .ZN(n4339) );
  NAND2_X1 U2815 ( .A1(n2291), .A2(n4323), .ZN(n2290) );
  NAND2_X1 U2816 ( .A1(n3282), .A2(REG2_REG_4__SCAN_IN), .ZN(n2292) );
  INV_X1 U2817 ( .A(n3284), .ZN(n2291) );
  NAND2_X1 U2818 ( .A1(n4339), .A2(n4340), .ZN(n4338) );
  AND2_X1 U2819 ( .A1(n3265), .A2(n2333), .ZN(n4335) );
  NAND2_X1 U2820 ( .A1(n3266), .A2(n4323), .ZN(n2333) );
  AND2_X1 U2821 ( .A1(n2329), .A2(n4525), .ZN(n3267) );
  XNOR2_X1 U2822 ( .A(n3291), .B(n4522), .ZN(n4368) );
  XNOR2_X1 U2823 ( .A(n3274), .B(n4517), .ZN(n4413) );
  NAND2_X1 U2824 ( .A1(n4406), .A2(n3299), .ZN(n3872) );
  OR2_X1 U2825 ( .A1(n2695), .A2(n2694), .ZN(n3870) );
  XNOR2_X1 U2826 ( .A(n3862), .B(n2208), .ZN(n4422) );
  XNOR2_X1 U2827 ( .A(n3879), .B(n3878), .ZN(n4437) );
  NAND2_X1 U2828 ( .A1(n4437), .A2(n4435), .ZN(n4436) );
  NOR2_X1 U2829 ( .A1(n4441), .A2(n3865), .ZN(n3869) );
  AND2_X1 U2830 ( .A1(n3070), .A2(n3069), .ZN(n4451) );
  INV_X1 U2831 ( .A(n3892), .ZN(n2325) );
  NOR2_X1 U2832 ( .A1(n2315), .A2(n2313), .ZN(n2312) );
  NAND2_X1 U2833 ( .A1(n3924), .A2(n2310), .ZN(n2309) );
  OR2_X1 U2834 ( .A1(n3924), .A2(n2314), .ZN(n2311) );
  NOR2_X1 U2835 ( .A1(n3516), .A2(n2316), .ZN(n4181) );
  OR2_X1 U2836 ( .A1(n2879), .A2(n3904), .ZN(n3519) );
  NAND2_X1 U2837 ( .A1(n2376), .A2(n2382), .ZN(n3968) );
  NAND2_X1 U2838 ( .A1(n4024), .A2(n2383), .ZN(n2376) );
  NOR2_X1 U2839 ( .A1(n4212), .A2(n2385), .ZN(n3987) );
  NAND2_X1 U2840 ( .A1(n4108), .A2(n2992), .ZN(n4079) );
  NAND2_X1 U2841 ( .A1(n2344), .A2(n2346), .ZN(n3429) );
  NAND2_X1 U2842 ( .A1(n2354), .A2(n2348), .ZN(n2344) );
  INV_X1 U2843 ( .A(n2975), .ZN(n2350) );
  NAND2_X1 U2844 ( .A1(n2354), .A2(n2172), .ZN(n2353) );
  AOI21_X1 U2845 ( .B1(n4159), .B2(n3196), .A(n4507), .ZN(n4131) );
  NAND2_X1 U2846 ( .A1(n3055), .A2(n3038), .ZN(n4166) );
  NAND2_X1 U2847 ( .A1(n3098), .A2(n2960), .ZN(n4474) );
  INV_X1 U2848 ( .A(n4166), .ZN(n4503) );
  AND2_X1 U2849 ( .A1(n4147), .A2(n3116), .ZN(n4504) );
  OR2_X1 U2850 ( .A1(n4228), .A2(n4227), .ZN(n4294) );
  AND2_X1 U2851 ( .A1(n4576), .A2(n4575), .ZN(n4600) );
  NAND2_X1 U2852 ( .A1(n3055), .A2(n3054), .ZN(n4508) );
  INV_X1 U2853 ( .A(n2452), .ZN(n3061) );
  AND2_X1 U2854 ( .A1(n2467), .A2(n2466), .ZN(n3058) );
  CLKBUF_X1 U2855 ( .A(n2462), .Z(n2464) );
  NOR2_X1 U2856 ( .A1(n2463), .A2(n2444), .ZN(n4315) );
  NAND2_X1 U2857 ( .A1(n2768), .A2(n2442), .ZN(n2460) );
  OR2_X1 U2858 ( .A1(n2458), .A2(n2459), .ZN(n2461) );
  XNOR2_X1 U2859 ( .A(n2469), .B(IR_REG_24__SCAN_IN), .ZN(n4316) );
  NAND2_X1 U2860 ( .A1(n2911), .A2(IR_REG_31__SCAN_IN), .ZN(n2469) );
  NAND2_X1 U2861 ( .A1(n3066), .A2(STATE_REG_SCAN_IN), .ZN(n4510) );
  XNOR2_X1 U2862 ( .A(n2483), .B(IR_REG_22__SCAN_IN), .ZN(n4317) );
  NOR2_X1 U2863 ( .A1(n2473), .A2(n2211), .ZN(n4318) );
  INV_X1 U2864 ( .A(n2482), .ZN(n2211) );
  INV_X1 U2865 ( .A(n2472), .ZN(n2473) );
  INV_X1 U2866 ( .A(n3898), .ZN(n4320) );
  AND2_X1 U2867 ( .A1(n2544), .A2(n2529), .ZN(n4324) );
  NAND2_X1 U2868 ( .A1(n2498), .A2(IR_REG_31__SCAN_IN), .ZN(n2513) );
  AOI211_X1 U2869 ( .C1(ADDR_REG_18__SCAN_IN), .C2(n4451), .A(n4450), .B(n4449), .ZN(n4457) );
  XNOR2_X1 U2870 ( .A(n2326), .B(n2325), .ZN(n3902) );
  OR2_X1 U2871 ( .A1(n3906), .A2(n4247), .ZN(n3046) );
  OAI21_X1 U2872 ( .B1(n3903), .B2(n2367), .A(n2363), .ZN(n3047) );
  OR2_X1 U2873 ( .A1(n3908), .A2(n4601), .ZN(n2367) );
  NAND2_X1 U2874 ( .A1(n2255), .A2(n2254), .ZN(U3515) );
  AND2_X1 U2875 ( .A1(n3051), .A2(n2203), .ZN(n2254) );
  INV_X1 U2876 ( .A(n2256), .ZN(n2255) );
  NOR2_X1 U2877 ( .A1(n2470), .A2(n2184), .ZN(n2458) );
  NAND2_X1 U2878 ( .A1(n2249), .A2(n2430), .ZN(n2557) );
  NOR2_X1 U2879 ( .A1(n3370), .A2(n2974), .ZN(n2172) );
  INV_X1 U2880 ( .A(n2349), .ZN(n2348) );
  NAND2_X1 U2881 ( .A1(n2172), .A2(n2355), .ZN(n2349) );
  NAND2_X1 U2882 ( .A1(n2445), .A2(n2391), .ZN(n2174) );
  NAND2_X1 U2883 ( .A1(n3407), .A2(n3404), .ZN(n2175) );
  AND3_X1 U2884 ( .A1(n2277), .A2(n2189), .A3(n2276), .ZN(n2176) );
  AND2_X1 U2885 ( .A1(n2322), .A2(n4066), .ZN(n2177) );
  INV_X1 U2886 ( .A(n3278), .ZN(n4518) );
  AND2_X1 U2887 ( .A1(n2661), .A2(n2671), .ZN(n3278) );
  AND2_X1 U2888 ( .A1(n3052), .A2(n3115), .ZN(n2533) );
  AND2_X1 U2889 ( .A1(n3061), .A2(n2453), .ZN(n2521) );
  INV_X1 U2890 ( .A(n2462), .ZN(n2444) );
  NAND4_X1 U2891 ( .A1(n2496), .A2(n2495), .A3(n2494), .A4(n2493), .ZN(n2956)
         );
  AND4_X1 U2892 ( .A1(n2512), .A2(n2511), .A3(n2510), .A4(n2509), .ZN(n2959)
         );
  OR2_X1 U2893 ( .A1(n4018), .A2(n4002), .ZN(n2178) );
  NAND2_X1 U2894 ( .A1(n2250), .A2(n3036), .ZN(n3908) );
  INV_X1 U2895 ( .A(n3675), .ZN(n2271) );
  INV_X1 U2896 ( .A(n2976), .ZN(n2355) );
  AND2_X1 U2897 ( .A1(n3016), .A2(n3446), .ZN(n2179) );
  AND2_X1 U2898 ( .A1(n3621), .A2(n4085), .ZN(n2180) );
  AND2_X1 U2899 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2181)
         );
  OR2_X1 U2900 ( .A1(n3606), .A2(n2414), .ZN(n2182) );
  INV_X1 U2901 ( .A(n2347), .ZN(n2346) );
  NOR2_X1 U2902 ( .A1(n2351), .A2(n2976), .ZN(n2347) );
  AND2_X1 U2903 ( .A1(n2238), .A2(n2418), .ZN(n2183) );
  OR2_X1 U2904 ( .A1(n2441), .A2(n2173), .ZN(n2184) );
  INV_X1 U2905 ( .A(IR_REG_26__SCAN_IN), .ZN(n2443) );
  NOR2_X1 U2906 ( .A1(n3974), .A2(n4006), .ZN(n2185) );
  NAND2_X1 U2907 ( .A1(n2497), .A2(n2433), .ZN(n2526) );
  NAND2_X1 U2908 ( .A1(n3815), .A2(n3413), .ZN(n2186) );
  AND2_X1 U2909 ( .A1(n2386), .A2(n2253), .ZN(n2187) );
  AND2_X1 U2910 ( .A1(n2405), .A2(n2404), .ZN(n2188) );
  NAND2_X1 U2911 ( .A1(n3735), .A2(n2282), .ZN(n2189) );
  INV_X1 U2912 ( .A(n2735), .ZN(n2230) );
  XOR2_X1 U2913 ( .A(n2707), .B(n2888), .Z(n2190) );
  INV_X1 U2914 ( .A(n2237), .ZN(n2691) );
  INV_X1 U2915 ( .A(n3767), .ZN(n2374) );
  AND2_X1 U2916 ( .A1(n3314), .A2(n3352), .ZN(n2191) );
  AND2_X1 U2917 ( .A1(n2353), .A2(n2350), .ZN(n2192) );
  OR2_X1 U2918 ( .A1(n2865), .A2(n2864), .ZN(n2193) );
  NOR2_X1 U2919 ( .A1(n3436), .A2(n2431), .ZN(n2194) );
  AND2_X1 U2920 ( .A1(n2738), .A2(n2737), .ZN(n2195) );
  AND2_X1 U2921 ( .A1(n3451), .A2(n2190), .ZN(n2196) );
  AND2_X1 U2922 ( .A1(n2323), .A2(n3382), .ZN(n2197) );
  INV_X1 U2923 ( .A(n3564), .ZN(n2222) );
  INV_X1 U2924 ( .A(IR_REG_25__SCAN_IN), .ZN(n2442) );
  INV_X1 U2925 ( .A(n2224), .ZN(n2223) );
  NAND2_X1 U2926 ( .A1(n2193), .A2(n3565), .ZN(n2224) );
  NAND2_X1 U2927 ( .A1(n2289), .A2(n4136), .ZN(n2198) );
  INV_X1 U2928 ( .A(n2842), .ZN(n2413) );
  INV_X1 U2929 ( .A(IR_REG_27__SCAN_IN), .ZN(n2391) );
  OR2_X1 U2930 ( .A1(n3479), .A2(n3478), .ZN(n2199) );
  NOR2_X1 U2931 ( .A1(n3194), .A2(n2273), .ZN(n2272) );
  NAND2_X1 U2932 ( .A1(n2243), .A2(n2596), .ZN(n3333) );
  INV_X1 U2933 ( .A(n3334), .ZN(n2419) );
  INV_X1 U2934 ( .A(n3782), .ZN(n2336) );
  INV_X1 U2935 ( .A(n3472), .ZN(n3478) );
  NOR3_X1 U2936 ( .A1(n3479), .A2(n2306), .A3(n4142), .ZN(n2305) );
  NAND2_X1 U2937 ( .A1(n2343), .A2(n3005), .ZN(n3098) );
  INV_X1 U2938 ( .A(n4101), .ZN(n4112) );
  OR2_X1 U2939 ( .A1(n3479), .A2(n2306), .ZN(n2200) );
  AND2_X1 U2940 ( .A1(n3716), .A2(DATAI_20_), .ZN(n4071) );
  INV_X1 U2941 ( .A(n3874), .ZN(n2208) );
  AND2_X2 U2942 ( .A1(n3113), .A2(n4166), .ZN(n4507) );
  INV_X1 U2943 ( .A(n4561), .ZN(n2366) );
  AND2_X1 U2944 ( .A1(n4553), .A2(n3314), .ZN(n2201) );
  AND2_X2 U2945 ( .A1(n3049), .A2(n3048), .ZN(n4585) );
  AND2_X2 U2946 ( .A1(n3049), .A2(n3111), .ZN(n4604) );
  AND2_X1 U2947 ( .A1(n3032), .A2(n3031), .ZN(n4483) );
  INV_X1 U2948 ( .A(n3633), .ZN(n3942) );
  NOR2_X1 U2949 ( .A1(n2466), .A2(IR_REG_27__SCAN_IN), .ZN(n2929) );
  NAND2_X1 U2950 ( .A1(n3091), .A2(n3092), .ZN(n3090) );
  OR2_X1 U2951 ( .A1(n3870), .A2(n3860), .ZN(n2202) );
  OR2_X1 U2952 ( .A1(n4585), .A2(n3050), .ZN(n2203) );
  AND2_X1 U2953 ( .A1(n3877), .A2(REG2_REG_15__SCAN_IN), .ZN(n2204) );
  AND2_X1 U2954 ( .A1(n3716), .A2(DATAI_25_), .ZN(n3959) );
  AND2_X1 U2955 ( .A1(n2319), .A2(n3942), .ZN(n2205) );
  AND2_X1 U2956 ( .A1(n3894), .A2(REG2_REG_18__SCAN_IN), .ZN(n2206) );
  OR2_X1 U2957 ( .A1(n4513), .A2(n3891), .ZN(n2207) );
  INV_X1 U2958 ( .A(IR_REG_30__SCAN_IN), .ZN(n2446) );
  INV_X1 U2959 ( .A(U4043), .ZN(n3823) );
  NAND2_X1 U2960 ( .A1(n3893), .A2(n2298), .ZN(n4447) );
  NOR2_X1 U2961 ( .A1(n4425), .A2(n2204), .ZN(n3879) );
  AOI21_X1 U2962 ( .B1(n4325), .B2(REG2_REG_2__SCAN_IN), .A(n3846), .ZN(n3168)
         );
  NAND2_X1 U2963 ( .A1(n2538), .A2(n2214), .ZN(n3229) );
  NAND2_X1 U2964 ( .A1(n3567), .A2(n2223), .ZN(n2216) );
  AOI21_X1 U2965 ( .B1(n3567), .B2(n3565), .A(n3564), .ZN(n3630) );
  OAI21_X1 U2966 ( .B1(n3567), .B2(n2219), .A(n2217), .ZN(n2923) );
  NAND4_X1 U2967 ( .A1(n2233), .A2(n2437), .A3(n2234), .A4(n2248), .ZN(n2470)
         );
  NOR2_X2 U2968 ( .A1(n2237), .A2(n2235), .ZN(n2440) );
  INV_X1 U2969 ( .A(n2440), .ZN(n2474) );
  NAND2_X1 U2970 ( .A1(n2444), .A2(n2386), .ZN(n2932) );
  NAND2_X1 U2971 ( .A1(n2444), .A2(n2187), .ZN(n2449) );
  OAI21_X1 U2972 ( .B1(n3184), .B2(n2265), .A(n2267), .ZN(n3010) );
  OAI21_X1 U2973 ( .B1(n2271), .B2(n2272), .A(n3677), .ZN(n2268) );
  INV_X1 U2974 ( .A(n3661), .ZN(n2273) );
  NAND2_X1 U2975 ( .A1(n3505), .A2(n2281), .ZN(n2287) );
  MUX2_X1 U2976 ( .A(n3063), .B(REG2_REG_1__SCAN_IN), .S(n3072), .Z(n3837) );
  NAND2_X1 U2977 ( .A1(n2300), .A2(n2440), .ZN(n2466) );
  NAND2_X1 U2978 ( .A1(n2440), .A2(n2426), .ZN(n2462) );
  INV_X1 U2979 ( .A(n2305), .ZN(n4240) );
  NAND3_X1 U2980 ( .A1(n2311), .A2(n2312), .A3(n2309), .ZN(n4328) );
  NOR2_X1 U2981 ( .A1(n3875), .A2(n4417), .ZN(n4427) );
  XNOR2_X2 U2982 ( .A(n2513), .B(IR_REG_2__SCAN_IN), .ZN(n4325) );
  MUX2_X1 U2983 ( .A(n4326), .B(DATAI_1_), .S(n3716), .Z(n3136) );
  NAND2_X1 U2984 ( .A1(n3765), .A2(n2335), .ZN(n3124) );
  INV_X1 U2985 ( .A(n3123), .ZN(n2335) );
  NAND2_X1 U2986 ( .A1(n3765), .A2(n2336), .ZN(n3127) );
  NAND2_X1 U2987 ( .A1(n2334), .A2(n3782), .ZN(n3126) );
  INV_X1 U2988 ( .A(n2960), .ZN(n2341) );
  NAND3_X1 U2989 ( .A1(n2339), .A2(n2342), .A3(n2337), .ZN(n3182) );
  NAND4_X1 U2990 ( .A1(n2338), .A2(n2960), .A3(n3655), .A4(n3652), .ZN(n2337)
         );
  INV_X1 U2991 ( .A(n2961), .ZN(n2338) );
  NOR2_X1 U2992 ( .A1(n2961), .A2(n2341), .ZN(n2340) );
  INV_X1 U2993 ( .A(n3371), .ZN(n2354) );
  NAND2_X1 U2994 ( .A1(n2991), .A2(n2358), .ZN(n2357) );
  NAND2_X1 U2995 ( .A1(n3515), .A2(n2370), .ZN(n2361) );
  OR2_X1 U2996 ( .A1(n4604), .A2(REG1_REG_29__SCAN_IN), .ZN(n2372) );
  INV_X1 U2997 ( .A(n3908), .ZN(n2373) );
  OAI21_X1 U2998 ( .B1(n4024), .B2(n2380), .A(n2377), .ZN(n3949) );
  OAI21_X2 U2999 ( .B1(n3195), .B2(n2964), .A(n2965), .ZN(n3326) );
  NAND2_X1 U3000 ( .A1(n2963), .A2(n2962), .ZN(n3195) );
  OAI21_X2 U3001 ( .B1(n3502), .B2(n2984), .A(n2986), .ZN(n4134) );
  NAND2_X2 U3002 ( .A1(n2983), .A2(n2982), .ZN(n3502) );
  NAND3_X1 U3003 ( .A1(n2388), .A2(n3143), .A3(n2387), .ZN(n2538) );
  NAND2_X1 U3004 ( .A1(n3154), .A2(n2519), .ZN(n2387) );
  NAND2_X1 U3005 ( .A1(n3153), .A2(n2519), .ZN(n2388) );
  NAND2_X1 U3006 ( .A1(n3151), .A2(n2519), .ZN(n3144) );
  NAND2_X1 U3007 ( .A1(n2390), .A2(n2389), .ZN(n3151) );
  INV_X1 U3008 ( .A(n3209), .ZN(n2395) );
  NAND2_X1 U3009 ( .A1(n3210), .A2(n2394), .ZN(n2397) );
  NAND2_X1 U3010 ( .A1(n3237), .A2(n3238), .ZN(n2399) );
  INV_X1 U3011 ( .A(n3607), .ZN(n2400) );
  OAI21_X1 U3012 ( .B1(n2400), .B2(n2188), .A(n2401), .ZN(n3567) );
  OAI21_X1 U3013 ( .B1(n3333), .B2(n3335), .A(n3334), .ZN(n3388) );
  NAND2_X1 U3014 ( .A1(n3335), .A2(n3334), .ZN(n2422) );
  OAI21_X1 U3015 ( .B1(n3451), .B2(n2190), .A(n3493), .ZN(n2425) );
  NOR2_X1 U3016 ( .A1(n2470), .A2(n2441), .ZN(n2468) );
  MUX2_X2 U3017 ( .A(REG0_REG_28__SCAN_IN), .B(n4263), .S(n4585), .Z(n4264) );
  MUX2_X2 U3018 ( .A(REG1_REG_28__SCAN_IN), .B(n4263), .S(n4604), .Z(n4190) );
  NAND2_X1 U3019 ( .A1(n2957), .A2(n3097), .ZN(n3650) );
  NAND2_X1 U3020 ( .A1(n4501), .A2(n3136), .ZN(n3651) );
  AND2_X1 U3021 ( .A1(n4312), .A2(n3061), .ZN(n2507) );
  CLKBUF_X1 U3022 ( .A(n2956), .Z(n2957) );
  OAI22_X2 U3023 ( .A1(n3949), .A2(n2999), .B1(n3935), .B2(n3954), .ZN(n3932)
         );
  NOR2_X1 U3024 ( .A1(n2431), .A2(n2682), .ZN(n2428) );
  NAND2_X1 U3025 ( .A1(n3441), .A2(n3440), .ZN(n2429) );
  AND2_X1 U3026 ( .A1(n2527), .A2(n2434), .ZN(n2430) );
  AND2_X1 U3027 ( .A1(n2677), .A2(n2676), .ZN(n2431) );
  AND2_X1 U3028 ( .A1(n2922), .A2(n2921), .ZN(n2432) );
  AND2_X1 U3029 ( .A1(n4080), .A2(n4081), .ZN(n4110) );
  INV_X1 U3030 ( .A(n4110), .ZN(n2990) );
  INV_X1 U3031 ( .A(IR_REG_4__SCAN_IN), .ZN(n2434) );
  INV_X1 U3032 ( .A(IR_REG_17__SCAN_IN), .ZN(n2436) );
  NAND2_X1 U3033 ( .A1(n3136), .A2(n2885), .ZN(n2499) );
  INV_X1 U3034 ( .A(n4102), .ZN(n3621) );
  INV_X1 U3035 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2663) );
  OR2_X1 U3036 ( .A1(n2740), .A2(n2739), .ZN(n2761) );
  INV_X1 U3037 ( .A(n3959), .ZN(n3954) );
  NOR2_X1 U3038 ( .A1(n2710), .A2(n2709), .ZN(n2725) );
  INV_X1 U3039 ( .A(n3413), .ZN(n3382) );
  INV_X1 U3040 ( .A(n4047), .ZN(n4039) );
  AND2_X1 U3041 ( .A1(n4313), .A2(n3065), .ZN(n4088) );
  INV_X1 U3042 ( .A(n3005), .ZN(n3764) );
  INV_X1 U3043 ( .A(n4316), .ZN(n2897) );
  AND2_X1 U3044 ( .A1(n2626), .A2(n2625), .ZN(n2639) );
  INV_X1 U3045 ( .A(n3320), .ZN(n3314) );
  INV_X1 U3046 ( .A(n4091), .ZN(n4085) );
  OR2_X1 U3047 ( .A1(n2801), .A2(n2800), .ZN(n2815) );
  INV_X1 U3048 ( .A(n4142), .ZN(n3580) );
  INV_X1 U3049 ( .A(n3815), .ZN(n4461) );
  INV_X1 U3050 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2615) );
  OR2_X1 U3051 ( .A1(n2684), .A2(n3276), .ZN(n2710) );
  INV_X1 U3052 ( .A(n3041), .ZN(n4469) );
  NOR2_X1 U3053 ( .A1(n2761), .A2(n2760), .ZN(n2774) );
  NOR2_X1 U3054 ( .A1(n2568), .A2(n3241), .ZN(n2580) );
  AND2_X1 U3055 ( .A1(n4318), .A2(n4317), .ZN(n3065) );
  OR2_X1 U3056 ( .A1(n3963), .A2(n2884), .ZN(n2850) );
  NOR2_X1 U3057 ( .A1(n2815), .A2(n4835), .ZN(n2825) );
  INV_X1 U3058 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3241) );
  INV_X1 U3059 ( .A(n4477), .ZN(n4182) );
  AOI21_X1 U3060 ( .B1(n3790), .B2(n3942), .A(n3000), .ZN(n3911) );
  INV_X1 U3061 ( .A(n3810), .ZN(n4005) );
  AND4_X1 U3062 ( .A1(n2745), .A2(n2744), .A3(n2743), .A4(n2742), .ZN(n4104)
         );
  INV_X1 U3063 ( .A(n4088), .ZN(n4478) );
  OR2_X1 U3064 ( .A1(n4115), .A2(n4577), .ZN(n4096) );
  AND2_X1 U3065 ( .A1(n2898), .A2(n2897), .ZN(n2899) );
  NAND2_X1 U3066 ( .A1(n3716), .A2(DATAI_22_), .ZN(n4026) );
  AND2_X1 U3067 ( .A1(n3657), .A2(n3654), .ZN(n4476) );
  AND2_X1 U3068 ( .A1(n2825), .A2(REG3_REG_23__SCAN_IN), .ZN(n2835) );
  OR2_X1 U3069 ( .A1(n2844), .A2(n3569), .ZN(n2854) );
  NAND2_X1 U3070 ( .A1(n2835), .A2(REG3_REG_24__SCAN_IN), .ZN(n2844) );
  INV_X1 U3071 ( .A(n3648), .ZN(n4939) );
  AOI21_X1 U3072 ( .B1(n2683), .B2(n2194), .A(n2428), .ZN(n3455) );
  AND2_X1 U3073 ( .A1(n3716), .A2(DATAI_26_), .ZN(n3633) );
  INV_X1 U3074 ( .A(n2856), .ZN(n2884) );
  AND4_X1 U3075 ( .A1(n2767), .A2(n2766), .A3(n2765), .A4(n2764), .ZN(n4120)
         );
  AND2_X1 U3076 ( .A1(n3070), .A2(n3068), .ZN(n3826) );
  AND2_X1 U3077 ( .A1(n3727), .A2(n3696), .ZN(n4136) );
  INV_X1 U3078 ( .A(n4483), .ZN(n4497) );
  INV_X1 U3079 ( .A(n4096), .ZN(n4491) );
  AOI21_X1 U3080 ( .B1(n2910), .B2(n3060), .A(n2899), .ZN(n3111) );
  NAND2_X1 U3081 ( .A1(n3716), .A2(DATAI_21_), .ZN(n4047) );
  INV_X1 U3082 ( .A(n4253), .ZN(n4583) );
  NAND2_X1 U3083 ( .A1(n2896), .A2(n3058), .ZN(n3054) );
  NAND2_X1 U3084 ( .A1(n2461), .A2(n2460), .ZN(n2463) );
  AND2_X1 U3085 ( .A1(n2719), .A2(n2731), .ZN(n3877) );
  AND2_X1 U3086 ( .A1(n2603), .A2(n2591), .ZN(n3280) );
  NAND2_X1 U3087 ( .A1(n2917), .A2(n2916), .ZN(n2955) );
  NAND2_X1 U3088 ( .A1(n2928), .A2(n2915), .ZN(n3648) );
  OAI21_X1 U3089 ( .B1(n3519), .B2(n2884), .A(n2883), .ZN(n3913) );
  OAI211_X1 U3090 ( .C1(n2884), .C2(n4029), .A(n2818), .B(n2817), .ZN(n4040)
         );
  INV_X1 U3091 ( .A(n4407), .ZN(n4445) );
  NAND2_X1 U3092 ( .A1(n3826), .A2(n3163), .ZN(n4458) );
  AND2_X1 U3093 ( .A1(n3381), .A2(n3380), .ZN(n4576) );
  INV_X1 U3094 ( .A(n4131), .ZN(n4150) );
  NAND2_X1 U3095 ( .A1(n4604), .A2(n4570), .ZN(n4247) );
  INV_X1 U3096 ( .A(n4604), .ZN(n4601) );
  OR2_X1 U3097 ( .A1(n3906), .A2(n4308), .ZN(n3051) );
  NAND2_X1 U3098 ( .A1(n4585), .A2(n4570), .ZN(n4308) );
  INV_X1 U3099 ( .A(n4585), .ZN(n4584) );
  INV_X1 U3100 ( .A(n4508), .ZN(n4509) );
  INV_X1 U3101 ( .A(n3297), .ZN(n4517) );
  INV_X1 U3102 ( .A(n3280), .ZN(n4524) );
  INV_X1 U3103 ( .A(n2453), .ZN(n4312) );
  INV_X1 U3104 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2451) );
  OR2_X1 U3105 ( .A1(n2171), .A2(n2451), .ZN(n2457) );
  NAND2_X1 U3106 ( .A1(n2506), .A2(REG0_REG_0__SCAN_IN), .ZN(n2456) );
  NAND2_X1 U3107 ( .A1(n2507), .A2(REG3_REG_0__SCAN_IN), .ZN(n2455) );
  NAND2_X1 U3108 ( .A1(n2521), .A2(REG1_REG_0__SCAN_IN), .ZN(n2454) );
  NAND2_X1 U3109 ( .A1(n2464), .A2(IR_REG_31__SCAN_IN), .ZN(n2465) );
  MUX2_X1 U3110 ( .A(IR_REG_31__SCAN_IN), .B(n2465), .S(IR_REG_26__SCAN_IN), 
        .Z(n2467) );
  OR2_X1 U3111 ( .A1(n2468), .A2(n2768), .ZN(n2913) );
  NAND2_X1 U3112 ( .A1(n2470), .A2(IR_REG_31__SCAN_IN), .ZN(n2471) );
  MUX2_X1 U3113 ( .A(IR_REG_31__SCAN_IN), .B(n2471), .S(IR_REG_21__SCAN_IN), 
        .Z(n2472) );
  NAND2_X1 U3114 ( .A1(n2474), .A2(IR_REG_31__SCAN_IN), .ZN(n2487) );
  NAND2_X1 U3115 ( .A1(n2487), .A2(n2486), .ZN(n2489) );
  NAND2_X1 U3116 ( .A1(n2489), .A2(IR_REG_31__SCAN_IN), .ZN(n2476) );
  INV_X1 U3117 ( .A(n3003), .ZN(n3115) );
  NAND2_X1 U3118 ( .A1(n2391), .A2(IR_REG_28__SCAN_IN), .ZN(n2477) );
  MUX2_X1 U3119 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n3716), .Z(n3135) );
  AND2_X1 U3120 ( .A1(n3135), .A2(n2885), .ZN(n2480) );
  INV_X1 U3121 ( .A(n3052), .ZN(n2484) );
  NAND2_X1 U3122 ( .A1(n2484), .A2(REG1_REG_0__SCAN_IN), .ZN(n2481) );
  NAND2_X1 U3123 ( .A1(n2490), .A2(n2481), .ZN(n3082) );
  INV_X1 U3124 ( .A(n4318), .ZN(n3763) );
  NAND2_X1 U3125 ( .A1(n2482), .A2(IR_REG_31__SCAN_IN), .ZN(n2483) );
  AOI22_X1 U3126 ( .A1(n3135), .A2(n2533), .B1(n2484), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2485) );
  OR2_X1 U3127 ( .A1(n2487), .A2(n2486), .ZN(n2488) );
  NAND2_X1 U3128 ( .A1(n4317), .A2(n3898), .ZN(n2934) );
  NAND2_X1 U3129 ( .A1(n2490), .A2(n2888), .ZN(n2491) );
  NAND2_X1 U3130 ( .A1(n3080), .A2(n2491), .ZN(n3091) );
  NAND2_X1 U3131 ( .A1(n2492), .A2(REG2_REG_1__SCAN_IN), .ZN(n2496) );
  NAND2_X1 U3132 ( .A1(n2507), .A2(REG3_REG_1__SCAN_IN), .ZN(n2495) );
  NAND2_X1 U3133 ( .A1(n2521), .A2(REG1_REG_1__SCAN_IN), .ZN(n2493) );
  NAND2_X1 U3134 ( .A1(n2956), .A2(n2533), .ZN(n2500) );
  INV_X1 U3135 ( .A(n3072), .ZN(n4326) );
  NAND2_X1 U3136 ( .A1(n2500), .A2(n2499), .ZN(n2501) );
  INV_X1 U3137 ( .A(n2956), .ZN(n4501) );
  INV_X1 U3138 ( .A(n2502), .ZN(n2504) );
  NAND2_X1 U3139 ( .A1(n2504), .A2(n2503), .ZN(n2505) );
  NAND2_X1 U3140 ( .A1(n2506), .A2(REG0_REG_2__SCAN_IN), .ZN(n2512) );
  NAND2_X1 U3141 ( .A1(n2507), .A2(REG3_REG_2__SCAN_IN), .ZN(n2511) );
  NAND2_X1 U3142 ( .A1(n2521), .A2(REG1_REG_2__SCAN_IN), .ZN(n2510) );
  INV_X1 U3143 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2508) );
  OR2_X1 U3144 ( .A1(n2539), .A2(n2508), .ZN(n2509) );
  MUX2_X1 U3145 ( .A(n4325), .B(DATAI_2_), .S(n3716), .Z(n3117) );
  INV_X1 U3146 ( .A(n3117), .ZN(n3156) );
  OAI22_X1 U3147 ( .A1(n2959), .A2(n2873), .B1(n2872), .B2(n3156), .ZN(n2514)
         );
  XNOR2_X1 U31480 ( .A(n2514), .B(n2862), .ZN(n2515) );
  OAI22_X1 U31490 ( .A1(n2959), .A2(n2875), .B1(n2873), .B2(n3156), .ZN(n2516)
         );
  XNOR2_X1 U3150 ( .A(n2515), .B(n2516), .ZN(n3154) );
  INV_X1 U3151 ( .A(n2515), .ZN(n2518) );
  INV_X1 U3152 ( .A(n2516), .ZN(n2517) );
  NAND2_X1 U3153 ( .A1(n2518), .A2(n2517), .ZN(n2519) );
  INV_X1 U3154 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2520) );
  OR2_X1 U3155 ( .A1(n2171), .A2(n2520), .ZN(n2525) );
  INV_X1 U3156 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4486) );
  NAND2_X1 U3157 ( .A1(n2507), .A2(n4486), .ZN(n2524) );
  NAND2_X1 U3158 ( .A1(n2506), .A2(REG0_REG_3__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U3159 ( .A1(n2521), .A2(REG1_REG_3__SCAN_IN), .ZN(n2522) );
  NAND2_X1 U3160 ( .A1(n3821), .A2(n2533), .ZN(n2531) );
  NAND2_X1 U3161 ( .A1(n2526), .A2(IR_REG_31__SCAN_IN), .ZN(n2528) );
  NAND2_X1 U3162 ( .A1(n2528), .A2(n2527), .ZN(n2544) );
  OR2_X1 U3163 ( .A1(n2528), .A2(n2527), .ZN(n2529) );
  MUX2_X1 U3164 ( .A(n4324), .B(DATAI_3_), .S(n3716), .Z(n3007) );
  NAND2_X1 U3165 ( .A1(n3007), .A2(n2885), .ZN(n2530) );
  NAND2_X1 U3166 ( .A1(n2531), .A2(n2530), .ZN(n2532) );
  AOI22_X1 U3167 ( .A1(n3821), .A2(n2891), .B1(n2890), .B2(n3007), .ZN(n2535)
         );
  XNOR2_X1 U3168 ( .A(n2534), .B(n2535), .ZN(n3143) );
  INV_X1 U3169 ( .A(n2534), .ZN(n2536) );
  NAND2_X1 U3170 ( .A1(n2536), .A2(n2535), .ZN(n2537) );
  NAND2_X1 U3171 ( .A1(n2506), .A2(REG0_REG_4__SCAN_IN), .ZN(n2543) );
  INV_X1 U3172 ( .A(REG3_REG_4__SCAN_IN), .ZN(n4728) );
  XNOR2_X1 U3173 ( .A(n4728), .B(REG3_REG_3__SCAN_IN), .ZN(n3235) );
  NAND2_X1 U3174 ( .A1(n2856), .A2(n3235), .ZN(n2542) );
  NAND2_X1 U3175 ( .A1(n3712), .A2(REG1_REG_4__SCAN_IN), .ZN(n2541) );
  INV_X1 U3176 ( .A(REG2_REG_4__SCAN_IN), .ZN(n3285) );
  OR2_X1 U3177 ( .A1(n2171), .A2(n3285), .ZN(n2540) );
  NAND2_X1 U3178 ( .A1(n2544), .A2(IR_REG_31__SCAN_IN), .ZN(n2545) );
  XNOR2_X1 U3179 ( .A(n2545), .B(IR_REG_4__SCAN_IN), .ZN(n4323) );
  MUX2_X1 U3180 ( .A(n4323), .B(DATAI_4_), .S(n3716), .Z(n3180) );
  INV_X1 U3181 ( .A(n3180), .ZN(n3228) );
  XNOR2_X1 U3182 ( .A(n2546), .B(n2862), .ZN(n2548) );
  OAI22_X1 U3183 ( .A1(n3213), .A2(n2875), .B1(n2873), .B2(n3228), .ZN(n2547)
         );
  XNOR2_X1 U3184 ( .A(n2548), .B(n2547), .ZN(n3232) );
  NAND2_X1 U3185 ( .A1(n2548), .A2(n2547), .ZN(n2549) );
  INV_X1 U3186 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2550) );
  OR2_X1 U3187 ( .A1(n2171), .A2(n2550), .ZN(n2556) );
  NAND2_X1 U3188 ( .A1(n2506), .A2(REG0_REG_5__SCAN_IN), .ZN(n2555) );
  OAI21_X1 U3189 ( .B1(n2551), .B2(REG3_REG_5__SCAN_IN), .A(n2568), .ZN(n3218)
         );
  INV_X1 U3190 ( .A(n3218), .ZN(n2552) );
  NAND2_X1 U3191 ( .A1(n2856), .A2(n2552), .ZN(n2554) );
  NAND2_X1 U3192 ( .A1(n2521), .A2(REG1_REG_5__SCAN_IN), .ZN(n2553) );
  NAND4_X1 U3193 ( .A1(n2556), .A2(n2555), .A3(n2554), .A4(n2553), .ZN(n3820)
         );
  NAND2_X1 U3194 ( .A1(n3820), .A2(n2890), .ZN(n2562) );
  NAND2_X1 U3195 ( .A1(n2557), .A2(IR_REG_31__SCAN_IN), .ZN(n2558) );
  MUX2_X1 U3196 ( .A(IR_REG_31__SCAN_IN), .B(n2558), .S(IR_REG_5__SCAN_IN), 
        .Z(n2560) );
  INV_X1 U3197 ( .A(n2626), .ZN(n2559) );
  MUX2_X1 U3198 ( .A(n3281), .B(DATAI_5_), .S(n3716), .Z(n3215) );
  NAND2_X1 U3199 ( .A1(n3215), .A2(n2885), .ZN(n2561) );
  NAND2_X1 U3200 ( .A1(n2562), .A2(n2561), .ZN(n2563) );
  XNOR2_X1 U3201 ( .A(n2563), .B(n2862), .ZN(n2566) );
  AOI22_X1 U3202 ( .A1(n3820), .A2(n2891), .B1(n2890), .B2(n3215), .ZN(n2564)
         );
  XNOR2_X1 U3203 ( .A(n2566), .B(n2564), .ZN(n3209) );
  INV_X1 U3204 ( .A(n2564), .ZN(n2565) );
  NAND2_X1 U3205 ( .A1(n2566), .A2(n2565), .ZN(n2567) );
  INV_X1 U3206 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3259) );
  OR2_X1 U3207 ( .A1(n2171), .A2(n3259), .ZN(n2573) );
  NAND2_X1 U3208 ( .A1(n2506), .A2(REG0_REG_6__SCAN_IN), .ZN(n2572) );
  AND2_X1 U3209 ( .A1(n2568), .A2(n3241), .ZN(n2569) );
  NOR2_X1 U32100 ( .A1(n2580), .A2(n2569), .ZN(n3257) );
  NAND2_X1 U32110 ( .A1(n2856), .A2(n3257), .ZN(n2571) );
  NAND2_X1 U32120 ( .A1(n2521), .A2(REG1_REG_6__SCAN_IN), .ZN(n2570) );
  NAND4_X1 U32130 ( .A1(n2573), .A2(n2572), .A3(n2571), .A4(n2570), .ZN(n3819)
         );
  NAND2_X1 U32140 ( .A1(n3819), .A2(n2891), .ZN(n2576) );
  OR2_X1 U32150 ( .A1(n2626), .A2(n2768), .ZN(n2574) );
  XNOR2_X1 U32160 ( .A(n2574), .B(IR_REG_6__SCAN_IN), .ZN(n4525) );
  MUX2_X1 U32170 ( .A(n4525), .B(DATAI_6_), .S(n3716), .Z(n3248) );
  NAND2_X1 U32180 ( .A1(n3248), .A2(n2890), .ZN(n2575) );
  NAND2_X1 U32190 ( .A1(n2576), .A2(n2575), .ZN(n3238) );
  NAND2_X1 U32200 ( .A1(n3819), .A2(n2890), .ZN(n2578) );
  NAND2_X1 U32210 ( .A1(n3248), .A2(n2885), .ZN(n2577) );
  NAND2_X1 U32220 ( .A1(n2578), .A2(n2577), .ZN(n2579) );
  XNOR2_X1 U32230 ( .A(n2579), .B(n2862), .ZN(n3237) );
  NAND2_X1 U32240 ( .A1(n2506), .A2(REG0_REG_7__SCAN_IN), .ZN(n2586) );
  NAND2_X1 U32250 ( .A1(n2580), .A2(REG3_REG_7__SCAN_IN), .ZN(n2597) );
  OR2_X1 U32260 ( .A1(n2580), .A2(REG3_REG_7__SCAN_IN), .ZN(n2581) );
  AND2_X1 U32270 ( .A1(n2597), .A2(n2581), .ZN(n3321) );
  NAND2_X1 U32280 ( .A1(n2856), .A2(n3321), .ZN(n2585) );
  NAND2_X1 U32290 ( .A1(n2521), .A2(REG1_REG_7__SCAN_IN), .ZN(n2584) );
  INV_X1 U32300 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2582) );
  OR2_X1 U32310 ( .A1(n2171), .A2(n2582), .ZN(n2583) );
  INV_X1 U32320 ( .A(IR_REG_6__SCAN_IN), .ZN(n2587) );
  NAND2_X1 U32330 ( .A1(n2626), .A2(n2587), .ZN(n2588) );
  NAND2_X1 U32340 ( .A1(n2588), .A2(IR_REG_31__SCAN_IN), .ZN(n2590) );
  INV_X1 U32350 ( .A(IR_REG_7__SCAN_IN), .ZN(n2589) );
  NAND2_X1 U32360 ( .A1(n2590), .A2(n2589), .ZN(n2603) );
  OR2_X1 U32370 ( .A1(n2590), .A2(n2589), .ZN(n2591) );
  MUX2_X1 U32380 ( .A(n3280), .B(DATAI_7_), .S(n3716), .Z(n3320) );
  OAI22_X1 U32390 ( .A1(n3347), .A2(n2873), .B1(n2872), .B2(n3314), .ZN(n2592)
         );
  XNOR2_X1 U32400 ( .A(n2592), .B(n2888), .ZN(n2593) );
  OAI22_X1 U32410 ( .A1(n3347), .A2(n2875), .B1(n2873), .B2(n3314), .ZN(n2594)
         );
  XNOR2_X1 U32420 ( .A(n2593), .B(n2594), .ZN(n3306) );
  INV_X1 U32430 ( .A(n2593), .ZN(n2595) );
  NAND2_X1 U32440 ( .A1(n2595), .A2(n2594), .ZN(n2596) );
  INV_X1 U32450 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3355) );
  OR2_X1 U32460 ( .A1(n2171), .A2(n3355), .ZN(n2602) );
  NAND2_X1 U32470 ( .A1(n2506), .A2(REG0_REG_8__SCAN_IN), .ZN(n2601) );
  NAND2_X1 U32480 ( .A1(n2597), .A2(n3337), .ZN(n2598) );
  AND2_X1 U32490 ( .A1(n2616), .A2(n2598), .ZN(n3353) );
  NAND2_X1 U32500 ( .A1(n2856), .A2(n3353), .ZN(n2600) );
  NAND2_X1 U32510 ( .A1(n3712), .A2(REG1_REG_8__SCAN_IN), .ZN(n2599) );
  NAND4_X1 U32520 ( .A1(n2602), .A2(n2601), .A3(n2600), .A4(n2599), .ZN(n3817)
         );
  NAND2_X1 U32530 ( .A1(n3817), .A2(n2533), .ZN(n2606) );
  NAND2_X1 U32540 ( .A1(n2603), .A2(IR_REG_31__SCAN_IN), .ZN(n2604) );
  XNOR2_X1 U32550 ( .A(n2604), .B(IR_REG_8__SCAN_IN), .ZN(n3290) );
  MUX2_X1 U32560 ( .A(n3290), .B(DATAI_8_), .S(n3716), .Z(n3345) );
  NAND2_X1 U32570 ( .A1(n3345), .A2(n2885), .ZN(n2605) );
  NAND2_X1 U32580 ( .A1(n2606), .A2(n2605), .ZN(n2607) );
  XNOR2_X1 U32590 ( .A(n2607), .B(n2862), .ZN(n2610) );
  NAND2_X1 U32600 ( .A1(n3817), .A2(n2891), .ZN(n2609) );
  NAND2_X1 U32610 ( .A1(n3345), .A2(n2533), .ZN(n2608) );
  NAND2_X1 U32620 ( .A1(n2609), .A2(n2608), .ZN(n2611) );
  AND2_X1 U32630 ( .A1(n2610), .A2(n2611), .ZN(n3335) );
  INV_X1 U32640 ( .A(n2610), .ZN(n2613) );
  INV_X1 U32650 ( .A(n2611), .ZN(n2612) );
  NAND2_X1 U32660 ( .A1(n2613), .A2(n2612), .ZN(n3334) );
  INV_X1 U32670 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2614) );
  OR2_X1 U32680 ( .A1(n2171), .A2(n2614), .ZN(n2622) );
  AND2_X1 U32690 ( .A1(n2616), .A2(n2615), .ZN(n2617) );
  OR2_X1 U32700 ( .A1(n2617), .A2(n2631), .ZN(n3397) );
  INV_X1 U32710 ( .A(n3397), .ZN(n2618) );
  NAND2_X1 U32720 ( .A1(n2856), .A2(n2618), .ZN(n2621) );
  NAND2_X1 U32730 ( .A1(n2506), .A2(REG0_REG_9__SCAN_IN), .ZN(n2620) );
  NAND2_X1 U32740 ( .A1(n3712), .A2(REG1_REG_9__SCAN_IN), .ZN(n2619) );
  NAND4_X1 U32750 ( .A1(n2622), .A2(n2621), .A3(n2620), .A4(n2619), .ZN(n3816)
         );
  NAND2_X1 U32760 ( .A1(n3816), .A2(n2533), .ZN(n2629) );
  INV_X1 U32770 ( .A(IR_REG_8__SCAN_IN), .ZN(n2623) );
  AND2_X1 U32780 ( .A1(n2624), .A2(n2623), .ZN(n2625) );
  OR2_X1 U32790 ( .A1(n2639), .A2(n2768), .ZN(n2627) );
  XNOR2_X1 U32800 ( .A(n2627), .B(IR_REG_9__SCAN_IN), .ZN(n3279) );
  MUX2_X1 U32810 ( .A(n3279), .B(DATAI_9_), .S(n3716), .Z(n3394) );
  NAND2_X1 U32820 ( .A1(n3394), .A2(n2885), .ZN(n2628) );
  NAND2_X1 U32830 ( .A1(n2629), .A2(n2628), .ZN(n2630) );
  XNOR2_X1 U32840 ( .A(n2630), .B(n2862), .ZN(n2644) );
  AOI22_X1 U32850 ( .A1(n3816), .A2(n2891), .B1(n2890), .B2(n3394), .ZN(n2645)
         );
  XNOR2_X1 U32860 ( .A(n2644), .B(n2645), .ZN(n3389) );
  INV_X1 U32870 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3384) );
  OR2_X1 U32880 ( .A1(n2171), .A2(n3384), .ZN(n2637) );
  NAND2_X1 U32890 ( .A1(n2506), .A2(REG0_REG_10__SCAN_IN), .ZN(n2636) );
  NOR2_X1 U32900 ( .A1(n2631), .A2(REG3_REG_10__SCAN_IN), .ZN(n2632) );
  OR2_X1 U32910 ( .A1(n2651), .A2(n2632), .ZN(n3416) );
  INV_X1 U32920 ( .A(n3416), .ZN(n2633) );
  NAND2_X1 U32930 ( .A1(n2856), .A2(n2633), .ZN(n2635) );
  NAND2_X1 U32940 ( .A1(n2521), .A2(REG1_REG_10__SCAN_IN), .ZN(n2634) );
  NAND4_X1 U32950 ( .A1(n2637), .A2(n2636), .A3(n2635), .A4(n2634), .ZN(n3815)
         );
  NAND2_X1 U32960 ( .A1(n3815), .A2(n2890), .ZN(n2642) );
  INV_X1 U32970 ( .A(IR_REG_9__SCAN_IN), .ZN(n2638) );
  NAND2_X1 U32980 ( .A1(n2639), .A2(n2638), .ZN(n2658) );
  NAND2_X1 U32990 ( .A1(n2658), .A2(IR_REG_31__SCAN_IN), .ZN(n2640) );
  XNOR2_X1 U33000 ( .A(n2640), .B(IR_REG_10__SCAN_IN), .ZN(n4519) );
  MUX2_X1 U33010 ( .A(n4519), .B(DATAI_10_), .S(n3716), .Z(n3413) );
  NAND2_X1 U33020 ( .A1(n3413), .A2(n2885), .ZN(n2641) );
  NAND2_X1 U33030 ( .A1(n2642), .A2(n2641), .ZN(n2643) );
  XNOR2_X1 U33040 ( .A(n2643), .B(n2862), .ZN(n2649) );
  AOI22_X1 U33050 ( .A1(n3815), .A2(n2891), .B1(n2890), .B2(n3413), .ZN(n2647)
         );
  XNOR2_X1 U33060 ( .A(n2649), .B(n2647), .ZN(n3407) );
  INV_X1 U33070 ( .A(n2644), .ZN(n2646) );
  NAND2_X1 U33080 ( .A1(n2646), .A2(n2645), .ZN(n3404) );
  INV_X1 U33090 ( .A(n2647), .ZN(n2648) );
  NAND2_X1 U33100 ( .A1(n2649), .A2(n2648), .ZN(n2650) );
  INV_X1 U33110 ( .A(n3437), .ZN(n2683) );
  NAND2_X1 U33120 ( .A1(n2506), .A2(REG0_REG_11__SCAN_IN), .ZN(n2657) );
  OR2_X1 U33130 ( .A1(n2651), .A2(REG3_REG_11__SCAN_IN), .ZN(n2652) );
  AND2_X1 U33140 ( .A1(n2664), .A2(n2652), .ZN(n4467) );
  NAND2_X1 U33150 ( .A1(n2507), .A2(n4467), .ZN(n2656) );
  NAND2_X1 U33160 ( .A1(n3712), .A2(REG1_REG_11__SCAN_IN), .ZN(n2655) );
  INV_X1 U33170 ( .A(REG2_REG_11__SCAN_IN), .ZN(n2653) );
  OR2_X1 U33180 ( .A1(n2171), .A2(n2653), .ZN(n2654) );
  NAND2_X1 U33190 ( .A1(n2659), .A2(IR_REG_31__SCAN_IN), .ZN(n2660) );
  OR2_X1 U33200 ( .A1(n2660), .A2(n4763), .ZN(n2661) );
  NAND2_X1 U33210 ( .A1(n2660), .A2(n4763), .ZN(n2671) );
  MUX2_X1 U33220 ( .A(n3278), .B(DATAI_11_), .S(n3716), .Z(n3041) );
  OAI22_X1 U33230 ( .A1(n3411), .A2(n2873), .B1(n2872), .B2(n4469), .ZN(n2662)
         );
  XNOR2_X1 U33240 ( .A(n2662), .B(n2862), .ZN(n2678) );
  OAI22_X1 U33250 ( .A1(n3411), .A2(n2875), .B1(n2873), .B2(n4469), .ZN(n2679)
         );
  AND2_X1 U33260 ( .A1(n2678), .A2(n2679), .ZN(n3436) );
  NAND2_X1 U33270 ( .A1(n2506), .A2(REG0_REG_12__SCAN_IN), .ZN(n2670) );
  NAND2_X1 U33280 ( .A1(n2664), .A2(n2663), .ZN(n2665) );
  AND2_X1 U33290 ( .A1(n2684), .A2(n2665), .ZN(n3448) );
  NAND2_X1 U33300 ( .A1(n2856), .A2(n3448), .ZN(n2669) );
  NAND2_X1 U33310 ( .A1(n3712), .A2(REG1_REG_12__SCAN_IN), .ZN(n2668) );
  INV_X1 U33320 ( .A(REG2_REG_12__SCAN_IN), .ZN(n2666) );
  OR2_X1 U33330 ( .A1(n2171), .A2(n2666), .ZN(n2667) );
  NAND2_X1 U33340 ( .A1(n2671), .A2(IR_REG_31__SCAN_IN), .ZN(n2672) );
  XNOR2_X1 U33350 ( .A(n2672), .B(IR_REG_12__SCAN_IN), .ZN(n3297) );
  INV_X1 U33360 ( .A(DATAI_12_), .ZN(n2673) );
  MUX2_X1 U33370 ( .A(n4517), .B(n2673), .S(n3716), .Z(n3446) );
  OAI22_X1 U33380 ( .A1(n3016), .A2(n2873), .B1(n2872), .B2(n3446), .ZN(n2674)
         );
  XNOR2_X1 U33390 ( .A(n2674), .B(n2888), .ZN(n3441) );
  INV_X1 U33400 ( .A(n3441), .ZN(n2677) );
  NOR2_X1 U33410 ( .A1(n3446), .A2(n2873), .ZN(n2675) );
  AOI21_X1 U33420 ( .B1(n4463), .B2(n2891), .A(n2675), .ZN(n3440) );
  INV_X1 U33430 ( .A(n3440), .ZN(n2676) );
  INV_X1 U33440 ( .A(n2678), .ZN(n2681) );
  INV_X1 U33450 ( .A(n2679), .ZN(n2680) );
  NAND2_X1 U33460 ( .A1(n2681), .A2(n2680), .ZN(n3438) );
  AND2_X1 U33470 ( .A1(n2429), .A2(n3438), .ZN(n2682) );
  NAND2_X1 U33480 ( .A1(n2506), .A2(REG0_REG_13__SCAN_IN), .ZN(n2690) );
  NAND2_X1 U33490 ( .A1(n2684), .A2(n3276), .ZN(n2685) );
  AND2_X1 U33500 ( .A1(n2710), .A2(n2685), .ZN(n3481) );
  NAND2_X1 U33510 ( .A1(n2856), .A2(n3481), .ZN(n2689) );
  NAND2_X1 U33520 ( .A1(n3712), .A2(REG1_REG_13__SCAN_IN), .ZN(n2688) );
  INV_X1 U3353 ( .A(REG2_REG_13__SCAN_IN), .ZN(n2686) );
  OR2_X1 U33540 ( .A1(n2171), .A2(n2686), .ZN(n2687) );
  NOR2_X1 U3355 ( .A1(n2691), .A2(n2768), .ZN(n2692) );
  MUX2_X1 U3356 ( .A(n2768), .B(n2692), .S(IR_REG_13__SCAN_IN), .Z(n2695) );
  NAND2_X1 U3357 ( .A1(n2691), .A2(n2693), .ZN(n2749) );
  INV_X1 U3358 ( .A(n2749), .ZN(n2694) );
  INV_X1 U3359 ( .A(DATAI_13_), .ZN(n4711) );
  MUX2_X1 U3360 ( .A(n3870), .B(n4711), .S(n3716), .Z(n3472) );
  OAI22_X1 U3361 ( .A1(n4155), .A2(n2873), .B1(n2872), .B2(n3472), .ZN(n2696)
         );
  XNOR2_X1 U3362 ( .A(n2696), .B(n2862), .ZN(n2697) );
  OAI22_X1 U3363 ( .A1(n4155), .A2(n2875), .B1(n2873), .B2(n3472), .ZN(n2698)
         );
  AND2_X1 U3364 ( .A1(n2697), .A2(n2698), .ZN(n3452) );
  INV_X1 U3365 ( .A(n2697), .ZN(n2700) );
  INV_X1 U3366 ( .A(n2698), .ZN(n2699) );
  NAND2_X1 U3367 ( .A1(n2700), .A2(n2699), .ZN(n3451) );
  NAND2_X1 U3368 ( .A1(n2506), .A2(REG0_REG_14__SCAN_IN), .ZN(n2705) );
  XNOR2_X1 U3369 ( .A(n2710), .B(REG3_REG_14__SCAN_IN), .ZN(n4165) );
  NAND2_X1 U3370 ( .A1(n2856), .A2(n4165), .ZN(n2704) );
  NAND2_X1 U3371 ( .A1(n3712), .A2(REG1_REG_14__SCAN_IN), .ZN(n2703) );
  INV_X1 U3372 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4168) );
  OR2_X1 U3373 ( .A1(n2171), .A2(n4168), .ZN(n2702) );
  NAND2_X1 U3374 ( .A1(n2749), .A2(IR_REG_31__SCAN_IN), .ZN(n2706) );
  XNOR2_X1 U3375 ( .A(n2706), .B(IR_REG_14__SCAN_IN), .ZN(n3874) );
  MUX2_X1 U3376 ( .A(n3874), .B(DATAI_14_), .S(n3716), .Z(n4164) );
  OAI22_X1 U3377 ( .A1(n3473), .A2(n2873), .B1(n2872), .B2(n3498), .ZN(n2707)
         );
  OAI22_X1 U3378 ( .A1(n3473), .A2(n2875), .B1(n2873), .B2(n3498), .ZN(n3493)
         );
  INV_X1 U3379 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3510) );
  OR2_X1 U3380 ( .A1(n2171), .A2(n3510), .ZN(n2715) );
  NAND2_X1 U3381 ( .A1(n2506), .A2(REG0_REG_15__SCAN_IN), .ZN(n2714) );
  INV_X1 U3382 ( .A(n2710), .ZN(n2708) );
  AOI21_X1 U3383 ( .B1(n2708), .B2(REG3_REG_14__SCAN_IN), .A(
        REG3_REG_15__SCAN_IN), .ZN(n2711) );
  NAND2_X1 U3384 ( .A1(REG3_REG_14__SCAN_IN), .A2(REG3_REG_15__SCAN_IN), .ZN(
        n2709) );
  OR2_X1 U3385 ( .A1(n2711), .A2(n2725), .ZN(n3509) );
  INV_X1 U3386 ( .A(n3509), .ZN(n3646) );
  NAND2_X1 U3387 ( .A1(n2856), .A2(n3646), .ZN(n2713) );
  NAND2_X1 U3388 ( .A1(n3712), .A2(REG1_REG_15__SCAN_IN), .ZN(n2712) );
  NAND4_X1 U3389 ( .A1(n2715), .A2(n2714), .A3(n2713), .A4(n2712), .ZN(n4153)
         );
  NAND2_X1 U3390 ( .A1(n4153), .A2(n2890), .ZN(n2721) );
  NAND2_X1 U3391 ( .A1(n2716), .A2(IR_REG_31__SCAN_IN), .ZN(n2718) );
  INV_X1 U3392 ( .A(IR_REG_15__SCAN_IN), .ZN(n2717) );
  OR2_X1 U3393 ( .A1(n2718), .A2(n2717), .ZN(n2719) );
  NAND2_X1 U3394 ( .A1(n2718), .A2(n2717), .ZN(n2731) );
  MUX2_X1 U3395 ( .A(n3877), .B(DATAI_15_), .S(n3716), .Z(n3019) );
  NAND2_X1 U3396 ( .A1(n3019), .A2(n2885), .ZN(n2720) );
  NAND2_X1 U3397 ( .A1(n2721), .A2(n2720), .ZN(n2722) );
  XNOR2_X1 U3398 ( .A(n2722), .B(n2888), .ZN(n2735) );
  NAND2_X1 U3399 ( .A1(n4153), .A2(n2891), .ZN(n2724) );
  NAND2_X1 U3400 ( .A1(n3019), .A2(n2890), .ZN(n2723) );
  NAND2_X1 U3401 ( .A1(n2724), .A2(n2723), .ZN(n3640) );
  NAND2_X1 U3402 ( .A1(n2506), .A2(REG0_REG_16__SCAN_IN), .ZN(n2730) );
  OR2_X1 U3403 ( .A1(n2725), .A2(REG3_REG_16__SCAN_IN), .ZN(n2726) );
  NAND2_X1 U3404 ( .A1(n2725), .A2(REG3_REG_16__SCAN_IN), .ZN(n2740) );
  AND2_X1 U3405 ( .A1(n2726), .A2(n2740), .ZN(n4143) );
  NAND2_X1 U3406 ( .A1(n2856), .A2(n4143), .ZN(n2729) );
  NAND2_X1 U3407 ( .A1(n3712), .A2(REG1_REG_16__SCAN_IN), .ZN(n2728) );
  OR2_X1 U3408 ( .A1(n2171), .A2(n4435), .ZN(n2727) );
  NAND2_X1 U3409 ( .A1(n2731), .A2(IR_REG_31__SCAN_IN), .ZN(n2732) );
  XNOR2_X1 U3410 ( .A(n2732), .B(IR_REG_16__SCAN_IN), .ZN(n3878) );
  MUX2_X1 U3411 ( .A(n3878), .B(DATAI_16_), .S(n3716), .Z(n4142) );
  OAI22_X1 U3412 ( .A1(n4927), .A2(n2873), .B1(n2872), .B2(n3580), .ZN(n2733)
         );
  XNOR2_X1 U3413 ( .A(n2733), .B(n2888), .ZN(n2738) );
  OAI22_X1 U3414 ( .A1(n4927), .A2(n2875), .B1(n2873), .B2(n3580), .ZN(n2736)
         );
  XNOR2_X1 U3415 ( .A(n2738), .B(n2736), .ZN(n3576) );
  INV_X1 U3416 ( .A(n2736), .ZN(n2737) );
  INV_X1 U3417 ( .A(n4925), .ZN(n2759) );
  NAND2_X1 U3418 ( .A1(n2506), .A2(REG0_REG_17__SCAN_IN), .ZN(n2745) );
  INV_X1 U3419 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2739) );
  NAND2_X1 U3420 ( .A1(n2740), .A2(n2739), .ZN(n2741) );
  AND2_X1 U3421 ( .A1(n2761), .A2(n2741), .ZN(n4932) );
  NAND2_X1 U3422 ( .A1(n2507), .A2(n4932), .ZN(n2744) );
  NAND2_X1 U3423 ( .A1(n3712), .A2(REG1_REG_17__SCAN_IN), .ZN(n2743) );
  INV_X1 U3424 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4855) );
  OR2_X1 U3425 ( .A1(n2539), .A2(n4855), .ZN(n2742) );
  NAND2_X1 U3426 ( .A1(n2747), .A2(n2746), .ZN(n2748) );
  OAI21_X1 U3427 ( .B1(n2749), .B2(n2748), .A(IR_REG_31__SCAN_IN), .ZN(n2750)
         );
  MUX2_X1 U3428 ( .A(IR_REG_31__SCAN_IN), .B(n2750), .S(IR_REG_17__SCAN_IN), 
        .Z(n2753) );
  INV_X1 U3429 ( .A(n2751), .ZN(n2752) );
  NAND2_X1 U3430 ( .A1(n2753), .A2(n2752), .ZN(n3884) );
  INV_X1 U3431 ( .A(DATAI_17_), .ZN(n2754) );
  MUX2_X1 U3432 ( .A(n3884), .B(n2754), .S(n3716), .Z(n4936) );
  NOR2_X1 U3433 ( .A1(n4936), .A2(n2873), .ZN(n2755) );
  AOI21_X1 U3434 ( .B1(n4137), .B2(n2891), .A(n2755), .ZN(n2757) );
  INV_X1 U3435 ( .A(n2757), .ZN(n4922) );
  OAI22_X1 U3436 ( .A1(n4104), .A2(n2873), .B1(n2872), .B2(n4936), .ZN(n2756)
         );
  XOR2_X1 U3437 ( .A(n2862), .B(n2756), .Z(n4923) );
  AOI21_X1 U3438 ( .B1(n4925), .B2(n2757), .A(n4923), .ZN(n2758) );
  AOI21_X1 U3439 ( .B1(n2759), .B2(n4922), .A(n2758), .ZN(n3619) );
  NAND2_X1 U3440 ( .A1(n2506), .A2(REG0_REG_18__SCAN_IN), .ZN(n2767) );
  INV_X1 U3441 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2760) );
  AND2_X1 U3442 ( .A1(n2761), .A2(n2760), .ZN(n2762) );
  NOR2_X1 U3443 ( .A1(n2774), .A2(n2762), .ZN(n4113) );
  NAND2_X1 U3444 ( .A1(n2856), .A2(n4113), .ZN(n2766) );
  NAND2_X1 U3445 ( .A1(n3712), .A2(REG1_REG_18__SCAN_IN), .ZN(n2765) );
  INV_X1 U3446 ( .A(REG2_REG_18__SCAN_IN), .ZN(n2763) );
  OR2_X1 U3447 ( .A1(n2171), .A2(n2763), .ZN(n2764) );
  OR2_X1 U3448 ( .A1(n2751), .A2(n2768), .ZN(n2769) );
  XNOR2_X1 U3449 ( .A(n2769), .B(IR_REG_18__SCAN_IN), .ZN(n3894) );
  MUX2_X1 U3450 ( .A(n3894), .B(DATAI_18_), .S(n3716), .Z(n4101) );
  OAI22_X1 U3451 ( .A1(n4120), .A2(n2873), .B1(n2872), .B2(n4112), .ZN(n2770)
         );
  XNOR2_X1 U3452 ( .A(n2770), .B(n2862), .ZN(n2772) );
  OAI22_X1 U3453 ( .A1(n4120), .A2(n2875), .B1(n2873), .B2(n4112), .ZN(n2771)
         );
  NAND2_X1 U3454 ( .A1(n2772), .A2(n2771), .ZN(n3616) );
  NOR2_X1 U3455 ( .A1(n2772), .A2(n2771), .ZN(n3615) );
  AOI21_X1 U3456 ( .B1(n3619), .B2(n3616), .A(n3615), .ZN(n3548) );
  INV_X1 U3457 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2773) );
  OR2_X1 U34580 ( .A1(n2171), .A2(n2773), .ZN(n2779) );
  NAND2_X1 U34590 ( .A1(n2506), .A2(REG0_REG_19__SCAN_IN), .ZN(n2778) );
  NOR2_X1 U3460 ( .A1(n2774), .A2(REG3_REG_19__SCAN_IN), .ZN(n2775) );
  NOR2_X1 U3461 ( .A1(n2785), .A2(n2775), .ZN(n4094) );
  NAND2_X1 U3462 ( .A1(n2856), .A2(n4094), .ZN(n2777) );
  NAND2_X1 U3463 ( .A1(n3712), .A2(REG1_REG_19__SCAN_IN), .ZN(n2776) );
  NAND2_X1 U3464 ( .A1(n4102), .A2(n2890), .ZN(n2781) );
  MUX2_X1 U3465 ( .A(n4320), .B(DATAI_19_), .S(n3716), .Z(n4091) );
  NAND2_X1 U3466 ( .A1(n4091), .A2(n2885), .ZN(n2780) );
  NAND2_X1 U34670 ( .A1(n2781), .A2(n2780), .ZN(n2782) );
  XNOR2_X1 U3468 ( .A(n2782), .B(n2862), .ZN(n2784) );
  OAI22_X1 U34690 ( .A1(n3621), .A2(n2875), .B1(n2873), .B2(n4085), .ZN(n2783)
         );
  XNOR2_X1 U3470 ( .A(n2784), .B(n2783), .ZN(n3549) );
  OAI22_X1 U34710 ( .A1(n3548), .A2(n3549), .B1(n2784), .B2(n2783), .ZN(n3596)
         );
  INV_X1 U3472 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4074) );
  OR2_X1 U34730 ( .A1(n2171), .A2(n4074), .ZN(n2790) );
  NAND2_X1 U3474 ( .A1(n2506), .A2(REG0_REG_20__SCAN_IN), .ZN(n2789) );
  OR2_X1 U34750 ( .A1(n2785), .A2(REG3_REG_20__SCAN_IN), .ZN(n2786) );
  AND2_X1 U3476 ( .A1(n2801), .A2(n2786), .ZN(n4072) );
  NAND2_X1 U34770 ( .A1(n2856), .A2(n4072), .ZN(n2788) );
  NAND2_X1 U3478 ( .A1(n3712), .A2(REG1_REG_20__SCAN_IN), .ZN(n2787) );
  NAND2_X1 U34790 ( .A1(n4041), .A2(n2890), .ZN(n2792) );
  NAND2_X1 U3480 ( .A1(n4071), .A2(n2885), .ZN(n2791) );
  NAND2_X1 U34810 ( .A1(n2792), .A2(n2791), .ZN(n2793) );
  XNOR2_X1 U3482 ( .A(n2793), .B(n2862), .ZN(n2796) );
  NAND2_X1 U34830 ( .A1(n4041), .A2(n2891), .ZN(n2795) );
  NAND2_X1 U3484 ( .A1(n4071), .A2(n2890), .ZN(n2794) );
  NAND2_X1 U34850 ( .A1(n2795), .A2(n2794), .ZN(n2797) );
  NAND2_X1 U3486 ( .A1(n2796), .A2(n2797), .ZN(n3597) );
  NAND2_X1 U34870 ( .A1(n3596), .A2(n3597), .ZN(n3595) );
  INV_X1 U3488 ( .A(n2796), .ZN(n2799) );
  INV_X1 U34890 ( .A(n2797), .ZN(n2798) );
  NAND2_X1 U3490 ( .A1(n2799), .A2(n2798), .ZN(n3599) );
  NAND2_X1 U34910 ( .A1(n3595), .A2(n3599), .ZN(n3558) );
  INV_X1 U3492 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4051) );
  OR2_X1 U34930 ( .A1(n2171), .A2(n4051), .ZN(n2806) );
  NAND2_X1 U3494 ( .A1(n2506), .A2(REG0_REG_21__SCAN_IN), .ZN(n2805) );
  INV_X1 U34950 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2800) );
  NAND2_X1 U3496 ( .A1(n2801), .A2(n2800), .ZN(n2802) );
  AND2_X1 U34970 ( .A1(n2815), .A2(n2802), .ZN(n4049) );
  NAND2_X1 U3498 ( .A1(n2856), .A2(n4049), .ZN(n2804) );
  NAND2_X1 U34990 ( .A1(n3712), .A2(REG1_REG_21__SCAN_IN), .ZN(n2803) );
  NAND2_X1 U3500 ( .A1(n4063), .A2(n2890), .ZN(n2808) );
  NAND2_X1 U35010 ( .A1(n4039), .A2(n2885), .ZN(n2807) );
  NAND2_X1 U3502 ( .A1(n2808), .A2(n2807), .ZN(n2809) );
  XNOR2_X1 U35030 ( .A(n2809), .B(n2862), .ZN(n3556) );
  NAND2_X1 U3504 ( .A1(n4063), .A2(n2891), .ZN(n2811) );
  NAND2_X1 U35050 ( .A1(n4039), .A2(n2890), .ZN(n2810) );
  NAND2_X1 U35060 ( .A1(n2811), .A2(n2810), .ZN(n3555) );
  NOR2_X1 U35070 ( .A1(n3556), .A2(n3555), .ZN(n2814) );
  INV_X1 U35080 ( .A(n3556), .ZN(n2813) );
  INV_X1 U35090 ( .A(n3555), .ZN(n2812) );
  INV_X1 U35100 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4835) );
  AND2_X1 U35110 ( .A1(n2815), .A2(n4835), .ZN(n2816) );
  OR2_X1 U35120 ( .A1(n2816), .A2(n2825), .ZN(n4029) );
  AOI22_X1 U35130 ( .A1(n2492), .A2(REG2_REG_22__SCAN_IN), .B1(n2506), .B2(
        REG0_REG_22__SCAN_IN), .ZN(n2818) );
  NAND2_X1 U35140 ( .A1(n3712), .A2(REG1_REG_22__SCAN_IN), .ZN(n2817) );
  INV_X1 U35150 ( .A(n4026), .ZN(n2997) );
  AOI22_X1 U35160 ( .A1(n4040), .A2(n2891), .B1(n2890), .B2(n2997), .ZN(n2822)
         );
  NAND2_X1 U35170 ( .A1(n4040), .A2(n2890), .ZN(n2820) );
  NAND2_X1 U35180 ( .A1(n2997), .A2(n2885), .ZN(n2819) );
  NAND2_X1 U35190 ( .A1(n2820), .A2(n2819), .ZN(n2821) );
  XNOR2_X1 U35200 ( .A(n2821), .B(n2862), .ZN(n2824) );
  XOR2_X1 U35210 ( .A(n2822), .B(n2824), .Z(n3608) );
  INV_X1 U35220 ( .A(n2822), .ZN(n2823) );
  NOR2_X1 U35230 ( .A1(n2824), .A2(n2823), .ZN(n3542) );
  NOR2_X1 U35240 ( .A1(n2825), .A2(REG3_REG_23__SCAN_IN), .ZN(n2826) );
  OR2_X1 U35250 ( .A1(n2835), .A2(n2826), .ZN(n4009) );
  AOI22_X1 U35260 ( .A1(n2492), .A2(REG2_REG_23__SCAN_IN), .B1(n2506), .B2(
        REG0_REG_23__SCAN_IN), .ZN(n2828) );
  NAND2_X1 U35270 ( .A1(n3712), .A2(REG1_REG_23__SCAN_IN), .ZN(n2827) );
  NAND2_X1 U35280 ( .A1(n4018), .A2(n2890), .ZN(n2830) );
  INV_X1 U35290 ( .A(n4006), .ZN(n4002) );
  NAND2_X1 U35300 ( .A1(n4002), .A2(n2885), .ZN(n2829) );
  NAND2_X1 U35310 ( .A1(n2830), .A2(n2829), .ZN(n2831) );
  XNOR2_X1 U35320 ( .A(n2831), .B(n2888), .ZN(n2834) );
  NOR2_X1 U35330 ( .A1(n4006), .A2(n2873), .ZN(n2832) );
  AOI21_X1 U35340 ( .B1(n4018), .B2(n2891), .A(n2832), .ZN(n2833) );
  XNOR2_X1 U35350 ( .A(n2834), .B(n2833), .ZN(n3541) );
  NOR2_X1 U35360 ( .A1(n2834), .A2(n2833), .ZN(n2843) );
  OR2_X1 U35370 ( .A1(n2835), .A2(REG3_REG_24__SCAN_IN), .ZN(n2836) );
  NAND2_X1 U35380 ( .A1(n2844), .A2(n2836), .ZN(n3982) );
  AOI22_X1 U35390 ( .A1(n2492), .A2(REG2_REG_24__SCAN_IN), .B1(n2506), .B2(
        REG0_REG_24__SCAN_IN), .ZN(n2838) );
  NAND2_X1 U35400 ( .A1(n3712), .A2(REG1_REG_24__SCAN_IN), .ZN(n2837) );
  NAND2_X1 U35410 ( .A1(n3810), .A2(n2891), .ZN(n2840) );
  INV_X1 U35420 ( .A(n3980), .ZN(n3592) );
  NAND2_X1 U35430 ( .A1(n3592), .A2(n2890), .ZN(n2839) );
  NAND2_X1 U35440 ( .A1(n2840), .A2(n2839), .ZN(n2842) );
  OAI22_X1 U35450 ( .A1(n4005), .A2(n2873), .B1(n2872), .B2(n3980), .ZN(n2841)
         );
  XOR2_X1 U35460 ( .A(n2862), .B(n2841), .Z(n3587) );
  INV_X1 U35470 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3569) );
  NAND2_X1 U35480 ( .A1(n2844), .A2(n3569), .ZN(n2845) );
  NAND2_X1 U35490 ( .A1(n2854), .A2(n2845), .ZN(n3963) );
  INV_X1 U35500 ( .A(REG2_REG_25__SCAN_IN), .ZN(n3962) );
  NAND2_X1 U35510 ( .A1(n3712), .A2(REG1_REG_25__SCAN_IN), .ZN(n2847) );
  NAND2_X1 U35520 ( .A1(n2506), .A2(REG0_REG_25__SCAN_IN), .ZN(n2846) );
  OAI211_X1 U35530 ( .C1(n2539), .C2(n3962), .A(n2847), .B(n2846), .ZN(n2848)
         );
  INV_X1 U35540 ( .A(n2848), .ZN(n2849) );
  OAI22_X1 U35550 ( .A1(n3935), .A2(n2873), .B1(n2872), .B2(n3954), .ZN(n2851)
         );
  XNOR2_X1 U35560 ( .A(n2851), .B(n2862), .ZN(n2853) );
  OAI22_X1 U35570 ( .A1(n3935), .A2(n2875), .B1(n2873), .B2(n3954), .ZN(n2852)
         );
  OR2_X1 U35580 ( .A1(n2853), .A2(n2852), .ZN(n3565) );
  AND2_X1 U35590 ( .A1(n2853), .A2(n2852), .ZN(n3564) );
  INV_X1 U35600 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4810) );
  NAND2_X1 U35610 ( .A1(n2854), .A2(n4810), .ZN(n2855) );
  NAND2_X1 U35620 ( .A1(n3944), .A2(n2856), .ZN(n2861) );
  NAND2_X1 U35630 ( .A1(n3712), .A2(REG1_REG_26__SCAN_IN), .ZN(n2858) );
  NAND2_X1 U35640 ( .A1(n2506), .A2(REG0_REG_26__SCAN_IN), .ZN(n2857) );
  OAI211_X1 U35650 ( .C1(n2171), .C2(n4834), .A(n2858), .B(n2857), .ZN(n2859)
         );
  INV_X1 U35660 ( .A(n2859), .ZN(n2860) );
  OAI22_X1 U35670 ( .A1(n3790), .A2(n2873), .B1(n2872), .B2(n3942), .ZN(n2863)
         );
  XNOR2_X1 U35680 ( .A(n2863), .B(n2862), .ZN(n2865) );
  OAI22_X1 U35690 ( .A1(n3790), .A2(n2875), .B1(n2873), .B2(n3942), .ZN(n2864)
         );
  NAND2_X1 U35700 ( .A1(n2865), .A2(n2864), .ZN(n3628) );
  XNOR2_X1 U35710 ( .A(n2878), .B(REG3_REG_27__SCAN_IN), .ZN(n3927) );
  NAND2_X1 U35720 ( .A1(n3927), .A2(n2856), .ZN(n2871) );
  INV_X1 U35730 ( .A(REG2_REG_27__SCAN_IN), .ZN(n2868) );
  NAND2_X1 U35740 ( .A1(n3712), .A2(REG1_REG_27__SCAN_IN), .ZN(n2867) );
  NAND2_X1 U35750 ( .A1(n2506), .A2(REG0_REG_27__SCAN_IN), .ZN(n2866) );
  OAI211_X1 U35760 ( .C1(n2171), .C2(n2868), .A(n2867), .B(n2866), .ZN(n2869)
         );
  INV_X1 U35770 ( .A(n2869), .ZN(n2870) );
  OAI22_X1 U35780 ( .A1(n3523), .A2(n2873), .B1(n3926), .B2(n2872), .ZN(n2874)
         );
  XNOR2_X1 U35790 ( .A(n2874), .B(n2888), .ZN(n2920) );
  OAI22_X1 U35800 ( .A1(n3523), .A2(n2875), .B1(n3926), .B2(n2873), .ZN(n2918)
         );
  XNOR2_X1 U35810 ( .A(n2920), .B(n2918), .ZN(n3532) );
  INV_X1 U3582 ( .A(n2878), .ZN(n2876) );
  AOI21_X1 U3583 ( .B1(n2876), .B2(REG3_REG_27__SCAN_IN), .A(
        REG3_REG_28__SCAN_IN), .ZN(n2879) );
  NAND2_X1 U3584 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_28__SCAN_IN), .ZN(
        n2877) );
  NOR2_X1 U3585 ( .A1(n2878), .A2(n2877), .ZN(n3904) );
  INV_X1 U3586 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3518) );
  NAND2_X1 U3587 ( .A1(n3712), .A2(REG1_REG_28__SCAN_IN), .ZN(n2881) );
  NAND2_X1 U3588 ( .A1(n2506), .A2(REG0_REG_28__SCAN_IN), .ZN(n2880) );
  OAI211_X1 U3589 ( .C1(n2539), .C2(n3518), .A(n2881), .B(n2880), .ZN(n2882)
         );
  INV_X1 U3590 ( .A(n2882), .ZN(n2883) );
  NAND2_X1 U3591 ( .A1(n3913), .A2(n2890), .ZN(n2887) );
  NAND2_X1 U3592 ( .A1(n3716), .A2(DATAI_28_), .ZN(n3517) );
  INV_X1 U3593 ( .A(n3517), .ZN(n3521) );
  NAND2_X1 U3594 ( .A1(n3521), .A2(n2885), .ZN(n2886) );
  NAND2_X1 U3595 ( .A1(n2887), .A2(n2886), .ZN(n2889) );
  XNOR2_X1 U3596 ( .A(n2889), .B(n2888), .ZN(n2893) );
  AOI22_X1 U3597 ( .A1(n3913), .A2(n2891), .B1(n2890), .B2(n3521), .ZN(n2892)
         );
  XNOR2_X1 U3598 ( .A(n2893), .B(n2892), .ZN(n2926) );
  INV_X1 U3599 ( .A(n4315), .ZN(n2894) );
  NAND2_X1 U3600 ( .A1(n2894), .A2(n2897), .ZN(n2895) );
  MUX2_X1 U3601 ( .A(n2897), .B(n2895), .S(B_REG_SCAN_IN), .Z(n2896) );
  OAI22_X1 U3602 ( .A1(n3054), .A2(D_REG_1__SCAN_IN), .B1(n4315), .B2(n3058), 
        .ZN(n3039) );
  INV_X1 U3603 ( .A(n3039), .ZN(n3110) );
  INV_X1 U3604 ( .A(D_REG_0__SCAN_IN), .ZN(n3060) );
  INV_X1 U3605 ( .A(n3058), .ZN(n2898) );
  NOR4_X1 U3606 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_2__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n2908) );
  NOR4_X1 U3607 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2907) );
  INV_X1 U3608 ( .A(D_REG_8__SCAN_IN), .ZN(n4743) );
  INV_X1 U3609 ( .A(D_REG_24__SCAN_IN), .ZN(n4742) );
  INV_X1 U3610 ( .A(D_REG_9__SCAN_IN), .ZN(n4770) );
  INV_X1 U3611 ( .A(D_REG_12__SCAN_IN), .ZN(n4769) );
  NAND4_X1 U3612 ( .A1(n4743), .A2(n4742), .A3(n4770), .A4(n4769), .ZN(n2905)
         );
  NOR4_X1 U3613 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_7__SCAN_IN), .ZN(n2903) );
  NOR4_X1 U3614 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2902) );
  NOR4_X1 U3615 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2901) );
  NOR4_X1 U3616 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2900) );
  NAND4_X1 U3617 ( .A1(n2903), .A2(n2902), .A3(n2901), .A4(n2900), .ZN(n2904)
         );
  NOR4_X1 U3618 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(n2905), 
        .A4(n2904), .ZN(n2906) );
  NAND3_X1 U3619 ( .A1(n2908), .A2(n2907), .A3(n2906), .ZN(n2909) );
  NAND2_X1 U3620 ( .A1(n2910), .A2(n2909), .ZN(n3109) );
  NAND3_X1 U3621 ( .A1(n3110), .A2(n3111), .A3(n3109), .ZN(n2947) );
  OAI21_X1 U3622 ( .B1(n2913), .B2(n2912), .A(n2911), .ZN(n3066) );
  INV_X1 U3623 ( .A(n4510), .ZN(n2914) );
  INV_X1 U3624 ( .A(n3055), .ZN(n3064) );
  NAND2_X1 U3625 ( .A1(n2927), .A2(n3898), .ZN(n2938) );
  AOI21_X1 U3626 ( .B1(n4494), .B2(n2938), .A(n3065), .ZN(n2915) );
  AND2_X1 U3627 ( .A1(n2926), .A2(n4939), .ZN(n2916) );
  INV_X1 U3628 ( .A(n2926), .ZN(n2922) );
  INV_X1 U3629 ( .A(n2918), .ZN(n2919) );
  OR2_X1 U3630 ( .A1(n2920), .A2(n2919), .ZN(n2924) );
  AND2_X1 U3631 ( .A1(n2924), .A2(n4939), .ZN(n2921) );
  NAND2_X1 U3632 ( .A1(n2923), .A2(n2432), .ZN(n2954) );
  INV_X1 U3633 ( .A(n2924), .ZN(n2925) );
  NAND3_X1 U3634 ( .A1(n2926), .A2(n4939), .A3(n2925), .ZN(n2953) );
  INV_X1 U3635 ( .A(n2927), .ZN(n4319) );
  NAND2_X1 U3636 ( .A1(n2927), .A2(n4320), .ZN(n4502) );
  NOR2_X1 U3637 ( .A1(n4253), .A2(n4318), .ZN(n3038) );
  INV_X1 U3638 ( .A(n3624), .ZN(n3632) );
  NOR2_X1 U3639 ( .A1(n2929), .A2(n2768), .ZN(n2930) );
  MUX2_X1 U3640 ( .A(n2768), .B(n2930), .S(IR_REG_28__SCAN_IN), .Z(n2931) );
  INV_X1 U3641 ( .A(n2931), .ZN(n2933) );
  NAND2_X1 U3642 ( .A1(n2933), .A2(n2932), .ZN(n3163) );
  INV_X1 U3643 ( .A(n3163), .ZN(n4313) );
  NOR2_X1 U3644 ( .A1(n4510), .A2(n2934), .ZN(n2935) );
  NAND2_X1 U3645 ( .A1(n4313), .A2(n3803), .ZN(n2936) );
  OR2_X1 U3646 ( .A1(n2947), .A2(n2936), .ZN(n4926) );
  NAND2_X1 U3647 ( .A1(n4494), .A2(n4320), .ZN(n2937) );
  OAI21_X1 U3648 ( .B1(n4182), .B2(n2937), .A(n2947), .ZN(n3084) );
  NAND2_X1 U3649 ( .A1(n3065), .A2(n2938), .ZN(n3037) );
  NAND4_X1 U3650 ( .A1(n3084), .A2(n3066), .A3(n3052), .A4(n3037), .ZN(n2939)
         );
  NAND2_X1 U3651 ( .A1(n2939), .A2(STATE_REG_SCAN_IN), .ZN(n2940) );
  INV_X1 U3652 ( .A(n2940), .ZN(n4933) );
  OAI22_X1 U3653 ( .A1(n3523), .A2(n4926), .B1(n2940), .B2(n3519), .ZN(n2951)
         );
  NAND2_X1 U3654 ( .A1(n3904), .A2(n2856), .ZN(n2945) );
  NAND2_X1 U3655 ( .A1(n3712), .A2(REG1_REG_29__SCAN_IN), .ZN(n2942) );
  NAND2_X1 U3656 ( .A1(n2506), .A2(REG0_REG_29__SCAN_IN), .ZN(n2941) );
  OAI211_X1 U3657 ( .C1(n2539), .C2(n4811), .A(n2942), .B(n2941), .ZN(n2943)
         );
  INV_X1 U3658 ( .A(n2943), .ZN(n2944) );
  NAND2_X1 U3659 ( .A1(n2945), .A2(n2944), .ZN(n3809) );
  INV_X1 U3660 ( .A(n3809), .ZN(n2949) );
  NAND2_X1 U3661 ( .A1(n3803), .A2(n3163), .ZN(n2946) );
  INV_X1 U3662 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2948) );
  OAI22_X1 U3663 ( .A1(n2949), .A2(n3620), .B1(STATE_REG_SCAN_IN), .B2(n2948), 
        .ZN(n2950) );
  AOI211_X1 U3664 ( .C1(n3521), .C2(n3632), .A(n2951), .B(n2950), .ZN(n2952)
         );
  NAND4_X1 U3665 ( .A1(n2955), .A2(n2954), .A3(n2953), .A4(n2952), .ZN(U3217)
         );
  AND2_X1 U3666 ( .A1(n3824), .A2(n3135), .ZN(n3123) );
  NAND2_X1 U3667 ( .A1(n2957), .A2(n3136), .ZN(n2958) );
  NAND2_X1 U3668 ( .A1(n3125), .A2(n2958), .ZN(n3099) );
  NAND2_X1 U3669 ( .A1(n3822), .A2(n3156), .ZN(n3655) );
  NAND2_X1 U3670 ( .A1(n2959), .A2(n3117), .ZN(n3652) );
  NAND2_X1 U3671 ( .A1(n2959), .A2(n3156), .ZN(n2960) );
  NOR2_X1 U3672 ( .A1(n3821), .A2(n3007), .ZN(n2961) );
  INV_X1 U3673 ( .A(n3821), .ZN(n3155) );
  NAND2_X1 U3674 ( .A1(n3213), .A2(n3180), .ZN(n3658) );
  NAND2_X1 U3675 ( .A1(n3658), .A2(n3661), .ZN(n3776) );
  NAND2_X1 U3676 ( .A1(n3182), .A2(n3776), .ZN(n2963) );
  NAND2_X1 U3677 ( .A1(n4480), .A2(n3180), .ZN(n2962) );
  AND2_X1 U3678 ( .A1(n3820), .A2(n3215), .ZN(n2964) );
  INV_X1 U3679 ( .A(n3820), .ZN(n3250) );
  INV_X1 U3680 ( .A(n3215), .ZN(n3200) );
  NAND2_X1 U3681 ( .A1(n3250), .A2(n3200), .ZN(n2965) );
  NOR2_X1 U3682 ( .A1(n3819), .A2(n3248), .ZN(n3325) );
  NAND2_X1 U3683 ( .A1(n3818), .A2(n3320), .ZN(n2967) );
  INV_X1 U3684 ( .A(n2967), .ZN(n2966) );
  NAND2_X1 U3685 ( .A1(n3347), .A2(n3320), .ZN(n3011) );
  NAND2_X1 U3686 ( .A1(n3818), .A2(n3314), .ZN(n3674) );
  NAND2_X1 U3687 ( .A1(n3011), .A2(n3674), .ZN(n3784) );
  NOR2_X1 U3688 ( .A1(n2966), .A2(n3784), .ZN(n2969) );
  OR2_X1 U3689 ( .A1(n3325), .A2(n2969), .ZN(n2971) );
  NAND2_X1 U3690 ( .A1(n3819), .A2(n3248), .ZN(n3327) );
  AND2_X1 U3691 ( .A1(n3327), .A2(n2967), .ZN(n2968) );
  OR2_X1 U3692 ( .A1(n2969), .A2(n2968), .ZN(n2970) );
  AND2_X1 U3693 ( .A1(n3817), .A2(n3345), .ZN(n2972) );
  NOR2_X1 U3694 ( .A1(n3816), .A2(n3394), .ZN(n3370) );
  AND2_X1 U3695 ( .A1(n4461), .A2(n3382), .ZN(n2974) );
  NAND2_X1 U3696 ( .A1(n3816), .A2(n3394), .ZN(n3372) );
  AND2_X1 U3697 ( .A1(n2186), .A2(n3372), .ZN(n2973) );
  NOR2_X1 U3698 ( .A1(n2974), .A2(n2973), .ZN(n2975) );
  NAND2_X1 U3699 ( .A1(n3411), .A2(n3041), .ZN(n3424) );
  NAND2_X1 U3700 ( .A1(n3814), .A2(n4469), .ZN(n3687) );
  NAND2_X1 U3701 ( .A1(n3424), .A2(n3687), .ZN(n4459) );
  NOR2_X1 U3702 ( .A1(n3814), .A2(n3041), .ZN(n2976) );
  NAND2_X1 U3703 ( .A1(n4463), .A2(n3430), .ZN(n2977) );
  NAND2_X1 U3704 ( .A1(n2978), .A2(n2977), .ZN(n3463) );
  NAND2_X1 U3705 ( .A1(n4155), .A2(n3472), .ZN(n2979) );
  NAND2_X1 U3706 ( .A1(n3463), .A2(n2979), .ZN(n2981) );
  NAND2_X1 U3707 ( .A1(n3813), .A2(n3478), .ZN(n2980) );
  NAND2_X1 U3708 ( .A1(n2981), .A2(n2980), .ZN(n4157) );
  INV_X1 U3709 ( .A(n4157), .ZN(n2983) );
  NAND2_X1 U3710 ( .A1(n3473), .A2(n4164), .ZN(n3691) );
  NAND2_X1 U3711 ( .A1(n3812), .A2(n3498), .ZN(n3670) );
  AND2_X1 U3712 ( .A1(n4153), .A2(n3019), .ZN(n2984) );
  NOR2_X1 U3713 ( .A1(n3812), .A2(n4164), .ZN(n3503) );
  INV_X1 U3714 ( .A(n2984), .ZN(n2985) );
  INV_X1 U3715 ( .A(n4153), .ZN(n4139) );
  AOI22_X1 U3716 ( .A1(n3503), .A2(n2985), .B1(n4139), .B2(n3644), .ZN(n2986)
         );
  NAND2_X1 U3717 ( .A1(n4927), .A2(n4142), .ZN(n3727) );
  INV_X1 U3718 ( .A(n4927), .ZN(n3811) );
  NAND2_X1 U3719 ( .A1(n3811), .A2(n3580), .ZN(n3696) );
  OAI22_X2 U3720 ( .A1(n4134), .A2(n4136), .B1(n4927), .B2(n3580), .ZN(n4130)
         );
  NAND2_X1 U3721 ( .A1(n4104), .A2(n4936), .ZN(n2987) );
  NAND2_X1 U3722 ( .A1(n4130), .A2(n2987), .ZN(n2989) );
  NAND2_X1 U3723 ( .A1(n4137), .A2(n3042), .ZN(n2988) );
  NAND2_X1 U3724 ( .A1(n2989), .A2(n2988), .ZN(n4107) );
  INV_X1 U3725 ( .A(n4107), .ZN(n2991) );
  NAND2_X1 U3726 ( .A1(n4120), .A2(n4101), .ZN(n4080) );
  INV_X1 U3727 ( .A(n4120), .ZN(n4930) );
  NAND2_X1 U3728 ( .A1(n4930), .A2(n4112), .ZN(n4081) );
  NAND2_X1 U3729 ( .A1(n4120), .A2(n4112), .ZN(n2992) );
  NAND2_X1 U3730 ( .A1(n4102), .A2(n4091), .ZN(n2993) );
  NAND2_X1 U3731 ( .A1(n4041), .A2(n4071), .ZN(n3756) );
  NAND2_X1 U3732 ( .A1(n4056), .A2(n3756), .ZN(n2994) );
  INV_X1 U3733 ( .A(n4041), .ZN(n4086) );
  INV_X1 U3734 ( .A(n4071), .ZN(n4066) );
  NAND2_X1 U3735 ( .A1(n4086), .A2(n4066), .ZN(n3757) );
  NAND2_X1 U3736 ( .A1(n2994), .A2(n3757), .ZN(n4034) );
  NAND2_X1 U3737 ( .A1(n4063), .A2(n4039), .ZN(n2996) );
  NOR2_X1 U3738 ( .A1(n4063), .A2(n4039), .ZN(n2995) );
  AOI21_X1 U3739 ( .B1(n4034), .B2(n2996), .A(n2995), .ZN(n4024) );
  OR2_X1 U3740 ( .A1(n4040), .A2(n4026), .ZN(n3998) );
  NAND2_X1 U3741 ( .A1(n4040), .A2(n4026), .ZN(n3025) );
  NAND2_X1 U3742 ( .A1(n3998), .A2(n3025), .ZN(n4023) );
  INV_X1 U3743 ( .A(n4018), .ZN(n3974) );
  NOR2_X1 U3744 ( .A1(n4005), .A2(n3980), .ZN(n2998) );
  NOR2_X1 U3745 ( .A1(n3976), .A2(n3959), .ZN(n2999) );
  AOI21_X1 U3746 ( .B1(n3633), .B2(n3956), .A(n3932), .ZN(n3000) );
  OAI21_X1 U3747 ( .B1(n3920), .B2(n3937), .A(n3911), .ZN(n3002) );
  NAND2_X1 U3748 ( .A1(n3937), .A2(n3920), .ZN(n3001) );
  OR2_X1 U3749 ( .A1(n3913), .A2(n3517), .ZN(n3711) );
  NAND2_X1 U3750 ( .A1(n3913), .A2(n3517), .ZN(n3740) );
  NAND2_X1 U3751 ( .A1(n3711), .A2(n3740), .ZN(n3762) );
  NAND2_X1 U3752 ( .A1(n3716), .A2(DATAI_29_), .ZN(n3044) );
  OR2_X1 U3753 ( .A1(n3809), .A2(n3044), .ZN(n3718) );
  NAND2_X1 U3754 ( .A1(n3809), .A2(n3044), .ZN(n3741) );
  NAND2_X1 U3755 ( .A1(n3718), .A2(n3741), .ZN(n3767) );
  XNOR2_X1 U3756 ( .A(n3003), .B(n4317), .ZN(n3004) );
  NAND2_X1 U3757 ( .A1(n3004), .A2(n3898), .ZN(n4159) );
  NAND2_X1 U3758 ( .A1(n4159), .A2(n4253), .ZN(n4561) );
  INV_X1 U3759 ( .A(n3824), .ZN(n3093) );
  NAND2_X1 U3760 ( .A1(n3093), .A2(n3135), .ZN(n3782) );
  NAND2_X1 U3761 ( .A1(n3127), .A2(n3651), .ZN(n3101) );
  NAND2_X1 U3762 ( .A1(n3101), .A2(n3764), .ZN(n3006) );
  NAND2_X1 U3763 ( .A1(n3006), .A2(n3652), .ZN(n4475) );
  NAND2_X1 U3764 ( .A1(n3155), .A2(n3007), .ZN(n3657) );
  NAND2_X1 U3765 ( .A1(n3821), .A2(n4488), .ZN(n3654) );
  NAND2_X1 U3766 ( .A1(n4475), .A2(n4476), .ZN(n3008) );
  NAND2_X1 U3767 ( .A1(n3008), .A2(n3657), .ZN(n3184) );
  INV_X1 U3768 ( .A(n3658), .ZN(n3009) );
  AND2_X1 U3769 ( .A1(n3820), .A2(n3200), .ZN(n3194) );
  NAND2_X1 U3770 ( .A1(n3250), .A2(n3215), .ZN(n3675) );
  NAND2_X1 U3771 ( .A1(n3819), .A2(n3255), .ZN(n3677) );
  INV_X1 U3772 ( .A(n3819), .ZN(n3201) );
  NAND2_X1 U3773 ( .A1(n3201), .A2(n3248), .ZN(n3663) );
  NAND2_X1 U3774 ( .A1(n3010), .A2(n3663), .ZN(n3313) );
  INV_X1 U3775 ( .A(n3011), .ZN(n3012) );
  OR2_X1 U3776 ( .A1(n3313), .A2(n3012), .ZN(n3013) );
  NAND2_X1 U3777 ( .A1(n3013), .A2(n3674), .ZN(n3344) );
  INV_X1 U3778 ( .A(n3817), .ZN(n3315) );
  NAND2_X1 U3779 ( .A1(n3315), .A2(n3345), .ZN(n3667) );
  INV_X1 U3780 ( .A(n3345), .ZN(n3352) );
  NAND2_X1 U3781 ( .A1(n3817), .A2(n3352), .ZN(n3678) );
  INV_X1 U3782 ( .A(n3394), .ZN(n3361) );
  AND2_X1 U3783 ( .A1(n3816), .A2(n3361), .ZN(n3672) );
  INV_X1 U3784 ( .A(n3816), .ZN(n3014) );
  NAND2_X1 U3785 ( .A1(n3014), .A2(n3394), .ZN(n3668) );
  NAND2_X1 U3786 ( .A1(n3815), .A2(n3382), .ZN(n3686) );
  NAND2_X1 U3787 ( .A1(n3375), .A2(n3686), .ZN(n3015) );
  NAND2_X1 U3788 ( .A1(n4461), .A2(n3413), .ZN(n3681) );
  NAND2_X1 U3789 ( .A1(n4463), .A2(n3446), .ZN(n3468) );
  NAND2_X1 U3790 ( .A1(n3813), .A2(n3472), .ZN(n3464) );
  NAND2_X1 U3791 ( .A1(n3468), .A2(n3464), .ZN(n3017) );
  NAND2_X1 U3792 ( .A1(n3016), .A2(n3430), .ZN(n3467) );
  NAND2_X1 U3793 ( .A1(n3424), .A2(n3467), .ZN(n3018) );
  INV_X1 U3794 ( .A(n3017), .ZN(n3688) );
  NOR2_X1 U3795 ( .A1(n3813), .A2(n3472), .ZN(n3466) );
  AOI21_X1 U3796 ( .B1(n3018), .B2(n3688), .A(n3466), .ZN(n3689) );
  NAND2_X1 U3797 ( .A1(n4152), .A2(n4158), .ZN(n4151) );
  NAND2_X1 U3798 ( .A1(n4151), .A2(n3691), .ZN(n3505) );
  NAND2_X1 U3799 ( .A1(n4139), .A2(n3019), .ZN(n3690) );
  NAND2_X1 U3800 ( .A1(n4153), .A2(n3644), .ZN(n3671) );
  NAND2_X1 U3801 ( .A1(n3690), .A2(n3671), .ZN(n3779) );
  INV_X1 U3802 ( .A(n3696), .ZN(n3726) );
  NAND2_X1 U3803 ( .A1(n4102), .A2(n4085), .ZN(n3020) );
  NAND2_X1 U3804 ( .A1(n4081), .A2(n3020), .ZN(n3021) );
  INV_X1 U3805 ( .A(n3021), .ZN(n3992) );
  NOR2_X1 U3806 ( .A1(n4137), .A2(n4936), .ZN(n3989) );
  OAI22_X1 U3807 ( .A1(n3021), .A2(n4080), .B1(n4102), .B2(n4085), .ZN(n4057)
         );
  NOR2_X1 U3808 ( .A1(n4041), .A2(n4066), .ZN(n3022) );
  OR2_X1 U3809 ( .A1(n4057), .A2(n3022), .ZN(n3993) );
  AOI21_X1 U3810 ( .B1(n3992), .B2(n3989), .A(n3993), .ZN(n3023) );
  INV_X1 U3811 ( .A(n3023), .ZN(n3730) );
  NAND2_X1 U3812 ( .A1(n4137), .A2(n4936), .ZN(n3988) );
  NAND2_X1 U3813 ( .A1(n3992), .A2(n3988), .ZN(n3698) );
  AND2_X1 U3814 ( .A1(n4041), .A2(n4066), .ZN(n3701) );
  AOI21_X1 U3815 ( .B1(n3023), .B2(n3698), .A(n3701), .ZN(n3729) );
  INV_X1 U3816 ( .A(n3998), .ZN(n3024) );
  NOR2_X1 U3817 ( .A1(n4063), .A2(n4047), .ZN(n3794) );
  NOR2_X1 U3818 ( .A1(n3024), .A2(n3794), .ZN(n3735) );
  NAND2_X1 U3819 ( .A1(n4018), .A2(n4006), .ZN(n3755) );
  AND2_X1 U3820 ( .A1(n3755), .A2(n3025), .ZN(n3706) );
  AND2_X1 U3821 ( .A1(n4063), .A2(n4047), .ZN(n3700) );
  NAND2_X1 U3822 ( .A1(n3998), .A2(n3700), .ZN(n3026) );
  NAND2_X1 U3823 ( .A1(n3706), .A2(n3026), .ZN(n3733) );
  NAND2_X1 U3824 ( .A1(n3976), .A2(n3954), .ZN(n3759) );
  NAND2_X1 U3825 ( .A1(n3810), .A2(n3980), .ZN(n3950) );
  NAND2_X1 U3826 ( .A1(n3759), .A2(n3950), .ZN(n3732) );
  INV_X1 U3827 ( .A(n3732), .ZN(n3028) );
  OR2_X1 U3828 ( .A1(n3810), .A2(n3980), .ZN(n3754) );
  OR2_X1 U3829 ( .A1(n4018), .A2(n4006), .ZN(n3969) );
  AND2_X1 U3830 ( .A1(n3754), .A2(n3969), .ZN(n3704) );
  OR2_X1 U3831 ( .A1(n3732), .A2(n3704), .ZN(n3027) );
  NAND2_X1 U3832 ( .A1(n3935), .A2(n3959), .ZN(n3758) );
  NAND2_X1 U3833 ( .A1(n3027), .A2(n3758), .ZN(n3737) );
  AOI21_X1 U3834 ( .B1(n3971), .B2(n3028), .A(n3737), .ZN(n3934) );
  NAND2_X1 U3835 ( .A1(n3790), .A2(n3633), .ZN(n3723) );
  NAND2_X1 U3836 ( .A1(n3934), .A2(n3723), .ZN(n3917) );
  NAND2_X1 U3837 ( .A1(n3937), .A2(n3926), .ZN(n3709) );
  NAND2_X1 U3838 ( .A1(n3523), .A2(n3920), .ZN(n3710) );
  NAND2_X1 U3839 ( .A1(n3709), .A2(n3710), .ZN(n3912) );
  NAND2_X1 U3840 ( .A1(n3956), .A2(n3942), .ZN(n3916) );
  INV_X1 U3841 ( .A(n3916), .ZN(n3029) );
  NOR2_X1 U3842 ( .A1(n3912), .A2(n3029), .ZN(n3742) );
  NAND2_X1 U3843 ( .A1(n3917), .A2(n3742), .ZN(n3914) );
  INV_X1 U3844 ( .A(n3711), .ZN(n3030) );
  NAND2_X1 U3845 ( .A1(n4318), .A2(n4319), .ZN(n3032) );
  NAND2_X1 U3846 ( .A1(n4317), .A2(n4320), .ZN(n3031) );
  AOI222_X1 U3847 ( .A1(n3712), .A2(REG1_REG_30__SCAN_IN), .B1(n2492), .B2(
        REG2_REG_30__SCAN_IN), .C1(n2506), .C2(REG0_REG_30__SCAN_IN), .ZN(
        n3747) );
  NAND2_X1 U3848 ( .A1(n3163), .A2(n3065), .ZN(n4500) );
  XNOR2_X1 U3849 ( .A(n3033), .B(IR_REG_27__SCAN_IN), .ZN(n4314) );
  AND2_X1 U3850 ( .A1(n4314), .A2(B_REG_SCAN_IN), .ZN(n3034) );
  OR2_X1 U3851 ( .A1(n4500), .A2(n3034), .ZN(n4173) );
  OAI22_X1 U3852 ( .A1(n3747), .A2(n4173), .B1(n4477), .B2(n3044), .ZN(n3035)
         );
  AOI21_X1 U3853 ( .B1(n3913), .B2(n4088), .A(n3035), .ZN(n3036) );
  NAND2_X1 U3854 ( .A1(n3055), .A2(n3037), .ZN(n3108) );
  NOR2_X1 U3855 ( .A1(n3108), .A2(n3038), .ZN(n3040) );
  INV_X1 U3856 ( .A(n3516), .ZN(n3045) );
  INV_X1 U3857 ( .A(n3044), .ZN(n3043) );
  NAND2_X1 U3858 ( .A1(n3047), .A2(n3046), .ZN(U3547) );
  INV_X1 U3859 ( .A(REG0_REG_29__SCAN_IN), .ZN(n3050) );
  INV_X1 U3860 ( .A(n3111), .ZN(n3048) );
  INV_X2 U3861 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3862 ( .A(DATAI_26_), .ZN(n4699) );
  NAND2_X1 U3863 ( .A1(n3058), .A2(STATE_REG_SCAN_IN), .ZN(n3053) );
  OAI21_X1 U3864 ( .B1(STATE_REG_SCAN_IN), .B2(n4699), .A(n3053), .ZN(U3326)
         );
  INV_X1 U3865 ( .A(D_REG_1__SCAN_IN), .ZN(n3057) );
  NOR3_X1 U3866 ( .A1(n4315), .A2(n3058), .A3(n4510), .ZN(n3056) );
  AOI21_X1 U3867 ( .B1(n4508), .B2(n3057), .A(n3056), .ZN(U3459) );
  NOR3_X1 U3868 ( .A1(n3058), .A2(n4316), .A3(n4510), .ZN(n3059) );
  AOI21_X1 U3869 ( .B1(n4508), .B2(n3060), .A(n3059), .ZN(U3458) );
  INV_X1 U3870 ( .A(DATAI_29_), .ZN(n4840) );
  NAND2_X1 U3871 ( .A1(n3061), .A2(STATE_REG_SCAN_IN), .ZN(n3062) );
  OAI21_X1 U3872 ( .B1(STATE_REG_SCAN_IN), .B2(n4840), .A(n3062), .ZN(U3323)
         );
  INV_X1 U3873 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3063) );
  AND2_X1 U3874 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3838)
         );
  NAND2_X1 U3875 ( .A1(n4326), .A2(REG2_REG_1__SCAN_IN), .ZN(n3848) );
  MUX2_X1 U3876 ( .A(n2508), .B(REG2_REG_2__SCAN_IN), .S(n4325), .Z(n3847) );
  AOI21_X1 U3877 ( .B1(n3849), .B2(n3848), .A(n3847), .ZN(n3846) );
  XNOR2_X1 U3878 ( .A(n3168), .B(n4324), .ZN(n3170) );
  XNOR2_X1 U3879 ( .A(n3170), .B(REG2_REG_3__SCAN_IN), .ZN(n3079) );
  OR2_X1 U3880 ( .A1(n3066), .A2(U3149), .ZN(n3807) );
  NAND2_X1 U3881 ( .A1(n3064), .A2(n3807), .ZN(n3070) );
  NAND2_X1 U3882 ( .A1(n3066), .A2(n3065), .ZN(n3067) );
  AND2_X1 U3883 ( .A1(n3716), .A2(n3067), .ZN(n3068) );
  INV_X1 U3884 ( .A(n4314), .ZN(n3164) );
  NOR2_X1 U3885 ( .A1(n3163), .A2(n3164), .ZN(n3804) );
  INV_X1 U3886 ( .A(n3068), .ZN(n3069) );
  NOR2_X1 U3887 ( .A1(STATE_REG_SCAN_IN), .A2(n4486), .ZN(n3145) );
  INV_X1 U3888 ( .A(n4324), .ZN(n3075) );
  NOR2_X1 U3889 ( .A1(n4458), .A2(n3075), .ZN(n3071) );
  AOI211_X1 U3890 ( .C1(n4451), .C2(ADDR_REG_3__SCAN_IN), .A(n3145), .B(n3071), 
        .ZN(n3078) );
  XNOR2_X1 U3891 ( .A(n3072), .B(REG1_REG_1__SCAN_IN), .ZN(n3836) );
  AND2_X1 U3892 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3835)
         );
  NAND2_X1 U3893 ( .A1(n3836), .A2(n3835), .ZN(n3834) );
  NAND2_X1 U3894 ( .A1(n4326), .A2(REG1_REG_1__SCAN_IN), .ZN(n3073) );
  NAND2_X1 U3895 ( .A1(n3834), .A2(n3073), .ZN(n3853) );
  INV_X1 U3896 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4850) );
  MUX2_X1 U3897 ( .A(REG1_REG_2__SCAN_IN), .B(n4850), .S(n4325), .Z(n3854) );
  NAND2_X1 U3898 ( .A1(n3853), .A2(n3854), .ZN(n3852) );
  NAND2_X1 U3899 ( .A1(n4325), .A2(REG1_REG_2__SCAN_IN), .ZN(n3074) );
  NAND2_X1 U3900 ( .A1(n3852), .A2(n3074), .ZN(n3171) );
  XNOR2_X1 U3901 ( .A(n3171), .B(n3075), .ZN(n3076) );
  NAND2_X1 U3902 ( .A1(n3076), .A2(REG1_REG_3__SCAN_IN), .ZN(n3173) );
  OAI211_X1 U3903 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3076), .A(n4453), .B(n3173), 
        .ZN(n3077) );
  OAI211_X1 U3904 ( .C1(n3079), .C2(n4445), .A(n3078), .B(n3077), .ZN(U3243)
         );
  NOR2_X1 U3905 ( .A1(n4451), .A2(U4043), .ZN(U3148) );
  OAI21_X1 U3906 ( .B1(n3082), .B2(n3081), .A(n3080), .ZN(n3165) );
  INV_X1 U3907 ( .A(n3108), .ZN(n3083) );
  NAND2_X1 U3908 ( .A1(n3084), .A2(n3083), .ZN(n3159) );
  AOI22_X1 U3909 ( .A1(n2957), .A2(n4931), .B1(n3159), .B2(REG3_REG_0__SCAN_IN), .ZN(n3086) );
  OR2_X1 U3910 ( .A1(n3624), .A2(n4496), .ZN(n3085) );
  OAI211_X1 U3911 ( .C1(n3165), .C2(n3648), .A(n3086), .B(n3085), .ZN(U3229)
         );
  INV_X1 U3912 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4793) );
  NAND2_X1 U3913 ( .A1(n4137), .A2(U4043), .ZN(n3087) );
  OAI21_X1 U3914 ( .B1(U4043), .B2(n4793), .A(n3087), .ZN(U3567) );
  INV_X1 U3915 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4764) );
  INV_X1 U3916 ( .A(n3747), .ZN(n3088) );
  NAND2_X1 U3917 ( .A1(n3088), .A2(U4043), .ZN(n3089) );
  OAI21_X1 U3918 ( .B1(U4043), .B2(n4764), .A(n3089), .ZN(U3580) );
  CLKBUF_X1 U3919 ( .A(n3624), .Z(n4937) );
  OAI211_X1 U3920 ( .C1(n3092), .C2(n3091), .A(n3090), .B(n4939), .ZN(n3096)
         );
  OAI22_X1 U3921 ( .A1(n3093), .A2(n4926), .B1(n2959), .B2(n3620), .ZN(n3094)
         );
  AOI21_X1 U3922 ( .B1(REG3_REG_1__SCAN_IN), .B2(n3159), .A(n3094), .ZN(n3095)
         );
  OAI211_X1 U3923 ( .C1(n4937), .C2(n3097), .A(n3096), .B(n3095), .ZN(U3219)
         );
  NAND2_X1 U3924 ( .A1(n3099), .A2(n3764), .ZN(n3100) );
  NAND2_X1 U3925 ( .A1(n3098), .A2(n3100), .ZN(n4541) );
  NAND2_X1 U3926 ( .A1(n4541), .A2(n4498), .ZN(n3107) );
  XNOR2_X1 U3927 ( .A(n3101), .B(n3764), .ZN(n3102) );
  NAND2_X1 U3928 ( .A1(n3102), .A2(n4497), .ZN(n3106) );
  AOI22_X1 U3929 ( .A1(n3821), .A2(n4481), .B1(n3117), .B2(n4182), .ZN(n3103)
         );
  OAI21_X1 U3930 ( .B1(n4501), .B2(n4478), .A(n3103), .ZN(n3104) );
  INV_X1 U3931 ( .A(n3104), .ZN(n3105) );
  NAND3_X1 U3932 ( .A1(n3107), .A2(n3106), .A3(n3105), .ZN(n4539) );
  NAND3_X1 U3933 ( .A1(n3110), .A2(n3083), .A3(n3109), .ZN(n3112) );
  OR2_X1 U3934 ( .A1(n3112), .A2(n3111), .ZN(n3113) );
  MUX2_X1 U3935 ( .A(n4539), .B(REG2_REG_2__SCAN_IN), .S(n4507), .Z(n3114) );
  INV_X1 U3936 ( .A(n3114), .ZN(n3122) );
  NAND2_X1 U3937 ( .A1(n3115), .A2(n4320), .ZN(n3196) );
  INV_X1 U3938 ( .A(n3196), .ZN(n3116) );
  INV_X2 U3939 ( .A(n4507), .ZN(n4147) );
  NAND2_X1 U3940 ( .A1(n4147), .A2(n3898), .ZN(n4115) );
  INV_X1 U3941 ( .A(n4489), .ZN(n4538) );
  NAND2_X1 U3942 ( .A1(n3138), .A2(n3117), .ZN(n4537) );
  NAND2_X1 U3943 ( .A1(n4538), .A2(n4537), .ZN(n3119) );
  INV_X1 U3944 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3118) );
  OAI22_X1 U3945 ( .A1(n4096), .A2(n3119), .B1(n3118), .B2(n4166), .ZN(n3120)
         );
  AOI21_X1 U3946 ( .B1(n4541), .B2(n4504), .A(n3120), .ZN(n3121) );
  NAND2_X1 U3947 ( .A1(n3122), .A2(n3121), .ZN(U3288) );
  AND2_X1 U3948 ( .A1(n3125), .A2(n3124), .ZN(n4534) );
  INV_X1 U3949 ( .A(n4534), .ZN(n3142) );
  INV_X1 U3950 ( .A(n4504), .ZN(n3141) );
  NAND2_X1 U3951 ( .A1(n3127), .A2(n3126), .ZN(n3131) );
  NAND2_X1 U3952 ( .A1(n3136), .A2(n4182), .ZN(n3129) );
  NAND2_X1 U3953 ( .A1(n3824), .A2(n4088), .ZN(n3128) );
  OAI211_X1 U3954 ( .C1(n2959), .C2(n4500), .A(n3129), .B(n3128), .ZN(n3130)
         );
  AOI21_X1 U3955 ( .B1(n3131), .B2(n4497), .A(n3130), .ZN(n3133) );
  NAND2_X1 U3956 ( .A1(n4534), .A2(n4498), .ZN(n3132) );
  NAND2_X1 U3957 ( .A1(n3133), .A2(n3132), .ZN(n4533) );
  MUX2_X1 U3958 ( .A(n4533), .B(REG2_REG_1__SCAN_IN), .S(n4507), .Z(n3134) );
  INV_X1 U3959 ( .A(n3134), .ZN(n3140) );
  NAND2_X1 U3960 ( .A1(n3136), .A2(n3135), .ZN(n3137) );
  AND2_X1 U3961 ( .A1(n3138), .A2(n3137), .ZN(n4588) );
  AOI22_X1 U3962 ( .A1(n4491), .A2(n4588), .B1(REG3_REG_1__SCAN_IN), .B2(n4503), .ZN(n3139) );
  OAI211_X1 U3963 ( .C1(n3142), .C2(n3141), .A(n3140), .B(n3139), .ZN(U3289)
         );
  XOR2_X1 U3964 ( .A(n3144), .B(n3143), .Z(n3150) );
  AOI21_X1 U3965 ( .B1(n4480), .B2(n4931), .A(n3145), .ZN(n3147) );
  NAND2_X1 U3966 ( .A1(n3822), .A2(n3641), .ZN(n3146) );
  OAI211_X1 U3967 ( .C1(n4937), .C2(n4488), .A(n3147), .B(n3146), .ZN(n3148)
         );
  AOI21_X1 U3968 ( .B1(n4486), .B2(n4933), .A(n3148), .ZN(n3149) );
  OAI21_X1 U3969 ( .B1(n3150), .B2(n3648), .A(n3149), .ZN(U3215) );
  INV_X1 U3970 ( .A(n3151), .ZN(n3152) );
  AOI21_X1 U3971 ( .B1(n3154), .B2(n3153), .A(n3152), .ZN(n3161) );
  OAI22_X1 U3972 ( .A1(n3155), .A2(n3620), .B1(n4501), .B2(n4926), .ZN(n3158)
         );
  NOR2_X1 U3973 ( .A1(n4937), .A2(n3156), .ZN(n3157) );
  AOI211_X1 U3974 ( .C1(REG3_REG_2__SCAN_IN), .C2(n3159), .A(n3158), .B(n3157), 
        .ZN(n3160) );
  OAI21_X1 U3975 ( .B1(n3161), .B2(n3648), .A(n3160), .ZN(U3234) );
  AND2_X1 U3976 ( .A1(n4314), .A2(n2451), .ZN(n3162) );
  NOR2_X1 U3977 ( .A1(n3163), .A2(n3162), .ZN(n3828) );
  NAND3_X1 U3978 ( .A1(n3165), .A2(n4313), .A3(n3164), .ZN(n3167) );
  AOI21_X1 U3979 ( .B1(n3804), .B2(n3838), .A(n3823), .ZN(n3166) );
  OAI211_X1 U3980 ( .C1(IR_REG_0__SCAN_IN), .C2(n3828), .A(n3167), .B(n3166), 
        .ZN(n3858) );
  INV_X1 U3981 ( .A(n3168), .ZN(n3169) );
  XOR2_X1 U3982 ( .A(n3282), .B(REG2_REG_4__SCAN_IN), .Z(n3178) );
  INV_X1 U3983 ( .A(n4323), .ZN(n3283) );
  NAND2_X1 U3984 ( .A1(n3171), .A2(n4324), .ZN(n3172) );
  NAND2_X1 U3985 ( .A1(n3173), .A2(n3172), .ZN(n3266) );
  OAI211_X1 U3986 ( .C1(REG1_REG_4__SCAN_IN), .C2(n3174), .A(n4453), .B(n3265), 
        .ZN(n3176) );
  NOR2_X1 U3987 ( .A1(STATE_REG_SCAN_IN), .A2(n4728), .ZN(n3225) );
  AOI21_X1 U3988 ( .B1(n4451), .B2(ADDR_REG_4__SCAN_IN), .A(n3225), .ZN(n3175)
         );
  OAI211_X1 U3989 ( .C1(n4458), .C2(n3283), .A(n3176), .B(n3175), .ZN(n3177)
         );
  AOI21_X1 U3990 ( .B1(n4407), .B2(n3178), .A(n3177), .ZN(n3179) );
  NAND2_X1 U3991 ( .A1(n3858), .A2(n3179), .ZN(U3244) );
  AOI21_X1 U3992 ( .B1(n4487), .B2(n3180), .A(n4577), .ZN(n3181) );
  NAND2_X1 U3993 ( .A1(n3181), .A2(n3197), .ZN(n4549) );
  NOR2_X1 U3994 ( .A1(n4549), .A2(n4320), .ZN(n3191) );
  INV_X1 U3995 ( .A(n3776), .ZN(n3183) );
  XNOR2_X1 U3996 ( .A(n3182), .B(n3183), .ZN(n4548) );
  NAND2_X1 U3997 ( .A1(n4548), .A2(n4498), .ZN(n3190) );
  XNOR2_X1 U3998 ( .A(n3184), .B(n3183), .ZN(n3188) );
  NAND2_X1 U3999 ( .A1(n3821), .A2(n4088), .ZN(n3186) );
  NAND2_X1 U4000 ( .A1(n3820), .A2(n4481), .ZN(n3185) );
  OAI211_X1 U4001 ( .C1(n4477), .C2(n3228), .A(n3186), .B(n3185), .ZN(n3187)
         );
  AOI21_X1 U4002 ( .B1(n3188), .B2(n4497), .A(n3187), .ZN(n3189) );
  NAND2_X1 U4003 ( .A1(n3190), .A2(n3189), .ZN(n4552) );
  AOI211_X1 U4004 ( .C1(n4503), .C2(n3235), .A(n3191), .B(n4552), .ZN(n3193)
         );
  AOI22_X1 U4005 ( .A1(n4548), .A2(n4504), .B1(REG2_REG_4__SCAN_IN), .B2(n4507), .ZN(n3192) );
  OAI21_X1 U4006 ( .B1(n3193), .B2(n4507), .A(n3192), .ZN(U3286) );
  INV_X1 U4007 ( .A(n3194), .ZN(n3660) );
  NAND2_X1 U4008 ( .A1(n3660), .A2(n3675), .ZN(n3775) );
  XOR2_X1 U4009 ( .A(n3195), .B(n3775), .Z(n3220) );
  INV_X1 U4010 ( .A(n3220), .ZN(n3207) );
  AOI21_X1 U4011 ( .B1(n3215), .B2(n3197), .A(n3256), .ZN(n3222) );
  OAI22_X1 U4012 ( .A1(n3218), .A2(n4166), .B1(n2550), .B2(n4147), .ZN(n3198)
         );
  AOI21_X1 U4013 ( .B1(n3222), .B2(n4491), .A(n3198), .ZN(n3206) );
  XOR2_X1 U4014 ( .A(n3775), .B(n3199), .Z(n3204) );
  OAI22_X1 U4015 ( .A1(n3201), .A2(n4500), .B1(n4477), .B2(n3200), .ZN(n3202)
         );
  AOI21_X1 U4016 ( .B1(n4088), .B2(n4480), .A(n3202), .ZN(n3203) );
  OAI21_X1 U4017 ( .B1(n3204), .B2(n4483), .A(n3203), .ZN(n3219) );
  NAND2_X1 U4018 ( .A1(n3219), .A2(n4147), .ZN(n3205) );
  OAI211_X1 U4019 ( .C1(n3207), .C2(n4150), .A(n3206), .B(n3205), .ZN(U3285)
         );
  OAI211_X1 U4020 ( .C1(n3210), .C2(n3209), .A(n3208), .B(n4939), .ZN(n3217)
         );
  NAND2_X1 U4021 ( .A1(n4931), .A2(n3819), .ZN(n3212) );
  INV_X1 U4022 ( .A(REG3_REG_5__SCAN_IN), .ZN(n4683) );
  NOR2_X1 U4023 ( .A1(STATE_REG_SCAN_IN), .A2(n4683), .ZN(n4337) );
  INV_X1 U4024 ( .A(n4337), .ZN(n3211) );
  OAI211_X1 U4025 ( .C1(n3213), .C2(n4926), .A(n3212), .B(n3211), .ZN(n3214)
         );
  AOI21_X1 U4026 ( .B1(n3632), .B2(n3215), .A(n3214), .ZN(n3216) );
  OAI211_X1 U4027 ( .C1(n2940), .C2(n3218), .A(n3217), .B(n3216), .ZN(U3224)
         );
  AOI21_X1 U4028 ( .B1(n3220), .B2(n4561), .A(n3219), .ZN(n3224) );
  INV_X1 U4029 ( .A(n4247), .ZN(n4589) );
  AOI22_X1 U4030 ( .A1(n3222), .A2(n4589), .B1(REG1_REG_5__SCAN_IN), .B2(n4601), .ZN(n3221) );
  OAI21_X1 U4031 ( .B1(n3224), .B2(n4601), .A(n3221), .ZN(U3523) );
  INV_X1 U4032 ( .A(n4308), .ZN(n4535) );
  AOI22_X1 U4033 ( .A1(n3222), .A2(n4535), .B1(REG0_REG_5__SCAN_IN), .B2(n4584), .ZN(n3223) );
  OAI21_X1 U4034 ( .B1(n3224), .B2(n4584), .A(n3223), .ZN(U3477) );
  AOI21_X1 U4035 ( .B1(n4931), .B2(n3820), .A(n3225), .ZN(n3227) );
  NAND2_X1 U4036 ( .A1(n3641), .A2(n3821), .ZN(n3226) );
  OAI211_X1 U4037 ( .C1(n4937), .C2(n3228), .A(n3227), .B(n3226), .ZN(n3234)
         );
  INV_X1 U4038 ( .A(n3229), .ZN(n3230) );
  AOI211_X1 U4039 ( .C1(n3232), .C2(n3231), .A(n3648), .B(n3230), .ZN(n3233)
         );
  AOI211_X1 U4040 ( .C1(n3235), .C2(n4933), .A(n3234), .B(n3233), .ZN(n3236)
         );
  INV_X1 U4041 ( .A(n3236), .ZN(U3227) );
  XOR2_X1 U4042 ( .A(n3238), .B(n3237), .Z(n3239) );
  XNOR2_X1 U40430 ( .A(n3240), .B(n3239), .ZN(n3246) );
  NOR2_X1 U4044 ( .A1(STATE_REG_SCAN_IN), .A2(n3241), .ZN(n4347) );
  AOI21_X1 U4045 ( .B1(n3818), .B2(n4931), .A(n4347), .ZN(n3243) );
  NAND2_X1 U4046 ( .A1(n3641), .A2(n3820), .ZN(n3242) );
  OAI211_X1 U4047 ( .C1(n3624), .C2(n3255), .A(n3243), .B(n3242), .ZN(n3244)
         );
  AOI21_X1 U4048 ( .B1(n3257), .B2(n4933), .A(n3244), .ZN(n3245) );
  OAI21_X1 U4049 ( .B1(n3246), .B2(n3648), .A(n3245), .ZN(U3236) );
  NAND2_X1 U4050 ( .A1(n3663), .A2(n3677), .ZN(n3783) );
  XOR2_X1 U4051 ( .A(n3783), .B(n3326), .Z(n3254) );
  XOR2_X1 U4052 ( .A(n3783), .B(n3247), .Z(n3252) );
  AOI22_X1 U4053 ( .A1(n3818), .A2(n4481), .B1(n3248), .B2(n4182), .ZN(n3249)
         );
  OAI21_X1 U4054 ( .B1(n3250), .B2(n4478), .A(n3249), .ZN(n3251) );
  AOI21_X1 U4055 ( .B1(n3252), .B2(n4497), .A(n3251), .ZN(n3253) );
  OAI21_X1 U4056 ( .B1(n3254), .B2(n4159), .A(n3253), .ZN(n4555) );
  INV_X1 U4057 ( .A(n4555), .ZN(n3263) );
  INV_X1 U4058 ( .A(n3254), .ZN(n4557) );
  NOR2_X1 U4059 ( .A1(n3256), .A2(n3255), .ZN(n4554) );
  NOR3_X1 U4060 ( .A1(n4554), .A2(n4553), .A3(n4096), .ZN(n3261) );
  INV_X1 U4061 ( .A(n3257), .ZN(n3258) );
  OAI22_X1 U4062 ( .A1(n4147), .A2(n3259), .B1(n3258), .B2(n4166), .ZN(n3260)
         );
  AOI211_X1 U4063 ( .C1(n4557), .C2(n4504), .A(n3261), .B(n3260), .ZN(n3262)
         );
  OAI21_X1 U4064 ( .B1(n3263), .B2(n4507), .A(n3262), .ZN(U3284) );
  INV_X1 U4065 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4602) );
  AOI22_X1 U4066 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3278), .B1(n4518), .B2(
        n4602), .ZN(n4397) );
  NAND2_X1 U4067 ( .A1(n3279), .A2(REG1_REG_9__SCAN_IN), .ZN(n3271) );
  INV_X1 U4068 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3264) );
  INV_X1 U4069 ( .A(n3279), .ZN(n4521) );
  AOI22_X1 U4070 ( .A1(n3279), .A2(REG1_REG_9__SCAN_IN), .B1(n3264), .B2(n4521), .ZN(n4376) );
  INV_X1 U4071 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4849) );
  INV_X1 U4072 ( .A(n3281), .ZN(n4528) );
  AOI22_X1 U4073 ( .A1(n3281), .A2(n4849), .B1(REG1_REG_5__SCAN_IN), .B2(n4528), .ZN(n4334) );
  NOR2_X1 U4074 ( .A1(n4335), .A2(n4334), .ZN(n4333) );
  INV_X1 U4075 ( .A(n4525), .ZN(n4352) );
  INV_X1 U4076 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4868) );
  NOR2_X1 U4077 ( .A1(n4868), .A2(n4345), .ZN(n4344) );
  NOR2_X1 U4078 ( .A1(n3267), .A2(n4344), .ZN(n4357) );
  NAND2_X1 U4079 ( .A1(REG1_REG_7__SCAN_IN), .A2(n3280), .ZN(n4353) );
  INV_X1 U4080 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4596) );
  NAND2_X1 U4081 ( .A1(n4596), .A2(n4524), .ZN(n4354) );
  INV_X1 U4082 ( .A(n4354), .ZN(n3268) );
  AOI21_X1 U4083 ( .B1(n4357), .B2(n4353), .A(n3268), .ZN(n3269) );
  NAND2_X1 U4084 ( .A1(n3290), .A2(n3269), .ZN(n3270) );
  INV_X1 U4085 ( .A(n3290), .ZN(n4522) );
  XNOR2_X1 U4086 ( .A(n4522), .B(n3269), .ZN(n4366) );
  NAND2_X1 U4087 ( .A1(REG1_REG_8__SCAN_IN), .A2(n4366), .ZN(n4365) );
  NAND2_X1 U4088 ( .A1(n3270), .A2(n4365), .ZN(n4375) );
  NAND2_X1 U4089 ( .A1(n4376), .A2(n4375), .ZN(n4374) );
  NAND2_X1 U4090 ( .A1(n3271), .A2(n4374), .ZN(n3272) );
  NAND2_X1 U4091 ( .A1(n4519), .A2(n3272), .ZN(n3273) );
  INV_X1 U4092 ( .A(n4519), .ZN(n4391) );
  XNOR2_X1 U4093 ( .A(n3272), .B(n4391), .ZN(n4386) );
  NAND2_X1 U4094 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4386), .ZN(n4385) );
  NAND2_X1 U4095 ( .A1(n3297), .A2(n3274), .ZN(n3275) );
  NAND2_X1 U4096 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4413), .ZN(n4412) );
  XOR2_X1 U4097 ( .A(REG1_REG_13__SCAN_IN), .B(n3870), .Z(n3861) );
  XNOR2_X1 U4098 ( .A(n3859), .B(n3861), .ZN(n3304) );
  NOR2_X1 U4099 ( .A1(n3276), .A2(STATE_REG_SCAN_IN), .ZN(n3456) );
  AOI21_X1 U4100 ( .B1(n4451), .B2(ADDR_REG_13__SCAN_IN), .A(n3456), .ZN(n3277) );
  OAI21_X1 U4101 ( .B1(n4458), .B2(n3870), .A(n3277), .ZN(n3303) );
  NOR2_X1 U4102 ( .A1(n3870), .A2(n2686), .ZN(n3871) );
  AOI21_X1 U4103 ( .B1(n2686), .B2(n3870), .A(n3871), .ZN(n3301) );
  NAND2_X1 U4104 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3278), .ZN(n3296) );
  AOI22_X1 U4105 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3278), .B1(n4518), .B2(
        n2653), .ZN(n4400) );
  NAND2_X1 U4106 ( .A1(n3279), .A2(REG2_REG_9__SCAN_IN), .ZN(n3293) );
  AOI22_X1 U4107 ( .A1(n3279), .A2(REG2_REG_9__SCAN_IN), .B1(n2614), .B2(n4521), .ZN(n4379) );
  NAND2_X1 U4108 ( .A1(REG2_REG_7__SCAN_IN), .A2(n3280), .ZN(n3289) );
  AOI22_X1 U4109 ( .A1(REG2_REG_7__SCAN_IN), .A2(n3280), .B1(n4524), .B2(n2582), .ZN(n4362) );
  NAND2_X1 U4110 ( .A1(n3281), .A2(REG2_REG_5__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4111 ( .A1(n3281), .A2(REG2_REG_5__SCAN_IN), .B1(n2550), .B2(n4528), .ZN(n4340) );
  NAND2_X1 U4112 ( .A1(n4525), .A2(n3287), .ZN(n3288) );
  XNOR2_X1 U4113 ( .A(n3287), .B(n4352), .ZN(n4349) );
  NAND2_X1 U4114 ( .A1(REG2_REG_6__SCAN_IN), .A2(n4349), .ZN(n4348) );
  NAND2_X1 U4115 ( .A1(n3288), .A2(n4348), .ZN(n4361) );
  NAND2_X1 U4116 ( .A1(n4362), .A2(n4361), .ZN(n4360) );
  NAND2_X1 U4117 ( .A1(n3290), .A2(n3291), .ZN(n3292) );
  NAND2_X1 U4118 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4368), .ZN(n4367) );
  NAND2_X1 U4119 ( .A1(n3292), .A2(n4367), .ZN(n4378) );
  NAND2_X1 U4120 ( .A1(n4379), .A2(n4378), .ZN(n4377) );
  NAND2_X1 U4121 ( .A1(n4519), .A2(n3294), .ZN(n3295) );
  XNOR2_X1 U4122 ( .A(n3294), .B(n4391), .ZN(n4388) );
  NAND2_X1 U4123 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4388), .ZN(n4387) );
  NAND2_X1 U4124 ( .A1(n3295), .A2(n4387), .ZN(n4399) );
  NAND2_X1 U4125 ( .A1(n4400), .A2(n4399), .ZN(n4398) );
  NAND2_X1 U4126 ( .A1(n3297), .A2(n3298), .ZN(n3299) );
  OAI21_X1 U4127 ( .B1(n3301), .B2(n3872), .A(n4407), .ZN(n3300) );
  AOI21_X1 U4128 ( .B1(n3301), .B2(n3872), .A(n3300), .ZN(n3302) );
  AOI211_X1 U4129 ( .C1(n3304), .C2(n4453), .A(n3303), .B(n3302), .ZN(n3305)
         );
  INV_X1 U4130 ( .A(n3305), .ZN(U3253) );
  XNOR2_X1 U4131 ( .A(n3307), .B(n3306), .ZN(n3312) );
  INV_X1 U4132 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4684) );
  NOR2_X1 U4133 ( .A1(STATE_REG_SCAN_IN), .A2(n4684), .ZN(n4359) );
  AOI21_X1 U4134 ( .B1(n4931), .B2(n3817), .A(n4359), .ZN(n3309) );
  NAND2_X1 U4135 ( .A1(n3641), .A2(n3819), .ZN(n3308) );
  OAI211_X1 U4136 ( .C1(n3624), .C2(n3314), .A(n3309), .B(n3308), .ZN(n3310)
         );
  AOI21_X1 U4137 ( .B1(n3321), .B2(n4933), .A(n3310), .ZN(n3311) );
  OAI21_X1 U4138 ( .B1(n3312), .B2(n3648), .A(n3311), .ZN(U3210) );
  XNOR2_X1 U4139 ( .A(n3313), .B(n3784), .ZN(n3318) );
  OAI22_X1 U4140 ( .A1(n3315), .A2(n4500), .B1(n4477), .B2(n3314), .ZN(n3316)
         );
  AOI21_X1 U4141 ( .B1(n4088), .B2(n3819), .A(n3316), .ZN(n3317) );
  OAI21_X1 U4142 ( .B1(n3318), .B2(n4483), .A(n3317), .ZN(n4559) );
  INV_X1 U4143 ( .A(n4559), .ZN(n3332) );
  INV_X1 U4144 ( .A(n4553), .ZN(n3319) );
  AOI211_X1 U4145 ( .C1(n3320), .C2(n3319), .A(n4577), .B(n2201), .ZN(n4560)
         );
  INV_X1 U4146 ( .A(n4115), .ZN(n3324) );
  INV_X1 U4147 ( .A(n3321), .ZN(n3322) );
  OAI22_X1 U4148 ( .A1(n4147), .A2(n2582), .B1(n3322), .B2(n4166), .ZN(n3323)
         );
  AOI21_X1 U4149 ( .B1(n4560), .B2(n3324), .A(n3323), .ZN(n3331) );
  OR2_X1 U4150 ( .A1(n3326), .A2(n3325), .ZN(n3328) );
  NAND2_X1 U4151 ( .A1(n3328), .A2(n3327), .ZN(n3329) );
  XOR2_X1 U4152 ( .A(n3784), .B(n3329), .Z(n4562) );
  NAND2_X1 U4153 ( .A1(n4562), .A2(n4131), .ZN(n3330) );
  OAI211_X1 U4154 ( .C1(n3332), .C2(n4507), .A(n3331), .B(n3330), .ZN(U3283)
         );
  NOR2_X1 U4155 ( .A1(n2419), .A2(n3335), .ZN(n3336) );
  XNOR2_X1 U4156 ( .A(n3333), .B(n3336), .ZN(n3342) );
  NOR2_X1 U4157 ( .A1(STATE_REG_SCAN_IN), .A2(n3337), .ZN(n4372) );
  AOI21_X1 U4158 ( .B1(n4931), .B2(n3816), .A(n4372), .ZN(n3339) );
  NAND2_X1 U4159 ( .A1(n3818), .A2(n3641), .ZN(n3338) );
  OAI211_X1 U4160 ( .C1(n4937), .C2(n3352), .A(n3339), .B(n3338), .ZN(n3340)
         );
  AOI21_X1 U4161 ( .B1(n3353), .B2(n4933), .A(n3340), .ZN(n3341) );
  OAI21_X1 U4162 ( .B1(n3342), .B2(n3648), .A(n3341), .ZN(U3218) );
  NAND2_X1 U4163 ( .A1(n3667), .A2(n3678), .ZN(n3777) );
  XNOR2_X1 U4164 ( .A(n3343), .B(n3777), .ZN(n3351) );
  XNOR2_X1 U4165 ( .A(n3344), .B(n3777), .ZN(n3349) );
  AOI22_X1 U4166 ( .A1(n3816), .A2(n4481), .B1(n3345), .B2(n4182), .ZN(n3346)
         );
  OAI21_X1 U4167 ( .B1(n3347), .B2(n4478), .A(n3346), .ZN(n3348) );
  AOI21_X1 U4168 ( .B1(n3349), .B2(n4497), .A(n3348), .ZN(n3350) );
  OAI21_X1 U4169 ( .B1(n3351), .B2(n4159), .A(n3350), .ZN(n4566) );
  INV_X1 U4170 ( .A(n4566), .ZN(n3359) );
  INV_X1 U4171 ( .A(n3351), .ZN(n4568) );
  NOR2_X1 U4172 ( .A1(n2201), .A2(n3352), .ZN(n4565) );
  INV_X1 U4173 ( .A(n3365), .ZN(n4564) );
  NOR3_X1 U4174 ( .A1(n4565), .A2(n4564), .A3(n4096), .ZN(n3357) );
  INV_X1 U4175 ( .A(n3353), .ZN(n3354) );
  OAI22_X1 U4176 ( .A1(n4147), .A2(n3355), .B1(n3354), .B2(n4166), .ZN(n3356)
         );
  AOI211_X1 U4177 ( .C1(n4568), .C2(n4504), .A(n3357), .B(n3356), .ZN(n3358)
         );
  OAI21_X1 U4178 ( .B1(n3359), .B2(n4507), .A(n3358), .ZN(U3282) );
  INV_X1 U4179 ( .A(n3672), .ZN(n3679) );
  NAND2_X1 U4180 ( .A1(n3679), .A2(n3668), .ZN(n3778) );
  XNOR2_X1 U4181 ( .A(n3371), .B(n3778), .ZN(n3399) );
  INV_X1 U4182 ( .A(n3399), .ZN(n3369) );
  XOR2_X1 U4183 ( .A(n3778), .B(n3360), .Z(n3364) );
  OAI22_X1 U4184 ( .A1(n4461), .A2(n4500), .B1(n4477), .B2(n3361), .ZN(n3362)
         );
  AOI21_X1 U4185 ( .B1(n4088), .B2(n3817), .A(n3362), .ZN(n3363) );
  OAI21_X1 U4186 ( .B1(n3364), .B2(n4483), .A(n3363), .ZN(n3398) );
  NAND2_X1 U4187 ( .A1(n3398), .A2(n4147), .ZN(n3368) );
  AOI21_X1 U4188 ( .B1(n3394), .B2(n3365), .A(n3383), .ZN(n3401) );
  OAI22_X1 U4189 ( .A1(n3397), .A2(n4166), .B1(n2614), .B2(n4147), .ZN(n3366)
         );
  AOI21_X1 U4190 ( .B1(n3401), .B2(n4491), .A(n3366), .ZN(n3367) );
  OAI211_X1 U4191 ( .C1(n3369), .C2(n4150), .A(n3368), .B(n3367), .ZN(U3281)
         );
  OR2_X1 U4192 ( .A1(n3371), .A2(n3370), .ZN(n3373) );
  NAND2_X1 U4193 ( .A1(n3373), .A2(n3372), .ZN(n3374) );
  AND2_X1 U4194 ( .A1(n3681), .A2(n3686), .ZN(n3772) );
  XNOR2_X1 U4195 ( .A(n3374), .B(n3772), .ZN(n4574) );
  NAND2_X1 U4196 ( .A1(n4574), .A2(n4498), .ZN(n3381) );
  XNOR2_X1 U4197 ( .A(n3375), .B(n3772), .ZN(n3379) );
  NAND2_X1 U4198 ( .A1(n3413), .A2(n4182), .ZN(n3377) );
  NAND2_X1 U4199 ( .A1(n3816), .A2(n4088), .ZN(n3376) );
  OAI211_X1 U4200 ( .C1(n3411), .C2(n4500), .A(n3377), .B(n3376), .ZN(n3378)
         );
  AOI21_X1 U4201 ( .B1(n3379), .B2(n4497), .A(n3378), .ZN(n3380) );
  OR2_X1 U4202 ( .A1(n3383), .A2(n3382), .ZN(n4571) );
  AND3_X1 U4203 ( .A1(n4572), .A2(n4571), .A3(n4491), .ZN(n3386) );
  OAI22_X1 U4204 ( .A1(n4147), .A2(n3384), .B1(n3416), .B2(n4166), .ZN(n3385)
         );
  AOI211_X1 U4205 ( .C1(n4574), .C2(n4504), .A(n3386), .B(n3385), .ZN(n3387)
         );
  OAI21_X1 U4206 ( .B1(n4576), .B2(n4507), .A(n3387), .ZN(U3280) );
  OAI21_X1 U4207 ( .B1(n3389), .B2(n3388), .A(n3405), .ZN(n3390) );
  NAND2_X1 U4208 ( .A1(n3390), .A2(n4939), .ZN(n3396) );
  NAND2_X1 U4209 ( .A1(n3641), .A2(n3817), .ZN(n3392) );
  AND2_X1 U4210 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4383) );
  INV_X1 U4211 ( .A(n4383), .ZN(n3391) );
  OAI211_X1 U4212 ( .C1(n4461), .C2(n3620), .A(n3392), .B(n3391), .ZN(n3393)
         );
  AOI21_X1 U4213 ( .B1(n3632), .B2(n3394), .A(n3393), .ZN(n3395) );
  OAI211_X1 U4214 ( .C1(n2940), .C2(n3397), .A(n3396), .B(n3395), .ZN(U3228)
         );
  AOI21_X1 U4215 ( .B1(n4561), .B2(n3399), .A(n3398), .ZN(n3403) );
  AOI22_X1 U4216 ( .A1(n3401), .A2(n4535), .B1(REG0_REG_9__SCAN_IN), .B2(n4584), .ZN(n3400) );
  OAI21_X1 U4217 ( .B1(n3403), .B2(n4584), .A(n3400), .ZN(U3485) );
  AOI22_X1 U4218 ( .A1(n3401), .A2(n4589), .B1(REG1_REG_9__SCAN_IN), .B2(n4601), .ZN(n3402) );
  OAI21_X1 U4219 ( .B1(n3403), .B2(n4601), .A(n3402), .ZN(U3527) );
  AND2_X1 U4220 ( .A1(n3405), .A2(n3404), .ZN(n3408) );
  OAI211_X1 U4221 ( .C1(n3408), .C2(n3407), .A(n4939), .B(n3406), .ZN(n3415)
         );
  NAND2_X1 U4222 ( .A1(n3641), .A2(n3816), .ZN(n3410) );
  INV_X1 U4223 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4731) );
  NOR2_X1 U4224 ( .A1(STATE_REG_SCAN_IN), .A2(n4731), .ZN(n4393) );
  INV_X1 U4225 ( .A(n4393), .ZN(n3409) );
  OAI211_X1 U4226 ( .C1(n3411), .C2(n3620), .A(n3410), .B(n3409), .ZN(n3412)
         );
  AOI21_X1 U4227 ( .B1(n3632), .B2(n3413), .A(n3412), .ZN(n3414) );
  OAI211_X1 U4228 ( .C1(n2940), .C2(n3416), .A(n3415), .B(n3414), .ZN(U3214)
         );
  INV_X1 U4229 ( .A(n3438), .ZN(n3417) );
  NOR2_X1 U4230 ( .A1(n3417), .A2(n3436), .ZN(n3418) );
  XNOR2_X1 U4231 ( .A(n3437), .B(n3418), .ZN(n3423) );
  INV_X1 U4232 ( .A(REG3_REG_11__SCAN_IN), .ZN(n4701) );
  NOR2_X1 U4233 ( .A1(STATE_REG_SCAN_IN), .A2(n4701), .ZN(n4404) );
  AOI21_X1 U4234 ( .B1(n4463), .B2(n4931), .A(n4404), .ZN(n3420) );
  NAND2_X1 U4235 ( .A1(n3641), .A2(n3815), .ZN(n3419) );
  OAI211_X1 U4236 ( .C1(n3624), .C2(n4469), .A(n3420), .B(n3419), .ZN(n3421)
         );
  AOI21_X1 U4237 ( .B1(n4467), .B2(n4933), .A(n3421), .ZN(n3422) );
  OAI21_X1 U4238 ( .B1(n3423), .B2(n3648), .A(n3422), .ZN(U3233) );
  NAND2_X1 U4239 ( .A1(n3425), .A2(n3424), .ZN(n3470) );
  NAND2_X1 U4240 ( .A1(n3467), .A2(n3468), .ZN(n3771) );
  XNOR2_X1 U4241 ( .A(n3470), .B(n3771), .ZN(n3428) );
  OAI22_X1 U4242 ( .A1(n4155), .A2(n4500), .B1(n4477), .B2(n3446), .ZN(n3426)
         );
  AOI21_X1 U4243 ( .B1(n4088), .B2(n3814), .A(n3426), .ZN(n3427) );
  OAI21_X1 U4244 ( .B1(n3428), .B2(n4483), .A(n3427), .ZN(n3485) );
  INV_X1 U4245 ( .A(n3485), .ZN(n3435) );
  XOR2_X1 U4246 ( .A(n3771), .B(n3429), .Z(n3486) );
  NAND2_X1 U4247 ( .A1(n4468), .A2(n3430), .ZN(n3431) );
  NAND2_X1 U4248 ( .A1(n3479), .A2(n3431), .ZN(n3492) );
  AOI22_X1 U4249 ( .A1(n4507), .A2(REG2_REG_12__SCAN_IN), .B1(n3448), .B2(
        n4503), .ZN(n3432) );
  OAI21_X1 U4250 ( .B1(n3492), .B2(n4096), .A(n3432), .ZN(n3433) );
  AOI21_X1 U4251 ( .B1(n3486), .B2(n4131), .A(n3433), .ZN(n3434) );
  OAI21_X1 U4252 ( .B1(n4507), .B2(n3435), .A(n3434), .ZN(U3278) );
  OR2_X1 U4253 ( .A1(n3437), .A2(n3436), .ZN(n3439) );
  NAND2_X1 U4254 ( .A1(n3439), .A2(n3438), .ZN(n3443) );
  XNOR2_X1 U4255 ( .A(n3441), .B(n3440), .ZN(n3442) );
  XNOR2_X1 U4256 ( .A(n3443), .B(n3442), .ZN(n3450) );
  NAND2_X1 U4257 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4409) );
  OAI21_X1 U4258 ( .B1(n4155), .B2(n3620), .A(n4409), .ZN(n3444) );
  AOI21_X1 U4259 ( .B1(n3641), .B2(n3814), .A(n3444), .ZN(n3445) );
  OAI21_X1 U4260 ( .B1(n4937), .B2(n3446), .A(n3445), .ZN(n3447) );
  AOI21_X1 U4261 ( .B1(n3448), .B2(n4933), .A(n3447), .ZN(n3449) );
  OAI21_X1 U4262 ( .B1(n3450), .B2(n3648), .A(n3449), .ZN(U3221) );
  INV_X1 U4263 ( .A(n3451), .ZN(n3453) );
  NOR2_X1 U4264 ( .A1(n3453), .A2(n3452), .ZN(n3454) );
  XNOR2_X1 U4265 ( .A(n3455), .B(n3454), .ZN(n3462) );
  INV_X1 U4266 ( .A(n3456), .ZN(n3457) );
  OAI21_X1 U4267 ( .B1(n3473), .B2(n3620), .A(n3457), .ZN(n3458) );
  AOI21_X1 U4268 ( .B1(n3641), .B2(n4463), .A(n3458), .ZN(n3459) );
  OAI21_X1 U4269 ( .B1(n3624), .B2(n3472), .A(n3459), .ZN(n3460) );
  AOI21_X1 U4270 ( .B1(n3481), .B2(n4933), .A(n3460), .ZN(n3461) );
  OAI21_X1 U4271 ( .B1(n3462), .B2(n3648), .A(n3461), .ZN(U3231) );
  INV_X1 U4272 ( .A(n3464), .ZN(n3465) );
  NOR2_X1 U4273 ( .A1(n3466), .A2(n3465), .ZN(n3774) );
  XNOR2_X1 U4274 ( .A(n3463), .B(n3774), .ZN(n4254) );
  INV_X1 U4275 ( .A(n3467), .ZN(n3469) );
  OAI21_X1 U4276 ( .B1(n3470), .B2(n3469), .A(n3468), .ZN(n3471) );
  XNOR2_X1 U4277 ( .A(n3471), .B(n3774), .ZN(n3476) );
  OAI22_X1 U4278 ( .A1(n3473), .A2(n4500), .B1(n4477), .B2(n3472), .ZN(n3474)
         );
  AOI21_X1 U4279 ( .B1(n4088), .B2(n4463), .A(n3474), .ZN(n3475) );
  OAI21_X1 U4280 ( .B1(n3476), .B2(n4483), .A(n3475), .ZN(n3477) );
  AOI21_X1 U4281 ( .B1(n4498), .B2(n4254), .A(n3477), .ZN(n4256) );
  NAND2_X1 U4282 ( .A1(n3479), .A2(n3478), .ZN(n3480) );
  NAND2_X1 U4283 ( .A1(n2199), .A2(n3480), .ZN(n4257) );
  AOI22_X1 U4284 ( .A1(n4507), .A2(REG2_REG_13__SCAN_IN), .B1(n3481), .B2(
        n4503), .ZN(n3482) );
  OAI21_X1 U4285 ( .B1(n4257), .B2(n4096), .A(n3482), .ZN(n3483) );
  AOI21_X1 U4286 ( .B1(n4254), .B2(n4504), .A(n3483), .ZN(n3484) );
  OAI21_X1 U4287 ( .B1(n4256), .B2(n4507), .A(n3484), .ZN(U3277) );
  INV_X1 U4288 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3487) );
  AOI21_X1 U4289 ( .B1(n3486), .B2(n4561), .A(n3485), .ZN(n3489) );
  MUX2_X1 U4290 ( .A(n3487), .B(n3489), .S(n4604), .Z(n3488) );
  OAI21_X1 U4291 ( .B1(n3492), .B2(n4247), .A(n3488), .ZN(U3530) );
  INV_X1 U4292 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3490) );
  MUX2_X1 U4293 ( .A(n3490), .B(n3489), .S(n4585), .Z(n3491) );
  OAI21_X1 U4294 ( .B1(n3492), .B2(n4308), .A(n3491), .ZN(U3491) );
  XNOR2_X1 U4295 ( .A(n2190), .B(n3493), .ZN(n3494) );
  XNOR2_X1 U4296 ( .A(n3495), .B(n3494), .ZN(n3501) );
  NAND2_X1 U4297 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4416) );
  OAI21_X1 U4298 ( .B1(n4139), .B2(n3620), .A(n4416), .ZN(n3496) );
  AOI21_X1 U4299 ( .B1(n3641), .B2(n3813), .A(n3496), .ZN(n3497) );
  OAI21_X1 U4300 ( .B1(n4937), .B2(n3498), .A(n3497), .ZN(n3499) );
  AOI21_X1 U4301 ( .B1(n4165), .B2(n4933), .A(n3499), .ZN(n3500) );
  OAI21_X1 U4302 ( .B1(n3501), .B2(n3648), .A(n3500), .ZN(U3212) );
  INV_X1 U4303 ( .A(n3502), .ZN(n4156) );
  NOR2_X1 U4304 ( .A1(n4156), .A2(n3503), .ZN(n3504) );
  XOR2_X1 U4305 ( .A(n3779), .B(n3504), .Z(n4245) );
  INV_X1 U4306 ( .A(n4245), .ZN(n3514) );
  XNOR2_X1 U4307 ( .A(n3505), .B(n3779), .ZN(n3508) );
  OAI22_X1 U4308 ( .A1(n4927), .A2(n4500), .B1(n4477), .B2(n3644), .ZN(n3506)
         );
  AOI21_X1 U4309 ( .B1(n4088), .B2(n3812), .A(n3506), .ZN(n3507) );
  OAI21_X1 U4310 ( .B1(n3508), .B2(n4483), .A(n3507), .ZN(n4244) );
  OAI21_X1 U4311 ( .B1(n4163), .B2(n3644), .A(n2200), .ZN(n4309) );
  NOR2_X1 U4312 ( .A1(n4309), .A2(n4096), .ZN(n3512) );
  OAI22_X1 U4313 ( .A1(n4147), .A2(n3510), .B1(n3509), .B2(n4166), .ZN(n3511)
         );
  AOI211_X1 U4314 ( .C1(n4244), .C2(n4147), .A(n3512), .B(n3511), .ZN(n3513)
         );
  OAI21_X1 U4315 ( .B1(n3514), .B2(n4150), .A(n3513), .ZN(U3275) );
  XNOR2_X1 U4316 ( .A(n3515), .B(n3762), .ZN(n4189) );
  OAI21_X1 U4317 ( .B1(n3924), .B2(n3517), .A(n3516), .ZN(n4266) );
  INV_X1 U4318 ( .A(n4266), .ZN(n3528) );
  OAI22_X1 U4319 ( .A1(n3519), .A2(n4166), .B1(n3518), .B2(n4147), .ZN(n3527)
         );
  XOR2_X1 U4320 ( .A(n3762), .B(n3520), .Z(n3525) );
  AOI22_X1 U4321 ( .A1(n3809), .A2(n4481), .B1(n4182), .B2(n3521), .ZN(n3522)
         );
  OAI21_X1 U4322 ( .B1(n3523), .B2(n4478), .A(n3522), .ZN(n3524) );
  AOI21_X1 U4323 ( .B1(n3525), .B2(n4497), .A(n3524), .ZN(n4188) );
  NOR2_X1 U4324 ( .A1(n4188), .A2(n4507), .ZN(n3526) );
  AOI211_X1 U4325 ( .C1(n4491), .C2(n3528), .A(n3527), .B(n3526), .ZN(n3529)
         );
  OAI21_X1 U4326 ( .B1(n4189), .B2(n4150), .A(n3529), .ZN(U3262) );
  NAND3_X1 U4327 ( .A1(n2446), .A2(STATE_REG_SCAN_IN), .A3(IR_REG_31__SCAN_IN), 
        .ZN(n3531) );
  INV_X1 U4328 ( .A(DATAI_31_), .ZN(n3530) );
  OAI22_X1 U4329 ( .A1(n2449), .A2(n3531), .B1(STATE_REG_SCAN_IN), .B2(n3530), 
        .ZN(U3321) );
  XNOR2_X1 U4330 ( .A(n3533), .B(n3532), .ZN(n3540) );
  INV_X1 U4331 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3534) );
  OAI22_X1 U4332 ( .A1(n3790), .A2(n4926), .B1(STATE_REG_SCAN_IN), .B2(n3534), 
        .ZN(n3535) );
  AOI21_X1 U4333 ( .B1(n3913), .B2(n4931), .A(n3535), .ZN(n3537) );
  NAND2_X1 U4334 ( .A1(n3927), .A2(n4933), .ZN(n3536) );
  OAI211_X1 U4335 ( .C1(n4937), .C2(n3926), .A(n3537), .B(n3536), .ZN(n3538)
         );
  INV_X1 U4336 ( .A(n3538), .ZN(n3539) );
  OAI21_X1 U4337 ( .B1(n3540), .B2(n3648), .A(n3539), .ZN(U3211) );
  OAI21_X1 U4338 ( .B1(n3606), .B2(n3542), .A(n3541), .ZN(n3543) );
  NAND3_X1 U4339 ( .A1(n2182), .A2(n4939), .A3(n3543), .ZN(n3547) );
  NOR2_X1 U4340 ( .A1(n4937), .A2(n4006), .ZN(n3545) );
  INV_X1 U4341 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4808) );
  OAI22_X1 U4342 ( .A1(n4005), .A2(n3620), .B1(STATE_REG_SCAN_IN), .B2(n4808), 
        .ZN(n3544) );
  AOI211_X1 U4343 ( .C1(n3641), .C2(n4040), .A(n3545), .B(n3544), .ZN(n3546)
         );
  OAI211_X1 U4344 ( .C1(n2940), .C2(n4009), .A(n3547), .B(n3546), .ZN(U3213)
         );
  XOR2_X1 U4345 ( .A(n3549), .B(n3548), .Z(n3554) );
  NAND2_X1 U4346 ( .A1(n4931), .A2(n4041), .ZN(n3550) );
  NAND2_X1 U4347 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3897) );
  OAI211_X1 U4348 ( .C1(n4120), .C2(n4926), .A(n3550), .B(n3897), .ZN(n3552)
         );
  NOR2_X1 U4349 ( .A1(n4937), .A2(n4085), .ZN(n3551) );
  AOI211_X1 U4350 ( .C1(n4094), .C2(n4933), .A(n3552), .B(n3551), .ZN(n3553)
         );
  OAI21_X1 U4351 ( .B1(n3554), .B2(n3648), .A(n3553), .ZN(U3216) );
  XNOR2_X1 U4352 ( .A(n3556), .B(n3555), .ZN(n3557) );
  XNOR2_X1 U4353 ( .A(n3558), .B(n3557), .ZN(n3563) );
  AOI22_X1 U4354 ( .A1(n4040), .A2(n4931), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3560) );
  NAND2_X1 U4355 ( .A1(n3641), .A2(n4041), .ZN(n3559) );
  OAI211_X1 U4356 ( .C1(n3624), .C2(n4047), .A(n3560), .B(n3559), .ZN(n3561)
         );
  AOI21_X1 U4357 ( .B1(n4049), .B2(n4933), .A(n3561), .ZN(n3562) );
  OAI21_X1 U4358 ( .B1(n3563), .B2(n3648), .A(n3562), .ZN(U3220) );
  NAND2_X1 U4359 ( .A1(n2222), .A2(n3565), .ZN(n3566) );
  XNOR2_X1 U4360 ( .A(n3567), .B(n3566), .ZN(n3568) );
  NAND2_X1 U4361 ( .A1(n3568), .A2(n4939), .ZN(n3573) );
  NOR2_X1 U4362 ( .A1(n4005), .A2(n4926), .ZN(n3571) );
  OAI22_X1 U4363 ( .A1(n3790), .A2(n3620), .B1(STATE_REG_SCAN_IN), .B2(n3569), 
        .ZN(n3570) );
  AOI211_X1 U4364 ( .C1(n3959), .C2(n3632), .A(n3571), .B(n3570), .ZN(n3572)
         );
  OAI211_X1 U4365 ( .C1(n2940), .C2(n3963), .A(n3573), .B(n3572), .ZN(U3222)
         );
  INV_X1 U4366 ( .A(n3637), .ZN(n3574) );
  OAI21_X1 U4367 ( .B1(n3574), .B2(n3640), .A(n3638), .ZN(n3575) );
  XOR2_X1 U4368 ( .A(n3576), .B(n3575), .Z(n3583) );
  INV_X1 U4369 ( .A(REG3_REG_16__SCAN_IN), .ZN(n3577) );
  NOR2_X1 U4370 ( .A1(STATE_REG_SCAN_IN), .A2(n3577), .ZN(n4439) );
  AOI21_X1 U4371 ( .B1(n4137), .B2(n4931), .A(n4439), .ZN(n3579) );
  NAND2_X1 U4372 ( .A1(n3641), .A2(n4153), .ZN(n3578) );
  OAI211_X1 U4373 ( .C1(n3624), .C2(n3580), .A(n3579), .B(n3578), .ZN(n3581)
         );
  AOI21_X1 U4374 ( .B1(n4143), .B2(n4933), .A(n3581), .ZN(n3582) );
  OAI21_X1 U4375 ( .B1(n3583), .B2(n3648), .A(n3582), .ZN(U3223) );
  INV_X1 U4376 ( .A(n3584), .ZN(n3585) );
  NOR2_X1 U4377 ( .A1(n3586), .A2(n3585), .ZN(n3588) );
  XNOR2_X1 U4378 ( .A(n3588), .B(n3587), .ZN(n3589) );
  NAND2_X1 U4379 ( .A1(n3589), .A2(n4939), .ZN(n3594) );
  NOR2_X1 U4380 ( .A1(n3974), .A2(n4926), .ZN(n3591) );
  INV_X1 U4381 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4807) );
  OAI22_X1 U4382 ( .A1(n3935), .A2(n3620), .B1(STATE_REG_SCAN_IN), .B2(n4807), 
        .ZN(n3590) );
  AOI211_X1 U4383 ( .C1(n3592), .C2(n3632), .A(n3591), .B(n3590), .ZN(n3593)
         );
  OAI211_X1 U4384 ( .C1(n2940), .C2(n3982), .A(n3594), .B(n3593), .ZN(U3226)
         );
  INV_X1 U4385 ( .A(n3595), .ZN(n3600) );
  AOI21_X1 U4386 ( .B1(n3599), .B2(n3597), .A(n3596), .ZN(n3598) );
  AOI21_X1 U4387 ( .B1(n3600), .B2(n3599), .A(n3598), .ZN(n3605) );
  AOI22_X1 U4388 ( .A1(n4931), .A2(n4063), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n3602) );
  NAND2_X1 U4389 ( .A1(n3641), .A2(n4102), .ZN(n3601) );
  OAI211_X1 U4390 ( .C1(n3624), .C2(n4066), .A(n3602), .B(n3601), .ZN(n3603)
         );
  AOI21_X1 U4391 ( .B1(n4072), .B2(n4933), .A(n3603), .ZN(n3604) );
  OAI21_X1 U4392 ( .B1(n3605), .B2(n3648), .A(n3604), .ZN(U3230) );
  AOI21_X1 U4393 ( .B1(n3608), .B2(n3607), .A(n3606), .ZN(n3614) );
  INV_X1 U4394 ( .A(n4029), .ZN(n3612) );
  AOI22_X1 U4395 ( .A1(n4018), .A2(n4931), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n3610) );
  NAND2_X1 U4396 ( .A1(n3641), .A2(n4063), .ZN(n3609) );
  OAI211_X1 U4397 ( .C1(n4937), .C2(n4026), .A(n3610), .B(n3609), .ZN(n3611)
         );
  AOI21_X1 U4398 ( .B1(n3612), .B2(n4933), .A(n3611), .ZN(n3613) );
  OAI21_X1 U4399 ( .B1(n3614), .B2(n3648), .A(n3613), .ZN(U3232) );
  INV_X1 U4400 ( .A(n3615), .ZN(n3617) );
  NAND2_X1 U4401 ( .A1(n3617), .A2(n3616), .ZN(n3618) );
  XNOR2_X1 U4402 ( .A(n3619), .B(n3618), .ZN(n3627) );
  NAND2_X1 U4403 ( .A1(REG3_REG_18__SCAN_IN), .A2(U3149), .ZN(n4444) );
  OAI21_X1 U4404 ( .B1(n3621), .B2(n3620), .A(n4444), .ZN(n3622) );
  AOI21_X1 U4405 ( .B1(n3641), .B2(n4137), .A(n3622), .ZN(n3623) );
  OAI21_X1 U4406 ( .B1(n3624), .B2(n4112), .A(n3623), .ZN(n3625) );
  AOI21_X1 U4407 ( .B1(n4113), .B2(n4933), .A(n3625), .ZN(n3626) );
  OAI21_X1 U4408 ( .B1(n3627), .B2(n3648), .A(n3626), .ZN(U3235) );
  NAND2_X1 U4409 ( .A1(n2193), .A2(n3628), .ZN(n3629) );
  XNOR2_X1 U4410 ( .A(n3630), .B(n3629), .ZN(n3636) );
  OAI22_X1 U4411 ( .A1(n3935), .A2(n4926), .B1(STATE_REG_SCAN_IN), .B2(n4810), 
        .ZN(n3631) );
  AOI21_X1 U4412 ( .B1(n3633), .B2(n3632), .A(n3631), .ZN(n3635) );
  AOI22_X1 U4413 ( .A1(n3937), .A2(n4931), .B1(n3944), .B2(n4933), .ZN(n3634)
         );
  OAI211_X1 U4414 ( .C1(n3636), .C2(n3648), .A(n3635), .B(n3634), .ZN(U3237)
         );
  NAND2_X1 U4415 ( .A1(n3638), .A2(n3637), .ZN(n3639) );
  XOR2_X1 U4416 ( .A(n3640), .B(n3639), .Z(n3649) );
  AND2_X1 U4417 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4429) );
  AOI21_X1 U4418 ( .B1(n3811), .B2(n4931), .A(n4429), .ZN(n3643) );
  NAND2_X1 U4419 ( .A1(n3812), .A2(n3641), .ZN(n3642) );
  OAI211_X1 U4420 ( .C1(n4937), .C2(n3644), .A(n3643), .B(n3642), .ZN(n3645)
         );
  AOI21_X1 U4421 ( .B1(n3646), .B2(n4933), .A(n3645), .ZN(n3647) );
  OAI21_X1 U4422 ( .B1(n3649), .B2(n3648), .A(n3647), .ZN(U3238) );
  AND2_X1 U4423 ( .A1(n3741), .A2(n3740), .ZN(n3719) );
  NAND2_X1 U4424 ( .A1(n3824), .A2(n4496), .ZN(n3781) );
  OAI211_X1 U4425 ( .C1(n2336), .C2(n4318), .A(n3781), .B(n3650), .ZN(n3653)
         );
  NAND3_X1 U4426 ( .A1(n3653), .A2(n3652), .A3(n3651), .ZN(n3656) );
  NAND3_X1 U4427 ( .A1(n3656), .A2(n3655), .A3(n3654), .ZN(n3659) );
  NAND3_X1 U4428 ( .A1(n3659), .A2(n3658), .A3(n3657), .ZN(n3662) );
  NAND4_X1 U4429 ( .A1(n3662), .A2(n3661), .A3(n3677), .A4(n3660), .ZN(n3665)
         );
  INV_X1 U4430 ( .A(n3784), .ZN(n3664) );
  NAND3_X1 U4431 ( .A1(n3665), .A2(n3664), .A3(n3663), .ZN(n3666) );
  NAND3_X1 U4432 ( .A1(n3666), .A2(n3674), .A3(n3678), .ZN(n3669) );
  NAND3_X1 U4433 ( .A1(n3669), .A2(n3668), .A3(n3667), .ZN(n3685) );
  NAND2_X1 U4434 ( .A1(n3671), .A2(n3670), .ZN(n3673) );
  NOR2_X1 U4435 ( .A1(n3673), .A2(n3672), .ZN(n3684) );
  NAND2_X1 U4436 ( .A1(n3673), .A2(n3690), .ZN(n3724) );
  INV_X1 U4437 ( .A(n3674), .ZN(n3676) );
  NOR2_X1 U4438 ( .A1(n3676), .A2(n3675), .ZN(n3680) );
  NAND4_X1 U4439 ( .A1(n3680), .A2(n3679), .A3(n3678), .A4(n3677), .ZN(n3682)
         );
  NAND2_X1 U4440 ( .A1(n3682), .A2(n3681), .ZN(n3683) );
  AOI22_X1 U4441 ( .A1(n3685), .A2(n3684), .B1(n3724), .B2(n3683), .ZN(n3695)
         );
  NAND3_X1 U4442 ( .A1(n3688), .A2(n3687), .A3(n3686), .ZN(n3694) );
  INV_X1 U4443 ( .A(n3689), .ZN(n3692) );
  NAND2_X1 U4444 ( .A1(n3691), .A2(n3690), .ZN(n3725) );
  OAI21_X1 U4445 ( .B1(n3692), .B2(n3725), .A(n3724), .ZN(n3693) );
  OAI21_X1 U4446 ( .B1(n3695), .B2(n3694), .A(n3693), .ZN(n3697) );
  NAND2_X1 U4447 ( .A1(n3697), .A2(n3696), .ZN(n3699) );
  AOI21_X1 U4448 ( .B1(n3699), .B2(n3727), .A(n3698), .ZN(n3702) );
  INV_X1 U4449 ( .A(n3700), .ZN(n3795) );
  INV_X1 U4450 ( .A(n3701), .ZN(n3995) );
  OAI211_X1 U4451 ( .C1(n3702), .C2(n3730), .A(n3795), .B(n3995), .ZN(n3703)
         );
  NAND2_X1 U4452 ( .A1(n3735), .A2(n3703), .ZN(n3705) );
  INV_X1 U4453 ( .A(n3704), .ZN(n3951) );
  AOI21_X1 U4454 ( .B1(n3706), .B2(n3705), .A(n3951), .ZN(n3707) );
  OAI211_X1 U4455 ( .C1(n3707), .C2(n3732), .A(n3723), .B(n3758), .ZN(n3708)
         );
  NAND4_X1 U4456 ( .A1(n3719), .A2(n3709), .A3(n3916), .A4(n3708), .ZN(n3721)
         );
  NAND2_X1 U4457 ( .A1(n3711), .A2(n3710), .ZN(n3722) );
  AND2_X1 U4458 ( .A1(n3716), .A2(DATAI_30_), .ZN(n4183) );
  INV_X1 U4459 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3715) );
  NAND2_X1 U4460 ( .A1(n3712), .A2(REG1_REG_31__SCAN_IN), .ZN(n3714) );
  NAND2_X1 U4461 ( .A1(n2506), .A2(REG0_REG_31__SCAN_IN), .ZN(n3713) );
  OAI211_X1 U4462 ( .C1(n2171), .C2(n3715), .A(n3714), .B(n3713), .ZN(n4175)
         );
  NAND2_X1 U4463 ( .A1(n3716), .A2(DATAI_31_), .ZN(n4176) );
  NAND2_X1 U4464 ( .A1(n4175), .A2(n4176), .ZN(n3720) );
  INV_X1 U4465 ( .A(n3720), .ZN(n3717) );
  AOI21_X1 U4466 ( .B1(n3747), .B2(n4183), .A(n3717), .ZN(n3793) );
  NAND2_X1 U4467 ( .A1(n3793), .A2(n3718), .ZN(n3736) );
  AOI21_X1 U4468 ( .B1(n3719), .B2(n3722), .A(n3736), .ZN(n3744) );
  OR2_X1 U4469 ( .A1(n4175), .A2(n4176), .ZN(n3748) );
  OAI21_X1 U4470 ( .B1(n3747), .B2(n4183), .A(n3748), .ZN(n3760) );
  AOI22_X1 U4471 ( .A1(n3721), .A2(n3744), .B1(n3760), .B2(n3720), .ZN(n3801)
         );
  INV_X1 U4472 ( .A(n4183), .ZN(n3753) );
  INV_X1 U4473 ( .A(n3722), .ZN(n3746) );
  INV_X1 U4474 ( .A(n3723), .ZN(n3739) );
  OAI21_X1 U4475 ( .B1(n4152), .B2(n3725), .A(n3724), .ZN(n3728) );
  AOI21_X1 U4476 ( .B1(n3728), .B2(n3727), .A(n3726), .ZN(n3731) );
  OAI21_X1 U4477 ( .B1(n3731), .B2(n3730), .A(n3729), .ZN(n3734) );
  AOI211_X1 U4478 ( .C1(n3735), .C2(n3734), .A(n3733), .B(n3732), .ZN(n3738)
         );
  NOR4_X1 U4479 ( .A1(n3739), .A2(n3738), .A3(n3737), .A4(n3736), .ZN(n3745)
         );
  NAND3_X1 U4480 ( .A1(n3742), .A2(n3741), .A3(n3740), .ZN(n3743) );
  AOI22_X1 U4481 ( .A1(n3746), .A2(n3745), .B1(n3744), .B2(n3743), .ZN(n3750)
         );
  OAI21_X1 U4482 ( .B1(n3747), .B2(n4176), .A(n3750), .ZN(n3752) );
  INV_X1 U4483 ( .A(n4175), .ZN(n3749) );
  OAI211_X1 U4484 ( .C1(n3750), .C2(n3749), .A(n4318), .B(n3748), .ZN(n3751)
         );
  AOI21_X1 U4485 ( .B1(n3753), .B2(n3752), .A(n3751), .ZN(n3799) );
  AND2_X1 U4486 ( .A1(n3754), .A2(n3950), .ZN(n3972) );
  AND2_X1 U4487 ( .A1(n3969), .A2(n3755), .ZN(n3999) );
  AND2_X1 U4488 ( .A1(n3757), .A2(n3756), .ZN(n4060) );
  NAND2_X1 U4489 ( .A1(n3759), .A2(n3758), .ZN(n3953) );
  XNOR2_X1 U4490 ( .A(n4102), .B(n4085), .ZN(n4084) );
  NOR4_X1 U4491 ( .A1(n4060), .A2(n3953), .A3(n4084), .A4(n3760), .ZN(n3761)
         );
  NAND3_X1 U4492 ( .A1(n3972), .A2(n3999), .A3(n3761), .ZN(n3797) );
  INV_X1 U4493 ( .A(n3762), .ZN(n3769) );
  INV_X1 U4494 ( .A(n3912), .ZN(n3915) );
  NAND4_X1 U4495 ( .A1(n3765), .A2(n4158), .A3(n3764), .A4(n3763), .ZN(n3766)
         );
  NOR2_X1 U4496 ( .A1(n3767), .A2(n3766), .ZN(n3768) );
  AND3_X1 U4497 ( .A1(n3769), .A2(n3915), .A3(n3768), .ZN(n3792) );
  INV_X1 U4498 ( .A(n3988), .ZN(n3770) );
  NOR2_X1 U4499 ( .A1(n3989), .A2(n3770), .ZN(n4129) );
  INV_X1 U4500 ( .A(n3771), .ZN(n3773) );
  AND4_X1 U4501 ( .A1(n4129), .A2(n3774), .A3(n3773), .A4(n3772), .ZN(n3789)
         );
  NOR4_X1 U4502 ( .A1(n2990), .A2(n4459), .A3(n3776), .A4(n3775), .ZN(n3788)
         );
  INV_X1 U4503 ( .A(n4476), .ZN(n3780) );
  NOR4_X1 U4504 ( .A1(n3780), .A2(n3779), .A3(n3778), .A4(n3777), .ZN(n3787)
         );
  INV_X1 U4505 ( .A(n4136), .ZN(n3785) );
  NAND2_X1 U4506 ( .A1(n3782), .A2(n3781), .ZN(n4531) );
  NOR4_X1 U4507 ( .A1(n3785), .A2(n3784), .A3(n3783), .A4(n4531), .ZN(n3786)
         );
  AND4_X1 U4508 ( .A1(n3789), .A2(n3788), .A3(n3787), .A4(n3786), .ZN(n3791)
         );
  XNOR2_X1 U4509 ( .A(n3790), .B(n3942), .ZN(n3933) );
  NAND4_X1 U4510 ( .A1(n3793), .A2(n3792), .A3(n3791), .A4(n3933), .ZN(n3796)
         );
  INV_X1 U4511 ( .A(n3794), .ZN(n3997) );
  NAND2_X1 U4512 ( .A1(n3997), .A2(n3795), .ZN(n4037) );
  NOR4_X1 U4513 ( .A1(n3797), .A2(n3796), .A3(n4037), .A4(n4023), .ZN(n3798)
         );
  OR2_X1 U4514 ( .A1(n3799), .A2(n3798), .ZN(n3800) );
  MUX2_X1 U4515 ( .A(n3801), .B(n3800), .S(n4319), .Z(n3802) );
  XNOR2_X1 U4516 ( .A(n3802), .B(n4320), .ZN(n3808) );
  NAND2_X1 U4517 ( .A1(n3804), .A2(n3803), .ZN(n3805) );
  OAI211_X1 U4518 ( .C1(n4317), .C2(n3807), .A(n3805), .B(B_REG_SCAN_IN), .ZN(
        n3806) );
  OAI21_X1 U4519 ( .B1(n3808), .B2(n3807), .A(n3806), .ZN(U3239) );
  MUX2_X1 U4520 ( .A(n4175), .B(DATAO_REG_31__SCAN_IN), .S(n3823), .Z(U3581)
         );
  MUX2_X1 U4521 ( .A(n3809), .B(DATAO_REG_29__SCAN_IN), .S(n3823), .Z(U3579)
         );
  MUX2_X1 U4522 ( .A(DATAO_REG_28__SCAN_IN), .B(n3913), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4523 ( .A(n3937), .B(DATAO_REG_27__SCAN_IN), .S(n3823), .Z(U3577)
         );
  MUX2_X1 U4524 ( .A(n3956), .B(DATAO_REG_26__SCAN_IN), .S(n3823), .Z(U3576)
         );
  MUX2_X1 U4525 ( .A(n3976), .B(DATAO_REG_25__SCAN_IN), .S(n3823), .Z(U3575)
         );
  MUX2_X1 U4526 ( .A(DATAO_REG_24__SCAN_IN), .B(n3810), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4527 ( .A(n4018), .B(DATAO_REG_23__SCAN_IN), .S(n3823), .Z(U3573)
         );
  MUX2_X1 U4528 ( .A(DATAO_REG_22__SCAN_IN), .B(n4040), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4529 ( .A(n4063), .B(DATAO_REG_21__SCAN_IN), .S(n3823), .Z(U3571)
         );
  MUX2_X1 U4530 ( .A(n4041), .B(DATAO_REG_20__SCAN_IN), .S(n3823), .Z(U3570)
         );
  MUX2_X1 U4531 ( .A(n4102), .B(DATAO_REG_19__SCAN_IN), .S(n3823), .Z(U3569)
         );
  MUX2_X1 U4532 ( .A(DATAO_REG_18__SCAN_IN), .B(n4930), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4533 ( .A(DATAO_REG_16__SCAN_IN), .B(n3811), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4534 ( .A(n4153), .B(DATAO_REG_15__SCAN_IN), .S(n3823), .Z(U3565)
         );
  MUX2_X1 U4535 ( .A(DATAO_REG_14__SCAN_IN), .B(n3812), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4536 ( .A(DATAO_REG_13__SCAN_IN), .B(n3813), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4537 ( .A(DATAO_REG_12__SCAN_IN), .B(n4463), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4538 ( .A(DATAO_REG_11__SCAN_IN), .B(n3814), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4539 ( .A(n3815), .B(DATAO_REG_10__SCAN_IN), .S(n3823), .Z(U3560)
         );
  MUX2_X1 U4540 ( .A(n3816), .B(DATAO_REG_9__SCAN_IN), .S(n3823), .Z(U3559) );
  MUX2_X1 U4541 ( .A(n3817), .B(DATAO_REG_8__SCAN_IN), .S(n3823), .Z(U3558) );
  MUX2_X1 U4542 ( .A(DATAO_REG_7__SCAN_IN), .B(n3818), .S(U4043), .Z(U3557) );
  MUX2_X1 U4543 ( .A(n3819), .B(DATAO_REG_6__SCAN_IN), .S(n3823), .Z(U3556) );
  MUX2_X1 U4544 ( .A(n3820), .B(DATAO_REG_5__SCAN_IN), .S(n3823), .Z(U3555) );
  MUX2_X1 U4545 ( .A(DATAO_REG_4__SCAN_IN), .B(n4480), .S(U4043), .Z(U3554) );
  MUX2_X1 U4546 ( .A(n3821), .B(DATAO_REG_3__SCAN_IN), .S(n3823), .Z(U3553) );
  MUX2_X1 U4547 ( .A(DATAO_REG_2__SCAN_IN), .B(n3822), .S(U4043), .Z(U3552) );
  MUX2_X1 U4548 ( .A(DATAO_REG_1__SCAN_IN), .B(n2956), .S(U4043), .Z(U3551) );
  MUX2_X1 U4549 ( .A(n3824), .B(DATAO_REG_0__SCAN_IN), .S(n3823), .Z(U3550) );
  INV_X1 U4550 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4586) );
  NAND3_X1 U4551 ( .A1(n4453), .A2(IR_REG_0__SCAN_IN), .A3(n4586), .ZN(n3832)
         );
  NAND2_X1 U4552 ( .A1(n4451), .A2(ADDR_REG_0__SCAN_IN), .ZN(n3831) );
  NAND2_X1 U4553 ( .A1(U3149), .A2(REG3_REG_0__SCAN_IN), .ZN(n3830) );
  NOR2_X1 U4554 ( .A1(n4314), .A2(REG1_REG_0__SCAN_IN), .ZN(n3825) );
  OAI21_X1 U4555 ( .B1(IR_REG_0__SCAN_IN), .B2(n3825), .A(n3828), .ZN(n3827)
         );
  OAI211_X1 U4556 ( .C1(IR_REG_0__SCAN_IN), .C2(n3828), .A(n3827), .B(n3826), 
        .ZN(n3829) );
  NAND4_X1 U4557 ( .A1(n3832), .A2(n3831), .A3(n3830), .A4(n3829), .ZN(U3240)
         );
  INV_X1 U4558 ( .A(n4458), .ZN(n3833) );
  NAND2_X1 U4559 ( .A1(n3833), .A2(n4326), .ZN(n3842) );
  OAI211_X1 U4560 ( .C1(n3836), .C2(n3835), .A(n4453), .B(n3834), .ZN(n3841)
         );
  OAI211_X1 U4561 ( .C1(n3838), .C2(n3837), .A(n4407), .B(n3849), .ZN(n3840)
         );
  AOI22_X1 U4562 ( .A1(n4451), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3839) );
  NAND4_X1 U4563 ( .A1(n3842), .A2(n3841), .A3(n3840), .A4(n3839), .ZN(U3241)
         );
  INV_X1 U4564 ( .A(n4325), .ZN(n3844) );
  AOI22_X1 U4565 ( .A1(n4451), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3843) );
  OAI21_X1 U4566 ( .B1(n4458), .B2(n3844), .A(n3843), .ZN(n3845) );
  INV_X1 U4567 ( .A(n3845), .ZN(n3857) );
  INV_X1 U4568 ( .A(n3846), .ZN(n3851) );
  NAND3_X1 U4569 ( .A1(n3849), .A2(n3848), .A3(n3847), .ZN(n3850) );
  NAND3_X1 U4570 ( .A1(n4407), .A2(n3851), .A3(n3850), .ZN(n3856) );
  OAI211_X1 U4571 ( .C1(n3854), .C2(n3853), .A(n4453), .B(n3852), .ZN(n3855)
         );
  NAND4_X1 U4572 ( .A1(n3858), .A2(n3857), .A3(n3856), .A4(n3855), .ZN(U3242)
         );
  INV_X1 U4573 ( .A(n3877), .ZN(n4516) );
  INV_X1 U4574 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4852) );
  AOI22_X1 U4575 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3877), .B1(n4516), .B2(
        n4852), .ZN(n4432) );
  INV_X1 U4576 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3860) );
  NAND2_X1 U4577 ( .A1(n3874), .A2(n3862), .ZN(n3863) );
  NAND2_X1 U4578 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4422), .ZN(n4421) );
  NAND2_X1 U4579 ( .A1(n3863), .A2(n4421), .ZN(n4431) );
  NAND2_X1 U4580 ( .A1(n4432), .A2(n4431), .ZN(n4430) );
  NOR2_X1 U4581 ( .A1(n3878), .A2(n3864), .ZN(n3865) );
  INV_X1 U4582 ( .A(n3878), .ZN(n4515) );
  INV_X1 U4583 ( .A(REG1_REG_17__SCAN_IN), .ZN(n3867) );
  INV_X1 U4584 ( .A(n3884), .ZN(n4321) );
  NOR2_X1 U4585 ( .A1(n4321), .A2(REG1_REG_17__SCAN_IN), .ZN(n3890) );
  INV_X1 U4586 ( .A(n3890), .ZN(n3866) );
  OAI21_X1 U4587 ( .B1(n3867), .B2(n3884), .A(n3866), .ZN(n3868) );
  NOR2_X1 U4588 ( .A1(n3869), .A2(n3868), .ZN(n3889) );
  AOI21_X1 U4589 ( .B1(n3869), .B2(n3868), .A(n3889), .ZN(n3888) );
  INV_X1 U4590 ( .A(n4453), .ZN(n4343) );
  XNOR2_X1 U4591 ( .A(n3884), .B(REG2_REG_17__SCAN_IN), .ZN(n3882) );
  INV_X1 U4592 ( .A(n3870), .ZN(n4322) );
  NOR2_X1 U4593 ( .A1(n2208), .A2(n3873), .ZN(n3875) );
  NOR2_X1 U4594 ( .A1(n4168), .A2(n4418), .ZN(n4417) );
  NAND2_X1 U4595 ( .A1(REG2_REG_15__SCAN_IN), .A2(n3877), .ZN(n3876) );
  OAI21_X1 U4596 ( .B1(REG2_REG_15__SCAN_IN), .B2(n3877), .A(n3876), .ZN(n4426) );
  NOR2_X1 U4597 ( .A1(n4427), .A2(n4426), .ZN(n4425) );
  NAND2_X1 U4598 ( .A1(n3879), .A2(n4515), .ZN(n3880) );
  INV_X1 U4599 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4435) );
  NAND2_X1 U4600 ( .A1(n3881), .A2(n3882), .ZN(n3893) );
  AOI221_X1 U4601 ( .B1(n3882), .B2(n3893), .C1(n3881), .C2(n3893), .A(n4445), 
        .ZN(n3886) );
  NOR2_X1 U4602 ( .A1(STATE_REG_SCAN_IN), .A2(n2739), .ZN(n4929) );
  AOI21_X1 U4603 ( .B1(n4451), .B2(ADDR_REG_17__SCAN_IN), .A(n4929), .ZN(n3883) );
  OAI21_X1 U4604 ( .B1(n4458), .B2(n3884), .A(n3883), .ZN(n3885) );
  NOR2_X1 U4605 ( .A1(n3886), .A2(n3885), .ZN(n3887) );
  OAI21_X1 U4606 ( .B1(n3888), .B2(n4343), .A(n3887), .ZN(U3257) );
  INV_X1 U4607 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4790) );
  MUX2_X1 U4608 ( .A(REG1_REG_19__SCAN_IN), .B(n4790), .S(n3898), .Z(n3892) );
  INV_X1 U4609 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3891) );
  INV_X1 U4610 ( .A(n3894), .ZN(n4513) );
  AOI22_X1 U4611 ( .A1(REG1_REG_18__SCAN_IN), .A2(n3894), .B1(n4513), .B2(
        n3891), .ZN(n4455) );
  AOI22_X1 U4612 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4513), .B1(n3894), .B2(
        n2763), .ZN(n4448) );
  MUX2_X1 U4613 ( .A(n2773), .B(REG2_REG_19__SCAN_IN), .S(n3898), .Z(n3895) );
  NAND2_X1 U4614 ( .A1(n4451), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3896) );
  OAI211_X1 U4615 ( .C1(n4458), .C2(n3898), .A(n3897), .B(n3896), .ZN(n3899)
         );
  AOI21_X1 U4616 ( .B1(n3900), .B2(n4407), .A(n3899), .ZN(n3901) );
  OAI21_X1 U4617 ( .B1(n3902), .B2(n4343), .A(n3901), .ZN(U3259) );
  NAND2_X1 U4618 ( .A1(n3903), .A2(n4131), .ZN(n3910) );
  INV_X1 U4619 ( .A(n3904), .ZN(n3905) );
  OAI22_X1 U4620 ( .A1(n3906), .A2(n4096), .B1(n4166), .B2(n3905), .ZN(n3907)
         );
  OAI21_X1 U4621 ( .B1(n3908), .B2(n3907), .A(n4147), .ZN(n3909) );
  OAI211_X1 U4622 ( .C1(n4147), .C2(n4811), .A(n3910), .B(n3909), .ZN(U3354)
         );
  XOR2_X1 U4623 ( .A(n3912), .B(n3911), .Z(n4193) );
  INV_X1 U4624 ( .A(n4193), .ZN(n3931) );
  INV_X1 U4625 ( .A(n3913), .ZN(n3923) );
  INV_X1 U4626 ( .A(n3914), .ZN(n3919) );
  AOI21_X1 U4627 ( .B1(n3917), .B2(n3916), .A(n3915), .ZN(n3918) );
  OAI21_X1 U4628 ( .B1(n3919), .B2(n3918), .A(n4497), .ZN(n3922) );
  AOI22_X1 U4629 ( .A1(n3956), .A2(n4088), .B1(n3920), .B2(n4182), .ZN(n3921)
         );
  OAI211_X1 U4630 ( .C1(n3923), .C2(n4500), .A(n3922), .B(n3921), .ZN(n4192)
         );
  INV_X1 U4631 ( .A(n3924), .ZN(n3925) );
  OAI21_X1 U4632 ( .B1(n3940), .B2(n3926), .A(n3925), .ZN(n4270) );
  AOI22_X1 U4633 ( .A1(n3927), .A2(n4503), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4507), .ZN(n3928) );
  OAI21_X1 U4634 ( .B1(n4270), .B2(n4096), .A(n3928), .ZN(n3929) );
  AOI21_X1 U4635 ( .B1(n4192), .B2(n4147), .A(n3929), .ZN(n3930) );
  OAI21_X1 U4636 ( .B1(n3931), .B2(n4150), .A(n3930), .ZN(U3263) );
  XNOR2_X1 U4637 ( .A(n3932), .B(n3933), .ZN(n4197) );
  INV_X1 U4638 ( .A(n4197), .ZN(n3948) );
  XNOR2_X1 U4639 ( .A(n3934), .B(n3933), .ZN(n3939) );
  OAI22_X1 U4640 ( .A1(n3935), .A2(n4478), .B1(n3942), .B2(n4477), .ZN(n3936)
         );
  AOI21_X1 U4641 ( .B1(n3937), .B2(n4481), .A(n3936), .ZN(n3938) );
  OAI21_X1 U4642 ( .B1(n3939), .B2(n4483), .A(n3938), .ZN(n4196) );
  INV_X1 U4643 ( .A(n3961), .ZN(n3943) );
  INV_X1 U4644 ( .A(n3940), .ZN(n3941) );
  OAI21_X1 U4645 ( .B1(n3943), .B2(n3942), .A(n3941), .ZN(n4274) );
  AOI22_X1 U4646 ( .A1(n3944), .A2(n4503), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4507), .ZN(n3945) );
  OAI21_X1 U4647 ( .B1(n4274), .B2(n4096), .A(n3945), .ZN(n3946) );
  AOI21_X1 U4648 ( .B1(n4196), .B2(n4147), .A(n3946), .ZN(n3947) );
  OAI21_X1 U4649 ( .B1(n3948), .B2(n4150), .A(n3947), .ZN(U3264) );
  XNOR2_X1 U4650 ( .A(n3949), .B(n3953), .ZN(n4201) );
  INV_X1 U4651 ( .A(n4201), .ZN(n3967) );
  OAI21_X1 U4652 ( .B1(n3971), .B2(n3951), .A(n3950), .ZN(n3952) );
  XOR2_X1 U4653 ( .A(n3953), .B(n3952), .Z(n3958) );
  OAI22_X1 U4654 ( .A1(n4005), .A2(n4478), .B1(n3954), .B2(n4477), .ZN(n3955)
         );
  AOI21_X1 U4655 ( .B1(n3956), .B2(n4481), .A(n3955), .ZN(n3957) );
  OAI21_X1 U4656 ( .B1(n3958), .B2(n4483), .A(n3957), .ZN(n4200) );
  NAND2_X1 U4657 ( .A1(n3979), .A2(n3959), .ZN(n3960) );
  NAND2_X1 U4658 ( .A1(n3961), .A2(n3960), .ZN(n4278) );
  NOR2_X1 U4659 ( .A1(n4278), .A2(n4096), .ZN(n3965) );
  OAI22_X1 U4660 ( .A1(n3963), .A2(n4166), .B1(n3962), .B2(n4147), .ZN(n3964)
         );
  AOI211_X1 U4661 ( .C1(n4200), .C2(n4147), .A(n3965), .B(n3964), .ZN(n3966)
         );
  OAI21_X1 U4662 ( .B1(n3967), .B2(n4150), .A(n3966), .ZN(U3265) );
  XNOR2_X1 U4663 ( .A(n3968), .B(n3972), .ZN(n4205) );
  INV_X1 U4664 ( .A(n4205), .ZN(n3986) );
  INV_X1 U4665 ( .A(n3969), .ZN(n3970) );
  NOR2_X1 U4666 ( .A1(n3971), .A2(n3970), .ZN(n3973) );
  XNOR2_X1 U4667 ( .A(n3973), .B(n3972), .ZN(n3978) );
  OAI22_X1 U4668 ( .A1(n3974), .A2(n4478), .B1(n4477), .B2(n3980), .ZN(n3975)
         );
  AOI21_X1 U4669 ( .B1(n4481), .B2(n3976), .A(n3975), .ZN(n3977) );
  OAI21_X1 U4670 ( .B1(n3978), .B2(n4483), .A(n3977), .ZN(n4204) );
  OAI21_X1 U4671 ( .B1(n4008), .B2(n3980), .A(n3979), .ZN(n4281) );
  NOR2_X1 U4672 ( .A1(n4281), .A2(n4096), .ZN(n3984) );
  INV_X1 U4673 ( .A(REG2_REG_24__SCAN_IN), .ZN(n3981) );
  OAI22_X1 U4674 ( .A1(n3982), .A2(n4166), .B1(n4147), .B2(n3981), .ZN(n3983)
         );
  AOI211_X1 U4675 ( .C1(n4204), .C2(n4147), .A(n3984), .B(n3983), .ZN(n3985)
         );
  OAI21_X1 U4676 ( .B1(n3986), .B2(n4150), .A(n3985), .ZN(U3266) );
  XOR2_X1 U4677 ( .A(n3999), .B(n3987), .Z(n4208) );
  INV_X1 U4678 ( .A(n4208), .ZN(n4014) );
  NAND2_X1 U4679 ( .A1(n4119), .A2(n3988), .ZN(n3991) );
  INV_X1 U4680 ( .A(n3989), .ZN(n3990) );
  NAND2_X1 U4681 ( .A1(n3991), .A2(n3990), .ZN(n4100) );
  NAND2_X1 U4682 ( .A1(n4100), .A2(n3992), .ZN(n4059) );
  INV_X1 U4683 ( .A(n3993), .ZN(n3994) );
  NAND2_X1 U4684 ( .A1(n4059), .A2(n3994), .ZN(n3996) );
  NAND2_X1 U4685 ( .A1(n3996), .A2(n3995), .ZN(n4038) );
  NAND2_X1 U4686 ( .A1(n4035), .A2(n3997), .ZN(n4016) );
  INV_X1 U4687 ( .A(n4023), .ZN(n4017) );
  NAND2_X1 U4688 ( .A1(n4016), .A2(n4017), .ZN(n4015) );
  NAND2_X1 U4689 ( .A1(n4015), .A2(n3998), .ZN(n4000) );
  XNOR2_X1 U4690 ( .A(n4000), .B(n3999), .ZN(n4001) );
  NAND2_X1 U4691 ( .A1(n4001), .A2(n4497), .ZN(n4004) );
  AOI22_X1 U4692 ( .A1(n4040), .A2(n4088), .B1(n4182), .B2(n4002), .ZN(n4003)
         );
  OAI211_X1 U4693 ( .C1(n4005), .C2(n4500), .A(n4004), .B(n4003), .ZN(n4207)
         );
  NOR2_X1 U4694 ( .A1(n4028), .A2(n4006), .ZN(n4007) );
  OR2_X1 U4695 ( .A1(n4008), .A2(n4007), .ZN(n4285) );
  INV_X1 U4696 ( .A(n4009), .ZN(n4010) );
  AOI22_X1 U4697 ( .A1(n4507), .A2(REG2_REG_23__SCAN_IN), .B1(n4010), .B2(
        n4503), .ZN(n4011) );
  OAI21_X1 U4698 ( .B1(n4285), .B2(n4096), .A(n4011), .ZN(n4012) );
  AOI21_X1 U4699 ( .B1(n4207), .B2(n4147), .A(n4012), .ZN(n4013) );
  OAI21_X1 U4700 ( .B1(n4014), .B2(n4150), .A(n4013), .ZN(U3267) );
  OAI21_X1 U4701 ( .B1(n4017), .B2(n4016), .A(n4015), .ZN(n4022) );
  NAND2_X1 U4702 ( .A1(n4018), .A2(n4481), .ZN(n4020) );
  NAND2_X1 U4703 ( .A1(n4063), .A2(n4088), .ZN(n4019) );
  OAI211_X1 U4704 ( .C1(n4477), .C2(n4026), .A(n4020), .B(n4019), .ZN(n4021)
         );
  AOI21_X1 U4705 ( .B1(n4022), .B2(n4497), .A(n4021), .ZN(n4214) );
  INV_X1 U4706 ( .A(n4212), .ZN(n4025) );
  OR2_X1 U4707 ( .A1(n4024), .A2(n4023), .ZN(n4211) );
  NAND3_X1 U4708 ( .A1(n4025), .A2(n4131), .A3(n4211), .ZN(n4033) );
  NOR2_X1 U4709 ( .A1(n4045), .A2(n4026), .ZN(n4027) );
  OR2_X1 U4710 ( .A1(n4028), .A2(n4027), .ZN(n4289) );
  INV_X1 U4711 ( .A(n4289), .ZN(n4031) );
  OAI22_X1 U4712 ( .A1(n4147), .A2(n4842), .B1(n4029), .B2(n4166), .ZN(n4030)
         );
  AOI21_X1 U4713 ( .B1(n4031), .B2(n4491), .A(n4030), .ZN(n4032) );
  OAI211_X1 U4714 ( .C1(n4507), .C2(n4214), .A(n4033), .B(n4032), .ZN(U3268)
         );
  XNOR2_X1 U4715 ( .A(n4034), .B(n4037), .ZN(n4219) );
  INV_X1 U4716 ( .A(n4219), .ZN(n4055) );
  INV_X1 U4717 ( .A(n4035), .ZN(n4036) );
  AOI21_X1 U4718 ( .B1(n4038), .B2(n4037), .A(n4036), .ZN(n4044) );
  AOI22_X1 U4719 ( .A1(n4040), .A2(n4481), .B1(n4182), .B2(n4039), .ZN(n4043)
         );
  NAND2_X1 U4720 ( .A1(n4041), .A2(n4088), .ZN(n4042) );
  OAI211_X1 U4721 ( .C1(n4044), .C2(n4483), .A(n4043), .B(n4042), .ZN(n4218)
         );
  INV_X1 U4722 ( .A(n4224), .ZN(n4048) );
  INV_X1 U4723 ( .A(n4045), .ZN(n4046) );
  OAI21_X1 U4724 ( .B1(n4048), .B2(n4047), .A(n4046), .ZN(n4293) );
  NOR2_X1 U4725 ( .A1(n4293), .A2(n4096), .ZN(n4053) );
  INV_X1 U4726 ( .A(n4049), .ZN(n4050) );
  OAI22_X1 U4727 ( .A1(n4147), .A2(n4051), .B1(n4050), .B2(n4166), .ZN(n4052)
         );
  AOI211_X1 U4728 ( .C1(n4218), .C2(n4147), .A(n4053), .B(n4052), .ZN(n4054)
         );
  OAI21_X1 U4729 ( .B1(n4055), .B2(n4150), .A(n4054), .ZN(U3269) );
  XNOR2_X1 U4730 ( .A(n4056), .B(n4060), .ZN(n4222) );
  NAND2_X1 U4731 ( .A1(n4222), .A2(n4498), .ZN(n4070) );
  INV_X1 U4732 ( .A(n4057), .ZN(n4058) );
  NAND2_X1 U4733 ( .A1(n4059), .A2(n4058), .ZN(n4062) );
  INV_X1 U4734 ( .A(n4060), .ZN(n4061) );
  XNOR2_X1 U4735 ( .A(n4062), .B(n4061), .ZN(n4068) );
  NAND2_X1 U4736 ( .A1(n4102), .A2(n4088), .ZN(n4065) );
  NAND2_X1 U4737 ( .A1(n4063), .A2(n4481), .ZN(n4064) );
  OAI211_X1 U4738 ( .C1(n4477), .C2(n4066), .A(n4065), .B(n4064), .ZN(n4067)
         );
  AOI21_X1 U4739 ( .B1(n4068), .B2(n4497), .A(n4067), .ZN(n4069) );
  NAND2_X1 U4740 ( .A1(n4070), .A2(n4069), .ZN(n4228) );
  INV_X1 U4741 ( .A(n4228), .ZN(n4078) );
  NAND2_X1 U4742 ( .A1(n4093), .A2(n4071), .ZN(n4223) );
  AND3_X1 U4743 ( .A1(n4224), .A2(n4491), .A3(n4223), .ZN(n4076) );
  INV_X1 U4744 ( .A(n4072), .ZN(n4073) );
  OAI22_X1 U4745 ( .A1(n4147), .A2(n4074), .B1(n4073), .B2(n4166), .ZN(n4075)
         );
  AOI211_X1 U4746 ( .C1(n4222), .C2(n4504), .A(n4076), .B(n4075), .ZN(n4077)
         );
  OAI21_X1 U4747 ( .B1(n4078), .B2(n4507), .A(n4077), .ZN(U3270) );
  XNOR2_X1 U4748 ( .A(n4079), .B(n4084), .ZN(n4230) );
  INV_X1 U4749 ( .A(n4230), .ZN(n4099) );
  INV_X1 U4750 ( .A(n4080), .ZN(n4082) );
  OAI21_X1 U4751 ( .B1(n4100), .B2(n4082), .A(n4081), .ZN(n4083) );
  XOR2_X1 U4752 ( .A(n4084), .B(n4083), .Z(n4090) );
  OAI22_X1 U4753 ( .A1(n4086), .A2(n4500), .B1(n4477), .B2(n4085), .ZN(n4087)
         );
  AOI21_X1 U4754 ( .B1(n4088), .B2(n4930), .A(n4087), .ZN(n4089) );
  OAI21_X1 U4755 ( .B1(n4090), .B2(n4483), .A(n4089), .ZN(n4229) );
  NAND2_X1 U4756 ( .A1(n4111), .A2(n4091), .ZN(n4092) );
  NAND2_X1 U4757 ( .A1(n4093), .A2(n4092), .ZN(n4298) );
  AOI22_X1 U4758 ( .A1(n4507), .A2(REG2_REG_19__SCAN_IN), .B1(n4094), .B2(
        n4503), .ZN(n4095) );
  OAI21_X1 U4759 ( .B1(n4298), .B2(n4096), .A(n4095), .ZN(n4097) );
  AOI21_X1 U4760 ( .B1(n4229), .B2(n4147), .A(n4097), .ZN(n4098) );
  OAI21_X1 U4761 ( .B1(n4099), .B2(n4150), .A(n4098), .ZN(U3271) );
  XNOR2_X1 U4762 ( .A(n4100), .B(n4110), .ZN(n4106) );
  AOI22_X1 U4763 ( .A1(n4102), .A2(n4481), .B1(n4101), .B2(n4182), .ZN(n4103)
         );
  OAI21_X1 U4764 ( .B1(n4104), .B2(n4478), .A(n4103), .ZN(n4105) );
  AOI21_X1 U4765 ( .B1(n4106), .B2(n4497), .A(n4105), .ZN(n4233) );
  INV_X1 U4766 ( .A(n4108), .ZN(n4109) );
  AOI21_X1 U4767 ( .B1(n4110), .B2(n4107), .A(n4109), .ZN(n4234) );
  INV_X1 U4768 ( .A(n4234), .ZN(n4117) );
  OAI211_X1 U4769 ( .C1(n4124), .C2(n4112), .A(n4111), .B(n4570), .ZN(n4232)
         );
  AOI22_X1 U4770 ( .A1(n4507), .A2(REG2_REG_18__SCAN_IN), .B1(n4113), .B2(
        n4503), .ZN(n4114) );
  OAI21_X1 U4771 ( .B1(n4232), .B2(n4115), .A(n4114), .ZN(n4116) );
  AOI21_X1 U4772 ( .B1(n4117), .B2(n4131), .A(n4116), .ZN(n4118) );
  OAI21_X1 U4773 ( .B1(n4507), .B2(n4233), .A(n4118), .ZN(U3272) );
  XNOR2_X1 U4774 ( .A(n4119), .B(n4129), .ZN(n4123) );
  NOR2_X1 U4775 ( .A1(n4927), .A2(n4478), .ZN(n4122) );
  OAI22_X1 U4776 ( .A1(n4120), .A2(n4500), .B1(n4477), .B2(n4936), .ZN(n4121)
         );
  AOI211_X1 U4777 ( .C1(n4123), .C2(n4497), .A(n4122), .B(n4121), .ZN(n4235)
         );
  INV_X1 U4778 ( .A(n4124), .ZN(n4125) );
  OAI21_X1 U4779 ( .B1(n2305), .B2(n4936), .A(n4125), .ZN(n4303) );
  INV_X1 U4780 ( .A(n4303), .ZN(n4128) );
  INV_X1 U4781 ( .A(n4932), .ZN(n4126) );
  OAI22_X1 U4782 ( .A1(n4147), .A2(n4855), .B1(n4126), .B2(n4166), .ZN(n4127)
         );
  AOI21_X1 U4783 ( .B1(n4128), .B2(n4491), .A(n4127), .ZN(n4133) );
  XNOR2_X1 U4784 ( .A(n4130), .B(n4129), .ZN(n4237) );
  NAND2_X1 U4785 ( .A1(n4237), .A2(n4131), .ZN(n4132) );
  OAI211_X1 U4786 ( .C1(n4235), .C2(n4507), .A(n4133), .B(n4132), .ZN(U3273)
         );
  XNOR2_X1 U4787 ( .A(n4134), .B(n4136), .ZN(n4243) );
  XOR2_X1 U4788 ( .A(n4136), .B(n4135), .Z(n4141) );
  AOI22_X1 U4789 ( .A1(n4137), .A2(n4481), .B1(n4142), .B2(n4182), .ZN(n4138)
         );
  OAI21_X1 U4790 ( .B1(n4139), .B2(n4478), .A(n4138), .ZN(n4140) );
  AOI21_X1 U4791 ( .B1(n4141), .B2(n4497), .A(n4140), .ZN(n4242) );
  INV_X1 U4792 ( .A(n4242), .ZN(n4148) );
  NAND2_X1 U4793 ( .A1(n2200), .A2(n4142), .ZN(n4239) );
  AND3_X1 U4794 ( .A1(n4240), .A2(n4491), .A3(n4239), .ZN(n4146) );
  INV_X1 U4795 ( .A(n4143), .ZN(n4144) );
  OAI22_X1 U4796 ( .A1(n4147), .A2(n4435), .B1(n4144), .B2(n4166), .ZN(n4145)
         );
  AOI211_X1 U4797 ( .C1(n4148), .C2(n4147), .A(n4146), .B(n4145), .ZN(n4149)
         );
  OAI21_X1 U4798 ( .B1(n4243), .B2(n4150), .A(n4149), .ZN(U3274) );
  OAI21_X1 U4799 ( .B1(n4158), .B2(n4152), .A(n4151), .ZN(n4162) );
  AOI22_X1 U4800 ( .A1(n4153), .A2(n4481), .B1(n4182), .B2(n4164), .ZN(n4154)
         );
  OAI21_X1 U4801 ( .B1(n4155), .B2(n4478), .A(n4154), .ZN(n4161) );
  AOI21_X1 U4802 ( .B1(n4158), .B2(n4157), .A(n4156), .ZN(n4252) );
  NOR2_X1 U4803 ( .A1(n4252), .A2(n4159), .ZN(n4160) );
  AOI211_X1 U4804 ( .C1(n4497), .C2(n4162), .A(n4161), .B(n4160), .ZN(n4251)
         );
  INV_X1 U4805 ( .A(n4252), .ZN(n4171) );
  INV_X1 U4806 ( .A(n4163), .ZN(n4249) );
  NAND2_X1 U4807 ( .A1(n2199), .A2(n4164), .ZN(n4248) );
  AND3_X1 U4808 ( .A1(n4249), .A2(n4491), .A3(n4248), .ZN(n4170) );
  INV_X1 U4809 ( .A(n4165), .ZN(n4167) );
  OAI22_X1 U4810 ( .A1(n4147), .A2(n4168), .B1(n4167), .B2(n4166), .ZN(n4169)
         );
  AOI211_X1 U4811 ( .C1(n4171), .C2(n4504), .A(n4170), .B(n4169), .ZN(n4172)
         );
  OAI21_X1 U4812 ( .B1(n4251), .B2(n4507), .A(n4172), .ZN(U3276) );
  INV_X1 U4813 ( .A(n4328), .ZN(n4260) );
  INV_X1 U4814 ( .A(n4173), .ZN(n4174) );
  NAND2_X1 U4815 ( .A1(n4175), .A2(n4174), .ZN(n4185) );
  OAI21_X1 U4816 ( .B1(n4176), .B2(n4477), .A(n4185), .ZN(n4327) );
  NAND2_X1 U4817 ( .A1(n4327), .A2(n4604), .ZN(n4178) );
  NAND2_X1 U4818 ( .A1(n4601), .A2(REG1_REG_31__SCAN_IN), .ZN(n4177) );
  OAI211_X1 U4819 ( .C1(n4260), .C2(n4247), .A(n4178), .B(n4177), .ZN(U3549)
         );
  AND2_X1 U4820 ( .A1(n4179), .A2(n4183), .ZN(n4180) );
  NOR2_X1 U4821 ( .A1(n4181), .A2(n4180), .ZN(n4330) );
  INV_X1 U4822 ( .A(n4330), .ZN(n4262) );
  NAND2_X1 U4823 ( .A1(n4183), .A2(n4182), .ZN(n4184) );
  AND2_X1 U4824 ( .A1(n4185), .A2(n4184), .ZN(n4332) );
  INV_X1 U4825 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4186) );
  MUX2_X1 U4826 ( .A(n4332), .B(n4186), .S(n4601), .Z(n4187) );
  OAI21_X1 U4827 ( .B1(n4262), .B2(n4247), .A(n4187), .ZN(U3548) );
  OAI21_X1 U4828 ( .B1(n4189), .B2(n2366), .A(n4188), .ZN(n4263) );
  INV_X1 U4829 ( .A(n4190), .ZN(n4191) );
  OAI21_X1 U4830 ( .B1(n4247), .B2(n4266), .A(n4191), .ZN(U3546) );
  INV_X1 U4831 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4194) );
  AOI21_X1 U4832 ( .B1(n4193), .B2(n4561), .A(n4192), .ZN(n4267) );
  MUX2_X1 U4833 ( .A(n4194), .B(n4267), .S(n4604), .Z(n4195) );
  OAI21_X1 U4834 ( .B1(n4247), .B2(n4270), .A(n4195), .ZN(U3545) );
  INV_X1 U4835 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4198) );
  AOI21_X1 U4836 ( .B1(n4197), .B2(n4561), .A(n4196), .ZN(n4271) );
  MUX2_X1 U4837 ( .A(n4198), .B(n4271), .S(n4604), .Z(n4199) );
  OAI21_X1 U4838 ( .B1(n4247), .B2(n4274), .A(n4199), .ZN(U3544) );
  INV_X1 U4839 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4202) );
  AOI21_X1 U4840 ( .B1(n4201), .B2(n4561), .A(n4200), .ZN(n4275) );
  MUX2_X1 U4841 ( .A(n4202), .B(n4275), .S(n4604), .Z(n4203) );
  OAI21_X1 U4842 ( .B1(n4247), .B2(n4278), .A(n4203), .ZN(U3543) );
  INV_X1 U4843 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4887) );
  AOI21_X1 U4844 ( .B1(n4205), .B2(n4561), .A(n4204), .ZN(n4279) );
  MUX2_X1 U4845 ( .A(n4887), .B(n4279), .S(n4604), .Z(n4206) );
  OAI21_X1 U4846 ( .B1(n4247), .B2(n4281), .A(n4206), .ZN(U3542) );
  INV_X1 U4847 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4209) );
  AOI21_X1 U4848 ( .B1(n4208), .B2(n4561), .A(n4207), .ZN(n4282) );
  MUX2_X1 U4849 ( .A(n4209), .B(n4282), .S(n4604), .Z(n4210) );
  OAI21_X1 U4850 ( .B1(n4247), .B2(n4285), .A(n4210), .ZN(U3541) );
  NAND2_X1 U4851 ( .A1(n4211), .A2(n4561), .ZN(n4213) );
  OR2_X1 U4852 ( .A1(n4213), .A2(n4212), .ZN(n4215) );
  NAND2_X1 U4853 ( .A1(n4215), .A2(n4214), .ZN(n4286) );
  MUX2_X1 U4854 ( .A(n4286), .B(REG1_REG_22__SCAN_IN), .S(n4601), .Z(n4216) );
  INV_X1 U4855 ( .A(n4216), .ZN(n4217) );
  OAI21_X1 U4856 ( .B1(n4247), .B2(n4289), .A(n4217), .ZN(U3540) );
  INV_X1 U4857 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4220) );
  AOI21_X1 U4858 ( .B1(n4219), .B2(n4561), .A(n4218), .ZN(n4290) );
  MUX2_X1 U4859 ( .A(n4220), .B(n4290), .S(n4604), .Z(n4221) );
  OAI21_X1 U4860 ( .B1(n4247), .B2(n4293), .A(n4221), .ZN(U3539) );
  INV_X1 U4861 ( .A(n4222), .ZN(n4226) );
  NAND3_X1 U4862 ( .A1(n4224), .A2(n4570), .A3(n4223), .ZN(n4225) );
  OAI21_X1 U4863 ( .B1(n4226), .B2(n4253), .A(n4225), .ZN(n4227) );
  MUX2_X1 U4864 ( .A(REG1_REG_20__SCAN_IN), .B(n4294), .S(n4604), .Z(U3538) );
  AOI21_X1 U4865 ( .B1(n4561), .B2(n4230), .A(n4229), .ZN(n4295) );
  MUX2_X1 U4866 ( .A(n4790), .B(n4295), .S(n4604), .Z(n4231) );
  OAI21_X1 U4867 ( .B1(n4247), .B2(n4298), .A(n4231), .ZN(U3537) );
  OAI211_X1 U4868 ( .C1(n4234), .C2(n2366), .A(n4233), .B(n4232), .ZN(n4299)
         );
  MUX2_X1 U4869 ( .A(REG1_REG_18__SCAN_IN), .B(n4299), .S(n4604), .Z(U3536) );
  INV_X1 U4870 ( .A(n4235), .ZN(n4236) );
  AOI21_X1 U4871 ( .B1(n4237), .B2(n4561), .A(n4236), .ZN(n4300) );
  MUX2_X1 U4872 ( .A(n3867), .B(n4300), .S(n4604), .Z(n4238) );
  OAI21_X1 U4873 ( .B1(n4247), .B2(n4303), .A(n4238), .ZN(U3535) );
  NAND3_X1 U4874 ( .A1(n4240), .A2(n4570), .A3(n4239), .ZN(n4241) );
  OAI211_X1 U4875 ( .C1(n4243), .C2(n2366), .A(n4242), .B(n4241), .ZN(n4304)
         );
  MUX2_X1 U4876 ( .A(n4304), .B(REG1_REG_16__SCAN_IN), .S(n4601), .Z(U3534) );
  AOI21_X1 U4877 ( .B1(n4245), .B2(n4561), .A(n4244), .ZN(n4305) );
  MUX2_X1 U4878 ( .A(n4852), .B(n4305), .S(n4604), .Z(n4246) );
  OAI21_X1 U4879 ( .B1(n4247), .B2(n4309), .A(n4246), .ZN(U3533) );
  NAND3_X1 U4880 ( .A1(n4249), .A2(n4570), .A3(n4248), .ZN(n4250) );
  OAI211_X1 U4881 ( .C1(n4252), .C2(n4253), .A(n4251), .B(n4250), .ZN(n4310)
         );
  MUX2_X1 U4882 ( .A(REG1_REG_14__SCAN_IN), .B(n4310), .S(n4604), .Z(U3532) );
  NAND2_X1 U4883 ( .A1(n4254), .A2(n4583), .ZN(n4255) );
  OAI211_X1 U4884 ( .C1(n4577), .C2(n4257), .A(n4256), .B(n4255), .ZN(n4311)
         );
  MUX2_X1 U4885 ( .A(REG1_REG_13__SCAN_IN), .B(n4311), .S(n4604), .Z(U3531) );
  NAND2_X1 U4886 ( .A1(n4327), .A2(n4585), .ZN(n4259) );
  NAND2_X1 U4887 ( .A1(n4584), .A2(REG0_REG_31__SCAN_IN), .ZN(n4258) );
  OAI211_X1 U4888 ( .C1(n4260), .C2(n4308), .A(n4259), .B(n4258), .ZN(U3517)
         );
  INV_X1 U4889 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4760) );
  MUX2_X1 U4890 ( .A(n4332), .B(n4760), .S(n4584), .Z(n4261) );
  OAI21_X1 U4891 ( .B1(n4262), .B2(n4308), .A(n4261), .ZN(U3516) );
  INV_X1 U4892 ( .A(n4264), .ZN(n4265) );
  OAI21_X1 U4893 ( .B1(n4266), .B2(n4308), .A(n4265), .ZN(U3514) );
  INV_X1 U4894 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4268) );
  MUX2_X1 U4895 ( .A(n4268), .B(n4267), .S(n4585), .Z(n4269) );
  OAI21_X1 U4896 ( .B1(n4270), .B2(n4308), .A(n4269), .ZN(U3513) );
  INV_X1 U4897 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4272) );
  MUX2_X1 U4898 ( .A(n4272), .B(n4271), .S(n4585), .Z(n4273) );
  OAI21_X1 U4899 ( .B1(n4274), .B2(n4308), .A(n4273), .ZN(U3512) );
  INV_X1 U4900 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4276) );
  MUX2_X1 U4901 ( .A(n4276), .B(n4275), .S(n4585), .Z(n4277) );
  OAI21_X1 U4902 ( .B1(n4278), .B2(n4308), .A(n4277), .ZN(U3511) );
  INV_X1 U4903 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4886) );
  MUX2_X1 U4904 ( .A(n4886), .B(n4279), .S(n4585), .Z(n4280) );
  OAI21_X1 U4905 ( .B1(n4281), .B2(n4308), .A(n4280), .ZN(U3510) );
  INV_X1 U4906 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4283) );
  MUX2_X1 U4907 ( .A(n4283), .B(n4282), .S(n4585), .Z(n4284) );
  OAI21_X1 U4908 ( .B1(n4285), .B2(n4308), .A(n4284), .ZN(U3509) );
  MUX2_X1 U4909 ( .A(n4286), .B(REG0_REG_22__SCAN_IN), .S(n4584), .Z(n4287) );
  INV_X1 U4910 ( .A(n4287), .ZN(n4288) );
  OAI21_X1 U4911 ( .B1(n4289), .B2(n4308), .A(n4288), .ZN(U3508) );
  INV_X1 U4912 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4291) );
  MUX2_X1 U4913 ( .A(n4291), .B(n4290), .S(n4585), .Z(n4292) );
  OAI21_X1 U4914 ( .B1(n4293), .B2(n4308), .A(n4292), .ZN(U3507) );
  MUX2_X1 U4915 ( .A(n4294), .B(REG0_REG_20__SCAN_IN), .S(n4584), .Z(U3506) );
  INV_X1 U4916 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4296) );
  MUX2_X1 U4917 ( .A(n4296), .B(n4295), .S(n4585), .Z(n4297) );
  OAI21_X1 U4918 ( .B1(n4298), .B2(n4308), .A(n4297), .ZN(U3505) );
  MUX2_X1 U4919 ( .A(REG0_REG_18__SCAN_IN), .B(n4299), .S(n4585), .Z(U3503) );
  INV_X1 U4920 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4301) );
  MUX2_X1 U4921 ( .A(n4301), .B(n4300), .S(n4585), .Z(n4302) );
  OAI21_X1 U4922 ( .B1(n4303), .B2(n4308), .A(n4302), .ZN(U3501) );
  MUX2_X1 U4923 ( .A(n4304), .B(REG0_REG_16__SCAN_IN), .S(n4584), .Z(U3499) );
  INV_X1 U4924 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4306) );
  MUX2_X1 U4925 ( .A(n4306), .B(n4305), .S(n4585), .Z(n4307) );
  OAI21_X1 U4926 ( .B1(n4309), .B2(n4308), .A(n4307), .ZN(U3497) );
  MUX2_X1 U4927 ( .A(REG0_REG_14__SCAN_IN), .B(n4310), .S(n4585), .Z(U3495) );
  MUX2_X1 U4928 ( .A(REG0_REG_13__SCAN_IN), .B(n4311), .S(n4585), .Z(U3493) );
  MUX2_X1 U4929 ( .A(DATAI_30_), .B(n4312), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4930 ( .A(DATAI_28_), .B(n4313), .S(STATE_REG_SCAN_IN), .Z(U3324)
         );
  MUX2_X1 U4931 ( .A(n4314), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U4932 ( .A(DATAI_25_), .B(n4315), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U4933 ( .A(n4316), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U4934 ( .A(n4317), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U4935 ( .A(n4318), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U4936 ( .A(DATAI_20_), .B(n4319), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4937 ( .A(DATAI_19_), .B(n4320), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U4938 ( .A(DATAI_17_), .B(n4321), .S(STATE_REG_SCAN_IN), .Z(U3335)
         );
  MUX2_X1 U4939 ( .A(n4322), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U4940 ( .A(DATAI_4_), .B(n4323), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4941 ( .A(n4324), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4942 ( .A(n4325), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4943 ( .A(n4326), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U4944 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(STATE_REG_SCAN_IN), 
        .Z(U3352) );
  AOI22_X1 U4945 ( .A1(n4328), .A2(n4491), .B1(n4147), .B2(n4327), .ZN(n4329)
         );
  OAI21_X1 U4946 ( .B1(n4147), .B2(n3715), .A(n4329), .ZN(U3260) );
  AOI22_X1 U4947 ( .A1(n4330), .A2(n4491), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4507), .ZN(n4331) );
  OAI21_X1 U4948 ( .B1(n4507), .B2(n4332), .A(n4331), .ZN(U3261) );
  AOI211_X1 U4949 ( .C1(n4335), .C2(n4334), .A(n4333), .B(n4343), .ZN(n4336)
         );
  AOI211_X1 U4950 ( .C1(n4451), .C2(ADDR_REG_5__SCAN_IN), .A(n4337), .B(n4336), 
        .ZN(n4342) );
  OAI211_X1 U4951 ( .C1(n4340), .C2(n4339), .A(n4407), .B(n4338), .ZN(n4341)
         );
  OAI211_X1 U4952 ( .C1(n4458), .C2(n4528), .A(n4342), .B(n4341), .ZN(U3245)
         );
  AOI211_X1 U4953 ( .C1(n4868), .C2(n4345), .A(n4344), .B(n4343), .ZN(n4346)
         );
  AOI211_X1 U4954 ( .C1(n4451), .C2(ADDR_REG_6__SCAN_IN), .A(n4347), .B(n4346), 
        .ZN(n4351) );
  OAI211_X1 U4955 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4349), .A(n4407), .B(n4348), 
        .ZN(n4350) );
  OAI211_X1 U4956 ( .C1(n4458), .C2(n4352), .A(n4351), .B(n4350), .ZN(U3246)
         );
  NAND2_X1 U4957 ( .A1(n4354), .A2(n4353), .ZN(n4356) );
  OAI21_X1 U4958 ( .B1(n4357), .B2(n4356), .A(n4453), .ZN(n4355) );
  AOI21_X1 U4959 ( .B1(n4357), .B2(n4356), .A(n4355), .ZN(n4358) );
  AOI211_X1 U4960 ( .C1(n4451), .C2(ADDR_REG_7__SCAN_IN), .A(n4359), .B(n4358), 
        .ZN(n4364) );
  OAI211_X1 U4961 ( .C1(n4362), .C2(n4361), .A(n4407), .B(n4360), .ZN(n4363)
         );
  OAI211_X1 U4962 ( .C1(n4458), .C2(n4524), .A(n4364), .B(n4363), .ZN(U3247)
         );
  OAI211_X1 U4963 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4366), .A(n4453), .B(n4365), 
        .ZN(n4370) );
  OAI211_X1 U4964 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4368), .A(n4407), .B(n4367), 
        .ZN(n4369) );
  OAI211_X1 U4965 ( .C1(n4458), .C2(n4522), .A(n4370), .B(n4369), .ZN(n4371)
         );
  AOI211_X1 U4966 ( .C1(n4451), .C2(ADDR_REG_8__SCAN_IN), .A(n4372), .B(n4371), 
        .ZN(n4373) );
  INV_X1 U4967 ( .A(n4373), .ZN(U3248) );
  OAI211_X1 U4968 ( .C1(n4376), .C2(n4375), .A(n4453), .B(n4374), .ZN(n4381)
         );
  OAI211_X1 U4969 ( .C1(n4379), .C2(n4378), .A(n4407), .B(n4377), .ZN(n4380)
         );
  OAI211_X1 U4970 ( .C1(n4458), .C2(n4521), .A(n4381), .B(n4380), .ZN(n4382)
         );
  AOI211_X1 U4971 ( .C1(n4451), .C2(ADDR_REG_9__SCAN_IN), .A(n4383), .B(n4382), 
        .ZN(n4384) );
  INV_X1 U4972 ( .A(n4384), .ZN(U3249) );
  OAI211_X1 U4973 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4386), .A(n4453), .B(n4385), .ZN(n4390) );
  OAI211_X1 U4974 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4388), .A(n4407), .B(n4387), .ZN(n4389) );
  OAI211_X1 U4975 ( .C1(n4458), .C2(n4391), .A(n4390), .B(n4389), .ZN(n4392)
         );
  AOI211_X1 U4976 ( .C1(n4451), .C2(ADDR_REG_10__SCAN_IN), .A(n4393), .B(n4392), .ZN(n4394) );
  INV_X1 U4977 ( .A(n4394), .ZN(U3250) );
  OAI211_X1 U4978 ( .C1(n4397), .C2(n4396), .A(n4453), .B(n4395), .ZN(n4402)
         );
  OAI211_X1 U4979 ( .C1(n4400), .C2(n4399), .A(n4407), .B(n4398), .ZN(n4401)
         );
  OAI211_X1 U4980 ( .C1(n4458), .C2(n4518), .A(n4402), .B(n4401), .ZN(n4403)
         );
  AOI211_X1 U4981 ( .C1(n4451), .C2(ADDR_REG_11__SCAN_IN), .A(n4404), .B(n4403), .ZN(n4405) );
  INV_X1 U4982 ( .A(n4405), .ZN(U3251) );
  OAI211_X1 U4983 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4408), .A(n4407), .B(n4406), .ZN(n4410) );
  NAND2_X1 U4984 ( .A1(n4410), .A2(n4409), .ZN(n4411) );
  AOI21_X1 U4985 ( .B1(n4451), .B2(ADDR_REG_12__SCAN_IN), .A(n4411), .ZN(n4415) );
  OAI211_X1 U4986 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4413), .A(n4453), .B(n4412), .ZN(n4414) );
  OAI211_X1 U4987 ( .C1(n4458), .C2(n4517), .A(n4415), .B(n4414), .ZN(U3252)
         );
  INV_X1 U4988 ( .A(n4416), .ZN(n4420) );
  AOI211_X1 U4989 ( .C1(n4168), .C2(n4418), .A(n4417), .B(n4445), .ZN(n4419)
         );
  AOI211_X1 U4990 ( .C1(ADDR_REG_14__SCAN_IN), .C2(n4451), .A(n4420), .B(n4419), .ZN(n4424) );
  OAI211_X1 U4991 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4422), .A(n4453), .B(n4421), .ZN(n4423) );
  OAI211_X1 U4992 ( .C1(n4458), .C2(n2208), .A(n4424), .B(n4423), .ZN(U3254)
         );
  AOI211_X1 U4993 ( .C1(n4427), .C2(n4426), .A(n4425), .B(n4445), .ZN(n4428)
         );
  AOI211_X1 U4994 ( .C1(n4451), .C2(ADDR_REG_15__SCAN_IN), .A(n4429), .B(n4428), .ZN(n4434) );
  OAI211_X1 U4995 ( .C1(n4432), .C2(n4431), .A(n4453), .B(n4430), .ZN(n4433)
         );
  OAI211_X1 U4996 ( .C1(n4458), .C2(n4516), .A(n4434), .B(n4433), .ZN(U3255)
         );
  AOI221_X1 U4997 ( .B1(n4437), .B2(n4436), .C1(n4435), .C2(n4436), .A(n4445), 
        .ZN(n4438) );
  AOI211_X1 U4998 ( .C1(ADDR_REG_16__SCAN_IN), .C2(n4451), .A(n4439), .B(n4438), .ZN(n4443) );
  OAI221_X1 U4999 ( .B1(n4441), .B2(REG1_REG_16__SCAN_IN), .C1(n4441), .C2(
        n4440), .A(n4453), .ZN(n4442) );
  OAI211_X1 U5000 ( .C1(n4458), .C2(n4515), .A(n4443), .B(n4442), .ZN(U3256)
         );
  INV_X1 U5001 ( .A(n4444), .ZN(n4450) );
  AOI211_X1 U5002 ( .C1(n4448), .C2(n4447), .A(n4446), .B(n4445), .ZN(n4449)
         );
  OAI211_X1 U5003 ( .C1(n4455), .C2(n4454), .A(n4453), .B(n4452), .ZN(n4456)
         );
  OAI211_X1 U5004 ( .C1(n4458), .C2(n4513), .A(n4457), .B(n4456), .ZN(U3258)
         );
  XNOR2_X1 U5005 ( .A(n2192), .B(n4459), .ZN(n4582) );
  XNOR2_X1 U5006 ( .A(n4460), .B(n4459), .ZN(n4465) );
  OAI22_X1 U5007 ( .A1(n4461), .A2(n4478), .B1(n4469), .B2(n4477), .ZN(n4462)
         );
  AOI21_X1 U5008 ( .B1(n4481), .B2(n4463), .A(n4462), .ZN(n4464) );
  OAI21_X1 U5009 ( .B1(n4465), .B2(n4483), .A(n4464), .ZN(n4466) );
  AOI21_X1 U5010 ( .B1(n4498), .B2(n4582), .A(n4466), .ZN(n4579) );
  AOI22_X1 U5011 ( .A1(n4467), .A2(n4503), .B1(REG2_REG_11__SCAN_IN), .B2(
        n4507), .ZN(n4473) );
  INV_X1 U5012 ( .A(n4572), .ZN(n4470) );
  OAI21_X1 U5013 ( .B1(n4470), .B2(n4469), .A(n4468), .ZN(n4578) );
  INV_X1 U5014 ( .A(n4578), .ZN(n4471) );
  AOI22_X1 U5015 ( .A1(n4582), .A2(n4504), .B1(n4491), .B2(n4471), .ZN(n4472)
         );
  OAI211_X1 U5016 ( .C1(n4507), .C2(n4579), .A(n4473), .B(n4472), .ZN(U3279)
         );
  XOR2_X1 U5017 ( .A(n4476), .B(n4474), .Z(n4547) );
  XOR2_X1 U5018 ( .A(n4476), .B(n4475), .Z(n4484) );
  OAI22_X1 U5019 ( .A1(n2959), .A2(n4478), .B1(n4477), .B2(n4488), .ZN(n4479)
         );
  AOI21_X1 U5020 ( .B1(n4481), .B2(n4480), .A(n4479), .ZN(n4482) );
  OAI21_X1 U5021 ( .B1(n4484), .B2(n4483), .A(n4482), .ZN(n4485) );
  AOI21_X1 U5022 ( .B1(n4498), .B2(n4547), .A(n4485), .ZN(n4544) );
  AOI22_X1 U5023 ( .A1(n4507), .A2(REG2_REG_3__SCAN_IN), .B1(n4503), .B2(n4486), .ZN(n4493) );
  OAI21_X1 U5024 ( .B1(n4489), .B2(n4488), .A(n4487), .ZN(n4543) );
  INV_X1 U5025 ( .A(n4543), .ZN(n4490) );
  AOI22_X1 U5026 ( .A1(n4547), .A2(n4504), .B1(n4491), .B2(n4490), .ZN(n4492)
         );
  OAI211_X1 U5027 ( .C1(n4507), .C2(n4544), .A(n4493), .B(n4492), .ZN(U3287)
         );
  INV_X1 U5028 ( .A(n4494), .ZN(n4495) );
  NOR2_X1 U5029 ( .A1(n4496), .A2(n4495), .ZN(n4530) );
  OAI21_X1 U5030 ( .B1(n4498), .B2(n4497), .A(n4531), .ZN(n4499) );
  OAI21_X1 U5031 ( .B1(n4501), .B2(n4500), .A(n4499), .ZN(n4529) );
  AOI21_X1 U5032 ( .B1(n4530), .B2(n4502), .A(n4529), .ZN(n4506) );
  AOI22_X1 U5033 ( .A1(n4531), .A2(n4504), .B1(REG3_REG_0__SCAN_IN), .B2(n4503), .ZN(n4505) );
  OAI221_X1 U5034 ( .B1(n4507), .B2(n4506), .C1(n4147), .C2(n2451), .A(n4505), 
        .ZN(U3290) );
  AND2_X1 U5035 ( .A1(D_REG_31__SCAN_IN), .A2(n4508), .ZN(U3291) );
  AND2_X1 U5036 ( .A1(D_REG_30__SCAN_IN), .A2(n4508), .ZN(U3292) );
  AND2_X1 U5037 ( .A1(D_REG_29__SCAN_IN), .A2(n4508), .ZN(U3293) );
  AND2_X1 U5038 ( .A1(D_REG_28__SCAN_IN), .A2(n4508), .ZN(U3294) );
  INV_X1 U5039 ( .A(D_REG_27__SCAN_IN), .ZN(n4675) );
  NOR2_X1 U5040 ( .A1(n4509), .A2(n4675), .ZN(U3295) );
  AND2_X1 U5041 ( .A1(D_REG_26__SCAN_IN), .A2(n4508), .ZN(U3296) );
  AND2_X1 U5042 ( .A1(D_REG_25__SCAN_IN), .A2(n4508), .ZN(U3297) );
  NOR2_X1 U5043 ( .A1(n4509), .A2(n4742), .ZN(U3298) );
  INV_X1 U5044 ( .A(D_REG_23__SCAN_IN), .ZN(n4773) );
  NOR2_X1 U5045 ( .A1(n4509), .A2(n4773), .ZN(U3299) );
  INV_X1 U5046 ( .A(D_REG_22__SCAN_IN), .ZN(n4672) );
  NOR2_X1 U5047 ( .A1(n4509), .A2(n4672), .ZN(U3300) );
  AND2_X1 U5048 ( .A1(D_REG_21__SCAN_IN), .A2(n4508), .ZN(U3301) );
  AND2_X1 U5049 ( .A1(D_REG_20__SCAN_IN), .A2(n4508), .ZN(U3302) );
  INV_X1 U5050 ( .A(D_REG_19__SCAN_IN), .ZN(n4677) );
  NOR2_X1 U5051 ( .A1(n4509), .A2(n4677), .ZN(U3303) );
  AND2_X1 U5052 ( .A1(D_REG_18__SCAN_IN), .A2(n4508), .ZN(U3304) );
  INV_X1 U5053 ( .A(D_REG_17__SCAN_IN), .ZN(n4678) );
  NOR2_X1 U5054 ( .A1(n4509), .A2(n4678), .ZN(U3305) );
  AND2_X1 U5055 ( .A1(D_REG_16__SCAN_IN), .A2(n4508), .ZN(U3306) );
  INV_X1 U5056 ( .A(D_REG_15__SCAN_IN), .ZN(n4776) );
  NOR2_X1 U5057 ( .A1(n4509), .A2(n4776), .ZN(U3307) );
  INV_X1 U5058 ( .A(D_REG_14__SCAN_IN), .ZN(n4669) );
  NOR2_X1 U5059 ( .A1(n4509), .A2(n4669), .ZN(U3308) );
  INV_X1 U5060 ( .A(D_REG_13__SCAN_IN), .ZN(n4668) );
  NOR2_X1 U5061 ( .A1(n4509), .A2(n4668), .ZN(U3309) );
  NOR2_X1 U5062 ( .A1(n4509), .A2(n4769), .ZN(U3310) );
  INV_X1 U5063 ( .A(D_REG_11__SCAN_IN), .ZN(n4778) );
  NOR2_X1 U5064 ( .A1(n4509), .A2(n4778), .ZN(U3311) );
  INV_X1 U5065 ( .A(D_REG_10__SCAN_IN), .ZN(n4671) );
  NOR2_X1 U5066 ( .A1(n4509), .A2(n4671), .ZN(U3312) );
  NOR2_X1 U5067 ( .A1(n4509), .A2(n4770), .ZN(U3313) );
  NOR2_X1 U5068 ( .A1(n4509), .A2(n4743), .ZN(U3314) );
  AND2_X1 U5069 ( .A1(D_REG_7__SCAN_IN), .A2(n4508), .ZN(U3315) );
  INV_X1 U5070 ( .A(D_REG_6__SCAN_IN), .ZN(n4775) );
  NOR2_X1 U5071 ( .A1(n4509), .A2(n4775), .ZN(U3316) );
  INV_X1 U5072 ( .A(D_REG_5__SCAN_IN), .ZN(n4779) );
  NOR2_X1 U5073 ( .A1(n4509), .A2(n4779), .ZN(U3317) );
  AND2_X1 U5074 ( .A1(D_REG_4__SCAN_IN), .A2(n4508), .ZN(U3318) );
  INV_X1 U5075 ( .A(D_REG_3__SCAN_IN), .ZN(n4674) );
  NOR2_X1 U5076 ( .A1(n4509), .A2(n4674), .ZN(U3319) );
  INV_X1 U5077 ( .A(D_REG_2__SCAN_IN), .ZN(n4772) );
  NOR2_X1 U5078 ( .A1(n4509), .A2(n4772), .ZN(U3320) );
  OAI21_X1 U5079 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4510), .ZN(
        n4511) );
  INV_X1 U5080 ( .A(n4511), .ZN(U3329) );
  INV_X1 U5081 ( .A(DATAI_18_), .ZN(n4512) );
  AOI22_X1 U5082 ( .A1(STATE_REG_SCAN_IN), .A2(n4513), .B1(n4512), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U5083 ( .A(DATAI_16_), .ZN(n4514) );
  AOI22_X1 U5084 ( .A1(STATE_REG_SCAN_IN), .A2(n4515), .B1(n4514), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5085 ( .A(DATAI_15_), .ZN(n4714) );
  AOI22_X1 U5086 ( .A1(STATE_REG_SCAN_IN), .A2(n4516), .B1(n4714), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5087 ( .A(DATAI_14_), .ZN(n4703) );
  AOI22_X1 U5088 ( .A1(STATE_REG_SCAN_IN), .A2(n2208), .B1(n4703), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U5089 ( .A1(STATE_REG_SCAN_IN), .A2(n4517), .B1(n2673), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5090 ( .A(DATAI_11_), .ZN(n4715) );
  AOI22_X1 U5091 ( .A1(STATE_REG_SCAN_IN), .A2(n4518), .B1(n4715), .B2(U3149), 
        .ZN(U3341) );
  OAI22_X1 U5092 ( .A1(U3149), .A2(n4519), .B1(DATAI_10_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4520) );
  INV_X1 U5093 ( .A(n4520), .ZN(U3342) );
  INV_X1 U5094 ( .A(DATAI_9_), .ZN(n4702) );
  AOI22_X1 U5095 ( .A1(STATE_REG_SCAN_IN), .A2(n4521), .B1(n4702), .B2(U3149), 
        .ZN(U3343) );
  INV_X1 U5096 ( .A(DATAI_8_), .ZN(n4712) );
  AOI22_X1 U5097 ( .A1(STATE_REG_SCAN_IN), .A2(n4522), .B1(n4712), .B2(U3149), 
        .ZN(U3344) );
  INV_X1 U5098 ( .A(DATAI_7_), .ZN(n4523) );
  AOI22_X1 U5099 ( .A1(STATE_REG_SCAN_IN), .A2(n4524), .B1(n4523), .B2(U3149), 
        .ZN(U3345) );
  OAI22_X1 U5100 ( .A1(U3149), .A2(n4525), .B1(DATAI_6_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4526) );
  INV_X1 U5101 ( .A(n4526), .ZN(U3346) );
  INV_X1 U5102 ( .A(DATAI_5_), .ZN(n4527) );
  AOI22_X1 U5103 ( .A1(STATE_REG_SCAN_IN), .A2(n4528), .B1(n4527), .B2(U3149), 
        .ZN(U3347) );
  AOI211_X1 U5104 ( .C1(n4583), .C2(n4531), .A(n4530), .B(n4529), .ZN(n4587)
         );
  INV_X1 U5105 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4532) );
  AOI22_X1 U5106 ( .A1(n4585), .A2(n4587), .B1(n4532), .B2(n4584), .ZN(U3467)
         );
  AOI21_X1 U5107 ( .B1(n4583), .B2(n4534), .A(n4533), .ZN(n4591) );
  AOI22_X1 U5108 ( .A1(n4535), .A2(n4588), .B1(REG0_REG_1__SCAN_IN), .B2(n4584), .ZN(n4536) );
  OAI21_X1 U5109 ( .B1(n4591), .B2(n4584), .A(n4536), .ZN(U3469) );
  AND3_X1 U5110 ( .A1(n4538), .A2(n4570), .A3(n4537), .ZN(n4540) );
  AOI211_X1 U5111 ( .C1(n4583), .C2(n4541), .A(n4540), .B(n4539), .ZN(n4592)
         );
  INV_X1 U5112 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4542) );
  AOI22_X1 U5113 ( .A1(n4585), .A2(n4592), .B1(n4542), .B2(n4584), .ZN(U3471)
         );
  NOR2_X1 U5114 ( .A1(n4543), .A2(n4577), .ZN(n4546) );
  INV_X1 U5115 ( .A(n4544), .ZN(n4545) );
  AOI211_X1 U5116 ( .C1(n4583), .C2(n4547), .A(n4546), .B(n4545), .ZN(n4593)
         );
  INV_X1 U5117 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4733) );
  AOI22_X1 U5118 ( .A1(n4585), .A2(n4593), .B1(n4733), .B2(n4584), .ZN(U3473)
         );
  NAND2_X1 U5119 ( .A1(n4548), .A2(n4583), .ZN(n4550) );
  NAND2_X1 U5120 ( .A1(n4550), .A2(n4549), .ZN(n4551) );
  NOR2_X1 U5121 ( .A1(n4552), .A2(n4551), .ZN(n4594) );
  INV_X1 U5122 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4729) );
  AOI22_X1 U5123 ( .A1(n4585), .A2(n4594), .B1(n4729), .B2(n4584), .ZN(U3475)
         );
  NOR3_X1 U5124 ( .A1(n4554), .A2(n4553), .A3(n4577), .ZN(n4556) );
  AOI211_X1 U5125 ( .C1(n4583), .C2(n4557), .A(n4556), .B(n4555), .ZN(n4595)
         );
  INV_X1 U5126 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4558) );
  AOI22_X1 U5127 ( .A1(n4585), .A2(n4595), .B1(n4558), .B2(n4584), .ZN(U3479)
         );
  AOI211_X1 U5128 ( .C1(n4562), .C2(n4561), .A(n4560), .B(n4559), .ZN(n4597)
         );
  INV_X1 U5129 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4563) );
  AOI22_X1 U5130 ( .A1(n4585), .A2(n4597), .B1(n4563), .B2(n4584), .ZN(U3481)
         );
  NOR3_X1 U5131 ( .A1(n4565), .A2(n4564), .A3(n4577), .ZN(n4567) );
  AOI211_X1 U5132 ( .C1(n4568), .C2(n4583), .A(n4567), .B(n4566), .ZN(n4599)
         );
  INV_X1 U5133 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4569) );
  AOI22_X1 U5134 ( .A1(n4585), .A2(n4599), .B1(n4569), .B2(n4584), .ZN(U3483)
         );
  AND3_X1 U5135 ( .A1(n4572), .A2(n4571), .A3(n4570), .ZN(n4573) );
  AOI21_X1 U5136 ( .B1(n4574), .B2(n4583), .A(n4573), .ZN(n4575) );
  INV_X1 U5137 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4732) );
  AOI22_X1 U5138 ( .A1(n4585), .A2(n4600), .B1(n4732), .B2(n4584), .ZN(U3487)
         );
  NOR2_X1 U5139 ( .A1(n4578), .A2(n4577), .ZN(n4581) );
  INV_X1 U5140 ( .A(n4579), .ZN(n4580) );
  AOI211_X1 U5141 ( .C1(n4583), .C2(n4582), .A(n4581), .B(n4580), .ZN(n4603)
         );
  INV_X1 U5142 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4747) );
  AOI22_X1 U5143 ( .A1(n4585), .A2(n4603), .B1(n4747), .B2(n4584), .ZN(U3489)
         );
  AOI22_X1 U5144 ( .A1(n4604), .A2(n4587), .B1(n4586), .B2(n4601), .ZN(U3518)
         );
  AOI22_X1 U5145 ( .A1(n4589), .A2(n4588), .B1(REG1_REG_1__SCAN_IN), .B2(n4601), .ZN(n4590) );
  OAI21_X1 U5146 ( .B1(n4591), .B2(n4601), .A(n4590), .ZN(U3519) );
  AOI22_X1 U5147 ( .A1(n4604), .A2(n4592), .B1(n4850), .B2(n4601), .ZN(U3520)
         );
  INV_X1 U5148 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4789) );
  AOI22_X1 U5149 ( .A1(n4604), .A2(n4593), .B1(n4789), .B2(n4601), .ZN(U3521)
         );
  INV_X1 U5150 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4826) );
  AOI22_X1 U5151 ( .A1(n4604), .A2(n4594), .B1(n4826), .B2(n4601), .ZN(U3522)
         );
  AOI22_X1 U5152 ( .A1(n4604), .A2(n4595), .B1(n4868), .B2(n4601), .ZN(U3524)
         );
  AOI22_X1 U5153 ( .A1(n4604), .A2(n4597), .B1(n4596), .B2(n4601), .ZN(U3525)
         );
  INV_X1 U5154 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4598) );
  AOI22_X1 U5155 ( .A1(n4604), .A2(n4599), .B1(n4598), .B2(n4601), .ZN(U3526)
         );
  INV_X1 U5156 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4762) );
  AOI22_X1 U5157 ( .A1(n4604), .A2(n4600), .B1(n4762), .B2(n4601), .ZN(U3528)
         );
  AOI22_X1 U5158 ( .A1(n4604), .A2(n4603), .B1(n4602), .B2(n4601), .ZN(U3529)
         );
  NOR4_X1 U5159 ( .A1(keyinput16), .A2(keyinput67), .A3(keyinput78), .A4(
        keyinput38), .ZN(n4632) );
  NAND2_X1 U5160 ( .A1(keyinput5), .A2(keyinput49), .ZN(n4605) );
  NOR3_X1 U5161 ( .A1(keyinput36), .A2(keyinput109), .A3(n4605), .ZN(n4631) );
  NAND2_X1 U5162 ( .A1(keyinput43), .A2(keyinput0), .ZN(n4606) );
  NOR3_X1 U5163 ( .A1(keyinput84), .A2(keyinput64), .A3(n4606), .ZN(n4607) );
  NAND3_X1 U5164 ( .A1(keyinput17), .A2(keyinput114), .A3(n4607), .ZN(n4616)
         );
  NAND3_X1 U5165 ( .A1(keyinput69), .A2(keyinput122), .A3(keyinput39), .ZN(
        n4608) );
  NOR2_X1 U5166 ( .A1(keyinput24), .A2(n4608), .ZN(n4614) );
  NAND2_X1 U5167 ( .A1(keyinput46), .A2(keyinput106), .ZN(n4609) );
  NOR3_X1 U5168 ( .A1(keyinput52), .A2(keyinput51), .A3(n4609), .ZN(n4613) );
  NOR4_X1 U5169 ( .A1(keyinput104), .A2(keyinput100), .A3(keyinput80), .A4(
        keyinput88), .ZN(n4612) );
  INV_X1 U5170 ( .A(keyinput112), .ZN(n4610) );
  NOR4_X1 U5171 ( .A1(keyinput93), .A2(keyinput119), .A3(keyinput118), .A4(
        n4610), .ZN(n4611) );
  NAND4_X1 U5172 ( .A1(n4614), .A2(n4613), .A3(n4612), .A4(n4611), .ZN(n4615)
         );
  NOR4_X1 U5173 ( .A1(keyinput20), .A2(keyinput53), .A3(n4616), .A4(n4615), 
        .ZN(n4630) );
  NAND4_X1 U5174 ( .A1(keyinput31), .A2(keyinput30), .A3(keyinput42), .A4(
        keyinput66), .ZN(n4628) );
  NAND4_X1 U5175 ( .A1(keyinput89), .A2(keyinput27), .A3(keyinput11), .A4(
        keyinput14), .ZN(n4627) );
  NAND4_X1 U5176 ( .A1(keyinput113), .A2(keyinput117), .A3(keyinput21), .A4(
        keyinput9), .ZN(n4617) );
  NOR3_X1 U5177 ( .A1(keyinput81), .A2(keyinput65), .A3(n4617), .ZN(n4618) );
  NAND3_X1 U5178 ( .A1(keyinput82), .A2(keyinput70), .A3(n4618), .ZN(n4626) );
  NOR4_X1 U5179 ( .A1(keyinput45), .A2(keyinput76), .A3(keyinput72), .A4(
        keyinput4), .ZN(n4624) );
  NAND2_X1 U5180 ( .A1(keyinput8), .A2(keyinput13), .ZN(n4619) );
  NOR3_X1 U5181 ( .A1(keyinput57), .A2(keyinput32), .A3(n4619), .ZN(n4623) );
  NAND2_X1 U5182 ( .A1(keyinput91), .A2(keyinput47), .ZN(n4620) );
  NOR3_X1 U5183 ( .A1(keyinput87), .A2(keyinput59), .A3(n4620), .ZN(n4622) );
  NOR4_X1 U5184 ( .A1(keyinput40), .A2(keyinput2), .A3(keyinput7), .A4(
        keyinput18), .ZN(n4621) );
  NAND4_X1 U5185 ( .A1(n4624), .A2(n4623), .A3(n4622), .A4(n4621), .ZN(n4625)
         );
  NOR4_X1 U5186 ( .A1(n4628), .A2(n4627), .A3(n4626), .A4(n4625), .ZN(n4629)
         );
  NAND4_X1 U5187 ( .A1(n4632), .A2(n4631), .A3(n4630), .A4(n4629), .ZN(n4666)
         );
  NOR2_X1 U5188 ( .A1(keyinput127), .A2(keyinput85), .ZN(n4633) );
  NAND3_X1 U5189 ( .A1(keyinput26), .A2(keyinput28), .A3(n4633), .ZN(n4634) );
  NOR4_X1 U5190 ( .A1(keyinput99), .A2(keyinput75), .A3(keyinput73), .A4(n4634), .ZN(n4664) );
  NAND2_X1 U5191 ( .A1(keyinput33), .A2(keyinput101), .ZN(n4635) );
  NOR3_X1 U5192 ( .A1(keyinput6), .A2(keyinput48), .A3(n4635), .ZN(n4637) );
  INV_X1 U5193 ( .A(keyinput35), .ZN(n4636) );
  NAND3_X1 U5194 ( .A1(keyinput3), .A2(n4637), .A3(n4636), .ZN(n4645) );
  NAND2_X1 U5195 ( .A1(keyinput107), .A2(keyinput125), .ZN(n4638) );
  NOR3_X1 U5196 ( .A1(keyinput74), .A2(keyinput29), .A3(n4638), .ZN(n4643) );
  NOR4_X1 U5197 ( .A1(keyinput19), .A2(keyinput50), .A3(keyinput102), .A4(
        keyinput10), .ZN(n4642) );
  NAND2_X1 U5198 ( .A1(keyinput34), .A2(keyinput126), .ZN(n4639) );
  NOR3_X1 U5199 ( .A1(keyinput98), .A2(keyinput77), .A3(n4639), .ZN(n4641) );
  INV_X1 U5200 ( .A(keyinput120), .ZN(n4823) );
  NOR4_X1 U5201 ( .A1(keyinput111), .A2(keyinput54), .A3(keyinput55), .A4(
        n4823), .ZN(n4640) );
  NAND4_X1 U5202 ( .A1(n4643), .A2(n4642), .A3(n4641), .A4(n4640), .ZN(n4644)
         );
  NOR4_X1 U5203 ( .A1(keyinput23), .A2(keyinput90), .A3(n4645), .A4(n4644), 
        .ZN(n4663) );
  NOR2_X1 U5204 ( .A1(keyinput103), .A2(keyinput1), .ZN(n4646) );
  NAND3_X1 U5205 ( .A1(keyinput22), .A2(keyinput79), .A3(n4646), .ZN(n4652) );
  INV_X1 U5206 ( .A(keyinput61), .ZN(n4647) );
  NAND4_X1 U5207 ( .A1(keyinput123), .A2(keyinput60), .A3(keyinput121), .A4(
        n4647), .ZN(n4651) );
  NOR2_X1 U5208 ( .A1(keyinput62), .A2(keyinput97), .ZN(n4648) );
  NAND3_X1 U5209 ( .A1(keyinput83), .A2(keyinput94), .A3(n4648), .ZN(n4650) );
  NAND4_X1 U5210 ( .A1(keyinput108), .A2(keyinput96), .A3(keyinput41), .A4(
        keyinput44), .ZN(n4649) );
  NOR4_X1 U5211 ( .A1(n4652), .A2(n4651), .A3(n4650), .A4(n4649), .ZN(n4662)
         );
  NOR2_X1 U5212 ( .A1(keyinput37), .A2(keyinput56), .ZN(n4653) );
  NAND3_X1 U5213 ( .A1(keyinput25), .A2(keyinput71), .A3(n4653), .ZN(n4660) );
  NOR3_X1 U5214 ( .A1(keyinput95), .A2(keyinput58), .A3(keyinput63), .ZN(n4654) );
  NAND2_X1 U5215 ( .A1(keyinput92), .A2(n4654), .ZN(n4659) );
  NOR2_X1 U5216 ( .A1(keyinput12), .A2(keyinput116), .ZN(n4655) );
  NAND3_X1 U5217 ( .A1(keyinput105), .A2(keyinput86), .A3(n4655), .ZN(n4658)
         );
  NOR2_X1 U5218 ( .A1(keyinput68), .A2(keyinput124), .ZN(n4656) );
  NAND3_X1 U5219 ( .A1(keyinput115), .A2(keyinput15), .A3(n4656), .ZN(n4657)
         );
  NOR4_X1 U5220 ( .A1(n4660), .A2(n4659), .A3(n4658), .A4(n4657), .ZN(n4661)
         );
  NAND4_X1 U5221 ( .A1(n4664), .A2(n4663), .A3(n4662), .A4(n4661), .ZN(n4665)
         );
  OAI21_X1 U5222 ( .B1(n4666), .B2(n4665), .A(keyinput110), .ZN(n4921) );
  AOI22_X1 U5223 ( .A1(n4669), .A2(keyinput27), .B1(keyinput11), .B2(n4668), 
        .ZN(n4667) );
  OAI221_X1 U5224 ( .B1(n4669), .B2(keyinput27), .C1(n4668), .C2(keyinput11), 
        .A(n4667), .ZN(n4682) );
  AOI22_X1 U5225 ( .A1(n4672), .A2(keyinput14), .B1(keyinput31), .B2(n4671), 
        .ZN(n4670) );
  OAI221_X1 U5226 ( .B1(n4672), .B2(keyinput14), .C1(n4671), .C2(keyinput31), 
        .A(n4670), .ZN(n4681) );
  AOI22_X1 U5227 ( .A1(n4675), .A2(keyinput30), .B1(keyinput42), .B2(n4674), 
        .ZN(n4673) );
  OAI221_X1 U5228 ( .B1(n4675), .B2(keyinput30), .C1(n4674), .C2(keyinput42), 
        .A(n4673), .ZN(n4680) );
  AOI22_X1 U5229 ( .A1(n4678), .A2(keyinput66), .B1(keyinput82), .B2(n4677), 
        .ZN(n4676) );
  OAI221_X1 U5230 ( .B1(n4678), .B2(keyinput66), .C1(n4677), .C2(keyinput82), 
        .A(n4676), .ZN(n4679) );
  NOR4_X1 U5231 ( .A1(n4682), .A2(n4681), .A3(n4680), .A4(n4679), .ZN(n4726)
         );
  XOR2_X1 U5232 ( .A(n4683), .B(keyinput21), .Z(n4688) );
  XOR2_X1 U5233 ( .A(n4684), .B(keyinput81), .Z(n4687) );
  XOR2_X1 U5234 ( .A(n2673), .B(keyinput113), .Z(n4686) );
  XNOR2_X1 U5235 ( .A(IR_REG_30__SCAN_IN), .B(keyinput13), .ZN(n4685) );
  NAND4_X1 U5236 ( .A1(n4688), .A2(n4687), .A3(n4686), .A4(n4685), .ZN(n4694)
         );
  XNOR2_X1 U5237 ( .A(IR_REG_4__SCAN_IN), .B(keyinput65), .ZN(n4692) );
  XNOR2_X1 U5238 ( .A(IR_REG_19__SCAN_IN), .B(keyinput70), .ZN(n4691) );
  XNOR2_X1 U5239 ( .A(REG3_REG_13__SCAN_IN), .B(keyinput9), .ZN(n4690) );
  XNOR2_X1 U5240 ( .A(IR_REG_20__SCAN_IN), .B(keyinput117), .ZN(n4689) );
  NAND4_X1 U5241 ( .A1(n4692), .A2(n4691), .A3(n4690), .A4(n4689), .ZN(n4693)
         );
  NOR2_X1 U5242 ( .A1(n4694), .A2(n4693), .ZN(n4725) );
  INV_X1 U5243 ( .A(DATAI_2_), .ZN(n4696) );
  AOI22_X1 U5244 ( .A1(n4696), .A2(keyinput4), .B1(n2739), .B2(keyinput8), 
        .ZN(n4695) );
  OAI221_X1 U5245 ( .B1(n4696), .B2(keyinput4), .C1(n2739), .C2(keyinput8), 
        .A(n4695), .ZN(n4709) );
  INV_X1 U5246 ( .A(B_REG_SCAN_IN), .ZN(n4698) );
  AOI22_X1 U5247 ( .A1(n4699), .A2(keyinput76), .B1(n4698), .B2(keyinput72), 
        .ZN(n4697) );
  OAI221_X1 U5248 ( .B1(n4699), .B2(keyinput76), .C1(n4698), .C2(keyinput72), 
        .A(n4697), .ZN(n4708) );
  AOI22_X1 U5249 ( .A1(n4702), .A2(keyinput32), .B1(n4701), .B2(keyinput40), 
        .ZN(n4700) );
  OAI221_X1 U5250 ( .B1(n4702), .B2(keyinput32), .C1(n4701), .C2(keyinput40), 
        .A(n4700), .ZN(n4707) );
  XOR2_X1 U5251 ( .A(n4703), .B(keyinput57), .Z(n4705) );
  XNOR2_X1 U5252 ( .A(IR_REG_26__SCAN_IN), .B(keyinput45), .ZN(n4704) );
  NAND2_X1 U5253 ( .A1(n4705), .A2(n4704), .ZN(n4706) );
  NOR4_X1 U5254 ( .A1(n4709), .A2(n4708), .A3(n4707), .A4(n4706), .ZN(n4724)
         );
  AOI22_X1 U5255 ( .A1(n4712), .A2(keyinput18), .B1(n4711), .B2(keyinput47), 
        .ZN(n4710) );
  OAI221_X1 U5256 ( .B1(n4712), .B2(keyinput18), .C1(n4711), .C2(keyinput47), 
        .A(n4710), .ZN(n4722) );
  AOI22_X1 U5257 ( .A1(n4715), .A2(keyinput59), .B1(keyinput87), .B2(n4714), 
        .ZN(n4713) );
  OAI221_X1 U5258 ( .B1(n4715), .B2(keyinput59), .C1(n4714), .C2(keyinput87), 
        .A(n4713), .ZN(n4721) );
  XNOR2_X1 U5259 ( .A(IR_REG_17__SCAN_IN), .B(keyinput2), .ZN(n4719) );
  XNOR2_X1 U5260 ( .A(IR_REG_21__SCAN_IN), .B(keyinput7), .ZN(n4718) );
  XNOR2_X1 U5261 ( .A(IR_REG_13__SCAN_IN), .B(keyinput99), .ZN(n4717) );
  XNOR2_X1 U5262 ( .A(DATAI_19_), .B(keyinput91), .ZN(n4716) );
  NAND4_X1 U5263 ( .A1(n4719), .A2(n4718), .A3(n4717), .A4(n4716), .ZN(n4720)
         );
  NOR3_X1 U5264 ( .A1(n4722), .A2(n4721), .A3(n4720), .ZN(n4723) );
  NAND4_X1 U5265 ( .A1(n4726), .A2(n4725), .A3(n4724), .A4(n4723), .ZN(n4920)
         );
  AOI22_X1 U5266 ( .A1(n4729), .A2(keyinput67), .B1(n4728), .B2(keyinput78), 
        .ZN(n4727) );
  OAI221_X1 U5267 ( .B1(n4729), .B2(keyinput67), .C1(n4728), .C2(keyinput78), 
        .A(n4727), .ZN(n4740) );
  AOI22_X1 U5268 ( .A1(n4732), .A2(keyinput109), .B1(n4731), .B2(keyinput36), 
        .ZN(n4730) );
  OAI221_X1 U5269 ( .B1(n4732), .B2(keyinput109), .C1(n4731), .C2(keyinput36), 
        .A(n4730), .ZN(n4739) );
  XOR2_X1 U5270 ( .A(n4733), .B(keyinput16), .Z(n4737) );
  XNOR2_X1 U5271 ( .A(keyinput38), .B(DATAI_4_), .ZN(n4736) );
  XNOR2_X1 U5272 ( .A(DATAI_0_), .B(keyinput5), .ZN(n4735) );
  XNOR2_X1 U5273 ( .A(IR_REG_3__SCAN_IN), .B(keyinput52), .ZN(n4734) );
  NAND4_X1 U5274 ( .A1(n4737), .A2(n4736), .A3(n4735), .A4(n4734), .ZN(n4738)
         );
  NOR3_X1 U5275 ( .A1(n4740), .A2(n4739), .A3(n4738), .ZN(n4918) );
  AOI22_X1 U5276 ( .A1(n4743), .A2(keyinput24), .B1(keyinput93), .B2(n4742), 
        .ZN(n4741) );
  OAI221_X1 U5277 ( .B1(n4743), .B2(keyinput24), .C1(n4742), .C2(keyinput93), 
        .A(n4741), .ZN(n4754) );
  INV_X1 U5278 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4745) );
  AOI22_X1 U5279 ( .A1(n4745), .A2(keyinput46), .B1(keyinput122), .B2(n4168), 
        .ZN(n4744) );
  OAI221_X1 U5280 ( .B1(n4745), .B2(keyinput46), .C1(n4168), .C2(keyinput122), 
        .A(n4744), .ZN(n4753) );
  INV_X1 U5281 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4748) );
  AOI22_X1 U5282 ( .A1(n4748), .A2(keyinput106), .B1(n4747), .B2(keyinput51), 
        .ZN(n4746) );
  OAI221_X1 U5283 ( .B1(n4748), .B2(keyinput106), .C1(n4747), .C2(keyinput51), 
        .A(n4746), .ZN(n4752) );
  XNOR2_X1 U5284 ( .A(REG0_REG_16__SCAN_IN), .B(keyinput39), .ZN(n4750) );
  XNOR2_X1 U5285 ( .A(IR_REG_27__SCAN_IN), .B(keyinput69), .ZN(n4749) );
  NAND2_X1 U5286 ( .A1(n4750), .A2(n4749), .ZN(n4751) );
  NOR4_X1 U5287 ( .A1(n4754), .A2(n4753), .A3(n4752), .A4(n4751), .ZN(n4917)
         );
  INV_X1 U5288 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4757) );
  INV_X1 U5289 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4756) );
  AOI22_X1 U5290 ( .A1(n4757), .A2(keyinput0), .B1(n4756), .B2(keyinput20), 
        .ZN(n4755) );
  OAI221_X1 U5291 ( .B1(n4757), .B2(keyinput0), .C1(n4756), .C2(keyinput20), 
        .A(n4755), .ZN(n4787) );
  INV_X1 U5292 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4759) );
  AOI22_X1 U5293 ( .A1(n4760), .A2(keyinput114), .B1(keyinput64), .B2(n4759), 
        .ZN(n4758) );
  OAI221_X1 U5294 ( .B1(n4760), .B2(keyinput114), .C1(n4759), .C2(keyinput64), 
        .A(n4758), .ZN(n4786) );
  OAI22_X1 U5295 ( .A1(n4763), .A2(keyinput43), .B1(n4762), .B2(keyinput49), 
        .ZN(n4761) );
  AOI221_X1 U5296 ( .B1(n4763), .B2(keyinput43), .C1(keyinput49), .C2(n4762), 
        .A(n4761), .ZN(n4767) );
  XNOR2_X1 U5297 ( .A(DATAO_REG_29__SCAN_IN), .B(keyinput53), .ZN(n4766) );
  XOR2_X1 U5298 ( .A(keyinput17), .B(n4764), .Z(n4765) );
  NAND3_X1 U5299 ( .A1(n4767), .A2(n4766), .A3(n4765), .ZN(n4785) );
  OAI22_X1 U5300 ( .A1(n4770), .A2(keyinput119), .B1(n4769), .B2(keyinput118), 
        .ZN(n4768) );
  AOI221_X1 U5301 ( .B1(n4770), .B2(keyinput119), .C1(keyinput118), .C2(n4769), 
        .A(n4768), .ZN(n4783) );
  OAI22_X1 U5302 ( .A1(n4773), .A2(keyinput112), .B1(n4772), .B2(keyinput104), 
        .ZN(n4771) );
  AOI221_X1 U5303 ( .B1(n4773), .B2(keyinput112), .C1(keyinput104), .C2(n4772), 
        .A(n4771), .ZN(n4782) );
  OAI22_X1 U5304 ( .A1(n4776), .A2(keyinput100), .B1(n4775), .B2(keyinput80), 
        .ZN(n4774) );
  AOI221_X1 U5305 ( .B1(n4776), .B2(keyinput100), .C1(keyinput80), .C2(n4775), 
        .A(n4774), .ZN(n4781) );
  OAI22_X1 U5306 ( .A1(n4779), .A2(keyinput88), .B1(n4778), .B2(keyinput89), 
        .ZN(n4777) );
  AOI221_X1 U5307 ( .B1(n4779), .B2(keyinput88), .C1(keyinput89), .C2(n4778), 
        .A(n4777), .ZN(n4780) );
  NAND4_X1 U5308 ( .A1(n4783), .A2(n4782), .A3(n4781), .A4(n4780), .ZN(n4784)
         );
  NOR4_X1 U5309 ( .A1(n4787), .A2(n4786), .A3(n4785), .A4(n4784), .ZN(n4916)
         );
  XOR2_X1 U5310 ( .A(keyinput75), .B(ADDR_REG_3__SCAN_IN), .Z(n4792) );
  AOI22_X1 U5311 ( .A1(n4790), .A2(keyinput127), .B1(keyinput26), .B2(n4789), 
        .ZN(n4788) );
  OAI221_X1 U5312 ( .B1(n4790), .B2(keyinput127), .C1(n4789), .C2(keyinput26), 
        .A(n4788), .ZN(n4791) );
  AOI211_X1 U5313 ( .C1(keyinput110), .C2(n4793), .A(n4792), .B(n4791), .ZN(
        n4819) );
  INV_X1 U5314 ( .A(keyinput28), .ZN(n4796) );
  INV_X1 U5315 ( .A(keyinput19), .ZN(n4795) );
  OAI22_X1 U5316 ( .A1(n4796), .A2(DATAO_REG_6__SCAN_IN), .B1(n4795), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n4794) );
  AOI221_X1 U5317 ( .B1(n4796), .B2(DATAO_REG_6__SCAN_IN), .C1(
        DATAO_REG_1__SCAN_IN), .C2(n4795), .A(n4794), .ZN(n4818) );
  INV_X1 U5318 ( .A(REG3_REG_0__SCAN_IN), .ZN(n4799) );
  INV_X1 U5319 ( .A(keyinput85), .ZN(n4798) );
  OAI22_X1 U5320 ( .A1(n4799), .A2(keyinput73), .B1(n4798), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n4797) );
  AOI221_X1 U5321 ( .B1(n4799), .B2(keyinput73), .C1(DATAO_REG_10__SCAN_IN), 
        .C2(n4798), .A(n4797), .ZN(n4817) );
  INV_X1 U5322 ( .A(keyinput29), .ZN(n4802) );
  INV_X1 U5323 ( .A(keyinput102), .ZN(n4801) );
  AOI22_X1 U5324 ( .A1(n4802), .A2(DATAO_REG_15__SCAN_IN), .B1(
        DATAO_REG_14__SCAN_IN), .B2(n4801), .ZN(n4800) );
  OAI221_X1 U5325 ( .B1(n4802), .B2(DATAO_REG_15__SCAN_IN), .C1(n4801), .C2(
        DATAO_REG_14__SCAN_IN), .A(n4800), .ZN(n4815) );
  INV_X1 U5326 ( .A(keyinput50), .ZN(n4805) );
  INV_X1 U5327 ( .A(keyinput125), .ZN(n4804) );
  AOI22_X1 U5328 ( .A1(n4805), .A2(DATAO_REG_2__SCAN_IN), .B1(
        DATAO_REG_9__SCAN_IN), .B2(n4804), .ZN(n4803) );
  OAI221_X1 U5329 ( .B1(n4805), .B2(DATAO_REG_2__SCAN_IN), .C1(n4804), .C2(
        DATAO_REG_9__SCAN_IN), .A(n4803), .ZN(n4814) );
  AOI22_X1 U5330 ( .A1(n4808), .A2(keyinput107), .B1(n4807), .B2(keyinput23), 
        .ZN(n4806) );
  OAI221_X1 U5331 ( .B1(n4808), .B2(keyinput107), .C1(n4807), .C2(keyinput23), 
        .A(n4806), .ZN(n4813) );
  INV_X1 U5332 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4811) );
  AOI22_X1 U5333 ( .A1(n4811), .A2(keyinput10), .B1(keyinput74), .B2(n4810), 
        .ZN(n4809) );
  OAI221_X1 U5334 ( .B1(n4811), .B2(keyinput10), .C1(n4810), .C2(keyinput74), 
        .A(n4809), .ZN(n4812) );
  NOR4_X1 U5335 ( .A1(n4815), .A2(n4814), .A3(n4813), .A4(n4812), .ZN(n4816)
         );
  NAND4_X1 U5336 ( .A1(n4819), .A2(n4818), .A3(n4817), .A4(n4816), .ZN(n4914)
         );
  INV_X1 U5337 ( .A(keyinput98), .ZN(n4821) );
  OAI22_X1 U5338 ( .A1(n2451), .A2(keyinput34), .B1(n4821), .B2(
        ADDR_REG_4__SCAN_IN), .ZN(n4820) );
  AOI221_X1 U5339 ( .B1(n2451), .B2(keyinput34), .C1(ADDR_REG_4__SCAN_IN), 
        .C2(n4821), .A(n4820), .ZN(n4832) );
  OAI22_X1 U5340 ( .A1(n3285), .A2(keyinput126), .B1(n4823), .B2(
        ADDR_REG_2__SCAN_IN), .ZN(n4822) );
  AOI221_X1 U5341 ( .B1(n3285), .B2(keyinput126), .C1(ADDR_REG_2__SCAN_IN), 
        .C2(n4823), .A(n4822), .ZN(n4831) );
  INV_X1 U5342 ( .A(keyinput77), .ZN(n4825) );
  OAI22_X1 U5343 ( .A1(n3259), .A2(keyinput95), .B1(n4825), .B2(
        ADDR_REG_5__SCAN_IN), .ZN(n4824) );
  AOI221_X1 U5344 ( .B1(n3259), .B2(keyinput95), .C1(ADDR_REG_5__SCAN_IN), 
        .C2(n4825), .A(n4824), .ZN(n4830) );
  XOR2_X1 U5345 ( .A(IR_REG_0__SCAN_IN), .B(keyinput54), .Z(n4828) );
  XNOR2_X1 U5346 ( .A(keyinput55), .B(n4826), .ZN(n4827) );
  NOR2_X1 U5347 ( .A1(n4828), .A2(n4827), .ZN(n4829) );
  NAND4_X1 U5348 ( .A1(n4832), .A2(n4831), .A3(n4830), .A4(n4829), .ZN(n4913)
         );
  INV_X1 U5349 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4834) );
  OAI22_X1 U5350 ( .A1(n4835), .A2(keyinput3), .B1(n4834), .B2(keyinput101), 
        .ZN(n4833) );
  AOI221_X1 U5351 ( .B1(n4835), .B2(keyinput3), .C1(keyinput101), .C2(n4834), 
        .A(n4833), .ZN(n4847) );
  INV_X1 U5352 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4837) );
  OAI22_X1 U5353 ( .A1(n4837), .A2(keyinput90), .B1(n3715), .B2(keyinput35), 
        .ZN(n4836) );
  AOI221_X1 U5354 ( .B1(n4837), .B2(keyinput90), .C1(keyinput35), .C2(n3715), 
        .A(n4836), .ZN(n4846) );
  INV_X1 U5355 ( .A(REG3_REG_1__SCAN_IN), .ZN(n4839) );
  OAI22_X1 U5356 ( .A1(n4840), .A2(keyinput48), .B1(n4839), .B2(keyinput111), 
        .ZN(n4838) );
  AOI221_X1 U5357 ( .B1(n4840), .B2(keyinput48), .C1(keyinput111), .C2(n4839), 
        .A(n4838), .ZN(n4845) );
  INV_X1 U5358 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4843) );
  INV_X1 U5359 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4842) );
  OAI22_X1 U5360 ( .A1(n4843), .A2(keyinput6), .B1(n4842), .B2(keyinput33), 
        .ZN(n4841) );
  AOI221_X1 U5361 ( .B1(n4843), .B2(keyinput6), .C1(keyinput33), .C2(n4842), 
        .A(n4841), .ZN(n4844) );
  NAND4_X1 U5362 ( .A1(n4847), .A2(n4846), .A3(n4845), .A4(n4844), .ZN(n4912)
         );
  AOI22_X1 U5363 ( .A1(n4850), .A2(keyinput105), .B1(n4849), .B2(keyinput116), 
        .ZN(n4848) );
  OAI221_X1 U5364 ( .B1(n4850), .B2(keyinput105), .C1(n4849), .C2(keyinput116), 
        .A(n4848), .ZN(n4862) );
  AOI22_X1 U5365 ( .A1(n2686), .A2(keyinput124), .B1(keyinput12), .B2(n4852), 
        .ZN(n4851) );
  OAI221_X1 U5366 ( .B1(n2686), .B2(keyinput124), .C1(n4852), .C2(keyinput12), 
        .A(n4851), .ZN(n4861) );
  INV_X1 U5367 ( .A(keyinput68), .ZN(n4854) );
  AOI22_X1 U5368 ( .A1(n4855), .A2(keyinput15), .B1(ADDR_REG_16__SCAN_IN), 
        .B2(n4854), .ZN(n4853) );
  OAI221_X1 U5369 ( .B1(n4855), .B2(keyinput15), .C1(n4854), .C2(
        ADDR_REG_16__SCAN_IN), .A(n4853), .ZN(n4860) );
  INV_X1 U5370 ( .A(keyinput86), .ZN(n4856) );
  XOR2_X1 U5371 ( .A(ADDR_REG_18__SCAN_IN), .B(n4856), .Z(n4858) );
  XNOR2_X1 U5372 ( .A(IR_REG_31__SCAN_IN), .B(keyinput123), .ZN(n4857) );
  NAND2_X1 U5373 ( .A1(n4858), .A2(n4857), .ZN(n4859) );
  NOR4_X1 U5374 ( .A1(n4862), .A2(n4861), .A3(n4860), .A4(n4859), .ZN(n4910)
         );
  INV_X1 U5375 ( .A(keyinput58), .ZN(n4865) );
  INV_X1 U5376 ( .A(keyinput25), .ZN(n4864) );
  AOI22_X1 U5377 ( .A1(n4865), .A2(ADDR_REG_7__SCAN_IN), .B1(
        ADDR_REG_8__SCAN_IN), .B2(n4864), .ZN(n4863) );
  OAI221_X1 U5378 ( .B1(n4865), .B2(ADDR_REG_7__SCAN_IN), .C1(n4864), .C2(
        ADDR_REG_8__SCAN_IN), .A(n4863), .ZN(n4878) );
  INV_X1 U5379 ( .A(keyinput92), .ZN(n4867) );
  AOI22_X1 U5380 ( .A1(n4868), .A2(keyinput63), .B1(ADDR_REG_6__SCAN_IN), .B2(
        n4867), .ZN(n4866) );
  OAI221_X1 U5381 ( .B1(n4868), .B2(keyinput63), .C1(n4867), .C2(
        ADDR_REG_6__SCAN_IN), .A(n4866), .ZN(n4877) );
  INV_X1 U5382 ( .A(keyinput71), .ZN(n4871) );
  INV_X1 U5383 ( .A(keyinput115), .ZN(n4870) );
  AOI22_X1 U5384 ( .A1(n4871), .A2(ADDR_REG_13__SCAN_IN), .B1(
        ADDR_REG_14__SCAN_IN), .B2(n4870), .ZN(n4869) );
  OAI221_X1 U5385 ( .B1(n4871), .B2(ADDR_REG_13__SCAN_IN), .C1(n4870), .C2(
        ADDR_REG_14__SCAN_IN), .A(n4869), .ZN(n4876) );
  INV_X1 U5386 ( .A(keyinput56), .ZN(n4874) );
  INV_X1 U5387 ( .A(keyinput37), .ZN(n4873) );
  AOI22_X1 U5388 ( .A1(n4874), .A2(ADDR_REG_9__SCAN_IN), .B1(
        ADDR_REG_11__SCAN_IN), .B2(n4873), .ZN(n4872) );
  OAI221_X1 U5389 ( .B1(n4874), .B2(ADDR_REG_9__SCAN_IN), .C1(n4873), .C2(
        ADDR_REG_11__SCAN_IN), .A(n4872), .ZN(n4875) );
  NOR4_X1 U5390 ( .A1(n4878), .A2(n4877), .A3(n4876), .A4(n4875), .ZN(n4909)
         );
  INV_X1 U5391 ( .A(keyinput62), .ZN(n4880) );
  AOI22_X1 U5392 ( .A1(n4283), .A2(keyinput97), .B1(DATAO_REG_24__SCAN_IN), 
        .B2(n4880), .ZN(n4879) );
  OAI221_X1 U5393 ( .B1(n4283), .B2(keyinput97), .C1(n4880), .C2(
        DATAO_REG_24__SCAN_IN), .A(n4879), .ZN(n4891) );
  INV_X1 U5394 ( .A(keyinput96), .ZN(n4882) );
  AOI22_X1 U5395 ( .A1(n4209), .A2(keyinput83), .B1(DATAO_REG_23__SCAN_IN), 
        .B2(n4882), .ZN(n4881) );
  OAI221_X1 U5396 ( .B1(n4209), .B2(keyinput83), .C1(n4882), .C2(
        DATAO_REG_23__SCAN_IN), .A(n4881), .ZN(n4890) );
  INV_X1 U5397 ( .A(keyinput44), .ZN(n4884) );
  AOI22_X1 U5398 ( .A1(n4276), .A2(keyinput84), .B1(DATAO_REG_25__SCAN_IN), 
        .B2(n4884), .ZN(n4883) );
  OAI221_X1 U5399 ( .B1(n4276), .B2(keyinput84), .C1(n4884), .C2(
        DATAO_REG_25__SCAN_IN), .A(n4883), .ZN(n4889) );
  AOI22_X1 U5400 ( .A1(n4887), .A2(keyinput94), .B1(n4886), .B2(keyinput41), 
        .ZN(n4885) );
  OAI221_X1 U5401 ( .B1(n4887), .B2(keyinput94), .C1(n4886), .C2(keyinput41), 
        .A(n4885), .ZN(n4888) );
  NOR4_X1 U5402 ( .A1(n4891), .A2(n4890), .A3(n4889), .A4(n4888), .ZN(n4908)
         );
  INV_X1 U5403 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4894) );
  INV_X1 U5404 ( .A(keyinput103), .ZN(n4893) );
  AOI22_X1 U5405 ( .A1(n4894), .A2(keyinput121), .B1(DATAO_REG_20__SCAN_IN), 
        .B2(n4893), .ZN(n4892) );
  OAI221_X1 U5406 ( .B1(n4894), .B2(keyinput121), .C1(n4893), .C2(
        DATAO_REG_20__SCAN_IN), .A(n4892), .ZN(n4906) );
  INV_X1 U5407 ( .A(keyinput60), .ZN(n4896) );
  AOI22_X1 U5408 ( .A1(n3057), .A2(keyinput61), .B1(DATAO_REG_16__SCAN_IN), 
        .B2(n4896), .ZN(n4895) );
  OAI221_X1 U5409 ( .B1(n3057), .B2(keyinput61), .C1(n4896), .C2(
        DATAO_REG_16__SCAN_IN), .A(n4895), .ZN(n4905) );
  INV_X1 U5410 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4899) );
  INV_X1 U5411 ( .A(keyinput1), .ZN(n4898) );
  AOI22_X1 U5412 ( .A1(n4899), .A2(keyinput108), .B1(DATAO_REG_22__SCAN_IN), 
        .B2(n4898), .ZN(n4897) );
  OAI221_X1 U5413 ( .B1(n4899), .B2(keyinput108), .C1(n4898), .C2(
        DATAO_REG_22__SCAN_IN), .A(n4897), .ZN(n4904) );
  INV_X1 U5414 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4902) );
  INV_X1 U5415 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4901) );
  AOI22_X1 U5416 ( .A1(n4902), .A2(keyinput22), .B1(n4901), .B2(keyinput79), 
        .ZN(n4900) );
  OAI221_X1 U5417 ( .B1(n4902), .B2(keyinput22), .C1(n4901), .C2(keyinput79), 
        .A(n4900), .ZN(n4903) );
  NOR4_X1 U5418 ( .A1(n4906), .A2(n4905), .A3(n4904), .A4(n4903), .ZN(n4907)
         );
  NAND4_X1 U5419 ( .A1(n4910), .A2(n4909), .A3(n4908), .A4(n4907), .ZN(n4911)
         );
  NOR4_X1 U5420 ( .A1(n4914), .A2(n4913), .A3(n4912), .A4(n4911), .ZN(n4915)
         );
  NAND4_X1 U5421 ( .A1(n4918), .A2(n4917), .A3(n4916), .A4(n4915), .ZN(n4919)
         );
  AOI211_X1 U5422 ( .C1(DATAO_REG_17__SCAN_IN), .C2(n4921), .A(n4920), .B(
        n4919), .ZN(n4942) );
  XNOR2_X1 U5423 ( .A(n4923), .B(n4922), .ZN(n4924) );
  XNOR2_X1 U5424 ( .A(n4925), .B(n4924), .ZN(n4940) );
  NOR2_X1 U5425 ( .A1(n4927), .A2(n4926), .ZN(n4928) );
  AOI211_X1 U5426 ( .C1(n4931), .C2(n4930), .A(n4929), .B(n4928), .ZN(n4935)
         );
  NAND2_X1 U5427 ( .A1(n4933), .A2(n4932), .ZN(n4934) );
  OAI211_X1 U5428 ( .C1(n4937), .C2(n4936), .A(n4935), .B(n4934), .ZN(n4938)
         );
  AOI21_X1 U5429 ( .B1(n4940), .B2(n4939), .A(n4938), .ZN(n4941) );
  XNOR2_X1 U5430 ( .A(n4942), .B(n4941), .ZN(U3225) );
endmodule

