

module b15_C_AntiSAT_k_256_1 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
         keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
         keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
         keyinput139, keyinput140, keyinput141, keyinput142, keyinput143,
         keyinput144, keyinput145, keyinput146, keyinput147, keyinput148,
         keyinput149, keyinput150, keyinput151, keyinput152, keyinput153,
         keyinput154, keyinput155, keyinput156, keyinput157, keyinput158,
         keyinput159, keyinput160, keyinput161, keyinput162, keyinput163,
         keyinput164, keyinput165, keyinput166, keyinput167, keyinput168,
         keyinput169, keyinput170, keyinput171, keyinput172, keyinput173,
         keyinput174, keyinput175, keyinput176, keyinput177, keyinput178,
         keyinput179, keyinput180, keyinput181, keyinput182, keyinput183,
         keyinput184, keyinput185, keyinput186, keyinput187, keyinput188,
         keyinput189, keyinput190, keyinput191, keyinput192, keyinput193,
         keyinput194, keyinput195, keyinput196, keyinput197, keyinput198,
         keyinput199, keyinput200, keyinput201, keyinput202, keyinput203,
         keyinput204, keyinput205, keyinput206, keyinput207, keyinput208,
         keyinput209, keyinput210, keyinput211, keyinput212, keyinput213,
         keyinput214, keyinput215, keyinput216, keyinput217, keyinput218,
         keyinput219, keyinput220, keyinput221, keyinput222, keyinput223,
         keyinput224, keyinput225, keyinput226, keyinput227, keyinput228,
         keyinput229, keyinput230, keyinput231, keyinput232, keyinput233,
         keyinput234, keyinput235, keyinput236, keyinput237, keyinput238,
         keyinput239, keyinput240, keyinput241, keyinput242, keyinput243,
         keyinput244, keyinput245, keyinput246, keyinput247, keyinput248,
         keyinput249, keyinput250, keyinput251, keyinput252, keyinput253,
         keyinput254, keyinput255;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124;

  AND2_X1 U3635 ( .A1(n5773), .A2(n4863), .ZN(n5939) );
  AND2_X1 U3636 ( .A1(n3573), .A2(n4595), .ZN(n4597) );
  CLKBUF_X2 U3637 ( .A(n4246), .Z(n5641) );
  CLKBUF_X2 U3638 ( .A(n3606), .Z(n3526) );
  CLKBUF_X1 U3640 ( .A(n3348), .Z(n4941) );
  CLKBUF_X2 U3641 ( .A(n3476), .Z(n4423) );
  INV_X1 U3643 ( .A(n3433), .ZN(n3454) );
  AND2_X2 U3644 ( .A1(n4517), .A2(n4659), .ZN(n3481) );
  AND2_X2 U3645 ( .A1(n4659), .A2(n4516), .ZN(n3476) );
  AND2_X1 U3646 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4673) );
  CLKBUF_X3 U3647 ( .A(n3407), .Z(n4167) );
  INV_X1 U3648 ( .A(n5963), .ZN(n5932) );
  OR3_X1 U3649 ( .A1(n6711), .A2(n6607), .A3(n4471), .ZN(n5773) );
  NAND2_X2 U3650 ( .A1(n3201), .A2(n3191), .ZN(n3428) );
  INV_X1 U3651 ( .A(n5929), .ZN(n5776) );
  INV_X1 U3652 ( .A(n5939), .ZN(n5973) );
  OR2_X1 U3653 ( .A1(n4588), .A2(n4237), .ZN(n6092) );
  INV_X2 U3654 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3223) );
  NAND2_X2 U3655 ( .A1(n3348), .A2(n3433), .ZN(n3421) );
  AND2_X4 U3656 ( .A1(n3199), .A2(n3324), .ZN(n3455) );
  AND2_X2 U3657 ( .A1(n4321), .A2(n4246), .ZN(n4601) );
  BUF_X2 U3658 ( .A(n4781), .Z(n3187) );
  XNOR2_X1 U3659 ( .A(n3575), .B(n3551), .ZN(n4781) );
  AND4_X2 U3660 ( .A1(n3309), .A2(n3308), .A3(n3307), .A4(n3306), .ZN(n3201)
         );
  OAI22_X2 U3661 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n5474), .B1(n5484), .B2(n5466), .ZN(n5467) );
  AOI21_X1 U3662 ( .B1(n5234), .B2(n4400), .A(n5221), .ZN(n5446) );
  CLKBUF_X1 U3663 ( .A(n5512), .Z(n5513) );
  INV_X4 U3664 ( .A(n5534), .ZN(n5514) );
  NOR2_X1 U3665 ( .A1(n5683), .A2(n5684), .ZN(n5671) );
  NAND2_X1 U3666 ( .A1(n3596), .A2(n4693), .ZN(n3652) );
  OAI21_X1 U3667 ( .B1(n4509), .B2(STATE2_REG_0__SCAN_IN), .A(n3505), .ZN(
        n3549) );
  AND2_X1 U3668 ( .A1(n3488), .A2(n4240), .ZN(n4190) );
  NOR2_X1 U3670 ( .A1(n3434), .A2(n3279), .ZN(n3401) );
  CLKBUF_X1 U3671 ( .A(n3409), .Z(n4933) );
  NAND2_X1 U3672 ( .A1(n3295), .A2(n3294), .ZN(n3407) );
  AND4_X2 U3673 ( .A1(n3372), .A2(n3371), .A3(n3370), .A4(n3369), .ZN(n4854)
         );
  AND4_X1 U3674 ( .A1(n3299), .A2(n3298), .A3(n3297), .A4(n3296), .ZN(n3305)
         );
  CLKBUF_X2 U3675 ( .A(n3587), .Z(n3512) );
  CLKBUF_X2 U3676 ( .A(n3391), .Z(n3640) );
  BUF_X2 U3677 ( .A(n3385), .Z(n3987) );
  BUF_X2 U3678 ( .A(n3384), .Z(n4408) );
  BUF_X2 U3679 ( .A(n3507), .Z(n4428) );
  BUF_X2 U3680 ( .A(n3481), .Z(n4388) );
  BUF_X2 U3681 ( .A(n3377), .Z(n3475) );
  CLKBUF_X2 U3682 ( .A(n3355), .Z(n3867) );
  BUF_X2 U3683 ( .A(n3378), .Z(n3506) );
  CLKBUF_X2 U3684 ( .A(n3383), .Z(n3929) );
  AND2_X2 U3685 ( .A1(n4516), .A2(n3289), .ZN(n3606) );
  AND2_X2 U3686 ( .A1(n3289), .A2(n4517), .ZN(n3355) );
  XNOR2_X1 U3687 ( .A(n5424), .B(n5423), .ZN(n5561) );
  XNOR2_X1 U3688 ( .A(n4467), .B(n4466), .ZN(n5191) );
  NAND2_X1 U3689 ( .A1(n5490), .A2(n5489), .ZN(n5488) );
  NOR3_X1 U3690 ( .A1(n4211), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5534), 
        .ZN(n5440) );
  AND2_X1 U3691 ( .A1(n3229), .A2(n3228), .ZN(n5552) );
  AND2_X1 U3692 ( .A1(n5023), .A2(n3781), .ZN(n3783) );
  INV_X1 U3693 ( .A(n4725), .ZN(n3261) );
  XNOR2_X1 U3694 ( .A(n4103), .B(n3683), .ZN(n4114) );
  NAND2_X2 U3695 ( .A1(n4103), .A2(n4125), .ZN(n5534) );
  AND2_X1 U3696 ( .A1(n5671), .A2(n3210), .ZN(n5374) );
  NAND2_X1 U3697 ( .A1(n3240), .A2(n3239), .ZN(n5683) );
  NAND2_X1 U3698 ( .A1(n6010), .A2(n4651), .ZN(n6011) );
  NAND2_X2 U3699 ( .A1(n5989), .A2(n3428), .ZN(n5389) );
  CLKBUF_X1 U3700 ( .A(n4055), .Z(n5723) );
  AOI21_X1 U3701 ( .B1(n3553), .B2(n3552), .A(n3550), .ZN(n3574) );
  AOI21_X1 U3702 ( .B1(n5104), .B2(n3561), .A(n6505), .ZN(n4552) );
  NAND2_X1 U3703 ( .A1(n4197), .A2(n4196), .ZN(n5209) );
  XNOR2_X1 U3704 ( .A(n3549), .B(n3547), .ZN(n3553) );
  AOI21_X1 U3705 ( .B1(n3559), .B2(n3558), .A(n3546), .ZN(n3552) );
  NAND2_X1 U3706 ( .A1(n3581), .A2(n3580), .ZN(n5031) );
  AOI21_X1 U3707 ( .B1(n3577), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3472), 
        .ZN(n3474) );
  NAND2_X1 U3708 ( .A1(n3416), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3442) );
  NAND2_X1 U3709 ( .A1(n3544), .A2(n3543), .ZN(n3558) );
  OR2_X1 U3710 ( .A1(n3682), .A2(n6919), .ZN(n3544) );
  AND2_X1 U3711 ( .A1(n4513), .A2(n3438), .ZN(n3458) );
  AND2_X1 U3712 ( .A1(n3436), .A2(n3460), .ZN(n3426) );
  AND2_X1 U3713 ( .A1(n3425), .A2(n3424), .ZN(n3459) );
  INV_X1 U3714 ( .A(n3455), .ZN(n4240) );
  OR2_X1 U3715 ( .A1(n3537), .A2(n3536), .ZN(n4069) );
  OR2_X1 U3716 ( .A1(n3433), .A2(n4854), .ZN(n4321) );
  OR2_X1 U3717 ( .A1(n3335), .A2(n3334), .ZN(n4221) );
  AND4_X1 U3718 ( .A1(n3323), .A2(n3322), .A3(n3321), .A4(n3320), .ZN(n3324)
         );
  AND4_X1 U3719 ( .A1(n3314), .A2(n3313), .A3(n3312), .A4(n3311), .ZN(n3191)
         );
  NAND2_X2 U3720 ( .A1(n3305), .A2(n3304), .ZN(n3406) );
  AND4_X1 U3721 ( .A1(n3288), .A2(n3287), .A3(n3286), .A4(n3285), .ZN(n3295)
         );
  AND4_X1 U3722 ( .A1(n3354), .A2(n3353), .A3(n3352), .A4(n3351), .ZN(n3372)
         );
  AND4_X1 U3723 ( .A1(n3360), .A2(n3359), .A3(n3358), .A4(n3357), .ZN(n3371)
         );
  AND4_X1 U3724 ( .A1(n3364), .A2(n3363), .A3(n3362), .A4(n3361), .ZN(n3370)
         );
  AND4_X1 U3725 ( .A1(n3382), .A2(n3381), .A3(n3380), .A4(n3379), .ZN(n3399)
         );
  AND4_X1 U3726 ( .A1(n3368), .A2(n3367), .A3(n3366), .A4(n3365), .ZN(n3369)
         );
  AND4_X1 U3727 ( .A1(n3396), .A2(n3395), .A3(n3394), .A4(n3393), .ZN(n3397)
         );
  AND4_X1 U3728 ( .A1(n3376), .A2(n3375), .A3(n3374), .A4(n3373), .ZN(n3400)
         );
  AND4_X1 U3729 ( .A1(n3293), .A2(n3292), .A3(n3291), .A4(n3290), .ZN(n3294)
         );
  AND2_X1 U3730 ( .A1(n3189), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3337) );
  AND2_X2 U3731 ( .A1(n4657), .A2(n4516), .ZN(n3378) );
  AND2_X2 U3732 ( .A1(n3223), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4659)
         );
  NOR2_X2 U3733 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4657) );
  NAND2_X1 U3734 ( .A1(n3216), .A2(n3473), .ZN(n3188) );
  NAND2_X1 U3735 ( .A1(n3216), .A2(n3473), .ZN(n3576) );
  XNOR2_X1 U3736 ( .A(n3188), .B(n5031), .ZN(n4655) );
  AND2_X2 U3737 ( .A1(n4533), .A2(n3289), .ZN(n3384) );
  AND2_X2 U3738 ( .A1(n3414), .A2(n3430), .ZN(n4223) );
  OAI21_X1 U3739 ( .B1(n4694), .B2(n3605), .A(n3604), .ZN(n4611) );
  AND2_X2 U3740 ( .A1(n3409), .A2(n3407), .ZN(n3448) );
  NOR2_X1 U3741 ( .A1(n3652), .A2(n3653), .ZN(n3649) );
  AND2_X1 U3742 ( .A1(n4516), .A2(n3289), .ZN(n3189) );
  INV_X2 U3743 ( .A(n4221), .ZN(n3348) );
  AND2_X2 U3744 ( .A1(n4533), .A2(n4659), .ZN(n3507) );
  AND2_X2 U3745 ( .A1(n4533), .A2(n4673), .ZN(n3356) );
  OAI21_X1 U3746 ( .B1(n5533), .B2(n4137), .A(n4136), .ZN(n5512) );
  NAND2_X2 U3747 ( .A1(n4223), .A2(n4926), .ZN(n4238) );
  OR2_X1 U3748 ( .A1(n4926), .A2(n4854), .ZN(n4271) );
  NAND2_X2 U3749 ( .A1(n3652), .A2(n3597), .ZN(n4694) );
  NOR2_X2 U3750 ( .A1(n5298), .A2(n3267), .ZN(n5378) );
  AOI221_X2 U3751 ( .B1(REIP_REG_23__SCAN_IN), .B2(n5743), .C1(n5742), .C2(
        n5743), .A(n5741), .ZN(n5744) );
  AOI21_X2 U3752 ( .B1(n4114), .B2(n3808), .A(n3685), .ZN(n4745) );
  OAI21_X2 U3753 ( .B1(n5542), .B2(n5543), .A(n5544), .ZN(n5533) );
  AND2_X4 U3754 ( .A1(n4657), .A2(n4517), .ZN(n3383) );
  AND2_X4 U3755 ( .A1(n4517), .A2(n4673), .ZN(n3392) );
  AND2_X4 U3756 ( .A1(n4659), .A2(n4508), .ZN(n3587) );
  OAI21_X2 U3757 ( .B1(n5357), .B2(n5355), .A(n5356), .ZN(n5740) );
  NOR2_X4 U3758 ( .A1(n5365), .A2(n5367), .ZN(n5355) );
  OAI22_X2 U3759 ( .A1(n5495), .A2(n5496), .B1(n5514), .B2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5490) );
  NOR2_X4 U3760 ( .A1(n4143), .A2(n3277), .ZN(n5420) );
  AND2_X2 U3761 ( .A1(n3250), .A2(n3206), .ZN(n4143) );
  NOR2_X1 U3762 ( .A1(n5519), .A2(n5800), .ZN(n3269) );
  NAND2_X1 U3763 ( .A1(n5209), .A2(n6616), .ZN(n4588) );
  INV_X1 U3764 ( .A(n5025), .ZN(n3262) );
  INV_X1 U3765 ( .A(n3633), .ZN(n3653) );
  OR2_X1 U3766 ( .A1(n3504), .A2(n3503), .ZN(n4070) );
  AOI22_X1 U3767 ( .A1(n3476), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3378), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3333) );
  INV_X1 U3768 ( .A(n4415), .ZN(n4442) );
  NOR2_X1 U3769 ( .A1(n5195), .A2(n6609), .ZN(n4415) );
  CLKBUF_X1 U3770 ( .A(n4395), .Z(n4439) );
  OR2_X1 U3771 ( .A1(n3487), .A2(n3486), .ZN(n4071) );
  NAND2_X1 U3772 ( .A1(n3433), .A2(n3434), .ZN(n4246) );
  AND2_X1 U3773 ( .A1(n6505), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4464) );
  AND2_X1 U3774 ( .A1(n4422), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4472)
         );
  NAND2_X1 U3775 ( .A1(n3269), .A2(n3268), .ZN(n3267) );
  INV_X1 U3776 ( .A(n5380), .ZN(n3268) );
  NAND2_X1 U3777 ( .A1(n3195), .A2(n3208), .ZN(n3251) );
  INV_X1 U3778 ( .A(n5375), .ZN(n3235) );
  NOR2_X1 U3779 ( .A1(n4124), .A2(n4123), .ZN(n4125) );
  INV_X2 U3780 ( .A(n3434), .ZN(n4926) );
  INV_X1 U3781 ( .A(n4195), .ZN(n4196) );
  AOI21_X1 U3782 ( .B1(n4194), .B2(n4218), .A(n4193), .ZN(n4195) );
  NAND3_X1 U3783 ( .A1(n4448), .A2(n3428), .A3(n3455), .ZN(n3437) );
  NAND2_X1 U3784 ( .A1(n3618), .A2(n3617), .ZN(n3633) );
  NAND2_X1 U3785 ( .A1(n3668), .A2(n3667), .ZN(n3679) );
  AOI21_X1 U3786 ( .B1(n6710), .B2(n6288), .A(n3417), .ZN(n3441) );
  AND4_X1 U3787 ( .A1(n3458), .A2(n4341), .A3(n3457), .A4(n6617), .ZN(n3465)
         );
  AND2_X1 U3788 ( .A1(n3522), .A2(n3521), .ZN(n3547) );
  OR2_X1 U3789 ( .A1(n3682), .A2(n4930), .ZN(n3521) );
  OR2_X1 U3790 ( .A1(n4123), .A2(n3519), .ZN(n3505) );
  AND2_X1 U3791 ( .A1(n5192), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3619) );
  NOR2_X1 U3792 ( .A1(n5234), .A2(n3273), .ZN(n3272) );
  INV_X1 U3793 ( .A(n4053), .ZN(n3273) );
  NAND2_X1 U3794 ( .A1(n4850), .A2(n3197), .ZN(n3784) );
  AND2_X1 U3795 ( .A1(n3780), .A2(n5148), .ZN(n3779) );
  NOR2_X1 U3796 ( .A1(n4301), .A2(n3237), .ZN(n3236) );
  INV_X1 U3797 ( .A(n5385), .ZN(n3237) );
  INV_X1 U3798 ( .A(n3247), .ZN(n3246) );
  OAI21_X1 U3799 ( .B1(n4131), .B2(n3248), .A(n5076), .ZN(n3247) );
  NAND2_X1 U3800 ( .A1(n4843), .A2(n3192), .ZN(n3221) );
  INV_X1 U3801 ( .A(n4709), .ZN(n3232) );
  INV_X1 U3802 ( .A(n4190), .ZN(n3682) );
  INV_X1 U3803 ( .A(n3469), .ZN(n3577) );
  AOI22_X1 U3804 ( .A1(n3355), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3498), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3292) );
  AOI22_X1 U3805 ( .A1(n4190), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3489), 
        .B2(n4071), .ZN(n3490) );
  INV_X1 U3806 ( .A(n3447), .ZN(n6713) );
  INV_X1 U3807 ( .A(n4601), .ZN(n4327) );
  NOR2_X1 U3808 ( .A1(n3242), .A2(n3241), .ZN(n4594) );
  CLKBUF_X1 U3809 ( .A(n3436), .Z(n4591) );
  OAI21_X1 U3810 ( .B1(n4445), .B2(n5426), .A(n4444), .ZN(n4447) );
  AND2_X1 U3811 ( .A1(n4052), .A2(n3270), .ZN(n4467) );
  AND2_X1 U3812 ( .A1(n3203), .A2(n3271), .ZN(n3270) );
  INV_X1 U3813 ( .A(n4447), .ZN(n3271) );
  NAND2_X1 U3814 ( .A1(n4029), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4375)
         );
  OR2_X1 U3815 ( .A1(n5869), .A2(n4445), .ZN(n3865) );
  NAND2_X1 U3816 ( .A1(n3828), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3859)
         );
  NAND2_X1 U3817 ( .A1(n3734), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3761)
         );
  INV_X1 U3818 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5909) );
  AND4_X1 U3819 ( .A1(n3701), .A2(n3700), .A3(n3699), .A4(n3698), .ZN(n4797)
         );
  INV_X1 U3820 ( .A(n5457), .ZN(n3249) );
  NAND2_X1 U3821 ( .A1(n5362), .A2(n5288), .ZN(n5287) );
  INV_X1 U3822 ( .A(n3219), .ZN(n3218) );
  OAI21_X1 U3823 ( .B1(n4142), .B2(n5504), .A(n5503), .ZN(n3219) );
  NOR2_X1 U3824 ( .A1(n5315), .A2(n5300), .ZN(n3239) );
  INV_X1 U3825 ( .A(n5715), .ZN(n3240) );
  AOI21_X1 U3826 ( .B1(n5804), .B2(n5170), .A(n3193), .ZN(n3244) );
  OR2_X1 U3827 ( .A1(n5084), .A2(n4353), .ZN(n5706) );
  NOR2_X1 U3828 ( .A1(n4709), .A2(n4710), .ZN(n4714) );
  NAND2_X1 U3829 ( .A1(n4235), .A2(n4234), .ZN(n4348) );
  OR2_X1 U3830 ( .A1(n4588), .A2(n4233), .ZN(n4234) );
  NAND2_X1 U3831 ( .A1(n4655), .A2(n6609), .ZN(n3595) );
  AND2_X1 U3832 ( .A1(n4682), .A2(n4681), .ZN(n4685) );
  NAND2_X1 U3833 ( .A1(n5220), .A2(n3227), .ZN(n3226) );
  NAND2_X1 U3834 ( .A1(n5968), .A2(EBX_REG_30__SCAN_IN), .ZN(n3227) );
  AND2_X1 U3835 ( .A1(n5773), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U3836 ( .A1(n4856), .A2(n4476), .ZN(n5958) );
  INV_X1 U3837 ( .A(n4459), .ZN(n3228) );
  NAND2_X1 U3838 ( .A1(n4461), .A2(n4460), .ZN(n3229) );
  AND2_X2 U3839 ( .A1(n4453), .A2(n6616), .ZN(n5989) );
  INV_X1 U3840 ( .A(n6009), .ZN(n6005) );
  NAND2_X1 U3841 ( .A1(n4650), .A2(n6079), .ZN(n6010) );
  OAI21_X1 U3842 ( .B1(n4649), .B2(n4648), .A(n6616), .ZN(n4650) );
  OR2_X1 U3843 ( .A1(n6030), .A2(n6041), .ZN(n6023) );
  NAND2_X1 U3844 ( .A1(n6925), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4147) );
  NAND2_X1 U3845 ( .A1(n3421), .A2(n4591), .ZN(n3457) );
  AND2_X1 U3846 ( .A1(n3356), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3325) );
  AOI22_X1 U3847 ( .A1(n3385), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3377), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3332) );
  AOI22_X1 U3848 ( .A1(n3378), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3300) );
  NAND2_X1 U3849 ( .A1(n4162), .A2(n4147), .ZN(n4181) );
  AND2_X1 U3850 ( .A1(n4149), .A2(n4148), .ZN(n4180) );
  NAND2_X1 U3851 ( .A1(n4181), .A2(n4180), .ZN(n4179) );
  NAND2_X1 U3852 ( .A1(n4179), .A2(n4149), .ZN(n4154) );
  AND2_X1 U3853 ( .A1(n4154), .A2(n4153), .ZN(n4156) );
  INV_X1 U3854 ( .A(n3652), .ZN(n3655) );
  OR2_X1 U3855 ( .A1(n3666), .A2(n3665), .ZN(n4116) );
  OR2_X1 U3856 ( .A1(n3616), .A2(n3615), .ZN(n4106) );
  OAI21_X1 U3857 ( .B1(n3469), .B2(n3283), .A(n3446), .ZN(n3523) );
  AND2_X1 U3858 ( .A1(n3455), .A2(n4221), .ZN(n3410) );
  NAND2_X1 U3859 ( .A1(n3435), .A2(n3408), .ZN(n4513) );
  INV_X1 U3860 ( .A(n4246), .ZN(n3435) );
  AOI22_X1 U3861 ( .A1(n3606), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3322) );
  AOI22_X1 U3862 ( .A1(n3476), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3378), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3320) );
  AOI22_X1 U3863 ( .A1(n3385), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3384), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3323) );
  AOI21_X1 U3864 ( .B1(n3391), .B2(INSTQUEUE_REG_1__4__SCAN_IN), .A(n3315), 
        .ZN(n3316) );
  AND2_X1 U3865 ( .A1(n3356), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3315) );
  AOI22_X1 U3866 ( .A1(n3587), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3481), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3288) );
  AOI22_X1 U3867 ( .A1(n3606), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3336), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3290) );
  AOI22_X1 U3868 ( .A1(n3378), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3291) );
  NAND2_X1 U3869 ( .A1(n4854), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3582) );
  AOI21_X1 U3870 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n6589), .A(n4156), 
        .ZN(n4152) );
  NOR2_X1 U3871 ( .A1(n3421), .A2(n4167), .ZN(n3349) );
  AOI21_X1 U3872 ( .B1(n3392), .B2(INSTQUEUE_REG_12__7__SCAN_IN), .A(n3310), 
        .ZN(n3312) );
  AND2_X1 U3873 ( .A1(n3507), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3310) );
  AOI21_X1 U3874 ( .B1(n3336), .B2(INSTQUEUE_REG_2__3__SCAN_IN), .A(n3337), 
        .ZN(n3341) );
  NAND2_X1 U3875 ( .A1(n4006), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4027)
         );
  NAND2_X1 U3876 ( .A1(n3764), .A2(n3763), .ZN(n3780) );
  NOR2_X1 U3877 ( .A1(n3598), .A2(n4616), .ZN(n3621) );
  OAI211_X1 U3878 ( .C1(n3602), .C2(n3223), .A(n3568), .B(n3567), .ZN(n3571)
         );
  OR2_X1 U3879 ( .A1(n3518), .A2(n3517), .ZN(n4127) );
  INV_X1 U3880 ( .A(n5171), .ZN(n3245) );
  INV_X1 U3881 ( .A(n4318), .ZN(n4305) );
  NOR2_X1 U3882 ( .A1(n3234), .A2(n4710), .ZN(n3233) );
  INV_X1 U3883 ( .A(n4713), .ZN(n3234) );
  NAND2_X1 U3884 ( .A1(n4295), .A2(n4246), .ZN(n4318) );
  AND3_X1 U3885 ( .A1(n3348), .A2(n3402), .A3(n3454), .ZN(n3405) );
  NAND2_X1 U3886 ( .A1(n3455), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4123) );
  INV_X1 U3887 ( .A(n4127), .ZN(n3545) );
  OR2_X1 U3888 ( .A1(n3418), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3419)
         );
  AND2_X1 U3889 ( .A1(n3336), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3390) );
  AND2_X2 U3890 ( .A1(n3284), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3289)
         );
  OR2_X1 U3891 ( .A1(n5723), .A2(n6832), .ZN(n6410) );
  OR2_X1 U3892 ( .A1(n6514), .A2(n3470), .ZN(n4767) );
  INV_X1 U3893 ( .A(n3406), .ZN(n3409) );
  OR2_X1 U3894 ( .A1(n3593), .A2(n3592), .ZN(n4088) );
  NOR2_X1 U3895 ( .A1(n4854), .A2(n6609), .ZN(n3488) );
  AOI21_X1 U3896 ( .B1(n6611), .B2(n4684), .A(n4654), .ZN(n4770) );
  INV_X1 U3897 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6925) );
  INV_X1 U3898 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6363) );
  AND2_X1 U3899 ( .A1(n4190), .A2(n4151), .ZN(n4171) );
  NAND2_X1 U3900 ( .A1(n4123), .A2(n3582), .ZN(n4194) );
  OR2_X1 U3901 ( .A1(n4588), .A2(n5210), .ZN(n4559) );
  INV_X1 U3902 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3796) );
  NOR2_X1 U3903 ( .A1(n5237), .A2(n5225), .ZN(n4457) );
  INV_X1 U3904 ( .A(n4246), .ZN(n5382) );
  NAND2_X1 U3905 ( .A1(n5253), .A2(n5235), .ZN(n5237) );
  INV_X1 U3906 ( .A(n4321), .ZN(n4450) );
  NAND2_X1 U3907 ( .A1(n4552), .A2(n4551), .ZN(n3566) );
  AOI22_X1 U3908 ( .A1(n4420), .A2(n4419), .B1(n4439), .B2(n5433), .ZN(n5222)
         );
  OAI21_X1 U3909 ( .B1(n4445), .B2(n5444), .A(n4399), .ZN(n5234) );
  AOI21_X1 U3910 ( .B1(n4051), .B2(n4050), .A(n4049), .ZN(n4053) );
  OR2_X1 U3911 ( .A1(n4033), .A2(n4032), .ZN(n5263) );
  NOR2_X1 U3912 ( .A1(n3265), .A2(n3264), .ZN(n3263) );
  INV_X1 U3913 ( .A(n5357), .ZN(n3265) );
  INV_X1 U3914 ( .A(n5286), .ZN(n3264) );
  NAND2_X1 U3915 ( .A1(n3982), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4005)
         );
  INV_X1 U3916 ( .A(n3981), .ZN(n3982) );
  NAND2_X1 U3917 ( .A1(n3940), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3981)
         );
  INV_X1 U3918 ( .A(n3918), .ZN(n3919) );
  CLKBUF_X1 U3919 ( .A(n5365), .Z(n5366) );
  AND2_X1 U3920 ( .A1(n3904), .A2(n3903), .ZN(n5498) );
  NAND2_X1 U3921 ( .A1(n3901), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3918)
         );
  AND2_X1 U3922 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n3860), .ZN(n3899)
         );
  INV_X1 U3923 ( .A(n3269), .ZN(n3266) );
  NAND2_X1 U3924 ( .A1(n3843), .A2(n3842), .ZN(n5800) );
  AND2_X1 U3925 ( .A1(n3814), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3828)
         );
  CLKBUF_X1 U3926 ( .A(n5298), .Z(n5799) );
  AND3_X1 U3927 ( .A1(n3813), .A2(n3812), .A3(n3811), .ZN(n5314) );
  CLKBUF_X1 U3928 ( .A(n5312), .Z(n5313) );
  AND2_X1 U3929 ( .A1(n3775), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3762)
         );
  AOI21_X1 U3930 ( .B1(n3749), .B2(n4439), .A(n3748), .ZN(n5025) );
  CLKBUF_X1 U3931 ( .A(n5023), .Z(n5024) );
  NAND2_X1 U3932 ( .A1(n3702), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3703)
         );
  INV_X1 U3933 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6997) );
  NAND2_X1 U3934 ( .A1(n4835), .A2(n3258), .ZN(n3257) );
  INV_X1 U3935 ( .A(n4797), .ZN(n3258) );
  AND2_X1 U3936 ( .A1(n3697), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3702)
         );
  NAND2_X1 U3937 ( .A1(n3670), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3672)
         );
  INV_X1 U3938 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3671) );
  NOR2_X1 U3939 ( .A1(n3672), .A2(n3671), .ZN(n3697) );
  INV_X1 U3940 ( .A(n3629), .ZN(n3630) );
  CLKBUF_X1 U3941 ( .A(n4705), .Z(n4706) );
  OR2_X1 U3942 ( .A1(n5732), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4200) );
  NAND2_X1 U3943 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3598) );
  AOI21_X1 U3944 ( .B1(n3187), .B2(n4151), .A(n4074), .ZN(n6109) );
  OR2_X1 U3945 ( .A1(n4236), .A2(n3450), .ZN(n4237) );
  NOR2_X1 U3946 ( .A1(n5553), .A2(n5423), .ZN(n3254) );
  NOR2_X1 U3947 ( .A1(n5251), .A2(n5264), .ZN(n5253) );
  NAND2_X1 U3948 ( .A1(n3238), .A2(n3212), .ZN(n5264) );
  AND2_X1 U3949 ( .A1(n5374), .A2(n4309), .ZN(n5362) );
  NAND2_X1 U3950 ( .A1(n5671), .A2(n3236), .ZN(n5376) );
  OR2_X1 U3951 ( .A1(n5534), .A2(n4140), .ZN(n4141) );
  NAND2_X1 U3952 ( .A1(n3198), .A2(n4285), .ZN(n5715) );
  AND2_X1 U3953 ( .A1(n4348), .A2(n4343), .ZN(n5703) );
  NOR2_X1 U3954 ( .A1(n5027), .A2(n5026), .ZN(n5150) );
  NAND2_X1 U3955 ( .A1(n3221), .A2(n3194), .ZN(n5181) );
  INV_X1 U3956 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3220) );
  OR2_X1 U3957 ( .A1(n4852), .A2(n4853), .ZN(n5027) );
  AND2_X1 U3958 ( .A1(n4828), .A2(n4829), .ZN(n4838) );
  NAND2_X1 U3959 ( .A1(n4838), .A2(n4837), .ZN(n4852) );
  OR2_X1 U3960 ( .A1(n4734), .A2(n4352), .ZN(n5084) );
  NOR2_X1 U3961 ( .A1(n4754), .A2(n4747), .ZN(n4828) );
  NAND2_X1 U3962 ( .A1(n3232), .A2(n3230), .ZN(n4754) );
  AND2_X1 U3963 ( .A1(n3233), .A2(n3231), .ZN(n3230) );
  INV_X1 U3964 ( .A(n4751), .ZN(n3231) );
  NAND2_X1 U3965 ( .A1(n6095), .A2(n6094), .ZN(n3214) );
  NAND2_X1 U3966 ( .A1(n3232), .A2(n3233), .ZN(n4752) );
  NAND2_X1 U3967 ( .A1(n4254), .A2(n4253), .ZN(n4709) );
  INV_X1 U3968 ( .A(n4689), .ZN(n4253) );
  INV_X1 U3969 ( .A(n3474), .ZN(n3473) );
  OR2_X1 U3970 ( .A1(n3460), .A2(n3823), .ZN(n5195) );
  AND2_X1 U3971 ( .A1(n6367), .A2(n6442), .ZN(n6232) );
  AND2_X1 U3972 ( .A1(n4694), .A2(n5727), .ZN(n6231) );
  NAND2_X1 U3973 ( .A1(n3187), .A2(n4695), .ZN(n6338) );
  OR2_X1 U3974 ( .A1(n5723), .A2(n5104), .ZN(n6413) );
  OR2_X1 U3975 ( .A1(n4694), .A2(n3187), .ZN(n6471) );
  INV_X1 U3976 ( .A(n6230), .ZN(n6337) );
  AND2_X1 U3977 ( .A1(n6925), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6514)
         );
  OR3_X1 U3978 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4770), .A3(n4054), .ZN(n4942) );
  AND2_X1 U3979 ( .A1(n5723), .A2(n4061), .ZN(n6230) );
  NOR2_X1 U3980 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4770), .ZN(n4940) );
  AND2_X1 U3981 ( .A1(n3187), .A2(n4760), .ZN(n4882) );
  AND3_X1 U3982 ( .A1(n4679), .A2(n4678), .A3(n5837), .ZN(n6597) );
  AND2_X1 U3983 ( .A1(n6858), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4198) );
  INV_X2 U3984 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6505) );
  INV_X1 U3985 ( .A(n4200), .ZN(n6710) );
  NAND2_X1 U3986 ( .A1(n4559), .A2(n5736), .ZN(n6711) );
  NOR2_X2 U3987 ( .A1(n4907), .A2(n4478), .ZN(n5963) );
  XNOR2_X1 U3988 ( .A(n4600), .B(n3242), .ZN(n4577) );
  AND2_X1 U3989 ( .A1(n6010), .A2(n5192), .ZN(n5997) );
  AND2_X1 U3990 ( .A1(n6010), .A2(n5390), .ZN(n6000) );
  INV_X1 U3991 ( .A(n6011), .ZN(n6006) );
  INV_X1 U3992 ( .A(n6010), .ZN(n5999) );
  NAND2_X1 U3993 ( .A1(n6010), .A2(n4652), .ZN(n6009) );
  AND2_X1 U3994 ( .A1(n4590), .A2(n6602), .ZN(n6030) );
  INV_X2 U3995 ( .A(n6023), .ZN(n6040) );
  INV_X1 U3996 ( .A(n6045), .ZN(n6083) );
  INV_X1 U3997 ( .A(n6054), .ZN(n6045) );
  XNOR2_X1 U3998 ( .A(n4474), .B(n4491), .ZN(n4862) );
  OR2_X1 U3999 ( .A1(n4473), .A2(n5216), .ZN(n4474) );
  INV_X1 U4000 ( .A(n4472), .ZN(n4473) );
  OAI21_X1 U4001 ( .B1(n5221), .B2(n5222), .A(n4446), .ZN(n5438) );
  AOI21_X1 U4002 ( .B1(n6088), .B2(n5254), .A(n4207), .ZN(n4208) );
  OAI21_X1 U4003 ( .B1(n4052), .B2(n4053), .A(n4400), .ZN(n5401) );
  NAND2_X1 U4004 ( .A1(n3243), .A2(n5169), .ZN(n5805) );
  OR2_X1 U4005 ( .A1(n5168), .A2(n5171), .ZN(n3243) );
  INV_X1 U4006 ( .A(n4745), .ZN(n3259) );
  INV_X1 U4007 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4616) );
  INV_X1 U4008 ( .A(n6117), .ZN(n6088) );
  INV_X1 U4009 ( .A(n5528), .ZN(n6108) );
  INV_X2 U4010 ( .A(n5494), .ZN(n6113) );
  XNOR2_X1 U4011 ( .A(n3255), .B(n4213), .ZN(n4503) );
  NAND2_X1 U4012 ( .A1(n3280), .A2(n3252), .ZN(n3255) );
  NOR2_X1 U4013 ( .A1(n5422), .A2(n5421), .ZN(n5424) );
  NOR2_X1 U4014 ( .A1(n5439), .A2(n5553), .ZN(n5422) );
  NAND2_X1 U4015 ( .A1(n4143), .A2(n5448), .ZN(n4144) );
  OR2_X1 U4016 ( .A1(n5604), .A2(n4368), .ZN(n5599) );
  NAND2_X1 U4017 ( .A1(n3250), .A2(n3251), .ZN(n5458) );
  NAND2_X1 U4018 ( .A1(n5671), .A2(n5385), .ZN(n5640) );
  NOR2_X1 U4019 ( .A1(n5699), .A2(n5823), .ZN(n5689) );
  NAND2_X1 U4020 ( .A1(n4841), .A2(n4131), .ZN(n5077) );
  AND2_X1 U4021 ( .A1(n4348), .A2(n4346), .ZN(n6190) );
  OR2_X1 U4022 ( .A1(n5829), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4582)
         );
  AND2_X1 U4023 ( .A1(n4348), .A2(n6581), .ZN(n5829) );
  INV_X1 U4024 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6580) );
  CLKBUF_X1 U4025 ( .A(n4509), .Z(n4510) );
  INV_X1 U4026 ( .A(n3187), .ZN(n5727) );
  CLKBUF_X1 U4027 ( .A(n4655), .Z(n6441) );
  INV_X1 U4028 ( .A(n6519), .ZN(n6506) );
  AND2_X1 U4029 ( .A1(n4223), .A2(n3434), .ZN(n6581) );
  INV_X1 U4030 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6858) );
  INV_X1 U4031 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5840) );
  INV_X1 U4032 ( .A(n6725), .ZN(n6253) );
  OR2_X1 U4033 ( .A1(n6338), .A2(n6413), .ZN(n6293) );
  INV_X1 U4034 ( .A(n6293), .ZN(n6323) );
  INV_X1 U4035 ( .A(n6405), .ZN(n6366) );
  INV_X1 U4036 ( .A(n6538), .ZN(n6379) );
  INV_X1 U4037 ( .A(n6544), .ZN(n6383) );
  INV_X1 U4038 ( .A(n6550), .ZN(n6387) );
  INV_X1 U4039 ( .A(n6556), .ZN(n6391) );
  INV_X1 U4040 ( .A(n6562), .ZN(n6395) );
  NOR2_X2 U4041 ( .A1(n6471), .A2(n6413), .ZN(n6466) );
  INV_X1 U4042 ( .A(n6390), .ZN(n6547) );
  INV_X1 U4043 ( .A(n6394), .ZN(n6551) );
  NOR2_X1 U4044 ( .A1(n6065), .A2(n4881), .ZN(n6364) );
  INV_X1 U4045 ( .A(n4946), .ZN(n5002) );
  INV_X1 U4046 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6609) );
  NAND2_X1 U4047 ( .A1(n5209), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6610) );
  INV_X1 U4048 ( .A(n6714), .ZN(n6611) );
  AND2_X1 U4049 ( .A1(n4198), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6616) );
  INV_X1 U4050 ( .A(n6622), .ZN(n6698) );
  OAI21_X1 U4051 ( .B1(n5552), .B2(n5958), .A(n3224), .ZN(U2797) );
  AOI21_X1 U4052 ( .B1(n5428), .B2(n5929), .A(n3225), .ZN(n3224) );
  OR2_X1 U4053 ( .A1(n5217), .A2(n3226), .ZN(n3225) );
  OAI22_X1 U4054 ( .A1(n5552), .A2(n5984), .B1(n6860), .B2(n5989), .ZN(n4462)
         );
  INV_X1 U4055 ( .A(n4854), .ZN(n3436) );
  AND2_X1 U4056 ( .A1(n5773), .A2(n4475), .ZN(n5929) );
  NAND2_X1 U4057 ( .A1(n4854), .A2(n3434), .ZN(n3449) );
  AND2_X1 U4058 ( .A1(n4842), .A2(n5075), .ZN(n3192) );
  OAI211_X1 U4059 ( .C1(n3469), .C2(n3282), .A(n3442), .B(n3441), .ZN(n3467)
         );
  AND2_X1 U4060 ( .A1(n5534), .A2(n4135), .ZN(n3193) );
  AND2_X1 U4061 ( .A1(n3246), .A2(n3220), .ZN(n3194) );
  NAND2_X1 U4062 ( .A1(n3275), .A2(n4142), .ZN(n3195) );
  NAND2_X1 U4063 ( .A1(n4850), .A2(n3733), .ZN(n4849) );
  AND2_X1 U4064 ( .A1(n3733), .A2(n3262), .ZN(n3196) );
  NAND2_X1 U4065 ( .A1(n3261), .A2(n3259), .ZN(n4795) );
  AND2_X1 U4066 ( .A1(n3196), .A2(n3779), .ZN(n3197) );
  NOR2_X1 U4067 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4395) );
  NOR2_X2 U4068 ( .A1(n3406), .A2(n6505), .ZN(n3808) );
  AOI21_X1 U4069 ( .B1(n4781), .B2(n3808), .A(n4464), .ZN(n4596) );
  AND2_X2 U4070 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4516) );
  AND2_X1 U4071 ( .A1(n5150), .A2(n5149), .ZN(n3198) );
  AND4_X1 U4072 ( .A1(n3319), .A2(n3318), .A3(n3317), .A4(n3316), .ZN(n3199)
         );
  AND3_X1 U4073 ( .A1(n4224), .A2(n3453), .A3(n3452), .ZN(n3200) );
  AND2_X2 U4074 ( .A1(n4533), .A2(n4657), .ZN(n3336) );
  NAND2_X1 U4075 ( .A1(n3440), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3469) );
  INV_X1 U4076 ( .A(n4143), .ZN(n4211) );
  OR2_X1 U4077 ( .A1(n5401), .A2(n5494), .ZN(n3202) );
  AND2_X1 U4078 ( .A1(n3455), .A2(n4167), .ZN(n3408) );
  NAND2_X1 U4079 ( .A1(n5355), .A2(n3263), .ZN(n5272) );
  OR2_X1 U4080 ( .A1(n5298), .A2(n5800), .ZN(n5517) );
  AND2_X1 U4081 ( .A1(n5222), .A2(n3272), .ZN(n3203) );
  NAND2_X1 U4082 ( .A1(n5420), .A2(n5449), .ZN(n5439) );
  INV_X1 U4083 ( .A(n5075), .ZN(n3248) );
  NAND2_X1 U4084 ( .A1(n5534), .A2(n5089), .ZN(n5075) );
  AOI21_X1 U4085 ( .B1(n4446), .B2(n4447), .A(n4467), .ZN(n5428) );
  OR2_X1 U4086 ( .A1(n5298), .A2(n3266), .ZN(n5379) );
  AND2_X1 U4087 ( .A1(n3245), .A2(n5804), .ZN(n3204) );
  NAND2_X1 U4088 ( .A1(n5476), .A2(n4142), .ZN(n3205) );
  AND2_X1 U4089 ( .A1(n3251), .A2(n3249), .ZN(n3206) );
  OR2_X1 U4090 ( .A1(n3428), .A2(n6505), .ZN(n3281) );
  NAND2_X1 U4091 ( .A1(n3595), .A2(n3594), .ZN(n4693) );
  NAND2_X1 U4092 ( .A1(n3221), .A2(n3246), .ZN(n4132) );
  AND2_X1 U4093 ( .A1(n3214), .A2(n3213), .ZN(n3207) );
  NAND2_X1 U4094 ( .A1(n5534), .A2(n4368), .ZN(n3208) );
  INV_X1 U4095 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3282) );
  NAND2_X1 U4096 ( .A1(n3222), .A2(n3244), .ZN(n5542) );
  NAND2_X1 U4097 ( .A1(n4134), .A2(n4133), .ZN(n5168) );
  NAND2_X1 U4098 ( .A1(n4843), .A2(n4842), .ZN(n4841) );
  INV_X1 U4099 ( .A(n3238), .ZN(n5277) );
  NOR2_X1 U4100 ( .A1(n5287), .A2(n5275), .ZN(n3238) );
  AND2_X1 U4101 ( .A1(n3261), .A2(n3260), .ZN(n4796) );
  AND2_X1 U4102 ( .A1(n3278), .A2(n3208), .ZN(n3209) );
  AND2_X1 U4103 ( .A1(n3236), .A2(n3235), .ZN(n3210) );
  AND2_X1 U4104 ( .A1(n3263), .A2(n4009), .ZN(n3211) );
  NAND2_X1 U4105 ( .A1(n3261), .A2(n3256), .ZN(n4834) );
  INV_X1 U4106 ( .A(n4271), .ZN(n4295) );
  NOR2_X1 U4107 ( .A1(n4230), .A2(n4854), .ZN(n4468) );
  INV_X1 U4108 ( .A(n4395), .ZN(n4445) );
  AND2_X1 U4109 ( .A1(n4574), .A2(n4575), .ZN(n3570) );
  NAND2_X1 U4110 ( .A1(n4573), .A2(n3572), .ZN(n4595) );
  NAND2_X1 U4111 ( .A1(n4317), .A2(n4316), .ZN(n3212) );
  AND2_X2 U4112 ( .A1(n3282), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4508)
         );
  AND2_X2 U4113 ( .A1(n3283), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4533)
         );
  NAND2_X1 U4114 ( .A1(n3214), .A2(n4113), .ZN(n4822) );
  OR2_X1 U4115 ( .A1(n6095), .A2(n6094), .ZN(n3213) );
  NAND2_X1 U4116 ( .A1(n3468), .A2(n3467), .ZN(n3217) );
  NAND2_X2 U4117 ( .A1(n3576), .A2(n3215), .ZN(n4536) );
  NAND2_X1 U4118 ( .A1(n3217), .A2(n3474), .ZN(n3215) );
  INV_X1 U4119 ( .A(n3217), .ZN(n3216) );
  OAI21_X2 U4120 ( .B1(n5476), .B2(n5504), .A(n3218), .ZN(n5495) );
  NAND3_X1 U4121 ( .A1(n4134), .A2(n3204), .A3(n4133), .ZN(n3222) );
  NAND2_X1 U4122 ( .A1(n4594), .A2(n4593), .ZN(n4690) );
  NOR2_X1 U4123 ( .A1(n4600), .A2(n3190), .ZN(n3241) );
  NAND2_X1 U4124 ( .A1(n4245), .A2(n4244), .ZN(n3242) );
  NAND2_X1 U4125 ( .A1(n4139), .A2(n3209), .ZN(n3250) );
  NAND2_X1 U4126 ( .A1(n4139), .A2(n3278), .ZN(n5476) );
  INV_X1 U4127 ( .A(n5439), .ZN(n3253) );
  NAND2_X1 U4128 ( .A1(n3253), .A2(n3254), .ZN(n3252) );
  NOR2_X1 U4129 ( .A1(n4745), .A2(n4797), .ZN(n3260) );
  NOR2_X1 U4130 ( .A1(n4745), .A2(n3257), .ZN(n3256) );
  AND2_X1 U4131 ( .A1(n4850), .A2(n3196), .ZN(n5023) );
  NAND2_X1 U4132 ( .A1(n3784), .A2(n3780), .ZN(n5807) );
  NAND2_X1 U4133 ( .A1(n5355), .A2(n3211), .ZN(n5262) );
  AND2_X1 U4134 ( .A1(n5355), .A2(n5357), .ZN(n5285) );
  NAND2_X1 U4135 ( .A1(n4052), .A2(n3203), .ZN(n4446) );
  AND2_X1 U4136 ( .A1(n4052), .A2(n3272), .ZN(n5221) );
  NAND2_X1 U4137 ( .A1(n4052), .A2(n4053), .ZN(n4400) );
  NAND2_X1 U4138 ( .A1(n3403), .A2(n4854), .ZN(n3431) );
  AND2_X1 U4139 ( .A1(n3648), .A2(n3647), .ZN(n3274) );
  OR2_X1 U4140 ( .A1(n3276), .A2(n5534), .ZN(n3275) );
  AND4_X1 U4141 ( .A1(n5627), .A2(n5608), .A3(n5664), .A4(n6933), .ZN(n3276)
         );
  AND2_X1 U4142 ( .A1(n5534), .A2(n6887), .ZN(n3277) );
  NOR2_X1 U4143 ( .A1(n5523), .A2(n4138), .ZN(n3278) );
  XOR2_X1 U4144 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .Z(n3279) );
  NAND2_X1 U4145 ( .A1(n3455), .A2(n4167), .ZN(n3450) );
  NAND2_X1 U4146 ( .A1(n5440), .A2(n4212), .ZN(n3280) );
  NAND2_X1 U4147 ( .A1(n5989), .A2(n5189), .ZN(n5984) );
  INV_X1 U4148 ( .A(n6092), .ZN(n4502) );
  OR2_X1 U4149 ( .A1(n4532), .A2(n4649), .ZN(n6577) );
  INV_X1 U4150 ( .A(n4230), .ZN(n4521) );
  INV_X1 U4151 ( .A(n4703), .ZN(n4704) );
  INV_X1 U4152 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n4054) );
  AND2_X2 U4153 ( .A1(n4508), .A2(n3289), .ZN(n3385) );
  INV_X1 U4154 ( .A(n4194), .ZN(n4182) );
  NOR2_X1 U4155 ( .A1(n4182), .A2(n4215), .ZN(n4184) );
  NOR2_X1 U4156 ( .A1(n3653), .A2(n3274), .ZN(n3654) );
  OR2_X1 U4157 ( .A1(n3682), .A2(n4923), .ZN(n3648) );
  INV_X1 U4158 ( .A(n4070), .ZN(n3519) );
  NAND2_X1 U4159 ( .A1(n6580), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4165) );
  NAND2_X1 U4160 ( .A1(n6363), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4149) );
  OR2_X1 U4161 ( .A1(n3682), .A2(n4937), .ZN(n3668) );
  OR2_X1 U4162 ( .A1(n3682), .A2(n4919), .ZN(n3618) );
  OR2_X1 U4163 ( .A1(n4160), .A2(n4165), .ZN(n4162) );
  INV_X1 U4164 ( .A(n3434), .ZN(n3403) );
  INV_X1 U4165 ( .A(n3678), .ZN(n3680) );
  INV_X1 U4166 ( .A(n4071), .ZN(n4079) );
  AND3_X1 U4167 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n4152), .A3(n5840), 
        .ZN(n4158) );
  INV_X1 U4168 ( .A(n4005), .ZN(n4006) );
  OR2_X1 U4169 ( .A1(n3646), .A2(n3645), .ZN(n4105) );
  NOR2_X1 U4170 ( .A1(n4158), .A2(n4157), .ZN(n4217) );
  INV_X1 U4171 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3858) );
  INV_X1 U4172 ( .A(n5274), .ZN(n4009) );
  AND2_X1 U4173 ( .A1(n4376), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4377)
         );
  AND2_X1 U4174 ( .A1(n4028), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4029)
         );
  INV_X1 U4175 ( .A(n5372), .ZN(n3923) );
  INV_X1 U4176 ( .A(n4848), .ZN(n3733) );
  INV_X1 U4177 ( .A(n3603), .ZN(n3604) );
  AND2_X1 U4178 ( .A1(n4279), .A2(n4278), .ZN(n5149) );
  AND2_X1 U4179 ( .A1(n4167), .A2(n3434), .ZN(n4151) );
  AOI221_X1 U4180 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n4152), .C1(
        n5840), .C2(n4152), .A(n4150), .ZN(n4218) );
  NOR2_X1 U4181 ( .A1(n3859), .A2(n3858), .ZN(n3860) );
  NOR2_X1 U4182 ( .A1(n4907), .A2(n6601), .ZN(n4856) );
  AND2_X1 U4183 ( .A1(n4252), .A2(n4251), .ZN(n4689) );
  OR2_X1 U4184 ( .A1(n4551), .A2(n4445), .ZN(n3565) );
  OR2_X1 U4185 ( .A1(n4588), .A2(n4587), .ZN(n4589) );
  NAND2_X1 U4186 ( .A1(n4377), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4421)
         );
  AND2_X1 U4187 ( .A1(n3899), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3901)
         );
  AND2_X1 U4188 ( .A1(n3784), .A2(n5148), .ZN(n5806) );
  AND2_X1 U4189 ( .A1(n5524), .A2(n4141), .ZN(n4142) );
  INV_X1 U4190 ( .A(n6722), .ZN(n5137) );
  INV_X1 U4191 ( .A(n4468), .ZN(n5210) );
  NAND2_X1 U4192 ( .A1(n5773), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4907) );
  NOR2_X1 U4193 ( .A1(n3796), .A2(n3795), .ZN(n3814) );
  NOR2_X1 U4194 ( .A1(n6997), .A2(n3703), .ZN(n3734) );
  INV_X1 U4195 ( .A(n5960), .ZN(n5934) );
  AND2_X1 U4196 ( .A1(n4862), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4863) );
  AND2_X1 U4197 ( .A1(n4265), .A2(n4264), .ZN(n4747) );
  NAND2_X1 U4198 ( .A1(n6085), .A2(n4589), .ZN(n4590) );
  AND2_X1 U4199 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n3919), .ZN(n3940)
         );
  NOR2_X1 U4200 ( .A1(n3761), .A2(n5909), .ZN(n3775) );
  CLKBUF_X1 U4201 ( .A(n4725), .Z(n4746) );
  AND2_X1 U4202 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3621), .ZN(n3670)
         );
  INV_X1 U4203 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4213) );
  AND2_X1 U4204 ( .A1(n5651), .A2(n5185), .ZN(n6125) );
  INV_X1 U4205 ( .A(n4733), .ZN(n5694) );
  OR2_X1 U4206 ( .A1(n5732), .A2(n6624), .ZN(n6177) );
  INV_X1 U4207 ( .A(n6189), .ZN(n6119) );
  INV_X1 U4208 ( .A(n6365), .ZN(n5036) );
  OR2_X1 U4209 ( .A1(n5723), .A2(n4061), .ZN(n6365) );
  INV_X1 U4210 ( .A(n6563), .ZN(n5018) );
  INV_X1 U4211 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6589) );
  AOI21_X1 U4212 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6580), .A(n4881), .ZN(
        n6521) );
  NAND2_X1 U4213 ( .A1(n4054), .A2(n6505), .ZN(n6519) );
  OAI21_X1 U4214 ( .B1(n5347), .B2(n5958), .A(n4495), .ZN(n4496) );
  NOR2_X1 U4215 ( .A1(n5932), .A2(n4479), .ZN(n5767) );
  INV_X1 U4216 ( .A(n5958), .ZN(n5904) );
  INV_X1 U4217 ( .A(n5984), .ZN(n5980) );
  AND2_X1 U4218 ( .A1(n6010), .A2(n5189), .ZN(n5190) );
  OAI21_X1 U4219 ( .B1(n3447), .B2(n6635), .A(n5735), .ZN(n6054) );
  NAND2_X1 U4220 ( .A1(n3762), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3795)
         );
  NAND2_X1 U4221 ( .A1(n6092), .A2(n4202), .ZN(n5528) );
  INV_X1 U4222 ( .A(n5721), .ZN(n4243) );
  NOR2_X1 U4223 ( .A1(n5599), .A2(n5590), .ZN(n5585) );
  OR2_X1 U4224 ( .A1(n5619), .A2(n4362), .ZN(n5606) );
  OR2_X1 U4225 ( .A1(n5829), .A2(n5703), .ZN(n5653) );
  OR2_X1 U4226 ( .A1(n5653), .A2(n6190), .ZN(n4733) );
  AND2_X1 U4227 ( .A1(n5653), .A2(n4582), .ZN(n6196) );
  AND2_X1 U4228 ( .A1(n4348), .A2(n4331), .ZN(n6189) );
  INV_X1 U4229 ( .A(n4940), .ZN(n4881) );
  INV_X1 U4230 ( .A(n6610), .ZN(n4654) );
  AND2_X1 U4231 ( .A1(n6231), .A2(n5036), .ZN(n6225) );
  AND2_X1 U4232 ( .A1(n6231), .A2(n5106), .ZN(n6724) );
  AND2_X1 U4233 ( .A1(n6329), .A2(n5036), .ZN(n6283) );
  AND2_X1 U4234 ( .A1(n5030), .A2(n6506), .ZN(n6264) );
  INV_X1 U4235 ( .A(n6327), .ZN(n6354) );
  INV_X1 U4236 ( .A(n6532), .ZN(n6375) );
  INV_X1 U4237 ( .A(n6572), .ZN(n6401) );
  NOR2_X2 U4238 ( .A1(n6471), .A2(n6365), .ZN(n6432) );
  AND2_X1 U4239 ( .A1(n6442), .A2(n6441), .ZN(n6474) );
  AND2_X1 U4240 ( .A1(n4799), .A2(n5104), .ZN(n6563) );
  INV_X1 U4241 ( .A(n6386), .ZN(n6539) );
  INV_X1 U4242 ( .A(n4815), .ZN(n6567) );
  OR2_X1 U4243 ( .A1(n6599), .A2(n6598), .ZN(n6600) );
  INV_X1 U4244 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6636) );
  INV_X1 U4245 ( .A(n6689), .ZN(n6690) );
  INV_X1 U4246 ( .A(n4496), .ZN(n4497) );
  INV_X1 U4247 ( .A(n5968), .ZN(n5746) );
  INV_X1 U4248 ( .A(n4825), .ZN(n5345) );
  NAND2_X1 U4249 ( .A1(n6030), .A2(n4591), .ZN(n4644) );
  OR2_X1 U4250 ( .A1(n4684), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6708) );
  INV_X1 U4251 ( .A(n6030), .ZN(n6043) );
  OR2_X1 U4252 ( .A1(n4588), .A2(n6604), .ZN(n6085) );
  OR3_X2 U4253 ( .A1(n4588), .A2(READY_N), .A3(n4560), .ZN(n6079) );
  NAND2_X1 U4254 ( .A1(n5528), .A2(n4205), .ZN(n6117) );
  XNOR2_X1 U4255 ( .A(n4145), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5587)
         );
  NAND2_X1 U4256 ( .A1(n4348), .A2(n4242), .ZN(n5721) );
  INV_X1 U4257 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6202) );
  AOI21_X1 U4258 ( .B1(n6207), .B2(n4786), .A(n4785), .ZN(n4950) );
  NAND2_X1 U4259 ( .A1(n6231), .A2(n5105), .ZN(n6725) );
  NAND2_X1 U4260 ( .A1(n6231), .A2(n6230), .ZN(n6287) );
  AOI21_X1 U4261 ( .B1(n6264), .B2(n5034), .A(n5033), .ZN(n5071) );
  OR2_X1 U4262 ( .A1(n6338), .A2(n6438), .ZN(n6327) );
  OR2_X1 U4263 ( .A1(n6338), .A2(n6337), .ZN(n6405) );
  INV_X1 U4264 ( .A(n6412), .ZN(n6437) );
  AOI22_X1 U4265 ( .A1(n6444), .A2(n6474), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6443), .ZN(n6470) );
  NOR2_X1 U4266 ( .A1(n4804), .A2(n4803), .ZN(n5022) );
  INV_X1 U4267 ( .A(n6364), .ZN(n6723) );
  NOR2_X1 U4268 ( .A1(n4765), .A2(n4764), .ZN(n4982) );
  OR2_X1 U4269 ( .A1(n4761), .A2(n4061), .ZN(n5006) );
  AND2_X1 U4270 ( .A1(n6606), .A2(n6605), .ZN(n6622) );
  INV_X1 U4271 ( .A(n6696), .ZN(n6627) );
  AND2_X1 U4272 ( .A1(n6636), .A2(STATE_REG_1__SCAN_IN), .ZN(n6678) );
  INV_X1 U4273 ( .A(n6687), .ZN(n6692) );
  OAI21_X1 U4274 ( .B1(n5393), .B2(n5389), .A(n4463), .ZN(U2829) );
  NOR2_X4 U4275 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4517) );
  INV_X1 U4276 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3283) );
  AOI22_X1 U4277 ( .A1(n3507), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3287) );
  INV_X1 U4278 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3284) );
  AOI22_X1 U4279 ( .A1(n3384), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3383), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3286) );
  AND2_X4 U4280 ( .A1(n4657), .A2(n4508), .ZN(n3391) );
  AOI22_X1 U4281 ( .A1(n3391), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3285) );
  AND2_X2 U4282 ( .A1(n4508), .A2(n4673), .ZN(n3377) );
  AOI22_X1 U4283 ( .A1(n3377), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3385), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3293) );
  AND2_X4 U4284 ( .A1(n4516), .A2(n4673), .ZN(n3498) );
  INV_X1 U4285 ( .A(n3407), .ZN(n3402) );
  AOI22_X1 U4286 ( .A1(n3507), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U4287 ( .A1(n3391), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4288 ( .A1(n3587), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3355), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3297) );
  AOI22_X1 U4289 ( .A1(n3481), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3498), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3296) );
  AOI22_X1 U4290 ( .A1(n3385), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3384), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3303) );
  AOI22_X1 U4291 ( .A1(n3606), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3336), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3302) );
  AOI22_X1 U4292 ( .A1(n3377), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3383), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3301) );
  AND4_X2 U4293 ( .A1(n3303), .A2(n3302), .A3(n3301), .A4(n3300), .ZN(n3304)
         );
  NAND2_X1 U4294 ( .A1(n3402), .A2(n3406), .ZN(n4448) );
  BUF_X4 U4295 ( .A(n3336), .Z(n4383) );
  AOI22_X1 U4296 ( .A1(n3606), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4297 ( .A1(n3385), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3384), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3308) );
  AOI22_X1 U4298 ( .A1(n3377), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3383), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3307) );
  AOI22_X1 U4299 ( .A1(n3476), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3378), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3306) );
  AOI22_X1 U4300 ( .A1(n3391), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4301 ( .A1(n3587), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3355), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4302 ( .A1(n3481), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3498), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3311) );
  AOI22_X1 U4303 ( .A1(n3507), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3319) );
  AOI22_X1 U4304 ( .A1(n3481), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3498), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3318) );
  AOI22_X1 U4305 ( .A1(n3587), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3355), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3317) );
  AOI22_X1 U4306 ( .A1(n3377), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3383), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3321) );
  INV_X1 U4307 ( .A(n3437), .ZN(n3350) );
  AOI21_X1 U4308 ( .B1(n3391), .B2(INSTQUEUE_REG_1__2__SCAN_IN), .A(n3325), 
        .ZN(n3329) );
  AOI22_X1 U4309 ( .A1(n3587), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3481), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3328) );
  AOI22_X1 U4310 ( .A1(n3606), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3336), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3327) );
  AOI22_X1 U4311 ( .A1(n3384), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3383), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3326) );
  NAND4_X1 U4312 ( .A1(n3329), .A2(n3328), .A3(n3327), .A4(n3326), .ZN(n3335)
         );
  AOI22_X1 U4313 ( .A1(n3507), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3331) );
  AOI22_X1 U4314 ( .A1(n3355), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3498), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3330) );
  NAND4_X1 U4315 ( .A1(n3333), .A2(n3332), .A3(n3331), .A4(n3330), .ZN(n3334)
         );
  AOI22_X1 U4316 ( .A1(n3385), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3384), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3340) );
  AOI22_X1 U4317 ( .A1(n3377), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3383), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3339) );
  AOI22_X1 U4318 ( .A1(n3476), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3378), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3338) );
  NAND4_X1 U4319 ( .A1(n3341), .A2(n3340), .A3(n3339), .A4(n3338), .ZN(n3347)
         );
  AOI22_X1 U4320 ( .A1(n3587), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3355), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3345) );
  AOI22_X1 U4321 ( .A1(n3391), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3344) );
  AOI22_X1 U4322 ( .A1(n3507), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3343) );
  AOI22_X1 U4323 ( .A1(n3481), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3498), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3342) );
  NAND4_X1 U4324 ( .A1(n3345), .A2(n3344), .A3(n3343), .A4(n3342), .ZN(n3346)
         );
  OR2_X2 U4325 ( .A1(n3347), .A2(n3346), .ZN(n3433) );
  NAND2_X1 U4326 ( .A1(n3350), .A2(n3349), .ZN(n4230) );
  NAND2_X1 U4327 ( .A1(n3476), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3354)
         );
  NAND2_X1 U4328 ( .A1(n3385), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3353) );
  NAND2_X1 U4329 ( .A1(n3384), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3352) );
  NAND2_X1 U4330 ( .A1(n3378), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3351) );
  NAND2_X1 U4331 ( .A1(n3587), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3360) );
  NAND2_X1 U4332 ( .A1(n3355), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3359) );
  NAND2_X1 U4333 ( .A1(n3391), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3358) );
  NAND2_X1 U4334 ( .A1(n3356), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3357)
         );
  NAND2_X1 U4335 ( .A1(n3377), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3364)
         );
  NAND2_X1 U4336 ( .A1(n3606), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3363) );
  NAND2_X1 U4337 ( .A1(n3336), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3362) );
  NAND2_X1 U4338 ( .A1(n3383), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3361) );
  NAND2_X1 U4339 ( .A1(n3507), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3368)
         );
  NAND2_X1 U4340 ( .A1(n3481), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3367) );
  NAND2_X1 U4341 ( .A1(n3392), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3366)
         );
  NAND2_X1 U4342 ( .A1(n3498), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3365)
         );
  NAND2_X1 U4343 ( .A1(n3507), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3376)
         );
  NAND2_X1 U4344 ( .A1(n3587), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3375) );
  NAND2_X1 U4345 ( .A1(n3355), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3374) );
  NAND2_X1 U4346 ( .A1(n3356), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3373)
         );
  NAND2_X1 U4347 ( .A1(n3476), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3382)
         );
  NAND2_X1 U4348 ( .A1(n3606), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3381) );
  NAND2_X1 U4349 ( .A1(n3377), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3380)
         );
  NAND2_X1 U4350 ( .A1(n3378), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3379) );
  NAND2_X1 U4351 ( .A1(n3383), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3388) );
  NAND2_X1 U4352 ( .A1(n3384), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3387) );
  NAND2_X1 U4353 ( .A1(n3385), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3386) );
  NAND3_X1 U4354 ( .A1(n3388), .A2(n3387), .A3(n3386), .ZN(n3389) );
  NOR2_X2 U4355 ( .A1(n3390), .A2(n3389), .ZN(n3398) );
  NAND2_X1 U4356 ( .A1(n3481), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3396) );
  NAND2_X1 U4357 ( .A1(n3391), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3395) );
  NAND2_X1 U4358 ( .A1(n3392), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3394)
         );
  NAND2_X1 U4359 ( .A1(n3498), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3393)
         );
  NAND4_X4 U4360 ( .A1(n3400), .A2(n3399), .A3(n3398), .A4(n3397), .ZN(n3434)
         );
  INV_X1 U4361 ( .A(n3401), .ZN(n3422) );
  INV_X1 U4362 ( .A(n3431), .ZN(n3404) );
  NAND2_X1 U4363 ( .A1(n3405), .A2(n3404), .ZN(n4512) );
  NAND2_X1 U4364 ( .A1(n3406), .A2(n3428), .ZN(n4332) );
  NOR2_X1 U4365 ( .A1(n4512), .A2(n4332), .ZN(n4239) );
  AOI21_X1 U4366 ( .B1(n4468), .B2(n3422), .A(n4239), .ZN(n3415) );
  OR2_X2 U4367 ( .A1(n3448), .A2(n3454), .ZN(n3429) );
  AND4_X2 U4368 ( .A1(n3429), .A2(n4854), .A3(n3408), .A4(n3428), .ZN(n3414)
         );
  NAND2_X1 U4369 ( .A1(n3428), .A2(n4933), .ZN(n3456) );
  NAND3_X1 U4370 ( .A1(n3410), .A2(n4448), .A3(n3456), .ZN(n3413) );
  OAI21_X1 U4371 ( .B1(n3455), .B2(n3406), .A(n4448), .ZN(n3411) );
  NAND2_X1 U4372 ( .A1(n3411), .A2(n3348), .ZN(n3412) );
  NAND2_X1 U4373 ( .A1(n3413), .A2(n3412), .ZN(n3430) );
  NAND2_X1 U4374 ( .A1(n3415), .A2(n4238), .ZN(n3416) );
  INV_X1 U4375 ( .A(n3442), .ZN(n3420) );
  NAND2_X1 U4376 ( .A1(n4054), .A2(n6858), .ZN(n5732) );
  XNOR2_X1 U4377 ( .A(n6925), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6288)
         );
  INV_X1 U4378 ( .A(n4198), .ZN(n3444) );
  AND2_X1 U4379 ( .A1(n3444), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3417)
         );
  INV_X1 U4380 ( .A(n3441), .ZN(n3418) );
  NAND2_X1 U4381 ( .A1(n3420), .A2(n3419), .ZN(n3443) );
  OAI21_X1 U4382 ( .B1(n3401), .B2(n4167), .A(n3449), .ZN(n3423) );
  NOR2_X1 U4383 ( .A1(n3421), .A2(n3423), .ZN(n3427) );
  NAND2_X1 U4384 ( .A1(n3448), .A2(n3455), .ZN(n3425) );
  AND2_X1 U4385 ( .A1(n4448), .A2(n3428), .ZN(n3424) );
  INV_X1 U4386 ( .A(n3448), .ZN(n3460) );
  NAND2_X1 U4387 ( .A1(n3437), .A2(n3426), .ZN(n4334) );
  AND3_X1 U4388 ( .A1(n3427), .A2(n3459), .A3(n4334), .ZN(n3439) );
  NAND3_X1 U4389 ( .A1(n3430), .A2(n3428), .A3(n3429), .ZN(n3432) );
  NAND2_X1 U4390 ( .A1(n3432), .A2(n3404), .ZN(n3452) );
  AND2_X2 U4391 ( .A1(n3436), .A2(n4926), .ZN(n3447) );
  NAND2_X1 U4392 ( .A1(n3447), .A2(n3437), .ZN(n3438) );
  NAND3_X1 U4393 ( .A1(n3439), .A2(n3452), .A3(n3458), .ZN(n3440) );
  NAND2_X1 U4394 ( .A1(n3443), .A2(n3467), .ZN(n3493) );
  INV_X1 U4395 ( .A(n3493), .ZN(n3466) );
  MUX2_X1 U4396 ( .A(n3444), .B(n6710), .S(n6580), .Z(n3445) );
  INV_X1 U4397 ( .A(n3445), .ZN(n3446) );
  NAND2_X1 U4398 ( .A1(n3447), .A2(n3448), .ZN(n4224) );
  INV_X1 U4399 ( .A(n3449), .ZN(n3451) );
  NAND2_X1 U4400 ( .A1(n3451), .A2(n3450), .ZN(n3453) );
  INV_X1 U4401 ( .A(n3456), .ZN(n3561) );
  NAND4_X1 U4402 ( .A1(n3454), .A2(n4941), .A3(n4240), .A4(n3561), .ZN(n4341)
         );
  INV_X1 U4403 ( .A(n3421), .ZN(n4056) );
  NOR2_X1 U4404 ( .A1(n5732), .A2(n6609), .ZN(n6617) );
  INV_X1 U4405 ( .A(n3459), .ZN(n3463) );
  NAND2_X1 U4406 ( .A1(n3460), .A2(n4240), .ZN(n3461) );
  NAND2_X1 U4407 ( .A1(n3461), .A2(n3433), .ZN(n3462) );
  OAI21_X1 U4408 ( .B1(n3463), .B2(n3462), .A(n3434), .ZN(n3464) );
  NAND3_X1 U4409 ( .A1(n3200), .A2(n3465), .A3(n3464), .ZN(n3524) );
  NAND2_X1 U4410 ( .A1(n3523), .A2(n3524), .ZN(n3492) );
  NAND2_X1 U4411 ( .A1(n3466), .A2(n3492), .ZN(n3468) );
  NOR2_X1 U4412 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6925), .ZN(n6445)
         );
  NAND2_X1 U4413 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6445), .ZN(n6475) );
  OAI21_X1 U4414 ( .B1(n6363), .B2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n6475), 
        .ZN(n3470) );
  NAND2_X1 U4415 ( .A1(n6710), .A2(n4767), .ZN(n3471) );
  OAI21_X1 U4416 ( .B1(n4198), .B2(n6363), .A(n3471), .ZN(n3472) );
  AOI22_X1 U4417 ( .A1(n3987), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3480) );
  AOI22_X1 U4418 ( .A1(n3606), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3479) );
  AOI22_X1 U4419 ( .A1(n3475), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3478) );
  AOI22_X1 U4420 ( .A1(n4423), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3477) );
  NAND4_X1 U4421 ( .A1(n3480), .A2(n3479), .A3(n3478), .A4(n3477), .ZN(n3487)
         );
  AOI22_X1 U4422 ( .A1(n3512), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3485) );
  INV_X1 U4423 ( .A(n3356), .ZN(n3639) );
  AOI22_X1 U4424 ( .A1(n3391), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3690), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3484) );
  AOI22_X1 U4425 ( .A1(n4428), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3483) );
  AOI22_X1 U4426 ( .A1(n4388), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3482) );
  NAND4_X1 U4427 ( .A1(n3485), .A2(n3484), .A3(n3483), .A4(n3482), .ZN(n3486)
         );
  OAI22_X2 U4428 ( .A1(n4536), .A2(STATE2_REG_0__SCAN_IN), .B1(n4079), .B2(
        n4123), .ZN(n3491) );
  INV_X1 U4429 ( .A(n3582), .ZN(n3489) );
  XNOR2_X2 U4430 ( .A(n3491), .B(n3490), .ZN(n3575) );
  XNOR2_X1 U4431 ( .A(n3493), .B(n3492), .ZN(n4509) );
  AOI22_X1 U4432 ( .A1(n4408), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3497) );
  AOI22_X1 U4433 ( .A1(n4428), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3496) );
  AOI22_X1 U4434 ( .A1(n4388), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3690), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3495) );
  AOI22_X1 U4435 ( .A1(n3987), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3494) );
  NAND4_X1 U4436 ( .A1(n3497), .A2(n3496), .A3(n3495), .A4(n3494), .ZN(n3504)
         );
  AOI22_X1 U4437 ( .A1(n3512), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3502) );
  AOI22_X1 U4438 ( .A1(n4423), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3383), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3501) );
  AOI22_X1 U4439 ( .A1(n3606), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3500) );
  BUF_X1 U4440 ( .A(n3498), .Z(n3531) );
  AOI22_X1 U4441 ( .A1(n3867), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3499) );
  NAND4_X1 U4442 ( .A1(n3502), .A2(n3501), .A3(n3500), .A4(n3499), .ZN(n3503)
         );
  AOI22_X1 U4443 ( .A1(n3867), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3640), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3511) );
  AOI22_X1 U4444 ( .A1(n3606), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3510) );
  AOI22_X1 U4445 ( .A1(n4423), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3509) );
  AOI22_X1 U4446 ( .A1(n4428), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3508) );
  NAND4_X1 U4447 ( .A1(n3511), .A2(n3510), .A3(n3509), .A4(n3508), .ZN(n3518)
         );
  AOI22_X1 U4448 ( .A1(n3987), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3516) );
  AOI22_X1 U4449 ( .A1(n3512), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3690), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3515) );
  AOI22_X1 U4450 ( .A1(n3475), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U4451 ( .A1(n4388), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3513) );
  NAND4_X1 U4452 ( .A1(n3516), .A2(n3515), .A3(n3514), .A4(n3513), .ZN(n3517)
         );
  OAI22_X1 U4453 ( .A1(n4123), .A2(n4127), .B1(n3582), .B2(n3519), .ZN(n3520)
         );
  INV_X1 U4454 ( .A(n3520), .ZN(n3522) );
  INV_X1 U4455 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4930) );
  INV_X1 U4456 ( .A(n3523), .ZN(n3525) );
  XNOR2_X1 U4457 ( .A(n3525), .B(n3524), .ZN(n3562) );
  NAND2_X1 U4458 ( .A1(n3562), .A2(n6609), .ZN(n3540) );
  INV_X1 U4459 ( .A(n4123), .ZN(n3539) );
  AOI22_X1 U4460 ( .A1(n3987), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3530) );
  AOI22_X1 U4461 ( .A1(n3475), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3606), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3529) );
  AOI22_X1 U4462 ( .A1(n3512), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3690), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3528) );
  BUF_X1 U4463 ( .A(n3392), .Z(n4403) );
  AOI22_X1 U4464 ( .A1(n3867), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3527) );
  NAND4_X1 U4465 ( .A1(n3530), .A2(n3529), .A3(n3528), .A4(n3527), .ZN(n3537)
         );
  AOI22_X1 U4466 ( .A1(n4428), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3535) );
  AOI22_X1 U4467 ( .A1(n4423), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3534) );
  AOI22_X1 U4468 ( .A1(n4383), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3533) );
  AOI22_X1 U4469 ( .A1(n3640), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3532) );
  NAND4_X1 U4470 ( .A1(n3535), .A2(n3534), .A3(n3533), .A4(n3532), .ZN(n3536)
         );
  XNOR2_X1 U4471 ( .A(n3545), .B(n4069), .ZN(n3538) );
  NAND2_X1 U4472 ( .A1(n3539), .A2(n3538), .ZN(n3560) );
  NAND2_X1 U4473 ( .A1(n3540), .A2(n3560), .ZN(n3559) );
  INV_X1 U4474 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n6919) );
  NAND2_X1 U4475 ( .A1(n4854), .A2(n4069), .ZN(n3541) );
  OAI211_X1 U4476 ( .C1(n3545), .C2(n4240), .A(STATE2_REG_0__SCAN_IN), .B(
        n3541), .ZN(n3542) );
  INV_X1 U4477 ( .A(n3542), .ZN(n3543) );
  NOR2_X1 U4478 ( .A1(n4123), .A2(n3545), .ZN(n3546) );
  INV_X1 U4479 ( .A(n3547), .ZN(n3548) );
  NOR2_X1 U4480 ( .A1(n3549), .A2(n3548), .ZN(n3550) );
  INV_X1 U4481 ( .A(n3574), .ZN(n3551) );
  XNOR2_X1 U4482 ( .A(n3553), .B(n3552), .ZN(n4055) );
  NAND2_X1 U4483 ( .A1(n4055), .A2(n3808), .ZN(n3557) );
  INV_X2 U4484 ( .A(n3281), .ZN(n4465) );
  AOI22_X1 U4485 ( .A1(n4465), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6505), .ZN(n3555) );
  INV_X1 U4486 ( .A(n4332), .ZN(n5192) );
  NAND2_X1 U4487 ( .A1(n3619), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3554) );
  AND2_X1 U4488 ( .A1(n3555), .A2(n3554), .ZN(n3556) );
  NAND2_X1 U4489 ( .A1(n3557), .A2(n3556), .ZN(n4574) );
  MUX2_X2 U4490 ( .A(n3560), .B(n3559), .S(n3558), .Z(n5104) );
  INV_X1 U4491 ( .A(n3619), .ZN(n3602) );
  NAND2_X1 U4493 ( .A1(n4686), .A2(n3808), .ZN(n3564) );
  AOI22_X1 U4494 ( .A1(n4465), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6505), .ZN(n3563) );
  OAI211_X1 U4495 ( .C1(n3602), .C2(n3283), .A(n3564), .B(n3563), .ZN(n4551)
         );
  NAND2_X1 U4496 ( .A1(n3566), .A2(n3565), .ZN(n4575) );
  OAI21_X1 U4497 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3598), .ZN(n6116) );
  AOI22_X1 U4498 ( .A1(n4464), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n4439), 
        .B2(n6116), .ZN(n3568) );
  NAND2_X1 U4499 ( .A1(n4465), .A2(EAX_REG_2__SCAN_IN), .ZN(n3567) );
  NAND2_X1 U4500 ( .A1(n3570), .A2(n3571), .ZN(n3569) );
  NAND2_X1 U4501 ( .A1(n4596), .A2(n3569), .ZN(n3573) );
  INV_X1 U4502 ( .A(n3570), .ZN(n4573) );
  INV_X1 U4503 ( .A(n3571), .ZN(n3572) );
  AND2_X2 U4504 ( .A1(n3575), .A2(n3574), .ZN(n3596) );
  NAND2_X1 U4505 ( .A1(n3577), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3581) );
  NOR3_X1 U4506 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6363), .A3(n6925), 
        .ZN(n6336) );
  NAND2_X1 U4507 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6336), .ZN(n6330) );
  NAND2_X1 U4508 ( .A1(n6589), .A2(n6330), .ZN(n3578) );
  NOR3_X1 U4509 ( .A1(n6589), .A2(n6363), .A3(n6925), .ZN(n4886) );
  NAND2_X1 U4510 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4886), .ZN(n4999) );
  NAND2_X1 U4511 ( .A1(n3578), .A2(n4999), .ZN(n4802) );
  OAI22_X1 U4512 ( .A1(n4200), .A2(n4802), .B1(n4198), .B2(n6589), .ZN(n3579)
         );
  INV_X1 U4513 ( .A(n3579), .ZN(n3580) );
  AOI22_X1 U4514 ( .A1(n3987), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3526), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4515 ( .A1(n4408), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3585) );
  AOI22_X1 U4516 ( .A1(n4428), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3584) );
  AOI22_X1 U4517 ( .A1(n3634), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3583) );
  NAND4_X1 U4518 ( .A1(n3586), .A2(n3585), .A3(n3584), .A4(n3583), .ZN(n3593)
         );
  AOI22_X1 U4519 ( .A1(n3512), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4520 ( .A1(n4423), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3590) );
  INV_X1 U4521 ( .A(n3639), .ZN(n3690) );
  AOI22_X1 U4522 ( .A1(n3690), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3589) );
  AOI22_X1 U4523 ( .A1(n4388), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3588) );
  NAND4_X1 U4524 ( .A1(n3591), .A2(n3590), .A3(n3589), .A4(n3588), .ZN(n3592)
         );
  AOI22_X1 U4525 ( .A1(n4190), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4194), 
        .B2(n4088), .ZN(n3594) );
  OR2_X2 U4526 ( .A1(n3596), .A2(n4693), .ZN(n3597) );
  INV_X1 U4527 ( .A(n3808), .ZN(n3605) );
  INV_X1 U4528 ( .A(n3598), .ZN(n3599) );
  INV_X1 U4529 ( .A(n3621), .ZN(n3622) );
  OAI21_X1 U4530 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3599), .A(n3622), 
        .ZN(n4614) );
  AOI22_X1 U4531 ( .A1(n4439), .A2(n4614), .B1(n4464), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3601) );
  NAND2_X1 U4532 ( .A1(n4465), .A2(EAX_REG_3__SCAN_IN), .ZN(n3600) );
  OAI211_X1 U4533 ( .C1(n3602), .C2(n3284), .A(n3601), .B(n3600), .ZN(n3603)
         );
  NAND2_X1 U4534 ( .A1(n4597), .A2(n4611), .ZN(n4612) );
  INV_X1 U4535 ( .A(n4612), .ZN(n3632) );
  INV_X1 U4536 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4919) );
  AOI22_X1 U4537 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3987), .B1(n4408), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3610) );
  AOI22_X1 U4538 ( .A1(n3526), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3609) );
  AOI22_X1 U4539 ( .A1(n3475), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3608) );
  AOI22_X1 U4540 ( .A1(n4423), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3607) );
  NAND4_X1 U4541 ( .A1(n3610), .A2(n3609), .A3(n3608), .A4(n3607), .ZN(n3616)
         );
  AOI22_X1 U4542 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n3512), .B1(n3867), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4543 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n3640), .B1(n3690), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3613) );
  AOI22_X1 U4544 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4428), .B1(n4403), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3612) );
  AOI22_X1 U4545 ( .A1(n4388), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3611) );
  NAND4_X1 U4546 ( .A1(n3614), .A2(n3613), .A3(n3612), .A4(n3611), .ZN(n3615)
         );
  NAND2_X1 U4547 ( .A1(n4194), .A2(n4106), .ZN(n3617) );
  XNOR2_X1 U4548 ( .A(n3652), .B(n3633), .ZN(n4087) );
  NAND2_X1 U4549 ( .A1(n4087), .A2(n3808), .ZN(n3631) );
  NAND2_X1 U4550 ( .A1(n3619), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3628) );
  INV_X1 U4551 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3623) );
  AOI21_X1 U4552 ( .B1(n3623), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3620) );
  AOI21_X1 U4553 ( .B1(n4465), .B2(EAX_REG_4__SCAN_IN), .A(n3620), .ZN(n3627)
         );
  INV_X1 U4554 ( .A(n3670), .ZN(n3625) );
  NAND2_X1 U4555 ( .A1(n3623), .A2(n3622), .ZN(n3624) );
  NAND2_X1 U4556 ( .A1(n3625), .A2(n3624), .ZN(n6107) );
  NOR2_X1 U4557 ( .A1(n6107), .A2(n4445), .ZN(n3626) );
  AOI21_X1 U4558 ( .B1(n3628), .B2(n3627), .A(n3626), .ZN(n3629) );
  NAND2_X1 U4559 ( .A1(n3631), .A2(n3630), .ZN(n4703) );
  NAND2_X1 U4560 ( .A1(n3632), .A2(n4703), .ZN(n4705) );
  INV_X1 U4561 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4923) );
  AOI22_X1 U4562 ( .A1(n3987), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3638) );
  INV_X1 U4563 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n6942) );
  AOI22_X1 U4564 ( .A1(n3526), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3637) );
  AOI22_X1 U4565 ( .A1(n3475), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3636) );
  AOI22_X1 U4566 ( .A1(n4423), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3635) );
  NAND4_X1 U4567 ( .A1(n3638), .A2(n3637), .A3(n3636), .A4(n3635), .ZN(n3646)
         );
  AOI22_X1 U4568 ( .A1(n3512), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3644) );
  INV_X1 U4569 ( .A(n3639), .ZN(n3660) );
  AOI22_X1 U4570 ( .A1(n3640), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4571 ( .A1(n4428), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4572 ( .A1(n4388), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3641) );
  NAND4_X1 U4573 ( .A1(n3644), .A2(n3643), .A3(n3642), .A4(n3641), .ZN(n3645)
         );
  NAND2_X1 U4574 ( .A1(n4194), .A2(n4105), .ZN(n3647) );
  XNOR2_X1 U4575 ( .A(n3649), .B(n3274), .ZN(n4095) );
  INV_X1 U4576 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4742) );
  XNOR2_X1 U4577 ( .A(n3670), .B(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5938) );
  AOI22_X1 U4578 ( .A1(n5938), .A2(n4439), .B1(n4464), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3650) );
  OAI21_X1 U4579 ( .B1(n3281), .B2(n4742), .A(n3650), .ZN(n3651) );
  AOI21_X1 U4580 ( .B1(n4095), .B2(n3808), .A(n3651), .ZN(n4712) );
  NOR2_X2 U4581 ( .A1(n4705), .A2(n4712), .ZN(n4727) );
  NAND2_X1 U4582 ( .A1(n3655), .A2(n3654), .ZN(n3678) );
  INV_X1 U4583 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4937) );
  AOI22_X1 U4584 ( .A1(n3987), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3659) );
  AOI22_X1 U4585 ( .A1(n3526), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U4586 ( .A1(n3475), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3657) );
  AOI22_X1 U4587 ( .A1(n4423), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3656) );
  NAND4_X1 U4588 ( .A1(n3659), .A2(n3658), .A3(n3657), .A4(n3656), .ZN(n3666)
         );
  AOI22_X1 U4589 ( .A1(n3512), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3664) );
  AOI22_X1 U4590 ( .A1(n3640), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4591 ( .A1(n4428), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U4592 ( .A1(n4388), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3661) );
  NAND4_X1 U4593 ( .A1(n3664), .A2(n3663), .A3(n3662), .A4(n3661), .ZN(n3665)
         );
  NAND2_X1 U4594 ( .A1(n4194), .A2(n4116), .ZN(n3667) );
  INV_X1 U4595 ( .A(n3679), .ZN(n3669) );
  NAND2_X1 U4596 ( .A1(n3678), .A2(n3669), .ZN(n4104) );
  NAND2_X1 U4597 ( .A1(n4104), .A2(n3808), .ZN(n3677) );
  AND2_X1 U4598 ( .A1(n3672), .A2(n3671), .ZN(n3673) );
  OR2_X1 U4599 ( .A1(n3673), .A2(n3697), .ZN(n6099) );
  INV_X1 U4600 ( .A(n6099), .ZN(n3675) );
  AOI22_X1 U4601 ( .A1(n4465), .A2(EAX_REG_6__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6505), .ZN(n3674) );
  MUX2_X1 U4602 ( .A(n3675), .B(n3674), .S(n4445), .Z(n3676) );
  NAND2_X1 U4603 ( .A1(n3677), .A2(n3676), .ZN(n4726) );
  NAND2_X1 U4604 ( .A1(n4727), .A2(n4726), .ZN(n4725) );
  NAND2_X1 U4605 ( .A1(n3680), .A2(n3679), .ZN(n4103) );
  INV_X1 U4606 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4791) );
  NAND2_X1 U4607 ( .A1(n4194), .A2(n4127), .ZN(n3681) );
  OAI21_X1 U4608 ( .B1(n3682), .B2(n4791), .A(n3681), .ZN(n3683) );
  INV_X1 U4609 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4757) );
  XNOR2_X1 U4610 ( .A(n3697), .B(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5335) );
  AOI22_X1 U4611 ( .A1(n5335), .A2(n4439), .B1(n4464), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3684) );
  OAI21_X1 U4612 ( .B1(n3281), .B2(n4757), .A(n3684), .ZN(n3685) );
  AOI22_X1 U4613 ( .A1(n4408), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4614 ( .A1(n3512), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3640), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4615 ( .A1(n3634), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4616 ( .A1(n4428), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3686) );
  NAND4_X1 U4617 ( .A1(n3689), .A2(n3688), .A3(n3687), .A4(n3686), .ZN(n3696)
         );
  AOI22_X1 U4618 ( .A1(n3987), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3526), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3694) );
  AOI22_X1 U4619 ( .A1(n3867), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3690), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3693) );
  AOI22_X1 U4620 ( .A1(n4423), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3692) );
  AOI22_X1 U4621 ( .A1(n4388), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3691) );
  NAND4_X1 U4622 ( .A1(n3694), .A2(n3693), .A3(n3692), .A4(n3691), .ZN(n3695)
         );
  OAI21_X1 U4623 ( .B1(n3696), .B2(n3695), .A(n3808), .ZN(n3701) );
  NAND2_X1 U4624 ( .A1(n4465), .A2(EAX_REG_8__SCAN_IN), .ZN(n3700) );
  XNOR2_X1 U4625 ( .A(n3702), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5325) );
  NAND2_X1 U4626 ( .A1(n5325), .A2(n4439), .ZN(n3699) );
  NAND2_X1 U4627 ( .A1(n4464), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3698)
         );
  AOI21_X1 U4628 ( .B1(n6997), .B2(n3703), .A(n3734), .ZN(n5918) );
  OR2_X1 U4629 ( .A1(n5918), .A2(n4445), .ZN(n3718) );
  AOI22_X1 U4630 ( .A1(n3987), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4423), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3707) );
  AOI22_X1 U4631 ( .A1(n3867), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4632 ( .A1(n4408), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4633 ( .A1(n4388), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3704) );
  NAND4_X1 U4634 ( .A1(n3707), .A2(n3706), .A3(n3705), .A4(n3704), .ZN(n3713)
         );
  AOI22_X1 U4635 ( .A1(n3512), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3640), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3711) );
  AOI22_X1 U4636 ( .A1(n3526), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3710) );
  AOI22_X1 U4637 ( .A1(n3475), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3709) );
  AOI22_X1 U4638 ( .A1(n4428), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3708) );
  NAND4_X1 U4639 ( .A1(n3711), .A2(n3710), .A3(n3709), .A4(n3708), .ZN(n3712)
         );
  OAI21_X1 U4640 ( .B1(n3713), .B2(n3712), .A(n3808), .ZN(n3716) );
  NAND2_X1 U4641 ( .A1(n4465), .A2(EAX_REG_9__SCAN_IN), .ZN(n3715) );
  NAND2_X1 U4642 ( .A1(n4464), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3714)
         );
  AND3_X1 U4643 ( .A1(n3716), .A2(n3715), .A3(n3714), .ZN(n3717) );
  NAND2_X1 U4644 ( .A1(n3718), .A2(n3717), .ZN(n4835) );
  XNOR2_X1 U4645 ( .A(n3734), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5143)
         );
  AOI22_X1 U4646 ( .A1(n4423), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4647 ( .A1(n3526), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4428), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4648 ( .A1(n3640), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4649 ( .A1(n3867), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3719) );
  NAND4_X1 U4650 ( .A1(n3722), .A2(n3721), .A3(n3720), .A4(n3719), .ZN(n3728)
         );
  AOI22_X1 U4651 ( .A1(n4388), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4652 ( .A1(n3475), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3725) );
  AOI22_X1 U4653 ( .A1(n3987), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4654 ( .A1(n3512), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3723) );
  NAND4_X1 U4655 ( .A1(n3726), .A2(n3725), .A3(n3724), .A4(n3723), .ZN(n3727)
         );
  OAI21_X1 U4656 ( .B1(n3728), .B2(n3727), .A(n3808), .ZN(n3731) );
  NAND2_X1 U4657 ( .A1(n4465), .A2(EAX_REG_10__SCAN_IN), .ZN(n3730) );
  NAND2_X1 U4658 ( .A1(n4464), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3729)
         );
  NAND3_X1 U4659 ( .A1(n3731), .A2(n3730), .A3(n3729), .ZN(n3732) );
  AOI21_X1 U4660 ( .B1(n5143), .B2(n4395), .A(n3732), .ZN(n4848) );
  XOR2_X1 U4661 ( .A(n5909), .B(n3761), .Z(n6087) );
  INV_X1 U4662 ( .A(n6087), .ZN(n3749) );
  AOI22_X1 U4663 ( .A1(n3987), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4428), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4664 ( .A1(n3512), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4665 ( .A1(n3640), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3736) );
  AOI22_X1 U4666 ( .A1(n4388), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3735) );
  NAND4_X1 U4667 ( .A1(n3738), .A2(n3737), .A3(n3736), .A4(n3735), .ZN(n3744)
         );
  AOI22_X1 U4668 ( .A1(n4408), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3742) );
  AOI22_X1 U4669 ( .A1(n4423), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3741) );
  AOI22_X1 U4670 ( .A1(n4383), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3740) );
  AOI22_X1 U4671 ( .A1(n3526), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3739) );
  NAND4_X1 U4672 ( .A1(n3742), .A2(n3741), .A3(n3740), .A4(n3739), .ZN(n3743)
         );
  OAI21_X1 U4673 ( .B1(n3744), .B2(n3743), .A(n3808), .ZN(n3747) );
  NAND2_X1 U4674 ( .A1(n4465), .A2(EAX_REG_11__SCAN_IN), .ZN(n3746) );
  NAND2_X1 U4675 ( .A1(n4464), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3745)
         );
  NAND3_X1 U4676 ( .A1(n3747), .A2(n3746), .A3(n3745), .ZN(n3748) );
  AOI22_X1 U4677 ( .A1(n4408), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4678 ( .A1(n3512), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4679 ( .A1(n3987), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4680 ( .A1(n4388), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3750) );
  NAND4_X1 U4681 ( .A1(n3753), .A2(n3752), .A3(n3751), .A4(n3750), .ZN(n3759)
         );
  AOI22_X1 U4682 ( .A1(n3526), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4683 ( .A1(n3640), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4684 ( .A1(n4423), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4685 ( .A1(n4428), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3754) );
  NAND4_X1 U4686 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n3758)
         );
  OR2_X1 U4687 ( .A1(n3759), .A2(n3758), .ZN(n3760) );
  NAND2_X1 U4688 ( .A1(n3808), .A2(n3760), .ZN(n5810) );
  INV_X1 U4689 ( .A(n5810), .ZN(n3781) );
  NAND2_X1 U4690 ( .A1(n4465), .A2(EAX_REG_13__SCAN_IN), .ZN(n3764) );
  OAI21_X1 U4691 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3762), .A(n3795), 
        .ZN(n5902) );
  AOI22_X1 U4692 ( .A1(n4439), .A2(n5902), .B1(n4464), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4693 ( .A1(n4423), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4694 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3512), .B1(n3867), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4695 ( .A1(n3526), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4696 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4428), .B1(n4403), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3765) );
  NAND4_X1 U4697 ( .A1(n3768), .A2(n3767), .A3(n3766), .A4(n3765), .ZN(n3774)
         );
  AOI22_X1 U4698 ( .A1(n3475), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4699 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n3640), .B1(n3660), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4700 ( .A1(n3987), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4701 ( .A1(n4388), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3769) );
  NAND4_X1 U4702 ( .A1(n3772), .A2(n3771), .A3(n3770), .A4(n3769), .ZN(n3773)
         );
  NOR2_X1 U4703 ( .A1(n3774), .A2(n3773), .ZN(n3778) );
  XNOR2_X1 U4704 ( .A(n3775), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5174)
         );
  NAND2_X1 U4705 ( .A1(n5174), .A2(n4395), .ZN(n3777) );
  AOI22_X1 U4706 ( .A1(n4465), .A2(EAX_REG_12__SCAN_IN), .B1(n4464), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3776) );
  OAI211_X1 U4707 ( .C1(n3778), .C2(n3605), .A(n3777), .B(n3776), .ZN(n5148)
         );
  NOR2_X1 U4708 ( .A1(n5807), .A2(n5810), .ZN(n3782) );
  AOI21_X1 U4709 ( .B1(n3783), .B2(n5806), .A(n3782), .ZN(n5813) );
  NAND2_X1 U4710 ( .A1(n5813), .A2(n3784), .ZN(n5418) );
  AOI22_X1 U4711 ( .A1(n4408), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4712 ( .A1(n3512), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4713 ( .A1(n3640), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4714 ( .A1(n3526), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3785) );
  NAND4_X1 U4715 ( .A1(n3788), .A2(n3787), .A3(n3786), .A4(n3785), .ZN(n3794)
         );
  AOI22_X1 U4716 ( .A1(n4428), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4717 ( .A1(n3987), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4718 ( .A1(n4423), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4719 ( .A1(n3867), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3789) );
  NAND4_X1 U4720 ( .A1(n3792), .A2(n3791), .A3(n3790), .A4(n3789), .ZN(n3793)
         );
  NOR2_X1 U4721 ( .A1(n3794), .A2(n3793), .ZN(n3799) );
  AOI21_X1 U4722 ( .B1(n3796), .B2(n3795), .A(n3814), .ZN(n5889) );
  INV_X1 U4723 ( .A(n5889), .ZN(n5549) );
  AOI22_X1 U4724 ( .A1(n4464), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n4439), 
        .B2(n5549), .ZN(n3798) );
  NAND2_X1 U4725 ( .A1(n4465), .A2(EAX_REG_14__SCAN_IN), .ZN(n3797) );
  OAI211_X1 U4726 ( .C1(n3605), .C2(n3799), .A(n3798), .B(n3797), .ZN(n5419)
         );
  NAND2_X1 U4727 ( .A1(n5418), .A2(n5419), .ZN(n5312) );
  AOI22_X1 U4728 ( .A1(n3867), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4729 ( .A1(n4388), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4730 ( .A1(n3475), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3801) );
  AOI22_X1 U4731 ( .A1(n4423), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3800) );
  NAND4_X1 U4732 ( .A1(n3803), .A2(n3802), .A3(n3801), .A4(n3800), .ZN(n3810)
         );
  AOI22_X1 U4733 ( .A1(n3987), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4734 ( .A1(n3526), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4428), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4735 ( .A1(n3587), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4736 ( .A1(n3392), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3804) );
  NAND4_X1 U4737 ( .A1(n3807), .A2(n3806), .A3(n3805), .A4(n3804), .ZN(n3809)
         );
  OAI21_X1 U4738 ( .B1(n3810), .B2(n3809), .A(n3808), .ZN(n3813) );
  XNOR2_X1 U4739 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3814), .ZN(n5537)
         );
  AOI22_X1 U4740 ( .A1(n4395), .A2(n5537), .B1(n4464), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3812) );
  NAND2_X1 U4741 ( .A1(n4465), .A2(EAX_REG_15__SCAN_IN), .ZN(n3811) );
  NOR2_X2 U4742 ( .A1(n5312), .A2(n5314), .ZN(n5297) );
  XOR2_X1 U4743 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3828), .Z(n5531) );
  AOI22_X1 U4744 ( .A1(n4465), .A2(EAX_REG_16__SCAN_IN), .B1(n4464), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4745 ( .A1(n4408), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4746 ( .A1(n3587), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4747 ( .A1(n3987), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3816) );
  AOI22_X1 U4748 ( .A1(n3867), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3815) );
  NAND4_X1 U4749 ( .A1(n3818), .A2(n3817), .A3(n3816), .A4(n3815), .ZN(n3825)
         );
  AOI22_X1 U4750 ( .A1(n4428), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4751 ( .A1(n3526), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4752 ( .A1(n4423), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4753 ( .A1(n3640), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3498), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3819) );
  NAND4_X1 U4754 ( .A1(n3822), .A2(n3821), .A3(n3820), .A4(n3819), .ZN(n3824)
         );
  NAND2_X1 U4755 ( .A1(n4240), .A2(n3428), .ZN(n3823) );
  OAI21_X1 U4756 ( .B1(n3825), .B2(n3824), .A(n4415), .ZN(n3826) );
  OAI211_X1 U4757 ( .C1(n5531), .C2(n4445), .A(n3827), .B(n3826), .ZN(n5299)
         );
  NAND2_X1 U4758 ( .A1(n5297), .A2(n5299), .ZN(n5298) );
  XNOR2_X1 U4759 ( .A(n3859), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5879)
         );
  NAND2_X1 U4760 ( .A1(n5879), .A2(n4395), .ZN(n3843) );
  AOI22_X1 U4761 ( .A1(n4408), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4762 ( .A1(n4428), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4763 ( .A1(n3512), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3830) );
  AOI22_X1 U4764 ( .A1(n3987), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3829) );
  NAND4_X1 U4765 ( .A1(n3832), .A2(n3831), .A3(n3830), .A4(n3829), .ZN(n3838)
         );
  AOI22_X1 U4766 ( .A1(n3526), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4767 ( .A1(n3867), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4768 ( .A1(n4423), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3834) );
  AOI22_X1 U4769 ( .A1(n4403), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3833) );
  NAND4_X1 U4770 ( .A1(n3836), .A2(n3835), .A3(n3834), .A4(n3833), .ZN(n3837)
         );
  NOR2_X1 U4771 ( .A1(n3838), .A2(n3837), .ZN(n3841) );
  AOI21_X1 U4772 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n3858), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3839) );
  AOI21_X1 U4773 ( .B1(n4465), .B2(EAX_REG_17__SCAN_IN), .A(n3839), .ZN(n3840)
         );
  OAI21_X1 U4774 ( .B1(n4442), .B2(n3841), .A(n3840), .ZN(n3842) );
  AOI22_X1 U4775 ( .A1(n4423), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4776 ( .A1(n3526), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4777 ( .A1(n3475), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4778 ( .A1(n3867), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3844) );
  NAND4_X1 U4779 ( .A1(n3847), .A2(n3846), .A3(n3845), .A4(n3844), .ZN(n3853)
         );
  AOI22_X1 U4780 ( .A1(n3640), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4781 ( .A1(n3987), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4782 ( .A1(n4428), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4783 ( .A1(n3512), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3848) );
  NAND4_X1 U4784 ( .A1(n3851), .A2(n3850), .A3(n3849), .A4(n3848), .ZN(n3852)
         );
  NOR2_X1 U4785 ( .A1(n3853), .A2(n3852), .ZN(n3857) );
  INV_X1 U4786 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6832) );
  OAI21_X1 U4787 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6832), .A(n6505), 
        .ZN(n3854) );
  INV_X1 U4788 ( .A(n3854), .ZN(n3855) );
  AOI21_X1 U4789 ( .B1(n4465), .B2(EAX_REG_18__SCAN_IN), .A(n3855), .ZN(n3856)
         );
  OAI21_X1 U4790 ( .B1(n4442), .B2(n3857), .A(n3856), .ZN(n3866) );
  INV_X1 U4791 ( .A(n3899), .ZN(n3864) );
  INV_X1 U4792 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3862) );
  INV_X1 U4793 ( .A(n3860), .ZN(n3861) );
  NAND2_X1 U4794 ( .A1(n3862), .A2(n3861), .ZN(n3863) );
  NAND2_X1 U4795 ( .A1(n3864), .A2(n3863), .ZN(n5869) );
  NAND2_X1 U4796 ( .A1(n3866), .A2(n3865), .ZN(n5519) );
  AOI22_X1 U4797 ( .A1(n3526), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4798 ( .A1(n3475), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4799 ( .A1(n4408), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3869) );
  AOI22_X1 U4800 ( .A1(n3867), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3868) );
  NAND4_X1 U4801 ( .A1(n3871), .A2(n3870), .A3(n3869), .A4(n3868), .ZN(n3877)
         );
  AOI22_X1 U4802 ( .A1(n3987), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4423), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4803 ( .A1(n3640), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4804 ( .A1(n4428), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4805 ( .A1(n3512), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3872) );
  NAND4_X1 U4806 ( .A1(n3875), .A2(n3874), .A3(n3873), .A4(n3872), .ZN(n3876)
         );
  NOR2_X1 U4807 ( .A1(n3877), .A2(n3876), .ZN(n3881) );
  NAND2_X1 U4808 ( .A1(n6505), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3878)
         );
  NAND2_X1 U4809 ( .A1(n4445), .A2(n3878), .ZN(n3879) );
  AOI21_X1 U4810 ( .B1(n4465), .B2(EAX_REG_19__SCAN_IN), .A(n3879), .ZN(n3880)
         );
  OAI21_X1 U4811 ( .B1(n4442), .B2(n3881), .A(n3880), .ZN(n3884) );
  INV_X1 U4812 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3882) );
  XNOR2_X1 U4813 ( .A(n3899), .B(n3882), .ZN(n5780) );
  NAND2_X1 U4814 ( .A1(n5780), .A2(n4439), .ZN(n3883) );
  NAND2_X1 U4815 ( .A1(n3884), .A2(n3883), .ZN(n5380) );
  AOI22_X1 U4816 ( .A1(n3987), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4423), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4817 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3587), .B1(n4388), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4818 ( .A1(n4408), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4819 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4428), .B1(n4403), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3885) );
  NAND4_X1 U4820 ( .A1(n3888), .A2(n3887), .A3(n3886), .A4(n3885), .ZN(n3894)
         );
  AOI22_X1 U4821 ( .A1(n3526), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4822 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n3640), .B1(n3660), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4823 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n3475), .B1(n3506), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4824 ( .A1(n3867), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3498), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3889) );
  NAND4_X1 U4825 ( .A1(n3892), .A2(n3891), .A3(n3890), .A4(n3889), .ZN(n3893)
         );
  NOR2_X1 U4826 ( .A1(n3894), .A2(n3893), .ZN(n3898) );
  OAI21_X1 U4827 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6832), .A(n6505), 
        .ZN(n3895) );
  INV_X1 U4828 ( .A(n3895), .ZN(n3896) );
  AOI21_X1 U4829 ( .B1(n4465), .B2(EAX_REG_20__SCAN_IN), .A(n3896), .ZN(n3897)
         );
  OAI21_X1 U4830 ( .B1(n4442), .B2(n3898), .A(n3897), .ZN(n3904) );
  INV_X1 U4831 ( .A(n3901), .ZN(n3900) );
  INV_X1 U4832 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U4833 ( .A1(n3900), .A2(n5497), .ZN(n3902) );
  AND2_X1 U4834 ( .A1(n3902), .A2(n3918), .ZN(n5768) );
  NAND2_X1 U4835 ( .A1(n5768), .A2(n4395), .ZN(n3903) );
  NAND2_X1 U4836 ( .A1(n5378), .A2(n5498), .ZN(n5371) );
  INV_X1 U4837 ( .A(n5371), .ZN(n3924) );
  AOI22_X1 U4838 ( .A1(n3987), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4423), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4839 ( .A1(n3526), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4840 ( .A1(n3587), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4841 ( .A1(n3867), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3905) );
  NAND4_X1 U4842 ( .A1(n3908), .A2(n3907), .A3(n3906), .A4(n3905), .ZN(n3914)
         );
  AOI22_X1 U4843 ( .A1(n4428), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4844 ( .A1(n4408), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4845 ( .A1(n3475), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4846 ( .A1(n3640), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3498), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3909) );
  NAND4_X1 U4847 ( .A1(n3912), .A2(n3911), .A3(n3910), .A4(n3909), .ZN(n3913)
         );
  NOR2_X1 U4848 ( .A1(n3914), .A2(n3913), .ZN(n3917) );
  INV_X1 U4849 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6864) );
  OAI21_X1 U4850 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6864), .A(n4445), .ZN(
        n3915) );
  AOI21_X1 U4851 ( .B1(n4465), .B2(EAX_REG_21__SCAN_IN), .A(n3915), .ZN(n3916)
         );
  OAI21_X1 U4852 ( .B1(n4442), .B2(n3917), .A(n3916), .ZN(n3922) );
  NOR2_X1 U4853 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n3919), .ZN(n3920)
         );
  NOR2_X1 U4854 ( .A1(n3940), .A2(n3920), .ZN(n5758) );
  NAND2_X1 U4855 ( .A1(n5758), .A2(n4439), .ZN(n3921) );
  NAND2_X1 U4856 ( .A1(n3922), .A2(n3921), .ZN(n5372) );
  NAND2_X1 U4857 ( .A1(n3924), .A2(n3923), .ZN(n5365) );
  AOI22_X1 U4858 ( .A1(n4408), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4859 ( .A1(n3640), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3690), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4860 ( .A1(n4423), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3926) );
  AOI22_X1 U4861 ( .A1(n4428), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3925) );
  NAND4_X1 U4862 ( .A1(n3928), .A2(n3927), .A3(n3926), .A4(n3925), .ZN(n3935)
         );
  AOI22_X1 U4863 ( .A1(n3512), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4864 ( .A1(n3526), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4865 ( .A1(n3987), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4866 ( .A1(n4388), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3498), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3930) );
  NAND4_X1 U4867 ( .A1(n3933), .A2(n3932), .A3(n3931), .A4(n3930), .ZN(n3934)
         );
  NOR2_X1 U4868 ( .A1(n3935), .A2(n3934), .ZN(n3939) );
  NAND2_X1 U4869 ( .A1(n6505), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3936)
         );
  NAND2_X1 U4870 ( .A1(n4445), .A2(n3936), .ZN(n3937) );
  AOI21_X1 U4871 ( .B1(n4465), .B2(EAX_REG_22__SCAN_IN), .A(n3937), .ZN(n3938)
         );
  OAI21_X1 U4872 ( .B1(n4442), .B2(n3939), .A(n3938), .ZN(n3942) );
  OAI21_X1 U4873 ( .B1(n3940), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n3981), 
        .ZN(n5747) );
  OR2_X1 U4874 ( .A1(n5747), .A2(n4445), .ZN(n3941) );
  NAND2_X1 U4875 ( .A1(n3942), .A2(n3941), .ZN(n5367) );
  AOI22_X1 U4876 ( .A1(n4408), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4877 ( .A1(n3526), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4428), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4878 ( .A1(n4423), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4879 ( .A1(n4403), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3943) );
  NAND4_X1 U4880 ( .A1(n3946), .A2(n3945), .A3(n3944), .A4(n3943), .ZN(n3952)
         );
  AOI22_X1 U4881 ( .A1(n4388), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3950) );
  AOI22_X1 U4882 ( .A1(n3512), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4883 ( .A1(n3640), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4884 ( .A1(n3987), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3947) );
  NAND4_X1 U4885 ( .A1(n3950), .A2(n3949), .A3(n3948), .A4(n3947), .ZN(n3951)
         );
  NOR2_X1 U4886 ( .A1(n3952), .A2(n3951), .ZN(n3969) );
  AOI22_X1 U4887 ( .A1(n3987), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4888 ( .A1(n4408), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4889 ( .A1(n3526), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4890 ( .A1(n3640), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3953) );
  NAND4_X1 U4891 ( .A1(n3956), .A2(n3955), .A3(n3954), .A4(n3953), .ZN(n3962)
         );
  AOI22_X1 U4892 ( .A1(n4423), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4893 ( .A1(n4388), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4894 ( .A1(n4428), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4895 ( .A1(n3512), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3957) );
  NAND4_X1 U4896 ( .A1(n3960), .A2(n3959), .A3(n3958), .A4(n3957), .ZN(n3961)
         );
  NOR2_X1 U4897 ( .A1(n3962), .A2(n3961), .ZN(n3970) );
  XOR2_X1 U4898 ( .A(n3969), .B(n3970), .Z(n3963) );
  NAND2_X1 U4899 ( .A1(n3963), .A2(n4415), .ZN(n3968) );
  NAND2_X1 U4900 ( .A1(n6505), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3964)
         );
  NAND2_X1 U4901 ( .A1(n4445), .A2(n3964), .ZN(n3965) );
  AOI21_X1 U4902 ( .B1(n4465), .B2(EAX_REG_23__SCAN_IN), .A(n3965), .ZN(n3967)
         );
  XNOR2_X1 U4903 ( .A(n3981), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5738)
         );
  AND2_X1 U4904 ( .A1(n5738), .A2(n4395), .ZN(n3966) );
  AOI21_X1 U4905 ( .B1(n3968), .B2(n3967), .A(n3966), .ZN(n5357) );
  OR2_X1 U4906 ( .A1(n3970), .A2(n3969), .ZN(n3999) );
  AOI22_X1 U4907 ( .A1(n4408), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3974) );
  INV_X1 U4908 ( .A(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n6987) );
  AOI22_X1 U4909 ( .A1(n3512), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3526), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4910 ( .A1(n4388), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4911 ( .A1(n3987), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3971) );
  NAND4_X1 U4912 ( .A1(n3974), .A2(n3973), .A3(n3972), .A4(n3971), .ZN(n3980)
         );
  AOI22_X1 U4913 ( .A1(n4423), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4914 ( .A1(n3867), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4915 ( .A1(n4428), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4916 ( .A1(n4383), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3975) );
  NAND4_X1 U4917 ( .A1(n3978), .A2(n3977), .A3(n3976), .A4(n3975), .ZN(n3979)
         );
  NOR2_X1 U4918 ( .A1(n3980), .A2(n3979), .ZN(n3998) );
  XNOR2_X1 U4919 ( .A(n3999), .B(n3998), .ZN(n3986) );
  XNOR2_X1 U4920 ( .A(n4005), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5470)
         );
  INV_X1 U4921 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5468) );
  INV_X1 U4922 ( .A(n4464), .ZN(n3983) );
  OAI22_X1 U4923 ( .A1(n5470), .A2(n4445), .B1(n5468), .B2(n3983), .ZN(n3984)
         );
  AOI21_X1 U4924 ( .B1(n4465), .B2(EAX_REG_24__SCAN_IN), .A(n3984), .ZN(n3985)
         );
  OAI21_X1 U4925 ( .B1(n3986), .B2(n4442), .A(n3985), .ZN(n5286) );
  AOI22_X1 U4926 ( .A1(n3987), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U4927 ( .A1(n3526), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3990) );
  AOI22_X1 U4928 ( .A1(n3475), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U4929 ( .A1(n4423), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3988) );
  NAND4_X1 U4930 ( .A1(n3991), .A2(n3990), .A3(n3989), .A4(n3988), .ZN(n3997)
         );
  AOI22_X1 U4931 ( .A1(n3512), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U4932 ( .A1(n3640), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U4933 ( .A1(n4428), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U4934 ( .A1(n4388), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3992) );
  NAND4_X1 U4935 ( .A1(n3995), .A2(n3994), .A3(n3993), .A4(n3992), .ZN(n3996)
         );
  NOR2_X1 U4936 ( .A1(n3997), .A2(n3996), .ZN(n4011) );
  OR2_X1 U4937 ( .A1(n3999), .A2(n3998), .ZN(n4010) );
  XOR2_X1 U4938 ( .A(n4011), .B(n4010), .Z(n4003) );
  INV_X1 U4939 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4001) );
  NAND2_X1 U4940 ( .A1(n6505), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4000)
         );
  OAI211_X1 U4941 ( .C1(n3281), .C2(n4001), .A(n4445), .B(n4000), .ZN(n4002)
         );
  AOI21_X1 U4942 ( .B1(n4003), .B2(n4415), .A(n4002), .ZN(n4004) );
  INV_X1 U4943 ( .A(n4004), .ZN(n4008) );
  XNOR2_X1 U4944 ( .A(n4027), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5459)
         );
  NAND2_X1 U4945 ( .A1(n5459), .A2(n4395), .ZN(n4007) );
  NAND2_X1 U4946 ( .A1(n4008), .A2(n4007), .ZN(n5274) );
  NOR2_X1 U4947 ( .A1(n4011), .A2(n4010), .ZN(n4035) );
  AOI22_X1 U4948 ( .A1(n3987), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U4949 ( .A1(n3526), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U4950 ( .A1(n3475), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3929), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4951 ( .A1(n4423), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4012) );
  NAND4_X1 U4952 ( .A1(n4015), .A2(n4014), .A3(n4013), .A4(n4012), .ZN(n4021)
         );
  AOI22_X1 U4953 ( .A1(n3512), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U4954 ( .A1(n3640), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U4955 ( .A1(n4428), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4956 ( .A1(n4388), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3531), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4016) );
  NAND4_X1 U4957 ( .A1(n4019), .A2(n4018), .A3(n4017), .A4(n4016), .ZN(n4020)
         );
  OR2_X1 U4958 ( .A1(n4021), .A2(n4020), .ZN(n4034) );
  INV_X1 U4959 ( .A(n4034), .ZN(n4022) );
  XNOR2_X1 U4960 ( .A(n4035), .B(n4022), .ZN(n4026) );
  INV_X1 U4961 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4024) );
  NAND2_X1 U4962 ( .A1(n6505), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4023)
         );
  OAI211_X1 U4963 ( .C1(n3281), .C2(n4024), .A(n4445), .B(n4023), .ZN(n4025)
         );
  AOI21_X1 U4964 ( .B1(n4026), .B2(n4415), .A(n4025), .ZN(n4033) );
  INV_X1 U4965 ( .A(n4027), .ZN(n4028) );
  INV_X1 U4966 ( .A(n4029), .ZN(n4030) );
  INV_X1 U4967 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U4968 ( .A1(n4030), .A2(n5452), .ZN(n4031) );
  NAND2_X1 U4969 ( .A1(n4375), .A2(n4031), .ZN(n5451) );
  NOR2_X1 U4970 ( .A1(n5451), .A2(n4445), .ZN(n4032) );
  NOR2_X2 U4971 ( .A1(n5262), .A2(n5263), .ZN(n4052) );
  NAND2_X1 U4972 ( .A1(n4035), .A2(n4034), .ZN(n4381) );
  AOI22_X1 U4973 ( .A1(n4408), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U4974 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3526), .B1(n4388), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4038) );
  AOI22_X1 U4975 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n3640), .B1(n3867), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U4976 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3634), .B1(n3383), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4036) );
  NAND4_X1 U4977 ( .A1(n4039), .A2(n4038), .A3(n4037), .A4(n4036), .ZN(n4045)
         );
  AOI22_X1 U4978 ( .A1(n3987), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4428), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U4979 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3512), .B1(n3660), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U4980 ( .A1(n4423), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U4981 ( .A1(n3392), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3498), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4040) );
  NAND4_X1 U4982 ( .A1(n4043), .A2(n4042), .A3(n4041), .A4(n4040), .ZN(n4044)
         );
  NOR2_X1 U4983 ( .A1(n4045), .A2(n4044), .ZN(n4382) );
  XOR2_X1 U4984 ( .A(n4381), .B(n4382), .Z(n4046) );
  NAND2_X1 U4985 ( .A1(n4046), .A2(n4415), .ZN(n4051) );
  NAND2_X1 U4986 ( .A1(n6505), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4047)
         );
  NAND2_X1 U4987 ( .A1(n4445), .A2(n4047), .ZN(n4048) );
  AOI21_X1 U4988 ( .B1(n4465), .B2(EAX_REG_27__SCAN_IN), .A(n4048), .ZN(n4050)
         );
  XNOR2_X1 U4989 ( .A(n4375), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5254)
         );
  AND2_X1 U4990 ( .A1(n5254), .A2(n4395), .ZN(n4049) );
  NAND3_X1 U4991 ( .A1(n6609), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6625) );
  OR2_X2 U4992 ( .A1(n6625), .A2(n6519), .ZN(n5494) );
  NAND2_X1 U4993 ( .A1(n4055), .A2(n4151), .ZN(n4060) );
  XNOR2_X1 U4994 ( .A(n4070), .B(n4069), .ZN(n4057) );
  OAI211_X1 U4995 ( .C1(n4057), .C2(n6713), .A(n4056), .B(n4167), .ZN(n4058)
         );
  INV_X1 U4996 ( .A(n4058), .ZN(n4059) );
  NAND2_X1 U4997 ( .A1(n4060), .A2(n4059), .ZN(n4580) );
  INV_X1 U4998 ( .A(n5104), .ZN(n4061) );
  NAND2_X1 U4999 ( .A1(n4061), .A2(n4151), .ZN(n4064) );
  NAND2_X1 U5000 ( .A1(n4854), .A2(n3433), .ZN(n4072) );
  OAI21_X1 U5001 ( .B1(n6713), .B2(n4069), .A(n4072), .ZN(n4062) );
  INV_X1 U5002 ( .A(n4062), .ZN(n4063) );
  NAND2_X1 U5003 ( .A1(n4064), .A2(n4063), .ZN(n4553) );
  NAND2_X1 U5004 ( .A1(n4553), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4065)
         );
  INV_X1 U5005 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6848) );
  NAND2_X1 U5006 ( .A1(n4065), .A2(n6848), .ZN(n4066) );
  AND2_X1 U5007 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6191) );
  NAND2_X1 U5008 ( .A1(n4553), .A2(n6191), .ZN(n4067) );
  AND2_X1 U5009 ( .A1(n4066), .A2(n4067), .ZN(n4581) );
  NAND2_X1 U5010 ( .A1(n4580), .A2(n4581), .ZN(n4068) );
  NAND2_X1 U5011 ( .A1(n4068), .A2(n4067), .ZN(n6111) );
  NAND2_X1 U5012 ( .A1(n6111), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4075)
         );
  NAND2_X1 U5013 ( .A1(n4070), .A2(n4069), .ZN(n4080) );
  XNOR2_X1 U5014 ( .A(n4080), .B(n4071), .ZN(n4073) );
  OAI21_X1 U5015 ( .B1(n4073), .B2(n6713), .A(n4072), .ZN(n4074) );
  NAND2_X1 U5016 ( .A1(n4075), .A2(n6109), .ZN(n4078) );
  INV_X1 U5017 ( .A(n6111), .ZN(n4076) );
  NAND2_X1 U5018 ( .A1(n4076), .A2(n6195), .ZN(n4077) );
  AND2_X1 U5019 ( .A1(n4078), .A2(n4077), .ZN(n4618) );
  INV_X1 U5020 ( .A(n4151), .ZN(n4084) );
  NAND2_X1 U5021 ( .A1(n4080), .A2(n4079), .ZN(n4089) );
  INV_X1 U5022 ( .A(n4088), .ZN(n4081) );
  XNOR2_X1 U5023 ( .A(n4089), .B(n4081), .ZN(n4082) );
  NAND2_X1 U5024 ( .A1(n4082), .A2(n3447), .ZN(n4083) );
  OAI21_X2 U5025 ( .B1(n4694), .B2(n4084), .A(n4083), .ZN(n4085) );
  INV_X1 U5026 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6184) );
  XNOR2_X1 U5027 ( .A(n4085), .B(n6184), .ZN(n4619) );
  NAND2_X1 U5028 ( .A1(n4618), .A2(n4619), .ZN(n4620) );
  NAND2_X1 U5029 ( .A1(n4085), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4086)
         );
  NAND2_X1 U5030 ( .A1(n4620), .A2(n4086), .ZN(n6102) );
  NAND2_X1 U5031 ( .A1(n4087), .A2(n4151), .ZN(n4092) );
  NAND2_X1 U5032 ( .A1(n4089), .A2(n4088), .ZN(n4108) );
  XNOR2_X1 U5033 ( .A(n4108), .B(n4106), .ZN(n4090) );
  NAND2_X1 U5034 ( .A1(n4090), .A2(n3447), .ZN(n4091) );
  NAND2_X1 U5035 ( .A1(n4092), .A2(n4091), .ZN(n4093) );
  INV_X1 U5036 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6174) );
  XNOR2_X1 U5037 ( .A(n4093), .B(n6174), .ZN(n6101) );
  NAND2_X1 U5038 ( .A1(n6102), .A2(n6101), .ZN(n6100) );
  NAND2_X1 U5039 ( .A1(n4093), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4094)
         );
  NAND2_X1 U5040 ( .A1(n6100), .A2(n4094), .ZN(n4719) );
  NAND2_X1 U5041 ( .A1(n4095), .A2(n4151), .ZN(n4100) );
  INV_X1 U5042 ( .A(n4106), .ZN(n4096) );
  OR2_X1 U5043 ( .A1(n4108), .A2(n4096), .ZN(n4097) );
  XNOR2_X1 U5044 ( .A(n4097), .B(n4105), .ZN(n4098) );
  NAND2_X1 U5045 ( .A1(n4098), .A2(n3447), .ZN(n4099) );
  NAND2_X1 U5046 ( .A1(n4100), .A2(n4099), .ZN(n4101) );
  INV_X1 U5047 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n7026) );
  XNOR2_X1 U5048 ( .A(n4101), .B(n7026), .ZN(n4718) );
  NAND2_X1 U5049 ( .A1(n4719), .A2(n4718), .ZN(n4717) );
  NAND2_X1 U5050 ( .A1(n4101), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4102)
         );
  NAND2_X1 U5051 ( .A1(n4717), .A2(n4102), .ZN(n6095) );
  NAND3_X1 U5052 ( .A1(n4103), .A2(n4151), .A3(n4104), .ZN(n4111) );
  NAND2_X1 U5053 ( .A1(n4106), .A2(n4105), .ZN(n4107) );
  OR2_X1 U5054 ( .A1(n4108), .A2(n4107), .ZN(n4115) );
  XNOR2_X1 U5055 ( .A(n4115), .B(n4116), .ZN(n4109) );
  NAND2_X1 U5056 ( .A1(n4109), .A2(n3447), .ZN(n4110) );
  NAND2_X1 U5057 ( .A1(n4111), .A2(n4110), .ZN(n4112) );
  INV_X1 U5058 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6166) );
  XNOR2_X1 U5059 ( .A(n4112), .B(n6166), .ZN(n6094) );
  NAND2_X1 U5060 ( .A1(n4112), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4113)
         );
  NAND2_X1 U5061 ( .A1(n4114), .A2(n4151), .ZN(n4120) );
  INV_X1 U5062 ( .A(n4115), .ZN(n4117) );
  NAND2_X1 U5063 ( .A1(n4117), .A2(n4116), .ZN(n4126) );
  XNOR2_X1 U5064 ( .A(n4126), .B(n4127), .ZN(n4118) );
  NAND2_X1 U5065 ( .A1(n4118), .A2(n3447), .ZN(n4119) );
  NAND2_X1 U5066 ( .A1(n4120), .A2(n4119), .ZN(n4121) );
  INV_X1 U5067 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6159) );
  XNOR2_X1 U5068 ( .A(n4121), .B(n6159), .ZN(n4821) );
  NAND2_X1 U5069 ( .A1(n4822), .A2(n4821), .ZN(n4820) );
  NAND2_X1 U5070 ( .A1(n4121), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4122)
         );
  NAND2_X1 U5071 ( .A1(n4820), .A2(n4122), .ZN(n4843) );
  NAND2_X1 U5072 ( .A1(n4151), .A2(n4127), .ZN(n4124) );
  INV_X1 U5073 ( .A(n4126), .ZN(n4128) );
  NAND3_X1 U5074 ( .A1(n4128), .A2(n3447), .A3(n4127), .ZN(n4129) );
  NAND2_X1 U5075 ( .A1(n5534), .A2(n4129), .ZN(n4130) );
  INV_X1 U5076 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6153) );
  XNOR2_X1 U5077 ( .A(n4130), .B(n6153), .ZN(n4842) );
  NAND2_X1 U5078 ( .A1(n4130), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4131)
         );
  INV_X1 U5079 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5089) );
  NAND2_X1 U5080 ( .A1(n5514), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5076)
         );
  OAI21_X1 U5081 ( .B1(n5181), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n5514), 
        .ZN(n4134) );
  NAND3_X1 U5082 ( .A1(n4132), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4133) );
  INV_X1 U5083 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6130) );
  NOR2_X1 U5084 ( .A1(n5534), .A2(n6130), .ZN(n5171) );
  NAND2_X1 U5085 ( .A1(n5534), .A2(n6130), .ZN(n5169) );
  XNOR2_X1 U5086 ( .A(n5534), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5804)
         );
  INV_X1 U5087 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4135) );
  INV_X1 U5088 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n7004) );
  AND2_X1 U5089 ( .A1(n5534), .A2(n7004), .ZN(n5543) );
  NAND2_X1 U5090 ( .A1(n5514), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5544) );
  INV_X1 U5091 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5692) );
  NOR2_X1 U5092 ( .A1(n5534), .A2(n5692), .ZN(n4137) );
  NAND2_X1 U5093 ( .A1(n5534), .A2(n5692), .ZN(n4136) );
  INV_X1 U5094 ( .A(n5512), .ZN(n4139) );
  INV_X1 U5095 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5691) );
  AND2_X1 U5096 ( .A1(n5534), .A2(n5691), .ZN(n5523) );
  NAND2_X1 U5097 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4366) );
  AND2_X1 U5098 ( .A1(n5534), .A2(n4366), .ZN(n4138) );
  NAND2_X1 U5099 ( .A1(n5514), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5524) );
  NOR2_X1 U5100 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4140) );
  NOR2_X1 U5101 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5627) );
  NOR2_X1 U5102 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5608) );
  INV_X1 U5103 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5664) );
  INV_X1 U5104 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6933) );
  NAND2_X1 U5105 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4354) );
  NAND2_X1 U5106 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5625) );
  NOR2_X1 U5107 ( .A1(n4354), .A2(n5625), .ZN(n5605) );
  AND2_X1 U5108 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4359) );
  NAND2_X1 U5109 ( .A1(n5605), .A2(n4359), .ZN(n4368) );
  XOR2_X1 U5110 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(n5534), .Z(n5457) );
  INV_X1 U5111 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6887) );
  INV_X1 U5112 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5592) );
  NOR2_X1 U5113 ( .A1(n5514), .A2(n5592), .ZN(n5449) );
  NOR2_X1 U5114 ( .A1(n5534), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5448)
         );
  NAND2_X1 U5115 ( .A1(n5439), .A2(n4144), .ZN(n4145) );
  INV_X1 U5116 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6797) );
  NAND2_X1 U5117 ( .A1(n3282), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4146) );
  NAND2_X1 U5118 ( .A1(n4147), .A2(n4146), .ZN(n4160) );
  NAND2_X1 U5119 ( .A1(n3223), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4148) );
  XNOR2_X1 U5120 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4153) );
  NOR2_X1 U5121 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6202), .ZN(n4150)
         );
  NAND2_X1 U5122 ( .A1(n4218), .A2(n4171), .ZN(n4197) );
  NOR2_X1 U5123 ( .A1(n4154), .A2(n4153), .ZN(n4155) );
  OR2_X1 U5124 ( .A1(n4156), .A2(n4155), .ZN(n4157) );
  INV_X1 U5125 ( .A(n4217), .ZN(n4159) );
  AOI22_X1 U5126 ( .A1(n4171), .A2(n4159), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6609), .ZN(n4192) );
  NAND2_X1 U5127 ( .A1(n4160), .A2(n4165), .ZN(n4161) );
  NAND2_X1 U5128 ( .A1(n4162), .A2(n4161), .ZN(n4214) );
  NOR2_X1 U5129 ( .A1(n4214), .A2(n6609), .ZN(n4178) );
  NAND2_X1 U5130 ( .A1(n4194), .A2(n3434), .ZN(n4163) );
  NAND2_X1 U5131 ( .A1(n4163), .A2(n4167), .ZN(n4177) );
  NAND2_X1 U5132 ( .A1(n3283), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4164) );
  AND2_X1 U5133 ( .A1(n4165), .A2(n4164), .ZN(n4166) );
  INV_X1 U5134 ( .A(n4166), .ZN(n4170) );
  AOI21_X1 U5135 ( .B1(n3450), .B2(n4166), .A(n4854), .ZN(n4169) );
  NAND2_X1 U5136 ( .A1(n4926), .A2(n4167), .ZN(n4168) );
  NAND2_X1 U5137 ( .A1(n3431), .A2(n4168), .ZN(n4183) );
  OAI22_X1 U5138 ( .A1(n4177), .A2(n4178), .B1(n4169), .B2(n4183), .ZN(n4173)
         );
  NOR3_X1 U5139 ( .A1(n4182), .A2(n4170), .A3(n4173), .ZN(n4176) );
  INV_X1 U5140 ( .A(n4214), .ZN(n4174) );
  INV_X1 U5141 ( .A(n4171), .ZN(n4172) );
  AOI21_X1 U5142 ( .B1(n4174), .B2(n4173), .A(n4172), .ZN(n4175) );
  AOI211_X1 U5143 ( .C1(n4178), .C2(n4177), .A(n4176), .B(n4175), .ZN(n4188)
         );
  OAI21_X1 U5144 ( .B1(n4181), .B2(n4180), .A(n4179), .ZN(n4215) );
  AOI211_X1 U5145 ( .C1(n4190), .C2(n4215), .A(n4184), .B(n4183), .ZN(n4187)
         );
  INV_X1 U5146 ( .A(n4183), .ZN(n4186) );
  INV_X1 U5147 ( .A(n4184), .ZN(n4185) );
  OAI22_X1 U5148 ( .A1(n4188), .A2(n4187), .B1(n4186), .B2(n4185), .ZN(n4189)
         );
  OAI21_X1 U5149 ( .B1(n4190), .B2(n4217), .A(n4189), .ZN(n4191) );
  NAND2_X1 U5150 ( .A1(n4192), .A2(n4191), .ZN(n4193) );
  AOI21_X1 U5151 ( .B1(n5195), .B2(n4854), .A(n3421), .ZN(n4199) );
  NAND2_X1 U5152 ( .A1(n3459), .A2(n4199), .ZN(n4236) );
  NAND2_X1 U5153 ( .A1(n4200), .A2(n6519), .ZN(n4201) );
  NAND2_X1 U5154 ( .A1(n4201), .A2(n6609), .ZN(n4202) );
  NAND2_X1 U5155 ( .A1(n6609), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4204) );
  NAND2_X1 U5156 ( .A1(n6832), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4203) );
  AND2_X1 U5157 ( .A1(n4204), .A2(n4203), .ZN(n4554) );
  INV_X1 U5158 ( .A(n4554), .ZN(n4205) );
  INV_X1 U5159 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4206) );
  NAND2_X1 U5160 ( .A1(n6609), .A2(n6505), .ZN(n6624) );
  INV_X2 U5161 ( .A(n6177), .ZN(n6187) );
  NAND2_X1 U5162 ( .A1(n6187), .A2(REIP_REG_27__SCAN_IN), .ZN(n5581) );
  OAI21_X1 U5163 ( .B1(n5528), .B2(n4206), .A(n5581), .ZN(n4207) );
  OAI21_X1 U5164 ( .B1(n5587), .B2(n6092), .A(n4208), .ZN(n4209) );
  INV_X1 U5165 ( .A(n4209), .ZN(n4210) );
  NAND2_X1 U5166 ( .A1(n3202), .A2(n4210), .ZN(U2959) );
  AND2_X1 U5167 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U5168 ( .A1(n5573), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5553) );
  NOR4_X1 U5169 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A3(INSTADDRPOINTER_REG_28__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4212) );
  NAND2_X1 U5170 ( .A1(n4941), .A2(n3434), .ZN(n4335) );
  NOR2_X1 U5171 ( .A1(n5195), .A2(n4335), .ZN(n4344) );
  INV_X1 U5172 ( .A(n4344), .ZN(n4228) );
  NAND2_X1 U5173 ( .A1(n3279), .A2(n6636), .ZN(n6633) );
  NAND2_X1 U5174 ( .A1(n3434), .A2(n6633), .ZN(n4222) );
  NOR2_X1 U5175 ( .A1(n4215), .A2(n4214), .ZN(n4216) );
  NAND2_X1 U5176 ( .A1(n4217), .A2(n4216), .ZN(n4220) );
  INV_X1 U5177 ( .A(n4218), .ZN(n4219) );
  NAND2_X1 U5178 ( .A1(n4220), .A2(n4219), .ZN(n5211) );
  NOR2_X1 U5179 ( .A1(READY_N), .A2(n5211), .ZN(n4528) );
  NAND3_X1 U5180 ( .A1(n4222), .A2(n4528), .A3(n4221), .ZN(n4227) );
  INV_X1 U5181 ( .A(n4223), .ZN(n5212) );
  NAND2_X1 U5182 ( .A1(n4334), .A2(n4224), .ZN(n4225) );
  OR2_X1 U5183 ( .A1(n4236), .A2(n4225), .ZN(n4226) );
  NAND2_X1 U5184 ( .A1(n5212), .A2(n4226), .ZN(n4523) );
  OAI211_X1 U5185 ( .C1(n5209), .C2(n4228), .A(n4227), .B(n4523), .ZN(n4229)
         );
  NAND2_X1 U5186 ( .A1(n4229), .A2(n6616), .ZN(n4235) );
  NAND2_X1 U5187 ( .A1(n4926), .A2(n6633), .ZN(n4477) );
  INV_X1 U5188 ( .A(READY_N), .ZN(n6635) );
  NAND3_X1 U5189 ( .A1(n4521), .A2(n4477), .A3(n6635), .ZN(n4231) );
  NAND3_X1 U5190 ( .A1(n4231), .A2(n4591), .A3(n4332), .ZN(n4232) );
  NAND2_X1 U5191 ( .A1(n4232), .A2(n4941), .ZN(n4233) );
  NOR2_X1 U5192 ( .A1(n4236), .A2(n3431), .ZN(n4537) );
  INV_X1 U5193 ( .A(n4237), .ZN(n6594) );
  NOR2_X1 U5194 ( .A1(n4537), .A2(n6594), .ZN(n5203) );
  INV_X1 U5195 ( .A(n4238), .ZN(n4529) );
  NAND2_X1 U5196 ( .A1(n4521), .A2(n4295), .ZN(n4560) );
  NAND2_X1 U5197 ( .A1(n4239), .A2(n4240), .ZN(n4241) );
  NAND4_X1 U5198 ( .A1(n5203), .A2(n4238), .A3(n4560), .A4(n4241), .ZN(n4242)
         );
  NAND2_X1 U5199 ( .A1(n4503), .A2(n4243), .ZN(n4374) );
  MUX2_X1 U5200 ( .A(n4318), .B(n5641), .S(EBX_REG_1__SCAN_IN), .Z(n4245) );
  NAND2_X1 U5201 ( .A1(n4601), .A2(n6848), .ZN(n4244) );
  INV_X1 U5202 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4911) );
  OAI22_X1 U5203 ( .A1(n4321), .A2(n4911), .B1(n5641), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n4600) );
  MUX2_X1 U5204 ( .A(n4305), .B(n5382), .S(EBX_REG_2__SCAN_IN), .Z(n4248) );
  NOR2_X1 U5205 ( .A1(n4327), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4247)
         );
  NOR2_X1 U5206 ( .A1(n4248), .A2(n4247), .ZN(n4593) );
  INV_X1 U5207 ( .A(n4690), .ZN(n4254) );
  NAND2_X1 U5208 ( .A1(n4321), .A2(n6184), .ZN(n4249) );
  OAI211_X1 U5209 ( .C1(n3190), .C2(EBX_REG_3__SCAN_IN), .A(n4249), .B(n5641), 
        .ZN(n4252) );
  INV_X1 U5210 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4250) );
  NAND2_X1 U5211 ( .A1(n5382), .A2(n4250), .ZN(n4251) );
  MUX2_X1 U5212 ( .A(n4318), .B(n5641), .S(EBX_REG_4__SCAN_IN), .Z(n4256) );
  NAND2_X1 U5213 ( .A1(n4601), .A2(n6174), .ZN(n4255) );
  NAND2_X1 U5214 ( .A1(n4256), .A2(n4255), .ZN(n4710) );
  NAND2_X1 U5215 ( .A1(n4321), .A2(n7026), .ZN(n4257) );
  OAI211_X1 U5216 ( .C1(n3190), .C2(EBX_REG_5__SCAN_IN), .A(n4257), .B(n5641), 
        .ZN(n4260) );
  INV_X1 U5217 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4258) );
  NAND2_X1 U5218 ( .A1(n5382), .A2(n4258), .ZN(n4259) );
  NAND2_X1 U5219 ( .A1(n4260), .A2(n4259), .ZN(n4713) );
  MUX2_X1 U5220 ( .A(n4318), .B(n5641), .S(EBX_REG_6__SCAN_IN), .Z(n4262) );
  NAND2_X1 U5221 ( .A1(n4601), .A2(n6166), .ZN(n4261) );
  NAND2_X1 U5222 ( .A1(n4262), .A2(n4261), .ZN(n4751) );
  NAND2_X1 U5223 ( .A1(n4321), .A2(n6159), .ZN(n4263) );
  OAI211_X1 U5224 ( .C1(n3190), .C2(EBX_REG_7__SCAN_IN), .A(n4263), .B(n5641), 
        .ZN(n4265) );
  INV_X1 U5225 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6871) );
  NAND2_X1 U5226 ( .A1(n5382), .A2(n6871), .ZN(n4264) );
  MUX2_X1 U5227 ( .A(n4305), .B(n5382), .S(EBX_REG_8__SCAN_IN), .Z(n4267) );
  NOR2_X1 U5228 ( .A1(n4327), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4266)
         );
  NOR2_X1 U5229 ( .A1(n4267), .A2(n4266), .ZN(n4829) );
  MUX2_X1 U5230 ( .A(n5382), .B(n4450), .S(EBX_REG_9__SCAN_IN), .Z(n4268) );
  INV_X1 U5231 ( .A(n4268), .ZN(n4270) );
  NAND2_X1 U5232 ( .A1(n3190), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4269)
         );
  NAND2_X1 U5233 ( .A1(n4270), .A2(n4269), .ZN(n4837) );
  INV_X1 U5234 ( .A(EBX_REG_10__SCAN_IN), .ZN(n7014) );
  NAND2_X1 U5235 ( .A1(n4305), .A2(n7014), .ZN(n4274) );
  NAND2_X1 U5236 ( .A1(n5641), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4272) );
  OAI211_X1 U5237 ( .C1(n3190), .C2(EBX_REG_10__SCAN_IN), .A(n4321), .B(n4272), 
        .ZN(n4273) );
  NAND2_X1 U5238 ( .A1(n4274), .A2(n4273), .ZN(n4853) );
  MUX2_X1 U5239 ( .A(n5382), .B(n4450), .S(EBX_REG_11__SCAN_IN), .Z(n4276) );
  AND2_X1 U5240 ( .A1(n3190), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4275)
         );
  NOR2_X1 U5241 ( .A1(n4276), .A2(n4275), .ZN(n5026) );
  INV_X1 U5242 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5165) );
  NAND2_X1 U5243 ( .A1(n4305), .A2(n5165), .ZN(n4279) );
  NAND2_X1 U5244 ( .A1(n5641), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4277) );
  OAI211_X1 U5245 ( .C1(n3190), .C2(EBX_REG_12__SCAN_IN), .A(n4321), .B(n4277), 
        .ZN(n4278) );
  MUX2_X1 U5246 ( .A(n5382), .B(n4450), .S(EBX_REG_13__SCAN_IN), .Z(n4281) );
  AND2_X1 U5247 ( .A1(n3190), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4280)
         );
  NOR2_X1 U5248 ( .A1(n4281), .A2(n4280), .ZN(n5712) );
  INV_X1 U5249 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5983) );
  NAND2_X1 U5250 ( .A1(n4305), .A2(n5983), .ZN(n4284) );
  NAND2_X1 U5251 ( .A1(n5641), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4282) );
  OAI211_X1 U5252 ( .C1(n3190), .C2(EBX_REG_14__SCAN_IN), .A(n4321), .B(n4282), 
        .ZN(n4283) );
  NAND2_X1 U5253 ( .A1(n4284), .A2(n4283), .ZN(n5713) );
  NOR2_X1 U5254 ( .A1(n5712), .A2(n5713), .ZN(n4285) );
  MUX2_X1 U5255 ( .A(n5382), .B(n4450), .S(EBX_REG_15__SCAN_IN), .Z(n4287) );
  AND2_X1 U5256 ( .A1(n3190), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4286)
         );
  NOR2_X1 U5257 ( .A1(n4287), .A2(n4286), .ZN(n5315) );
  INV_X1 U5258 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U5259 ( .A1(n4305), .A2(n5307), .ZN(n4290) );
  NAND2_X1 U5260 ( .A1(n5641), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4288) );
  OAI211_X1 U5261 ( .C1(n3190), .C2(EBX_REG_16__SCAN_IN), .A(n4321), .B(n4288), 
        .ZN(n4289) );
  NAND2_X1 U5262 ( .A1(n4290), .A2(n4289), .ZN(n5300) );
  MUX2_X1 U5263 ( .A(n5382), .B(n4450), .S(EBX_REG_17__SCAN_IN), .Z(n4292) );
  AND2_X1 U5264 ( .A1(n3190), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4291)
         );
  NOR2_X1 U5265 ( .A1(n4292), .A2(n4291), .ZN(n5684) );
  MUX2_X1 U5266 ( .A(n4305), .B(n5382), .S(EBX_REG_19__SCAN_IN), .Z(n4294) );
  NOR2_X1 U5267 ( .A1(n4327), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4293)
         );
  NOR2_X1 U5268 ( .A1(n4294), .A2(n4293), .ZN(n5385) );
  OAI22_X1 U5269 ( .A1(n4327), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n3190), .ZN(n5643) );
  INV_X1 U5270 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5675) );
  NAND2_X1 U5271 ( .A1(n4601), .A2(n5675), .ZN(n4297) );
  INV_X1 U5272 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5383) );
  NAND2_X1 U5273 ( .A1(n4295), .A2(n5383), .ZN(n4296) );
  NAND2_X1 U5274 ( .A1(n4297), .A2(n4296), .ZN(n5642) );
  INV_X1 U5275 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U5276 ( .A1(n5642), .A2(n5788), .ZN(n4298) );
  OAI21_X1 U5277 ( .B1(n5643), .B2(n5382), .A(n4298), .ZN(n4300) );
  NAND2_X1 U5278 ( .A1(n5642), .A2(n5641), .ZN(n4299) );
  NAND2_X1 U5279 ( .A1(n4300), .A2(n4299), .ZN(n4301) );
  MUX2_X1 U5280 ( .A(n4318), .B(n5641), .S(EBX_REG_21__SCAN_IN), .Z(n4302) );
  OAI21_X1 U5281 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n4327), .A(n4302), 
        .ZN(n5375) );
  MUX2_X1 U5282 ( .A(n5382), .B(n4450), .S(EBX_REG_22__SCAN_IN), .Z(n4304) );
  AND2_X1 U5283 ( .A1(n3190), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4303)
         );
  NOR2_X1 U5284 ( .A1(n4304), .A2(n4303), .ZN(n5358) );
  INV_X1 U5285 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6939) );
  NAND2_X1 U5286 ( .A1(n4305), .A2(n6939), .ZN(n4308) );
  NAND2_X1 U5287 ( .A1(n5641), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4306) );
  OAI211_X1 U5288 ( .C1(n3190), .C2(EBX_REG_23__SCAN_IN), .A(n4321), .B(n4306), 
        .ZN(n4307) );
  NAND2_X1 U5289 ( .A1(n4308), .A2(n4307), .ZN(n5359) );
  NOR2_X1 U5290 ( .A1(n5358), .A2(n5359), .ZN(n4309) );
  INV_X1 U5291 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U5292 ( .A1(n4321), .A2(n5609), .ZN(n4310) );
  OAI211_X1 U5293 ( .C1(n3190), .C2(EBX_REG_24__SCAN_IN), .A(n4310), .B(n5641), 
        .ZN(n4312) );
  INV_X1 U5294 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5292) );
  NAND2_X1 U5295 ( .A1(n5382), .A2(n5292), .ZN(n4311) );
  NAND2_X1 U5296 ( .A1(n4312), .A2(n4311), .ZN(n5288) );
  MUX2_X1 U5297 ( .A(n4318), .B(n5641), .S(EBX_REG_25__SCAN_IN), .Z(n4314) );
  NAND2_X1 U5298 ( .A1(n4601), .A2(n6887), .ZN(n4313) );
  NAND2_X1 U5299 ( .A1(n4314), .A2(n4313), .ZN(n5275) );
  NAND2_X1 U5300 ( .A1(n4321), .A2(n5592), .ZN(n4315) );
  OAI211_X1 U5301 ( .C1(n3190), .C2(EBX_REG_26__SCAN_IN), .A(n4315), .B(n5641), 
        .ZN(n4317) );
  INV_X1 U5302 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U5303 ( .A1(n5382), .A2(n5352), .ZN(n4316) );
  MUX2_X1 U5304 ( .A(n4318), .B(n5641), .S(EBX_REG_27__SCAN_IN), .Z(n4320) );
  NAND2_X1 U5305 ( .A1(n4601), .A2(n6797), .ZN(n4319) );
  NAND2_X1 U5306 ( .A1(n4320), .A2(n4319), .ZN(n5251) );
  INV_X1 U5307 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U5308 ( .A1(n4321), .A2(n5441), .ZN(n4322) );
  OAI211_X1 U5309 ( .C1(n3190), .C2(EBX_REG_28__SCAN_IN), .A(n4322), .B(n5641), 
        .ZN(n4324) );
  INV_X1 U5310 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5350) );
  NAND2_X1 U5311 ( .A1(n5382), .A2(n5350), .ZN(n4323) );
  NAND2_X1 U5312 ( .A1(n4324), .A2(n4323), .ZN(n5235) );
  OAI22_X1 U5313 ( .A1(n4327), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        EBX_REG_29__SCAN_IN), .B2(n3190), .ZN(n5225) );
  NOR2_X1 U5314 ( .A1(n5641), .A2(EBX_REG_29__SCAN_IN), .ZN(n5223) );
  INV_X1 U5315 ( .A(n5237), .ZN(n4454) );
  AOI22_X1 U5316 ( .A1(n4457), .A2(n5641), .B1(n5223), .B2(n4454), .ZN(n5227)
         );
  NAND2_X1 U5317 ( .A1(n4327), .A2(EBX_REG_30__SCAN_IN), .ZN(n4326) );
  NAND2_X1 U5318 ( .A1(n3190), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4325) );
  NAND2_X1 U5319 ( .A1(n4326), .A2(n4325), .ZN(n4456) );
  INV_X1 U5320 ( .A(n4457), .ZN(n4455) );
  NAND2_X1 U5321 ( .A1(n4455), .A2(n5641), .ZN(n4460) );
  OAI21_X1 U5322 ( .B1(n5227), .B2(n4456), .A(n4460), .ZN(n4329) );
  AOI22_X1 U5323 ( .A1(n4327), .A2(EBX_REG_31__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n3190), .ZN(n4328) );
  XNOR2_X1 U5324 ( .A(n4329), .B(n4328), .ZN(n5347) );
  INV_X1 U5325 ( .A(n5347), .ZN(n4372) );
  NAND2_X1 U5326 ( .A1(n4521), .A2(n3447), .ZN(n6604) );
  NAND2_X1 U5327 ( .A1(n4239), .A2(n3455), .ZN(n4330) );
  NAND2_X1 U5328 ( .A1(n6604), .A2(n4330), .ZN(n4331) );
  OAI21_X1 U5329 ( .B1(n4591), .B2(n4332), .A(n4221), .ZN(n4333) );
  AND2_X1 U5330 ( .A1(n4334), .A2(n4333), .ZN(n4338) );
  NAND2_X1 U5331 ( .A1(n4601), .A2(n4335), .ZN(n4336) );
  NAND2_X1 U5332 ( .A1(n4336), .A2(n3421), .ZN(n4337) );
  OAI211_X1 U5333 ( .C1(n3459), .C2(n5641), .A(n4338), .B(n4337), .ZN(n4339)
         );
  INV_X1 U5334 ( .A(n4339), .ZN(n4340) );
  NAND2_X1 U5335 ( .A1(n3200), .A2(n4340), .ZN(n4511) );
  OAI21_X1 U5336 ( .B1(n4513), .B2(n4591), .A(n4341), .ZN(n4342) );
  NOR2_X1 U5337 ( .A1(n4511), .A2(n4342), .ZN(n4345) );
  INV_X1 U5338 ( .A(n4345), .ZN(n4343) );
  NAND2_X1 U5339 ( .A1(n4345), .A2(n4344), .ZN(n5204) );
  INV_X1 U5340 ( .A(n5204), .ZN(n4346) );
  NAND2_X1 U5341 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4364) );
  INV_X1 U5342 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4545) );
  INV_X1 U5343 ( .A(n6190), .ZN(n4360) );
  INV_X1 U5344 ( .A(n5703), .ZN(n4347) );
  NAND2_X1 U5345 ( .A1(n4360), .A2(n4347), .ZN(n5707) );
  NAND2_X1 U5346 ( .A1(n4545), .A2(n5707), .ZN(n4610) );
  INV_X1 U5347 ( .A(n4610), .ZN(n4349) );
  NOR2_X1 U5348 ( .A1(n4348), .A2(n6187), .ZN(n4604) );
  NOR2_X1 U5349 ( .A1(n4349), .A2(n4604), .ZN(n4732) );
  NAND2_X1 U5350 ( .A1(n4732), .A2(n4360), .ZN(n5646) );
  NAND3_X1 U5351 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5710) );
  NOR2_X1 U5352 ( .A1(n7004), .A2(n5710), .ZN(n5693) );
  NAND2_X1 U5353 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5699) );
  INV_X1 U5354 ( .A(n5699), .ZN(n4350) );
  NAND2_X1 U5355 ( .A1(n5693), .A2(n4350), .ZN(n5647) );
  NOR2_X1 U5356 ( .A1(n6159), .A2(n6153), .ZN(n6148) );
  INV_X1 U5357 ( .A(n6148), .ZN(n5088) );
  NAND2_X1 U5358 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6138) );
  OR2_X1 U5359 ( .A1(n5088), .A2(n6138), .ZN(n4353) );
  NOR2_X1 U5360 ( .A1(n6184), .A2(n6174), .ZN(n4351) );
  INV_X1 U5361 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6195) );
  NOR2_X1 U5362 ( .A1(n6195), .A2(n6848), .ZN(n5086) );
  NAND4_X1 U5363 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n4351), .A4(n5086), .ZN(n5083) );
  NOR2_X1 U5364 ( .A1(n4353), .A2(n5083), .ZN(n4365) );
  INV_X1 U5365 ( .A(n4365), .ZN(n5826) );
  OR2_X1 U5366 ( .A1(n5647), .A2(n5826), .ZN(n5648) );
  AOI21_X1 U5367 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6192) );
  INV_X1 U5368 ( .A(n4351), .ZN(n6170) );
  NOR2_X1 U5369 ( .A1(n6192), .A2(n6170), .ZN(n4730) );
  NAND2_X1 U5370 ( .A1(n6190), .A2(n4730), .ZN(n4734) );
  NAND2_X1 U5371 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4352) );
  OAI22_X1 U5372 ( .A1(n5646), .A2(n5648), .B1(n5706), .B2(n5647), .ZN(n4355)
         );
  NOR2_X1 U5373 ( .A1(n4366), .A2(n4354), .ZN(n5624) );
  NAND2_X1 U5374 ( .A1(n4355), .A2(n5624), .ZN(n4357) );
  OR2_X1 U5375 ( .A1(n5646), .A2(n5653), .ZN(n4356) );
  NAND2_X1 U5376 ( .A1(n4357), .A2(n4356), .ZN(n5622) );
  NAND2_X1 U5377 ( .A1(n4733), .A2(n5625), .ZN(n4358) );
  NAND2_X1 U5378 ( .A1(n5622), .A2(n4358), .ZN(n5619) );
  INV_X1 U5379 ( .A(n6196), .ZN(n4361) );
  AOI21_X1 U5380 ( .B1(n4361), .B2(n4360), .A(n4359), .ZN(n4362) );
  NAND2_X1 U5381 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5590) );
  AND2_X1 U5382 ( .A1(n4733), .A2(n5590), .ZN(n4363) );
  NOR2_X1 U5383 ( .A1(n5606), .A2(n4363), .ZN(n5583) );
  OAI21_X1 U5384 ( .B1(n5573), .B2(n5694), .A(n5583), .ZN(n5567) );
  AOI21_X1 U5385 ( .B1(n4733), .B2(n4364), .A(n5567), .ZN(n5557) );
  NAND2_X1 U5386 ( .A1(n6187), .A2(REIP_REG_31__SCAN_IN), .ZN(n4500) );
  NAND2_X1 U5387 ( .A1(n6196), .A2(n4365), .ZN(n6123) );
  NAND2_X1 U5388 ( .A1(n5706), .A2(n6123), .ZN(n6129) );
  NAND2_X1 U5389 ( .A1(n5693), .A2(n6129), .ZN(n5823) );
  INV_X1 U5390 ( .A(n4366), .ZN(n4367) );
  NAND2_X1 U5391 ( .A1(n5689), .A2(n4367), .ZN(n5604) );
  INV_X1 U5392 ( .A(n5553), .ZN(n4369) );
  NAND4_X1 U5393 ( .A1(n5585), .A2(n4369), .A3(INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n4213), .ZN(n4370) );
  OAI211_X1 U5394 ( .C1(n5557), .C2(n4213), .A(n4500), .B(n4370), .ZN(n4371)
         );
  AOI21_X1 U5395 ( .B1(n4372), .B2(n6189), .A(n4371), .ZN(n4373) );
  NAND2_X1 U5396 ( .A1(n4374), .A2(n4373), .ZN(U2987) );
  INV_X1 U5397 ( .A(n4375), .ZN(n4376) );
  INV_X1 U5398 ( .A(n4377), .ZN(n4379) );
  INV_X1 U5399 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4378) );
  NAND2_X1 U5400 ( .A1(n4379), .A2(n4378), .ZN(n4380) );
  NAND2_X1 U5401 ( .A1(n4421), .A2(n4380), .ZN(n5444) );
  NOR2_X1 U5402 ( .A1(n4382), .A2(n4381), .ZN(n4402) );
  AOI22_X1 U5403 ( .A1(n3987), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4387) );
  AOI22_X1 U5404 ( .A1(n3526), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4383), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4386) );
  AOI22_X1 U5405 ( .A1(n3475), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3383), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4385) );
  AOI22_X1 U5406 ( .A1(n4423), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4384) );
  NAND4_X1 U5407 ( .A1(n4387), .A2(n4386), .A3(n4385), .A4(n4384), .ZN(n4394)
         );
  AOI22_X1 U5408 ( .A1(n3587), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4392) );
  AOI22_X1 U5409 ( .A1(n3640), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4391) );
  AOI22_X1 U5410 ( .A1(n4428), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4390) );
  AOI22_X1 U5411 ( .A1(n4388), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3498), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4389) );
  NAND4_X1 U5412 ( .A1(n4392), .A2(n4391), .A3(n4390), .A4(n4389), .ZN(n4393)
         );
  OR2_X1 U5413 ( .A1(n4394), .A2(n4393), .ZN(n4401) );
  XNOR2_X1 U5414 ( .A(n4402), .B(n4401), .ZN(n4398) );
  AOI21_X1 U5415 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6505), .A(n4395), 
        .ZN(n4397) );
  NAND2_X1 U5416 ( .A1(n4465), .A2(EAX_REG_28__SCAN_IN), .ZN(n4396) );
  OAI211_X1 U5417 ( .C1(n4398), .C2(n4442), .A(n4397), .B(n4396), .ZN(n4399)
         );
  NAND2_X1 U5418 ( .A1(n4402), .A2(n4401), .ZN(n4435) );
  AOI22_X1 U5419 ( .A1(n3987), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3526), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4407) );
  AOI22_X1 U5420 ( .A1(n3512), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4406) );
  AOI22_X1 U5421 ( .A1(n4423), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4405) );
  AOI22_X1 U5422 ( .A1(n3867), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4404) );
  NAND4_X1 U5423 ( .A1(n4407), .A2(n4406), .A3(n4405), .A4(n4404), .ZN(n4414)
         );
  AOI22_X1 U5424 ( .A1(n4408), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3475), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4412) );
  AOI22_X1 U5425 ( .A1(n4428), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4411) );
  AOI22_X1 U5426 ( .A1(n3634), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3383), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4410) );
  AOI22_X1 U5427 ( .A1(n3660), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3498), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4409) );
  NAND4_X1 U5428 ( .A1(n4412), .A2(n4411), .A3(n4410), .A4(n4409), .ZN(n4413)
         );
  NOR2_X1 U5429 ( .A1(n4414), .A2(n4413), .ZN(n4436) );
  XOR2_X1 U5430 ( .A(n4435), .B(n4436), .Z(n4416) );
  NAND2_X1 U5431 ( .A1(n4416), .A2(n4415), .ZN(n4420) );
  INV_X1 U5432 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4417) );
  AOI21_X1 U5433 ( .B1(n4417), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4418) );
  AOI21_X1 U5434 ( .B1(n4465), .B2(EAX_REG_29__SCAN_IN), .A(n4418), .ZN(n4419)
         );
  XNOR2_X1 U5435 ( .A(n4421), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5433)
         );
  INV_X1 U5436 ( .A(n4421), .ZN(n4422) );
  XNOR2_X1 U5437 ( .A(n4472), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5426)
         );
  AOI22_X1 U5438 ( .A1(n4423), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4408), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4427) );
  AOI22_X1 U5439 ( .A1(n3475), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3634), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4426) );
  AOI22_X1 U5440 ( .A1(n3640), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3660), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4425) );
  AOI22_X1 U5441 ( .A1(n4388), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3498), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4424) );
  NAND4_X1 U5442 ( .A1(n4427), .A2(n4426), .A3(n4425), .A4(n4424), .ZN(n4434)
         );
  AOI22_X1 U5443 ( .A1(n3512), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4432) );
  AOI22_X1 U5444 ( .A1(n3987), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3506), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4431) );
  AOI22_X1 U5445 ( .A1(n3526), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3383), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4430) );
  AOI22_X1 U5446 ( .A1(n4428), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4429) );
  NAND4_X1 U5447 ( .A1(n4432), .A2(n4431), .A3(n4430), .A4(n4429), .ZN(n4433)
         );
  NOR2_X1 U5448 ( .A1(n4434), .A2(n4433), .ZN(n4438) );
  NOR2_X1 U5449 ( .A1(n4436), .A2(n4435), .ZN(n4437) );
  XOR2_X1 U5450 ( .A(n4438), .B(n4437), .Z(n4443) );
  AOI21_X1 U5451 ( .B1(PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6505), .A(n4439), 
        .ZN(n4441) );
  NAND2_X1 U5452 ( .A1(n4465), .A2(EAX_REG_30__SCAN_IN), .ZN(n4440) );
  OAI211_X1 U5453 ( .C1(n4443), .C2(n4442), .A(n4441), .B(n4440), .ZN(n4444)
         );
  INV_X1 U5454 ( .A(n5428), .ZN(n5393) );
  OR2_X1 U5455 ( .A1(n5204), .A2(n5209), .ZN(n4527) );
  INV_X1 U5456 ( .A(n3428), .ZN(n5189) );
  NAND3_X1 U5457 ( .A1(n3455), .A2(n4941), .A3(n5189), .ZN(n4449) );
  OR2_X1 U5458 ( .A1(n4449), .A2(n4448), .ZN(n4647) );
  INV_X1 U5459 ( .A(n4647), .ZN(n4451) );
  NAND3_X1 U5460 ( .A1(n4451), .A2(n4450), .A3(n3434), .ZN(n4452) );
  NAND2_X1 U5461 ( .A1(n4527), .A2(n4452), .ZN(n4453) );
  AOI21_X1 U5462 ( .B1(n4455), .B2(n4454), .A(n4456), .ZN(n4461) );
  INV_X1 U5463 ( .A(n4456), .ZN(n4458) );
  AOI211_X1 U5464 ( .C1(n5382), .C2(n5237), .A(n4458), .B(n4457), .ZN(n4459)
         );
  INV_X1 U5465 ( .A(EBX_REG_30__SCAN_IN), .ZN(n6860) );
  INV_X1 U5466 ( .A(n4462), .ZN(n4463) );
  AOI22_X1 U5467 ( .A1(n4465), .A2(EAX_REG_31__SCAN_IN), .B1(n4464), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4466) );
  INV_X1 U5468 ( .A(n5211), .ZN(n4470) );
  AND2_X1 U5469 ( .A1(n4223), .A2(n6616), .ZN(n4469) );
  NAND2_X1 U5470 ( .A1(n4470), .A2(n4469), .ZN(n5736) );
  NOR2_X1 U5471 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6714) );
  NOR3_X1 U5472 ( .A1(n6609), .A2(n4054), .A3(n6611), .ZN(n6607) );
  OR3_X1 U5473 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n6624), .A3(n6858), .ZN(n6620) );
  NAND2_X1 U5474 ( .A1(n6177), .A2(n6620), .ZN(n4471) );
  INV_X1 U5475 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5216) );
  INV_X1 U5476 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4491) );
  NOR2_X1 U5477 ( .A1(n4862), .A2(n6858), .ZN(n4475) );
  NAND2_X1 U5478 ( .A1(n5191), .A2(n5929), .ZN(n4498) );
  NOR2_X1 U5479 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6601) );
  INV_X1 U5480 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5346) );
  NOR2_X1 U5481 ( .A1(n3190), .A2(n5346), .ZN(n4476) );
  NAND2_X1 U5482 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5752) );
  NAND3_X1 U5483 ( .A1(n4477), .A2(n4591), .A3(n6601), .ZN(n4478) );
  INV_X1 U5484 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6671) );
  INV_X1 U5485 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6666) );
  INV_X1 U5486 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6662) );
  INV_X1 U5487 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6661) );
  INV_X1 U5488 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6657) );
  INV_X1 U5489 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6647) );
  NAND2_X1 U5490 ( .A1(REIP_REG_3__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .ZN(
        n5931) );
  NOR2_X1 U5491 ( .A1(n6647), .A2(n5931), .ZN(n4987) );
  NAND3_X1 U5492 ( .A1(REIP_REG_4__SCAN_IN), .A2(REIP_REG_5__SCAN_IN), .A3(
        n4987), .ZN(n5333) );
  NAND2_X1 U5493 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .ZN(
        n5339) );
  NOR3_X1 U5494 ( .A1(n6657), .A2(n5333), .A3(n5339), .ZN(n4864) );
  NAND2_X1 U5495 ( .A1(REIP_REG_9__SCAN_IN), .A2(n4864), .ZN(n4865) );
  NOR2_X1 U5496 ( .A1(n6661), .A2(n4865), .ZN(n5906) );
  NAND2_X1 U5497 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5906), .ZN(n5157) );
  NOR2_X1 U5498 ( .A1(n6662), .A2(n5157), .ZN(n5893) );
  NAND2_X1 U5499 ( .A1(REIP_REG_13__SCAN_IN), .A2(n5893), .ZN(n5883) );
  NOR2_X1 U5500 ( .A1(n6666), .A2(n5883), .ZN(n5302) );
  NAND4_X1 U5501 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5302), .A3(
        REIP_REG_16__SCAN_IN), .A4(REIP_REG_15__SCAN_IN), .ZN(n5868) );
  NOR2_X1 U5502 ( .A1(n6671), .A2(n5868), .ZN(n5781) );
  NAND2_X1 U5503 ( .A1(REIP_REG_19__SCAN_IN), .A2(n5781), .ZN(n4479) );
  NAND2_X1 U5504 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5767), .ZN(n5751) );
  NOR2_X1 U5505 ( .A1(n5752), .A2(n5751), .ZN(n5742) );
  NAND2_X1 U5506 ( .A1(REIP_REG_23__SCAN_IN), .A2(n5742), .ZN(n5293) );
  NAND3_X1 U5507 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5243) );
  NOR2_X1 U5508 ( .A1(n5293), .A2(n5243), .ZN(n5259) );
  NAND3_X1 U5509 ( .A1(n5259), .A2(REIP_REG_28__SCAN_IN), .A3(
        REIP_REG_27__SCAN_IN), .ZN(n5228) );
  NAND2_X1 U5510 ( .A1(REIP_REG_30__SCAN_IN), .A2(REIP_REG_29__SCAN_IN), .ZN(
        n4492) );
  INV_X1 U5511 ( .A(n4492), .ZN(n4488) );
  INV_X1 U5512 ( .A(n4479), .ZN(n4480) );
  NAND2_X1 U5513 ( .A1(REIP_REG_20__SCAN_IN), .A2(n4480), .ZN(n4481) );
  NAND2_X1 U5514 ( .A1(n5963), .A2(n4481), .ZN(n4482) );
  NAND2_X1 U5515 ( .A1(n4482), .A2(n5773), .ZN(n5766) );
  INV_X1 U5516 ( .A(n5766), .ZN(n4484) );
  INV_X1 U5517 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6677) );
  INV_X1 U5518 ( .A(n5773), .ZN(n5959) );
  OR2_X1 U5519 ( .A1(n5963), .A2(n5959), .ZN(n4914) );
  OAI21_X1 U5520 ( .B1(n5752), .B2(n6677), .A(n4914), .ZN(n4483) );
  NAND2_X1 U5521 ( .A1(n4484), .A2(n4483), .ZN(n5743) );
  AND2_X1 U5522 ( .A1(n5963), .A2(n5243), .ZN(n4485) );
  OR2_X1 U5523 ( .A1(n5743), .A2(n4485), .ZN(n5268) );
  AND2_X1 U5524 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4486) );
  NOR2_X1 U5525 ( .A1(n5932), .A2(n4486), .ZN(n4487) );
  NOR2_X1 U5526 ( .A1(n5268), .A2(n4487), .ZN(n5241) );
  OAI21_X1 U5527 ( .B1(n5228), .B2(n4488), .A(n5241), .ZN(n5218) );
  INV_X1 U5528 ( .A(n6601), .ZN(n4489) );
  OAI21_X1 U5529 ( .B1(n6633), .B2(n4489), .A(n3447), .ZN(n4490) );
  OR2_X1 U5530 ( .A1(n4907), .A2(n4490), .ZN(n4857) );
  OAI22_X1 U5531 ( .A1(n5934), .A2(n4491), .B1(n4857), .B2(n5346), .ZN(n4494)
         );
  NOR3_X1 U5532 ( .A1(n5228), .A2(REIP_REG_31__SCAN_IN), .A3(n4492), .ZN(n4493) );
  AOI211_X1 U5533 ( .C1(REIP_REG_31__SCAN_IN), .C2(n5218), .A(n4494), .B(n4493), .ZN(n4495) );
  NAND2_X1 U5534 ( .A1(n4498), .A2(n4497), .ZN(U2796) );
  NAND2_X1 U5535 ( .A1(n6108), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4499)
         );
  OAI211_X1 U5536 ( .C1(n6117), .C2(n4862), .A(n4500), .B(n4499), .ZN(n4501)
         );
  AOI21_X1 U5537 ( .B1(n5191), .B2(n6113), .A(n4501), .ZN(n4505) );
  NAND2_X1 U5538 ( .A1(n4503), .A2(n4502), .ZN(n4504) );
  NAND2_X1 U5539 ( .A1(n4505), .A2(n4504), .ZN(U2955) );
  INV_X1 U5540 ( .A(n6711), .ZN(n4507) );
  NAND2_X1 U5541 ( .A1(n6713), .A2(n3449), .ZN(n5215) );
  OR2_X1 U5542 ( .A1(n6519), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5846) );
  INV_X1 U5543 ( .A(n5846), .ZN(n4859) );
  OAI21_X1 U5544 ( .B1(n4859), .B2(READREQUEST_REG_SCAN_IN), .A(n4507), .ZN(
        n4506) );
  OAI21_X1 U5545 ( .B1(n4507), .B2(n5215), .A(n4506), .ZN(U3474) );
  AOI22_X1 U5546 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4213), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6848), .ZN(n4544) );
  NOR2_X1 U5547 ( .A1(n6858), .A2(n4545), .ZN(n4520) );
  INV_X1 U5548 ( .A(n4511), .ZN(n4515) );
  AND4_X1 U5549 ( .A1(n4238), .A2(n4513), .A3(n4230), .A4(n4512), .ZN(n4514)
         );
  NAND2_X1 U5550 ( .A1(n4515), .A2(n4514), .ZN(n4656) );
  INV_X1 U5551 ( .A(n4656), .ZN(n5196) );
  NOR3_X1 U5552 ( .A1(n5195), .A2(n4516), .A3(n4517), .ZN(n4518) );
  AOI21_X1 U5553 ( .B1(n6581), .B2(n3282), .A(n4518), .ZN(n4519) );
  OAI21_X1 U5554 ( .B1(n4510), .B2(n5196), .A(n4519), .ZN(n6578) );
  INV_X1 U5555 ( .A(n5732), .ZN(n5199) );
  AOI222_X1 U5556 ( .A1(n4654), .A2(n4508), .B1(n4544), .B2(n4520), .C1(n6578), 
        .C2(n5199), .ZN(n4535) );
  INV_X1 U5557 ( .A(n6633), .ZN(n6602) );
  OAI21_X1 U5558 ( .B1(n6581), .B2(n4521), .A(n6602), .ZN(n4522) );
  AOI21_X1 U5559 ( .B1(n4522), .B2(n4560), .A(READY_N), .ZN(n4525) );
  OAI21_X1 U5560 ( .B1(n3449), .B2(n4221), .A(n4523), .ZN(n4524) );
  AOI21_X1 U5561 ( .B1(n5209), .B2(n4525), .A(n4524), .ZN(n4526) );
  NAND2_X1 U5562 ( .A1(n4527), .A2(n4526), .ZN(n4532) );
  NAND2_X1 U5563 ( .A1(n5209), .A2(n4537), .ZN(n4531) );
  NAND2_X1 U5564 ( .A1(n4529), .A2(n4528), .ZN(n4530) );
  NAND2_X1 U5565 ( .A1(n4531), .A2(n4530), .ZN(n4649) );
  NAND2_X1 U5566 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4684) );
  NOR2_X1 U5567 ( .A1(n6609), .A2(n4684), .ZN(n6623) );
  AOI22_X1 U5568 ( .A1(n6577), .A2(n6616), .B1(FLUSH_REG_SCAN_IN), .B2(n6623), 
        .ZN(n5842) );
  OAI21_X1 U5569 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n4054), .A(n5842), .ZN(
        n5839) );
  INV_X1 U5570 ( .A(n5839), .ZN(n5201) );
  AOI22_X1 U5571 ( .A1(n5201), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(n4533), .B2(n4654), .ZN(n4534) );
  OAI21_X1 U5572 ( .B1(n4535), .B2(n5201), .A(n4534), .ZN(U3460) );
  INV_X1 U5573 ( .A(n4516), .ZN(n4546) );
  AOI21_X1 U5574 ( .B1(n4546), .B2(n4654), .A(n5201), .ZN(n4550) );
  INV_X1 U5575 ( .A(n4537), .ZN(n4538) );
  NAND2_X1 U5576 ( .A1(n5204), .A2(n4538), .ZN(n4669) );
  XNOR2_X1 U5577 ( .A(n4516), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4542)
         );
  XNOR2_X1 U5578 ( .A(n3223), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4539)
         );
  NAND2_X1 U5579 ( .A1(n6581), .A2(n4539), .ZN(n4540) );
  OAI21_X1 U5580 ( .B1(n4542), .B2(n4341), .A(n4540), .ZN(n4541) );
  AOI21_X1 U5581 ( .B1(n4669), .B2(n4542), .A(n4541), .ZN(n4543) );
  OAI21_X1 U5582 ( .B1(n4536), .B2(n5196), .A(n4543), .ZN(n6576) );
  NOR3_X1 U5583 ( .A1(n6858), .A2(n4545), .A3(n4544), .ZN(n4548) );
  NOR3_X1 U5584 ( .A1(n4546), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n6610), 
        .ZN(n4547) );
  AOI211_X1 U5585 ( .C1(n6576), .C2(n5199), .A(n4548), .B(n4547), .ZN(n4549)
         );
  OAI22_X1 U5586 ( .A1(n4550), .A2(n3223), .B1(n5201), .B2(n4549), .ZN(U3459)
         );
  XNOR2_X1 U5587 ( .A(n4552), .B(n4551), .ZN(n6012) );
  XOR2_X1 U5588 ( .A(n4553), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n4608) );
  NAND2_X1 U5589 ( .A1(n4608), .A2(n4502), .ZN(n4558) );
  NAND2_X1 U5590 ( .A1(n4554), .A2(n5528), .ZN(n4556) );
  NAND2_X1 U5591 ( .A1(n6187), .A2(REIP_REG_0__SCAN_IN), .ZN(n4605) );
  INV_X1 U5592 ( .A(n4605), .ZN(n4555) );
  AOI21_X1 U5593 ( .B1(PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n4556), .A(n4555), 
        .ZN(n4557) );
  OAI211_X1 U5594 ( .C1(n6012), .C2(n5494), .A(n4558), .B(n4557), .ZN(U2986)
         );
  INV_X1 U5595 ( .A(n4559), .ZN(n5735) );
  INV_X1 U5596 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n7016) );
  INV_X2 U5597 ( .A(n6085), .ZN(n6077) );
  INV_X1 U5598 ( .A(DATAI_11_), .ZN(n5072) );
  NOR2_X1 U5599 ( .A1(n6079), .A2(n5072), .ZN(n6080) );
  AOI21_X1 U5600 ( .B1(n6077), .B2(EAX_REG_27__SCAN_IN), .A(n6080), .ZN(n4561)
         );
  OAI21_X1 U5601 ( .B1(n6045), .B2(n7016), .A(n4561), .ZN(U2935) );
  INV_X1 U5602 ( .A(LWORD_REG_9__SCAN_IN), .ZN(n6024) );
  INV_X1 U5603 ( .A(DATAI_9_), .ZN(n4562) );
  NOR2_X1 U5604 ( .A1(n6079), .A2(n4562), .ZN(n6056) );
  AOI21_X1 U5605 ( .B1(n6077), .B2(EAX_REG_9__SCAN_IN), .A(n6056), .ZN(n4563)
         );
  OAI21_X1 U5606 ( .B1(n6045), .B2(n6024), .A(n4563), .ZN(U2948) );
  INV_X1 U5607 ( .A(LWORD_REG_12__SCAN_IN), .ZN(n6873) );
  INV_X1 U5608 ( .A(DATAI_12_), .ZN(n5180) );
  NOR2_X1 U5609 ( .A1(n6079), .A2(n5180), .ZN(n4567) );
  AOI21_X1 U5610 ( .B1(n6077), .B2(EAX_REG_12__SCAN_IN), .A(n4567), .ZN(n4564)
         );
  OAI21_X1 U5611 ( .B1(n6045), .B2(n6873), .A(n4564), .ZN(U2951) );
  INV_X1 U5612 ( .A(LWORD_REG_13__SCAN_IN), .ZN(n6816) );
  INV_X1 U5613 ( .A(DATAI_13_), .ZN(n4565) );
  NOR2_X1 U5614 ( .A1(n6079), .A2(n4565), .ZN(n6058) );
  AOI21_X1 U5615 ( .B1(n6077), .B2(EAX_REG_13__SCAN_IN), .A(n6058), .ZN(n4566)
         );
  OAI21_X1 U5616 ( .B1(n6045), .B2(n6816), .A(n4566), .ZN(U2952) );
  INV_X1 U5617 ( .A(UWORD_REG_12__SCAN_IN), .ZN(n7020) );
  AOI21_X1 U5618 ( .B1(n6077), .B2(EAX_REG_28__SCAN_IN), .A(n4567), .ZN(n4568)
         );
  OAI21_X1 U5619 ( .B1(n6045), .B2(n7020), .A(n4568), .ZN(U2936) );
  INV_X1 U5620 ( .A(UWORD_REG_10__SCAN_IN), .ZN(n6917) );
  NAND2_X1 U5621 ( .A1(n6077), .A2(EAX_REG_26__SCAN_IN), .ZN(n4570) );
  INV_X1 U5622 ( .A(n6079), .ZN(n4569) );
  NAND2_X1 U5623 ( .A1(n4569), .A2(DATAI_10_), .ZN(n4571) );
  OAI211_X1 U5624 ( .C1(n6045), .C2(n6917), .A(n4570), .B(n4571), .ZN(U2934)
         );
  INV_X1 U5625 ( .A(LWORD_REG_10__SCAN_IN), .ZN(n6840) );
  NAND2_X1 U5626 ( .A1(n6077), .A2(EAX_REG_10__SCAN_IN), .ZN(n4572) );
  OAI211_X1 U5627 ( .C1(n6045), .C2(n6840), .A(n4572), .B(n4571), .ZN(U2949)
         );
  NOR2_X1 U5628 ( .A1(n4574), .A2(n4575), .ZN(n4576) );
  OR2_X1 U5629 ( .A1(n3570), .A2(n4576), .ZN(n4653) );
  INV_X1 U5630 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4578) );
  XNOR2_X1 U5631 ( .A(n4577), .B(n3190), .ZN(n5957) );
  OAI222_X1 U5632 ( .A1(n4653), .A2(n5389), .B1(n4578), .B2(n5989), .C1(n5957), 
        .C2(n5984), .ZN(U2858) );
  INV_X1 U5633 ( .A(DATAI_15_), .ZN(n5415) );
  INV_X1 U5634 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4579) );
  INV_X1 U5635 ( .A(EAX_REG_15__SCAN_IN), .ZN(n5416) );
  OAI222_X1 U5636 ( .A1(n5415), .A2(n6079), .B1(n4579), .B2(n6045), .C1(n5416), 
        .C2(n6085), .ZN(U2954) );
  XNOR2_X1 U5637 ( .A(n4580), .B(n4581), .ZN(n4626) );
  INV_X1 U5638 ( .A(n4732), .ZN(n4585) );
  AND3_X1 U5639 ( .A1(n4733), .A2(n6848), .A3(n4582), .ZN(n4584) );
  OAI22_X1 U5640 ( .A1(n6119), .A2(n5957), .B1(n6647), .B2(n6177), .ZN(n4583)
         );
  AOI211_X1 U5641 ( .C1(n4585), .C2(INSTADDRPOINTER_REG_1__SCAN_IN), .A(n4584), 
        .B(n4583), .ZN(n4586) );
  OAI21_X1 U5642 ( .B1(n4626), .B2(n5721), .A(n4586), .ZN(U3017) );
  INV_X1 U5643 ( .A(n6581), .ZN(n4587) );
  INV_X2 U5644 ( .A(n6708), .ZN(n6041) );
  INV_X1 U5645 ( .A(n4644), .ZN(n6015) );
  AOI222_X1 U5646 ( .A1(n6040), .A2(DATAO_REG_27__SCAN_IN), .B1(n6015), .B2(
        EAX_REG_27__SCAN_IN), .C1(n6041), .C2(UWORD_REG_11__SCAN_IN), .ZN(
        n4592) );
  INV_X1 U5647 ( .A(n4592), .ZN(U2896) );
  OAI21_X1 U5648 ( .B1(n4594), .B2(n4593), .A(n4690), .ZN(n6186) );
  INV_X1 U5649 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4599) );
  INV_X1 U5650 ( .A(n4595), .ZN(n4598) );
  CLKBUF_X1 U5651 ( .A(n4597), .Z(n4613) );
  AOI21_X1 U5652 ( .B1(n4598), .B2(n4596), .A(n4613), .ZN(n6112) );
  INV_X1 U5653 ( .A(n6112), .ZN(n5103) );
  OAI222_X1 U5654 ( .A1(n6186), .A2(n5984), .B1(n4599), .B2(n5989), .C1(n5103), 
        .C2(n5389), .ZN(U2857) );
  INV_X1 U5655 ( .A(n4600), .ZN(n4603) );
  NAND2_X1 U5656 ( .A1(n4601), .A2(n4545), .ZN(n4602) );
  NAND2_X1 U5657 ( .A1(n4603), .A2(n4602), .ZN(n4910) );
  OAI21_X1 U5658 ( .B1(n5829), .B2(n4604), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4606) );
  OAI211_X1 U5659 ( .C1(n6119), .C2(n4910), .A(n4606), .B(n4605), .ZN(n4607)
         );
  AOI21_X1 U5660 ( .B1(n4608), .B2(n4243), .A(n4607), .ZN(n4609) );
  NAND2_X1 U5661 ( .A1(n4610), .A2(n4609), .ZN(U3018) );
  CLKBUF_X1 U5662 ( .A(n4612), .Z(n4708) );
  OAI21_X1 U5663 ( .B1(n4613), .B2(n4611), .A(n4708), .ZN(n4995) );
  INV_X1 U5664 ( .A(n4614), .ZN(n4983) );
  INV_X1 U5665 ( .A(REIP_REG_3__SCAN_IN), .ZN(n4615) );
  OAI22_X1 U5666 ( .A1(n5528), .A2(n4616), .B1(n6177), .B2(n4615), .ZN(n4617)
         );
  AOI21_X1 U5667 ( .B1(n6088), .B2(n4983), .A(n4617), .ZN(n4622) );
  OR2_X1 U5668 ( .A1(n4619), .A2(n4618), .ZN(n6176) );
  NAND3_X1 U5669 ( .A1(n6176), .A2(n4502), .A3(n4620), .ZN(n4621) );
  OAI211_X1 U5670 ( .C1(n4995), .C2(n5494), .A(n4622), .B(n4621), .ZN(U2983)
         );
  INV_X1 U5671 ( .A(n4653), .ZN(n5970) );
  AOI22_X1 U5672 ( .A1(n6108), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6187), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4623) );
  OAI21_X1 U5673 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6117), .A(n4623), 
        .ZN(n4624) );
  AOI21_X1 U5674 ( .B1(n5970), .B2(n6113), .A(n4624), .ZN(n4625) );
  OAI21_X1 U5675 ( .B1(n4626), .B2(n6092), .A(n4625), .ZN(U2985) );
  INV_X1 U5676 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4628) );
  AOI22_X1 U5677 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n6041), .B1(n6040), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4627) );
  OAI21_X1 U5678 ( .B1(n4628), .B2(n4644), .A(n4627), .ZN(U2902) );
  INV_X1 U5679 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4630) );
  AOI22_X1 U5680 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n6041), .B1(n6040), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4629) );
  OAI21_X1 U5681 ( .B1(n4630), .B2(n4644), .A(n4629), .ZN(U2905) );
  INV_X1 U5682 ( .A(EAX_REG_28__SCAN_IN), .ZN(n7027) );
  AOI22_X1 U5683 ( .A1(UWORD_REG_12__SCAN_IN), .A2(n6041), .B1(n6040), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4631) );
  OAI21_X1 U5684 ( .B1(n7027), .B2(n4644), .A(n4631), .ZN(U2895) );
  INV_X1 U5685 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4633) );
  AOI22_X1 U5686 ( .A1(n6041), .A2(UWORD_REG_1__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4632) );
  OAI21_X1 U5687 ( .B1(n4633), .B2(n4644), .A(n4632), .ZN(U2906) );
  INV_X1 U5688 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6063) );
  AOI22_X1 U5689 ( .A1(n6041), .A2(UWORD_REG_14__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4634) );
  OAI21_X1 U5690 ( .B1(n6063), .B2(n4644), .A(n4634), .ZN(U2893) );
  INV_X1 U5691 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4636) );
  AOI22_X1 U5692 ( .A1(n6041), .A2(UWORD_REG_4__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4635) );
  OAI21_X1 U5693 ( .B1(n4636), .B2(n4644), .A(n4635), .ZN(U2903) );
  INV_X1 U5694 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4638) );
  AOI22_X1 U5695 ( .A1(n6041), .A2(UWORD_REG_7__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4637) );
  OAI21_X1 U5696 ( .B1(n4638), .B2(n4644), .A(n4637), .ZN(U2900) );
  INV_X1 U5697 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4640) );
  AOI22_X1 U5698 ( .A1(n6041), .A2(UWORD_REG_3__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4639) );
  OAI21_X1 U5699 ( .B1(n4640), .B2(n4644), .A(n4639), .ZN(U2904) );
  AOI22_X1 U5700 ( .A1(n6041), .A2(UWORD_REG_9__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4641) );
  OAI21_X1 U5701 ( .B1(n4001), .B2(n4644), .A(n4641), .ZN(U2898) );
  INV_X1 U5702 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6060) );
  AOI22_X1 U5703 ( .A1(n6041), .A2(UWORD_REG_13__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4642) );
  OAI21_X1 U5704 ( .B1(n6060), .B2(n4644), .A(n4642), .ZN(U2894) );
  INV_X1 U5705 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4645) );
  AOI22_X1 U5706 ( .A1(n6041), .A2(UWORD_REG_8__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4643) );
  OAI21_X1 U5707 ( .B1(n4645), .B2(n4644), .A(n4643), .ZN(U2899) );
  OR2_X1 U5708 ( .A1(n3431), .A2(n3433), .ZN(n4646) );
  NOR2_X1 U5709 ( .A1(n4647), .A2(n4646), .ZN(n4648) );
  NAND2_X1 U5710 ( .A1(n3460), .A2(n3428), .ZN(n4651) );
  INV_X1 U5711 ( .A(n4651), .ZN(n4652) );
  INV_X1 U5712 ( .A(DATAI_2_), .ZN(n6068) );
  INV_X1 U5713 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6037) );
  OAI222_X1 U5714 ( .A1(n5103), .A2(n6011), .B1(n6009), .B2(n6068), .C1(n6010), 
        .C2(n6037), .ZN(U2889) );
  INV_X1 U5715 ( .A(DATAI_1_), .ZN(n6961) );
  INV_X1 U5716 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6039) );
  OAI222_X1 U5717 ( .A1(n4653), .A2(n6011), .B1(n6009), .B2(n6961), .C1(n6010), 
        .C2(n6039), .ZN(U2890) );
  NAND2_X1 U5718 ( .A1(n6441), .A2(n4656), .ZN(n4671) );
  MUX2_X1 U5719 ( .A(n4657), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4516), 
        .Z(n4658) );
  NOR2_X1 U5720 ( .A1(n4658), .A2(n4673), .ZN(n4668) );
  INV_X1 U5721 ( .A(n4659), .ZN(n4660) );
  OAI21_X1 U5722 ( .B1(n4516), .B2(n3284), .A(n4660), .ZN(n4661) );
  NOR2_X1 U5723 ( .A1(n4661), .A2(n3526), .ZN(n5731) );
  AND2_X1 U5724 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4664) );
  INV_X1 U5725 ( .A(n4664), .ZN(n4663) );
  MUX2_X1 U5726 ( .A(n4664), .B(n4663), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4665) );
  NAND2_X1 U5727 ( .A1(n6581), .A2(n4665), .ZN(n4666) );
  OAI21_X1 U5728 ( .B1(n5731), .B2(n4341), .A(n4666), .ZN(n4667) );
  AOI21_X1 U5729 ( .B1(n4669), .B2(n4668), .A(n4667), .ZN(n4670) );
  NAND2_X1 U5730 ( .A1(n4671), .A2(n4670), .ZN(n6574) );
  NAND4_X1 U5731 ( .A1(n6574), .A2(n6858), .A3(n6576), .A4(n6577), .ZN(n4679)
         );
  INV_X1 U5732 ( .A(FLUSH_REG_SCAN_IN), .ZN(n7032) );
  NAND2_X1 U5733 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n7032), .ZN(n4672) );
  OAI21_X1 U5734 ( .B1(n6577), .B2(STATE2_REG_1__SCAN_IN), .A(n4672), .ZN(
        n4674) );
  NAND2_X1 U5735 ( .A1(n4674), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4680) );
  NAND2_X1 U5736 ( .A1(n4674), .A2(n4673), .ZN(n4675) );
  AND2_X1 U5737 ( .A1(n4680), .A2(n4675), .ZN(n4678) );
  INV_X1 U5738 ( .A(n5031), .ZN(n6295) );
  NOR2_X1 U5739 ( .A1(n3188), .A2(n6295), .ZN(n4676) );
  XNOR2_X1 U5740 ( .A(n4676), .B(n5840), .ZN(n5948) );
  NOR2_X1 U5741 ( .A1(n4238), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4677) );
  NAND2_X1 U5742 ( .A1(n5948), .A2(n4677), .ZN(n5837) );
  INV_X1 U5743 ( .A(n6597), .ZN(n4682) );
  NAND2_X1 U5744 ( .A1(n4680), .A2(n4517), .ZN(n4681) );
  OAI21_X1 U5745 ( .B1(n4685), .B2(FLUSH_REG_SCAN_IN), .A(n6623), .ZN(n4683)
         );
  NAND2_X1 U5746 ( .A1(n4881), .A2(n4683), .ZN(n6201) );
  NOR2_X1 U5747 ( .A1(n4685), .A2(n4684), .ZN(n6608) );
  INV_X1 U5748 ( .A(n4686), .ZN(n5197) );
  NAND2_X1 U5749 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n4054), .ZN(n4697) );
  INV_X1 U5750 ( .A(n4697), .ZN(n5728) );
  OAI22_X1 U5751 ( .A1(n5104), .A2(n6519), .B1(n5197), .B2(n5728), .ZN(n4687)
         );
  OAI21_X1 U5752 ( .B1(n6608), .B2(n4687), .A(n6201), .ZN(n4688) );
  OAI21_X1 U5753 ( .B1(n6201), .B2(n6580), .A(n4688), .ZN(U3465) );
  NAND2_X1 U5754 ( .A1(n4690), .A2(n4689), .ZN(n4691) );
  AND2_X1 U5755 ( .A1(n4709), .A2(n4691), .ZN(n6179) );
  INV_X1 U5756 ( .A(n5989), .ZN(n5387) );
  AOI22_X1 U5757 ( .A1(n5980), .A2(n6179), .B1(EBX_REG_3__SCAN_IN), .B2(n5387), 
        .ZN(n4692) );
  OAI21_X1 U5758 ( .B1(n4995), .B2(n5389), .A(n4692), .ZN(U2856) );
  OAI222_X1 U5759 ( .A1(n5984), .A2(n4910), .B1(n4911), .B2(n5989), .C1(n5389), 
        .C2(n6012), .ZN(U2859) );
  INV_X1 U5760 ( .A(n6201), .ZN(n4702) );
  INV_X1 U5761 ( .A(n4693), .ZN(n4695) );
  NAND2_X1 U5762 ( .A1(n5723), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5726) );
  NOR2_X1 U5763 ( .A1(n5723), .A2(n4695), .ZN(n4696) );
  NAND2_X1 U5764 ( .A1(n3187), .A2(n4696), .ZN(n6507) );
  OAI211_X1 U5765 ( .C1(n6338), .C2(n5726), .A(n6471), .B(n6507), .ZN(n4699)
         );
  INV_X1 U5766 ( .A(n4694), .ZN(n4698) );
  OR2_X1 U5767 ( .A1(n6519), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6508) );
  INV_X1 U5768 ( .A(n6508), .ZN(n6439) );
  AOI222_X1 U5769 ( .A1(n4699), .A2(n6506), .B1(n4698), .B2(n6439), .C1(n6441), 
        .C2(n4697), .ZN(n4701) );
  NAND2_X1 U5770 ( .A1(n4702), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4700) );
  OAI21_X1 U5771 ( .B1(n4702), .B2(n4701), .A(n4700), .ZN(U3462) );
  INV_X1 U5772 ( .A(n4706), .ZN(n4707) );
  AOI21_X1 U5773 ( .B1(n4704), .B2(n4708), .A(n4707), .ZN(n6104) );
  INV_X1 U5774 ( .A(n6104), .ZN(n4724) );
  AOI21_X1 U5775 ( .B1(n4710), .B2(n4709), .A(n4714), .ZN(n6168) );
  AOI22_X1 U5776 ( .A1(n6168), .A2(n5980), .B1(EBX_REG_4__SCAN_IN), .B2(n5387), 
        .ZN(n4711) );
  OAI21_X1 U5777 ( .B1(n4724), .B2(n5389), .A(n4711), .ZN(U2855) );
  XOR2_X1 U5778 ( .A(n4712), .B(n4706), .Z(n5941) );
  INV_X1 U5779 ( .A(n5941), .ZN(n4743) );
  OR2_X1 U5780 ( .A1(n4714), .A2(n4713), .ZN(n4715) );
  AND2_X1 U5781 ( .A1(n4715), .A2(n4752), .ZN(n5933) );
  AOI22_X1 U5782 ( .A1(n5980), .A2(n5933), .B1(EBX_REG_5__SCAN_IN), .B2(n5387), 
        .ZN(n4716) );
  OAI21_X1 U5783 ( .B1(n4743), .B2(n5389), .A(n4716), .ZN(U2854) );
  OAI21_X1 U5784 ( .B1(n4719), .B2(n4718), .A(n4717), .ZN(n4741) );
  INV_X1 U5785 ( .A(REIP_REG_5__SCAN_IN), .ZN(n4720) );
  NOR2_X1 U5786 ( .A1(n6177), .A2(n4720), .ZN(n4738) );
  AOI21_X1 U5787 ( .B1(n6108), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n4738), 
        .ZN(n4721) );
  OAI21_X1 U5788 ( .B1(n5938), .B2(n6117), .A(n4721), .ZN(n4722) );
  AOI21_X1 U5789 ( .B1(n5941), .B2(n6113), .A(n4722), .ZN(n4723) );
  OAI21_X1 U5790 ( .B1(n4741), .B2(n6092), .A(n4723), .ZN(U2981) );
  INV_X1 U5791 ( .A(DATAI_4_), .ZN(n6072) );
  INV_X1 U5792 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6033) );
  OAI222_X1 U5793 ( .A1(n4724), .A2(n6011), .B1(n6009), .B2(n6072), .C1(n6033), 
        .C2(n6010), .ZN(U2887) );
  OR2_X1 U5794 ( .A1(n4727), .A2(n4726), .ZN(n4728) );
  AND2_X1 U5795 ( .A1(n4746), .A2(n4728), .ZN(n6096) );
  INV_X1 U5796 ( .A(n6096), .ZN(n4755) );
  AOI22_X1 U5797 ( .A1(n6005), .A2(DATAI_6_), .B1(EAX_REG_6__SCAN_IN), .B2(
        n5999), .ZN(n4729) );
  OAI21_X1 U5798 ( .B1(n4755), .B2(n6011), .A(n4729), .ZN(U2885) );
  INV_X1 U5799 ( .A(DATAI_3_), .ZN(n6070) );
  INV_X1 U5800 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6035) );
  OAI222_X1 U5801 ( .A1(n4995), .A2(n6011), .B1(n6009), .B2(n6070), .C1(n6010), 
        .C2(n6035), .ZN(U2888) );
  NAND2_X1 U5802 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4730), .ZN(n5087)
         );
  INV_X1 U5803 ( .A(n5653), .ZN(n4731) );
  OAI22_X1 U5804 ( .A1(n4732), .A2(n6190), .B1(n4731), .B2(n5086), .ZN(n6194)
         );
  AOI21_X1 U5805 ( .B1(n4733), .B2(n5087), .A(n6194), .ZN(n6167) );
  AOI21_X1 U5806 ( .B1(n7026), .B2(n4734), .A(n6167), .ZN(n4739) );
  NAND2_X1 U5807 ( .A1(n5086), .A2(n6196), .ZN(n4735) );
  NOR3_X1 U5808 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6170), .A3(n4735), 
        .ZN(n4737) );
  AND2_X1 U5809 ( .A1(n5933), .A2(n6189), .ZN(n4736) );
  NOR4_X1 U5810 ( .A1(n4739), .A2(n4738), .A3(n4737), .A4(n4736), .ZN(n4740)
         );
  OAI21_X1 U5811 ( .B1(n5721), .B2(n4741), .A(n4740), .ZN(U3013) );
  INV_X1 U5812 ( .A(DATAI_5_), .ZN(n4744) );
  OAI222_X1 U5813 ( .A1(n4744), .A2(n6009), .B1(n6011), .B2(n4743), .C1(n4742), 
        .C2(n6010), .ZN(U2886) );
  XOR2_X1 U5814 ( .A(n4745), .B(n4746), .Z(n4825) );
  AND2_X1 U5815 ( .A1(n4754), .A2(n4747), .ZN(n4748) );
  NOR2_X1 U5816 ( .A1(n4828), .A2(n4748), .ZN(n6156) );
  NOR2_X1 U5817 ( .A1(n5989), .A2(n6871), .ZN(n4749) );
  AOI21_X1 U5818 ( .B1(n6156), .B2(n5980), .A(n4749), .ZN(n4750) );
  OAI21_X1 U5819 ( .B1(n5345), .B2(n5389), .A(n4750), .ZN(U2852) );
  NAND2_X1 U5820 ( .A1(n4752), .A2(n4751), .ZN(n4753) );
  NAND2_X1 U5821 ( .A1(n4754), .A2(n4753), .ZN(n6161) );
  INV_X1 U5822 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4756) );
  OAI222_X1 U5823 ( .A1(n6161), .A2(n5984), .B1(n4756), .B2(n5989), .C1(n4755), 
        .C2(n5389), .ZN(U2853) );
  INV_X1 U5824 ( .A(DATAI_7_), .ZN(n4758) );
  OAI222_X1 U5825 ( .A1(n6009), .A2(n4758), .B1(n6011), .B2(n5345), .C1(n4757), 
        .C2(n6010), .ZN(U2884) );
  INV_X1 U5826 ( .A(n4886), .ZN(n4879) );
  NOR2_X1 U5827 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4879), .ZN(n4976)
         );
  NOR2_X1 U5828 ( .A1(n4767), .A2(n6505), .ZN(n4787) );
  OAI21_X1 U5829 ( .B1(n6288), .B2(n6505), .A(n4940), .ZN(n5110) );
  NOR2_X1 U5830 ( .A1(n4787), .A2(n5110), .ZN(n6299) );
  NOR2_X1 U5831 ( .A1(n6505), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6446)
         );
  INV_X1 U5832 ( .A(n6446), .ZN(n4759) );
  OAI211_X1 U5833 ( .C1(n4054), .C2(n4976), .A(n6299), .B(n4759), .ZN(n4765)
         );
  OR2_X1 U5834 ( .A1(n6507), .A2(n5104), .ZN(n4815) );
  AND2_X1 U5835 ( .A1(n5723), .A2(n4693), .ZN(n4760) );
  INV_X1 U5836 ( .A(n4882), .ZN(n4761) );
  AOI21_X1 U5837 ( .B1(n4815), .B2(n5006), .A(n6832), .ZN(n4763) );
  NOR2_X1 U5838 ( .A1(n4536), .A2(n4510), .ZN(n6296) );
  NAND2_X1 U5839 ( .A1(n6296), .A2(n6441), .ZN(n4769) );
  INV_X1 U5840 ( .A(n4769), .ZN(n4762) );
  NOR3_X1 U5841 ( .A1(n4763), .A2(n4762), .A3(n6519), .ZN(n4764) );
  INV_X1 U5842 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4774) );
  INV_X1 U5843 ( .A(DATAI_31_), .ZN(n4766) );
  NOR2_X2 U5844 ( .A1(n5494), .A2(n4766), .ZN(n6564) );
  NAND2_X1 U5845 ( .A1(n6113), .A2(DATAI_23_), .ZN(n6328) );
  NAND2_X1 U5846 ( .A1(DATAI_7_), .A2(n4940), .ZN(n6572) );
  NAND2_X1 U5847 ( .A1(n4767), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6370) );
  INV_X1 U5848 ( .A(n6370), .ZN(n6289) );
  NAND3_X1 U5849 ( .A1(n6289), .A2(n6288), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4768) );
  OAI21_X1 U5850 ( .B1(n4769), .B2(n6519), .A(n4768), .ZN(n4977) );
  NOR2_X2 U5851 ( .A1(n4942), .A2(n5189), .ZN(n6566) );
  AOI22_X1 U5852 ( .A1(n6401), .A2(n4977), .B1(n6566), .B2(n4976), .ZN(n4771)
         );
  OAI21_X1 U5853 ( .B1(n6328), .B2(n5006), .A(n4771), .ZN(n4772) );
  AOI21_X1 U5854 ( .B1(n6564), .B2(n6567), .A(n4772), .ZN(n4773) );
  OAI21_X1 U5855 ( .B1(n4982), .B2(n4774), .A(n4773), .ZN(U3139) );
  INV_X1 U5856 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4779) );
  NAND2_X1 U5857 ( .A1(n6113), .A2(DATAI_27_), .ZN(n6386) );
  INV_X1 U5858 ( .A(DATAI_19_), .ZN(n4775) );
  NOR2_X1 U5859 ( .A1(n5494), .A2(n4775), .ZN(n6541) );
  INV_X1 U5860 ( .A(n6541), .ZN(n6311) );
  NAND2_X1 U5861 ( .A1(DATAI_3_), .A2(n4940), .ZN(n6544) );
  NOR2_X2 U5862 ( .A1(n4942), .A2(n3454), .ZN(n6540) );
  AOI22_X1 U5863 ( .A1(n6383), .A2(n4977), .B1(n6540), .B2(n4976), .ZN(n4776)
         );
  OAI21_X1 U5864 ( .B1(n6311), .B2(n5006), .A(n4776), .ZN(n4777) );
  AOI21_X1 U5865 ( .B1(n6539), .B2(n6567), .A(n4777), .ZN(n4778) );
  OAI21_X1 U5866 ( .B1(n4982), .B2(n4779), .A(n4778), .ZN(U3135) );
  INV_X1 U5867 ( .A(n6410), .ZN(n4780) );
  AOI21_X1 U5868 ( .B1(n6231), .B2(n4780), .A(n6519), .ZN(n6207) );
  NAND3_X1 U5869 ( .A1(n3187), .A2(n6230), .A3(n4693), .ZN(n4946) );
  NAND2_X1 U5870 ( .A1(n4536), .A2(n4510), .ZN(n6407) );
  NOR2_X1 U5871 ( .A1(n6441), .A2(n6407), .ZN(n6203) );
  AOI21_X1 U5872 ( .B1(n5002), .B2(n6508), .A(n6203), .ZN(n4786) );
  NAND3_X1 U5873 ( .A1(n6589), .A2(n6363), .A3(n6925), .ZN(n6204) );
  NOR2_X1 U5874 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6204), .ZN(n4943)
         );
  INV_X1 U5875 ( .A(n4943), .ZN(n4873) );
  INV_X1 U5876 ( .A(n4802), .ZN(n4782) );
  OR2_X1 U5877 ( .A1(n6288), .A2(n4782), .ZN(n6258) );
  INV_X1 U5878 ( .A(n6258), .ZN(n4783) );
  OAI21_X1 U5879 ( .B1(n4783), .B2(n6505), .A(n4940), .ZN(n6260) );
  AOI211_X1 U5880 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4873), .A(n6289), .B(
        n6260), .ZN(n4784) );
  INV_X1 U5881 ( .A(n4784), .ZN(n4785) );
  INV_X1 U5882 ( .A(n6328), .ZN(n6568) );
  INV_X1 U5883 ( .A(n6564), .ZN(n6406) );
  INV_X1 U5884 ( .A(n6441), .ZN(n6367) );
  NAND2_X1 U5885 ( .A1(n6367), .A2(n6506), .ZN(n6292) );
  INV_X1 U5886 ( .A(n4787), .ZN(n6361) );
  OAI22_X1 U5887 ( .A1(n6292), .A2(n6407), .B1(n6361), .B2(n6258), .ZN(n4944)
         );
  AOI22_X1 U5888 ( .A1(n6401), .A2(n4944), .B1(n6566), .B2(n4943), .ZN(n4788)
         );
  OAI21_X1 U5889 ( .B1(n6406), .B2(n4946), .A(n4788), .ZN(n4789) );
  AOI21_X1 U5890 ( .B1(n6568), .B2(n6225), .A(n4789), .ZN(n4790) );
  OAI21_X1 U5891 ( .B1(n4950), .B2(n4791), .A(n4790), .ZN(U3027) );
  INV_X1 U5892 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n6822) );
  AOI22_X1 U5893 ( .A1(n6383), .A2(n4944), .B1(n6540), .B2(n4943), .ZN(n4792)
         );
  OAI21_X1 U5894 ( .B1(n6386), .B2(n4946), .A(n4792), .ZN(n4793) );
  AOI21_X1 U5895 ( .B1(n6541), .B2(n6225), .A(n4793), .ZN(n4794) );
  OAI21_X1 U5896 ( .B1(n4950), .B2(n6822), .A(n4794), .ZN(U3023) );
  AOI21_X1 U5897 ( .B1(n4797), .B2(n4795), .A(n4796), .ZN(n4846) );
  INV_X1 U5898 ( .A(n4846), .ZN(n5332) );
  AOI22_X1 U5899 ( .A1(n6005), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n5999), .ZN(n4798) );
  OAI21_X1 U5900 ( .B1(n5332), .B2(n6011), .A(n4798), .ZN(U2883) );
  NOR2_X2 U5901 ( .A1(n6471), .A2(n6337), .ZN(n6499) );
  INV_X1 U5902 ( .A(n6499), .ZN(n4800) );
  INV_X1 U5903 ( .A(n6507), .ZN(n4799) );
  NAND3_X1 U5904 ( .A1(n4800), .A2(n6506), .A3(n5018), .ZN(n4801) );
  INV_X1 U5905 ( .A(n4536), .ZN(n5098) );
  NAND2_X1 U5906 ( .A1(n5098), .A2(n4510), .ZN(n6511) );
  INV_X1 U5907 ( .A(n6511), .ZN(n4805) );
  AOI22_X1 U5908 ( .A1(n4801), .A2(n6508), .B1(n4805), .B2(n5031), .ZN(n4804)
         );
  NAND2_X1 U5909 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6514), .ZN(n6518) );
  NOR2_X1 U5910 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6518), .ZN(n5015)
         );
  OR2_X1 U5911 ( .A1(n6288), .A2(n4802), .ZN(n6362) );
  AOI21_X1 U5912 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6362), .A(n4881), .ZN(
        n6371) );
  OAI211_X1 U5913 ( .C1(n4054), .C2(n5015), .A(n6371), .B(n6361), .ZN(n4803)
         );
  INV_X1 U5914 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4810) );
  NAND3_X1 U5915 ( .A1(n4805), .A2(n6506), .A3(n6441), .ZN(n4806) );
  OAI21_X1 U5916 ( .B1(n6370), .B2(n6362), .A(n4806), .ZN(n5016) );
  AOI22_X1 U5917 ( .A1(n6383), .A2(n5016), .B1(n5015), .B2(n6540), .ZN(n4807)
         );
  OAI21_X1 U5918 ( .B1(n6311), .B2(n5018), .A(n4807), .ZN(n4808) );
  AOI21_X1 U5919 ( .B1(n6539), .B2(n6499), .A(n4808), .ZN(n4809) );
  OAI21_X1 U5920 ( .B1(n5022), .B2(n4810), .A(n4809), .ZN(U3119) );
  INV_X1 U5921 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4814) );
  AOI22_X1 U5922 ( .A1(n6401), .A2(n5016), .B1(n5015), .B2(n6566), .ZN(n4811)
         );
  OAI21_X1 U5923 ( .B1(n6328), .B2(n5018), .A(n4811), .ZN(n4812) );
  AOI21_X1 U5924 ( .B1(n6564), .B2(n6499), .A(n4812), .ZN(n4813) );
  OAI21_X1 U5925 ( .B1(n5022), .B2(n4814), .A(n4813), .ZN(U3123) );
  INV_X1 U5926 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4819) );
  INV_X1 U5927 ( .A(DATAI_0_), .ZN(n6065) );
  NOR2_X2 U5928 ( .A1(n4942), .A2(n4854), .ZN(n6516) );
  AOI22_X1 U5929 ( .A1(n6364), .A2(n4977), .B1(n6516), .B2(n4976), .ZN(n4818)
         );
  INV_X1 U5930 ( .A(DATAI_24_), .ZN(n6828) );
  NOR2_X1 U5931 ( .A1(n5494), .A2(n6828), .ZN(n6524) );
  INV_X1 U5932 ( .A(n6524), .ZN(n6727) );
  INV_X1 U5933 ( .A(DATAI_16_), .ZN(n6923) );
  NOR2_X1 U5934 ( .A1(n5494), .A2(n6923), .ZN(n6515) );
  INV_X1 U5935 ( .A(n6515), .ZN(n6726) );
  OAI22_X1 U5936 ( .A1(n6727), .A2(n4815), .B1(n5006), .B2(n6726), .ZN(n4816)
         );
  INV_X1 U5937 ( .A(n4816), .ZN(n4817) );
  OAI211_X1 U5938 ( .C1(n4982), .C2(n4819), .A(n4818), .B(n4817), .ZN(U3132)
         );
  OAI21_X1 U5939 ( .B1(n4822), .B2(n4821), .A(n4820), .ZN(n6154) );
  AOI22_X1 U5940 ( .A1(n6108), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .B1(n6187), 
        .B2(REIP_REG_7__SCAN_IN), .ZN(n4823) );
  OAI21_X1 U5941 ( .B1(n5335), .B2(n6117), .A(n4823), .ZN(n4824) );
  AOI21_X1 U5942 ( .B1(n4825), .B2(n6113), .A(n4824), .ZN(n4826) );
  OAI21_X1 U5943 ( .B1(n6154), .B2(n6092), .A(n4826), .ZN(U2979) );
  INV_X1 U5944 ( .A(n4838), .ZN(n4827) );
  OAI21_X1 U5945 ( .B1(n4829), .B2(n4828), .A(n4827), .ZN(n6143) );
  INV_X1 U5946 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4830) );
  OAI222_X1 U5947 ( .A1(n6143), .A2(n5984), .B1(n5989), .B2(n4830), .C1(n5332), 
        .C2(n5389), .ZN(U2851) );
  INV_X1 U5948 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4833) );
  AOI22_X1 U5949 ( .A1(n6364), .A2(n5016), .B1(n5015), .B2(n6516), .ZN(n4832)
         );
  AOI22_X1 U5950 ( .A1(n6499), .A2(n6524), .B1(n6515), .B2(n6563), .ZN(n4831)
         );
  OAI211_X1 U5951 ( .C1(n5022), .C2(n4833), .A(n4832), .B(n4831), .ZN(U3116)
         );
  OR2_X1 U5952 ( .A1(n4796), .A2(n4835), .ZN(n4836) );
  AND2_X1 U5953 ( .A1(n4834), .A2(n4836), .ZN(n6007) );
  INV_X1 U5954 ( .A(n6007), .ZN(n4840) );
  INV_X1 U5955 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4839) );
  OAI21_X1 U5956 ( .B1(n4838), .B2(n4837), .A(n4852), .ZN(n5915) );
  OAI222_X1 U5957 ( .A1(n4840), .A2(n5389), .B1(n4839), .B2(n5989), .C1(n5984), 
        .C2(n5915), .ZN(U2850) );
  OAI21_X1 U5958 ( .B1(n4843), .B2(n4842), .A(n4841), .ZN(n6147) );
  NAND2_X1 U5959 ( .A1(n6187), .A2(REIP_REG_8__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U5960 ( .A1(n6108), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4844)
         );
  OAI211_X1 U5961 ( .C1(n6117), .C2(n5325), .A(n6144), .B(n4844), .ZN(n4845)
         );
  AOI21_X1 U5962 ( .B1(n4846), .B2(n6113), .A(n4845), .ZN(n4847) );
  OAI21_X1 U5963 ( .B1(n6147), .B2(n6092), .A(n4847), .ZN(U2978) );
  INV_X1 U5964 ( .A(n4834), .ZN(n4850) );
  OAI21_X1 U5965 ( .B1(n4850), .B2(n3733), .A(n4849), .ZN(n5147) );
  INV_X1 U5966 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4861) );
  INV_X1 U5967 ( .A(n5027), .ZN(n4851) );
  AOI21_X1 U5968 ( .B1(n4853), .B2(n4852), .A(n4851), .ZN(n6135) );
  NOR2_X1 U5969 ( .A1(n4854), .A2(EBX_REG_31__SCAN_IN), .ZN(n4855) );
  NAND2_X1 U5970 ( .A1(n4856), .A2(n4855), .ZN(n4858) );
  NAND2_X2 U5971 ( .A1(n4858), .A2(n4857), .ZN(n5968) );
  AOI22_X1 U5972 ( .A1(n6135), .A2(n5904), .B1(EBX_REG_10__SCAN_IN), .B2(n5968), .ZN(n4860) );
  NAND2_X1 U5973 ( .A1(n5773), .A2(n4859), .ZN(n5924) );
  OAI211_X1 U5974 ( .C1(n5934), .C2(n4861), .A(n4860), .B(n5924), .ZN(n4869)
         );
  OAI21_X1 U5975 ( .B1(n5932), .B2(n4864), .A(n5773), .ZN(n5914) );
  INV_X1 U5976 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6659) );
  AND3_X1 U5977 ( .A1(n5963), .A2(n6659), .A3(n4864), .ZN(n5917) );
  OAI21_X1 U5978 ( .B1(n5914), .B2(n5917), .A(REIP_REG_10__SCAN_IN), .ZN(n4867) );
  OR3_X1 U5979 ( .A1(n5932), .A2(REIP_REG_10__SCAN_IN), .A3(n4865), .ZN(n4866)
         );
  OAI211_X1 U5980 ( .C1(n5973), .C2(n5143), .A(n4867), .B(n4866), .ZN(n4868)
         );
  NOR2_X1 U5981 ( .A1(n4869), .A2(n4868), .ZN(n4870) );
  OAI21_X1 U5982 ( .B1(n5147), .B2(n5776), .A(n4870), .ZN(U2817) );
  AOI22_X1 U5983 ( .A1(n6005), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n5999), .ZN(n4871) );
  OAI21_X1 U5984 ( .B1(n5147), .B2(n6011), .A(n4871), .ZN(U2881) );
  AOI22_X1 U5985 ( .A1(n6135), .A2(n5980), .B1(EBX_REG_10__SCAN_IN), .B2(n5387), .ZN(n4872) );
  OAI21_X1 U5986 ( .B1(n5147), .B2(n5389), .A(n4872), .ZN(U2849) );
  INV_X1 U5987 ( .A(n6516), .ZN(n6721) );
  OAI22_X1 U5988 ( .A1(n6721), .A2(n4873), .B1(n6727), .B2(n4946), .ZN(n4874)
         );
  AOI21_X1 U5989 ( .B1(n6364), .B2(n4944), .A(n4874), .ZN(n4876) );
  NAND2_X1 U5990 ( .A1(n6225), .A2(n6515), .ZN(n4875) );
  OAI211_X1 U5991 ( .C1(n4950), .C2(n6919), .A(n4876), .B(n4875), .ZN(U3020)
         );
  NAND2_X1 U5992 ( .A1(n6441), .A2(n4686), .ZN(n6512) );
  INV_X1 U5993 ( .A(n6512), .ZN(n4878) );
  INV_X1 U5994 ( .A(n4999), .ZN(n4877) );
  AOI21_X1 U5995 ( .B1(n4878), .B2(n6296), .A(n4877), .ZN(n4883) );
  OAI22_X1 U5996 ( .A1(n4883), .A2(n6519), .B1(n6505), .B2(n4879), .ZN(n4893)
         );
  INV_X1 U5997 ( .A(n4893), .ZN(n5000) );
  INV_X1 U5998 ( .A(n6540), .ZN(n5114) );
  OAI22_X1 U5999 ( .A1(n6544), .A2(n5000), .B1(n4999), .B2(n5114), .ZN(n4880)
         );
  AOI21_X1 U6000 ( .B1(n6541), .B2(n5002), .A(n4880), .ZN(n4888) );
  OAI21_X1 U6001 ( .B1(n4882), .B2(n5494), .A(n6508), .ZN(n4884) );
  NAND2_X1 U6002 ( .A1(n4884), .A2(n4883), .ZN(n4885) );
  OAI211_X1 U6003 ( .C1(n4886), .C2(n6506), .A(n6521), .B(n4885), .ZN(n5003)
         );
  NAND2_X1 U6004 ( .A1(n5003), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4887)
         );
  OAI211_X1 U6005 ( .C1(n5006), .C2(n6386), .A(n4888), .B(n4887), .ZN(U3143)
         );
  INV_X1 U6006 ( .A(n6566), .ZN(n5126) );
  OAI22_X1 U6007 ( .A1(n6572), .A2(n5000), .B1(n4999), .B2(n5126), .ZN(n4889)
         );
  AOI21_X1 U6008 ( .B1(n6568), .B2(n5002), .A(n4889), .ZN(n4891) );
  NAND2_X1 U6009 ( .A1(n5003), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4890)
         );
  OAI211_X1 U6010 ( .C1(n5006), .C2(n6406), .A(n4891), .B(n4890), .ZN(U3147)
         );
  NAND2_X1 U6011 ( .A1(n5003), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4895)
         );
  OAI22_X1 U6012 ( .A1(n6721), .A2(n4999), .B1(n6726), .B2(n4946), .ZN(n4892)
         );
  AOI21_X1 U6013 ( .B1(n6364), .B2(n4893), .A(n4892), .ZN(n4894) );
  OAI211_X1 U6014 ( .C1(n5006), .C2(n6727), .A(n4895), .B(n4894), .ZN(U3140)
         );
  INV_X1 U6015 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4900) );
  NAND2_X1 U6016 ( .A1(n6113), .A2(DATAI_29_), .ZN(n6394) );
  INV_X1 U6017 ( .A(DATAI_21_), .ZN(n4896) );
  NOR2_X1 U6018 ( .A1(n5494), .A2(n4896), .ZN(n6553) );
  INV_X1 U6019 ( .A(n6553), .ZN(n6317) );
  NAND2_X1 U6020 ( .A1(DATAI_5_), .A2(n4940), .ZN(n6556) );
  NOR2_X2 U6021 ( .A1(n4942), .A2(n3402), .ZN(n6552) );
  AOI22_X1 U6022 ( .A1(n6391), .A2(n4977), .B1(n6552), .B2(n4976), .ZN(n4897)
         );
  OAI21_X1 U6023 ( .B1(n6317), .B2(n5006), .A(n4897), .ZN(n4898) );
  AOI21_X1 U6024 ( .B1(n6551), .B2(n6567), .A(n4898), .ZN(n4899) );
  OAI21_X1 U6025 ( .B1(n4982), .B2(n4900), .A(n4899), .ZN(U3137) );
  INV_X1 U6026 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4905) );
  NAND2_X1 U6027 ( .A1(n6113), .A2(DATAI_28_), .ZN(n6390) );
  INV_X1 U6028 ( .A(DATAI_20_), .ZN(n4901) );
  NOR2_X1 U6029 ( .A1(n5494), .A2(n4901), .ZN(n6545) );
  INV_X1 U6030 ( .A(n6545), .ZN(n6314) );
  NAND2_X1 U6031 ( .A1(DATAI_4_), .A2(n4940), .ZN(n6550) );
  NOR2_X2 U6032 ( .A1(n4942), .A2(n3455), .ZN(n6546) );
  AOI22_X1 U6033 ( .A1(n6387), .A2(n4977), .B1(n6546), .B2(n4976), .ZN(n4902)
         );
  OAI21_X1 U6034 ( .B1(n6314), .B2(n5006), .A(n4902), .ZN(n4903) );
  AOI21_X1 U6035 ( .B1(n6547), .B2(n6567), .A(n4903), .ZN(n4904) );
  OAI21_X1 U6036 ( .B1(n4982), .B2(n4905), .A(n4904), .ZN(U3136) );
  OR2_X1 U6037 ( .A1(n4907), .A2(n3431), .ZN(n4906) );
  NAND2_X1 U6038 ( .A1(n5776), .A2(n4906), .ZN(n5969) );
  INV_X1 U6039 ( .A(n5969), .ZN(n5102) );
  NOR2_X1 U6040 ( .A1(n4907), .A2(n3449), .ZN(n5962) );
  NAND2_X1 U6041 ( .A1(n5962), .A2(n4686), .ZN(n4909) );
  OAI21_X1 U6042 ( .B1(n5960), .B2(n5939), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4908) );
  OAI211_X1 U6043 ( .C1(n5958), .C2(n4910), .A(n4909), .B(n4908), .ZN(n4913)
         );
  NOR2_X1 U6044 ( .A1(n5746), .A2(n4911), .ZN(n4912) );
  AOI211_X1 U6045 ( .C1(REIP_REG_0__SCAN_IN), .C2(n4914), .A(n4913), .B(n4912), 
        .ZN(n4915) );
  OAI21_X1 U6046 ( .B1(n5102), .B2(n6012), .A(n4915), .ZN(U2827) );
  AOI22_X1 U6047 ( .A1(n6387), .A2(n4944), .B1(n6546), .B2(n4943), .ZN(n4916)
         );
  OAI21_X1 U6048 ( .B1(n6390), .B2(n4946), .A(n4916), .ZN(n4917) );
  AOI21_X1 U6049 ( .B1(n6545), .B2(n6225), .A(n4917), .ZN(n4918) );
  OAI21_X1 U6050 ( .B1(n4950), .B2(n4919), .A(n4918), .ZN(U3024) );
  AOI22_X1 U6051 ( .A1(n6391), .A2(n4944), .B1(n6552), .B2(n4943), .ZN(n4920)
         );
  OAI21_X1 U6052 ( .B1(n6394), .B2(n4946), .A(n4920), .ZN(n4921) );
  AOI21_X1 U6053 ( .B1(n6553), .B2(n6225), .A(n4921), .ZN(n4922) );
  OAI21_X1 U6054 ( .B1(n4950), .B2(n4923), .A(n4922), .ZN(U3025) );
  INV_X1 U6055 ( .A(DATAI_17_), .ZN(n4924) );
  NOR2_X1 U6056 ( .A1(n5494), .A2(n4924), .ZN(n6529) );
  INV_X1 U6057 ( .A(DATAI_25_), .ZN(n4925) );
  NOR2_X2 U6058 ( .A1(n5494), .A2(n4925), .ZN(n6527) );
  INV_X1 U6059 ( .A(n6527), .ZN(n6378) );
  NAND2_X1 U6060 ( .A1(DATAI_1_), .A2(n4940), .ZN(n6532) );
  NOR2_X2 U6061 ( .A1(n4942), .A2(n4926), .ZN(n6528) );
  AOI22_X1 U6062 ( .A1(n6375), .A2(n4944), .B1(n6528), .B2(n4943), .ZN(n4927)
         );
  OAI21_X1 U6063 ( .B1(n6378), .B2(n4946), .A(n4927), .ZN(n4928) );
  AOI21_X1 U6064 ( .B1(n6529), .B2(n6225), .A(n4928), .ZN(n4929) );
  OAI21_X1 U6065 ( .B1(n4950), .B2(n4930), .A(n4929), .ZN(U3021) );
  INV_X1 U6066 ( .A(DATAI_22_), .ZN(n4931) );
  NOR2_X1 U6067 ( .A1(n5494), .A2(n4931), .ZN(n6559) );
  INV_X1 U6068 ( .A(DATAI_30_), .ZN(n4932) );
  NOR2_X2 U6069 ( .A1(n5494), .A2(n4932), .ZN(n6557) );
  INV_X1 U6070 ( .A(n6557), .ZN(n6398) );
  NAND2_X1 U6071 ( .A1(DATAI_6_), .A2(n4940), .ZN(n6562) );
  NOR2_X2 U6072 ( .A1(n4942), .A2(n4933), .ZN(n6558) );
  AOI22_X1 U6073 ( .A1(n6395), .A2(n4944), .B1(n6558), .B2(n4943), .ZN(n4934)
         );
  OAI21_X1 U6074 ( .B1(n6398), .B2(n4946), .A(n4934), .ZN(n4935) );
  AOI21_X1 U6075 ( .B1(n6559), .B2(n6225), .A(n4935), .ZN(n4936) );
  OAI21_X1 U6076 ( .B1(n4950), .B2(n4937), .A(n4936), .ZN(U3026) );
  INV_X1 U6077 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4949) );
  INV_X1 U6078 ( .A(DATAI_18_), .ZN(n4938) );
  NOR2_X1 U6079 ( .A1(n5494), .A2(n4938), .ZN(n6535) );
  INV_X1 U6080 ( .A(DATAI_26_), .ZN(n4939) );
  NOR2_X2 U6081 ( .A1(n5494), .A2(n4939), .ZN(n6533) );
  INV_X1 U6082 ( .A(n6533), .ZN(n6382) );
  NAND2_X1 U6083 ( .A1(DATAI_2_), .A2(n4940), .ZN(n6538) );
  NOR2_X2 U6084 ( .A1(n4942), .A2(n4941), .ZN(n6534) );
  AOI22_X1 U6085 ( .A1(n6379), .A2(n4944), .B1(n6534), .B2(n4943), .ZN(n4945)
         );
  OAI21_X1 U6086 ( .B1(n6382), .B2(n4946), .A(n4945), .ZN(n4947) );
  AOI21_X1 U6087 ( .B1(n6535), .B2(n6225), .A(n4947), .ZN(n4948) );
  OAI21_X1 U6088 ( .B1(n4950), .B2(n4949), .A(n4948), .ZN(U3022) );
  INV_X1 U6089 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4954) );
  INV_X1 U6090 ( .A(n6535), .ZN(n6308) );
  AOI22_X1 U6091 ( .A1(n6379), .A2(n4977), .B1(n6534), .B2(n4976), .ZN(n4951)
         );
  OAI21_X1 U6092 ( .B1(n6308), .B2(n5006), .A(n4951), .ZN(n4952) );
  AOI21_X1 U6093 ( .B1(n6533), .B2(n6567), .A(n4952), .ZN(n4953) );
  OAI21_X1 U6094 ( .B1(n4982), .B2(n4954), .A(n4953), .ZN(U3134) );
  INV_X1 U6095 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4958) );
  INV_X1 U6096 ( .A(n6559), .ZN(n6320) );
  AOI22_X1 U6097 ( .A1(n6395), .A2(n4977), .B1(n6558), .B2(n4976), .ZN(n4955)
         );
  OAI21_X1 U6098 ( .B1(n6320), .B2(n5006), .A(n4955), .ZN(n4956) );
  AOI21_X1 U6099 ( .B1(n6557), .B2(n6567), .A(n4956), .ZN(n4957) );
  OAI21_X1 U6100 ( .B1(n4982), .B2(n4958), .A(n4957), .ZN(U3138) );
  INV_X1 U6101 ( .A(n6546), .ZN(n5122) );
  OAI22_X1 U6102 ( .A1(n6550), .A2(n5000), .B1(n4999), .B2(n5122), .ZN(n4959)
         );
  AOI21_X1 U6103 ( .B1(n6545), .B2(n5002), .A(n4959), .ZN(n4961) );
  NAND2_X1 U6104 ( .A1(n5003), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4960)
         );
  OAI211_X1 U6105 ( .C1(n5006), .C2(n6390), .A(n4961), .B(n4960), .ZN(U3144)
         );
  INV_X1 U6106 ( .A(n6552), .ZN(n5118) );
  OAI22_X1 U6107 ( .A1(n6556), .A2(n5000), .B1(n4999), .B2(n5118), .ZN(n4962)
         );
  AOI21_X1 U6108 ( .B1(n6553), .B2(n5002), .A(n4962), .ZN(n4964) );
  NAND2_X1 U6109 ( .A1(n5003), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4963)
         );
  OAI211_X1 U6110 ( .C1(n5006), .C2(n6394), .A(n4964), .B(n4963), .ZN(U3145)
         );
  INV_X1 U6111 ( .A(n6528), .ZN(n5139) );
  OAI22_X1 U6112 ( .A1(n6532), .A2(n5000), .B1(n4999), .B2(n5139), .ZN(n4965)
         );
  AOI21_X1 U6113 ( .B1(n6529), .B2(n5002), .A(n4965), .ZN(n4967) );
  NAND2_X1 U6114 ( .A1(n5003), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4966)
         );
  OAI211_X1 U6115 ( .C1(n5006), .C2(n6378), .A(n4967), .B(n4966), .ZN(U3141)
         );
  INV_X1 U6116 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4971) );
  AOI22_X1 U6117 ( .A1(n6387), .A2(n5016), .B1(n5015), .B2(n6546), .ZN(n4968)
         );
  OAI21_X1 U6118 ( .B1(n6314), .B2(n5018), .A(n4968), .ZN(n4969) );
  AOI21_X1 U6119 ( .B1(n6547), .B2(n6499), .A(n4969), .ZN(n4970) );
  OAI21_X1 U6120 ( .B1(n5022), .B2(n4971), .A(n4970), .ZN(U3120) );
  INV_X1 U6121 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4975) );
  AOI22_X1 U6122 ( .A1(n6391), .A2(n5016), .B1(n5015), .B2(n6552), .ZN(n4972)
         );
  OAI21_X1 U6123 ( .B1(n6317), .B2(n5018), .A(n4972), .ZN(n4973) );
  AOI21_X1 U6124 ( .B1(n6551), .B2(n6499), .A(n4973), .ZN(n4974) );
  OAI21_X1 U6125 ( .B1(n5022), .B2(n4975), .A(n4974), .ZN(U3121) );
  INV_X1 U6126 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4981) );
  INV_X1 U6127 ( .A(n6529), .ZN(n6305) );
  AOI22_X1 U6128 ( .A1(n6375), .A2(n4977), .B1(n6528), .B2(n4976), .ZN(n4978)
         );
  OAI21_X1 U6129 ( .B1(n6305), .B2(n5006), .A(n4978), .ZN(n4979) );
  AOI21_X1 U6130 ( .B1(n6527), .B2(n6567), .A(n4979), .ZN(n4980) );
  OAI21_X1 U6131 ( .B1(n4982), .B2(n4981), .A(n4980), .ZN(U3133) );
  INV_X1 U6132 ( .A(n6179), .ZN(n4986) );
  AOI22_X1 U6133 ( .A1(n4983), .A2(n5939), .B1(n5960), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4985) );
  NAND2_X1 U6134 ( .A1(n5962), .A2(n6441), .ZN(n4984) );
  OAI211_X1 U6135 ( .C1(n5958), .C2(n4986), .A(n4985), .B(n4984), .ZN(n4993)
         );
  INV_X1 U6136 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6649) );
  AOI211_X1 U6137 ( .C1(n5963), .C2(n6647), .A(n5959), .B(n6649), .ZN(n5093)
         );
  INV_X1 U6138 ( .A(n5093), .ZN(n4991) );
  INV_X1 U6139 ( .A(n4987), .ZN(n4988) );
  NAND2_X1 U6140 ( .A1(n5963), .A2(n4988), .ZN(n4990) );
  NAND2_X1 U6141 ( .A1(n4990), .A2(n5773), .ZN(n5953) );
  INV_X1 U6142 ( .A(n5953), .ZN(n4989) );
  OAI22_X1 U6143 ( .A1(n4991), .A2(n4990), .B1(n4615), .B2(n4989), .ZN(n4992)
         );
  AOI211_X1 U6144 ( .C1(EBX_REG_3__SCAN_IN), .C2(n5968), .A(n4993), .B(n4992), 
        .ZN(n4994) );
  OAI21_X1 U6145 ( .B1(n4995), .B2(n5102), .A(n4994), .ZN(U2824) );
  INV_X1 U6146 ( .A(n6558), .ZN(n5130) );
  OAI22_X1 U6147 ( .A1(n6562), .A2(n5000), .B1(n4999), .B2(n5130), .ZN(n4996)
         );
  AOI21_X1 U6148 ( .B1(n6559), .B2(n5002), .A(n4996), .ZN(n4998) );
  NAND2_X1 U6149 ( .A1(n5003), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4997)
         );
  OAI211_X1 U6150 ( .C1(n5006), .C2(n6398), .A(n4998), .B(n4997), .ZN(U3146)
         );
  INV_X1 U6151 ( .A(n6534), .ZN(n5134) );
  OAI22_X1 U6152 ( .A1(n6538), .A2(n5000), .B1(n4999), .B2(n5134), .ZN(n5001)
         );
  AOI21_X1 U6153 ( .B1(n6535), .B2(n5002), .A(n5001), .ZN(n5005) );
  NAND2_X1 U6154 ( .A1(n5003), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n5004)
         );
  OAI211_X1 U6155 ( .C1(n5006), .C2(n6382), .A(n5005), .B(n5004), .ZN(U3142)
         );
  INV_X1 U6156 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5010) );
  AOI22_X1 U6157 ( .A1(n6395), .A2(n5016), .B1(n5015), .B2(n6558), .ZN(n5007)
         );
  OAI21_X1 U6158 ( .B1(n6320), .B2(n5018), .A(n5007), .ZN(n5008) );
  AOI21_X1 U6159 ( .B1(n6557), .B2(n6499), .A(n5008), .ZN(n5009) );
  OAI21_X1 U6160 ( .B1(n5022), .B2(n5010), .A(n5009), .ZN(U3122) );
  INV_X1 U6161 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5014) );
  AOI22_X1 U6162 ( .A1(n6379), .A2(n5016), .B1(n5015), .B2(n6534), .ZN(n5011)
         );
  OAI21_X1 U6163 ( .B1(n6308), .B2(n5018), .A(n5011), .ZN(n5012) );
  AOI21_X1 U6164 ( .B1(n6533), .B2(n6499), .A(n5012), .ZN(n5013) );
  OAI21_X1 U6165 ( .B1(n5022), .B2(n5014), .A(n5013), .ZN(U3118) );
  INV_X1 U6166 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5021) );
  AOI22_X1 U6167 ( .A1(n6375), .A2(n5016), .B1(n5015), .B2(n6528), .ZN(n5017)
         );
  OAI21_X1 U6168 ( .B1(n6305), .B2(n5018), .A(n5017), .ZN(n5019) );
  AOI21_X1 U6169 ( .B1(n6527), .B2(n6499), .A(n5019), .ZN(n5020) );
  OAI21_X1 U6170 ( .B1(n5022), .B2(n5021), .A(n5020), .ZN(U3117) );
  AOI21_X1 U6171 ( .B1(n5025), .B2(n4849), .A(n5024), .ZN(n6089) );
  INV_X1 U6172 ( .A(n6089), .ZN(n5074) );
  AND2_X1 U6173 ( .A1(n5027), .A2(n5026), .ZN(n5028) );
  NOR2_X1 U6174 ( .A1(n5150), .A2(n5028), .ZN(n5905) );
  AOI22_X1 U6175 ( .A1(n5905), .A2(n5980), .B1(EBX_REG_11__SCAN_IN), .B2(n5387), .ZN(n5029) );
  OAI21_X1 U6176 ( .B1(n5074), .B2(n5389), .A(n5029), .ZN(U2848) );
  OR2_X1 U6177 ( .A1(n6410), .A2(n6338), .ZN(n5030) );
  NOR2_X1 U6178 ( .A1(n6511), .A2(n5031), .ZN(n6262) );
  NAND2_X1 U6179 ( .A1(n6514), .A2(n6589), .ZN(n6259) );
  NOR2_X1 U6180 ( .A1(n6580), .A2(n6259), .ZN(n5065) );
  AOI21_X1 U6181 ( .B1(n6262), .B2(n4686), .A(n5065), .ZN(n5034) );
  INV_X1 U6182 ( .A(n6259), .ZN(n5032) );
  OAI21_X1 U6183 ( .B1(n6506), .B2(n5032), .A(n6521), .ZN(n5033) );
  INV_X1 U6184 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n5040) );
  INV_X1 U6185 ( .A(n6264), .ZN(n5035) );
  OAI22_X1 U6186 ( .A1(n5035), .A2(n5034), .B1(n6505), .B2(n6259), .ZN(n5068)
         );
  INV_X1 U6187 ( .A(n6338), .ZN(n6329) );
  AOI22_X1 U6188 ( .A1(n6552), .A2(n5065), .B1(n6551), .B2(n6283), .ZN(n5037)
         );
  OAI21_X1 U6189 ( .B1(n6293), .B2(n6317), .A(n5037), .ZN(n5038) );
  AOI21_X1 U6190 ( .B1(n6391), .B2(n5068), .A(n5038), .ZN(n5039) );
  OAI21_X1 U6191 ( .B1(n5071), .B2(n5040), .A(n5039), .ZN(U3065) );
  INV_X1 U6192 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5044) );
  AOI22_X1 U6193 ( .A1(n6558), .A2(n5065), .B1(n6557), .B2(n6283), .ZN(n5041)
         );
  OAI21_X1 U6194 ( .B1(n6293), .B2(n6320), .A(n5041), .ZN(n5042) );
  AOI21_X1 U6195 ( .B1(n6395), .B2(n5068), .A(n5042), .ZN(n5043) );
  OAI21_X1 U6196 ( .B1(n5071), .B2(n5044), .A(n5043), .ZN(U3066) );
  INV_X1 U6197 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n5048) );
  AOI22_X1 U6198 ( .A1(n6534), .A2(n5065), .B1(n6533), .B2(n6283), .ZN(n5045)
         );
  OAI21_X1 U6199 ( .B1(n6293), .B2(n6308), .A(n5045), .ZN(n5046) );
  AOI21_X1 U6200 ( .B1(n6379), .B2(n5068), .A(n5046), .ZN(n5047) );
  OAI21_X1 U6201 ( .B1(n5071), .B2(n5048), .A(n5047), .ZN(U3062) );
  INV_X1 U6202 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n5052) );
  AOI22_X1 U6203 ( .A1(n6528), .A2(n5065), .B1(n6527), .B2(n6283), .ZN(n5049)
         );
  OAI21_X1 U6204 ( .B1(n6293), .B2(n6305), .A(n5049), .ZN(n5050) );
  AOI21_X1 U6205 ( .B1(n6375), .B2(n5068), .A(n5050), .ZN(n5051) );
  OAI21_X1 U6206 ( .B1(n5071), .B2(n5052), .A(n5051), .ZN(U3061) );
  INV_X1 U6207 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n5056) );
  AOI22_X1 U6208 ( .A1(n6546), .A2(n5065), .B1(n6547), .B2(n6283), .ZN(n5053)
         );
  OAI21_X1 U6209 ( .B1(n6293), .B2(n6314), .A(n5053), .ZN(n5054) );
  AOI21_X1 U6210 ( .B1(n6387), .B2(n5068), .A(n5054), .ZN(n5055) );
  OAI21_X1 U6211 ( .B1(n5071), .B2(n5056), .A(n5055), .ZN(U3064) );
  INV_X1 U6212 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n5060) );
  AOI22_X1 U6213 ( .A1(n6516), .A2(n5065), .B1(n6524), .B2(n6283), .ZN(n5057)
         );
  OAI21_X1 U6214 ( .B1(n6293), .B2(n6726), .A(n5057), .ZN(n5058) );
  AOI21_X1 U6215 ( .B1(n6364), .B2(n5068), .A(n5058), .ZN(n5059) );
  OAI21_X1 U6216 ( .B1(n5071), .B2(n5060), .A(n5059), .ZN(U3060) );
  INV_X1 U6217 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5064) );
  AOI22_X1 U6218 ( .A1(n6566), .A2(n5065), .B1(n6564), .B2(n6283), .ZN(n5061)
         );
  OAI21_X1 U6219 ( .B1(n6293), .B2(n6328), .A(n5061), .ZN(n5062) );
  AOI21_X1 U6220 ( .B1(n6401), .B2(n5068), .A(n5062), .ZN(n5063) );
  OAI21_X1 U6221 ( .B1(n5071), .B2(n5064), .A(n5063), .ZN(U3067) );
  INV_X1 U6222 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n5070) );
  AOI22_X1 U6223 ( .A1(n6540), .A2(n5065), .B1(n6539), .B2(n6283), .ZN(n5066)
         );
  OAI21_X1 U6224 ( .B1(n6293), .B2(n6311), .A(n5066), .ZN(n5067) );
  AOI21_X1 U6225 ( .B1(n6383), .B2(n5068), .A(n5067), .ZN(n5069) );
  OAI21_X1 U6226 ( .B1(n5071), .B2(n5070), .A(n5069), .ZN(U3063) );
  INV_X1 U6227 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5073) );
  OAI222_X1 U6228 ( .A1(n5074), .A2(n6011), .B1(n6010), .B2(n5073), .C1(n6009), 
        .C2(n5072), .ZN(U2880) );
  NAND2_X1 U6229 ( .A1(n5076), .A2(n5075), .ZN(n5078) );
  XOR2_X1 U6230 ( .A(n5078), .B(n5077), .Z(n5092) );
  INV_X1 U6231 ( .A(n5918), .ZN(n5080) );
  AOI22_X1 U6232 ( .A1(n6108), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .B1(n6187), 
        .B2(REIP_REG_9__SCAN_IN), .ZN(n5079) );
  OAI21_X1 U6233 ( .B1(n6117), .B2(n5080), .A(n5079), .ZN(n5081) );
  AOI21_X1 U6234 ( .B1(n6007), .B2(n6113), .A(n5081), .ZN(n5082) );
  OAI21_X1 U6235 ( .B1(n5092), .B2(n6092), .A(n5082), .ZN(U2977) );
  AOI22_X1 U6236 ( .A1(n5646), .A2(n5084), .B1(n5653), .B2(n5083), .ZN(n6158)
         );
  OAI21_X1 U6237 ( .B1(n5694), .B2(n6148), .A(n6158), .ZN(n6136) );
  OAI22_X1 U6238 ( .A1(n5915), .A2(n6119), .B1(n6659), .B2(n6177), .ZN(n5085)
         );
  AOI21_X1 U6239 ( .B1(n6136), .B2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n5085), 
        .ZN(n5091) );
  AOI21_X1 U6240 ( .B1(n5086), .B2(n6196), .A(n6190), .ZN(n6175) );
  NOR2_X1 U6241 ( .A1(n6175), .A2(n5087), .ZN(n6163) );
  NAND2_X1 U6242 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6163), .ZN(n6160)
         );
  NOR2_X1 U6243 ( .A1(n5088), .A2(n6160), .ZN(n6139) );
  NAND2_X1 U6244 ( .A1(n6139), .A2(n5089), .ZN(n5090) );
  OAI211_X1 U6245 ( .C1(n5092), .C2(n5721), .A(n5091), .B(n5090), .ZN(U3009)
         );
  NAND2_X1 U6246 ( .A1(n5963), .A2(REIP_REG_1__SCAN_IN), .ZN(n5094) );
  AOI21_X1 U6247 ( .B1(n6649), .B2(n5094), .A(n5093), .ZN(n5095) );
  AOI21_X1 U6248 ( .B1(n5960), .B2(PHYADDRPOINTER_REG_2__SCAN_IN), .A(n5095), 
        .ZN(n5096) );
  OAI21_X1 U6249 ( .B1(n5973), .B2(n6116), .A(n5096), .ZN(n5097) );
  AOI21_X1 U6250 ( .B1(n5098), .B2(n5962), .A(n5097), .ZN(n5099) );
  OAI21_X1 U6251 ( .B1(n5958), .B2(n6186), .A(n5099), .ZN(n5100) );
  AOI21_X1 U6252 ( .B1(EBX_REG_2__SCAN_IN), .B2(n5968), .A(n5100), .ZN(n5101)
         );
  OAI21_X1 U6253 ( .B1(n5103), .B2(n5102), .A(n5101), .ZN(U2825) );
  NAND2_X1 U6254 ( .A1(n5723), .A2(n5104), .ZN(n6438) );
  INV_X1 U6255 ( .A(n6438), .ZN(n5105) );
  INV_X1 U6256 ( .A(n6413), .ZN(n5106) );
  NAND2_X1 U6257 ( .A1(n6445), .A2(n6589), .ZN(n6235) );
  NOR2_X1 U6258 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6235), .ZN(n5112)
         );
  INV_X1 U6259 ( .A(n5112), .ZN(n6720) );
  INV_X1 U6260 ( .A(n4510), .ZN(n5961) );
  AND2_X1 U6261 ( .A1(n4536), .A2(n5961), .ZN(n6442) );
  INV_X1 U6262 ( .A(n6288), .ZN(n5107) );
  NOR2_X1 U6263 ( .A1(n6361), .A2(n5107), .ZN(n6443) );
  AOI22_X1 U6264 ( .A1(n6232), .A2(n6506), .B1(n6443), .B2(n6589), .ZN(n6722)
         );
  INV_X1 U6265 ( .A(n6232), .ZN(n5109) );
  OAI21_X1 U6266 ( .B1(n6724), .B2(n6253), .A(n6508), .ZN(n5108) );
  NAND2_X1 U6267 ( .A1(n5109), .A2(n5108), .ZN(n5111) );
  NOR2_X1 U6268 ( .A1(n6289), .A2(n5110), .ZN(n6449) );
  OAI221_X1 U6269 ( .B1(n5112), .B2(n4054), .C1(n5112), .C2(n5111), .A(n6449), 
        .ZN(n6731) );
  AOI22_X1 U6270 ( .A1(n6383), .A2(n5137), .B1(INSTQUEUE_REG_2__3__SCAN_IN), 
        .B2(n6731), .ZN(n5113) );
  OAI21_X1 U6271 ( .B1(n5114), .B2(n6720), .A(n5113), .ZN(n5115) );
  AOI21_X1 U6272 ( .B1(n6539), .B2(n6724), .A(n5115), .ZN(n5116) );
  OAI21_X1 U6273 ( .B1(n6311), .B2(n6725), .A(n5116), .ZN(U3039) );
  AOI22_X1 U6274 ( .A1(n6391), .A2(n5137), .B1(INSTQUEUE_REG_2__5__SCAN_IN), 
        .B2(n6731), .ZN(n5117) );
  OAI21_X1 U6275 ( .B1(n5118), .B2(n6720), .A(n5117), .ZN(n5119) );
  AOI21_X1 U6276 ( .B1(n6551), .B2(n6724), .A(n5119), .ZN(n5120) );
  OAI21_X1 U6277 ( .B1(n6317), .B2(n6725), .A(n5120), .ZN(U3041) );
  AOI22_X1 U6278 ( .A1(n6387), .A2(n5137), .B1(INSTQUEUE_REG_2__4__SCAN_IN), 
        .B2(n6731), .ZN(n5121) );
  OAI21_X1 U6279 ( .B1(n5122), .B2(n6720), .A(n5121), .ZN(n5123) );
  AOI21_X1 U6280 ( .B1(n6547), .B2(n6724), .A(n5123), .ZN(n5124) );
  OAI21_X1 U6281 ( .B1(n6314), .B2(n6725), .A(n5124), .ZN(U3040) );
  AOI22_X1 U6282 ( .A1(n6401), .A2(n5137), .B1(INSTQUEUE_REG_2__7__SCAN_IN), 
        .B2(n6731), .ZN(n5125) );
  OAI21_X1 U6283 ( .B1(n5126), .B2(n6720), .A(n5125), .ZN(n5127) );
  AOI21_X1 U6284 ( .B1(n6564), .B2(n6724), .A(n5127), .ZN(n5128) );
  OAI21_X1 U6285 ( .B1(n6328), .B2(n6725), .A(n5128), .ZN(U3043) );
  AOI22_X1 U6286 ( .A1(n6395), .A2(n5137), .B1(INSTQUEUE_REG_2__6__SCAN_IN), 
        .B2(n6731), .ZN(n5129) );
  OAI21_X1 U6287 ( .B1(n5130), .B2(n6720), .A(n5129), .ZN(n5131) );
  AOI21_X1 U6288 ( .B1(n6557), .B2(n6724), .A(n5131), .ZN(n5132) );
  OAI21_X1 U6289 ( .B1(n6320), .B2(n6725), .A(n5132), .ZN(U3042) );
  AOI22_X1 U6290 ( .A1(n6379), .A2(n5137), .B1(INSTQUEUE_REG_2__2__SCAN_IN), 
        .B2(n6731), .ZN(n5133) );
  OAI21_X1 U6291 ( .B1(n5134), .B2(n6720), .A(n5133), .ZN(n5135) );
  AOI21_X1 U6292 ( .B1(n6533), .B2(n6724), .A(n5135), .ZN(n5136) );
  OAI21_X1 U6293 ( .B1(n6308), .B2(n6725), .A(n5136), .ZN(U3038) );
  AOI22_X1 U6294 ( .A1(n6375), .A2(n5137), .B1(INSTQUEUE_REG_2__1__SCAN_IN), 
        .B2(n6731), .ZN(n5138) );
  OAI21_X1 U6295 ( .B1(n5139), .B2(n6720), .A(n5138), .ZN(n5140) );
  AOI21_X1 U6296 ( .B1(n6527), .B2(n6724), .A(n5140), .ZN(n5141) );
  OAI21_X1 U6297 ( .B1(n6305), .B2(n6725), .A(n5141), .ZN(U3037) );
  XNOR2_X1 U6298 ( .A(n5514), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5142)
         );
  XNOR2_X1 U6299 ( .A(n4132), .B(n5142), .ZN(n6137) );
  NAND2_X1 U6300 ( .A1(n6137), .A2(n4502), .ZN(n5146) );
  NOR2_X1 U6301 ( .A1(n6177), .A2(n6661), .ZN(n6134) );
  NOR2_X1 U6302 ( .A1(n6117), .A2(n5143), .ZN(n5144) );
  AOI211_X1 U6303 ( .C1(n6108), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6134), 
        .B(n5144), .ZN(n5145) );
  OAI211_X1 U6304 ( .C1(n5494), .C2(n5147), .A(n5146), .B(n5145), .ZN(U2976)
         );
  XOR2_X1 U6305 ( .A(n5148), .B(n5024), .Z(n5177) );
  NAND2_X1 U6306 ( .A1(n5963), .A2(n5157), .ZN(n5907) );
  NAND2_X1 U6307 ( .A1(n5907), .A2(n5773), .ZN(n5903) );
  NAND2_X1 U6308 ( .A1(n5903), .A2(REIP_REG_12__SCAN_IN), .ZN(n5162) );
  INV_X1 U6309 ( .A(n5174), .ZN(n5156) );
  NOR2_X1 U6310 ( .A1(n5150), .A2(n5149), .ZN(n5151) );
  OR2_X1 U6311 ( .A1(n3198), .A2(n5151), .ZN(n6120) );
  INV_X1 U6312 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5152) );
  OAI22_X1 U6313 ( .A1(n6120), .A2(n5958), .B1(n5152), .B2(n5934), .ZN(n5153)
         );
  INV_X1 U6314 ( .A(n5153), .ZN(n5154) );
  NAND2_X1 U6315 ( .A1(n5154), .A2(n5924), .ZN(n5155) );
  AOI21_X1 U6316 ( .B1(n5939), .B2(n5156), .A(n5155), .ZN(n5161) );
  NAND2_X1 U6317 ( .A1(n5968), .A2(EBX_REG_12__SCAN_IN), .ZN(n5160) );
  NOR2_X1 U6318 ( .A1(n5157), .A2(REIP_REG_12__SCAN_IN), .ZN(n5158) );
  AND2_X1 U6319 ( .A1(n5963), .A2(n5158), .ZN(n5899) );
  INV_X1 U6320 ( .A(n5899), .ZN(n5159) );
  NAND4_X1 U6321 ( .A1(n5162), .A2(n5161), .A3(n5160), .A4(n5159), .ZN(n5163)
         );
  AOI21_X1 U6322 ( .B1(n5177), .B2(n5929), .A(n5163), .ZN(n5164) );
  INV_X1 U6323 ( .A(n5164), .ZN(U2815) );
  INV_X1 U6324 ( .A(n5389), .ZN(n5987) );
  OAI22_X1 U6325 ( .A1(n6120), .A2(n5984), .B1(n5165), .B2(n5989), .ZN(n5166)
         );
  AOI21_X1 U6326 ( .B1(n5177), .B2(n5987), .A(n5166), .ZN(n5167) );
  INV_X1 U6327 ( .A(n5167), .ZN(U2847) );
  INV_X1 U6328 ( .A(n5169), .ZN(n5170) );
  NOR2_X1 U6329 ( .A1(n5171), .A2(n5170), .ZN(n5172) );
  XNOR2_X1 U6330 ( .A(n5168), .B(n5172), .ZN(n6122) );
  NAND2_X1 U6331 ( .A1(n6187), .A2(REIP_REG_12__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U6332 ( .A1(n6108), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5173)
         );
  OAI211_X1 U6333 ( .C1(n6117), .C2(n5174), .A(n6118), .B(n5173), .ZN(n5175)
         );
  AOI21_X1 U6334 ( .B1(n5177), .B2(n6113), .A(n5175), .ZN(n5176) );
  OAI21_X1 U6335 ( .B1(n6122), .B2(n6092), .A(n5176), .ZN(U2974) );
  INV_X1 U6336 ( .A(n5177), .ZN(n5179) );
  INV_X1 U6337 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5178) );
  OAI222_X1 U6338 ( .A1(n6009), .A2(n5180), .B1(n6011), .B2(n5179), .C1(n5178), 
        .C2(n6010), .ZN(U2879) );
  AOI22_X1 U6339 ( .A1(n5181), .A2(n5514), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n4132), .ZN(n5183) );
  XNOR2_X1 U6340 ( .A(n5514), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5182)
         );
  XNOR2_X1 U6341 ( .A(n5183), .B(n5182), .ZN(n6093) );
  INV_X1 U6342 ( .A(n6129), .ZN(n5711) );
  OAI22_X1 U6343 ( .A1(n6177), .A2(n6970), .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n5711), .ZN(n5184) );
  AOI21_X1 U6344 ( .B1(n5905), .B2(n6189), .A(n5184), .ZN(n5188) );
  NAND2_X1 U6345 ( .A1(n5646), .A2(n5706), .ZN(n5651) );
  NAND2_X1 U6346 ( .A1(n5653), .A2(n5826), .ZN(n5185) );
  INV_X1 U6347 ( .A(n6125), .ZN(n5186) );
  NAND2_X1 U6348 ( .A1(n5186), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5187) );
  OAI211_X1 U6349 ( .C1(n6093), .C2(n5721), .A(n5188), .B(n5187), .ZN(U3007)
         );
  NAND2_X1 U6350 ( .A1(n5191), .A2(n5190), .ZN(n5194) );
  AOI22_X1 U6351 ( .A1(n5997), .A2(DATAI_31_), .B1(n5999), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5193) );
  NAND2_X1 U6352 ( .A1(n5194), .A2(n5193), .ZN(U2860) );
  AOI21_X1 U6353 ( .B1(n6581), .B2(n5199), .A(n5201), .ZN(n5202) );
  OAI22_X1 U6354 ( .A1(n5197), .A2(n5196), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5195), .ZN(n6579) );
  OAI22_X1 U6355 ( .A1(n6858), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6610), .ZN(n5198) );
  AOI21_X1 U6356 ( .B1(n6579), .B2(n5199), .A(n5198), .ZN(n5200) );
  OAI22_X1 U6357 ( .A1(n5202), .A2(n3283), .B1(n5201), .B2(n5200), .ZN(U3461)
         );
  AND2_X1 U6358 ( .A1(n5203), .A2(n5210), .ZN(n5208) );
  INV_X1 U6359 ( .A(n5209), .ZN(n5205) );
  OR2_X1 U6360 ( .A1(n5205), .A2(n5204), .ZN(n5207) );
  NAND2_X1 U6361 ( .A1(n5211), .A2(n4223), .ZN(n5206) );
  OAI211_X1 U6362 ( .C1(n5208), .C2(n5209), .A(n5207), .B(n5206), .ZN(n6595)
         );
  OR2_X1 U6363 ( .A1(n5209), .A2(n3404), .ZN(n5214) );
  OAI21_X1 U6364 ( .B1(n5212), .B2(n5211), .A(n5210), .ZN(n5213) );
  NAND2_X1 U6365 ( .A1(n5214), .A2(n5213), .ZN(n5844) );
  AOI21_X1 U6366 ( .B1(n5215), .B2(n6633), .A(READY_N), .ZN(n6712) );
  NOR2_X1 U6367 ( .A1(n5844), .A2(n6712), .ZN(n6591) );
  INV_X1 U6368 ( .A(n6616), .ZN(n6614) );
  OR2_X1 U6369 ( .A1(n6591), .A2(n6614), .ZN(n5850) );
  MUX2_X1 U6370 ( .A(n6595), .B(MORE_REG_SCAN_IN), .S(n5850), .Z(U3471) );
  OAI22_X1 U6371 ( .A1(n5216), .A2(n5934), .B1(n5973), .B2(n5426), .ZN(n5217)
         );
  INV_X1 U6372 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6686) );
  NOR2_X1 U6373 ( .A1(n5228), .A2(n6686), .ZN(n5219) );
  OAI21_X1 U6374 ( .B1(n5219), .B2(REIP_REG_30__SCAN_IN), .A(n5218), .ZN(n5220) );
  INV_X1 U6375 ( .A(n5223), .ZN(n5224) );
  OAI211_X1 U6376 ( .C1(n5382), .C2(n5225), .A(n5237), .B(n5224), .ZN(n5226)
         );
  NAND2_X1 U6377 ( .A1(n5227), .A2(n5226), .ZN(n5348) );
  INV_X1 U6378 ( .A(n5348), .ZN(n5566) );
  NOR2_X1 U6379 ( .A1(n5228), .A2(REIP_REG_29__SCAN_IN), .ZN(n5232) );
  AOI22_X1 U6380 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n5960), .B1(n5939), 
        .B2(n5433), .ZN(n5230) );
  NAND2_X1 U6381 ( .A1(n5968), .A2(EBX_REG_29__SCAN_IN), .ZN(n5229) );
  OAI211_X1 U6382 ( .C1(n5241), .C2(n6686), .A(n5230), .B(n5229), .ZN(n5231)
         );
  AOI211_X1 U6383 ( .C1(n5566), .C2(n5904), .A(n5232), .B(n5231), .ZN(n5233)
         );
  OAI21_X1 U6384 ( .B1(n5438), .B2(n5776), .A(n5233), .ZN(U2798) );
  OR2_X1 U6385 ( .A1(n5253), .A2(n5235), .ZN(n5236) );
  NAND2_X1 U6386 ( .A1(n5237), .A2(n5236), .ZN(n5571) );
  INV_X1 U6387 ( .A(REIP_REG_28__SCAN_IN), .ZN(n5245) );
  INV_X1 U6388 ( .A(n5444), .ZN(n5238) );
  AOI22_X1 U6389 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n5960), .B1(n5939), 
        .B2(n5238), .ZN(n5240) );
  NAND2_X1 U6390 ( .A1(n5968), .A2(EBX_REG_28__SCAN_IN), .ZN(n5239) );
  OAI211_X1 U6391 ( .C1(n5241), .C2(n5245), .A(n5240), .B(n5239), .ZN(n5242)
         );
  INV_X1 U6392 ( .A(n5242), .ZN(n5248) );
  INV_X1 U6393 ( .A(n5293), .ZN(n5246) );
  INV_X1 U6394 ( .A(n5243), .ZN(n5244) );
  NAND4_X1 U6395 ( .A1(n5246), .A2(REIP_REG_27__SCAN_IN), .A3(n5245), .A4(
        n5244), .ZN(n5247) );
  OAI211_X1 U6396 ( .C1(n5571), .C2(n5958), .A(n5248), .B(n5247), .ZN(n5249)
         );
  AOI21_X1 U6397 ( .B1(n5446), .B2(n5929), .A(n5249), .ZN(n5250) );
  INV_X1 U6398 ( .A(n5250), .ZN(U2799) );
  AND2_X1 U6399 ( .A1(n5264), .A2(n5251), .ZN(n5252) );
  NOR2_X1 U6400 ( .A1(n5253), .A2(n5252), .ZN(n5580) );
  INV_X1 U6401 ( .A(n5268), .ZN(n5257) );
  INV_X1 U6402 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6684) );
  AOI22_X1 U6403 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n5960), .B1(n5939), 
        .B2(n5254), .ZN(n5256) );
  NAND2_X1 U6404 ( .A1(n5968), .A2(EBX_REG_27__SCAN_IN), .ZN(n5255) );
  OAI211_X1 U6405 ( .C1(n5257), .C2(n6684), .A(n5256), .B(n5255), .ZN(n5258)
         );
  AOI21_X1 U6406 ( .B1(n5580), .B2(n5904), .A(n5258), .ZN(n5261) );
  NAND2_X1 U6407 ( .A1(n5259), .A2(n6684), .ZN(n5260) );
  OAI211_X1 U6408 ( .C1(n5401), .C2(n5776), .A(n5261), .B(n5260), .ZN(U2800)
         );
  AOI21_X1 U6409 ( .B1(n5263), .B2(n5262), .A(n4052), .ZN(n5455) );
  INV_X1 U6410 ( .A(n5455), .ZN(n5404) );
  OAI22_X1 U6411 ( .A1(n5452), .A2(n5934), .B1(n5973), .B2(n5451), .ZN(n5266)
         );
  OAI21_X1 U6412 ( .B1(n3238), .B2(n3212), .A(n5264), .ZN(n5589) );
  NOR2_X1 U6413 ( .A1(n5589), .A2(n5958), .ZN(n5265) );
  AOI211_X1 U6414 ( .C1(EBX_REG_26__SCAN_IN), .C2(n5968), .A(n5266), .B(n5265), 
        .ZN(n5271) );
  INV_X1 U6415 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6984) );
  INV_X1 U6416 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5267) );
  NOR3_X1 U6417 ( .A1(n5293), .A2(n6984), .A3(n5267), .ZN(n5269) );
  OAI21_X1 U6418 ( .B1(n5269), .B2(REIP_REG_26__SCAN_IN), .A(n5268), .ZN(n5270) );
  OAI211_X1 U6419 ( .C1(n5404), .C2(n5776), .A(n5271), .B(n5270), .ZN(U2801)
         );
  XNOR2_X1 U6420 ( .A(REIP_REG_24__SCAN_IN), .B(REIP_REG_25__SCAN_IN), .ZN(
        n5284) );
  INV_X1 U6421 ( .A(n5262), .ZN(n5273) );
  AOI21_X1 U6422 ( .B1(n5274), .B2(n5272), .A(n5273), .ZN(n5463) );
  NAND2_X1 U6423 ( .A1(n5463), .A2(n5929), .ZN(n5283) );
  NAND2_X1 U6424 ( .A1(n5287), .A2(n5275), .ZN(n5276) );
  NAND2_X1 U6425 ( .A1(n5277), .A2(n5276), .ZN(n5598) );
  INV_X1 U6426 ( .A(n5598), .ZN(n5281) );
  INV_X1 U6427 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U6428 ( .A1(n5743), .A2(REIP_REG_25__SCAN_IN), .ZN(n5279) );
  AOI22_X1 U6429 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n5960), .B1(n5939), 
        .B2(n5459), .ZN(n5278) );
  OAI211_X1 U6430 ( .C1(n5746), .C2(n5353), .A(n5279), .B(n5278), .ZN(n5280)
         );
  AOI21_X1 U6431 ( .B1(n5281), .B2(n5904), .A(n5280), .ZN(n5282) );
  OAI211_X1 U6432 ( .C1(n5293), .C2(n5284), .A(n5283), .B(n5282), .ZN(U2802)
         );
  XOR2_X1 U6433 ( .A(n5286), .B(n5285), .Z(n5471) );
  INV_X1 U6434 ( .A(n5471), .ZN(n5410) );
  OAI21_X1 U6435 ( .B1(n5362), .B2(n5288), .A(n5287), .ZN(n5289) );
  INV_X1 U6436 ( .A(n5289), .ZN(n5612) );
  NAND2_X1 U6437 ( .A1(n5743), .A2(REIP_REG_24__SCAN_IN), .ZN(n5291) );
  AOI22_X1 U6438 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n5960), .B1(n5939), 
        .B2(n5470), .ZN(n5290) );
  OAI211_X1 U6439 ( .C1(n5292), .C2(n5746), .A(n5291), .B(n5290), .ZN(n5295)
         );
  NOR2_X1 U6440 ( .A1(n5293), .A2(REIP_REG_24__SCAN_IN), .ZN(n5294) );
  AOI211_X1 U6441 ( .C1(n5904), .C2(n5612), .A(n5295), .B(n5294), .ZN(n5296)
         );
  OAI21_X1 U6442 ( .B1(n5410), .B2(n5776), .A(n5296), .ZN(U2803) );
  OAI21_X1 U6443 ( .B1(n5297), .B2(n5299), .A(n5799), .ZN(n5996) );
  OAI21_X1 U6444 ( .B1(n5715), .B2(n5315), .A(n5300), .ZN(n5301) );
  NAND2_X1 U6445 ( .A1(n5301), .A2(n5683), .ZN(n5697) );
  INV_X1 U6446 ( .A(n5697), .ZN(n5310) );
  INV_X1 U6447 ( .A(n5531), .ZN(n5304) );
  NOR2_X1 U6448 ( .A1(n5932), .A2(n5302), .ZN(n5884) );
  OR2_X1 U6449 ( .A1(n5884), .A2(n5959), .ZN(n5886) );
  NAND2_X1 U6450 ( .A1(n5963), .A2(n5302), .ZN(n5875) );
  NOR2_X1 U6451 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5875), .ZN(n5318) );
  OAI21_X1 U6452 ( .B1(n5886), .B2(n5318), .A(REIP_REG_16__SCAN_IN), .ZN(n5303) );
  OAI21_X1 U6453 ( .B1(n5304), .B2(n5973), .A(n5303), .ZN(n5309) );
  NOR2_X1 U6454 ( .A1(REIP_REG_16__SCAN_IN), .A2(n5875), .ZN(n5305) );
  AOI22_X1 U6455 ( .A1(PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n5960), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5305), .ZN(n5306) );
  OAI211_X1 U6456 ( .C1(n5746), .C2(n5307), .A(n5306), .B(n5924), .ZN(n5308)
         );
  AOI211_X1 U6457 ( .C1(n5310), .C2(n5904), .A(n5309), .B(n5308), .ZN(n5311)
         );
  OAI21_X1 U6458 ( .B1(n5996), .B2(n5776), .A(n5311), .ZN(U2811) );
  AOI21_X1 U6459 ( .B1(n5314), .B2(n5313), .A(n5297), .ZN(n5539) );
  INV_X1 U6460 ( .A(n5539), .ZN(n5417) );
  XOR2_X1 U6461 ( .A(n5315), .B(n5715), .Z(n5818) );
  INV_X1 U6462 ( .A(n5886), .ZN(n5317) );
  INV_X1 U6463 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5316) );
  OAI22_X1 U6464 ( .A1(n5317), .A2(n5316), .B1(n5537), .B2(n5973), .ZN(n5322)
         );
  INV_X1 U6465 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5320) );
  AOI21_X1 U6466 ( .B1(EBX_REG_15__SCAN_IN), .B2(n5968), .A(n5318), .ZN(n5319)
         );
  OAI211_X1 U6467 ( .C1(n5934), .C2(n5320), .A(n5319), .B(n5924), .ZN(n5321)
         );
  AOI211_X1 U6468 ( .C1(n5904), .C2(n5818), .A(n5322), .B(n5321), .ZN(n5323)
         );
  OAI21_X1 U6469 ( .B1(n5417), .B2(n5776), .A(n5323), .ZN(U2812) );
  INV_X1 U6470 ( .A(n5333), .ZN(n5324) );
  NAND2_X1 U6471 ( .A1(n5963), .A2(n5324), .ZN(n5922) );
  OAI21_X1 U6472 ( .B1(n5339), .B2(n5922), .A(n6657), .ZN(n5330) );
  INV_X1 U6473 ( .A(n5924), .ZN(n5947) );
  NOR2_X1 U6474 ( .A1(n5973), .A2(n5325), .ZN(n5326) );
  AOI211_X1 U6475 ( .C1(n5960), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n5947), 
        .B(n5326), .ZN(n5328) );
  NAND2_X1 U6476 ( .A1(n5968), .A2(EBX_REG_8__SCAN_IN), .ZN(n5327) );
  OAI211_X1 U6477 ( .C1(n6143), .C2(n5958), .A(n5328), .B(n5327), .ZN(n5329)
         );
  AOI21_X1 U6478 ( .B1(n5330), .B2(n5914), .A(n5329), .ZN(n5331) );
  OAI21_X1 U6479 ( .B1(n5332), .B2(n5776), .A(n5331), .ZN(U2819) );
  NAND2_X1 U6480 ( .A1(n5963), .A2(n5333), .ZN(n5334) );
  AND2_X1 U6481 ( .A1(n5334), .A2(n5773), .ZN(n5944) );
  INV_X1 U6482 ( .A(n5944), .ZN(n5343) );
  INV_X1 U6483 ( .A(n6156), .ZN(n5338) );
  OAI21_X1 U6484 ( .B1(n5973), .B2(n5335), .A(n5924), .ZN(n5336) );
  AOI21_X1 U6485 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n5960), .A(n5336), 
        .ZN(n5337) );
  OAI21_X1 U6486 ( .B1(n5338), .B2(n5958), .A(n5337), .ZN(n5342) );
  OAI21_X1 U6487 ( .B1(REIP_REG_7__SCAN_IN), .B2(REIP_REG_6__SCAN_IN), .A(
        n5339), .ZN(n5340) );
  OAI22_X1 U6488 ( .A1(n5746), .A2(n6871), .B1(n5922), .B2(n5340), .ZN(n5341)
         );
  AOI211_X1 U6489 ( .C1(REIP_REG_7__SCAN_IN), .C2(n5343), .A(n5342), .B(n5341), 
        .ZN(n5344) );
  OAI21_X1 U6490 ( .B1(n5345), .B2(n5776), .A(n5344), .ZN(U2820) );
  OAI22_X1 U6491 ( .A1(n5347), .A2(n5984), .B1(n5989), .B2(n5346), .ZN(U2828)
         );
  INV_X1 U6492 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5349) );
  OAI222_X1 U6493 ( .A1(n5389), .A2(n5438), .B1(n5349), .B2(n5989), .C1(n5348), 
        .C2(n5984), .ZN(U2830) );
  INV_X1 U6494 ( .A(n5446), .ZN(n5398) );
  OAI222_X1 U6495 ( .A1(n5389), .A2(n5398), .B1(n5350), .B2(n5989), .C1(n5571), 
        .C2(n5984), .ZN(U2831) );
  AOI22_X1 U6496 ( .A1(n5580), .A2(n5980), .B1(EBX_REG_27__SCAN_IN), .B2(n5387), .ZN(n5351) );
  OAI21_X1 U6497 ( .B1(n5401), .B2(n5389), .A(n5351), .ZN(U2832) );
  OAI222_X1 U6498 ( .A1(n5389), .A2(n5404), .B1(n5352), .B2(n5989), .C1(n5589), 
        .C2(n5984), .ZN(U2833) );
  INV_X1 U6499 ( .A(n5463), .ZN(n5407) );
  OAI222_X1 U6500 ( .A1(n5407), .A2(n5389), .B1(n5353), .B2(n5989), .C1(n5598), 
        .C2(n5984), .ZN(U2834) );
  AOI22_X1 U6501 ( .A1(n5612), .A2(n5980), .B1(EBX_REG_24__SCAN_IN), .B2(n5387), .ZN(n5354) );
  OAI21_X1 U6502 ( .B1(n5410), .B2(n5389), .A(n5354), .ZN(U2835) );
  INV_X1 U6503 ( .A(n5285), .ZN(n5356) );
  INV_X1 U6504 ( .A(n5358), .ZN(n5368) );
  INV_X1 U6505 ( .A(n5359), .ZN(n5360) );
  AOI21_X1 U6506 ( .B1(n5374), .B2(n5368), .A(n5360), .ZN(n5361) );
  OR2_X1 U6507 ( .A1(n5362), .A2(n5361), .ZN(n5739) );
  OAI22_X1 U6508 ( .A1(n5739), .A2(n5984), .B1(n6939), .B2(n5989), .ZN(n5363)
         );
  INV_X1 U6509 ( .A(n5363), .ZN(n5364) );
  OAI21_X1 U6510 ( .B1(n5740), .B2(n5389), .A(n5364), .ZN(U2836) );
  AOI21_X1 U6511 ( .B1(n5367), .B2(n5366), .A(n5355), .ZN(n5789) );
  INV_X1 U6512 ( .A(n5789), .ZN(n5370) );
  INV_X1 U6513 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5369) );
  XNOR2_X1 U6514 ( .A(n5374), .B(n5368), .ZN(n5749) );
  OAI222_X1 U6515 ( .A1(n5389), .A2(n5370), .B1(n5369), .B2(n5989), .C1(n5984), 
        .C2(n5749), .ZN(U2837) );
  NAND2_X1 U6516 ( .A1(n5371), .A2(n5372), .ZN(n5373) );
  NAND2_X1 U6517 ( .A1(n5366), .A2(n5373), .ZN(n5759) );
  INV_X1 U6518 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5377) );
  AOI21_X1 U6519 ( .B1(n5376), .B2(n5375), .A(n5374), .ZN(n5760) );
  INV_X1 U6520 ( .A(n5760), .ZN(n5634) );
  OAI222_X1 U6521 ( .A1(n5389), .A2(n5759), .B1(n5377), .B2(n5989), .C1(n5634), 
        .C2(n5984), .ZN(U2838) );
  AND2_X1 U6522 ( .A1(n5379), .A2(n5380), .ZN(n5381) );
  NOR2_X1 U6523 ( .A1(n5378), .A2(n5381), .ZN(n5510) );
  INV_X1 U6524 ( .A(n5510), .ZN(n5777) );
  INV_X1 U6525 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5386) );
  INV_X1 U6526 ( .A(n5642), .ZN(n5384) );
  MUX2_X1 U6527 ( .A(n5384), .B(n5383), .S(n5382), .Z(n5670) );
  NAND2_X1 U6528 ( .A1(n5671), .A2(n5670), .ZN(n5669) );
  XNOR2_X1 U6529 ( .A(n5669), .B(n5385), .ZN(n5659) );
  INV_X1 U6530 ( .A(n5659), .ZN(n5775) );
  OAI222_X1 U6531 ( .A1(n5777), .A2(n5389), .B1(n5989), .B2(n5386), .C1(n5775), 
        .C2(n5984), .ZN(U2840) );
  OAI222_X1 U6532 ( .A1(n5697), .A2(n5984), .B1(n5307), .B2(n5989), .C1(n5996), 
        .C2(n5389), .ZN(U2843) );
  AOI22_X1 U6533 ( .A1(n5818), .A2(n5980), .B1(EBX_REG_15__SCAN_IN), .B2(n5387), .ZN(n5388) );
  OAI21_X1 U6534 ( .B1(n5417), .B2(n5389), .A(n5388), .ZN(U2844) );
  AOI22_X1 U6535 ( .A1(n5997), .A2(DATAI_30_), .B1(n5999), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5392) );
  AND2_X1 U6536 ( .A1(n3402), .A2(n3428), .ZN(n5390) );
  NAND2_X1 U6537 ( .A1(n6000), .A2(DATAI_14_), .ZN(n5391) );
  OAI211_X1 U6538 ( .C1(n5393), .C2(n6011), .A(n5392), .B(n5391), .ZN(U2861)
         );
  AOI22_X1 U6539 ( .A1(n5997), .A2(DATAI_29_), .B1(n5999), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U6540 ( .A1(n6000), .A2(DATAI_13_), .ZN(n5394) );
  OAI211_X1 U6541 ( .C1(n5438), .C2(n6011), .A(n5395), .B(n5394), .ZN(U2862)
         );
  AOI22_X1 U6542 ( .A1(n5997), .A2(DATAI_28_), .B1(n5999), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6543 ( .A1(n6000), .A2(DATAI_12_), .ZN(n5396) );
  OAI211_X1 U6544 ( .C1(n5398), .C2(n6011), .A(n5397), .B(n5396), .ZN(U2863)
         );
  AOI22_X1 U6545 ( .A1(n5997), .A2(DATAI_27_), .B1(n5999), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U6546 ( .A1(n6000), .A2(DATAI_11_), .ZN(n5399) );
  OAI211_X1 U6547 ( .C1(n5401), .C2(n6011), .A(n5400), .B(n5399), .ZN(U2864)
         );
  AOI22_X1 U6548 ( .A1(n5997), .A2(DATAI_26_), .B1(n5999), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U6549 ( .A1(n6000), .A2(DATAI_10_), .ZN(n5402) );
  OAI211_X1 U6550 ( .C1(n5404), .C2(n6011), .A(n5403), .B(n5402), .ZN(U2865)
         );
  AOI22_X1 U6551 ( .A1(n5997), .A2(DATAI_25_), .B1(n5999), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U6552 ( .A1(n6000), .A2(DATAI_9_), .ZN(n5405) );
  OAI211_X1 U6553 ( .C1(n5407), .C2(n6011), .A(n5406), .B(n5405), .ZN(U2866)
         );
  AOI22_X1 U6554 ( .A1(n5997), .A2(DATAI_24_), .B1(n5999), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5409) );
  NAND2_X1 U6555 ( .A1(n6000), .A2(DATAI_8_), .ZN(n5408) );
  OAI211_X1 U6556 ( .C1(n5410), .C2(n6011), .A(n5409), .B(n5408), .ZN(U2867)
         );
  AOI22_X1 U6557 ( .A1(n6000), .A2(DATAI_7_), .B1(n5999), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U6558 ( .A1(n5997), .A2(DATAI_23_), .ZN(n5411) );
  OAI211_X1 U6559 ( .C1(n5740), .C2(n6011), .A(n5412), .B(n5411), .ZN(U2868)
         );
  AOI22_X1 U6560 ( .A1(n6000), .A2(DATAI_3_), .B1(n5999), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5414) );
  NAND2_X1 U6561 ( .A1(n5997), .A2(DATAI_19_), .ZN(n5413) );
  OAI211_X1 U6562 ( .C1(n5777), .C2(n6011), .A(n5414), .B(n5413), .ZN(U2872)
         );
  OAI222_X1 U6563 ( .A1(n5417), .A2(n6011), .B1(n6010), .B2(n5416), .C1(n6009), 
        .C2(n5415), .ZN(U2876) );
  OAI21_X1 U6564 ( .B1(n5418), .B2(n5419), .A(n5313), .ZN(n5547) );
  INV_X1 U6565 ( .A(DATAI_14_), .ZN(n6061) );
  OAI222_X1 U6566 ( .A1(n5547), .A2(n6011), .B1(n6010), .B2(n6086), .C1(n6061), 
        .C2(n6009), .ZN(U2877) );
  NOR2_X1 U6567 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U6568 ( .A1(n5448), .A2(n5572), .ZN(n5430) );
  NOR3_X1 U6569 ( .A1(n5420), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5430), 
        .ZN(n5421) );
  INV_X1 U6570 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5423) );
  INV_X1 U6571 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6693) );
  NOR2_X1 U6572 ( .A1(n6177), .A2(n6693), .ZN(n5555) );
  AOI21_X1 U6573 ( .B1(n6108), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5555), 
        .ZN(n5425) );
  OAI21_X1 U6574 ( .B1(n5426), .B2(n6117), .A(n5425), .ZN(n5427) );
  AOI21_X1 U6575 ( .B1(n5428), .B2(n6113), .A(n5427), .ZN(n5429) );
  OAI21_X1 U6576 ( .B1(n5561), .B2(n6092), .A(n5429), .ZN(U2956) );
  INV_X1 U6577 ( .A(n5573), .ZN(n5563) );
  OAI22_X1 U6578 ( .A1(n5439), .A2(n5563), .B1(n5420), .B2(n5430), .ZN(n5431)
         );
  XNOR2_X1 U6579 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .B(n5431), .ZN(n5432)
         );
  INV_X1 U6580 ( .A(n5432), .ZN(n5562) );
  NAND2_X1 U6581 ( .A1(n5562), .A2(n4502), .ZN(n5437) );
  NOR2_X1 U6582 ( .A1(n6177), .A2(n6686), .ZN(n5565) );
  INV_X1 U6583 ( .A(n5433), .ZN(n5434) );
  NOR2_X1 U6584 ( .A1(n6117), .A2(n5434), .ZN(n5435) );
  AOI211_X1 U6585 ( .C1(n6108), .C2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5565), 
        .B(n5435), .ZN(n5436) );
  OAI211_X1 U6586 ( .C1(n5494), .C2(n5438), .A(n5437), .B(n5436), .ZN(U2957)
         );
  OAI22_X1 U6587 ( .A1(n3253), .A2(n5440), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5592), .ZN(n5442) );
  XNOR2_X1 U6588 ( .A(n5442), .B(n5441), .ZN(n5579) );
  NAND2_X1 U6589 ( .A1(n6187), .A2(REIP_REG_28__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U6590 ( .A1(n6108), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5443)
         );
  OAI211_X1 U6591 ( .C1(n6117), .C2(n5444), .A(n5570), .B(n5443), .ZN(n5445)
         );
  AOI21_X1 U6592 ( .B1(n5446), .B2(n6113), .A(n5445), .ZN(n5447) );
  OAI21_X1 U6593 ( .B1(n5579), .B2(n6092), .A(n5447), .ZN(U2958) );
  NOR2_X1 U6594 ( .A1(n5449), .A2(n5448), .ZN(n5450) );
  XOR2_X1 U6595 ( .A(n5450), .B(n5420), .Z(n5596) );
  NOR2_X1 U6596 ( .A1(n6117), .A2(n5451), .ZN(n5454) );
  NAND2_X1 U6597 ( .A1(n6187), .A2(REIP_REG_26__SCAN_IN), .ZN(n5588) );
  OAI21_X1 U6598 ( .B1(n5528), .B2(n5452), .A(n5588), .ZN(n5453) );
  AOI211_X1 U6599 ( .C1(n5455), .C2(n6113), .A(n5454), .B(n5453), .ZN(n5456)
         );
  OAI21_X1 U6600 ( .B1(n5596), .B2(n6092), .A(n5456), .ZN(U2960) );
  AOI21_X1 U6601 ( .B1(n5458), .B2(n5457), .A(n4143), .ZN(n5603) );
  INV_X1 U6602 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U6603 ( .A1(n6088), .A2(n5459), .ZN(n5460) );
  NAND2_X1 U6604 ( .A1(n6187), .A2(REIP_REG_25__SCAN_IN), .ZN(n5597) );
  OAI211_X1 U6605 ( .C1(n5528), .C2(n5461), .A(n5460), .B(n5597), .ZN(n5462)
         );
  AOI21_X1 U6606 ( .B1(n5463), .B2(n6113), .A(n5462), .ZN(n5464) );
  OAI21_X1 U6607 ( .B1(n5603), .B2(n6092), .A(n5464), .ZN(U2961) );
  AND2_X1 U6608 ( .A1(n5534), .A2(n5664), .ZN(n5504) );
  NAND2_X1 U6609 ( .A1(n5514), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5503) );
  XNOR2_X1 U6610 ( .A(n5534), .B(n6933), .ZN(n5496) );
  XNOR2_X1 U6611 ( .A(n5534), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5489)
         );
  INV_X1 U6612 ( .A(n5488), .ZN(n5465) );
  NOR2_X1 U6613 ( .A1(n5534), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5482)
         );
  NAND2_X1 U6614 ( .A1(n5465), .A2(n5482), .ZN(n5474) );
  OAI21_X1 U6615 ( .B1(n5514), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5488), 
        .ZN(n5484) );
  NAND3_X1 U6616 ( .A1(n5534), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5466) );
  XNOR2_X1 U6617 ( .A(n5467), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5614)
         );
  NOR2_X1 U6618 ( .A1(n6177), .A2(n6984), .ZN(n5611) );
  NOR2_X1 U6619 ( .A1(n5528), .A2(n5468), .ZN(n5469) );
  AOI211_X1 U6620 ( .C1(n6088), .C2(n5470), .A(n5611), .B(n5469), .ZN(n5473)
         );
  NAND2_X1 U6621 ( .A1(n5471), .A2(n6113), .ZN(n5472) );
  OAI211_X1 U6622 ( .C1(n5614), .C2(n6092), .A(n5473), .B(n5472), .ZN(U2962)
         );
  NAND2_X1 U6623 ( .A1(n5534), .A2(n5605), .ZN(n5475) );
  OAI21_X1 U6624 ( .B1(n5476), .B2(n5475), .A(n5474), .ZN(n5477) );
  XNOR2_X1 U6625 ( .A(n5477), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5621)
         );
  INV_X1 U6626 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U6627 ( .A1(n6187), .A2(REIP_REG_23__SCAN_IN), .ZN(n5615) );
  OAI21_X1 U6628 ( .B1(n5528), .B2(n5478), .A(n5615), .ZN(n5480) );
  NOR2_X1 U6629 ( .A1(n5740), .A2(n5494), .ZN(n5479) );
  AOI211_X1 U6630 ( .C1(n6088), .C2(n5738), .A(n5480), .B(n5479), .ZN(n5481)
         );
  OAI21_X1 U6631 ( .B1(n5621), .B2(n6092), .A(n5481), .ZN(U2963) );
  AOI21_X1 U6632 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5534), .A(n5482), 
        .ZN(n5483) );
  XNOR2_X1 U6633 ( .A(n5484), .B(n5483), .ZN(n5631) );
  NAND2_X1 U6634 ( .A1(n6187), .A2(REIP_REG_22__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U6635 ( .A1(n6108), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5485)
         );
  OAI211_X1 U6636 ( .C1(n6117), .C2(n5747), .A(n5623), .B(n5485), .ZN(n5486)
         );
  AOI21_X1 U6637 ( .B1(n5789), .B2(n6113), .A(n5486), .ZN(n5487) );
  OAI21_X1 U6638 ( .B1(n5631), .B2(n6092), .A(n5487), .ZN(U2964) );
  OAI21_X1 U6639 ( .B1(n5490), .B2(n5489), .A(n5488), .ZN(n5632) );
  NAND2_X1 U6640 ( .A1(n5632), .A2(n4502), .ZN(n5493) );
  NAND2_X1 U6641 ( .A1(n6187), .A2(REIP_REG_21__SCAN_IN), .ZN(n5633) );
  OAI21_X1 U6642 ( .B1(n5528), .B2(n6864), .A(n5633), .ZN(n5491) );
  AOI21_X1 U6643 ( .B1(n6088), .B2(n5758), .A(n5491), .ZN(n5492) );
  OAI211_X1 U6644 ( .C1(n5494), .C2(n5759), .A(n5493), .B(n5492), .ZN(U2965)
         );
  XOR2_X1 U6645 ( .A(n5496), .B(n5495), .Z(n5658) );
  NAND2_X1 U6646 ( .A1(n6187), .A2(REIP_REG_20__SCAN_IN), .ZN(n5645) );
  OAI21_X1 U6647 ( .B1(n5528), .B2(n5497), .A(n5645), .ZN(n5501) );
  OR2_X1 U6648 ( .A1(n5378), .A2(n5498), .ZN(n5499) );
  NAND2_X1 U6649 ( .A1(n5371), .A2(n5499), .ZN(n5795) );
  NOR2_X1 U6650 ( .A1(n5795), .A2(n5494), .ZN(n5500) );
  AOI211_X1 U6651 ( .C1(n6088), .C2(n5768), .A(n5501), .B(n5500), .ZN(n5502)
         );
  OAI21_X1 U6652 ( .B1(n5658), .B2(n6092), .A(n5502), .ZN(U2966) );
  INV_X1 U6653 ( .A(n5503), .ZN(n5505) );
  NOR2_X1 U6654 ( .A1(n5505), .A2(n5504), .ZN(n5506) );
  XNOR2_X1 U6655 ( .A(n3205), .B(n5506), .ZN(n5667) );
  INV_X1 U6656 ( .A(n5780), .ZN(n5508) );
  NAND2_X1 U6657 ( .A1(n6187), .A2(REIP_REG_19__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U6658 ( .A1(n6108), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5507)
         );
  OAI211_X1 U6659 ( .C1(n6117), .C2(n5508), .A(n5661), .B(n5507), .ZN(n5509)
         );
  AOI21_X1 U6660 ( .B1(n5510), .B2(n6113), .A(n5509), .ZN(n5511) );
  OAI21_X1 U6661 ( .B1(n5667), .B2(n6092), .A(n5511), .ZN(U2967) );
  NAND3_X1 U6662 ( .A1(n5513), .A2(n5514), .A3(n5691), .ZN(n5679) );
  NOR3_X1 U6663 ( .A1(n5513), .A2(n5514), .A3(n5691), .ZN(n5681) );
  NAND2_X1 U6664 ( .A1(n5681), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5515) );
  OAI21_X1 U6665 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5679), .A(n5515), 
        .ZN(n5516) );
  XNOR2_X1 U6666 ( .A(n5516), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5678)
         );
  INV_X1 U6667 ( .A(n5379), .ZN(n5518) );
  AOI21_X1 U6668 ( .B1(n5519), .B2(n5517), .A(n5518), .ZN(n5990) );
  NAND2_X1 U6669 ( .A1(n6187), .A2(REIP_REG_18__SCAN_IN), .ZN(n5672) );
  NAND2_X1 U6670 ( .A1(n6108), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5520)
         );
  OAI211_X1 U6671 ( .C1(n6117), .C2(n5869), .A(n5672), .B(n5520), .ZN(n5521)
         );
  AOI21_X1 U6672 ( .B1(n5990), .B2(n6113), .A(n5521), .ZN(n5522) );
  OAI21_X1 U6673 ( .B1(n5678), .B2(n6092), .A(n5522), .ZN(U2968) );
  INV_X1 U6674 ( .A(n5523), .ZN(n5525) );
  NAND2_X1 U6675 ( .A1(n5525), .A2(n5524), .ZN(n5526) );
  XNOR2_X1 U6676 ( .A(n5513), .B(n5526), .ZN(n5702) );
  INV_X1 U6677 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U6678 ( .A1(n6187), .A2(REIP_REG_16__SCAN_IN), .ZN(n5695) );
  OAI21_X1 U6679 ( .B1(n5528), .B2(n5527), .A(n5695), .ZN(n5530) );
  NOR2_X1 U6680 ( .A1(n5996), .A2(n5494), .ZN(n5529) );
  AOI211_X1 U6681 ( .C1(n6088), .C2(n5531), .A(n5530), .B(n5529), .ZN(n5532)
         );
  OAI21_X1 U6682 ( .B1(n6092), .B2(n5702), .A(n5532), .ZN(U2970) );
  XNOR2_X1 U6683 ( .A(n5534), .B(n5692), .ZN(n5535) );
  XNOR2_X1 U6684 ( .A(n5533), .B(n5535), .ZN(n5820) );
  INV_X1 U6685 ( .A(n5820), .ZN(n5541) );
  NAND2_X1 U6686 ( .A1(n6187), .A2(REIP_REG_15__SCAN_IN), .ZN(n5816) );
  NAND2_X1 U6687 ( .A1(n6108), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5536)
         );
  OAI211_X1 U6688 ( .C1(n6117), .C2(n5537), .A(n5816), .B(n5536), .ZN(n5538)
         );
  AOI21_X1 U6689 ( .B1(n5539), .B2(n6113), .A(n5538), .ZN(n5540) );
  OAI21_X1 U6690 ( .B1(n5541), .B2(n6092), .A(n5540), .ZN(U2971) );
  INV_X1 U6691 ( .A(n5543), .ZN(n5545) );
  NAND2_X1 U6692 ( .A1(n5545), .A2(n5544), .ZN(n5546) );
  XNOR2_X1 U6693 ( .A(n5542), .B(n5546), .ZN(n5722) );
  INV_X1 U6694 ( .A(n5547), .ZN(n5981) );
  AOI22_X1 U6695 ( .A1(n6108), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6187), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5548) );
  OAI21_X1 U6696 ( .B1(n6117), .B2(n5549), .A(n5548), .ZN(n5550) );
  AOI21_X1 U6697 ( .B1(n5981), .B2(n6113), .A(n5550), .ZN(n5551) );
  OAI21_X1 U6698 ( .B1(n5722), .B2(n6092), .A(n5551), .ZN(U2972) );
  INV_X1 U6699 ( .A(n5552), .ZN(n5556) );
  INV_X1 U6700 ( .A(n5585), .ZN(n5574) );
  NOR3_X1 U6701 ( .A1(n5574), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5553), 
        .ZN(n5554) );
  AOI211_X1 U6702 ( .C1(n5556), .C2(n6189), .A(n5555), .B(n5554), .ZN(n5560)
         );
  INV_X1 U6703 ( .A(n5557), .ZN(n5558) );
  NAND2_X1 U6704 ( .A1(n5558), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5559) );
  OAI211_X1 U6705 ( .C1(n5561), .C2(n5721), .A(n5560), .B(n5559), .ZN(U2988)
         );
  NOR3_X1 U6706 ( .A1(n5574), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5563), 
        .ZN(n5564) );
  AOI211_X1 U6707 ( .C1(n5566), .C2(n6189), .A(n5565), .B(n5564), .ZN(n5569)
         );
  NAND2_X1 U6708 ( .A1(n5567), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5568) );
  OAI211_X1 U6709 ( .C1(n5432), .C2(n5721), .A(n5569), .B(n5568), .ZN(U2989)
         );
  INV_X1 U6710 ( .A(n5583), .ZN(n5577) );
  OAI21_X1 U6711 ( .B1(n5571), .B2(n6119), .A(n5570), .ZN(n5576) );
  NOR3_X1 U6712 ( .A1(n5574), .A2(n5573), .A3(n5572), .ZN(n5575) );
  AOI211_X1 U6713 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n5577), .A(n5576), .B(n5575), .ZN(n5578) );
  OAI21_X1 U6714 ( .B1(n5579), .B2(n5721), .A(n5578), .ZN(U2990) );
  NAND2_X1 U6715 ( .A1(n5580), .A2(n6189), .ZN(n5582) );
  OAI211_X1 U6716 ( .C1(n5583), .C2(n6797), .A(n5582), .B(n5581), .ZN(n5584)
         );
  AOI21_X1 U6717 ( .B1(n5585), .B2(n6797), .A(n5584), .ZN(n5586) );
  OAI21_X1 U6718 ( .B1(n5587), .B2(n5721), .A(n5586), .ZN(U2991) );
  OAI21_X1 U6719 ( .B1(n5589), .B2(n6119), .A(n5588), .ZN(n5594) );
  INV_X1 U6720 ( .A(n5590), .ZN(n5591) );
  AOI211_X1 U6721 ( .C1(n6887), .C2(n5592), .A(n5591), .B(n5599), .ZN(n5593)
         );
  AOI211_X1 U6722 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n5606), .A(n5594), .B(n5593), .ZN(n5595) );
  OAI21_X1 U6723 ( .B1(n5596), .B2(n5721), .A(n5595), .ZN(U2992) );
  OAI21_X1 U6724 ( .B1(n5598), .B2(n6119), .A(n5597), .ZN(n5601) );
  NOR2_X1 U6725 ( .A1(n5599), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5600)
         );
  AOI211_X1 U6726 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5606), .A(n5601), .B(n5600), .ZN(n5602) );
  OAI21_X1 U6727 ( .B1(n5603), .B2(n5721), .A(n5602), .ZN(U2993) );
  INV_X1 U6728 ( .A(n5604), .ZN(n5665) );
  NAND2_X1 U6729 ( .A1(n5665), .A2(n5605), .ZN(n5616) );
  INV_X1 U6730 ( .A(n5606), .ZN(n5607) );
  AOI211_X1 U6731 ( .C1(n5609), .C2(n5616), .A(n5608), .B(n5607), .ZN(n5610)
         );
  AOI211_X1 U6732 ( .C1(n6189), .C2(n5612), .A(n5611), .B(n5610), .ZN(n5613)
         );
  OAI21_X1 U6733 ( .B1(n5614), .B2(n5721), .A(n5613), .ZN(U2994) );
  OAI21_X1 U6734 ( .B1(n5739), .B2(n6119), .A(n5615), .ZN(n5618) );
  NOR2_X1 U6735 ( .A1(n5616), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5617)
         );
  AOI211_X1 U6736 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5619), .A(n5618), .B(n5617), .ZN(n5620) );
  OAI21_X1 U6737 ( .B1(n5621), .B2(n5721), .A(n5620), .ZN(U2995) );
  INV_X1 U6738 ( .A(n5622), .ZN(n5636) );
  OAI21_X1 U6739 ( .B1(n5749), .B2(n6119), .A(n5623), .ZN(n5629) );
  NAND2_X1 U6740 ( .A1(n5689), .A2(n5624), .ZN(n5639) );
  INV_X1 U6741 ( .A(n5625), .ZN(n5626) );
  NOR3_X1 U6742 ( .A1(n5639), .A2(n5627), .A3(n5626), .ZN(n5628) );
  AOI211_X1 U6743 ( .C1(n5636), .C2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5629), .B(n5628), .ZN(n5630) );
  OAI21_X1 U6744 ( .B1(n5631), .B2(n5721), .A(n5630), .ZN(U2996) );
  NAND2_X1 U6745 ( .A1(n5632), .A2(n4243), .ZN(n5638) );
  OAI21_X1 U6746 ( .B1(n5634), .B2(n6119), .A(n5633), .ZN(n5635) );
  AOI21_X1 U6747 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5636), .A(n5635), 
        .ZN(n5637) );
  OAI211_X1 U6748 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5639), .A(n5638), .B(n5637), .ZN(U2997) );
  XNOR2_X1 U6749 ( .A(n5664), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5656)
         );
  MUX2_X1 U6750 ( .A(n5642), .B(n5641), .S(n5640), .Z(n5644) );
  XNOR2_X1 U6751 ( .A(n5644), .B(n5643), .ZN(n5785) );
  OAI21_X1 U6752 ( .B1(n5785), .B2(n6119), .A(n5645), .ZN(n5655) );
  INV_X1 U6753 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5688) );
  NOR2_X1 U6754 ( .A1(n5694), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5652)
         );
  OAI21_X1 U6755 ( .B1(n5647), .B2(n5688), .A(n5646), .ZN(n5650) );
  NAND2_X1 U6756 ( .A1(n5653), .A2(n5648), .ZN(n5649) );
  NAND3_X1 U6757 ( .A1(n5651), .A2(n5650), .A3(n5649), .ZN(n5668) );
  AOI211_X1 U6758 ( .C1(n5688), .C2(n5653), .A(n5652), .B(n5668), .ZN(n5662)
         );
  NOR2_X1 U6759 ( .A1(n5662), .A2(n6933), .ZN(n5654) );
  AOI211_X1 U6760 ( .C1(n5656), .C2(n5665), .A(n5655), .B(n5654), .ZN(n5657)
         );
  OAI21_X1 U6761 ( .B1(n5658), .B2(n5721), .A(n5657), .ZN(U2998) );
  NAND2_X1 U6762 ( .A1(n5659), .A2(n6189), .ZN(n5660) );
  OAI211_X1 U6763 ( .C1(n5662), .C2(n5664), .A(n5661), .B(n5660), .ZN(n5663)
         );
  AOI21_X1 U6764 ( .B1(n5665), .B2(n5664), .A(n5663), .ZN(n5666) );
  OAI21_X1 U6765 ( .B1(n5667), .B2(n5721), .A(n5666), .ZN(U2999) );
  INV_X1 U6766 ( .A(n5668), .ZN(n5686) );
  OAI21_X1 U6767 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n6123), .A(n5686), 
        .ZN(n5674) );
  OAI21_X1 U6768 ( .B1(n5671), .B2(n5670), .A(n5669), .ZN(n5871) );
  OAI21_X1 U6769 ( .B1(n5871), .B2(n6119), .A(n5672), .ZN(n5673) );
  AOI21_X1 U6770 ( .B1(n5674), .B2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n5673), 
        .ZN(n5677) );
  NAND3_X1 U6771 ( .A1(n5689), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5675), .ZN(n5676) );
  OAI211_X1 U6772 ( .C1(n5678), .C2(n5721), .A(n5677), .B(n5676), .ZN(U3000)
         );
  INV_X1 U6773 ( .A(n5679), .ZN(n5680) );
  NOR2_X1 U6774 ( .A1(n5681), .A2(n5680), .ZN(n5682) );
  XNOR2_X1 U6775 ( .A(n5682), .B(n5688), .ZN(n5803) );
  XOR2_X1 U6776 ( .A(n5684), .B(n5683), .Z(n5976) );
  AOI22_X1 U6777 ( .A1(n5976), .A2(n6189), .B1(n6187), .B2(
        REIP_REG_17__SCAN_IN), .ZN(n5685) );
  OAI21_X1 U6778 ( .B1(n5686), .B2(n5688), .A(n5685), .ZN(n5687) );
  AOI21_X1 U6779 ( .B1(n5689), .B2(n5688), .A(n5687), .ZN(n5690) );
  OAI21_X1 U6780 ( .B1(n5803), .B2(n5721), .A(n5690), .ZN(U3001) );
  AOI21_X1 U6781 ( .B1(n5692), .B2(n5691), .A(n5823), .ZN(n5700) );
  OAI21_X1 U6782 ( .B1(n5694), .B2(n5693), .A(n6125), .ZN(n5819) );
  NAND2_X1 U6783 ( .A1(n5819), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5696) );
  OAI211_X1 U6784 ( .C1(n6119), .C2(n5697), .A(n5696), .B(n5695), .ZN(n5698)
         );
  AOI21_X1 U6785 ( .B1(n5700), .B2(n5699), .A(n5698), .ZN(n5701) );
  OAI21_X1 U6786 ( .B1(n5702), .B2(n5721), .A(n5701), .ZN(U3002) );
  NAND2_X1 U6787 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5703), .ZN(n5705)
         );
  INV_X1 U6788 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6899) );
  OR3_X1 U6789 ( .A1(n6130), .A2(n6899), .A3(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5704) );
  AOI221_X1 U6790 ( .B1(n5826), .B2(n5706), .C1(n5705), .C2(n5706), .A(n5704), 
        .ZN(n5824) );
  NAND2_X1 U6791 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5827) );
  AOI22_X1 U6792 ( .A1(n5829), .A2(n5710), .B1(n5707), .B2(n5827), .ZN(n5708)
         );
  NAND2_X1 U6793 ( .A1(n6125), .A2(n5708), .ZN(n5831) );
  OAI21_X1 U6794 ( .B1(n5824), .B2(n5831), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5709) );
  INV_X1 U6795 ( .A(n5709), .ZN(n5719) );
  NOR3_X1 U6796 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5711), .A3(n5710), 
        .ZN(n5718) );
  INV_X1 U6797 ( .A(n5712), .ZN(n5825) );
  NAND2_X1 U6798 ( .A1(n3198), .A2(n5825), .ZN(n5714) );
  NAND2_X1 U6799 ( .A1(n5714), .A2(n5713), .ZN(n5716) );
  NAND2_X1 U6800 ( .A1(n5716), .A2(n5715), .ZN(n5978) );
  OAI22_X1 U6801 ( .A1(n5978), .A2(n6119), .B1(n6666), .B2(n6177), .ZN(n5717)
         );
  NOR3_X1 U6802 ( .A1(n5719), .A2(n5718), .A3(n5717), .ZN(n5720) );
  OAI21_X1 U6803 ( .B1(n5722), .B2(n5721), .A(n5720), .ZN(U3004) );
  NAND2_X1 U6804 ( .A1(n5726), .A2(n6506), .ZN(n6472) );
  NOR2_X1 U6805 ( .A1(n5723), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5724) );
  OAI22_X1 U6806 ( .A1(n6472), .A2(n5724), .B1(n4510), .B2(n5728), .ZN(n5725)
         );
  MUX2_X1 U6807 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5725), .S(n6201), 
        .Z(U3464) );
  XNOR2_X1 U6808 ( .A(n5727), .B(n5726), .ZN(n5729) );
  OAI22_X1 U6809 ( .A1(n5729), .A2(n6519), .B1(n4536), .B2(n5728), .ZN(n5730)
         );
  MUX2_X1 U6810 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5730), .S(n6201), 
        .Z(U3463) );
  INV_X1 U6811 ( .A(n6574), .ZN(n5733) );
  OAI22_X1 U6812 ( .A1(n5733), .A2(n5732), .B1(n5731), .B2(n6610), .ZN(n5734)
         );
  MUX2_X1 U6813 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5734), .S(n5839), 
        .Z(U3456) );
  AND2_X1 U6814 ( .A1(n6040), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI21_X1 U6815 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n5736), .A(n5735), .ZN(
        n5737) );
  NAND2_X1 U6816 ( .A1(n5846), .A2(n5737), .ZN(U2788) );
  AOI22_X1 U6817 ( .A1(PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n5960), .B1(n5738), 
        .B2(n5939), .ZN(n5745) );
  OAI22_X1 U6818 ( .A1(n5740), .A2(n5776), .B1(n5739), .B2(n5958), .ZN(n5741)
         );
  OAI211_X1 U6819 ( .C1(n5746), .C2(n6939), .A(n5745), .B(n5744), .ZN(U2804)
         );
  AOI22_X1 U6820 ( .A1(EBX_REG_22__SCAN_IN), .A2(n5968), .B1(
        REIP_REG_22__SCAN_IN), .B2(n5766), .ZN(n5756) );
  INV_X1 U6821 ( .A(n5747), .ZN(n5748) );
  AOI22_X1 U6822 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n5960), .B1(n5748), 
        .B2(n5939), .ZN(n5755) );
  INV_X1 U6823 ( .A(n5749), .ZN(n5750) );
  AOI22_X1 U6824 ( .A1(n5789), .A2(n5929), .B1(n5904), .B2(n5750), .ZN(n5754)
         );
  INV_X1 U6825 ( .A(n5751), .ZN(n5757) );
  OAI211_X1 U6826 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5757), .B(n5752), .ZN(n5753) );
  NAND4_X1 U6827 ( .A1(n5756), .A2(n5755), .A3(n5754), .A4(n5753), .ZN(U2805)
         );
  INV_X1 U6828 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6675) );
  AOI22_X1 U6829 ( .A1(EBX_REG_21__SCAN_IN), .A2(n5968), .B1(n5757), .B2(n6675), .ZN(n5764) );
  AOI22_X1 U6830 ( .A1(n5758), .A2(n5939), .B1(REIP_REG_21__SCAN_IN), .B2(
        n5766), .ZN(n5763) );
  INV_X1 U6831 ( .A(n5759), .ZN(n5792) );
  AOI22_X1 U6832 ( .A1(n5792), .A2(n5929), .B1(n5904), .B2(n5760), .ZN(n5762)
         );
  NAND2_X1 U6833 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n5960), .ZN(n5761)
         );
  NAND4_X1 U6834 ( .A1(n5764), .A2(n5763), .A3(n5762), .A4(n5761), .ZN(U2806)
         );
  AOI22_X1 U6835 ( .A1(EBX_REG_20__SCAN_IN), .A2(n5968), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n5960), .ZN(n5772) );
  OAI22_X1 U6836 ( .A1(n5795), .A2(n5776), .B1(n5958), .B2(n5785), .ZN(n5765)
         );
  INV_X1 U6837 ( .A(n5765), .ZN(n5771) );
  OAI21_X1 U6838 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5767), .A(n5766), .ZN(n5770) );
  NAND2_X1 U6839 ( .A1(n5768), .A2(n5939), .ZN(n5769) );
  NAND4_X1 U6840 ( .A1(n5772), .A2(n5771), .A3(n5770), .A4(n5769), .ZN(U2807)
         );
  AOI22_X1 U6841 ( .A1(EBX_REG_19__SCAN_IN), .A2(n5968), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n5960), .ZN(n5784) );
  NAND2_X1 U6842 ( .A1(n5963), .A2(n5868), .ZN(n5774) );
  AND2_X1 U6843 ( .A1(n5774), .A2(n5773), .ZN(n5866) );
  NAND2_X1 U6844 ( .A1(n5963), .A2(n6671), .ZN(n5867) );
  INV_X1 U6845 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6948) );
  AOI21_X1 U6846 ( .B1(n5866), .B2(n5867), .A(n6948), .ZN(n5779) );
  OAI22_X1 U6847 ( .A1(n5777), .A2(n5776), .B1(n5958), .B2(n5775), .ZN(n5778)
         );
  AOI211_X1 U6848 ( .C1(n5939), .C2(n5780), .A(n5779), .B(n5778), .ZN(n5783)
         );
  NAND3_X1 U6849 ( .A1(n5963), .A2(n6948), .A3(n5781), .ZN(n5782) );
  NAND4_X1 U6850 ( .A1(n5784), .A2(n5783), .A3(n5924), .A4(n5782), .ZN(U2808)
         );
  OAI22_X1 U6851 ( .A1(n5795), .A2(n5389), .B1(n5785), .B2(n5984), .ZN(n5786)
         );
  INV_X1 U6852 ( .A(n5786), .ZN(n5787) );
  OAI21_X1 U6853 ( .B1(n5989), .B2(n5788), .A(n5787), .ZN(U2839) );
  AOI22_X1 U6854 ( .A1(n5789), .A2(n6006), .B1(n5997), .B2(DATAI_22_), .ZN(
        n5791) );
  AOI22_X1 U6855 ( .A1(n6000), .A2(DATAI_6_), .B1(n5999), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U6856 ( .A1(n5791), .A2(n5790), .ZN(U2869) );
  AOI22_X1 U6857 ( .A1(n5792), .A2(n6006), .B1(n5997), .B2(DATAI_21_), .ZN(
        n5794) );
  AOI22_X1 U6858 ( .A1(n6000), .A2(DATAI_5_), .B1(n5999), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5793) );
  NAND2_X1 U6859 ( .A1(n5794), .A2(n5793), .ZN(U2870) );
  INV_X1 U6860 ( .A(n5795), .ZN(n5796) );
  AOI22_X1 U6861 ( .A1(n5796), .A2(n6006), .B1(n5997), .B2(DATAI_20_), .ZN(
        n5798) );
  AOI22_X1 U6862 ( .A1(n6000), .A2(DATAI_4_), .B1(n5999), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5797) );
  NAND2_X1 U6863 ( .A1(n5798), .A2(n5797), .ZN(U2871) );
  AOI22_X1 U6864 ( .A1(n6187), .A2(REIP_REG_17__SCAN_IN), .B1(n6108), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5802) );
  XOR2_X1 U6865 ( .A(n5800), .B(n5799), .Z(n5993) );
  AOI22_X1 U6866 ( .A1(n5993), .A2(n6113), .B1(n6088), .B2(n5879), .ZN(n5801)
         );
  OAI211_X1 U6867 ( .C1(n5803), .C2(n6092), .A(n5802), .B(n5801), .ZN(U2969)
         );
  AOI22_X1 U6868 ( .A1(n6187), .A2(REIP_REG_13__SCAN_IN), .B1(n6108), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5815) );
  XNOR2_X1 U6869 ( .A(n5805), .B(n5804), .ZN(n5832) );
  AND2_X1 U6870 ( .A1(n5806), .A2(n5024), .ZN(n5809) );
  INV_X1 U6871 ( .A(n5807), .ZN(n5808) );
  NOR2_X1 U6872 ( .A1(n5809), .A2(n5808), .ZN(n5811) );
  NAND2_X1 U6873 ( .A1(n5811), .A2(n5810), .ZN(n5812) );
  AND2_X1 U6874 ( .A1(n5813), .A2(n5812), .ZN(n6003) );
  AOI22_X1 U6875 ( .A1(n5832), .A2(n4502), .B1(n6113), .B2(n6003), .ZN(n5814)
         );
  OAI211_X1 U6876 ( .C1(n6117), .C2(n5902), .A(n5815), .B(n5814), .ZN(U2973)
         );
  INV_X1 U6877 ( .A(n5816), .ZN(n5817) );
  AOI21_X1 U6878 ( .B1(n5818), .B2(n6189), .A(n5817), .ZN(n5822) );
  AOI22_X1 U6879 ( .A1(n5820), .A2(n4243), .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n5819), .ZN(n5821) );
  OAI211_X1 U6880 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n5823), .A(n5822), .B(n5821), .ZN(U3003) );
  INV_X1 U6881 ( .A(n5824), .ZN(n5836) );
  XNOR2_X1 U6882 ( .A(n3198), .B(n5825), .ZN(n5985) );
  INV_X1 U6883 ( .A(n5985), .ZN(n5830) );
  NOR3_X1 U6884 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5827), .A3(n5826), 
        .ZN(n5828) );
  AOI22_X1 U6885 ( .A1(n5830), .A2(n6189), .B1(n5829), .B2(n5828), .ZN(n5835)
         );
  AOI22_X1 U6886 ( .A1(n5832), .A2(n4243), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5831), .ZN(n5834) );
  NAND2_X1 U6887 ( .A1(n6187), .A2(REIP_REG_13__SCAN_IN), .ZN(n5833) );
  NAND4_X1 U6888 ( .A1(n5836), .A2(n5835), .A3(n5834), .A4(n5833), .ZN(U3005)
         );
  INV_X1 U6889 ( .A(n5837), .ZN(n5838) );
  NAND2_X1 U6890 ( .A1(n5838), .A2(n4054), .ZN(n5841) );
  OAI22_X1 U6891 ( .A1(n5842), .A2(n5841), .B1(n5840), .B2(n5839), .ZN(U3455)
         );
  INV_X1 U6892 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6645) );
  AOI21_X1 U6893 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6645), .A(n6636), .ZN(n5848) );
  INV_X1 U6894 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5843) );
  AOI21_X1 U6895 ( .B1(n5848), .B2(n5843), .A(n6678), .ZN(U2789) );
  OAI21_X1 U6896 ( .B1(n5844), .B2(n6614), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5845) );
  OAI21_X1 U6897 ( .B1(n5846), .B2(n6609), .A(n5845), .ZN(U2790) );
  INV_X2 U6898 ( .A(n6678), .ZN(n6719) );
  NOR2_X1 U6899 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n5849) );
  OAI21_X1 U6900 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5849), .A(n6719), .ZN(n5847)
         );
  OAI21_X1 U6901 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6719), .A(n5847), .ZN(
        U2791) );
  NOR2_X2 U6902 ( .A1(n6678), .A2(n5848), .ZN(n6696) );
  OAI21_X1 U6903 ( .B1(BS16_N), .B2(n5849), .A(n6696), .ZN(n6695) );
  OAI21_X1 U6904 ( .B1(n6696), .B2(n6832), .A(n6695), .ZN(U2792) );
  INV_X1 U6905 ( .A(n5850), .ZN(n5851) );
  OAI21_X1 U6906 ( .B1(n5851), .B2(n7032), .A(n6092), .ZN(U2793) );
  NOR4_X1 U6907 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_31__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_20__SCAN_IN), .ZN(n5861) );
  AOI211_X1 U6908 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_16__SCAN_IN), .B(
        DATAWIDTH_REG_12__SCAN_IN), .ZN(n5860) );
  NOR4_X1 U6909 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_5__SCAN_IN), .ZN(n5852) );
  INV_X1 U6910 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n7010) );
  INV_X1 U6911 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6990) );
  NAND3_X1 U6912 ( .A1(n5852), .A2(n7010), .A3(n6990), .ZN(n5858) );
  NOR4_X1 U6913 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_17__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n5856) );
  NOR4_X1 U6914 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_9__SCAN_IN), .A4(DATAWIDTH_REG_10__SCAN_IN), .ZN(
        n5855) );
  NOR4_X1 U6915 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(
        DATAWIDTH_REG_26__SCAN_IN), .A3(DATAWIDTH_REG_27__SCAN_IN), .A4(
        DATAWIDTH_REG_28__SCAN_IN), .ZN(n5854) );
  NOR4_X1 U6916 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_24__SCAN_IN), .ZN(n5853) );
  NAND4_X1 U6917 ( .A1(n5856), .A2(n5855), .A3(n5854), .A4(n5853), .ZN(n5857)
         );
  NOR4_X1 U6918 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(
        DATAWIDTH_REG_11__SCAN_IN), .A3(n5858), .A4(n5857), .ZN(n5859) );
  NAND3_X1 U6919 ( .A1(n5861), .A2(n5860), .A3(n5859), .ZN(n6705) );
  NOR2_X1 U6920 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6705), .ZN(n6706) );
  INV_X1 U6921 ( .A(n6705), .ZN(n5862) );
  NOR2_X1 U6922 ( .A1(n5862), .A2(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5863) );
  INV_X1 U6923 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6699) );
  INV_X1 U6924 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6829) );
  INV_X1 U6925 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6700) );
  NAND4_X1 U6926 ( .A1(n5862), .A2(n6699), .A3(n6829), .A4(n6700), .ZN(n5864)
         );
  OAI21_X1 U6927 ( .B1(n6706), .B2(n5863), .A(n5864), .ZN(U2794) );
  AOI22_X1 U6928 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(n6705), .B1(n6706), 
        .B2(n6699), .ZN(n5865) );
  NAND2_X1 U6929 ( .A1(n5865), .A2(n5864), .ZN(U2795) );
  INV_X1 U6930 ( .A(n5866), .ZN(n5878) );
  AOI22_X1 U6931 ( .A1(EBX_REG_18__SCAN_IN), .A2(n5968), .B1(
        REIP_REG_18__SCAN_IN), .B2(n5878), .ZN(n5874) );
  OAI22_X1 U6932 ( .A1(n5869), .A2(n5973), .B1(n5868), .B2(n5867), .ZN(n5870)
         );
  AOI21_X1 U6933 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n5960), .A(n5870), 
        .ZN(n5873) );
  INV_X1 U6934 ( .A(n5871), .ZN(n5974) );
  AOI22_X1 U6935 ( .A1(n5990), .A2(n5929), .B1(n5904), .B2(n5974), .ZN(n5872)
         );
  NAND4_X1 U6936 ( .A1(n5874), .A2(n5873), .A3(n5872), .A4(n5924), .ZN(U2809)
         );
  NAND2_X1 U6937 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n5876) );
  INV_X1 U6938 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6669) );
  OAI21_X1 U6939 ( .B1(n5876), .B2(n5875), .A(n6669), .ZN(n5877) );
  AOI22_X1 U6940 ( .A1(n5879), .A2(n5939), .B1(n5878), .B2(n5877), .ZN(n5882)
         );
  AOI22_X1 U6941 ( .A1(EBX_REG_17__SCAN_IN), .A2(n5968), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n5960), .ZN(n5881) );
  AOI22_X1 U6942 ( .A1(n5993), .A2(n5929), .B1(n5904), .B2(n5976), .ZN(n5880)
         );
  NAND4_X1 U6943 ( .A1(n5882), .A2(n5881), .A3(n5880), .A4(n5924), .ZN(U2810)
         );
  INV_X1 U6944 ( .A(n5883), .ZN(n5885) );
  AOI22_X1 U6945 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5886), .B1(n5885), .B2(
        n5884), .ZN(n5892) );
  OR2_X1 U6946 ( .A1(n5978), .A2(n5958), .ZN(n5888) );
  AOI22_X1 U6947 ( .A1(n5968), .A2(EBX_REG_14__SCAN_IN), .B1(n5960), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5887) );
  AND2_X1 U6948 ( .A1(n5888), .A2(n5887), .ZN(n5891) );
  AOI22_X1 U6949 ( .A1(n5981), .A2(n5929), .B1(n5939), .B2(n5889), .ZN(n5890)
         );
  NAND4_X1 U6950 ( .A1(n5892), .A2(n5891), .A3(n5890), .A4(n5924), .ZN(U2813)
         );
  INV_X1 U6951 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5895) );
  INV_X1 U6952 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6664) );
  NAND3_X1 U6953 ( .A1(n5963), .A2(n6664), .A3(n5893), .ZN(n5894) );
  OAI211_X1 U6954 ( .C1(n5895), .C2(n5934), .A(n5894), .B(n5924), .ZN(n5896)
         );
  AOI21_X1 U6955 ( .B1(EBX_REG_13__SCAN_IN), .B2(n5968), .A(n5896), .ZN(n5897)
         );
  OAI21_X1 U6956 ( .B1(n5985), .B2(n5958), .A(n5897), .ZN(n5898) );
  AOI21_X1 U6957 ( .B1(n6003), .B2(n5929), .A(n5898), .ZN(n5901) );
  OAI21_X1 U6958 ( .B1(n5899), .B2(n5903), .A(REIP_REG_13__SCAN_IN), .ZN(n5900) );
  OAI211_X1 U6959 ( .C1(n5973), .C2(n5902), .A(n5901), .B(n5900), .ZN(U2814)
         );
  AOI22_X1 U6960 ( .A1(n5905), .A2(n5904), .B1(REIP_REG_11__SCAN_IN), .B2(
        n5903), .ZN(n5913) );
  INV_X1 U6961 ( .A(n5906), .ZN(n5908) );
  OAI22_X1 U6962 ( .A1(n5909), .A2(n5934), .B1(n5908), .B2(n5907), .ZN(n5910)
         );
  AOI21_X1 U6963 ( .B1(EBX_REG_11__SCAN_IN), .B2(n5968), .A(n5910), .ZN(n5912)
         );
  AOI22_X1 U6964 ( .A1(n6089), .A2(n5929), .B1(n5939), .B2(n6087), .ZN(n5911)
         );
  NAND4_X1 U6965 ( .A1(n5913), .A2(n5912), .A3(n5911), .A4(n5924), .ZN(U2816)
         );
  AOI22_X1 U6966 ( .A1(EBX_REG_9__SCAN_IN), .A2(n5968), .B1(
        REIP_REG_9__SCAN_IN), .B2(n5914), .ZN(n5921) );
  OAI21_X1 U6967 ( .B1(n5915), .B2(n5958), .A(n5924), .ZN(n5916) );
  AOI211_X1 U6968 ( .C1(n5960), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n5917), 
        .B(n5916), .ZN(n5920) );
  AOI22_X1 U6969 ( .A1(n6007), .A2(n5929), .B1(n5939), .B2(n5918), .ZN(n5919)
         );
  NAND3_X1 U6970 ( .A1(n5921), .A2(n5920), .A3(n5919), .ZN(U2818) );
  AND2_X1 U6971 ( .A1(n5968), .A2(EBX_REG_6__SCAN_IN), .ZN(n5927) );
  INV_X1 U6972 ( .A(REIP_REG_6__SCAN_IN), .ZN(n7017) );
  AOI22_X1 U6973 ( .A1(n5944), .A2(REIP_REG_6__SCAN_IN), .B1(n7017), .B2(n5922), .ZN(n5926) );
  NAND2_X1 U6974 ( .A1(n5960), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5923)
         );
  OAI211_X1 U6975 ( .C1(n5958), .C2(n6161), .A(n5924), .B(n5923), .ZN(n5925)
         );
  OR3_X1 U6976 ( .A1(n5927), .A2(n5926), .A3(n5925), .ZN(n5928) );
  AOI21_X1 U6977 ( .B1(n6096), .B2(n5929), .A(n5928), .ZN(n5930) );
  OAI21_X1 U6978 ( .B1(n6099), .B2(n5973), .A(n5930), .ZN(U2821) );
  NOR3_X1 U6979 ( .A1(n5932), .A2(n6647), .A3(n5931), .ZN(n5954) );
  AOI21_X1 U6980 ( .B1(REIP_REG_4__SCAN_IN), .B2(n5954), .A(
        REIP_REG_5__SCAN_IN), .ZN(n5945) );
  INV_X1 U6981 ( .A(n5933), .ZN(n5936) );
  INV_X1 U6982 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5935) );
  OAI22_X1 U6983 ( .A1(n5958), .A2(n5936), .B1(n5935), .B2(n5934), .ZN(n5937)
         );
  AOI211_X1 U6984 ( .C1(EBX_REG_5__SCAN_IN), .C2(n5968), .A(n5947), .B(n5937), 
        .ZN(n5943) );
  INV_X1 U6985 ( .A(n5938), .ZN(n5940) );
  AOI22_X1 U6986 ( .A1(n5941), .A2(n5969), .B1(n5940), .B2(n5939), .ZN(n5942)
         );
  OAI211_X1 U6987 ( .C1(n5945), .C2(n5944), .A(n5943), .B(n5942), .ZN(U2822)
         );
  INV_X1 U6988 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6986) );
  INV_X1 U6989 ( .A(n6168), .ZN(n5951) );
  AND2_X1 U6990 ( .A1(n5960), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5946)
         );
  AOI211_X1 U6991 ( .C1(n5948), .C2(n5962), .A(n5947), .B(n5946), .ZN(n5950)
         );
  NAND2_X1 U6992 ( .A1(n5968), .A2(EBX_REG_4__SCAN_IN), .ZN(n5949) );
  OAI211_X1 U6993 ( .C1(n5951), .C2(n5958), .A(n5950), .B(n5949), .ZN(n5952)
         );
  AOI221_X1 U6994 ( .B1(n5954), .B2(n6986), .C1(n5953), .C2(
        REIP_REG_4__SCAN_IN), .A(n5952), .ZN(n5956) );
  NAND2_X1 U6995 ( .A1(n6104), .A2(n5969), .ZN(n5955) );
  OAI211_X1 U6996 ( .C1(n5973), .C2(n6107), .A(n5956), .B(n5955), .ZN(U2823)
         );
  OR2_X1 U6997 ( .A1(n5958), .A2(n5957), .ZN(n5967) );
  AOI22_X1 U6998 ( .A1(n5960), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n5959), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5966) );
  NAND2_X1 U6999 ( .A1(n5962), .A2(n5961), .ZN(n5965) );
  NAND2_X1 U7000 ( .A1(n5963), .A2(n6647), .ZN(n5964) );
  AND4_X1 U7001 ( .A1(n5967), .A2(n5966), .A3(n5965), .A4(n5964), .ZN(n5972)
         );
  AOI22_X1 U7002 ( .A1(n5970), .A2(n5969), .B1(EBX_REG_1__SCAN_IN), .B2(n5968), 
        .ZN(n5971) );
  OAI211_X1 U7003 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n5973), .A(n5972), 
        .B(n5971), .ZN(U2826) );
  AOI22_X1 U7004 ( .A1(n5990), .A2(n5987), .B1(n5974), .B2(n5980), .ZN(n5975)
         );
  OAI21_X1 U7005 ( .B1(n5989), .B2(n5383), .A(n5975), .ZN(U2841) );
  INV_X1 U7006 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6982) );
  AOI22_X1 U7007 ( .A1(n5993), .A2(n5987), .B1(n5980), .B2(n5976), .ZN(n5977)
         );
  OAI21_X1 U7008 ( .B1(n5989), .B2(n6982), .A(n5977), .ZN(U2842) );
  INV_X1 U7009 ( .A(n5978), .ZN(n5979) );
  AOI22_X1 U7010 ( .A1(n5981), .A2(n5987), .B1(n5980), .B2(n5979), .ZN(n5982)
         );
  OAI21_X1 U7011 ( .B1(n5989), .B2(n5983), .A(n5982), .ZN(U2845) );
  INV_X1 U7012 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6820) );
  NOR2_X1 U7013 ( .A1(n5985), .A2(n5984), .ZN(n5986) );
  AOI21_X1 U7014 ( .B1(n6003), .B2(n5987), .A(n5986), .ZN(n5988) );
  OAI21_X1 U7015 ( .B1(n5989), .B2(n6820), .A(n5988), .ZN(U2846) );
  AOI22_X1 U7016 ( .A1(n5990), .A2(n6006), .B1(n5997), .B2(DATAI_18_), .ZN(
        n5992) );
  AOI22_X1 U7017 ( .A1(n6000), .A2(DATAI_2_), .B1(n5999), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U7018 ( .A1(n5992), .A2(n5991), .ZN(U2873) );
  AOI22_X1 U7019 ( .A1(n5993), .A2(n6006), .B1(n5997), .B2(DATAI_17_), .ZN(
        n5995) );
  AOI22_X1 U7020 ( .A1(n6000), .A2(DATAI_1_), .B1(n5999), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5994) );
  NAND2_X1 U7021 ( .A1(n5995), .A2(n5994), .ZN(U2874) );
  INV_X1 U7022 ( .A(n5996), .ZN(n5998) );
  AOI22_X1 U7023 ( .A1(n5998), .A2(n6006), .B1(n5997), .B2(DATAI_16_), .ZN(
        n6002) );
  AOI22_X1 U7024 ( .A1(n6000), .A2(DATAI_0_), .B1(n5999), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7025 ( .A1(n6002), .A2(n6001), .ZN(U2875) );
  INV_X1 U7026 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6870) );
  AOI22_X1 U7027 ( .A1(n6003), .A2(n6006), .B1(DATAI_13_), .B2(n6005), .ZN(
        n6004) );
  OAI21_X1 U7028 ( .B1(n6870), .B2(n6010), .A(n6004), .ZN(U2878) );
  INV_X1 U7029 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6971) );
  AOI22_X1 U7030 ( .A1(n6007), .A2(n6006), .B1(DATAI_9_), .B2(n6005), .ZN(
        n6008) );
  OAI21_X1 U7031 ( .B1(n6971), .B2(n6010), .A(n6008), .ZN(U2882) );
  INV_X1 U7032 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6044) );
  OAI222_X1 U7033 ( .A1(n6012), .A2(n6011), .B1(n6010), .B2(n6044), .C1(n6009), 
        .C2(n6065), .ZN(U2891) );
  AOI22_X1 U7034 ( .A1(n6040), .A2(DATAO_REG_26__SCAN_IN), .B1(n6015), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6013) );
  OAI21_X1 U7035 ( .B1(n6917), .B2(n6708), .A(n6013), .ZN(U2897) );
  INV_X1 U7036 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n6998) );
  AOI22_X1 U7037 ( .A1(n6015), .A2(EAX_REG_22__SCAN_IN), .B1(n6041), .B2(
        UWORD_REG_6__SCAN_IN), .ZN(n6014) );
  OAI21_X1 U7038 ( .B1(n6998), .B2(n6023), .A(n6014), .ZN(U2901) );
  INV_X1 U7039 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n6941) );
  AOI22_X1 U7040 ( .A1(n6015), .A2(EAX_REG_16__SCAN_IN), .B1(n6041), .B2(
        UWORD_REG_0__SCAN_IN), .ZN(n6016) );
  OAI21_X1 U7041 ( .B1(n6941), .B2(n6023), .A(n6016), .ZN(U2907) );
  AOI22_X1 U7042 ( .A1(EAX_REG_15__SCAN_IN), .A2(n6030), .B1(n6040), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6017) );
  OAI21_X1 U7043 ( .B1(n4579), .B2(n6708), .A(n6017), .ZN(U2908) );
  INV_X1 U7044 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6086) );
  AOI22_X1 U7045 ( .A1(DATAO_REG_14__SCAN_IN), .A2(n6040), .B1(n6041), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n6018) );
  OAI21_X1 U7046 ( .B1(n6086), .B2(n6043), .A(n6018), .ZN(U2909) );
  AOI22_X1 U7047 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n6041), .B1(n6040), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6019) );
  OAI21_X1 U7048 ( .B1(n6870), .B2(n6043), .A(n6019), .ZN(U2910) );
  AOI22_X1 U7049 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6030), .B1(n6040), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6020) );
  OAI21_X1 U7050 ( .B1(n6873), .B2(n6708), .A(n6020), .ZN(U2911) );
  AOI22_X1 U7051 ( .A1(n6041), .A2(LWORD_REG_11__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6021) );
  OAI21_X1 U7052 ( .B1(n5073), .B2(n6043), .A(n6021), .ZN(U2912) );
  AOI222_X1 U7053 ( .A1(n6041), .A2(LWORD_REG_10__SCAN_IN), .B1(n6030), .B2(
        EAX_REG_10__SCAN_IN), .C1(DATAO_REG_10__SCAN_IN), .C2(n6040), .ZN(
        n6022) );
  INV_X1 U7054 ( .A(n6022), .ZN(U2913) );
  INV_X1 U7055 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n7003) );
  OAI222_X1 U7056 ( .A1(n6024), .A2(n6708), .B1(n6043), .B2(n6971), .C1(n6023), 
        .C2(n7003), .ZN(U2914) );
  INV_X1 U7057 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6026) );
  AOI22_X1 U7058 ( .A1(n6041), .A2(LWORD_REG_8__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6025) );
  OAI21_X1 U7059 ( .B1(n6026), .B2(n6043), .A(n6025), .ZN(U2915) );
  AOI222_X1 U7060 ( .A1(n6041), .A2(LWORD_REG_7__SCAN_IN), .B1(n6030), .B2(
        EAX_REG_7__SCAN_IN), .C1(DATAO_REG_7__SCAN_IN), .C2(n6040), .ZN(n6027)
         );
  INV_X1 U7061 ( .A(n6027), .ZN(U2916) );
  INV_X1 U7062 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6029) );
  AOI22_X1 U7063 ( .A1(n6041), .A2(LWORD_REG_6__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6028) );
  OAI21_X1 U7064 ( .B1(n6029), .B2(n6043), .A(n6028), .ZN(U2917) );
  INV_X1 U7065 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n6952) );
  AOI22_X1 U7066 ( .A1(EAX_REG_5__SCAN_IN), .A2(n6030), .B1(n6040), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6031) );
  OAI21_X1 U7067 ( .B1(n6952), .B2(n6708), .A(n6031), .ZN(U2918) );
  AOI22_X1 U7068 ( .A1(n6041), .A2(LWORD_REG_4__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6032) );
  OAI21_X1 U7069 ( .B1(n6033), .B2(n6043), .A(n6032), .ZN(U2919) );
  AOI22_X1 U7070 ( .A1(DATAO_REG_3__SCAN_IN), .A2(n6040), .B1(n6041), .B2(
        LWORD_REG_3__SCAN_IN), .ZN(n6034) );
  OAI21_X1 U7071 ( .B1(n6035), .B2(n6043), .A(n6034), .ZN(U2920) );
  AOI22_X1 U7072 ( .A1(n6041), .A2(LWORD_REG_2__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6036) );
  OAI21_X1 U7073 ( .B1(n6037), .B2(n6043), .A(n6036), .ZN(U2921) );
  AOI22_X1 U7074 ( .A1(n6041), .A2(LWORD_REG_1__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6038) );
  OAI21_X1 U7075 ( .B1(n6039), .B2(n6043), .A(n6038), .ZN(U2922) );
  AOI22_X1 U7076 ( .A1(n6041), .A2(LWORD_REG_0__SCAN_IN), .B1(n6040), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6042) );
  OAI21_X1 U7077 ( .B1(n6044), .B2(n6043), .A(n6042), .ZN(U2923) );
  AOI22_X1 U7078 ( .A1(n6083), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n6077), .ZN(n6046) );
  OAI21_X1 U7079 ( .B1(n6079), .B2(n6065), .A(n6046), .ZN(U2924) );
  AOI22_X1 U7080 ( .A1(n6083), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n6077), .ZN(n6047) );
  OAI21_X1 U7081 ( .B1(n6079), .B2(n6961), .A(n6047), .ZN(U2925) );
  AOI22_X1 U7082 ( .A1(n6083), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n6077), .ZN(n6048) );
  OAI21_X1 U7083 ( .B1(n6079), .B2(n6068), .A(n6048), .ZN(U2926) );
  AOI22_X1 U7084 ( .A1(n6054), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n6077), .ZN(n6049) );
  OAI21_X1 U7085 ( .B1(n6079), .B2(n6070), .A(n6049), .ZN(U2927) );
  AOI22_X1 U7086 ( .A1(n6054), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n6077), .ZN(n6050) );
  OAI21_X1 U7087 ( .B1(n6079), .B2(n6072), .A(n6050), .ZN(U2928) );
  AOI22_X1 U7088 ( .A1(n6054), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n6077), .ZN(n6051) );
  OAI21_X1 U7089 ( .B1(n6079), .B2(n4744), .A(n6051), .ZN(U2929) );
  INV_X1 U7090 ( .A(DATAI_6_), .ZN(n6075) );
  AOI22_X1 U7091 ( .A1(n6054), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n6077), .ZN(n6052) );
  OAI21_X1 U7092 ( .B1(n6079), .B2(n6075), .A(n6052), .ZN(U2930) );
  AOI22_X1 U7093 ( .A1(n6054), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6077), .ZN(n6053) );
  OAI21_X1 U7094 ( .B1(n6079), .B2(n4758), .A(n6053), .ZN(U2931) );
  INV_X1 U7095 ( .A(DATAI_8_), .ZN(n7035) );
  AOI22_X1 U7096 ( .A1(n6054), .A2(UWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n6077), .ZN(n6055) );
  OAI21_X1 U7097 ( .B1(n6079), .B2(n7035), .A(n6055), .ZN(U2932) );
  AOI21_X1 U7098 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n6083), .A(n6056), .ZN(n6057) );
  OAI21_X1 U7099 ( .B1(n4001), .B2(n6085), .A(n6057), .ZN(U2933) );
  AOI21_X1 U7100 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n6083), .A(n6058), .ZN(
        n6059) );
  OAI21_X1 U7101 ( .B1(n6060), .B2(n6085), .A(n6059), .ZN(U2937) );
  NOR2_X1 U7102 ( .A1(n6079), .A2(n6061), .ZN(n6082) );
  AOI21_X1 U7103 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6083), .A(n6082), .ZN(
        n6062) );
  OAI21_X1 U7104 ( .B1(n6063), .B2(n6085), .A(n6062), .ZN(U2938) );
  AOI22_X1 U7105 ( .A1(n6083), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n6077), .ZN(n6064) );
  OAI21_X1 U7106 ( .B1(n6079), .B2(n6065), .A(n6064), .ZN(U2939) );
  AOI22_X1 U7107 ( .A1(n6083), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n6077), .ZN(n6066) );
  OAI21_X1 U7108 ( .B1(n6079), .B2(n6961), .A(n6066), .ZN(U2940) );
  AOI22_X1 U7109 ( .A1(n6083), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6077), .ZN(n6067) );
  OAI21_X1 U7110 ( .B1(n6079), .B2(n6068), .A(n6067), .ZN(U2941) );
  AOI22_X1 U7111 ( .A1(n6083), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6077), .ZN(n6069) );
  OAI21_X1 U7112 ( .B1(n6079), .B2(n6070), .A(n6069), .ZN(U2942) );
  AOI22_X1 U7113 ( .A1(n6083), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6077), .ZN(n6071) );
  OAI21_X1 U7114 ( .B1(n6079), .B2(n6072), .A(n6071), .ZN(U2943) );
  AOI22_X1 U7115 ( .A1(n6083), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6077), .ZN(n6073) );
  OAI21_X1 U7116 ( .B1(n6079), .B2(n4744), .A(n6073), .ZN(U2944) );
  AOI22_X1 U7117 ( .A1(n6083), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n6077), .ZN(n6074) );
  OAI21_X1 U7118 ( .B1(n6079), .B2(n6075), .A(n6074), .ZN(U2945) );
  AOI22_X1 U7119 ( .A1(n6083), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6077), .ZN(n6076) );
  OAI21_X1 U7120 ( .B1(n6079), .B2(n4758), .A(n6076), .ZN(U2946) );
  AOI22_X1 U7121 ( .A1(n6083), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n6077), .ZN(n6078) );
  OAI21_X1 U7122 ( .B1(n6079), .B2(n7035), .A(n6078), .ZN(U2947) );
  AOI21_X1 U7123 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n6083), .A(n6080), .ZN(
        n6081) );
  OAI21_X1 U7124 ( .B1(n5073), .B2(n6085), .A(n6081), .ZN(U2950) );
  AOI21_X1 U7125 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n6083), .A(n6082), .ZN(
        n6084) );
  OAI21_X1 U7126 ( .B1(n6086), .B2(n6085), .A(n6084), .ZN(U2953) );
  AOI22_X1 U7127 ( .A1(n6187), .A2(REIP_REG_11__SCAN_IN), .B1(n6108), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6091) );
  AOI22_X1 U7128 ( .A1(n6089), .A2(n6113), .B1(n6088), .B2(n6087), .ZN(n6090)
         );
  OAI211_X1 U7129 ( .C1(n6093), .C2(n6092), .A(n6091), .B(n6090), .ZN(U2975)
         );
  AOI22_X1 U7130 ( .A1(n6187), .A2(REIP_REG_6__SCAN_IN), .B1(n6108), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6098) );
  AOI22_X1 U7131 ( .A1(n3207), .A2(n4502), .B1(n6113), .B2(n6096), .ZN(n6097)
         );
  OAI211_X1 U7132 ( .C1(n6117), .C2(n6099), .A(n6098), .B(n6097), .ZN(U2980)
         );
  AOI22_X1 U7133 ( .A1(n6187), .A2(REIP_REG_4__SCAN_IN), .B1(n6108), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6106) );
  OAI21_X1 U7134 ( .B1(n6102), .B2(n6101), .A(n6100), .ZN(n6103) );
  INV_X1 U7135 ( .A(n6103), .ZN(n6169) );
  AOI22_X1 U7136 ( .A1(n4502), .A2(n6169), .B1(n6104), .B2(n6113), .ZN(n6105)
         );
  OAI211_X1 U7137 ( .C1(n6117), .C2(n6107), .A(n6106), .B(n6105), .ZN(U2982)
         );
  AOI22_X1 U7138 ( .A1(n6187), .A2(REIP_REG_2__SCAN_IN), .B1(n6108), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6115) );
  XOR2_X1 U7139 ( .A(n6109), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n6110) );
  XNOR2_X1 U7140 ( .A(n6111), .B(n6110), .ZN(n6193) );
  AOI22_X1 U7141 ( .A1(n6113), .A2(n6112), .B1(n6193), .B2(n4502), .ZN(n6114)
         );
  OAI211_X1 U7142 ( .C1(n6117), .C2(n6116), .A(n6115), .B(n6114), .ZN(U2984)
         );
  OAI21_X1 U7143 ( .B1(n6120), .B2(n6119), .A(n6118), .ZN(n6121) );
  INV_X1 U7144 ( .A(n6121), .ZN(n6133) );
  INV_X1 U7145 ( .A(n6122), .ZN(n6128) );
  INV_X1 U7146 ( .A(n6123), .ZN(n6124) );
  NOR2_X1 U7147 ( .A1(n6124), .A2(n6190), .ZN(n6126) );
  OAI21_X1 U7148 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6126), .A(n6125), 
        .ZN(n6127) );
  AOI22_X1 U7149 ( .A1(n6128), .A2(n4243), .B1(INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n6127), .ZN(n6132) );
  NAND3_X1 U7150 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6130), .A3(n6129), .ZN(n6131) );
  NAND3_X1 U7151 ( .A1(n6133), .A2(n6132), .A3(n6131), .ZN(U3006) );
  AOI21_X1 U7152 ( .B1(n6135), .B2(n6189), .A(n6134), .ZN(n6142) );
  AOI22_X1 U7153 ( .A1(n6137), .A2(n4243), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6136), .ZN(n6141) );
  OAI211_X1 U7154 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6139), .B(n6138), .ZN(n6140) );
  NAND3_X1 U7155 ( .A1(n6142), .A2(n6141), .A3(n6140), .ZN(U3008) );
  INV_X1 U7156 ( .A(n6143), .ZN(n6146) );
  INV_X1 U7157 ( .A(n6144), .ZN(n6145) );
  AOI21_X1 U7158 ( .B1(n6146), .B2(n6189), .A(n6145), .ZN(n6152) );
  INV_X1 U7159 ( .A(n6147), .ZN(n6150) );
  AOI211_X1 U7160 ( .C1(n6159), .C2(n6153), .A(n6148), .B(n6160), .ZN(n6149)
         );
  AOI21_X1 U7161 ( .B1(n6150), .B2(n4243), .A(n6149), .ZN(n6151) );
  OAI211_X1 U7162 ( .C1(n6158), .C2(n6153), .A(n6152), .B(n6151), .ZN(U3010)
         );
  INV_X1 U7163 ( .A(n6154), .ZN(n6155) );
  AOI222_X1 U7164 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6187), .B1(n6189), .B2(
        n6156), .C1(n4243), .C2(n6155), .ZN(n6157) );
  OAI221_X1 U7165 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n6160), .C1(n6159), .C2(n6158), .A(n6157), .ZN(U3011) );
  INV_X1 U7166 ( .A(n6161), .ZN(n6162) );
  AOI22_X1 U7167 ( .A1(n6162), .A2(n6189), .B1(n6187), .B2(REIP_REG_6__SCAN_IN), .ZN(n6165) );
  AOI22_X1 U7168 ( .A1(n3207), .A2(n4243), .B1(n6163), .B2(n6166), .ZN(n6164)
         );
  OAI211_X1 U7169 ( .C1(n6167), .C2(n6166), .A(n6165), .B(n6164), .ZN(U3012)
         );
  AOI21_X1 U7170 ( .B1(n6190), .B2(n6192), .A(n6194), .ZN(n6183) );
  AOI22_X1 U7171 ( .A1(n6168), .A2(n6189), .B1(n6187), .B2(REIP_REG_4__SCAN_IN), .ZN(n6173) );
  AOI211_X1 U7172 ( .C1(n6184), .C2(n6174), .A(n6175), .B(n6192), .ZN(n6171)
         );
  AOI22_X1 U7173 ( .A1(n6171), .A2(n6170), .B1(n4243), .B2(n6169), .ZN(n6172)
         );
  OAI211_X1 U7174 ( .C1(n6183), .C2(n6174), .A(n6173), .B(n6172), .ZN(U3014)
         );
  OR2_X1 U7175 ( .A1(n6192), .A2(n6175), .ZN(n6185) );
  NAND3_X1 U7176 ( .A1(n6176), .A2(n4243), .A3(n4620), .ZN(n6181) );
  NOR2_X1 U7177 ( .A1(n6177), .A2(n4615), .ZN(n6178) );
  AOI21_X1 U7178 ( .B1(n6189), .B2(n6179), .A(n6178), .ZN(n6180) );
  AND2_X1 U7179 ( .A1(n6181), .A2(n6180), .ZN(n6182) );
  OAI221_X1 U7180 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n6185), .C1(n6184), .C2(n6183), .A(n6182), .ZN(U3015) );
  INV_X1 U7181 ( .A(n6186), .ZN(n6188) );
  AOI22_X1 U7182 ( .A1(n6189), .A2(n6188), .B1(n6187), .B2(REIP_REG_2__SCAN_IN), .ZN(n6200) );
  OAI221_X1 U7183 ( .B1(n6192), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .C1(n6192), .C2(n6191), .A(n6190), .ZN(n6199) );
  AOI22_X1 U7184 ( .A1(n6194), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n4243), 
        .B2(n6193), .ZN(n6198) );
  NAND3_X1 U7185 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6196), .A3(n6195), 
        .ZN(n6197) );
  NAND4_X1 U7186 ( .A1(n6200), .A2(n6199), .A3(n6198), .A4(n6197), .ZN(U3016)
         );
  NOR2_X1 U7187 ( .A1(n6202), .A2(n6201), .ZN(U3019) );
  NOR2_X1 U7188 ( .A1(n6580), .A2(n6204), .ZN(n6224) );
  AOI21_X1 U7189 ( .B1(n6203), .B2(n4686), .A(n6224), .ZN(n6206) );
  INV_X1 U7190 ( .A(n6206), .ZN(n6205) );
  INV_X1 U7191 ( .A(n6204), .ZN(n6209) );
  AOI22_X1 U7192 ( .A1(n6207), .A2(n6205), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6209), .ZN(n6229) );
  AOI22_X1 U7193 ( .A1(n6516), .A2(n6224), .B1(n6724), .B2(n6515), .ZN(n6211)
         );
  NAND2_X1 U7194 ( .A1(n6207), .A2(n6206), .ZN(n6208) );
  OAI211_X1 U7195 ( .C1(n6506), .C2(n6209), .A(n6521), .B(n6208), .ZN(n6226)
         );
  AOI22_X1 U7196 ( .A1(n6226), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n6524), 
        .B2(n6225), .ZN(n6210) );
  OAI211_X1 U7197 ( .C1(n6229), .C2(n6723), .A(n6211), .B(n6210), .ZN(U3028)
         );
  AOI22_X1 U7198 ( .A1(n6528), .A2(n6224), .B1(n6724), .B2(n6529), .ZN(n6213)
         );
  AOI22_X1 U7199 ( .A1(n6226), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n6527), 
        .B2(n6225), .ZN(n6212) );
  OAI211_X1 U7200 ( .C1(n6229), .C2(n6532), .A(n6213), .B(n6212), .ZN(U3029)
         );
  AOI22_X1 U7201 ( .A1(n6534), .A2(n6224), .B1(n6724), .B2(n6535), .ZN(n6215)
         );
  AOI22_X1 U7202 ( .A1(n6226), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n6533), 
        .B2(n6225), .ZN(n6214) );
  OAI211_X1 U7203 ( .C1(n6229), .C2(n6538), .A(n6215), .B(n6214), .ZN(U3030)
         );
  AOI22_X1 U7204 ( .A1(n6540), .A2(n6224), .B1(n6724), .B2(n6541), .ZN(n6217)
         );
  AOI22_X1 U7205 ( .A1(n6226), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n6539), 
        .B2(n6225), .ZN(n6216) );
  OAI211_X1 U7206 ( .C1(n6229), .C2(n6544), .A(n6217), .B(n6216), .ZN(U3031)
         );
  AOI22_X1 U7207 ( .A1(n6546), .A2(n6224), .B1(n6724), .B2(n6545), .ZN(n6219)
         );
  AOI22_X1 U7208 ( .A1(n6226), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n6547), 
        .B2(n6225), .ZN(n6218) );
  OAI211_X1 U7209 ( .C1(n6229), .C2(n6550), .A(n6219), .B(n6218), .ZN(U3032)
         );
  AOI22_X1 U7210 ( .A1(n6552), .A2(n6224), .B1(n6724), .B2(n6553), .ZN(n6221)
         );
  AOI22_X1 U7211 ( .A1(n6226), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n6551), 
        .B2(n6225), .ZN(n6220) );
  OAI211_X1 U7212 ( .C1(n6229), .C2(n6556), .A(n6221), .B(n6220), .ZN(U3033)
         );
  AOI22_X1 U7213 ( .A1(n6558), .A2(n6224), .B1(n6724), .B2(n6559), .ZN(n6223)
         );
  AOI22_X1 U7214 ( .A1(n6226), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n6557), 
        .B2(n6225), .ZN(n6222) );
  OAI211_X1 U7215 ( .C1(n6229), .C2(n6562), .A(n6223), .B(n6222), .ZN(U3034)
         );
  AOI22_X1 U7216 ( .A1(n6566), .A2(n6224), .B1(n6724), .B2(n6568), .ZN(n6228)
         );
  AOI22_X1 U7217 ( .A1(n6226), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n6564), 
        .B2(n6225), .ZN(n6227) );
  OAI211_X1 U7218 ( .C1(n6229), .C2(n6572), .A(n6228), .B(n6227), .ZN(U3035)
         );
  NOR2_X1 U7219 ( .A1(n6475), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6252)
         );
  AOI22_X1 U7220 ( .A1(n6524), .A2(n6253), .B1(n6516), .B2(n6252), .ZN(n6239)
         );
  OAI21_X1 U7221 ( .B1(n6231), .B2(n6519), .A(n6472), .ZN(n6234) );
  AOI21_X1 U7222 ( .B1(n6232), .B2(n4686), .A(n6252), .ZN(n6236) );
  AOI22_X1 U7223 ( .A1(n6234), .A2(n6236), .B1(n6235), .B2(n6519), .ZN(n6233)
         );
  NAND2_X1 U7224 ( .A1(n6521), .A2(n6233), .ZN(n6255) );
  INV_X1 U7225 ( .A(n6234), .ZN(n6237) );
  OAI22_X1 U7226 ( .A1(n6237), .A2(n6236), .B1(n6235), .B2(n6505), .ZN(n6254)
         );
  AOI22_X1 U7227 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6255), .B1(n6364), 
        .B2(n6254), .ZN(n6238) );
  OAI211_X1 U7228 ( .C1(n6726), .C2(n6287), .A(n6239), .B(n6238), .ZN(U3044)
         );
  AOI22_X1 U7229 ( .A1(n6527), .A2(n6253), .B1(n6528), .B2(n6252), .ZN(n6241)
         );
  AOI22_X1 U7230 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6255), .B1(n6375), 
        .B2(n6254), .ZN(n6240) );
  OAI211_X1 U7231 ( .C1(n6305), .C2(n6287), .A(n6241), .B(n6240), .ZN(U3045)
         );
  AOI22_X1 U7232 ( .A1(n6533), .A2(n6253), .B1(n6534), .B2(n6252), .ZN(n6243)
         );
  AOI22_X1 U7233 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6255), .B1(n6379), 
        .B2(n6254), .ZN(n6242) );
  OAI211_X1 U7234 ( .C1(n6308), .C2(n6287), .A(n6243), .B(n6242), .ZN(U3046)
         );
  AOI22_X1 U7235 ( .A1(n6539), .A2(n6253), .B1(n6540), .B2(n6252), .ZN(n6245)
         );
  AOI22_X1 U7236 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6255), .B1(n6383), 
        .B2(n6254), .ZN(n6244) );
  OAI211_X1 U7237 ( .C1(n6311), .C2(n6287), .A(n6245), .B(n6244), .ZN(U3047)
         );
  AOI22_X1 U7238 ( .A1(n6547), .A2(n6253), .B1(n6546), .B2(n6252), .ZN(n6247)
         );
  AOI22_X1 U7239 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6255), .B1(n6387), 
        .B2(n6254), .ZN(n6246) );
  OAI211_X1 U7240 ( .C1(n6314), .C2(n6287), .A(n6247), .B(n6246), .ZN(U3048)
         );
  AOI22_X1 U7241 ( .A1(n6551), .A2(n6253), .B1(n6552), .B2(n6252), .ZN(n6249)
         );
  AOI22_X1 U7242 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6255), .B1(n6391), 
        .B2(n6254), .ZN(n6248) );
  OAI211_X1 U7243 ( .C1(n6317), .C2(n6287), .A(n6249), .B(n6248), .ZN(U3049)
         );
  AOI22_X1 U7244 ( .A1(n6557), .A2(n6253), .B1(n6558), .B2(n6252), .ZN(n6251)
         );
  AOI22_X1 U7245 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6255), .B1(n6395), 
        .B2(n6254), .ZN(n6250) );
  OAI211_X1 U7246 ( .C1(n6320), .C2(n6287), .A(n6251), .B(n6250), .ZN(U3050)
         );
  AOI22_X1 U7247 ( .A1(n6564), .A2(n6253), .B1(n6566), .B2(n6252), .ZN(n6257)
         );
  AOI22_X1 U7248 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6255), .B1(n6401), 
        .B2(n6254), .ZN(n6256) );
  OAI211_X1 U7249 ( .C1(n6328), .C2(n6287), .A(n6257), .B(n6256), .ZN(U3051)
         );
  OAI22_X1 U7250 ( .A1(n6292), .A2(n6511), .B1(n6370), .B2(n6258), .ZN(n6282)
         );
  NOR2_X1 U7251 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6259), .ZN(n6281)
         );
  AOI22_X1 U7252 ( .A1(n6364), .A2(n6282), .B1(n6516), .B2(n6281), .ZN(n6268)
         );
  INV_X1 U7253 ( .A(n6281), .ZN(n6261) );
  AOI21_X1 U7254 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6261), .A(n6260), .ZN(
        n6266) );
  INV_X1 U7255 ( .A(n6262), .ZN(n6263) );
  OAI211_X1 U7256 ( .C1(n6287), .C2(n6439), .A(n6264), .B(n6263), .ZN(n6265)
         );
  NAND3_X1 U7257 ( .A1(n6266), .A2(n6361), .A3(n6265), .ZN(n6284) );
  AOI22_X1 U7258 ( .A1(n6284), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n6515), 
        .B2(n6283), .ZN(n6267) );
  OAI211_X1 U7259 ( .C1(n6727), .C2(n6287), .A(n6268), .B(n6267), .ZN(U3052)
         );
  AOI22_X1 U7260 ( .A1(n6375), .A2(n6282), .B1(n6528), .B2(n6281), .ZN(n6270)
         );
  AOI22_X1 U7261 ( .A1(n6284), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n6529), 
        .B2(n6283), .ZN(n6269) );
  OAI211_X1 U7262 ( .C1(n6378), .C2(n6287), .A(n6270), .B(n6269), .ZN(U3053)
         );
  AOI22_X1 U7263 ( .A1(n6379), .A2(n6282), .B1(n6534), .B2(n6281), .ZN(n6272)
         );
  AOI22_X1 U7264 ( .A1(n6284), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n6535), 
        .B2(n6283), .ZN(n6271) );
  OAI211_X1 U7265 ( .C1(n6382), .C2(n6287), .A(n6272), .B(n6271), .ZN(U3054)
         );
  AOI22_X1 U7266 ( .A1(n6383), .A2(n6282), .B1(n6540), .B2(n6281), .ZN(n6274)
         );
  AOI22_X1 U7267 ( .A1(n6284), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n6541), 
        .B2(n6283), .ZN(n6273) );
  OAI211_X1 U7268 ( .C1(n6386), .C2(n6287), .A(n6274), .B(n6273), .ZN(U3055)
         );
  AOI22_X1 U7269 ( .A1(n6387), .A2(n6282), .B1(n6546), .B2(n6281), .ZN(n6276)
         );
  AOI22_X1 U7270 ( .A1(n6284), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n6545), 
        .B2(n6283), .ZN(n6275) );
  OAI211_X1 U7271 ( .C1(n6390), .C2(n6287), .A(n6276), .B(n6275), .ZN(U3056)
         );
  AOI22_X1 U7272 ( .A1(n6391), .A2(n6282), .B1(n6552), .B2(n6281), .ZN(n6278)
         );
  AOI22_X1 U7273 ( .A1(n6284), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n6553), 
        .B2(n6283), .ZN(n6277) );
  OAI211_X1 U7274 ( .C1(n6394), .C2(n6287), .A(n6278), .B(n6277), .ZN(U3057)
         );
  AOI22_X1 U7275 ( .A1(n6395), .A2(n6282), .B1(n6558), .B2(n6281), .ZN(n6280)
         );
  AOI22_X1 U7276 ( .A1(n6284), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n6559), 
        .B2(n6283), .ZN(n6279) );
  OAI211_X1 U7277 ( .C1(n6398), .C2(n6287), .A(n6280), .B(n6279), .ZN(U3058)
         );
  AOI22_X1 U7278 ( .A1(n6401), .A2(n6282), .B1(n6566), .B2(n6281), .ZN(n6286)
         );
  AOI22_X1 U7279 ( .A1(n6284), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n6568), 
        .B2(n6283), .ZN(n6285) );
  OAI211_X1 U7280 ( .C1(n6406), .C2(n6287), .A(n6286), .B(n6285), .ZN(U3059)
         );
  INV_X1 U7281 ( .A(n6296), .ZN(n6291) );
  NAND3_X1 U7282 ( .A1(n6289), .A2(n6288), .A3(n6589), .ZN(n6290) );
  OAI21_X1 U7283 ( .B1(n6292), .B2(n6291), .A(n6290), .ZN(n6322) );
  NAND2_X1 U7284 ( .A1(n6580), .A2(n6336), .ZN(n6297) );
  INV_X1 U7285 ( .A(n6297), .ZN(n6321) );
  AOI22_X1 U7286 ( .A1(n6364), .A2(n6322), .B1(n6516), .B2(n6321), .ZN(n6302)
         );
  NOR3_X1 U7287 ( .A1(n6354), .A2(n6323), .A3(n6519), .ZN(n6294) );
  NOR2_X1 U7288 ( .A1(n6294), .A2(n6439), .ZN(n6300) );
  AND2_X1 U7289 ( .A1(n6296), .A2(n6295), .ZN(n6331) );
  AOI21_X1 U7290 ( .B1(n6297), .B2(STATE2_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6298) );
  OAI211_X1 U7291 ( .C1(n6300), .C2(n6331), .A(n6299), .B(n6298), .ZN(n6324)
         );
  AOI22_X1 U7292 ( .A1(n6324), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6524), 
        .B2(n6323), .ZN(n6301) );
  OAI211_X1 U7293 ( .C1(n6726), .C2(n6327), .A(n6302), .B(n6301), .ZN(U3068)
         );
  AOI22_X1 U7294 ( .A1(n6375), .A2(n6322), .B1(n6528), .B2(n6321), .ZN(n6304)
         );
  AOI22_X1 U7295 ( .A1(n6324), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6527), 
        .B2(n6323), .ZN(n6303) );
  OAI211_X1 U7296 ( .C1(n6305), .C2(n6327), .A(n6304), .B(n6303), .ZN(U3069)
         );
  AOI22_X1 U7297 ( .A1(n6379), .A2(n6322), .B1(n6534), .B2(n6321), .ZN(n6307)
         );
  AOI22_X1 U7298 ( .A1(n6324), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6533), 
        .B2(n6323), .ZN(n6306) );
  OAI211_X1 U7299 ( .C1(n6308), .C2(n6327), .A(n6307), .B(n6306), .ZN(U3070)
         );
  AOI22_X1 U7300 ( .A1(n6383), .A2(n6322), .B1(n6540), .B2(n6321), .ZN(n6310)
         );
  AOI22_X1 U7301 ( .A1(n6324), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6539), 
        .B2(n6323), .ZN(n6309) );
  OAI211_X1 U7302 ( .C1(n6311), .C2(n6327), .A(n6310), .B(n6309), .ZN(U3071)
         );
  AOI22_X1 U7303 ( .A1(n6387), .A2(n6322), .B1(n6546), .B2(n6321), .ZN(n6313)
         );
  AOI22_X1 U7304 ( .A1(n6324), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6547), 
        .B2(n6323), .ZN(n6312) );
  OAI211_X1 U7305 ( .C1(n6314), .C2(n6327), .A(n6313), .B(n6312), .ZN(U3072)
         );
  AOI22_X1 U7306 ( .A1(n6391), .A2(n6322), .B1(n6552), .B2(n6321), .ZN(n6316)
         );
  AOI22_X1 U7307 ( .A1(n6324), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6551), 
        .B2(n6323), .ZN(n6315) );
  OAI211_X1 U7308 ( .C1(n6317), .C2(n6327), .A(n6316), .B(n6315), .ZN(U3073)
         );
  AOI22_X1 U7309 ( .A1(n6395), .A2(n6322), .B1(n6558), .B2(n6321), .ZN(n6319)
         );
  AOI22_X1 U7310 ( .A1(n6324), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6557), 
        .B2(n6323), .ZN(n6318) );
  OAI211_X1 U7311 ( .C1(n6320), .C2(n6327), .A(n6319), .B(n6318), .ZN(U3074)
         );
  AOI22_X1 U7312 ( .A1(n6401), .A2(n6322), .B1(n6566), .B2(n6321), .ZN(n6326)
         );
  AOI22_X1 U7313 ( .A1(n6324), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6564), 
        .B2(n6323), .ZN(n6325) );
  OAI211_X1 U7314 ( .C1(n6328), .C2(n6327), .A(n6326), .B(n6325), .ZN(U3075)
         );
  OAI21_X1 U7315 ( .B1(n6329), .B2(n6519), .A(n6472), .ZN(n6334) );
  INV_X1 U7316 ( .A(n6330), .ZN(n6353) );
  AOI21_X1 U7317 ( .B1(n6331), .B2(n4686), .A(n6353), .ZN(n6333) );
  INV_X1 U7318 ( .A(n6333), .ZN(n6332) );
  AOI22_X1 U7319 ( .A1(n6334), .A2(n6332), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6336), .ZN(n6358) );
  AOI22_X1 U7320 ( .A1(n6516), .A2(n6353), .B1(n6524), .B2(n6354), .ZN(n6340)
         );
  NAND2_X1 U7321 ( .A1(n6334), .A2(n6333), .ZN(n6335) );
  OAI211_X1 U7322 ( .C1(n6336), .C2(n6506), .A(n6521), .B(n6335), .ZN(n6355)
         );
  AOI22_X1 U7323 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6355), .B1(n6515), 
        .B2(n6366), .ZN(n6339) );
  OAI211_X1 U7324 ( .C1(n6358), .C2(n6723), .A(n6340), .B(n6339), .ZN(U3076)
         );
  AOI22_X1 U7325 ( .A1(n6528), .A2(n6353), .B1(n6366), .B2(n6529), .ZN(n6342)
         );
  AOI22_X1 U7326 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6355), .B1(n6527), 
        .B2(n6354), .ZN(n6341) );
  OAI211_X1 U7327 ( .C1(n6358), .C2(n6532), .A(n6342), .B(n6341), .ZN(U3077)
         );
  AOI22_X1 U7328 ( .A1(n6534), .A2(n6353), .B1(n6533), .B2(n6354), .ZN(n6344)
         );
  AOI22_X1 U7329 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6355), .B1(n6535), 
        .B2(n6366), .ZN(n6343) );
  OAI211_X1 U7330 ( .C1(n6358), .C2(n6538), .A(n6344), .B(n6343), .ZN(U3078)
         );
  AOI22_X1 U7331 ( .A1(n6540), .A2(n6353), .B1(n6539), .B2(n6354), .ZN(n6346)
         );
  AOI22_X1 U7332 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6355), .B1(n6541), 
        .B2(n6366), .ZN(n6345) );
  OAI211_X1 U7333 ( .C1(n6358), .C2(n6544), .A(n6346), .B(n6345), .ZN(U3079)
         );
  AOI22_X1 U7334 ( .A1(n6546), .A2(n6353), .B1(n6547), .B2(n6354), .ZN(n6348)
         );
  AOI22_X1 U7335 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6355), .B1(n6545), 
        .B2(n6366), .ZN(n6347) );
  OAI211_X1 U7336 ( .C1(n6358), .C2(n6550), .A(n6348), .B(n6347), .ZN(U3080)
         );
  AOI22_X1 U7337 ( .A1(n6552), .A2(n6353), .B1(n6551), .B2(n6354), .ZN(n6350)
         );
  AOI22_X1 U7338 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6355), .B1(n6553), 
        .B2(n6366), .ZN(n6349) );
  OAI211_X1 U7339 ( .C1(n6358), .C2(n6556), .A(n6350), .B(n6349), .ZN(U3081)
         );
  AOI22_X1 U7340 ( .A1(n6558), .A2(n6353), .B1(n6557), .B2(n6354), .ZN(n6352)
         );
  AOI22_X1 U7341 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6355), .B1(n6559), 
        .B2(n6366), .ZN(n6351) );
  OAI211_X1 U7342 ( .C1(n6358), .C2(n6562), .A(n6352), .B(n6351), .ZN(U3082)
         );
  AOI22_X1 U7343 ( .A1(n6566), .A2(n6353), .B1(n6366), .B2(n6568), .ZN(n6357)
         );
  AOI22_X1 U7344 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6355), .B1(n6564), 
        .B2(n6354), .ZN(n6356) );
  OAI211_X1 U7345 ( .C1(n6358), .C2(n6572), .A(n6357), .B(n6356), .ZN(U3083)
         );
  INV_X1 U7346 ( .A(n6407), .ZN(n6359) );
  NAND3_X1 U7347 ( .A1(n6359), .A2(n6506), .A3(n6441), .ZN(n6360) );
  OAI21_X1 U7348 ( .B1(n6362), .B2(n6361), .A(n6360), .ZN(n6400) );
  NAND3_X1 U7349 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6363), .A3(n6925), .ZN(n6414) );
  NOR2_X1 U7350 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6414), .ZN(n6399)
         );
  AOI22_X1 U7351 ( .A1(n6364), .A2(n6400), .B1(n6516), .B2(n6399), .ZN(n6374)
         );
  NOR3_X1 U7352 ( .A1(n6432), .A2(n6366), .A3(n6519), .ZN(n6368) );
  OAI22_X1 U7353 ( .A1(n6368), .A2(n6439), .B1(n6367), .B2(n6407), .ZN(n6372)
         );
  OR2_X1 U7354 ( .A1(n6399), .A2(n4054), .ZN(n6369) );
  NAND4_X1 U7355 ( .A1(n6372), .A2(n6371), .A3(n6370), .A4(n6369), .ZN(n6402)
         );
  AOI22_X1 U7356 ( .A1(n6402), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6515), 
        .B2(n6432), .ZN(n6373) );
  OAI211_X1 U7357 ( .C1(n6727), .C2(n6405), .A(n6374), .B(n6373), .ZN(U3084)
         );
  AOI22_X1 U7358 ( .A1(n6375), .A2(n6400), .B1(n6528), .B2(n6399), .ZN(n6377)
         );
  AOI22_X1 U7359 ( .A1(n6402), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6432), 
        .B2(n6529), .ZN(n6376) );
  OAI211_X1 U7360 ( .C1(n6378), .C2(n6405), .A(n6377), .B(n6376), .ZN(U3085)
         );
  AOI22_X1 U7361 ( .A1(n6379), .A2(n6400), .B1(n6534), .B2(n6399), .ZN(n6381)
         );
  AOI22_X1 U7362 ( .A1(n6402), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6432), 
        .B2(n6535), .ZN(n6380) );
  OAI211_X1 U7363 ( .C1(n6382), .C2(n6405), .A(n6381), .B(n6380), .ZN(U3086)
         );
  AOI22_X1 U7364 ( .A1(n6383), .A2(n6400), .B1(n6540), .B2(n6399), .ZN(n6385)
         );
  AOI22_X1 U7365 ( .A1(n6402), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6432), 
        .B2(n6541), .ZN(n6384) );
  OAI211_X1 U7366 ( .C1(n6386), .C2(n6405), .A(n6385), .B(n6384), .ZN(U3087)
         );
  AOI22_X1 U7367 ( .A1(n6387), .A2(n6400), .B1(n6546), .B2(n6399), .ZN(n6389)
         );
  AOI22_X1 U7368 ( .A1(n6402), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6432), 
        .B2(n6545), .ZN(n6388) );
  OAI211_X1 U7369 ( .C1(n6390), .C2(n6405), .A(n6389), .B(n6388), .ZN(U3088)
         );
  AOI22_X1 U7370 ( .A1(n6391), .A2(n6400), .B1(n6552), .B2(n6399), .ZN(n6393)
         );
  AOI22_X1 U7371 ( .A1(n6402), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6432), 
        .B2(n6553), .ZN(n6392) );
  OAI211_X1 U7372 ( .C1(n6394), .C2(n6405), .A(n6393), .B(n6392), .ZN(U3089)
         );
  AOI22_X1 U7373 ( .A1(n6395), .A2(n6400), .B1(n6558), .B2(n6399), .ZN(n6397)
         );
  AOI22_X1 U7374 ( .A1(n6402), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6432), 
        .B2(n6559), .ZN(n6396) );
  OAI211_X1 U7375 ( .C1(n6398), .C2(n6405), .A(n6397), .B(n6396), .ZN(U3090)
         );
  AOI22_X1 U7376 ( .A1(n6401), .A2(n6400), .B1(n6566), .B2(n6399), .ZN(n6404)
         );
  AOI22_X1 U7377 ( .A1(n6402), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6432), 
        .B2(n6568), .ZN(n6403) );
  OAI211_X1 U7378 ( .C1(n6406), .C2(n6405), .A(n6404), .B(n6403), .ZN(U3091)
         );
  OR2_X1 U7379 ( .A1(n6512), .A2(n6407), .ZN(n6409) );
  NOR2_X1 U7380 ( .A1(n6580), .A2(n6414), .ZN(n6433) );
  INV_X1 U7381 ( .A(n6433), .ZN(n6408) );
  NAND2_X1 U7382 ( .A1(n6409), .A2(n6408), .ZN(n6417) );
  INV_X1 U7383 ( .A(n6417), .ZN(n6411) );
  OAI21_X1 U7384 ( .B1(n6471), .B2(n6410), .A(n6506), .ZN(n6416) );
  OAI22_X1 U7385 ( .A1(n6505), .A2(n6414), .B1(n6411), .B2(n6416), .ZN(n6412)
         );
  AOI22_X1 U7386 ( .A1(n6516), .A2(n6433), .B1(n6466), .B2(n6515), .ZN(n6419)
         );
  NAND2_X1 U7387 ( .A1(n6519), .A2(n6414), .ZN(n6415) );
  OAI211_X1 U7388 ( .C1(n6417), .C2(n6416), .A(n6521), .B(n6415), .ZN(n6434)
         );
  AOI22_X1 U7389 ( .A1(n6434), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n6524), 
        .B2(n6432), .ZN(n6418) );
  OAI211_X1 U7390 ( .C1(n6437), .C2(n6723), .A(n6419), .B(n6418), .ZN(U3092)
         );
  AOI22_X1 U7391 ( .A1(n6528), .A2(n6433), .B1(n6432), .B2(n6527), .ZN(n6421)
         );
  AOI22_X1 U7392 ( .A1(n6434), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n6466), 
        .B2(n6529), .ZN(n6420) );
  OAI211_X1 U7393 ( .C1(n6437), .C2(n6532), .A(n6421), .B(n6420), .ZN(U3093)
         );
  AOI22_X1 U7394 ( .A1(n6534), .A2(n6433), .B1(n6466), .B2(n6535), .ZN(n6423)
         );
  AOI22_X1 U7395 ( .A1(n6434), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n6533), 
        .B2(n6432), .ZN(n6422) );
  OAI211_X1 U7396 ( .C1(n6437), .C2(n6538), .A(n6423), .B(n6422), .ZN(U3094)
         );
  AOI22_X1 U7397 ( .A1(n6540), .A2(n6433), .B1(n6432), .B2(n6539), .ZN(n6425)
         );
  AOI22_X1 U7398 ( .A1(n6434), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n6466), 
        .B2(n6541), .ZN(n6424) );
  OAI211_X1 U7399 ( .C1(n6437), .C2(n6544), .A(n6425), .B(n6424), .ZN(U3095)
         );
  AOI22_X1 U7400 ( .A1(n6546), .A2(n6433), .B1(n6432), .B2(n6547), .ZN(n6427)
         );
  AOI22_X1 U7401 ( .A1(n6434), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n6466), 
        .B2(n6545), .ZN(n6426) );
  OAI211_X1 U7402 ( .C1(n6437), .C2(n6550), .A(n6427), .B(n6426), .ZN(U3096)
         );
  AOI22_X1 U7403 ( .A1(n6552), .A2(n6433), .B1(n6466), .B2(n6553), .ZN(n6429)
         );
  AOI22_X1 U7404 ( .A1(n6434), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n6551), 
        .B2(n6432), .ZN(n6428) );
  OAI211_X1 U7405 ( .C1(n6437), .C2(n6556), .A(n6429), .B(n6428), .ZN(U3097)
         );
  AOI22_X1 U7406 ( .A1(n6558), .A2(n6433), .B1(n6466), .B2(n6559), .ZN(n6431)
         );
  AOI22_X1 U7407 ( .A1(n6434), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n6557), 
        .B2(n6432), .ZN(n6430) );
  OAI211_X1 U7408 ( .C1(n6437), .C2(n6562), .A(n6431), .B(n6430), .ZN(U3098)
         );
  AOI22_X1 U7409 ( .A1(n6566), .A2(n6433), .B1(n6432), .B2(n6564), .ZN(n6436)
         );
  AOI22_X1 U7410 ( .A1(n6434), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n6466), 
        .B2(n6568), .ZN(n6435) );
  OAI211_X1 U7411 ( .C1(n6437), .C2(n6572), .A(n6436), .B(n6435), .ZN(U3099)
         );
  NOR2_X2 U7412 ( .A1(n6471), .A2(n6438), .ZN(n6500) );
  NOR3_X1 U7413 ( .A1(n6500), .A2(n6466), .A3(n6519), .ZN(n6440) );
  NOR2_X1 U7414 ( .A1(n6440), .A2(n6439), .ZN(n6450) );
  INV_X1 U7415 ( .A(n6450), .ZN(n6444) );
  NAND2_X1 U7416 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6445), .ZN(n6480) );
  NOR2_X1 U7417 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6480), .ZN(n6465)
         );
  AOI22_X1 U7418 ( .A1(n6500), .A2(n6515), .B1(n6516), .B2(n6465), .ZN(n6452)
         );
  INV_X1 U7419 ( .A(n6465), .ZN(n6447) );
  AOI21_X1 U7420 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6447), .A(n6446), .ZN(
        n6448) );
  OAI211_X1 U7421 ( .C1(n6450), .C2(n6474), .A(n6449), .B(n6448), .ZN(n6467)
         );
  AOI22_X1 U7422 ( .A1(n6467), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n6524), 
        .B2(n6466), .ZN(n6451) );
  OAI211_X1 U7423 ( .C1(n6470), .C2(n6723), .A(n6452), .B(n6451), .ZN(U3100)
         );
  AOI22_X1 U7424 ( .A1(n6500), .A2(n6529), .B1(n6528), .B2(n6465), .ZN(n6454)
         );
  AOI22_X1 U7425 ( .A1(n6467), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n6466), 
        .B2(n6527), .ZN(n6453) );
  OAI211_X1 U7426 ( .C1(n6470), .C2(n6532), .A(n6454), .B(n6453), .ZN(U3101)
         );
  AOI22_X1 U7427 ( .A1(n6500), .A2(n6535), .B1(n6534), .B2(n6465), .ZN(n6456)
         );
  AOI22_X1 U7428 ( .A1(n6467), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n6466), 
        .B2(n6533), .ZN(n6455) );
  OAI211_X1 U7429 ( .C1(n6470), .C2(n6538), .A(n6456), .B(n6455), .ZN(U3102)
         );
  AOI22_X1 U7430 ( .A1(n6500), .A2(n6541), .B1(n6540), .B2(n6465), .ZN(n6458)
         );
  AOI22_X1 U7431 ( .A1(n6467), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n6466), 
        .B2(n6539), .ZN(n6457) );
  OAI211_X1 U7432 ( .C1(n6470), .C2(n6544), .A(n6458), .B(n6457), .ZN(U3103)
         );
  AOI22_X1 U7433 ( .A1(n6500), .A2(n6545), .B1(n6546), .B2(n6465), .ZN(n6460)
         );
  AOI22_X1 U7434 ( .A1(n6467), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n6466), 
        .B2(n6547), .ZN(n6459) );
  OAI211_X1 U7435 ( .C1(n6470), .C2(n6550), .A(n6460), .B(n6459), .ZN(U3104)
         );
  AOI22_X1 U7436 ( .A1(n6500), .A2(n6553), .B1(n6552), .B2(n6465), .ZN(n6462)
         );
  AOI22_X1 U7437 ( .A1(n6467), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n6466), 
        .B2(n6551), .ZN(n6461) );
  OAI211_X1 U7438 ( .C1(n6470), .C2(n6556), .A(n6462), .B(n6461), .ZN(U3105)
         );
  AOI22_X1 U7439 ( .A1(n6500), .A2(n6559), .B1(n6558), .B2(n6465), .ZN(n6464)
         );
  AOI22_X1 U7440 ( .A1(n6467), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n6466), 
        .B2(n6557), .ZN(n6463) );
  OAI211_X1 U7441 ( .C1(n6470), .C2(n6562), .A(n6464), .B(n6463), .ZN(U3106)
         );
  AOI22_X1 U7442 ( .A1(n6500), .A2(n6568), .B1(n6566), .B2(n6465), .ZN(n6469)
         );
  AOI22_X1 U7443 ( .A1(n6467), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n6466), 
        .B2(n6564), .ZN(n6468) );
  OAI211_X1 U7444 ( .C1(n6470), .C2(n6572), .A(n6469), .B(n6468), .ZN(U3107)
         );
  INV_X1 U7445 ( .A(n6471), .ZN(n6473) );
  OAI21_X1 U7446 ( .B1(n6473), .B2(n6519), .A(n6472), .ZN(n6482) );
  NAND2_X1 U7447 ( .A1(n6474), .A2(n4686), .ZN(n6477) );
  NOR2_X1 U7448 ( .A1(n6589), .A2(n6475), .ZN(n6498) );
  INV_X1 U7449 ( .A(n6498), .ZN(n6476) );
  NAND2_X1 U7450 ( .A1(n6477), .A2(n6476), .ZN(n6479) );
  INV_X1 U7451 ( .A(n6480), .ZN(n6478) );
  AOI22_X1 U7452 ( .A1(n6482), .A2(n6479), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6478), .ZN(n6504) );
  AOI22_X1 U7453 ( .A1(n6515), .A2(n6499), .B1(n6516), .B2(n6498), .ZN(n6485)
         );
  INV_X1 U7454 ( .A(n6479), .ZN(n6481) );
  AOI22_X1 U7455 ( .A1(n6482), .A2(n6481), .B1(n6480), .B2(n6519), .ZN(n6483)
         );
  NAND2_X1 U7456 ( .A1(n6521), .A2(n6483), .ZN(n6501) );
  AOI22_X1 U7457 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6501), .B1(n6524), 
        .B2(n6500), .ZN(n6484) );
  OAI211_X1 U7458 ( .C1(n6504), .C2(n6723), .A(n6485), .B(n6484), .ZN(U3108)
         );
  AOI22_X1 U7459 ( .A1(n6500), .A2(n6527), .B1(n6528), .B2(n6498), .ZN(n6487)
         );
  AOI22_X1 U7460 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6501), .B1(n6529), 
        .B2(n6499), .ZN(n6486) );
  OAI211_X1 U7461 ( .C1(n6504), .C2(n6532), .A(n6487), .B(n6486), .ZN(U3109)
         );
  AOI22_X1 U7462 ( .A1(n6535), .A2(n6499), .B1(n6534), .B2(n6498), .ZN(n6489)
         );
  AOI22_X1 U7463 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6501), .B1(n6533), 
        .B2(n6500), .ZN(n6488) );
  OAI211_X1 U7464 ( .C1(n6504), .C2(n6538), .A(n6489), .B(n6488), .ZN(U3110)
         );
  AOI22_X1 U7465 ( .A1(n6500), .A2(n6539), .B1(n6540), .B2(n6498), .ZN(n6491)
         );
  AOI22_X1 U7466 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6501), .B1(n6541), 
        .B2(n6499), .ZN(n6490) );
  OAI211_X1 U7467 ( .C1(n6504), .C2(n6544), .A(n6491), .B(n6490), .ZN(U3111)
         );
  AOI22_X1 U7468 ( .A1(n6500), .A2(n6547), .B1(n6546), .B2(n6498), .ZN(n6493)
         );
  AOI22_X1 U7469 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6501), .B1(n6545), 
        .B2(n6499), .ZN(n6492) );
  OAI211_X1 U7470 ( .C1(n6504), .C2(n6550), .A(n6493), .B(n6492), .ZN(U3112)
         );
  AOI22_X1 U7471 ( .A1(n6500), .A2(n6551), .B1(n6552), .B2(n6498), .ZN(n6495)
         );
  AOI22_X1 U7472 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6501), .B1(n6553), 
        .B2(n6499), .ZN(n6494) );
  OAI211_X1 U7473 ( .C1(n6504), .C2(n6556), .A(n6495), .B(n6494), .ZN(U3113)
         );
  AOI22_X1 U7474 ( .A1(n6559), .A2(n6499), .B1(n6558), .B2(n6498), .ZN(n6497)
         );
  AOI22_X1 U7475 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6501), .B1(n6557), 
        .B2(n6500), .ZN(n6496) );
  OAI211_X1 U7476 ( .C1(n6504), .C2(n6562), .A(n6497), .B(n6496), .ZN(U3114)
         );
  AOI22_X1 U7477 ( .A1(n6568), .A2(n6499), .B1(n6566), .B2(n6498), .ZN(n6503)
         );
  AOI22_X1 U7478 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6501), .B1(n6564), 
        .B2(n6500), .ZN(n6502) );
  OAI211_X1 U7479 ( .C1(n6504), .C2(n6572), .A(n6503), .B(n6502), .ZN(U3115)
         );
  NOR2_X1 U7480 ( .A1(n6505), .A2(n6589), .ZN(n6513) );
  NAND2_X1 U7481 ( .A1(n6507), .A2(n6506), .ZN(n6509) );
  NAND2_X1 U7482 ( .A1(n6509), .A2(n6508), .ZN(n6517) );
  NOR2_X1 U7483 ( .A1(n6580), .A2(n6518), .ZN(n6565) );
  INV_X1 U7484 ( .A(n6565), .ZN(n6510) );
  OAI21_X1 U7485 ( .B1(n6512), .B2(n6511), .A(n6510), .ZN(n6522) );
  AOI22_X1 U7486 ( .A1(n6514), .A2(n6513), .B1(n6517), .B2(n6522), .ZN(n6573)
         );
  AOI22_X1 U7487 ( .A1(n6516), .A2(n6565), .B1(n6515), .B2(n6567), .ZN(n6526)
         );
  INV_X1 U7488 ( .A(n6517), .ZN(n6523) );
  NAND2_X1 U7489 ( .A1(n6519), .A2(n6518), .ZN(n6520) );
  OAI211_X1 U7490 ( .C1(n6523), .C2(n6522), .A(n6521), .B(n6520), .ZN(n6569)
         );
  AOI22_X1 U7491 ( .A1(n6569), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n6524), 
        .B2(n6563), .ZN(n6525) );
  OAI211_X1 U7492 ( .C1(n6573), .C2(n6723), .A(n6526), .B(n6525), .ZN(U3124)
         );
  AOI22_X1 U7493 ( .A1(n6528), .A2(n6565), .B1(n6527), .B2(n6563), .ZN(n6531)
         );
  AOI22_X1 U7494 ( .A1(n6569), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n6529), 
        .B2(n6567), .ZN(n6530) );
  OAI211_X1 U7495 ( .C1(n6573), .C2(n6532), .A(n6531), .B(n6530), .ZN(U3125)
         );
  AOI22_X1 U7496 ( .A1(n6534), .A2(n6565), .B1(n6533), .B2(n6563), .ZN(n6537)
         );
  AOI22_X1 U7497 ( .A1(n6569), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n6535), 
        .B2(n6567), .ZN(n6536) );
  OAI211_X1 U7498 ( .C1(n6573), .C2(n6538), .A(n6537), .B(n6536), .ZN(U3126)
         );
  AOI22_X1 U7499 ( .A1(n6540), .A2(n6565), .B1(n6539), .B2(n6563), .ZN(n6543)
         );
  AOI22_X1 U7500 ( .A1(n6569), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n6541), 
        .B2(n6567), .ZN(n6542) );
  OAI211_X1 U7501 ( .C1(n6573), .C2(n6544), .A(n6543), .B(n6542), .ZN(U3127)
         );
  AOI22_X1 U7502 ( .A1(n6546), .A2(n6565), .B1(n6545), .B2(n6567), .ZN(n6549)
         );
  AOI22_X1 U7503 ( .A1(n6569), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n6547), 
        .B2(n6563), .ZN(n6548) );
  OAI211_X1 U7504 ( .C1(n6573), .C2(n6550), .A(n6549), .B(n6548), .ZN(U3128)
         );
  AOI22_X1 U7505 ( .A1(n6552), .A2(n6565), .B1(n6551), .B2(n6563), .ZN(n6555)
         );
  AOI22_X1 U7506 ( .A1(n6569), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n6553), 
        .B2(n6567), .ZN(n6554) );
  OAI211_X1 U7507 ( .C1(n6573), .C2(n6556), .A(n6555), .B(n6554), .ZN(U3129)
         );
  AOI22_X1 U7508 ( .A1(n6558), .A2(n6565), .B1(n6557), .B2(n6563), .ZN(n6561)
         );
  AOI22_X1 U7509 ( .A1(n6569), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n6559), 
        .B2(n6567), .ZN(n6560) );
  OAI211_X1 U7510 ( .C1(n6573), .C2(n6562), .A(n6561), .B(n6560), .ZN(U3130)
         );
  AOI22_X1 U7511 ( .A1(n6566), .A2(n6565), .B1(n6564), .B2(n6563), .ZN(n6571)
         );
  AOI22_X1 U7512 ( .A1(n6569), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n6568), 
        .B2(n6567), .ZN(n6570) );
  OAI211_X1 U7513 ( .C1(n6573), .C2(n6572), .A(n6571), .B(n6570), .ZN(U3131)
         );
  INV_X1 U7514 ( .A(n6577), .ZN(n6575) );
  NOR2_X1 U7515 ( .A1(n6575), .A2(n5733), .ZN(n6590) );
  NAND2_X1 U7516 ( .A1(n6577), .A2(n6576), .ZN(n6587) );
  NAND2_X1 U7517 ( .A1(n6578), .A2(n6577), .ZN(n6583) );
  INV_X1 U7518 ( .A(n6583), .ZN(n6585) );
  AOI211_X1 U7519 ( .C1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n6581), .A(n6580), .B(n6579), .ZN(n6582) );
  OAI21_X1 U7520 ( .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6583), .A(n6582), 
        .ZN(n6584) );
  OAI21_X1 U7521 ( .B1(n6585), .B2(n6925), .A(n6584), .ZN(n6586) );
  AOI222_X1 U7522 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6587), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6586), .C1(n6587), .C2(n6586), 
        .ZN(n6588) );
  AOI222_X1 U7523 ( .A1(n6590), .A2(n6589), .B1(n6590), .B2(n6588), .C1(n6589), 
        .C2(n6588), .ZN(n6593) );
  OAI21_X1 U7524 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6591), 
        .ZN(n6592) );
  OAI21_X1 U7525 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n6593), .A(n6592), 
        .ZN(n6599) );
  NOR2_X1 U7526 ( .A1(n6595), .A2(n6594), .ZN(n6596) );
  NAND2_X1 U7527 ( .A1(n6597), .A2(n6596), .ZN(n6598) );
  INV_X1 U7528 ( .A(n6600), .ZN(n6615) );
  OAI22_X1 U7529 ( .A1(n6600), .A2(n6614), .B1(n6635), .B2(n6708), .ZN(n6606)
         );
  NAND2_X1 U7530 ( .A1(n6602), .A2(n6601), .ZN(n6603) );
  OR2_X1 U7531 ( .A1(n6604), .A2(n6603), .ZN(n6605) );
  OAI21_X1 U7532 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6635), .A(n6698), .ZN(
        n6618) );
  AOI221_X1 U7533 ( .B1(n6608), .B2(STATE2_REG_0__SCAN_IN), .C1(n6618), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6607), .ZN(n6613) );
  OAI211_X1 U7534 ( .C1(n6611), .C2(n6610), .A(n6609), .B(n6698), .ZN(n6612)
         );
  OAI211_X1 U7535 ( .C1(n6615), .C2(n6614), .A(n6613), .B(n6612), .ZN(U3148)
         );
  AOI21_X1 U7536 ( .B1(n6617), .B2(n6635), .A(n6616), .ZN(n6621) );
  NAND3_X1 U7537 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6624), .A3(n6618), .ZN(
        n6619) );
  OAI211_X1 U7538 ( .C1(n6622), .C2(n6621), .A(n6620), .B(n6619), .ZN(U3149)
         );
  INV_X1 U7539 ( .A(n6623), .ZN(n6697) );
  OAI211_X1 U7540 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6635), .A(n6697), .B(
        n6624), .ZN(n6626) );
  OAI21_X1 U7541 ( .B1(n6714), .B2(n6626), .A(n6625), .ZN(U3150) );
  INV_X1 U7542 ( .A(DATAWIDTH_REG_31__SCAN_IN), .ZN(n6951) );
  NOR2_X1 U7543 ( .A1(n6696), .A2(n6951), .ZN(U3151) );
  INV_X1 U7544 ( .A(DATAWIDTH_REG_30__SCAN_IN), .ZN(n6968) );
  NOR2_X1 U7545 ( .A1(n6696), .A2(n6968), .ZN(U3152) );
  INV_X1 U7546 ( .A(DATAWIDTH_REG_29__SCAN_IN), .ZN(n7030) );
  NOR2_X1 U7547 ( .A1(n6696), .A2(n7030), .ZN(U3153) );
  AND2_X1 U7548 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6627), .ZN(U3154) );
  AND2_X1 U7549 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6627), .ZN(U3155) );
  AND2_X1 U7550 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6627), .ZN(U3156) );
  AND2_X1 U7551 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6627), .ZN(U3157) );
  AND2_X1 U7552 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6627), .ZN(U3158) );
  INV_X1 U7553 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n7029) );
  NOR2_X1 U7554 ( .A1(n6696), .A2(n7029), .ZN(U3159) );
  AND2_X1 U7555 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6627), .ZN(U3160) );
  AND2_X1 U7556 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6627), .ZN(U3161) );
  INV_X1 U7557 ( .A(DATAWIDTH_REG_20__SCAN_IN), .ZN(n6841) );
  NOR2_X1 U7558 ( .A1(n6696), .A2(n6841), .ZN(U3162) );
  AND2_X1 U7559 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6627), .ZN(U3163) );
  AND2_X1 U7560 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6627), .ZN(U3164) );
  AND2_X1 U7561 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6627), .ZN(U3165) );
  INV_X1 U7562 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6876) );
  NOR2_X1 U7563 ( .A1(n6696), .A2(n6876), .ZN(U3166) );
  AND2_X1 U7564 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6627), .ZN(U3167) );
  AND2_X1 U7565 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6627), .ZN(U3168) );
  AND2_X1 U7566 ( .A1(n6627), .A2(DATAWIDTH_REG_13__SCAN_IN), .ZN(U3169) );
  INV_X1 U7567 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6796) );
  NOR2_X1 U7568 ( .A1(n6696), .A2(n6796), .ZN(U3170) );
  INV_X1 U7569 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n7019) );
  NOR2_X1 U7570 ( .A1(n6696), .A2(n7019), .ZN(U3171) );
  AND2_X1 U7571 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6627), .ZN(U3172) );
  AND2_X1 U7572 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6627), .ZN(U3173) );
  NOR2_X1 U7573 ( .A1(n6696), .A2(n7010), .ZN(U3174) );
  AND2_X1 U7574 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6627), .ZN(U3175) );
  AND2_X1 U7575 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6627), .ZN(U3176) );
  AND2_X1 U7576 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6627), .ZN(U3177) );
  NOR2_X1 U7577 ( .A1(n6696), .A2(n6990), .ZN(U3178) );
  AND2_X1 U7578 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6627), .ZN(U3179) );
  AND2_X1 U7579 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6627), .ZN(U3180) );
  INV_X1 U7580 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6634) );
  NOR2_X1 U7581 ( .A1(n6645), .A2(n6634), .ZN(n6638) );
  AOI22_X1 U7582 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6642) );
  AND2_X1 U7583 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6631) );
  INV_X1 U7584 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6629) );
  INV_X1 U7585 ( .A(NA_N), .ZN(n6639) );
  AOI211_X1 U7586 ( .C1(STATE_REG_2__SCAN_IN), .C2(n6639), .A(
        STATE_REG_0__SCAN_IN), .B(n6638), .ZN(n6644) );
  AOI221_X1 U7587 ( .B1(n6631), .B2(n6719), .C1(n6629), .C2(n6719), .A(n6644), 
        .ZN(n6628) );
  OAI21_X1 U7588 ( .B1(n6638), .B2(n6642), .A(n6628), .ZN(U3181) );
  NOR2_X1 U7589 ( .A1(n6636), .A2(n6629), .ZN(n6640) );
  NAND2_X1 U7590 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6630) );
  OAI21_X1 U7591 ( .B1(n6640), .B2(n6631), .A(n6630), .ZN(n6632) );
  OAI211_X1 U7592 ( .C1(n6634), .C2(n6635), .A(n6633), .B(n6632), .ZN(U3182)
         );
  AOI221_X1 U7593 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6635), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6637) );
  AOI221_X1 U7594 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6637), .C2(HOLD), .A(n6636), .ZN(n6643) );
  AOI21_X1 U7595 ( .B1(n6640), .B2(n6639), .A(n6638), .ZN(n6641) );
  OAI22_X1 U7596 ( .A1(n6644), .A2(n6643), .B1(n6642), .B2(n6641), .ZN(U3183)
         );
  NOR2_X2 U7597 ( .A1(n6645), .A2(n6719), .ZN(n6687) );
  NAND2_X1 U7598 ( .A1(n6645), .A2(n6678), .ZN(n6689) );
  AOI22_X1 U7599 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6719), .ZN(n6646) );
  OAI21_X1 U7600 ( .B1(n6647), .B2(n6692), .A(n6646), .ZN(U3184) );
  AOI22_X1 U7601 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6719), .ZN(n6648) );
  OAI21_X1 U7602 ( .B1(n6649), .B2(n6692), .A(n6648), .ZN(U3185) );
  AOI22_X1 U7603 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6719), .ZN(n6650) );
  OAI21_X1 U7604 ( .B1(n4615), .B2(n6692), .A(n6650), .ZN(U3186) );
  AOI22_X1 U7605 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6719), .ZN(n6651) );
  OAI21_X1 U7606 ( .B1(n6986), .B2(n6692), .A(n6651), .ZN(U3187) );
  AOI222_X1 U7607 ( .A1(n6690), .A2(REIP_REG_6__SCAN_IN), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6719), .C1(REIP_REG_5__SCAN_IN), .C2(
        n6687), .ZN(n6652) );
  INV_X1 U7608 ( .A(n6652), .ZN(U3188) );
  AOI22_X1 U7609 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6719), .ZN(n6653) );
  OAI21_X1 U7610 ( .B1(n7017), .B2(n6692), .A(n6653), .ZN(U3189) );
  INV_X1 U7611 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6655) );
  AOI22_X1 U7612 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6719), .ZN(n6654) );
  OAI21_X1 U7613 ( .B1(n6655), .B2(n6692), .A(n6654), .ZN(U3190) );
  AOI22_X1 U7614 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6719), .ZN(n6656) );
  OAI21_X1 U7615 ( .B1(n6657), .B2(n6692), .A(n6656), .ZN(U3191) );
  AOI22_X1 U7616 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6719), .ZN(n6658) );
  OAI21_X1 U7617 ( .B1(n6659), .B2(n6692), .A(n6658), .ZN(U3192) );
  AOI22_X1 U7618 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6719), .ZN(n6660) );
  OAI21_X1 U7619 ( .B1(n6661), .B2(n6692), .A(n6660), .ZN(U3193) );
  INV_X1 U7620 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6970) );
  INV_X1 U7621 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n6897) );
  OAI222_X1 U7622 ( .A1(n6692), .A2(n6970), .B1(n6897), .B2(n6678), .C1(n6662), 
        .C2(n6689), .ZN(U3194) );
  AOI222_X1 U7623 ( .A1(n6687), .A2(REIP_REG_12__SCAN_IN), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6719), .C1(REIP_REG_13__SCAN_IN), .C2(
        n6690), .ZN(n6663) );
  INV_X1 U7624 ( .A(n6663), .ZN(U3195) );
  INV_X1 U7625 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n6920) );
  OAI222_X1 U7626 ( .A1(n6692), .A2(n6664), .B1(n6920), .B2(n6678), .C1(n6666), 
        .C2(n6689), .ZN(U3196) );
  AOI22_X1 U7627 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6719), .ZN(n6665) );
  OAI21_X1 U7628 ( .B1(n6666), .B2(n6692), .A(n6665), .ZN(U3197) );
  AOI22_X1 U7629 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6719), .ZN(n6667) );
  OAI21_X1 U7630 ( .B1(n5316), .B2(n6692), .A(n6667), .ZN(U3198) );
  AOI22_X1 U7631 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6687), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6719), .ZN(n6668) );
  OAI21_X1 U7632 ( .B1(n6669), .B2(n6689), .A(n6668), .ZN(U3199) );
  AOI22_X1 U7633 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6687), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6719), .ZN(n6670) );
  OAI21_X1 U7634 ( .B1(n6671), .B2(n6689), .A(n6670), .ZN(U3200) );
  AOI222_X1 U7635 ( .A1(n6687), .A2(REIP_REG_18__SCAN_IN), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6719), .C1(REIP_REG_19__SCAN_IN), .C2(
        n6690), .ZN(n6672) );
  INV_X1 U7636 ( .A(n6672), .ZN(U3201) );
  AOI22_X1 U7637 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6719), .ZN(n6673) );
  OAI21_X1 U7638 ( .B1(n6948), .B2(n6692), .A(n6673), .ZN(U3202) );
  AOI22_X1 U7639 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6687), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6719), .ZN(n6674) );
  OAI21_X1 U7640 ( .B1(n6675), .B2(n6689), .A(n6674), .ZN(U3203) );
  INV_X1 U7641 ( .A(REIP_REG_22__SCAN_IN), .ZN(n7036) );
  AOI22_X1 U7642 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6687), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6719), .ZN(n6676) );
  OAI21_X1 U7643 ( .B1(n7036), .B2(n6689), .A(n6676), .ZN(U3204) );
  INV_X1 U7644 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n7033) );
  OAI222_X1 U7645 ( .A1(n6692), .A2(n7036), .B1(n7033), .B2(n6678), .C1(n6677), 
        .C2(n6689), .ZN(U3205) );
  AOI22_X1 U7646 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6687), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6719), .ZN(n6679) );
  OAI21_X1 U7647 ( .B1(n6984), .B2(n6689), .A(n6679), .ZN(U3206) );
  AOI22_X1 U7648 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6719), .ZN(n6680) );
  OAI21_X1 U7649 ( .B1(n6984), .B2(n6692), .A(n6680), .ZN(U3207) );
  INV_X1 U7650 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6926) );
  AOI22_X1 U7651 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6687), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6719), .ZN(n6681) );
  OAI21_X1 U7652 ( .B1(n6926), .B2(n6689), .A(n6681), .ZN(U3208) );
  AOI22_X1 U7653 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6687), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6719), .ZN(n6682) );
  OAI21_X1 U7654 ( .B1(n6684), .B2(n6689), .A(n6682), .ZN(U3209) );
  AOI22_X1 U7655 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6719), .ZN(n6683) );
  OAI21_X1 U7656 ( .B1(n6684), .B2(n6692), .A(n6683), .ZN(U3210) );
  AOI22_X1 U7657 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6687), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6719), .ZN(n6685) );
  OAI21_X1 U7658 ( .B1(n6686), .B2(n6689), .A(n6685), .ZN(U3211) );
  AOI22_X1 U7659 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6687), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6719), .ZN(n6688) );
  OAI21_X1 U7660 ( .B1(n6693), .B2(n6689), .A(n6688), .ZN(U3212) );
  AOI22_X1 U7661 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6690), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6719), .ZN(n6691) );
  OAI21_X1 U7662 ( .B1(n6693), .B2(n6692), .A(n6691), .ZN(U3213) );
  MUX2_X1 U7663 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6719), .Z(U3445) );
  MUX2_X1 U7664 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6719), .Z(U3446) );
  MUX2_X1 U7665 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6719), .Z(U3447) );
  MUX2_X1 U7666 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6719), .Z(U3448) );
  OAI21_X1 U7667 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6696), .A(n6695), .ZN(
        n6694) );
  INV_X1 U7668 ( .A(n6694), .ZN(U3451) );
  OAI21_X1 U7669 ( .B1(n6696), .B2(n6699), .A(n6695), .ZN(U3452) );
  OAI221_X1 U7670 ( .B1(n4054), .B2(STATE2_REG_0__SCAN_IN), .C1(n4054), .C2(
        n6698), .A(n6697), .ZN(U3453) );
  OAI211_X1 U7671 ( .C1(n6700), .C2(n6829), .A(n6699), .B(n6706), .ZN(n6703)
         );
  NOR2_X1 U7672 ( .A1(n6705), .A2(n6829), .ZN(n6701) );
  AOI22_X1 U7673 ( .A1(BYTEENABLE_REG_2__SCAN_IN), .A2(n6705), .B1(
        REIP_REG_1__SCAN_IN), .B2(n6701), .ZN(n6702) );
  NAND2_X1 U7674 ( .A1(n6703), .A2(n6702), .ZN(U3468) );
  INV_X1 U7675 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6704) );
  AOI22_X1 U7676 ( .A1(n6706), .A2(n6829), .B1(n6705), .B2(n6704), .ZN(U3469)
         );
  NAND2_X1 U7677 ( .A1(n6719), .A2(W_R_N_REG_SCAN_IN), .ZN(n6707) );
  OAI21_X1 U7678 ( .B1(n6719), .B2(READREQUEST_REG_SCAN_IN), .A(n6707), .ZN(
        U3470) );
  OAI21_X1 U7679 ( .B1(READY_N), .B2(n6708), .A(n6519), .ZN(n6709) );
  NOR3_X1 U7680 ( .A1(n6711), .A2(n6710), .A3(n6709), .ZN(n6718) );
  OAI211_X1 U7681 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6713), .A(n6712), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6715) );
  AOI21_X1 U7682 ( .B1(n6715), .B2(STATE2_REG_0__SCAN_IN), .A(n6714), .ZN(
        n6717) );
  NAND2_X1 U7683 ( .A1(n6718), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6716) );
  OAI21_X1 U7684 ( .B1(n6718), .B2(n6717), .A(n6716), .ZN(U3472) );
  MUX2_X1 U7685 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6719), .Z(U3473) );
  OAI22_X1 U7686 ( .A1(n6723), .A2(n6722), .B1(n6721), .B2(n6720), .ZN(n6730)
         );
  INV_X1 U7687 ( .A(n6724), .ZN(n6728) );
  OAI22_X1 U7688 ( .A1(n6728), .A2(n6727), .B1(n6726), .B2(n6725), .ZN(n6729)
         );
  AOI211_X1 U7689 ( .C1(INSTQUEUE_REG_2__0__SCAN_IN), .C2(n6731), .A(n6730), 
        .B(n6729), .ZN(n7124) );
  AOI22_X1 U7690 ( .A1(REIP_REG_7__SCAN_IN), .A2(keyinput241), .B1(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(keyinput214), .ZN(n6732) );
  OAI221_X1 U7691 ( .B1(REIP_REG_7__SCAN_IN), .B2(keyinput241), .C1(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(keyinput214), .A(n6732), .ZN(
        n6739) );
  AOI22_X1 U7692 ( .A1(UWORD_REG_5__SCAN_IN), .A2(keyinput153), .B1(
        EBX_REG_17__SCAN_IN), .B2(keyinput191), .ZN(n6733) );
  OAI221_X1 U7693 ( .B1(UWORD_REG_5__SCAN_IN), .B2(keyinput153), .C1(
        EBX_REG_17__SCAN_IN), .C2(keyinput191), .A(n6733), .ZN(n6738) );
  AOI22_X1 U7694 ( .A1(INSTQUEUE_REG_6__6__SCAN_IN), .A2(keyinput148), .B1(
        INSTQUEUE_REG_7__7__SCAN_IN), .B2(keyinput253), .ZN(n6734) );
  OAI221_X1 U7695 ( .B1(INSTQUEUE_REG_6__6__SCAN_IN), .B2(keyinput148), .C1(
        INSTQUEUE_REG_7__7__SCAN_IN), .C2(keyinput253), .A(n6734), .ZN(n6737)
         );
  AOI22_X1 U7696 ( .A1(ADDRESS_REG_21__SCAN_IN), .A2(keyinput198), .B1(
        DATAWIDTH_REG_13__SCAN_IN), .B2(keyinput248), .ZN(n6735) );
  OAI221_X1 U7697 ( .B1(ADDRESS_REG_21__SCAN_IN), .B2(keyinput198), .C1(
        DATAWIDTH_REG_13__SCAN_IN), .C2(keyinput248), .A(n6735), .ZN(n6736) );
  NOR4_X1 U7698 ( .A1(n6739), .A2(n6738), .A3(n6737), .A4(n6736), .ZN(n6767)
         );
  AOI22_X1 U7699 ( .A1(ADS_N_REG_SCAN_IN), .A2(keyinput240), .B1(
        REIP_REG_19__SCAN_IN), .B2(keyinput144), .ZN(n6740) );
  OAI221_X1 U7700 ( .B1(ADS_N_REG_SCAN_IN), .B2(keyinput240), .C1(
        REIP_REG_19__SCAN_IN), .C2(keyinput144), .A(n6740), .ZN(n6747) );
  AOI22_X1 U7701 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(keyinput200), 
        .B1(INSTQUEUE_REG_3__5__SCAN_IN), .B2(keyinput163), .ZN(n6741) );
  OAI221_X1 U7702 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(keyinput200), 
        .C1(INSTQUEUE_REG_3__5__SCAN_IN), .C2(keyinput163), .A(n6741), .ZN(
        n6746) );
  AOI22_X1 U7703 ( .A1(DATAO_REG_10__SCAN_IN), .A2(keyinput152), .B1(
        INSTQUEUE_REG_12__0__SCAN_IN), .B2(keyinput139), .ZN(n6742) );
  OAI221_X1 U7704 ( .B1(DATAO_REG_10__SCAN_IN), .B2(keyinput152), .C1(
        INSTQUEUE_REG_12__0__SCAN_IN), .C2(keyinput139), .A(n6742), .ZN(n6745)
         );
  AOI22_X1 U7705 ( .A1(DATAWIDTH_REG_1__SCAN_IN), .A2(keyinput130), .B1(
        DATAI_1_), .B2(keyinput221), .ZN(n6743) );
  OAI221_X1 U7706 ( .B1(DATAWIDTH_REG_1__SCAN_IN), .B2(keyinput130), .C1(
        DATAI_1_), .C2(keyinput221), .A(n6743), .ZN(n6744) );
  NOR4_X1 U7707 ( .A1(n6747), .A2(n6746), .A3(n6745), .A4(n6744), .ZN(n6766)
         );
  AOI22_X1 U7708 ( .A1(UWORD_REG_10__SCAN_IN), .A2(keyinput162), .B1(
        INSTQUEUE_REG_14__1__SCAN_IN), .B2(keyinput213), .ZN(n6748) );
  OAI221_X1 U7709 ( .B1(UWORD_REG_10__SCAN_IN), .B2(keyinput162), .C1(
        INSTQUEUE_REG_14__1__SCAN_IN), .C2(keyinput213), .A(n6748), .ZN(n6755)
         );
  AOI22_X1 U7710 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(keyinput243), .B1(
        DATAWIDTH_REG_29__SCAN_IN), .B2(keyinput202), .ZN(n6749) );
  OAI221_X1 U7711 ( .B1(DATAWIDTH_REG_23__SCAN_IN), .B2(keyinput243), .C1(
        DATAWIDTH_REG_29__SCAN_IN), .C2(keyinput202), .A(n6749), .ZN(n6754) );
  AOI22_X1 U7712 ( .A1(INSTQUEUE_REG_8__6__SCAN_IN), .A2(keyinput197), .B1(
        INSTQUEUE_REG_13__7__SCAN_IN), .B2(keyinput217), .ZN(n6750) );
  OAI221_X1 U7713 ( .B1(INSTQUEUE_REG_8__6__SCAN_IN), .B2(keyinput197), .C1(
        INSTQUEUE_REG_13__7__SCAN_IN), .C2(keyinput217), .A(n6750), .ZN(n6753)
         );
  AOI22_X1 U7714 ( .A1(D_C_N_REG_SCAN_IN), .A2(keyinput231), .B1(
        PHYADDRPOINTER_REG_14__SCAN_IN), .B2(keyinput199), .ZN(n6751) );
  OAI221_X1 U7715 ( .B1(D_C_N_REG_SCAN_IN), .B2(keyinput231), .C1(
        PHYADDRPOINTER_REG_14__SCAN_IN), .C2(keyinput199), .A(n6751), .ZN(
        n6752) );
  NOR4_X1 U7716 ( .A1(n6755), .A2(n6754), .A3(n6753), .A4(n6752), .ZN(n6765)
         );
  AOI22_X1 U7717 ( .A1(REIP_REG_4__SCAN_IN), .A2(keyinput254), .B1(
        EBX_REG_16__SCAN_IN), .B2(keyinput194), .ZN(n6756) );
  OAI221_X1 U7718 ( .B1(REIP_REG_4__SCAN_IN), .B2(keyinput254), .C1(
        EBX_REG_16__SCAN_IN), .C2(keyinput194), .A(n6756), .ZN(n6763) );
  AOI22_X1 U7719 ( .A1(STATE2_REG_3__SCAN_IN), .A2(keyinput212), .B1(
        INSTQUEUE_REG_11__6__SCAN_IN), .B2(keyinput209), .ZN(n6757) );
  OAI221_X1 U7720 ( .B1(STATE2_REG_3__SCAN_IN), .B2(keyinput212), .C1(
        INSTQUEUE_REG_11__6__SCAN_IN), .C2(keyinput209), .A(n6757), .ZN(n6762)
         );
  AOI22_X1 U7721 ( .A1(INSTQUEUE_REG_4__6__SCAN_IN), .A2(keyinput136), .B1(
        INSTQUEUE_REG_5__7__SCAN_IN), .B2(keyinput211), .ZN(n6758) );
  OAI221_X1 U7722 ( .B1(INSTQUEUE_REG_4__6__SCAN_IN), .B2(keyinput136), .C1(
        INSTQUEUE_REG_5__7__SCAN_IN), .C2(keyinput211), .A(n6758), .ZN(n6761)
         );
  AOI22_X1 U7723 ( .A1(DATAO_REG_3__SCAN_IN), .A2(keyinput235), .B1(
        EAX_REG_28__SCAN_IN), .B2(keyinput179), .ZN(n6759) );
  OAI221_X1 U7724 ( .B1(DATAO_REG_3__SCAN_IN), .B2(keyinput235), .C1(
        EAX_REG_28__SCAN_IN), .C2(keyinput179), .A(n6759), .ZN(n6760) );
  NOR4_X1 U7725 ( .A1(n6763), .A2(n6762), .A3(n6761), .A4(n6760), .ZN(n6764)
         );
  NAND4_X1 U7726 ( .A1(n6767), .A2(n6766), .A3(n6765), .A4(n6764), .ZN(n6915)
         );
  AOI22_X1 U7727 ( .A1(REIP_REG_17__SCAN_IN), .A2(keyinput233), .B1(
        INSTQUEUE_REG_9__3__SCAN_IN), .B2(keyinput146), .ZN(n6768) );
  OAI221_X1 U7728 ( .B1(REIP_REG_17__SCAN_IN), .B2(keyinput233), .C1(
        INSTQUEUE_REG_9__3__SCAN_IN), .C2(keyinput146), .A(n6768), .ZN(n6775)
         );
  AOI22_X1 U7729 ( .A1(ADDRESS_REG_11__SCAN_IN), .A2(keyinput242), .B1(
        DATAI_31_), .B2(keyinput145), .ZN(n6769) );
  OAI221_X1 U7730 ( .B1(ADDRESS_REG_11__SCAN_IN), .B2(keyinput242), .C1(
        DATAI_31_), .C2(keyinput145), .A(n6769), .ZN(n6774) );
  AOI22_X1 U7731 ( .A1(REIP_REG_22__SCAN_IN), .A2(keyinput205), .B1(
        INSTQUEUE_REG_2__4__SCAN_IN), .B2(keyinput229), .ZN(n6770) );
  OAI221_X1 U7732 ( .B1(REIP_REG_22__SCAN_IN), .B2(keyinput205), .C1(
        INSTQUEUE_REG_2__4__SCAN_IN), .C2(keyinput229), .A(n6770), .ZN(n6773)
         );
  AOI22_X1 U7733 ( .A1(REIP_REG_27__SCAN_IN), .A2(keyinput239), .B1(
        INSTQUEUE_REG_15__5__SCAN_IN), .B2(keyinput245), .ZN(n6771) );
  OAI221_X1 U7734 ( .B1(REIP_REG_27__SCAN_IN), .B2(keyinput239), .C1(
        INSTQUEUE_REG_15__5__SCAN_IN), .C2(keyinput245), .A(n6771), .ZN(n6772)
         );
  NOR4_X1 U7735 ( .A1(n6775), .A2(n6774), .A3(n6773), .A4(n6772), .ZN(n6805)
         );
  AOI22_X1 U7736 ( .A1(DATAO_REG_14__SCAN_IN), .A2(keyinput220), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(keyinput222), .ZN(n6776) );
  OAI221_X1 U7737 ( .B1(DATAO_REG_14__SCAN_IN), .B2(keyinput220), .C1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .C2(keyinput222), .A(n6776), .ZN(
        n6783) );
  AOI22_X1 U7738 ( .A1(UWORD_REG_11__SCAN_IN), .A2(keyinput175), .B1(
        INSTQUEUE_REG_5__6__SCAN_IN), .B2(keyinput180), .ZN(n6777) );
  OAI221_X1 U7739 ( .B1(UWORD_REG_11__SCAN_IN), .B2(keyinput175), .C1(
        INSTQUEUE_REG_5__6__SCAN_IN), .C2(keyinput180), .A(n6777), .ZN(n6782)
         );
  AOI22_X1 U7740 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(keyinput159), .B1(
        INSTQUEUE_REG_4__2__SCAN_IN), .B2(keyinput227), .ZN(n6778) );
  OAI221_X1 U7741 ( .B1(INSTQUEUE_REG_1__3__SCAN_IN), .B2(keyinput159), .C1(
        INSTQUEUE_REG_4__2__SCAN_IN), .C2(keyinput227), .A(n6778), .ZN(n6781)
         );
  AOI22_X1 U7742 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(keyinput203), .B1(
        INSTQUEUE_REG_3__0__SCAN_IN), .B2(keyinput215), .ZN(n6779) );
  OAI221_X1 U7743 ( .B1(INSTQUEUE_REG_3__7__SCAN_IN), .B2(keyinput203), .C1(
        INSTQUEUE_REG_3__0__SCAN_IN), .C2(keyinput215), .A(n6779), .ZN(n6780)
         );
  NOR4_X1 U7744 ( .A1(n6783), .A2(n6782), .A3(n6781), .A4(n6780), .ZN(n6804)
         );
  AOI22_X1 U7745 ( .A1(ADDRESS_REG_17__SCAN_IN), .A2(keyinput234), .B1(
        DATAWIDTH_REG_8__SCAN_IN), .B2(keyinput216), .ZN(n6784) );
  OAI221_X1 U7746 ( .B1(ADDRESS_REG_17__SCAN_IN), .B2(keyinput234), .C1(
        DATAWIDTH_REG_8__SCAN_IN), .C2(keyinput216), .A(n6784), .ZN(n6791) );
  AOI22_X1 U7747 ( .A1(FLUSH_REG_SCAN_IN), .A2(keyinput154), .B1(
        INSTQUEUE_REG_6__7__SCAN_IN), .B2(keyinput244), .ZN(n6785) );
  OAI221_X1 U7748 ( .B1(FLUSH_REG_SCAN_IN), .B2(keyinput154), .C1(
        INSTQUEUE_REG_6__7__SCAN_IN), .C2(keyinput244), .A(n6785), .ZN(n6790)
         );
  AOI22_X1 U7749 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(keyinput250), .B1(
        PHYADDRPOINTER_REG_9__SCAN_IN), .B2(keyinput228), .ZN(n6786) );
  OAI221_X1 U7750 ( .B1(DATAWIDTH_REG_31__SCAN_IN), .B2(keyinput250), .C1(
        PHYADDRPOINTER_REG_9__SCAN_IN), .C2(keyinput228), .A(n6786), .ZN(n6789) );
  AOI22_X1 U7751 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(keyinput143), .B1(
        DATAI_8_), .B2(keyinput208), .ZN(n6787) );
  OAI221_X1 U7752 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(keyinput143), .C1(
        DATAI_8_), .C2(keyinput208), .A(n6787), .ZN(n6788) );
  NOR4_X1 U7753 ( .A1(n6791), .A2(n6790), .A3(n6789), .A4(n6788), .ZN(n6803)
         );
  AOI22_X1 U7754 ( .A1(EBX_REG_27__SCAN_IN), .A2(keyinput131), .B1(
        INSTQUEUE_REG_9__5__SCAN_IN), .B2(keyinput193), .ZN(n6792) );
  OAI221_X1 U7755 ( .B1(EBX_REG_27__SCAN_IN), .B2(keyinput131), .C1(
        INSTQUEUE_REG_9__5__SCAN_IN), .C2(keyinput193), .A(n6792), .ZN(n6801)
         );
  AOI22_X1 U7756 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(keyinput195), .B1(
        INSTQUEUE_REG_5__2__SCAN_IN), .B2(keyinput150), .ZN(n6793) );
  OAI221_X1 U7757 ( .B1(DATAWIDTH_REG_30__SCAN_IN), .B2(keyinput195), .C1(
        INSTQUEUE_REG_5__2__SCAN_IN), .C2(keyinput150), .A(n6793), .ZN(n6800)
         );
  AOI22_X1 U7758 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(keyinput206), .B1(
        n6939), .B2(keyinput247), .ZN(n6794) );
  OAI221_X1 U7759 ( .B1(INSTQUEUE_REG_10__5__SCAN_IN), .B2(keyinput206), .C1(
        n6939), .C2(keyinput247), .A(n6794), .ZN(n6799) );
  AOI22_X1 U7760 ( .A1(n6797), .A2(keyinput219), .B1(keyinput142), .B2(n6796), 
        .ZN(n6795) );
  OAI221_X1 U7761 ( .B1(n6797), .B2(keyinput219), .C1(n6796), .C2(keyinput142), 
        .A(n6795), .ZN(n6798) );
  NOR4_X1 U7762 ( .A1(n6801), .A2(n6800), .A3(n6799), .A4(n6798), .ZN(n6802)
         );
  NAND4_X1 U7763 ( .A1(n6805), .A2(n6804), .A3(n6803), .A4(n6802), .ZN(n6914)
         );
  INV_X1 U7764 ( .A(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n6807) );
  INV_X1 U7765 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n6981) );
  AOI22_X1 U7766 ( .A1(n6807), .A2(keyinput252), .B1(keyinput168), .B2(n6981), 
        .ZN(n6806) );
  OAI221_X1 U7767 ( .B1(n6807), .B2(keyinput252), .C1(n6981), .C2(keyinput168), 
        .A(n6806), .ZN(n6814) );
  INV_X1 U7768 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n6950) );
  AOI22_X1 U7769 ( .A1(n6950), .A2(keyinput185), .B1(n7026), .B2(keyinput151), 
        .ZN(n6808) );
  OAI221_X1 U7770 ( .B1(n6950), .B2(keyinput185), .C1(n7026), .C2(keyinput151), 
        .A(n6808), .ZN(n6813) );
  INV_X1 U7771 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n7013) );
  INV_X1 U7772 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n6965) );
  AOI22_X1 U7773 ( .A1(n7013), .A2(keyinput140), .B1(keyinput167), .B2(n6965), 
        .ZN(n6809) );
  OAI221_X1 U7774 ( .B1(n7013), .B2(keyinput140), .C1(n6965), .C2(keyinput167), 
        .A(n6809), .ZN(n6812) );
  AOI22_X1 U7775 ( .A1(n6919), .A2(keyinput255), .B1(keyinput164), .B2(n7020), 
        .ZN(n6810) );
  OAI221_X1 U7776 ( .B1(n6919), .B2(keyinput255), .C1(n7020), .C2(keyinput164), 
        .A(n6810), .ZN(n6811) );
  NOR4_X1 U7777 ( .A1(n6814), .A2(n6813), .A3(n6812), .A4(n6811), .ZN(n6856)
         );
  AOI22_X1 U7778 ( .A1(n6970), .A2(keyinput182), .B1(keyinput207), .B2(n6816), 
        .ZN(n6815) );
  OAI221_X1 U7779 ( .B1(n6970), .B2(keyinput182), .C1(n6816), .C2(keyinput207), 
        .A(n6815), .ZN(n6826) );
  AOI22_X1 U7780 ( .A1(n4938), .A2(keyinput137), .B1(n7014), .B2(keyinput225), 
        .ZN(n6817) );
  OAI221_X1 U7781 ( .B1(n4938), .B2(keyinput137), .C1(n7014), .C2(keyinput225), 
        .A(n6817), .ZN(n6825) );
  INV_X1 U7782 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n6819) );
  AOI22_X1 U7783 ( .A1(n6820), .A2(keyinput246), .B1(keyinput218), .B2(n6819), 
        .ZN(n6818) );
  OAI221_X1 U7784 ( .B1(n6820), .B2(keyinput246), .C1(n6819), .C2(keyinput218), 
        .A(n6818), .ZN(n6824) );
  INV_X1 U7785 ( .A(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n6967) );
  AOI22_X1 U7786 ( .A1(n6822), .A2(keyinput183), .B1(n6967), .B2(keyinput188), 
        .ZN(n6821) );
  OAI221_X1 U7787 ( .B1(n6822), .B2(keyinput183), .C1(n6967), .C2(keyinput188), 
        .A(n6821), .ZN(n6823) );
  NOR4_X1 U7788 ( .A1(n6826), .A2(n6825), .A3(n6824), .A4(n6823), .ZN(n6855)
         );
  AOI22_X1 U7789 ( .A1(n6829), .A2(keyinput132), .B1(n6828), .B2(keyinput184), 
        .ZN(n6827) );
  OAI221_X1 U7790 ( .B1(n6829), .B2(keyinput132), .C1(n6828), .C2(keyinput184), 
        .A(n6827), .ZN(n6838) );
  AOI22_X1 U7791 ( .A1(n6923), .A2(keyinput134), .B1(n4924), .B2(keyinput135), 
        .ZN(n6830) );
  OAI221_X1 U7792 ( .B1(n6923), .B2(keyinput134), .C1(n4924), .C2(keyinput135), 
        .A(n6830), .ZN(n6837) );
  INV_X1 U7793 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n6932) );
  AOI22_X1 U7794 ( .A1(n6832), .A2(keyinput165), .B1(keyinput147), .B2(n6932), 
        .ZN(n6831) );
  OAI221_X1 U7795 ( .B1(n6832), .B2(keyinput165), .C1(n6932), .C2(keyinput147), 
        .A(n6831), .ZN(n6836) );
  INV_X1 U7796 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6834) );
  AOI22_X1 U7797 ( .A1(n6834), .A2(keyinput232), .B1(keyinput177), .B2(n7017), 
        .ZN(n6833) );
  OAI221_X1 U7798 ( .B1(n6834), .B2(keyinput232), .C1(n7017), .C2(keyinput177), 
        .A(n6833), .ZN(n6835) );
  NOR4_X1 U7799 ( .A1(n6838), .A2(n6837), .A3(n6836), .A4(n6835), .ZN(n6854)
         );
  AOI22_X1 U7800 ( .A1(n6841), .A2(keyinput170), .B1(keyinput189), .B2(n6840), 
        .ZN(n6839) );
  OAI221_X1 U7801 ( .B1(n6841), .B2(keyinput170), .C1(n6840), .C2(keyinput189), 
        .A(n6839), .ZN(n6852) );
  INV_X1 U7802 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6843) );
  AOI22_X1 U7803 ( .A1(n6843), .A2(keyinput210), .B1(keyinput149), .B2(n6952), 
        .ZN(n6842) );
  OAI221_X1 U7804 ( .B1(n6843), .B2(keyinput210), .C1(n6952), .C2(keyinput149), 
        .A(n6842), .ZN(n6851) );
  INV_X1 U7805 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n6845) );
  AOI22_X1 U7806 ( .A1(n6845), .A2(keyinput171), .B1(keyinput186), .B2(n6920), 
        .ZN(n6844) );
  OAI221_X1 U7807 ( .B1(n6845), .B2(keyinput171), .C1(n6920), .C2(keyinput186), 
        .A(n6844), .ZN(n6850) );
  INV_X1 U7808 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n6847) );
  AOI22_X1 U7809 ( .A1(n6848), .A2(keyinput166), .B1(n6847), .B2(keyinput173), 
        .ZN(n6846) );
  OAI221_X1 U7810 ( .B1(n6848), .B2(keyinput166), .C1(n6847), .C2(keyinput173), 
        .A(n6846), .ZN(n6849) );
  NOR4_X1 U7811 ( .A1(n6852), .A2(n6851), .A3(n6850), .A4(n6849), .ZN(n6853)
         );
  NAND4_X1 U7812 ( .A1(n6856), .A2(n6855), .A3(n6854), .A4(n6853), .ZN(n6913)
         );
  AOI22_X1 U7813 ( .A1(n6926), .A2(keyinput190), .B1(n6858), .B2(keyinput141), 
        .ZN(n6857) );
  OAI221_X1 U7814 ( .B1(n6926), .B2(keyinput190), .C1(n6858), .C2(keyinput141), 
        .A(n6857), .ZN(n6868) );
  INV_X1 U7815 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n6861) );
  AOI22_X1 U7816 ( .A1(n6861), .A2(keyinput174), .B1(keyinput181), .B2(n6860), 
        .ZN(n6859) );
  OAI221_X1 U7817 ( .B1(n6861), .B2(keyinput174), .C1(n6860), .C2(keyinput181), 
        .A(n6859), .ZN(n6867) );
  AOI22_X1 U7818 ( .A1(n7003), .A2(keyinput169), .B1(n6984), .B2(keyinput192), 
        .ZN(n6862) );
  OAI221_X1 U7819 ( .B1(n7003), .B2(keyinput169), .C1(n6984), .C2(keyinput192), 
        .A(n6862), .ZN(n6866) );
  AOI22_X1 U7820 ( .A1(n6864), .A2(keyinput160), .B1(keyinput238), .B2(n6998), 
        .ZN(n6863) );
  OAI221_X1 U7821 ( .B1(n6864), .B2(keyinput160), .C1(n6998), .C2(keyinput238), 
        .A(n6863), .ZN(n6865) );
  NOR4_X1 U7822 ( .A1(n6868), .A2(n6867), .A3(n6866), .A4(n6865), .ZN(n6911)
         );
  AOI22_X1 U7823 ( .A1(n6871), .A2(keyinput157), .B1(keyinput237), .B2(n6870), 
        .ZN(n6869) );
  OAI221_X1 U7824 ( .B1(n6871), .B2(keyinput157), .C1(n6870), .C2(keyinput237), 
        .A(n6869), .ZN(n6880) );
  AOI22_X1 U7825 ( .A1(n6941), .A2(keyinput223), .B1(keyinput178), .B2(n6873), 
        .ZN(n6872) );
  OAI221_X1 U7826 ( .B1(n6941), .B2(keyinput223), .C1(n6873), .C2(keyinput178), 
        .A(n6872), .ZN(n6879) );
  AOI22_X1 U7827 ( .A1(n6990), .A2(keyinput129), .B1(n5383), .B2(keyinput224), 
        .ZN(n6874) );
  OAI221_X1 U7828 ( .B1(n6990), .B2(keyinput129), .C1(n5383), .C2(keyinput224), 
        .A(n6874), .ZN(n6878) );
  AOI22_X1 U7829 ( .A1(n6876), .A2(keyinput161), .B1(n4615), .B2(keyinput251), 
        .ZN(n6875) );
  OAI221_X1 U7830 ( .B1(n6876), .B2(keyinput161), .C1(n4615), .C2(keyinput251), 
        .A(n6875), .ZN(n6877) );
  NOR4_X1 U7831 ( .A1(n6880), .A2(n6879), .A3(n6878), .A4(n6877), .ZN(n6910)
         );
  INV_X1 U7832 ( .A(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n6962) );
  AOI22_X1 U7833 ( .A1(n5416), .A2(keyinput176), .B1(n6962), .B2(keyinput133), 
        .ZN(n6881) );
  OAI221_X1 U7834 ( .B1(n5416), .B2(keyinput176), .C1(n6962), .C2(keyinput133), 
        .A(n6881), .ZN(n6882) );
  INV_X1 U7835 ( .A(n6882), .ZN(n6895) );
  INV_X1 U7836 ( .A(BS16_N), .ZN(n6884) );
  AOI22_X1 U7837 ( .A1(n6987), .A2(keyinput128), .B1(keyinput187), .B2(n6884), 
        .ZN(n6883) );
  OAI221_X1 U7838 ( .B1(n6987), .B2(keyinput128), .C1(n6884), .C2(keyinput187), 
        .A(n6883), .ZN(n6885) );
  INV_X1 U7839 ( .A(n6885), .ZN(n6894) );
  AOI22_X1 U7840 ( .A1(n6887), .A2(keyinput204), .B1(keyinput138), .B2(n6933), 
        .ZN(n6886) );
  OAI221_X1 U7841 ( .B1(n6887), .B2(keyinput204), .C1(n6933), .C2(keyinput138), 
        .A(n6886), .ZN(n6890) );
  INV_X1 U7842 ( .A(keyinput155), .ZN(n6888) );
  XNOR2_X1 U7843 ( .A(n6888), .B(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n6889) );
  NOR2_X1 U7844 ( .A1(n6890), .A2(n6889), .ZN(n6893) );
  INV_X1 U7845 ( .A(keyinput156), .ZN(n6891) );
  XNOR2_X1 U7846 ( .A(n7019), .B(n6891), .ZN(n6892) );
  AND4_X1 U7847 ( .A1(n6895), .A2(n6894), .A3(n6893), .A4(n6892), .ZN(n6909)
         );
  INV_X1 U7848 ( .A(UWORD_REG_2__SCAN_IN), .ZN(n7011) );
  AOI22_X1 U7849 ( .A1(n6897), .A2(keyinput226), .B1(keyinput249), .B2(n7011), 
        .ZN(n6896) );
  OAI221_X1 U7850 ( .B1(n6897), .B2(keyinput226), .C1(n7011), .C2(keyinput249), 
        .A(n6896), .ZN(n6907) );
  INV_X1 U7851 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n6900) );
  AOI22_X1 U7852 ( .A1(n6900), .A2(keyinput158), .B1(keyinput230), .B2(n6899), 
        .ZN(n6898) );
  OAI221_X1 U7853 ( .B1(n6900), .B2(keyinput158), .C1(n6899), .C2(keyinput230), 
        .A(n6898), .ZN(n6906) );
  AOI22_X1 U7854 ( .A1(n4579), .A2(keyinput196), .B1(n4896), .B2(keyinput201), 
        .ZN(n6901) );
  OAI221_X1 U7855 ( .B1(n4579), .B2(keyinput196), .C1(n4896), .C2(keyinput201), 
        .A(n6901), .ZN(n6905) );
  XOR2_X1 U7856 ( .A(n6971), .B(keyinput172), .Z(n6903) );
  XNOR2_X1 U7857 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput236), .ZN(
        n6902) );
  NAND2_X1 U7858 ( .A1(n6903), .A2(n6902), .ZN(n6904) );
  NOR4_X1 U7859 ( .A1(n6907), .A2(n6906), .A3(n6905), .A4(n6904), .ZN(n6908)
         );
  NAND4_X1 U7860 ( .A1(n6911), .A2(n6910), .A3(n6909), .A4(n6908), .ZN(n6912)
         );
  NOR4_X1 U7861 ( .A1(n6915), .A2(n6914), .A3(n6913), .A4(n6912), .ZN(n7122)
         );
  AOI22_X1 U7862 ( .A1(n6917), .A2(keyinput34), .B1(n4896), .B2(keyinput73), 
        .ZN(n6916) );
  OAI221_X1 U7863 ( .B1(n6917), .B2(keyinput34), .C1(n4896), .C2(keyinput73), 
        .A(n6916), .ZN(n6930) );
  AOI22_X1 U7864 ( .A1(n6920), .A2(keyinput58), .B1(n6919), .B2(keyinput127), 
        .ZN(n6918) );
  OAI221_X1 U7865 ( .B1(n6920), .B2(keyinput58), .C1(n6919), .C2(keyinput127), 
        .A(n6918), .ZN(n6929) );
  INV_X1 U7866 ( .A(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n6922) );
  AOI22_X1 U7867 ( .A1(n6923), .A2(keyinput6), .B1(n6922), .B2(keyinput75), 
        .ZN(n6921) );
  OAI221_X1 U7868 ( .B1(n6923), .B2(keyinput6), .C1(n6922), .C2(keyinput75), 
        .A(n6921), .ZN(n6928) );
  AOI22_X1 U7869 ( .A1(n6926), .A2(keyinput62), .B1(n6925), .B2(keyinput86), 
        .ZN(n6924) );
  OAI221_X1 U7870 ( .B1(n6926), .B2(keyinput62), .C1(n6925), .C2(keyinput86), 
        .A(n6924), .ZN(n6927) );
  NOR4_X1 U7871 ( .A1(n6930), .A2(n6929), .A3(n6928), .A4(n6927), .ZN(n6979)
         );
  AOI22_X1 U7872 ( .A1(n6933), .A2(keyinput10), .B1(keyinput19), .B2(n6932), 
        .ZN(n6931) );
  OAI221_X1 U7873 ( .B1(n6933), .B2(keyinput10), .C1(n6932), .C2(keyinput19), 
        .A(n6931), .ZN(n6946) );
  INV_X1 U7874 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n6936) );
  INV_X1 U7875 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n6935) );
  AOI22_X1 U7876 ( .A1(n6936), .A2(keyinput99), .B1(n6935), .B2(keyinput81), 
        .ZN(n6934) );
  OAI221_X1 U7877 ( .B1(n6936), .B2(keyinput99), .C1(n6935), .C2(keyinput81), 
        .A(n6934), .ZN(n6945) );
  INV_X1 U7878 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n6938) );
  AOI22_X1 U7879 ( .A1(n6939), .A2(keyinput119), .B1(n6938), .B2(keyinput116), 
        .ZN(n6937) );
  OAI221_X1 U7880 ( .B1(n6939), .B2(keyinput119), .C1(n6938), .C2(keyinput116), 
        .A(n6937), .ZN(n6944) );
  AOI22_X1 U7881 ( .A1(n6942), .A2(keyinput35), .B1(keyinput95), .B2(n6941), 
        .ZN(n6940) );
  OAI221_X1 U7882 ( .B1(n6942), .B2(keyinput35), .C1(n6941), .C2(keyinput95), 
        .A(n6940), .ZN(n6943) );
  NOR4_X1 U7883 ( .A1(n6946), .A2(n6945), .A3(n6944), .A4(n6943), .ZN(n6978)
         );
  AOI22_X1 U7884 ( .A1(n5048), .A2(keyinput22), .B1(keyinput16), .B2(n6948), 
        .ZN(n6947) );
  OAI221_X1 U7885 ( .B1(n5048), .B2(keyinput22), .C1(n6948), .C2(keyinput16), 
        .A(n6947), .ZN(n6959) );
  AOI22_X1 U7886 ( .A1(n6951), .A2(keyinput122), .B1(keyinput57), .B2(n6950), 
        .ZN(n6949) );
  OAI221_X1 U7887 ( .B1(n6951), .B2(keyinput122), .C1(n6950), .C2(keyinput57), 
        .A(n6949), .ZN(n6958) );
  XOR2_X1 U7888 ( .A(n6952), .B(keyinput21), .Z(n6956) );
  XNOR2_X1 U7889 ( .A(keyinput71), .B(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n6955) );
  XNOR2_X1 U7890 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .B(keyinput101), .ZN(n6954) );
  XNOR2_X1 U7891 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput108), .ZN(
        n6953) );
  NAND4_X1 U7892 ( .A1(n6956), .A2(n6955), .A3(n6954), .A4(n6953), .ZN(n6957)
         );
  NOR3_X1 U7893 ( .A1(n6959), .A2(n6958), .A3(n6957), .ZN(n6977) );
  AOI22_X1 U7894 ( .A1(n6962), .A2(keyinput5), .B1(keyinput93), .B2(n6961), 
        .ZN(n6960) );
  OAI221_X1 U7895 ( .B1(n6962), .B2(keyinput5), .C1(n6961), .C2(keyinput93), 
        .A(n6960), .ZN(n6975) );
  INV_X1 U7896 ( .A(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n6964) );
  AOI22_X1 U7897 ( .A1(n6965), .A2(keyinput39), .B1(n6964), .B2(keyinput87), 
        .ZN(n6963) );
  OAI221_X1 U7898 ( .B1(n6965), .B2(keyinput39), .C1(n6964), .C2(keyinput87), 
        .A(n6963), .ZN(n6974) );
  AOI22_X1 U7899 ( .A1(n6968), .A2(keyinput67), .B1(n6967), .B2(keyinput60), 
        .ZN(n6966) );
  OAI221_X1 U7900 ( .B1(n6968), .B2(keyinput67), .C1(n6967), .C2(keyinput60), 
        .A(n6966), .ZN(n6973) );
  AOI22_X1 U7901 ( .A1(n6971), .A2(keyinput44), .B1(keyinput54), .B2(n6970), 
        .ZN(n6969) );
  OAI221_X1 U7902 ( .B1(n6971), .B2(keyinput44), .C1(n6970), .C2(keyinput54), 
        .A(n6969), .ZN(n6972) );
  NOR4_X1 U7903 ( .A1(n6975), .A2(n6974), .A3(n6973), .A4(n6972), .ZN(n6976)
         );
  NAND4_X1 U7904 ( .A1(n6979), .A2(n6978), .A3(n6977), .A4(n6976), .ZN(n7121)
         );
  AOI22_X1 U7905 ( .A1(n6982), .A2(keyinput63), .B1(keyinput40), .B2(n6981), 
        .ZN(n6980) );
  OAI221_X1 U7906 ( .B1(n6982), .B2(keyinput63), .C1(n6981), .C2(keyinput40), 
        .A(n6980), .ZN(n6994) );
  AOI22_X1 U7907 ( .A1(n4924), .A2(keyinput7), .B1(n6984), .B2(keyinput64), 
        .ZN(n6983) );
  OAI221_X1 U7908 ( .B1(n4924), .B2(keyinput7), .C1(n6984), .C2(keyinput64), 
        .A(n6983), .ZN(n6993) );
  AOI22_X1 U7909 ( .A1(n6987), .A2(keyinput0), .B1(keyinput126), .B2(n6986), 
        .ZN(n6985) );
  OAI221_X1 U7910 ( .B1(n6987), .B2(keyinput0), .C1(n6986), .C2(keyinput126), 
        .A(n6985), .ZN(n6992) );
  INV_X1 U7911 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n6989) );
  AOI22_X1 U7912 ( .A1(n6990), .A2(keyinput1), .B1(n6989), .B2(keyinput117), 
        .ZN(n6988) );
  OAI221_X1 U7913 ( .B1(n6990), .B2(keyinput1), .C1(n6989), .C2(keyinput117), 
        .A(n6988), .ZN(n6991) );
  NOR4_X1 U7914 ( .A1(n6994), .A2(n6993), .A3(n6992), .A4(n6991), .ZN(n7044)
         );
  AOI22_X1 U7915 ( .A1(n5383), .A2(keyinput96), .B1(keyinput9), .B2(n4938), 
        .ZN(n6995) );
  OAI221_X1 U7916 ( .B1(n5383), .B2(keyinput96), .C1(n4938), .C2(keyinput9), 
        .A(n6995), .ZN(n7008) );
  AOI22_X1 U7917 ( .A1(n6998), .A2(keyinput110), .B1(n6997), .B2(keyinput100), 
        .ZN(n6996) );
  OAI221_X1 U7918 ( .B1(n6998), .B2(keyinput110), .C1(n6997), .C2(keyinput100), 
        .A(n6996), .ZN(n7007) );
  INV_X1 U7919 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n7001) );
  INV_X1 U7920 ( .A(D_C_N_REG_SCAN_IN), .ZN(n7000) );
  AOI22_X1 U7921 ( .A1(n7001), .A2(keyinput125), .B1(keyinput103), .B2(n7000), 
        .ZN(n6999) );
  OAI221_X1 U7922 ( .B1(n7001), .B2(keyinput125), .C1(n7000), .C2(keyinput103), 
        .A(n6999), .ZN(n7006) );
  AOI22_X1 U7923 ( .A1(n7004), .A2(keyinput72), .B1(keyinput41), .B2(n7003), 
        .ZN(n7002) );
  OAI221_X1 U7924 ( .B1(n7004), .B2(keyinput72), .C1(n7003), .C2(keyinput41), 
        .A(n7002), .ZN(n7005) );
  NOR4_X1 U7925 ( .A1(n7008), .A2(n7007), .A3(n7006), .A4(n7005), .ZN(n7043)
         );
  AOI22_X1 U7926 ( .A1(n7011), .A2(keyinput121), .B1(n7010), .B2(keyinput88), 
        .ZN(n7009) );
  OAI221_X1 U7927 ( .B1(n7011), .B2(keyinput121), .C1(n7010), .C2(keyinput88), 
        .A(n7009), .ZN(n7024) );
  AOI22_X1 U7928 ( .A1(n7014), .A2(keyinput97), .B1(n7013), .B2(keyinput12), 
        .ZN(n7012) );
  OAI221_X1 U7929 ( .B1(n7014), .B2(keyinput97), .C1(n7013), .C2(keyinput12), 
        .A(n7012), .ZN(n7023) );
  AOI22_X1 U7930 ( .A1(n7017), .A2(keyinput49), .B1(keyinput47), .B2(n7016), 
        .ZN(n7015) );
  OAI221_X1 U7931 ( .B1(n7017), .B2(keyinput49), .C1(n7016), .C2(keyinput47), 
        .A(n7015), .ZN(n7022) );
  AOI22_X1 U7932 ( .A1(n7020), .A2(keyinput36), .B1(keyinput28), .B2(n7019), 
        .ZN(n7018) );
  OAI221_X1 U7933 ( .B1(n7020), .B2(keyinput36), .C1(n7019), .C2(keyinput28), 
        .A(n7018), .ZN(n7021) );
  NOR4_X1 U7934 ( .A1(n7024), .A2(n7023), .A3(n7022), .A4(n7021), .ZN(n7042)
         );
  AOI22_X1 U7935 ( .A1(n7027), .A2(keyinput51), .B1(n7026), .B2(keyinput23), 
        .ZN(n7025) );
  OAI221_X1 U7936 ( .B1(n7027), .B2(keyinput51), .C1(n7026), .C2(keyinput23), 
        .A(n7025), .ZN(n7040) );
  AOI22_X1 U7937 ( .A1(n7030), .A2(keyinput74), .B1(keyinput115), .B2(n7029), 
        .ZN(n7028) );
  OAI221_X1 U7938 ( .B1(n7030), .B2(keyinput74), .C1(n7029), .C2(keyinput115), 
        .A(n7028), .ZN(n7039) );
  AOI22_X1 U7939 ( .A1(n7033), .A2(keyinput70), .B1(keyinput26), .B2(n7032), 
        .ZN(n7031) );
  OAI221_X1 U7940 ( .B1(n7033), .B2(keyinput70), .C1(n7032), .C2(keyinput26), 
        .A(n7031), .ZN(n7038) );
  AOI22_X1 U7941 ( .A1(n7036), .A2(keyinput77), .B1(keyinput80), .B2(n7035), 
        .ZN(n7034) );
  OAI221_X1 U7942 ( .B1(n7036), .B2(keyinput77), .C1(n7035), .C2(keyinput80), 
        .A(n7034), .ZN(n7037) );
  NOR4_X1 U7943 ( .A1(n7040), .A2(n7039), .A3(n7038), .A4(n7037), .ZN(n7041)
         );
  NAND4_X1 U7944 ( .A1(n7044), .A2(n7043), .A3(n7042), .A4(n7041), .ZN(n7120)
         );
  OAI22_X1 U7945 ( .A1(INSTQUEUE_REG_4__6__SCAN_IN), .A2(keyinput8), .B1(
        INSTQUEUE_REG_8__6__SCAN_IN), .B2(keyinput69), .ZN(n7045) );
  AOI221_X1 U7946 ( .B1(INSTQUEUE_REG_4__6__SCAN_IN), .B2(keyinput8), .C1(
        keyinput69), .C2(INSTQUEUE_REG_8__6__SCAN_IN), .A(n7045), .ZN(n7052)
         );
  OAI22_X1 U7947 ( .A1(EBX_REG_27__SCAN_IN), .A2(keyinput3), .B1(keyinput37), 
        .B2(STATEBS16_REG_SCAN_IN), .ZN(n7046) );
  AOI221_X1 U7948 ( .B1(EBX_REG_27__SCAN_IN), .B2(keyinput3), .C1(
        STATEBS16_REG_SCAN_IN), .C2(keyinput37), .A(n7046), .ZN(n7051) );
  OAI22_X1 U7949 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(keyinput120), .B1(
        DATAO_REG_10__SCAN_IN), .B2(keyinput24), .ZN(n7047) );
  AOI221_X1 U7950 ( .B1(DATAWIDTH_REG_13__SCAN_IN), .B2(keyinput120), .C1(
        keyinput24), .C2(DATAO_REG_10__SCAN_IN), .A(n7047), .ZN(n7050) );
  OAI22_X1 U7951 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(keyinput89), .B1(
        keyinput56), .B2(DATAI_24_), .ZN(n7048) );
  AOI221_X1 U7952 ( .B1(INSTQUEUE_REG_13__7__SCAN_IN), .B2(keyinput89), .C1(
        DATAI_24_), .C2(keyinput56), .A(n7048), .ZN(n7049) );
  NAND4_X1 U7953 ( .A1(n7052), .A2(n7051), .A3(n7050), .A4(n7049), .ZN(n7080)
         );
  OAI22_X1 U7954 ( .A1(EAX_REG_10__SCAN_IN), .A2(keyinput104), .B1(keyinput59), 
        .B2(BS16_N), .ZN(n7053) );
  AOI221_X1 U7955 ( .B1(EAX_REG_10__SCAN_IN), .B2(keyinput104), .C1(BS16_N), 
        .C2(keyinput59), .A(n7053), .ZN(n7060) );
  OAI22_X1 U7956 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(keyinput55), .B1(
        keyinput109), .B2(EAX_REG_13__SCAN_IN), .ZN(n7054) );
  AOI221_X1 U7957 ( .B1(INSTQUEUE_REG_0__3__SCAN_IN), .B2(keyinput55), .C1(
        EAX_REG_13__SCAN_IN), .C2(keyinput109), .A(n7054), .ZN(n7059) );
  OAI22_X1 U7958 ( .A1(INSTQUEUE_REG_6__5__SCAN_IN), .A2(keyinput30), .B1(
        keyinput27), .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n7055) );
  AOI221_X1 U7959 ( .B1(INSTQUEUE_REG_6__5__SCAN_IN), .B2(keyinput30), .C1(
        INSTQUEUE_REG_0__6__SCAN_IN), .C2(keyinput27), .A(n7055), .ZN(n7058)
         );
  OAI22_X1 U7960 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(keyinput65), .B1(
        INSTQUEUE_REG_4__3__SCAN_IN), .B2(keyinput45), .ZN(n7056) );
  AOI221_X1 U7961 ( .B1(INSTQUEUE_REG_9__5__SCAN_IN), .B2(keyinput65), .C1(
        keyinput45), .C2(INSTQUEUE_REG_4__3__SCAN_IN), .A(n7056), .ZN(n7057)
         );
  NAND4_X1 U7962 ( .A1(n7060), .A2(n7059), .A3(n7058), .A4(n7057), .ZN(n7079)
         );
  OAI22_X1 U7963 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(keyinput38), .B1(
        keyinput17), .B2(DATAI_31_), .ZN(n7061) );
  AOI221_X1 U7964 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(keyinput38), .C1(
        DATAI_31_), .C2(keyinput17), .A(n7061), .ZN(n7068) );
  OAI22_X1 U7965 ( .A1(UWORD_REG_5__SCAN_IN), .A2(keyinput25), .B1(keyinput2), 
        .B2(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7062) );
  AOI221_X1 U7966 ( .B1(UWORD_REG_5__SCAN_IN), .B2(keyinput25), .C1(
        DATAWIDTH_REG_1__SCAN_IN), .C2(keyinput2), .A(n7062), .ZN(n7067) );
  OAI22_X1 U7967 ( .A1(n4833), .A2(keyinput11), .B1(keyinput85), .B2(
        INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n7063) );
  AOI221_X1 U7968 ( .B1(n4833), .B2(keyinput11), .C1(
        INSTQUEUE_REG_14__1__SCAN_IN), .C2(keyinput85), .A(n7063), .ZN(n7066)
         );
  OAI22_X1 U7969 ( .A1(LWORD_REG_10__SCAN_IN), .A2(keyinput61), .B1(
        BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput82), .ZN(n7064) );
  AOI221_X1 U7970 ( .B1(LWORD_REG_10__SCAN_IN), .B2(keyinput61), .C1(
        keyinput82), .C2(BYTEENABLE_REG_3__SCAN_IN), .A(n7064), .ZN(n7065) );
  NAND4_X1 U7971 ( .A1(n7068), .A2(n7067), .A3(n7066), .A4(n7065), .ZN(n7078)
         );
  OAI22_X1 U7972 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(keyinput83), .B1(
        keyinput42), .B2(DATAWIDTH_REG_20__SCAN_IN), .ZN(n7069) );
  AOI221_X1 U7973 ( .B1(INSTQUEUE_REG_5__7__SCAN_IN), .B2(keyinput83), .C1(
        DATAWIDTH_REG_20__SCAN_IN), .C2(keyinput42), .A(n7069), .ZN(n7076) );
  OAI22_X1 U7974 ( .A1(EBX_REG_30__SCAN_IN), .A2(keyinput53), .B1(keyinput15), 
        .B2(REQUESTPENDING_REG_SCAN_IN), .ZN(n7070) );
  AOI221_X1 U7975 ( .B1(EBX_REG_30__SCAN_IN), .B2(keyinput53), .C1(
        REQUESTPENDING_REG_SCAN_IN), .C2(keyinput15), .A(n7070), .ZN(n7075) );
  OAI22_X1 U7976 ( .A1(DATAO_REG_3__SCAN_IN), .A2(keyinput107), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(keyinput98), .ZN(n7071) );
  AOI221_X1 U7977 ( .B1(DATAO_REG_3__SCAN_IN), .B2(keyinput107), .C1(
        keyinput98), .C2(ADDRESS_REG_10__SCAN_IN), .A(n7071), .ZN(n7074) );
  OAI22_X1 U7978 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(keyinput76), .B1(
        keyinput79), .B2(LWORD_REG_13__SCAN_IN), .ZN(n7072) );
  AOI221_X1 U7979 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(keyinput76), 
        .C1(LWORD_REG_13__SCAN_IN), .C2(keyinput79), .A(n7072), .ZN(n7073) );
  NAND4_X1 U7980 ( .A1(n7076), .A2(n7075), .A3(n7074), .A4(n7073), .ZN(n7077)
         );
  NOR4_X1 U7981 ( .A1(n7080), .A2(n7079), .A3(n7078), .A4(n7077), .ZN(n7118)
         );
  OAI22_X1 U7982 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(keyinput43), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(keyinput94), .ZN(n7081) );
  AOI221_X1 U7983 ( .B1(INSTQUEUE_REG_10__4__SCAN_IN), .B2(keyinput43), .C1(
        keyinput94), .C2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n7081), .ZN(n7088) );
  OAI22_X1 U7984 ( .A1(REIP_REG_17__SCAN_IN), .A2(keyinput105), .B1(
        ADS_N_REG_SCAN_IN), .B2(keyinput112), .ZN(n7082) );
  AOI221_X1 U7985 ( .B1(REIP_REG_17__SCAN_IN), .B2(keyinput105), .C1(
        keyinput112), .C2(ADS_N_REG_SCAN_IN), .A(n7082), .ZN(n7087) );
  OAI22_X1 U7986 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(keyinput14), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(keyinput90), .ZN(n7083) );
  AOI221_X1 U7987 ( .B1(DATAWIDTH_REG_12__SCAN_IN), .B2(keyinput14), .C1(
        keyinput90), .C2(ADDRESS_REG_4__SCAN_IN), .A(n7083), .ZN(n7086) );
  OAI22_X1 U7988 ( .A1(ADDRESS_REG_11__SCAN_IN), .A2(keyinput114), .B1(
        keyinput106), .B2(ADDRESS_REG_17__SCAN_IN), .ZN(n7084) );
  AOI221_X1 U7989 ( .B1(ADDRESS_REG_11__SCAN_IN), .B2(keyinput114), .C1(
        ADDRESS_REG_17__SCAN_IN), .C2(keyinput106), .A(n7084), .ZN(n7085) );
  NAND4_X1 U7990 ( .A1(n7088), .A2(n7087), .A3(n7086), .A4(n7085), .ZN(n7116)
         );
  OAI22_X1 U7991 ( .A1(REIP_REG_27__SCAN_IN), .A2(keyinput111), .B1(
        keyinput113), .B2(REIP_REG_7__SCAN_IN), .ZN(n7089) );
  AOI221_X1 U7992 ( .B1(REIP_REG_27__SCAN_IN), .B2(keyinput111), .C1(
        REIP_REG_7__SCAN_IN), .C2(keyinput113), .A(n7089), .ZN(n7096) );
  OAI22_X1 U7993 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(keyinput32), .B1(
        DATAO_REG_14__SCAN_IN), .B2(keyinput92), .ZN(n7090) );
  AOI221_X1 U7994 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(keyinput32), .C1(
        keyinput92), .C2(DATAO_REG_14__SCAN_IN), .A(n7090), .ZN(n7095) );
  OAI22_X1 U7995 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(keyinput78), .B1(
        STATE2_REG_3__SCAN_IN), .B2(keyinput84), .ZN(n7091) );
  AOI221_X1 U7996 ( .B1(INSTQUEUE_REG_10__5__SCAN_IN), .B2(keyinput78), .C1(
        keyinput84), .C2(STATE2_REG_3__SCAN_IN), .A(n7091), .ZN(n7094) );
  OAI22_X1 U7997 ( .A1(EBX_REG_7__SCAN_IN), .A2(keyinput29), .B1(
        EAX_REG_15__SCAN_IN), .B2(keyinput48), .ZN(n7092) );
  AOI221_X1 U7998 ( .B1(EBX_REG_7__SCAN_IN), .B2(keyinput29), .C1(keyinput48), 
        .C2(EAX_REG_15__SCAN_IN), .A(n7092), .ZN(n7093) );
  NAND4_X1 U7999 ( .A1(n7096), .A2(n7095), .A3(n7094), .A4(n7093), .ZN(n7115)
         );
  OAI22_X1 U8000 ( .A1(REIP_REG_0__SCAN_IN), .A2(keyinput4), .B1(
        DATAWIDTH_REG_16__SCAN_IN), .B2(keyinput33), .ZN(n7097) );
  AOI221_X1 U8001 ( .B1(REIP_REG_0__SCAN_IN), .B2(keyinput4), .C1(keyinput33), 
        .C2(DATAWIDTH_REG_16__SCAN_IN), .A(n7097), .ZN(n7104) );
  OAI22_X1 U8002 ( .A1(INSTQUEUE_REG_6__6__SCAN_IN), .A2(keyinput20), .B1(
        REIP_REG_3__SCAN_IN), .B2(keyinput123), .ZN(n7098) );
  AOI221_X1 U8003 ( .B1(INSTQUEUE_REG_6__6__SCAN_IN), .B2(keyinput20), .C1(
        keyinput123), .C2(REIP_REG_3__SCAN_IN), .A(n7098), .ZN(n7103) );
  OAI22_X1 U8004 ( .A1(STATE2_REG_1__SCAN_IN), .A2(keyinput13), .B1(
        INSTADDRPOINTER_REG_11__SCAN_IN), .B2(keyinput102), .ZN(n7099) );
  AOI221_X1 U8005 ( .B1(STATE2_REG_1__SCAN_IN), .B2(keyinput13), .C1(
        keyinput102), .C2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n7099), .ZN(
        n7102) );
  OAI22_X1 U8006 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(keyinput124), .B1(
        keyinput66), .B2(EBX_REG_16__SCAN_IN), .ZN(n7100) );
  AOI221_X1 U8007 ( .B1(INSTQUEUE_REG_3__2__SCAN_IN), .B2(keyinput124), .C1(
        EBX_REG_16__SCAN_IN), .C2(keyinput66), .A(n7100), .ZN(n7101) );
  NAND4_X1 U8008 ( .A1(n7104), .A2(n7103), .A3(n7102), .A4(n7101), .ZN(n7114)
         );
  OAI22_X1 U8009 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(keyinput91), .B1(
        keyinput118), .B2(EBX_REG_13__SCAN_IN), .ZN(n7105) );
  AOI221_X1 U8010 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(keyinput91), 
        .C1(EBX_REG_13__SCAN_IN), .C2(keyinput118), .A(n7105), .ZN(n7112) );
  OAI22_X1 U8011 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(keyinput46), .B1(
        INSTQUEUE_REG_1__3__SCAN_IN), .B2(keyinput31), .ZN(n7106) );
  AOI221_X1 U8012 ( .B1(INSTQUEUE_REG_13__1__SCAN_IN), .B2(keyinput46), .C1(
        keyinput31), .C2(INSTQUEUE_REG_1__3__SCAN_IN), .A(n7106), .ZN(n7111)
         );
  OAI22_X1 U8013 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(keyinput18), .B1(
        LWORD_REG_12__SCAN_IN), .B2(keyinput50), .ZN(n7107) );
  AOI221_X1 U8014 ( .B1(INSTQUEUE_REG_9__3__SCAN_IN), .B2(keyinput18), .C1(
        keyinput50), .C2(LWORD_REG_12__SCAN_IN), .A(n7107), .ZN(n7110) );
  OAI22_X1 U8015 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(keyinput52), .B1(
        LWORD_REG_15__SCAN_IN), .B2(keyinput68), .ZN(n7108) );
  AOI221_X1 U8016 ( .B1(INSTQUEUE_REG_5__6__SCAN_IN), .B2(keyinput52), .C1(
        keyinput68), .C2(LWORD_REG_15__SCAN_IN), .A(n7108), .ZN(n7109) );
  NAND4_X1 U8017 ( .A1(n7112), .A2(n7111), .A3(n7110), .A4(n7109), .ZN(n7113)
         );
  NOR4_X1 U8018 ( .A1(n7116), .A2(n7115), .A3(n7114), .A4(n7113), .ZN(n7117)
         );
  NAND2_X1 U8019 ( .A1(n7118), .A2(n7117), .ZN(n7119) );
  NOR4_X1 U8020 ( .A1(n7122), .A2(n7121), .A3(n7120), .A4(n7119), .ZN(n7123)
         );
  XNOR2_X1 U8021 ( .A(n7124), .B(n7123), .ZN(U3036) );
  BUF_X1 U3642 ( .A(n4383), .Z(n3634) );
  CLKBUF_X1 U3639 ( .A(n3562), .Z(n4686) );
  CLKBUF_X2 U3669 ( .A(n4271), .Z(n3190) );
endmodule

