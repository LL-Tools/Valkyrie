

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2003, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684;

  OR2_X1 U2245 ( .A1(n4018), .A2(n4390), .ZN(n2741) );
  OR2_X1 U2246 ( .A1(n4018), .A2(n4471), .ZN(n2745) );
  NAND3_X1 U2247 ( .A1(n2147), .A2(n2146), .A3(n2045), .ZN(n2152) );
  BUF_X1 U2248 ( .A(n2959), .Z(n3436) );
  BUF_X1 U2249 ( .A(n2448), .Z(n2617) );
  INV_X1 U2250 ( .A(n3433), .ZN(n3396) );
  OR2_X1 U2251 ( .A1(n2615), .A2(n3762), .ZN(n2625) );
  AND2_X1 U2253 ( .A1(n2176), .A2(n2049), .ZN(n4511) );
  CLKBUF_X3 U2254 ( .A(n2338), .Z(n3850) );
  INV_X2 U2255 ( .A(n4623), .ZN(n4289) );
  AND4_X1 U2256 ( .A1(n2315), .A2(n2314), .A3(n2313), .A4(n2312), .ZN(n2003)
         );
  NAND2_X1 U2257 ( .A1(n3931), .A2(n2739), .ZN(n2981) );
  AND2_X2 U2258 ( .A1(n2402), .A2(n2672), .ZN(n3931) );
  AOI21_X2 U2259 ( .B1(n2912), .B2(n2911), .A(n2910), .ZN(n3729) );
  NOR3_X2 U2260 ( .A1(n4284), .A2(n2235), .A3(n4202), .ZN(n2233) );
  OAI21_X2 U2261 ( .B1(n4515), .B2(n4554), .A(n2177), .ZN(n2179) );
  BUF_X2 U2262 ( .A(n2007), .Z(n3846) );
  INV_X2 U2263 ( .A(IR_REG_31__SCAN_IN), .ZN(n2763) );
  AOI21_X1 U2264 ( .B1(n4016), .B2(n4289), .A(n4015), .ZN(n4017) );
  MUX2_X1 U2265 ( .A(n3569), .B(n2744), .S(n4675), .Z(n2746) );
  MUX2_X1 U2266 ( .A(n3570), .B(n2744), .S(n4684), .Z(n2742) );
  AND2_X1 U2267 ( .A1(n2668), .A2(n4011), .ZN(n2744) );
  AOI21_X1 U2268 ( .B1(n2074), .B2(n2073), .A(n2071), .ZN(n4602) );
  NOR2_X1 U2269 ( .A1(n4591), .A2(n2054), .ZN(n2172) );
  OAI21_X1 U2270 ( .B1(n4523), .B2(n4596), .A(n2066), .ZN(n2060) );
  NOR2_X1 U2271 ( .A1(n4592), .A2(n4593), .ZN(n4591) );
  XNOR2_X1 U2272 ( .A(n2133), .B(n4508), .ZN(n4523) );
  NAND2_X1 U2273 ( .A1(n4580), .A2(n2173), .ZN(n4592) );
  OR2_X1 U2274 ( .A1(n4019), .A2(n4029), .ZN(n4021) );
  OR2_X1 U2275 ( .A1(n4597), .A2(n4507), .ZN(n2133) );
  NAND2_X1 U2276 ( .A1(n3701), .A2(n2121), .ZN(n2296) );
  NAND2_X1 U2277 ( .A1(n2599), .A2(n2256), .ZN(n4061) );
  AOI21_X1 U2278 ( .B1(n4088), .B2(n2733), .A(n2047), .ZN(n4073) );
  NAND2_X1 U2279 ( .A1(n4503), .A2(n4566), .ZN(n4578) );
  NAND2_X1 U2280 ( .A1(n4568), .A2(n4567), .ZN(n4566) );
  OAI211_X1 U2281 ( .C1(n4552), .C2(n2143), .A(n2141), .B(n2140), .ZN(n4568)
         );
  NOR2_X1 U2282 ( .A1(n4550), .A2(n4501), .ZN(n4502) );
  NAND2_X1 U2283 ( .A1(n3993), .A2(REG1_REG_14__SCAN_IN), .ZN(n4515) );
  AND2_X1 U2284 ( .A1(n4499), .A2(n4498), .ZN(n4552) );
  NAND2_X1 U2285 ( .A1(n3987), .A2(REG2_REG_14__SCAN_IN), .ZN(n4499) );
  AOI21_X1 U2286 ( .B1(n3990), .B2(n4388), .A(n4539), .ZN(n2174) );
  NAND2_X1 U2287 ( .A1(n3974), .A2(n3973), .ZN(n3984) );
  NAND2_X1 U2288 ( .A1(n2164), .A2(n2166), .ZN(n3989) );
  NAND2_X1 U2289 ( .A1(n2464), .A2(n3804), .ZN(n3132) );
  NAND2_X1 U2290 ( .A1(n3286), .A2(n4487), .ZN(n3288) );
  NOR2_X1 U2291 ( .A1(n2099), .A2(n3322), .ZN(n2098) );
  OR2_X1 U2292 ( .A1(n2600), .A2(n3696), .ZN(n2608) );
  XNOR2_X1 U2293 ( .A(n3053), .B(n3055), .ZN(n3056) );
  AND4_X1 U2294 ( .A1(n2456), .A2(n2455), .A3(n2454), .A4(n2453), .ZN(n3046)
         );
  BUF_X4 U2295 ( .A(n2431), .Z(n3845) );
  AOI21_X1 U2296 ( .B1(n4525), .B2(REG1_REG_4__SCAN_IN), .A(n2069), .ZN(n2833)
         );
  AND2_X1 U2297 ( .A1(n3393), .A2(n4661), .ZN(n2936) );
  BUF_X2 U2298 ( .A(n2956), .Z(n3392) );
  INV_X2 U2299 ( .A(n2240), .ZN(n2432) );
  CLKBUF_X3 U2300 ( .A(n2867), .Z(n3431) );
  INV_X2 U2301 ( .A(n2867), .ZN(n3393) );
  INV_X1 U2302 ( .A(n2956), .ZN(n3337) );
  NAND2_X1 U2303 ( .A1(n2862), .A2(n2981), .ZN(n2867) );
  NAND2_X2 U2304 ( .A1(n3936), .A2(n2981), .ZN(n3433) );
  NAND2_X1 U2305 ( .A1(n2495), .A2(REG3_REG_11__SCAN_IN), .ZN(n2511) );
  XNOR2_X1 U2306 ( .A(n2675), .B(IR_REG_26__SCAN_IN), .ZN(n3415) );
  NAND3_X1 U2307 ( .A1(n2326), .A2(n2325), .A3(n2324), .ZN(n2338) );
  OR2_X1 U2308 ( .A1(n2662), .A2(IR_REG_27__SCAN_IN), .ZN(n2326) );
  OAI21_X1 U2309 ( .B1(n2669), .B2(n2220), .A(IR_REG_31__SCAN_IN), .ZN(n2662)
         );
  NOR2_X1 U2310 ( .A1(n2414), .A2(n2413), .ZN(n2416) );
  AND3_X2 U2311 ( .A1(n2307), .A2(n2330), .A3(n2329), .ZN(n4493) );
  NAND2_X1 U2312 ( .A1(n2180), .A2(n2311), .ZN(n2787) );
  NAND2_X1 U2313 ( .A1(n2311), .A2(n2056), .ZN(n2330) );
  AND2_X1 U2314 ( .A1(n2003), .A2(n2318), .ZN(n2415) );
  AND2_X1 U2315 ( .A1(n2183), .A2(n2181), .ZN(n2180) );
  AND4_X1 U2316 ( .A1(n2317), .A2(n2316), .A3(n2351), .A4(n2406), .ZN(n2318)
         );
  INV_X1 U2317 ( .A(IR_REG_21__SCAN_IN), .ZN(n2398) );
  INV_X1 U2318 ( .A(IR_REG_20__SCAN_IN), .ZN(n2406) );
  NOR2_X1 U2319 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2316)
         );
  INV_X1 U2320 ( .A(IR_REG_2__SCAN_IN), .ZN(n2328) );
  INV_X1 U2321 ( .A(IR_REG_8__SCAN_IN), .ZN(n2351) );
  NOR2_X1 U2322 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2315)
         );
  NOR2_X1 U2323 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2314)
         );
  NOR2_X1 U2324 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2313)
         );
  NOR2_X1 U2325 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2312)
         );
  OAI211_X1 U2326 ( .C1(n3984), .C2(n2155), .A(n2154), .B(1'b1), .ZN(n4496) );
  AOI21_X2 U2328 ( .B1(n4104), .B2(n4281), .A(n4103), .ZN(n4342) );
  AOI21_X2 U2329 ( .B1(n3112), .B2(n3802), .A(n3110), .ZN(n3045) );
  OAI21_X2 U2330 ( .B1(n3132), .B2(n2266), .A(n2263), .ZN(n3203) );
  NOR2_X2 U2331 ( .A1(n2310), .A2(n4172), .ZN(n4162) );
  NAND2_X1 U2332 ( .A1(n2607), .A2(REG3_REG_25__SCAN_IN), .ZN(n2615) );
  INV_X1 U2333 ( .A(n2608), .ZN(n2607) );
  NAND2_X1 U2334 ( .A1(n2322), .A2(n2415), .ZN(n2669) );
  NAND2_X1 U2335 ( .A1(n2145), .A2(n2148), .ZN(n2147) );
  INV_X1 U2336 ( .A(n3058), .ZN(n2148) );
  INV_X1 U2337 ( .A(n2153), .ZN(n2145) );
  AND2_X1 U2338 ( .A1(n2722), .A2(n4265), .ZN(n2724) );
  OAI21_X1 U2339 ( .B1(n2294), .B2(n2022), .A(n3385), .ZN(n2293) );
  INV_X1 U2340 ( .A(n3638), .ZN(n2104) );
  OAI21_X1 U2341 ( .B1(n2959), .B2(n2928), .A(n2915), .ZN(n2916) );
  NAND2_X1 U2342 ( .A1(n2518), .A2(REG3_REG_14__SCAN_IN), .ZN(n2526) );
  INV_X1 U2343 ( .A(n2519), .ZN(n2518) );
  AOI21_X1 U2344 ( .B1(n2209), .B2(n2029), .A(n2212), .ZN(n2208) );
  NOR2_X1 U2345 ( .A1(n4297), .A2(n3631), .ZN(n2212) );
  INV_X1 U2346 ( .A(n2718), .ZN(n2209) );
  AND2_X1 U2347 ( .A1(n2990), .A2(n2702), .ZN(n2222) );
  AND2_X1 U2348 ( .A1(n2367), .A2(n2366), .ZN(n2371) );
  NOR2_X1 U2349 ( .A1(n2305), .A2(n2030), .ZN(n2130) );
  NAND2_X1 U2350 ( .A1(n2130), .A2(n2128), .ZN(n2127) );
  INV_X1 U2351 ( .A(n3625), .ZN(n2128) );
  NAND2_X1 U2352 ( .A1(n2278), .A2(n2277), .ZN(n3242) );
  AND2_X1 U2353 ( .A1(n2870), .A2(n2869), .ZN(n2308) );
  INV_X1 U2354 ( .A(n3737), .ZN(n2945) );
  INV_X1 U2355 ( .A(n2217), .ZN(n2325) );
  NAND2_X1 U2356 ( .A1(n2625), .A2(n2616), .ZN(n2093) );
  INV_X1 U2357 ( .A(n3846), .ZN(n2620) );
  AND2_X1 U2358 ( .A1(n2446), .A2(n2026), .ZN(n2932) );
  OAI21_X1 U2359 ( .B1(n4527), .B2(n2136), .A(n2134), .ZN(n2138) );
  AOI21_X1 U2360 ( .B1(n2139), .B2(n2135), .A(n2829), .ZN(n2134) );
  NOR2_X1 U2361 ( .A1(n2967), .A2(n2966), .ZN(n3053) );
  AND2_X1 U2362 ( .A1(n4489), .A2(REG2_REG_7__SCAN_IN), .ZN(n2966) );
  INV_X1 U2363 ( .A(n3290), .ZN(n2170) );
  OR2_X1 U2364 ( .A1(n3283), .A2(n3282), .ZN(n3974) );
  AOI21_X1 U2365 ( .B1(n2191), .B2(n2190), .A(n2005), .ZN(n2189) );
  INV_X1 U2366 ( .A(n2735), .ZN(n2190) );
  NAND2_X1 U2367 ( .A1(n2356), .A2(n2182), .ZN(n2181) );
  NAND2_X1 U2368 ( .A1(n4578), .A2(n4579), .ZN(n4577) );
  NOR2_X1 U2369 ( .A1(n4109), .A2(n2088), .ZN(n2087) );
  NAND2_X1 U2370 ( .A1(n2042), .A2(n2089), .ZN(n2088) );
  NOR2_X1 U2371 ( .A1(n2091), .A2(n2090), .ZN(n2089) );
  INV_X1 U2372 ( .A(n2724), .ZN(n2205) );
  INV_X1 U2373 ( .A(n3469), .ZN(n2108) );
  AOI22_X1 U2374 ( .A1(n3947), .A2(n3399), .B1(n3392), .B2(n4311), .ZN(n3307)
         );
  AND2_X1 U2375 ( .A1(n4501), .A2(n4638), .ZN(n2142) );
  INV_X1 U2376 ( .A(n4638), .ZN(n2144) );
  INV_X1 U2377 ( .A(n2178), .ZN(n2177) );
  OAI21_X1 U2378 ( .B1(n4514), .B2(n4554), .A(n2046), .ZN(n2178) );
  NOR2_X1 U2379 ( .A1(n2254), .A2(n2253), .ZN(n2252) );
  NOR2_X1 U2380 ( .A1(n2256), .A2(n2255), .ZN(n2253) );
  NAND2_X1 U2381 ( .A1(n2011), .A2(n2025), .ZN(n2200) );
  NOR2_X1 U2382 ( .A1(n2211), .A2(n2718), .ZN(n2210) );
  INV_X1 U2383 ( .A(n2716), .ZN(n2211) );
  NAND2_X1 U2384 ( .A1(n3798), .A2(n3795), .ZN(n2990) );
  INV_X1 U2385 ( .A(n2200), .ZN(n2198) );
  NOR2_X1 U2386 ( .A1(n2730), .A2(n2202), .ZN(n2195) );
  INV_X1 U2387 ( .A(n3867), .ZN(n2197) );
  NAND2_X1 U2388 ( .A1(n2236), .A2(n3671), .ZN(n2235) );
  AND2_X1 U2389 ( .A1(n3820), .A2(n2249), .ZN(n2248) );
  NAND2_X1 U2390 ( .A1(n2008), .A2(n2027), .ZN(n2249) );
  INV_X1 U2391 ( .A(n3813), .ZN(n2250) );
  NAND2_X1 U2392 ( .A1(n2008), .A2(n3817), .ZN(n2251) );
  AND2_X1 U2393 ( .A1(n2009), .A2(n3272), .ZN(n2232) );
  INV_X1 U2394 ( .A(n3810), .ZN(n2268) );
  INV_X1 U2395 ( .A(n3806), .ZN(n2264) );
  NAND2_X1 U2396 ( .A1(n2708), .A2(n2214), .ZN(n2213) );
  NOR2_X1 U2397 ( .A1(n2709), .A2(n2215), .ZN(n2214) );
  INV_X1 U2398 ( .A(n2707), .ZN(n2215) );
  OR2_X1 U2399 ( .A1(n3114), .A2(n3051), .ZN(n2216) );
  INV_X1 U2400 ( .A(IR_REG_27__SCAN_IN), .ZN(n2661) );
  NAND2_X1 U2401 ( .A1(n2398), .A2(n2276), .ZN(n2275) );
  INV_X1 U2402 ( .A(n2275), .ZN(n2274) );
  OR2_X1 U2403 ( .A1(n2400), .A2(n2763), .ZN(n2269) );
  NOR2_X1 U2404 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2317)
         );
  NOR2_X2 U2405 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2327)
         );
  AOI21_X1 U2406 ( .B1(n2287), .B2(n2117), .A(n2116), .ZN(n2115) );
  NAND2_X1 U2407 ( .A1(n3477), .A2(n3381), .ZN(n3480) );
  NAND2_X1 U2408 ( .A1(n2081), .A2(n2033), .ZN(n2481) );
  AND2_X1 U2409 ( .A1(REG3_REG_7__SCAN_IN), .A2(REG3_REG_8__SCAN_IN), .ZN(
        n2471) );
  NAND2_X1 U2410 ( .A1(n3381), .A2(n2297), .ZN(n2291) );
  INV_X1 U2411 ( .A(n2293), .ZN(n2292) );
  AOI22_X1 U2412 ( .A1(n3953), .A2(n3399), .B1(n3000), .B2(n3263), .ZN(n2952)
         );
  XNOR2_X1 U2413 ( .A(n2906), .B(n3433), .ZN(n2937) );
  NAND2_X1 U2414 ( .A1(n3242), .A2(n3241), .ZN(n2131) );
  NAND2_X1 U2415 ( .A1(n3358), .A2(n3357), .ZN(n3359) );
  NAND2_X1 U2416 ( .A1(n2105), .A2(n2103), .ZN(n3360) );
  INV_X1 U2417 ( .A(n3356), .ZN(n3357) );
  NAND2_X1 U2418 ( .A1(n3702), .A2(n3703), .ZN(n3701) );
  NAND2_X1 U2419 ( .A1(n2296), .A2(n2022), .ZN(n3477) );
  NAND2_X1 U2420 ( .A1(n2126), .A2(n2124), .ZN(n3308) );
  NAND2_X1 U2421 ( .A1(n2127), .A2(n2023), .ZN(n2126) );
  AND2_X1 U2422 ( .A1(n2023), .A2(n3241), .ZN(n2125) );
  INV_X1 U2423 ( .A(n2497), .ZN(n2495) );
  NAND2_X1 U2424 ( .A1(n2081), .A2(REG3_REG_6__SCAN_IN), .ZN(n2473) );
  INV_X1 U2425 ( .A(n3656), .ZN(n2289) );
  INV_X1 U2426 ( .A(n4047), .ZN(n3763) );
  OR2_X1 U2428 ( .A1(n2891), .A2(n2881), .ZN(n2889) );
  AND2_X1 U2429 ( .A1(n2863), .A2(n2862), .ZN(n2956) );
  NOR2_X1 U2430 ( .A1(n2078), .A2(n3931), .ZN(n2077) );
  NOR2_X1 U2431 ( .A1(n3898), .A2(n2079), .ZN(n2078) );
  NAND2_X1 U2432 ( .A1(n3900), .A2(n2080), .ZN(n2079) );
  AND2_X1 U2433 ( .A1(n2432), .A2(REG1_REG_3__SCAN_IN), .ZN(n2436) );
  NAND2_X1 U2434 ( .A1(n2688), .A2(n2687), .ZN(n2862) );
  AND2_X1 U2435 ( .A1(n3415), .A2(n4481), .ZN(n2687) );
  NAND2_X1 U2436 ( .A1(n3967), .A2(n2805), .ZN(n2818) );
  OR3_X1 U2437 ( .A1(n2307), .A2(IR_REG_3__SCAN_IN), .A3(IR_REG_4__SCAN_IN), 
        .ZN(n2340) );
  NAND2_X1 U2438 ( .A1(n4491), .A2(REG2_REG_5__SCAN_IN), .ZN(n2137) );
  NAND2_X1 U2439 ( .A1(n3056), .A2(n2150), .ZN(n2146) );
  NOR2_X1 U2440 ( .A1(n3058), .A2(n2151), .ZN(n2150) );
  INV_X1 U2441 ( .A(REG2_REG_8__SCAN_IN), .ZN(n2151) );
  NAND2_X1 U2442 ( .A1(n3054), .A2(n3055), .ZN(n2153) );
  NAND2_X1 U2443 ( .A1(n3167), .A2(n2169), .ZN(n2166) );
  OAI21_X1 U2444 ( .B1(n3288), .B2(n2170), .A(n3978), .ZN(n2165) );
  NAND2_X1 U2445 ( .A1(n4486), .A2(REG2_REG_11__SCAN_IN), .ZN(n3973) );
  XNOR2_X1 U2446 ( .A(n2179), .B(n4638), .ZN(n4571) );
  NAND2_X1 U2447 ( .A1(n4571), .A2(n4570), .ZN(n4569) );
  INV_X1 U2448 ( .A(n4479), .ZN(n3935) );
  NAND2_X1 U2449 ( .A1(n4589), .A2(n4510), .ZN(n2173) );
  NAND2_X1 U2450 ( .A1(n2624), .A2(REG3_REG_27__SCAN_IN), .ZN(n2634) );
  NAND2_X1 U2451 ( .A1(n4061), .A2(n3914), .ZN(n4042) );
  AND2_X1 U2452 ( .A1(n3869), .A2(n3920), .ZN(n4044) );
  INV_X1 U2453 ( .A(n3945), .ZN(n4067) );
  NAND2_X1 U2454 ( .A1(n2566), .A2(REG3_REG_20__SCAN_IN), .ZN(n2583) );
  NAND2_X1 U2455 ( .A1(n2539), .A2(REG3_REG_18__SCAN_IN), .ZN(n2547) );
  INV_X1 U2456 ( .A(n2557), .ZN(n2539) );
  INV_X1 U2457 ( .A(n2092), .ZN(n2555) );
  AND2_X1 U2458 ( .A1(n2721), .A2(n2720), .ZN(n4265) );
  AND2_X1 U2459 ( .A1(n2037), .A2(n2208), .ZN(n2206) );
  NAND2_X1 U2460 ( .A1(n3201), .A2(n2210), .ZN(n2207) );
  INV_X1 U2461 ( .A(n3316), .ZN(n3421) );
  AND2_X1 U2462 ( .A1(n3805), .A2(n3807), .ZN(n3884) );
  NAND2_X1 U2463 ( .A1(n2994), .A2(n2704), .ZN(n3117) );
  INV_X1 U2464 ( .A(IR_REG_19__SCAN_IN), .ZN(n2403) );
  NAND2_X1 U2465 ( .A1(n2393), .A2(n2392), .ZN(n2410) );
  AND2_X1 U2466 ( .A1(n2003), .A2(n2391), .ZN(n2392) );
  AND2_X1 U2467 ( .A1(n2390), .A2(n2389), .ZN(n2391) );
  INV_X1 U2468 ( .A(IR_REG_18__SCAN_IN), .ZN(n2390) );
  INV_X1 U2469 ( .A(n2990), .ZN(n3883) );
  NAND2_X1 U2470 ( .A1(n2439), .A2(n3794), .ZN(n2991) );
  AND2_X1 U2471 ( .A1(n2692), .A2(n2693), .ZN(n2901) );
  AND2_X1 U2472 ( .A1(n2698), .A2(n2697), .ZN(n2880) );
  AND2_X1 U2473 ( .A1(n4082), .A2(n2226), .ZN(n4034) );
  NOR2_X1 U2474 ( .A1(n2227), .A2(n4032), .ZN(n2226) );
  INV_X1 U2475 ( .A(n2228), .ZN(n2227) );
  INV_X1 U2476 ( .A(n3446), .ZN(n3435) );
  NAND2_X1 U2477 ( .A1(n4034), .A2(n3435), .ZN(n2752) );
  NAND2_X1 U2478 ( .A1(n2188), .A2(n2186), .ZN(n4028) );
  AND2_X1 U2479 ( .A1(n2187), .A2(n2304), .ZN(n2186) );
  NAND2_X1 U2480 ( .A1(n4065), .A2(n2734), .ZN(n2735) );
  AOI21_X1 U2481 ( .B1(n4227), .B2(n2726), .A(n2306), .ZN(n4213) );
  INV_X1 U2482 ( .A(n2880), .ZN(n2979) );
  AOI21_X1 U2483 ( .B1(n2275), .B2(IR_REG_31__SCAN_IN), .A(IR_REG_23__SCAN_IN), 
        .ZN(n2273) );
  NAND2_X1 U2484 ( .A1(n2400), .A2(n2398), .ZN(n2672) );
  AND2_X1 U2485 ( .A1(n2415), .A2(n2397), .ZN(n2400) );
  AND2_X1 U2486 ( .A1(n2372), .A2(n2374), .ZN(n3992) );
  NAND2_X1 U2487 ( .A1(n2448), .A2(REG3_REG_2__SCAN_IN), .ZN(n2427) );
  INV_X1 U2488 ( .A(n3949), .ZN(n3627) );
  NAND2_X1 U2489 ( .A1(n3701), .A2(n3705), .ZN(n3648) );
  AND2_X1 U2490 ( .A1(n2238), .A2(n2237), .ZN(n3468) );
  INV_X1 U2491 ( .A(n4229), .ZN(n4203) );
  NAND4_X2 U2492 ( .A1(n2425), .A2(n2424), .A3(n2423), .A4(n2422), .ZN(n3956)
         );
  NAND2_X1 U2493 ( .A1(n2007), .A2(REG0_REG_0__SCAN_IN), .ZN(n2424) );
  NAND2_X1 U2494 ( .A1(n2789), .A2(n2788), .ZN(n2792) );
  OR2_X1 U2495 ( .A1(n2787), .A2(REG2_REG_1__SCAN_IN), .ZN(n2789) );
  OAI21_X1 U2496 ( .B1(n4493), .B2(n2802), .A(n2132), .ZN(n3969) );
  NAND2_X1 U2497 ( .A1(n4493), .A2(n2802), .ZN(n2132) );
  NAND2_X1 U2498 ( .A1(n3968), .A2(n3969), .ZN(n3967) );
  AND2_X1 U2499 ( .A1(n2815), .A2(n4529), .ZN(n2069) );
  NAND2_X1 U2500 ( .A1(n3167), .A2(REG1_REG_10__SCAN_IN), .ZN(n3289) );
  AOI21_X1 U2501 ( .B1(n3288), .B2(n2171), .A(n2170), .ZN(n2167) );
  INV_X1 U2502 ( .A(n3288), .ZN(n2168) );
  NAND2_X1 U2503 ( .A1(n3288), .A2(n3289), .ZN(n3291) );
  NAND2_X1 U2504 ( .A1(n3980), .A2(REG1_REG_12__SCAN_IN), .ZN(n3991) );
  AND2_X1 U2505 ( .A1(n4577), .A2(n2052), .ZN(n4597) );
  NAND2_X1 U2506 ( .A1(n4577), .A2(n4505), .ZN(n4598) );
  INV_X1 U2507 ( .A(n4591), .ZN(n2073) );
  AOI21_X1 U2508 ( .B1(n4592), .B2(n4593), .A(n4590), .ZN(n2074) );
  INV_X1 U2509 ( .A(n2072), .ZN(n2071) );
  AOI21_X1 U2510 ( .B1(n4595), .B2(ADDR_REG_18__SCAN_IN), .A(n4594), .ZN(n2072) );
  INV_X1 U2511 ( .A(n4586), .ZN(n4596) );
  AND2_X1 U2512 ( .A1(n2791), .A2(n3960), .ZN(n4584) );
  INV_X1 U2513 ( .A(n4618), .ZN(n4287) );
  INV_X1 U2514 ( .A(n4317), .ZN(n4608) );
  INV_X1 U2515 ( .A(IR_REG_29__SCAN_IN), .ZN(n2418) );
  INV_X1 U2516 ( .A(n4171), .ZN(n2090) );
  INV_X1 U2517 ( .A(n3914), .ZN(n2255) );
  NOR2_X1 U2518 ( .A1(n3861), .A2(n2257), .ZN(n2256) );
  AND2_X1 U2519 ( .A1(n3831), .A2(n2597), .ZN(n3910) );
  NAND2_X1 U2520 ( .A1(n2323), .A2(n2221), .ZN(n2220) );
  INV_X1 U2521 ( .A(IR_REG_24__SCAN_IN), .ZN(n2321) );
  INV_X1 U2522 ( .A(n3355), .ZN(n3358) );
  INV_X1 U2523 ( .A(n3722), .ZN(n2295) );
  AOI21_X1 U2524 ( .B1(n2669), .B2(IR_REG_31__SCAN_IN), .A(n2218), .ZN(n2217)
         );
  NAND2_X1 U2525 ( .A1(n2219), .A2(IR_REG_28__SCAN_IN), .ZN(n2218) );
  NAND2_X1 U2526 ( .A1(IR_REG_31__SCAN_IN), .A2(n2220), .ZN(n2219) );
  INV_X1 U2527 ( .A(IR_REG_28__SCAN_IN), .ZN(n3604) );
  INV_X1 U2528 ( .A(n2458), .ZN(n2081) );
  AND2_X1 U2529 ( .A1(n3899), .A2(n2632), .ZN(n2080) );
  AND2_X1 U2530 ( .A1(n3889), .A2(n2085), .ZN(n3896) );
  NOR2_X1 U2531 ( .A1(n4098), .A2(n2086), .ZN(n2085) );
  NAND2_X1 U2532 ( .A1(n2087), .A2(n4145), .ZN(n2086) );
  NAND2_X1 U2533 ( .A1(n4486), .A2(REG1_REG_11__SCAN_IN), .ZN(n3978) );
  NOR2_X1 U2534 ( .A1(n2170), .A2(n2171), .ZN(n2169) );
  AND2_X1 U2535 ( .A1(n3870), .A2(n4060), .ZN(n3914) );
  NOR2_X1 U2536 ( .A1(n2576), .A2(n2083), .ZN(n2082) );
  INV_X1 U2537 ( .A(n2567), .ZN(n2566) );
  NAND2_X1 U2538 ( .A1(n2538), .A2(n2258), .ZN(n2260) );
  NOR2_X1 U2539 ( .A1(n3904), .A2(n2259), .ZN(n2258) );
  NOR2_X1 U2540 ( .A1(n2533), .A2(n2532), .ZN(n2092) );
  INV_X1 U2541 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2525) );
  INV_X1 U2542 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2487) );
  NAND2_X1 U2543 ( .A1(n2479), .A2(REG3_REG_9__SCAN_IN), .ZN(n2488) );
  INV_X1 U2544 ( .A(n2481), .ZN(n2479) );
  AND2_X1 U2545 ( .A1(n2189), .A2(n2012), .ZN(n2184) );
  NOR2_X1 U2546 ( .A1(n2736), .A2(n4064), .ZN(n2228) );
  NOR2_X1 U2547 ( .A1(n4154), .A2(n4128), .ZN(n2224) );
  NOR2_X1 U2548 ( .A1(n4238), .A2(n4256), .ZN(n2236) );
  OAI21_X1 U2549 ( .B1(n2206), .B2(n2205), .A(n2035), .ZN(n2204) );
  INV_X1 U2550 ( .A(n2882), .ZN(n2660) );
  AND2_X1 U2551 ( .A1(n2898), .A2(n2864), .ZN(n2230) );
  INV_X1 U2552 ( .A(n2381), .ZN(n2393) );
  AND2_X1 U2553 ( .A1(n2359), .A2(n2358), .ZN(n2367) );
  NOR2_X1 U2554 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .ZN(n2320)
         );
  NOR2_X1 U2555 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2319)
         );
  OR2_X1 U2556 ( .A1(n3103), .A2(n2281), .ZN(n2280) );
  INV_X1 U2557 ( .A(n3100), .ZN(n2281) );
  NAND2_X1 U2558 ( .A1(n3472), .A2(n3470), .ZN(n3330) );
  AOI21_X1 U2559 ( .B1(n2032), .B2(n3351), .A(n2107), .ZN(n2106) );
  INV_X1 U2560 ( .A(n3742), .ZN(n2107) );
  OAI21_X1 U2561 ( .B1(n3046), .B2(n3432), .A(n2957), .ZN(n2958) );
  INV_X1 U2562 ( .A(n3000), .ZN(n2944) );
  NAND2_X1 U2563 ( .A1(n2308), .A2(n2301), .ZN(n3463) );
  NOR2_X1 U2564 ( .A1(n2100), .A2(n3419), .ZN(n2099) );
  INV_X1 U2565 ( .A(n2050), .ZN(n2100) );
  OR2_X1 U2566 ( .A1(n2511), .A2(n2505), .ZN(n2519) );
  NOR2_X1 U2567 ( .A1(n3376), .A2(n2122), .ZN(n2121) );
  INV_X1 U2568 ( .A(n3705), .ZN(n2122) );
  OR2_X1 U2569 ( .A1(n2488), .A2(n2487), .ZN(n2497) );
  NAND2_X1 U2570 ( .A1(n3330), .A2(n3469), .ZN(n3666) );
  NAND2_X1 U2571 ( .A1(n2449), .A2(REG3_REG_5__SCAN_IN), .ZN(n2458) );
  INV_X1 U2572 ( .A(n2451), .ZN(n2449) );
  AND2_X1 U2573 ( .A1(n3931), .A2(n4482), .ZN(n2882) );
  NAND2_X1 U2574 ( .A1(n2865), .A2(n4482), .ZN(n3936) );
  AND2_X1 U2575 ( .A1(n2545), .A2(n2544), .ZN(n4187) );
  NAND2_X1 U2576 ( .A1(n2799), .A2(n2798), .ZN(n3965) );
  INV_X1 U2577 ( .A(n2139), .ZN(n2136) );
  NAND2_X1 U2578 ( .A1(n2057), .A2(n2972), .ZN(n3064) );
  NAND2_X1 U2579 ( .A1(n2971), .A2(n4682), .ZN(n2972) );
  NAND2_X1 U2580 ( .A1(n2970), .A2(n2058), .ZN(n2057) );
  NAND2_X1 U2581 ( .A1(n4489), .A2(REG1_REG_7__SCAN_IN), .ZN(n2058) );
  INV_X1 U2582 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2171) );
  NAND2_X1 U2583 ( .A1(n4513), .A2(n4512), .ZN(n4514) );
  NAND2_X1 U2584 ( .A1(n2040), .A2(n2156), .ZN(n2154) );
  AOI21_X1 U2585 ( .B1(n2157), .B2(n2159), .A(n2040), .ZN(n2155) );
  OR2_X1 U2586 ( .A1(n4551), .A2(n2144), .ZN(n2143) );
  AOI21_X1 U2587 ( .B1(n2039), .B2(n4551), .A(n2142), .ZN(n2141) );
  NAND2_X1 U2588 ( .A1(n4552), .A2(n2039), .ZN(n2140) );
  NAND2_X1 U2589 ( .A1(n4569), .A2(n4518), .ZN(n4581) );
  NAND2_X1 U2590 ( .A1(n4581), .A2(n4582), .ZN(n4580) );
  AND2_X1 U2591 ( .A1(n3850), .A2(DATAI_27_), .ZN(n4032) );
  NAND2_X1 U2592 ( .A1(n2599), .A2(n3865), .ZN(n4075) );
  NAND2_X1 U2593 ( .A1(n2566), .A2(n2082), .ZN(n2589) );
  OR2_X1 U2594 ( .A1(n2547), .A2(n3639), .ZN(n2567) );
  NAND2_X1 U2595 ( .A1(n4212), .A2(n2201), .ZN(n2199) );
  NAND2_X1 U2596 ( .A1(n2092), .A2(REG3_REG_17__SCAN_IN), .ZN(n2557) );
  OR2_X1 U2597 ( .A1(n2526), .A2(n2525), .ZN(n2533) );
  INV_X1 U2598 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2532) );
  AND2_X1 U2599 ( .A1(n2232), .A2(n3421), .ZN(n2231) );
  NAND2_X1 U2600 ( .A1(n4295), .A2(n3817), .ZN(n3298) );
  AND2_X1 U2601 ( .A1(n3297), .A2(n3817), .ZN(n4302) );
  NAND2_X1 U2602 ( .A1(n2494), .A2(n3813), .ZN(n4295) );
  AND3_X1 U2603 ( .A1(n3072), .A2(n2230), .A3(n2229), .ZN(n3120) );
  AND2_X1 U2604 ( .A1(n3034), .A2(n2944), .ZN(n2229) );
  NAND2_X1 U2605 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2451) );
  NAND2_X1 U2606 ( .A1(n2703), .A2(n2702), .ZN(n2992) );
  OR2_X1 U2607 ( .A1(n3850), .A2(n2331), .ZN(n2333) );
  NOR2_X1 U2608 ( .A1(n3077), .A2(n3078), .ZN(n3076) );
  INV_X1 U2609 ( .A(n2892), .ZN(n2864) );
  INV_X1 U2610 ( .A(n3466), .ZN(n2898) );
  OR2_X1 U2611 ( .A1(n2752), .A2(n3835), .ZN(n4004) );
  NOR2_X1 U2612 ( .A1(n4004), .A2(n4005), .ZN(n4003) );
  NAND2_X1 U2613 ( .A1(n4082), .A2(n2228), .ZN(n4050) );
  AND2_X1 U2614 ( .A1(n4089), .A2(n4080), .ZN(n4082) );
  AND2_X1 U2615 ( .A1(n4162), .A2(n2223), .ZN(n4089) );
  AND2_X1 U2616 ( .A1(n2006), .A2(n3483), .ZN(n2223) );
  NAND2_X1 U2617 ( .A1(n4162), .A2(n2006), .ZN(n4346) );
  AND2_X1 U2618 ( .A1(n3850), .A2(DATAI_21_), .ZN(n4128) );
  AOI21_X1 U2619 ( .B1(n2203), .B2(n2031), .A(n2197), .ZN(n2196) );
  OR2_X1 U2620 ( .A1(n4190), .A2(n4184), .ZN(n2310) );
  INV_X1 U2621 ( .A(n3640), .ZN(n4172) );
  NAND2_X1 U2622 ( .A1(n2538), .A2(n3903), .ZN(n4164) );
  AND2_X1 U2623 ( .A1(n2552), .A2(n2551), .ZN(n4205) );
  NAND2_X1 U2624 ( .A1(n2247), .A2(n2246), .ZN(n4246) );
  AOI21_X1 U2625 ( .B1(n2248), .B2(n2251), .A(n4244), .ZN(n2246) );
  INV_X1 U2626 ( .A(n4276), .ZN(n4298) );
  INV_X1 U2627 ( .A(n4279), .ZN(n4306) );
  NOR2_X1 U2628 ( .A1(n4284), .A2(n2234), .ZN(n4237) );
  INV_X1 U2629 ( .A(n2236), .ZN(n2234) );
  OR2_X1 U2630 ( .A1(n3302), .A2(n2723), .ZN(n4284) );
  AND2_X1 U2631 ( .A1(n3207), .A2(n2232), .ZN(n4314) );
  NAND2_X1 U2632 ( .A1(n3207), .A2(n2009), .ZN(n4312) );
  NAND2_X1 U2633 ( .A1(n3207), .A2(n3249), .ZN(n3222) );
  AOI21_X1 U2634 ( .B1(n2267), .B2(n2265), .A(n2264), .ZN(n2263) );
  INV_X1 U2635 ( .A(n2267), .ZN(n2266) );
  INV_X1 U2636 ( .A(n3807), .ZN(n2265) );
  NAND2_X1 U2637 ( .A1(n4483), .A2(n2901), .ZN(n4279) );
  NOR2_X1 U2638 ( .A1(n3138), .A2(n3137), .ZN(n3156) );
  AND2_X1 U2639 ( .A1(n3156), .A2(n3184), .ZN(n3207) );
  NAND2_X1 U2640 ( .A1(n2213), .A2(n2216), .ZN(n3144) );
  OR2_X1 U2641 ( .A1(n3118), .A2(n3051), .ZN(n3138) );
  INV_X1 U2642 ( .A(n4668), .ZN(n4665) );
  NAND2_X1 U2643 ( .A1(n2230), .A2(n3034), .ZN(n3077) );
  NAND2_X1 U2644 ( .A1(n2898), .A2(n2864), .ZN(n3038) );
  INV_X1 U2645 ( .A(n4661), .ZN(n4653) );
  NAND2_X1 U2646 ( .A1(n2901), .A2(n2739), .ZN(n4661) );
  AND2_X1 U2647 ( .A1(n2862), .A2(n2691), .ZN(n2887) );
  NAND2_X1 U2648 ( .A1(n2669), .A2(IR_REG_31__SCAN_IN), .ZN(n2120) );
  NAND2_X1 U2649 ( .A1(n2272), .A2(IR_REG_31__SCAN_IN), .ZN(n2690) );
  NAND2_X1 U2650 ( .A1(n2269), .A2(n2273), .ZN(n2689) );
  NAND2_X1 U2651 ( .A1(n2400), .A2(n2274), .ZN(n2272) );
  XNOR2_X1 U2652 ( .A(n2399), .B(n2276), .ZN(n2692) );
  INV_X1 U2653 ( .A(IR_REG_17__SCAN_IN), .ZN(n2389) );
  OR2_X1 U2654 ( .A1(n2374), .A2(IR_REG_14__SCAN_IN), .ZN(n2375) );
  NOR2_X1 U2655 ( .A1(n2367), .A2(n2763), .ZN(n2360) );
  NOR2_X1 U2656 ( .A1(n2381), .A2(IR_REG_9__SCAN_IN), .ZN(n2359) );
  INV_X1 U2657 ( .A(IR_REG_7__SCAN_IN), .ZN(n2352) );
  NAND2_X1 U2658 ( .A1(n2282), .A2(n3100), .ZN(n3102) );
  AND2_X1 U2659 ( .A1(n2641), .A2(n2640), .ZN(n4025) );
  OR2_X1 U2660 ( .A1(n3456), .A2(n2643), .ZN(n2641) );
  INV_X1 U2661 ( .A(n2115), .ZN(n2111) );
  NAND2_X1 U2662 ( .A1(n3430), .A2(n2287), .ZN(n2114) );
  OR2_X1 U2663 ( .A1(n3695), .A2(n2643), .ZN(n2606) );
  NAND2_X1 U2664 ( .A1(n2131), .A2(n2130), .ZN(n3624) );
  AND2_X1 U2665 ( .A1(n2123), .A2(n2131), .ZN(n3623) );
  INV_X1 U2666 ( .A(n2127), .ZN(n2123) );
  OAI21_X1 U2667 ( .B1(n3658), .B2(n2288), .A(n2034), .ZN(n2309) );
  NAND2_X1 U2668 ( .A1(n2287), .A2(n2117), .ZN(n2285) );
  NOR2_X1 U2669 ( .A1(n3430), .A2(n2116), .ZN(n2286) );
  AND4_X1 U2670 ( .A1(n2468), .A2(n2467), .A3(n2466), .A4(n2465), .ZN(n3185)
         );
  AND4_X1 U2671 ( .A1(n2502), .A2(n2501), .A3(n2500), .A4(n2499), .ZN(n3626)
         );
  NAND2_X1 U2672 ( .A1(n3310), .A2(n3309), .ZN(n2101) );
  NAND2_X1 U2673 ( .A1(n3312), .A2(n3311), .ZN(n2102) );
  NAND2_X1 U2674 ( .A1(n2955), .A2(n2954), .ZN(n3007) );
  CLKBUF_X1 U2675 ( .A(n3690), .Z(n3691) );
  NAND2_X1 U2676 ( .A1(n2920), .A2(n2921), .ZN(n2941) );
  AND4_X1 U2677 ( .A1(n2478), .A2(n2477), .A3(n2476), .A4(n2475), .ZN(n3245)
         );
  INV_X1 U2678 ( .A(n2305), .ZN(n2129) );
  NAND3_X1 U2679 ( .A1(n2096), .A2(n2095), .A3(n2097), .ZN(n3715) );
  INV_X1 U2680 ( .A(n2099), .ZN(n2097) );
  AND2_X1 U2681 ( .A1(n2595), .A2(n2594), .ZN(n4115) );
  NAND2_X1 U2682 ( .A1(n2296), .A2(n3375), .ZN(n3721) );
  INV_X1 U2683 ( .A(n3948), .ZN(n4297) );
  CLKBUF_X1 U2684 ( .A(n3729), .Z(n3730) );
  INV_X1 U2685 ( .A(n3776), .ZN(n3750) );
  INV_X1 U2686 ( .A(n3777), .ZN(n3749) );
  OAI21_X1 U2687 ( .B1(n2889), .B2(n4279), .A(n4287), .ZN(n3754) );
  INV_X1 U2688 ( .A(n3754), .ZN(n3775) );
  INV_X1 U2689 ( .A(n2093), .ZN(n4052) );
  AND4_X1 U2690 ( .A1(n2524), .A2(n2523), .A3(n2522), .A4(n2521), .ZN(n4228)
         );
  AND3_X1 U2691 ( .A1(n2537), .A2(n2536), .A3(n2535), .ZN(n4229) );
  NAND2_X1 U2692 ( .A1(n2886), .A2(n4479), .ZN(n3777) );
  OAI21_X1 U2693 ( .B1(n2076), .B2(n2739), .A(n2075), .ZN(n3934) );
  NAND2_X1 U2694 ( .A1(n3933), .A2(n2739), .ZN(n2075) );
  AOI21_X1 U2695 ( .B1(n3932), .B2(n3931), .A(n2077), .ZN(n2076) );
  INV_X1 U2696 ( .A(n4025), .ZN(n3944) );
  NAND2_X1 U2697 ( .A1(n2631), .A2(n2630), .ZN(n4047) );
  OR2_X1 U2698 ( .A1(n4036), .A2(n2643), .ZN(n2631) );
  OAI21_X1 U2699 ( .B1(n2093), .B2(n2643), .A(n2622), .ZN(n3945) );
  OR2_X1 U2700 ( .A1(n3659), .A2(n2643), .ZN(n2614) );
  INV_X1 U2701 ( .A(n4115), .ZN(n2896) );
  NAND2_X1 U2702 ( .A1(n2573), .A2(n2572), .ZN(n4129) );
  INV_X1 U2703 ( .A(n4187), .ZN(n3946) );
  INV_X1 U2704 ( .A(n4205), .ZN(n4173) );
  INV_X1 U2705 ( .A(n4217), .ZN(n4185) );
  INV_X1 U2706 ( .A(n3185), .ZN(n3951) );
  NOR2_X1 U2707 ( .A1(n2436), .A2(n2435), .ZN(n2437) );
  XNOR2_X1 U2708 ( .A(n2787), .B(REG1_REG_1__SCAN_IN), .ZN(n2797) );
  NAND2_X1 U2709 ( .A1(n2804), .A2(n2803), .ZN(n3968) );
  XNOR2_X1 U2710 ( .A(n2818), .B(n2331), .ZN(n2817) );
  NAND2_X1 U2711 ( .A1(n2343), .A2(n2345), .ZN(n2835) );
  AOI21_X1 U2712 ( .B1(n4527), .B2(REG2_REG_4__SCAN_IN), .A(n2136), .ZN(n2830)
         );
  XNOR2_X1 U2713 ( .A(n2063), .B(n2062), .ZN(n2855) );
  AOI22_X1 U2714 ( .A1(n2855), .A2(REG2_REG_6__SCAN_IN), .B1(n4490), .B2(n2063), .ZN(n2857) );
  XNOR2_X1 U2715 ( .A(n3064), .B(n3055), .ZN(n2973) );
  NAND2_X1 U2716 ( .A1(n2973), .A2(REG1_REG_8__SCAN_IN), .ZN(n3062) );
  NAND2_X1 U2717 ( .A1(n3062), .A2(n2162), .ZN(n3066) );
  NAND2_X1 U2718 ( .A1(n2163), .A2(n3055), .ZN(n2162) );
  INV_X1 U2719 ( .A(n3064), .ZN(n2163) );
  NAND2_X1 U2720 ( .A1(n3066), .A2(n3065), .ZN(n3166) );
  NAND2_X1 U2721 ( .A1(n2146), .A2(n2147), .ZN(n3162) );
  NAND2_X1 U2722 ( .A1(n3056), .A2(REG2_REG_8__SCAN_IN), .ZN(n2149) );
  XNOR2_X1 U2723 ( .A(n2152), .B(n3287), .ZN(n3279) );
  OAI21_X1 U2724 ( .B1(n3986), .B2(n3985), .A(n2161), .ZN(n4546) );
  AND2_X1 U2725 ( .A1(n3991), .A2(n3990), .ZN(n4540) );
  XNOR2_X1 U2726 ( .A(n4496), .B(n4512), .ZN(n3987) );
  NOR2_X1 U2727 ( .A1(n4555), .A2(n4554), .ZN(n4553) );
  AND2_X1 U2728 ( .A1(n4515), .A2(n4514), .ZN(n4555) );
  NOR2_X1 U2729 ( .A1(n4552), .A2(n4551), .ZN(n4550) );
  AND2_X1 U2730 ( .A1(n2791), .A2(n2790), .ZN(n4586) );
  INV_X1 U2731 ( .A(n4522), .ZN(n2066) );
  OR2_X1 U2732 ( .A1(n2634), .A2(n2633), .ZN(n4012) );
  NAND2_X1 U2733 ( .A1(n2185), .A2(n2189), .ZN(n4040) );
  OR2_X1 U2734 ( .A1(n4073), .A2(n2192), .ZN(n2185) );
  NAND2_X1 U2735 ( .A1(n4162), .A2(n4147), .ZN(n4355) );
  NAND2_X1 U2736 ( .A1(n2207), .A2(n2206), .ZN(n4266) );
  OAI21_X1 U2737 ( .B1(n3201), .B2(n2717), .A(n2716), .ZN(n3220) );
  NAND2_X1 U2738 ( .A1(n2708), .A2(n2707), .ZN(n3044) );
  AND2_X1 U2739 ( .A1(n4289), .A2(n2982), .ZN(n4620) );
  XNOR2_X1 U2740 ( .A(n4003), .B(n4000), .ZN(n4399) );
  NAND2_X1 U2741 ( .A1(n2193), .A2(n2010), .ZN(n4057) );
  NAND2_X1 U2742 ( .A1(n4073), .A2(n2735), .ZN(n2193) );
  NAND2_X1 U2743 ( .A1(n4212), .A2(n2728), .ZN(n4198) );
  INV_X1 U2744 ( .A(n4476), .ZN(n4455) );
  NAND2_X1 U2745 ( .A1(n2764), .A2(IR_REG_31__SCAN_IN), .ZN(n2420) );
  NAND2_X1 U2746 ( .A1(n2655), .A2(IR_REG_31__SCAN_IN), .ZN(n2417) );
  AND2_X1 U2747 ( .A1(n2670), .A2(n2013), .ZN(n4481) );
  NAND2_X1 U2748 ( .A1(n2119), .A2(n2118), .ZN(n2670) );
  NAND2_X1 U2749 ( .A1(IR_REG_31__SCAN_IN), .A2(n2323), .ZN(n2118) );
  NAND2_X1 U2750 ( .A1(n2120), .A2(IR_REG_25__SCAN_IN), .ZN(n2119) );
  AOI21_X1 U2751 ( .B1(n2273), .B2(n2763), .A(n2763), .ZN(n2270) );
  INV_X1 U2752 ( .A(n2692), .ZN(n4482) );
  XNOR2_X1 U2753 ( .A(n2337), .B(IR_REG_4__SCAN_IN), .ZN(n4529) );
  NOR2_X1 U2754 ( .A1(n2763), .A2(n2328), .ZN(n2056) );
  OAI21_X1 U2755 ( .B1(n3167), .B2(n2168), .A(n2167), .ZN(n3979) );
  AOI211_X1 U2756 ( .C1(n4599), .C2(n4598), .A(n4597), .B(n4596), .ZN(n4600)
         );
  OAI21_X1 U2757 ( .B1(n3461), .B2(n4242), .A(n2065), .ZN(n2064) );
  AOI21_X1 U2758 ( .B1(n3460), .B2(n4608), .A(n3459), .ZN(n2065) );
  OR2_X1 U2759 ( .A1(n3454), .A2(n4395), .ZN(n2756) );
  NAND2_X1 U2760 ( .A1(n4681), .A2(n2638), .ZN(n2068) );
  OR2_X1 U2761 ( .A1(n3454), .A2(n4476), .ZN(n2753) );
  AND2_X1 U2762 ( .A1(n4077), .A2(n4064), .ZN(n2005) );
  INV_X1 U2763 ( .A(n4485), .ZN(n2157) );
  AND2_X1 U2764 ( .A1(n4112), .A2(n2224), .ZN(n2006) );
  INV_X1 U2765 ( .A(n4112), .ZN(n4120) );
  INV_X1 U2766 ( .A(IR_REG_31__SCAN_IN), .ZN(n2356) );
  AND2_X1 U2767 ( .A1(n2245), .A2(n2421), .ZN(n2007) );
  AND2_X1 U2768 ( .A1(n3891), .A2(n4269), .ZN(n2008) );
  AND2_X1 U2769 ( .A1(n3249), .A2(n3631), .ZN(n2009) );
  OR2_X1 U2770 ( .A1(n4065), .A2(n2734), .ZN(n2010) );
  NAND2_X1 U2771 ( .A1(n4185), .A2(n4202), .ZN(n2011) );
  OR2_X1 U2772 ( .A1(n4067), .A2(n4051), .ZN(n2012) );
  OR2_X1 U2773 ( .A1(n2669), .A2(IR_REG_25__SCAN_IN), .ZN(n2013) );
  INV_X1 U2774 ( .A(n2730), .ZN(n2203) );
  NAND2_X1 U2775 ( .A1(n2614), .A2(n2613), .ZN(n4077) );
  NAND2_X1 U2776 ( .A1(n4162), .A2(n2224), .ZN(n2225) );
  AND2_X1 U2777 ( .A1(n2050), .A2(n3311), .ZN(n2014) );
  AND2_X1 U2778 ( .A1(n2942), .A2(n2943), .ZN(n2015) );
  AND2_X1 U2779 ( .A1(n2115), .A2(n2288), .ZN(n2016) );
  AND2_X1 U2780 ( .A1(n2050), .A2(n3309), .ZN(n2017) );
  NOR2_X1 U2781 ( .A1(n4543), .A2(REG2_REG_12__SCAN_IN), .ZN(n2018) );
  OR2_X1 U2782 ( .A1(n4284), .A2(n2235), .ZN(n2019) );
  INV_X1 U2783 ( .A(n3655), .ZN(n2117) );
  NAND2_X1 U2784 ( .A1(n2160), .A2(n4485), .ZN(n2156) );
  INV_X2 U2785 ( .A(n4673), .ZN(n4675) );
  NAND2_X1 U2786 ( .A1(n2199), .A2(n2200), .ZN(n4137) );
  NAND2_X1 U2787 ( .A1(n3173), .A2(n3172), .ZN(n2020) );
  AND2_X1 U2788 ( .A1(n4082), .A2(n3661), .ZN(n2021) );
  AND2_X1 U2789 ( .A1(n2295), .A2(n3375), .ZN(n2022) );
  NAND2_X1 U2790 ( .A1(n2138), .A2(n2137), .ZN(n2063) );
  NAND4_X1 U2791 ( .A1(n2327), .A2(n2320), .A3(n2319), .A4(n2328), .ZN(n2413)
         );
  OR2_X1 U2792 ( .A1(n3268), .A2(n3267), .ZN(n2023) );
  AND3_X1 U2793 ( .A1(n3428), .A2(n4478), .A3(REG3_REG_1__SCAN_IN), .ZN(n2024)
         );
  NAND2_X1 U2794 ( .A1(n2333), .A2(n2332), .ZN(n3078) );
  AND2_X1 U2795 ( .A1(n4217), .A2(n3339), .ZN(n2025) );
  OAI21_X1 U2796 ( .B1(n3648), .B2(n2291), .A(n2292), .ZN(n3692) );
  AND3_X1 U2797 ( .A1(n2445), .A2(n2444), .A3(n2443), .ZN(n2026) );
  AND2_X1 U2798 ( .A1(n3817), .A2(n2250), .ZN(n2027) );
  OR2_X1 U2799 ( .A1(n4077), .A2(n4064), .ZN(n2028) );
  AND2_X1 U2800 ( .A1(n2717), .A2(n2716), .ZN(n2029) );
  INV_X1 U2801 ( .A(n2192), .ZN(n2191) );
  NAND2_X1 U2802 ( .A1(n2010), .A2(n2028), .ZN(n2192) );
  INV_X1 U2803 ( .A(n3917), .ZN(n2254) );
  NOR2_X1 U2804 ( .A1(n3261), .A2(n3260), .ZN(n2030) );
  OR2_X1 U2805 ( .A1(n2729), .A2(n2198), .ZN(n2031) );
  OR2_X1 U2806 ( .A1(n3745), .A2(n2108), .ZN(n2032) );
  NAND2_X1 U2807 ( .A1(n2207), .A2(n2208), .ZN(n3294) );
  INV_X1 U2808 ( .A(n3381), .ZN(n2294) );
  AND2_X1 U2809 ( .A1(n2471), .A2(REG3_REG_6__SCAN_IN), .ZN(n2033) );
  AND2_X1 U2810 ( .A1(n2286), .A2(n2285), .ZN(n2034) );
  NAND2_X1 U2811 ( .A1(n2723), .A2(n4249), .ZN(n2035) );
  INV_X1 U2812 ( .A(n2202), .ZN(n2201) );
  NAND2_X1 U2813 ( .A1(n2011), .A2(n2728), .ZN(n2202) );
  INV_X1 U2814 ( .A(IR_REG_25__SCAN_IN), .ZN(n2323) );
  INV_X1 U2815 ( .A(IR_REG_23__SCAN_IN), .ZN(n3507) );
  AND2_X1 U2816 ( .A1(n2283), .A2(n2020), .ZN(n2036) );
  NOR2_X1 U2817 ( .A1(n4302), .A2(n2719), .ZN(n2037) );
  AND2_X1 U2818 ( .A1(n2724), .A2(n2210), .ZN(n2038) );
  INV_X1 U2819 ( .A(IR_REG_26__SCAN_IN), .ZN(n2221) );
  XNOR2_X1 U2820 ( .A(n2673), .B(IR_REG_24__SCAN_IN), .ZN(n2688) );
  AND2_X1 U2821 ( .A1(n3905), .A2(n3903), .ZN(n4211) );
  NAND2_X1 U2822 ( .A1(n3984), .A2(n4485), .ZN(n2161) );
  NOR2_X1 U2823 ( .A1(n4501), .A2(n4638), .ZN(n2039) );
  OR2_X1 U2824 ( .A1(n2018), .A2(n2158), .ZN(n2040) );
  AND2_X1 U2825 ( .A1(n3850), .A2(DATAI_20_), .ZN(n4154) );
  INV_X1 U2826 ( .A(n3903), .ZN(n2259) );
  AND2_X1 U2827 ( .A1(n2102), .A2(n2101), .ZN(n3418) );
  INV_X1 U2828 ( .A(IR_REG_10__SCAN_IN), .ZN(n2358) );
  INV_X1 U2829 ( .A(n2617), .ZN(n2643) );
  AND2_X1 U2830 ( .A1(n3012), .A2(n3011), .ZN(n2041) );
  INV_X1 U2831 ( .A(IR_REG_22__SCAN_IN), .ZN(n2276) );
  AND4_X1 U2832 ( .A1(n3895), .A2(n3894), .A3(n4248), .A4(n3893), .ZN(n2042)
         );
  OR2_X1 U2833 ( .A1(n4284), .A2(n4256), .ZN(n2043) );
  AND2_X1 U2834 ( .A1(n2131), .A2(n2129), .ZN(n3262) );
  INV_X1 U2835 ( .A(n3865), .ZN(n2257) );
  INV_X1 U2836 ( .A(n3760), .ZN(n2116) );
  INV_X1 U2837 ( .A(n4543), .ZN(n2159) );
  AND2_X1 U2838 ( .A1(n2282), .A2(n2279), .ZN(n2044) );
  NAND2_X1 U2839 ( .A1(n4488), .A2(REG2_REG_9__SCAN_IN), .ZN(n2045) );
  INV_X1 U2840 ( .A(n2288), .ZN(n2287) );
  NAND2_X1 U2841 ( .A1(n3759), .A2(n2289), .ZN(n2288) );
  NAND2_X1 U2842 ( .A1(n4558), .A2(REG1_REG_15__SCAN_IN), .ZN(n2046) );
  AND2_X1 U2843 ( .A1(n2349), .A2(n2348), .ZN(n4489) );
  AND2_X1 U2844 ( .A1(n2896), .A2(n4099), .ZN(n2047) );
  INV_X1 U2845 ( .A(n2160), .ZN(n2158) );
  INV_X1 U2846 ( .A(n3483), .ZN(n4099) );
  AND2_X1 U2847 ( .A1(n2082), .A2(REG3_REG_23__SCAN_IN), .ZN(n2048) );
  INV_X1 U2848 ( .A(n4100), .ZN(n4131) );
  NAND2_X1 U2849 ( .A1(n2582), .A2(n2581), .ZN(n4100) );
  NAND2_X1 U2850 ( .A1(n3992), .A2(REG1_REG_13__SCAN_IN), .ZN(n2049) );
  INV_X1 U2851 ( .A(REG3_REG_20__SCAN_IN), .ZN(n2083) );
  INV_X1 U2852 ( .A(REG3_REG_23__SCAN_IN), .ZN(n2084) );
  INV_X1 U2853 ( .A(n4684), .ZN(n4681) );
  NAND2_X1 U2854 ( .A1(n3850), .A2(DATAI_22_), .ZN(n4112) );
  XNOR2_X1 U2855 ( .A(n2380), .B(n2379), .ZN(n4638) );
  INV_X1 U2856 ( .A(n4064), .ZN(n3661) );
  NAND2_X1 U2857 ( .A1(n3320), .A2(n3319), .ZN(n2050) );
  OR2_X1 U2858 ( .A1(n4675), .A2(REG0_REG_28__SCAN_IN), .ZN(n2051) );
  NOR2_X1 U2859 ( .A1(n4599), .A2(n4504), .ZN(n2052) );
  AND2_X1 U2860 ( .A1(n2149), .A2(n2153), .ZN(n2053) );
  XNOR2_X1 U2861 ( .A(n2346), .B(IR_REG_6__SCAN_IN), .ZN(n4490) );
  INV_X1 U2862 ( .A(n4490), .ZN(n2062) );
  AND2_X1 U2863 ( .A1(n4633), .A2(REG1_REG_18__SCAN_IN), .ZN(n2054) );
  INV_X1 U2864 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2135) );
  NAND2_X1 U2865 ( .A1(n2055), .A2(n2651), .ZN(n4281) );
  NAND2_X1 U2866 ( .A1(n3931), .A2(n4483), .ZN(n2055) );
  OAI211_X2 U2867 ( .C1(n2410), .C2(n2409), .A(n2408), .B(n2407), .ZN(n2739)
         );
  INV_X1 U2868 ( .A(n3931), .ZN(n2693) );
  AOI21_X1 U2869 ( .B1(n2067), .B2(n4281), .A(n2751), .ZN(n3457) );
  INV_X1 U2870 ( .A(n4281), .ZN(n4309) );
  NAND2_X1 U2871 ( .A1(n2061), .A2(n2059), .ZN(U3259) );
  INV_X1 U2872 ( .A(n2060), .ZN(n2059) );
  NAND2_X1 U2873 ( .A1(n2070), .A2(n4584), .ZN(n2061) );
  NOR2_X1 U2874 ( .A1(n2857), .A2(n2856), .ZN(n2967) );
  OAI21_X2 U2875 ( .B1(n3877), .B2(n3784), .A(n3788), .ZN(n3032) );
  OR2_X1 U2876 ( .A1(n3458), .A2(n2064), .ZN(U3262) );
  OAI21_X2 U2877 ( .B1(n3203), .B2(n3814), .A(n3811), .ZN(n3216) );
  XNOR2_X1 U2878 ( .A(n2748), .B(n3900), .ZN(n2067) );
  NAND2_X2 U2879 ( .A1(n2437), .A2(n2438), .ZN(n3737) );
  OAI21_X1 U2880 ( .B1(n2755), .B2(n4673), .A(n2051), .ZN(n2754) );
  OAI21_X1 U2881 ( .B1(n2755), .B2(n4681), .A(n2068), .ZN(n2757) );
  OAI21_X1 U2882 ( .B1(n2599), .B2(n2255), .A(n2252), .ZN(n2623) );
  XNOR2_X2 U2883 ( .A(n2815), .B(n2821), .ZN(n4525) );
  XNOR2_X1 U2884 ( .A(n2172), .B(n4519), .ZN(n2070) );
  NAND3_X1 U2885 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .A3(
        IR_REG_1__SCAN_IN), .ZN(n2183) );
  XNOR2_X2 U2886 ( .A(n4511), .B(n4512), .ZN(n3993) );
  NAND2_X1 U2887 ( .A1(n2566), .A2(n2048), .ZN(n2600) );
  NAND4_X1 U2888 ( .A1(n3887), .A2(n4231), .A3(n3888), .A4(n4211), .ZN(n2091)
         );
  NAND2_X1 U2889 ( .A1(n2941), .A2(n2015), .ZN(n2955) );
  XNOR2_X1 U2890 ( .A(n2951), .B(n2952), .ZN(n2942) );
  NAND2_X1 U2891 ( .A1(n3731), .A2(n2919), .ZN(n2920) );
  AOI22_X2 U2892 ( .A1(n3715), .A2(n3322), .B1(n2094), .B2(n3712), .ZN(n3472)
         );
  NAND3_X1 U2893 ( .A1(n2096), .A2(n2095), .A3(n2098), .ZN(n2094) );
  NAND2_X1 U2894 ( .A1(n3310), .A2(n2017), .ZN(n2095) );
  NAND2_X1 U2895 ( .A1(n3312), .A2(n2014), .ZN(n2096) );
  NAND2_X1 U2896 ( .A1(n3330), .A2(n2106), .ZN(n2105) );
  OAI21_X1 U2897 ( .B1(n3330), .B2(n3350), .A(n2106), .ZN(n3637) );
  AOI21_X1 U2898 ( .B1(n2106), .B2(n3350), .A(n2104), .ZN(n2103) );
  NAND2_X1 U2899 ( .A1(n3658), .A2(n3655), .ZN(n2290) );
  OAI211_X1 U2900 ( .C1(n3658), .C2(n2114), .A(n2112), .B(n2109), .ZN(n3413)
         );
  NAND2_X1 U2901 ( .A1(n3658), .A2(n2110), .ZN(n2109) );
  NOR2_X1 U2902 ( .A1(n2111), .A2(n3430), .ZN(n2110) );
  OAI21_X1 U2903 ( .B1(n2016), .B2(n3430), .A(n2113), .ZN(n2112) );
  NAND2_X1 U2904 ( .A1(n3430), .A2(n2115), .ZN(n2113) );
  NAND2_X1 U2905 ( .A1(n3242), .A2(n2125), .ZN(n2124) );
  INV_X1 U2906 ( .A(n2138), .ZN(n2828) );
  NAND2_X1 U2907 ( .A1(n2822), .A2(n4529), .ZN(n2139) );
  XNOR2_X1 U2908 ( .A(n3984), .B(n4485), .ZN(n3986) );
  OR2_X1 U2909 ( .A1(n3992), .A2(REG2_REG_13__SCAN_IN), .ZN(n2160) );
  NAND2_X2 U2910 ( .A1(n3166), .A2(n2298), .ZN(n3286) );
  INV_X1 U2911 ( .A(n2165), .ZN(n2164) );
  OAI21_X1 U2912 ( .B1(n3980), .B2(n2175), .A(n2174), .ZN(n2176) );
  INV_X1 U2913 ( .A(n3990), .ZN(n2175) );
  INV_X1 U2914 ( .A(n2176), .ZN(n4538) );
  INV_X1 U2915 ( .A(n2179), .ZN(n4517) );
  INV_X1 U2916 ( .A(IR_REG_1__SCAN_IN), .ZN(n2182) );
  XNOR2_X2 U2917 ( .A(n2850), .B(n4490), .ZN(n2852) );
  XNOR2_X2 U2918 ( .A(n2812), .B(n2331), .ZN(n2811) );
  NAND2_X1 U2919 ( .A1(n4073), .A2(n2184), .ZN(n2188) );
  NAND3_X1 U2920 ( .A1(n2189), .A2(n2192), .A3(n2012), .ZN(n2187) );
  NAND2_X1 U2921 ( .A1(n4212), .A2(n2195), .ZN(n2194) );
  NAND2_X1 U2922 ( .A1(n2194), .A2(n2196), .ZN(n4125) );
  AOI21_X1 U2923 ( .B1(n3201), .B2(n2038), .A(n2204), .ZN(n4245) );
  NAND3_X1 U2924 ( .A1(n2213), .A2(n2710), .A3(n2216), .ZN(n3143) );
  NAND2_X1 U2925 ( .A1(n2222), .A2(n2703), .ZN(n2994) );
  INV_X1 U2926 ( .A(n2225), .ZN(n4119) );
  NAND2_X1 U2927 ( .A1(n3207), .A2(n2231), .ZN(n3302) );
  INV_X1 U2928 ( .A(n2233), .ZN(n4190) );
  NAND2_X1 U2929 ( .A1(n2421), .A2(REG0_REG_1__SCAN_IN), .ZN(n2244) );
  NAND2_X1 U2930 ( .A1(n2242), .A2(n2245), .ZN(n2237) );
  AOI21_X1 U2931 ( .B1(n2241), .B2(n2421), .A(n2024), .ZN(n2238) );
  AND2_X1 U2932 ( .A1(n3428), .A2(n4478), .ZN(n2448) );
  INV_X1 U2933 ( .A(n2239), .ZN(n2431) );
  NAND2_X1 U2934 ( .A1(n2421), .A2(n3428), .ZN(n2239) );
  NAND2_X1 U2935 ( .A1(n2245), .A2(n4478), .ZN(n2240) );
  AND2_X1 U2936 ( .A1(n3428), .A2(REG2_REG_1__SCAN_IN), .ZN(n2241) );
  NAND2_X1 U2937 ( .A1(n2244), .A2(n2243), .ZN(n2242) );
  NAND2_X1 U2938 ( .A1(n4478), .A2(REG1_REG_1__SCAN_IN), .ZN(n2243) );
  XNOR2_X2 U2939 ( .A(n2417), .B(IR_REG_29__SCAN_IN), .ZN(n4478) );
  INV_X1 U2940 ( .A(n3428), .ZN(n2245) );
  OAI21_X1 U2941 ( .B1(n2494), .B2(n2251), .A(n2248), .ZN(n4247) );
  NAND2_X1 U2942 ( .A1(n2494), .A2(n2248), .ZN(n2247) );
  OAI21_X2 U2943 ( .B1(n2991), .B2(n2447), .A(n3798), .ZN(n3112) );
  NAND2_X1 U2944 ( .A1(n2260), .A2(n3829), .ZN(n2575) );
  INV_X1 U2945 ( .A(n2260), .ZN(n2561) );
  NAND2_X1 U2946 ( .A1(n4019), .A2(n3842), .ZN(n2261) );
  NAND2_X1 U2947 ( .A1(n2261), .A2(n2262), .ZN(n2642) );
  AOI21_X1 U2948 ( .B1(n4029), .B2(n3842), .A(n3837), .ZN(n2262) );
  NAND2_X1 U2949 ( .A1(n4021), .A2(n3842), .ZN(n2748) );
  OAI21_X1 U2950 ( .B1(n3132), .B2(n2469), .A(n3807), .ZN(n3151) );
  AOI21_X1 U2951 ( .B1(n2469), .B2(n3807), .A(n2268), .ZN(n2267) );
  NAND2_X2 U2952 ( .A1(n3785), .A2(n3788), .ZN(n3877) );
  NAND2_X1 U2953 ( .A1(n2400), .A2(n2273), .ZN(n2271) );
  NAND2_X1 U2954 ( .A1(n2271), .A2(n2270), .ZN(n2673) );
  NAND2_X1 U2955 ( .A1(n2280), .A2(n2020), .ZN(n2277) );
  NAND2_X1 U2956 ( .A1(n3012), .A2(n2036), .ZN(n2278) );
  INV_X1 U2957 ( .A(n2280), .ZN(n2279) );
  NAND2_X1 U2958 ( .A1(n3012), .A2(n2283), .ZN(n2282) );
  NOR2_X1 U2959 ( .A1(n2284), .A2(n3101), .ZN(n2283) );
  INV_X1 U2960 ( .A(n3011), .ZN(n2284) );
  AND2_X1 U2961 ( .A1(n2290), .A2(n2289), .ZN(n3758) );
  INV_X1 U2962 ( .A(n3376), .ZN(n2297) );
  AOI21_X1 U2963 ( .B1(n4005), .B2(n4004), .A(n4003), .ZN(n4400) );
  NAND2_X1 U2964 ( .A1(n2763), .A2(n2328), .ZN(n2329) );
  NAND2_X2 U2965 ( .A1(n2814), .A2(n2813), .ZN(n2815) );
  NAND2_X1 U2966 ( .A1(n2787), .A2(REG2_REG_1__SCAN_IN), .ZN(n2788) );
  INV_X4 U2967 ( .A(n2932), .ZN(n3953) );
  OR2_X1 U2968 ( .A1(n2400), .A2(n2763), .ZN(n2401) );
  INV_X1 U2969 ( .A(n4478), .ZN(n2421) );
  CLKBUF_X1 U2970 ( .A(n3308), .Z(n3271) );
  NAND2_X1 U2971 ( .A1(n2951), .A2(n2953), .ZN(n2954) );
  INV_X1 U2972 ( .A(n3468), .ZN(n2868) );
  AND2_X1 U2973 ( .A1(n2676), .A2(n3415), .ZN(n2694) );
  OR2_X1 U2974 ( .A1(n3165), .A2(n3576), .ZN(n2298) );
  AND2_X1 U2975 ( .A1(n2352), .A2(n2351), .ZN(n2299) );
  AND3_X1 U2976 ( .A1(n2221), .A2(n2661), .A3(n2323), .ZN(n2300) );
  OR2_X1 U2977 ( .A1(n2862), .A2(n2871), .ZN(n2301) );
  OR2_X1 U2978 ( .A1(n3936), .A2(n2981), .ZN(n2302) );
  AND2_X1 U2979 ( .A1(n2887), .A2(n2922), .ZN(n2303) );
  INV_X1 U2980 ( .A(n4029), .ZN(n2632) );
  AND2_X1 U2981 ( .A1(n2606), .A2(n2605), .ZN(n4102) );
  INV_X1 U2982 ( .A(n4102), .ZN(n4065) );
  OR2_X1 U2983 ( .A1(n3945), .A2(n2736), .ZN(n2304) );
  NOR2_X1 U2984 ( .A1(n3240), .A2(n3239), .ZN(n2305) );
  AND2_X1 U2985 ( .A1(n3774), .A2(n3672), .ZN(n2306) );
  AND2_X2 U2986 ( .A1(n2980), .A2(n4287), .ZN(n4623) );
  NAND2_X1 U2987 ( .A1(n2327), .A2(n2328), .ZN(n2307) );
  INV_X1 U2988 ( .A(n4080), .ZN(n2734) );
  INV_X1 U2989 ( .A(n2688), .ZN(n2696) );
  XNOR2_X1 U2990 ( .A(n2935), .B(n3433), .ZN(n2951) );
  AND2_X1 U2991 ( .A1(n2363), .A2(n2364), .ZN(n4486) );
  XNOR2_X1 U2992 ( .A(n2357), .B(IR_REG_10__SCAN_IN), .ZN(n4487) );
  OR2_X1 U2993 ( .A1(n2562), .A2(n4166), .ZN(n3904) );
  AND2_X1 U2994 ( .A1(n3388), .A2(n3387), .ZN(n3385) );
  AND2_X1 U2995 ( .A1(n3869), .A2(n4041), .ZN(n3917) );
  INV_X1 U2996 ( .A(n4492), .ZN(n2331) );
  NAND2_X1 U2997 ( .A1(n3010), .A2(n3009), .ZN(n3011) );
  OR2_X1 U2998 ( .A1(n3482), .A2(n2643), .ZN(n2595) );
  AND2_X1 U2999 ( .A1(n4491), .A2(REG1_REG_5__SCAN_IN), .ZN(n2816) );
  NAND2_X1 U3000 ( .A1(n3792), .A2(n3789), .ZN(n2699) );
  INV_X1 U3001 ( .A(n4275), .ZN(n4296) );
  NAND2_X1 U3002 ( .A1(n3850), .A2(DATAI_3_), .ZN(n2332) );
  INV_X1 U3003 ( .A(REG3_REG_19__SCAN_IN), .ZN(n3639) );
  INV_X1 U3004 ( .A(n4154), .ZN(n4147) );
  AND3_X1 U3005 ( .A1(n2560), .A2(n2559), .A3(n2558), .ZN(n4217) );
  INV_X1 U3006 ( .A(n2699), .ZN(n3880) );
  AND2_X1 U3007 ( .A1(n3850), .A2(DATAI_25_), .ZN(n4064) );
  NAND2_X1 U3008 ( .A1(n4100), .A2(n4120), .ZN(n2732) );
  INV_X1 U3009 ( .A(n4211), .ZN(n2727) );
  MUX2_X1 U3010 ( .A(n4558), .B(DATAI_15_), .S(n3850), .Z(n4238) );
  INV_X1 U3011 ( .A(n3233), .ZN(n3249) );
  NAND2_X1 U3012 ( .A1(n3120), .A2(n3119), .ZN(n3118) );
  AND2_X1 U3013 ( .A1(n2879), .A2(n2303), .ZN(n2978) );
  NAND2_X1 U3014 ( .A1(n2371), .A2(n2370), .ZN(n2374) );
  INV_X1 U3015 ( .A(n4191), .ZN(n4184) );
  INV_X1 U3016 ( .A(n3752), .ZN(n3780) );
  OR2_X1 U3017 ( .A1(n4012), .A2(n2643), .ZN(n2649) );
  OR2_X1 U3018 ( .A1(n4156), .A2(n2643), .ZN(n2573) );
  AND2_X1 U3019 ( .A1(n2776), .A2(n2774), .ZN(n2791) );
  AND2_X1 U3020 ( .A1(n2791), .A2(n3935), .ZN(n4559) );
  AND2_X1 U3021 ( .A1(n2888), .A2(n2887), .ZN(n4618) );
  INV_X1 U3022 ( .A(n4395), .ZN(n4372) );
  AND2_X1 U3023 ( .A1(n3863), .A2(n4093), .ZN(n4127) );
  AND2_X1 U3024 ( .A1(n4303), .A2(n4648), .ZN(n4668) );
  AND2_X1 U3025 ( .A1(n4613), .A2(n2692), .ZN(n4658) );
  AND3_X1 U3026 ( .A1(n2978), .A2(n2878), .A3(n2890), .ZN(n2743) );
  XNOR2_X1 U3027 ( .A(n2377), .B(IR_REG_15__SCAN_IN), .ZN(n4558) );
  AND2_X1 U3028 ( .A1(n2776), .A2(n2775), .ZN(n4595) );
  NAND2_X1 U3029 ( .A1(n2309), .A2(n3441), .ZN(n3452) );
  NAND2_X1 U3030 ( .A1(n2886), .A2(n3935), .ZN(n3776) );
  NAND2_X1 U3031 ( .A1(n2649), .A2(n2648), .ZN(n3943) );
  NAND2_X1 U3032 ( .A1(n2588), .A2(n2587), .ZN(n4149) );
  OAI211_X1 U3033 ( .C1(n2620), .C2(n4454), .A(n2529), .B(n2528), .ZN(n4250)
         );
  INV_X1 U3034 ( .A(n3245), .ZN(n3950) );
  OR2_X1 U3035 ( .A1(n2862), .A2(n4631), .ZN(n3955) );
  INV_X1 U3036 ( .A(n4584), .ZN(n4590) );
  INV_X1 U3037 ( .A(n4559), .ZN(n4604) );
  NAND2_X1 U3038 ( .A1(n4289), .A2(n3090), .ZN(n4242) );
  OR2_X1 U3039 ( .A1(n4192), .A2(n4661), .ZN(n4317) );
  AND2_X2 U3040 ( .A1(n2743), .A2(n2880), .ZN(n4684) );
  NAND2_X1 U3041 ( .A1(n4675), .A2(n4653), .ZN(n4476) );
  NAND2_X1 U3042 ( .A1(n2743), .A2(n2979), .ZN(n4673) );
  NAND2_X1 U3043 ( .A1(n2767), .A2(n2887), .ZN(n4628) );
  XNOR2_X1 U3044 ( .A(n2373), .B(IR_REG_14__SCAN_IN), .ZN(n4512) );
  INV_X1 U3045 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3570) );
  INV_X1 U3046 ( .A(n2327), .ZN(n2311) );
  INV_X1 U3047 ( .A(n2787), .ZN(n4494) );
  NAND4_X1 U3048 ( .A1(n3507), .A2(n2276), .A3(n2398), .A4(n2321), .ZN(n2411)
         );
  NOR2_X1 U3049 ( .A1(n2413), .A2(n2411), .ZN(n2322) );
  NAND2_X1 U3050 ( .A1(n3604), .A2(IR_REG_27__SCAN_IN), .ZN(n2324) );
  MUX2_X1 U3051 ( .A(n4494), .B(DATAI_1_), .S(n2338), .Z(n2892) );
  MUX2_X1 U3052 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2338), .Z(n3466) );
  MUX2_X1 U3053 ( .A(n4493), .B(DATAI_2_), .S(n2338), .Z(n3736) );
  NAND2_X1 U3054 ( .A1(n2307), .A2(IR_REG_31__SCAN_IN), .ZN(n2335) );
  XNOR2_X1 U3055 ( .A(n2335), .B(IR_REG_3__SCAN_IN), .ZN(n4492) );
  INV_X1 U3056 ( .A(IR_REG_3__SCAN_IN), .ZN(n2334) );
  NAND2_X1 U3057 ( .A1(n2335), .A2(n2334), .ZN(n2336) );
  NAND2_X1 U3058 ( .A1(n2336), .A2(IR_REG_31__SCAN_IN), .ZN(n2337) );
  MUX2_X1 U3059 ( .A(n4529), .B(DATAI_4_), .S(n2338), .Z(n3000) );
  NAND2_X1 U3060 ( .A1(n2340), .A2(IR_REG_31__SCAN_IN), .ZN(n2339) );
  MUX2_X1 U3061 ( .A(IR_REG_31__SCAN_IN), .B(n2339), .S(IR_REG_5__SCAN_IN), 
        .Z(n2343) );
  INV_X1 U3062 ( .A(n2340), .ZN(n2342) );
  INV_X1 U3063 ( .A(IR_REG_5__SCAN_IN), .ZN(n2341) );
  NAND2_X1 U3064 ( .A1(n2342), .A2(n2341), .ZN(n2345) );
  INV_X1 U3065 ( .A(DATAI_5_), .ZN(n2344) );
  MUX2_X1 U3066 ( .A(n2835), .B(n2344), .S(n3850), .Z(n3119) );
  NAND2_X1 U3067 ( .A1(n2345), .A2(IR_REG_31__SCAN_IN), .ZN(n2346) );
  MUX2_X1 U3068 ( .A(n4490), .B(DATAI_6_), .S(n3850), .Z(n3051) );
  NAND2_X1 U3069 ( .A1(n2413), .A2(IR_REG_31__SCAN_IN), .ZN(n2347) );
  NAND2_X1 U3070 ( .A1(n2347), .A2(n2352), .ZN(n2349) );
  OR2_X1 U3071 ( .A1(n2347), .A2(n2352), .ZN(n2348) );
  MUX2_X1 U3072 ( .A(n4489), .B(DATAI_7_), .S(n3850), .Z(n3137) );
  NAND2_X1 U3073 ( .A1(n2349), .A2(IR_REG_31__SCAN_IN), .ZN(n2350) );
  XNOR2_X1 U3074 ( .A(n2350), .B(n2351), .ZN(n3063) );
  INV_X1 U3075 ( .A(DATAI_8_), .ZN(n2758) );
  MUX2_X1 U3076 ( .A(n3063), .B(n2758), .S(n3850), .Z(n3184) );
  INV_X1 U3077 ( .A(n2413), .ZN(n2397) );
  NAND2_X1 U3078 ( .A1(n2397), .A2(n2299), .ZN(n2381) );
  NAND2_X1 U3079 ( .A1(n2381), .A2(IR_REG_31__SCAN_IN), .ZN(n2353) );
  MUX2_X1 U3080 ( .A(IR_REG_31__SCAN_IN), .B(n2353), .S(IR_REG_9__SCAN_IN), 
        .Z(n2354) );
  INV_X1 U3081 ( .A(n2354), .ZN(n2355) );
  NOR2_X1 U3082 ( .A1(n2355), .A2(n2359), .ZN(n4488) );
  MUX2_X1 U3083 ( .A(n4488), .B(DATAI_9_), .S(n3850), .Z(n3233) );
  OR2_X1 U3084 ( .A1(n2359), .A2(n2763), .ZN(n2357) );
  MUX2_X1 U3085 ( .A(n4487), .B(DATAI_10_), .S(n3850), .Z(n3264) );
  NAND2_X1 U3086 ( .A1(n2360), .A2(IR_REG_11__SCAN_IN), .ZN(n2363) );
  INV_X1 U3087 ( .A(n2360), .ZN(n2362) );
  INV_X1 U3088 ( .A(IR_REG_11__SCAN_IN), .ZN(n2361) );
  NAND2_X1 U3089 ( .A1(n2362), .A2(n2361), .ZN(n2364) );
  MUX2_X1 U3090 ( .A(n4486), .B(DATAI_11_), .S(n3850), .Z(n4311) );
  NAND2_X1 U3091 ( .A1(n2364), .A2(IR_REG_31__SCAN_IN), .ZN(n2365) );
  XNOR2_X1 U3092 ( .A(n2365), .B(IR_REG_12__SCAN_IN), .ZN(n4485) );
  MUX2_X1 U3093 ( .A(n4485), .B(DATAI_12_), .S(n3850), .Z(n3316) );
  NOR2_X1 U3094 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2366)
         );
  NOR2_X1 U3095 ( .A1(n2371), .A2(n2763), .ZN(n2368) );
  MUX2_X1 U3096 ( .A(n2763), .B(n2368), .S(IR_REG_13__SCAN_IN), .Z(n2369) );
  INV_X1 U3097 ( .A(n2369), .ZN(n2372) );
  INV_X1 U3098 ( .A(IR_REG_13__SCAN_IN), .ZN(n2370) );
  MUX2_X1 U3099 ( .A(n3992), .B(DATAI_13_), .S(n3850), .Z(n2723) );
  NAND2_X1 U3100 ( .A1(n2374), .A2(IR_REG_31__SCAN_IN), .ZN(n2373) );
  MUX2_X1 U3101 ( .A(n4512), .B(DATAI_14_), .S(n3850), .Z(n4256) );
  NAND2_X1 U3102 ( .A1(n2375), .A2(IR_REG_31__SCAN_IN), .ZN(n2377) );
  INV_X1 U3103 ( .A(IR_REG_15__SCAN_IN), .ZN(n2376) );
  NAND2_X1 U3104 ( .A1(n2377), .A2(n2376), .ZN(n2378) );
  NAND2_X1 U3105 ( .A1(n2378), .A2(IR_REG_31__SCAN_IN), .ZN(n2380) );
  INV_X1 U3106 ( .A(IR_REG_16__SCAN_IN), .ZN(n2379) );
  INV_X1 U3107 ( .A(DATAI_16_), .ZN(n4637) );
  MUX2_X1 U3108 ( .A(n4638), .B(n4637), .S(n3850), .Z(n3671) );
  NAND2_X1 U3109 ( .A1(n2393), .A2(n2003), .ZN(n2384) );
  NAND2_X1 U3110 ( .A1(n2384), .A2(IR_REG_31__SCAN_IN), .ZN(n2382) );
  XNOR2_X1 U3111 ( .A(n2382), .B(IR_REG_17__SCAN_IN), .ZN(n4635) );
  INV_X1 U3112 ( .A(n4635), .ZN(n4589) );
  INV_X1 U3113 ( .A(DATAI_17_), .ZN(n2383) );
  MUX2_X1 U3114 ( .A(n4589), .B(n2383), .S(n3850), .Z(n3339) );
  INV_X1 U3115 ( .A(n2384), .ZN(n2385) );
  NAND2_X1 U3116 ( .A1(n2385), .A2(n2389), .ZN(n2386) );
  NAND2_X1 U3117 ( .A1(n2386), .A2(IR_REG_31__SCAN_IN), .ZN(n2387) );
  XNOR2_X1 U3118 ( .A(n2387), .B(IR_REG_18__SCAN_IN), .ZN(n4633) );
  INV_X1 U3119 ( .A(n4633), .ZN(n4603) );
  INV_X1 U3120 ( .A(DATAI_18_), .ZN(n2388) );
  MUX2_X1 U3121 ( .A(n4603), .B(n2388), .S(n3850), .Z(n4191) );
  NAND2_X1 U3122 ( .A1(n2410), .A2(IR_REG_31__SCAN_IN), .ZN(n2394) );
  XNOR2_X2 U3123 ( .A(n2394), .B(n2403), .ZN(n2865) );
  INV_X1 U3124 ( .A(DATAI_19_), .ZN(n2395) );
  MUX2_X1 U3125 ( .A(n2865), .B(n2395), .S(n3850), .Z(n3640) );
  NAND2_X1 U3126 ( .A1(n3850), .A2(DATAI_23_), .ZN(n3483) );
  NAND2_X1 U3127 ( .A1(n3850), .A2(DATAI_24_), .ZN(n4080) );
  NAND2_X1 U3128 ( .A1(n3850), .A2(DATAI_26_), .ZN(n4051) );
  INV_X1 U3129 ( .A(n4051), .ZN(n2736) );
  AND2_X1 U3130 ( .A1(n3850), .A2(DATAI_28_), .ZN(n3446) );
  AND2_X1 U3131 ( .A1(n3850), .A2(DATAI_29_), .ZN(n3835) );
  NAND2_X1 U3132 ( .A1(n2752), .A2(n3835), .ZN(n2396) );
  NAND2_X1 U3133 ( .A1(n4004), .A2(n2396), .ZN(n4014) );
  NAND2_X1 U3134 ( .A1(n2672), .A2(IR_REG_31__SCAN_IN), .ZN(n2399) );
  MUX2_X1 U3135 ( .A(n2401), .B(IR_REG_31__SCAN_IN), .S(n2398), .Z(n2402) );
  NAND2_X1 U3136 ( .A1(n2406), .A2(n2403), .ZN(n2409) );
  NAND3_X1 U3137 ( .A1(n2410), .A2(IR_REG_31__SCAN_IN), .A3(IR_REG_20__SCAN_IN), .ZN(n2408) );
  NAND2_X1 U3138 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2404) );
  NAND2_X1 U3139 ( .A1(n2404), .A2(IR_REG_31__SCAN_IN), .ZN(n2405) );
  OAI21_X1 U3140 ( .B1(n2406), .B2(IR_REG_31__SCAN_IN), .A(n2405), .ZN(n2407)
         );
  OR2_X1 U3141 ( .A1(n4014), .A2(n4661), .ZN(n2668) );
  INV_X1 U3142 ( .A(n2411), .ZN(n2412) );
  NAND2_X1 U3143 ( .A1(n2412), .A2(n2300), .ZN(n2414) );
  NAND2_X1 U3144 ( .A1(n2416), .A2(n2415), .ZN(n2652) );
  NOR2_X2 U3145 ( .A1(n2652), .A2(IR_REG_28__SCAN_IN), .ZN(n2419) );
  INV_X1 U3146 ( .A(n2419), .ZN(n2655) );
  NAND2_X1 U3147 ( .A1(n2419), .A2(n2418), .ZN(n2764) );
  XNOR2_X2 U31480 ( .A(n2420), .B(IR_REG_30__SCAN_IN), .ZN(n3428) );
  NAND2_X1 U31490 ( .A1(n2868), .A2(n2864), .ZN(n3785) );
  NAND2_X1 U3150 ( .A1(n3468), .A2(n2892), .ZN(n3788) );
  NAND2_X1 U3151 ( .A1(n2448), .A2(REG3_REG_0__SCAN_IN), .ZN(n2425) );
  NAND2_X1 U3152 ( .A1(n2431), .A2(REG2_REG_0__SCAN_IN), .ZN(n2423) );
  NAND2_X1 U3153 ( .A1(n2432), .A2(REG1_REG_0__SCAN_IN), .ZN(n2422) );
  INV_X1 U3154 ( .A(n3956), .ZN(n2426) );
  NAND2_X1 U3155 ( .A1(n2426), .A2(n3466), .ZN(n3784) );
  NAND2_X1 U3156 ( .A1(n2007), .A2(REG0_REG_2__SCAN_IN), .ZN(n2430) );
  NAND2_X1 U3157 ( .A1(n2431), .A2(REG2_REG_2__SCAN_IN), .ZN(n2429) );
  NAND2_X1 U3158 ( .A1(n2432), .A2(REG1_REG_2__SCAN_IN), .ZN(n2428) );
  AND4_X2 U3159 ( .A1(n2430), .A2(n2429), .A3(n2428), .A4(n2427), .ZN(n2928)
         );
  OR2_X1 U3160 ( .A1(n3736), .A2(n2928), .ZN(n3792) );
  NAND2_X1 U3161 ( .A1(n2928), .A2(n3736), .ZN(n3789) );
  NAND2_X1 U3162 ( .A1(n3032), .A2(n3880), .ZN(n3031) );
  NAND2_X1 U3163 ( .A1(n3031), .A2(n3789), .ZN(n3070) );
  NAND2_X1 U3164 ( .A1(n3845), .A2(REG2_REG_3__SCAN_IN), .ZN(n2438) );
  NAND2_X1 U3165 ( .A1(n2007), .A2(REG0_REG_3__SCAN_IN), .ZN(n2434) );
  INV_X1 U3166 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2441) );
  NAND2_X1 U3167 ( .A1(n2448), .A2(n2441), .ZN(n2433) );
  NAND2_X1 U3168 ( .A1(n2434), .A2(n2433), .ZN(n2435) );
  NAND2_X1 U3169 ( .A1(n2945), .A2(n3078), .ZN(n3794) );
  INV_X1 U3170 ( .A(n3078), .ZN(n3072) );
  NAND2_X1 U3171 ( .A1(n3072), .A2(n3737), .ZN(n3791) );
  AND2_X2 U3172 ( .A1(n3794), .A2(n3791), .ZN(n3882) );
  NAND2_X1 U3173 ( .A1(n3070), .A2(n3882), .ZN(n2439) );
  NAND2_X1 U3174 ( .A1(n3845), .A2(REG2_REG_4__SCAN_IN), .ZN(n2446) );
  NAND2_X1 U3175 ( .A1(n2432), .A2(REG1_REG_4__SCAN_IN), .ZN(n2445) );
  NAND2_X1 U3176 ( .A1(n2007), .A2(REG0_REG_4__SCAN_IN), .ZN(n2444) );
  INV_X1 U3177 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2440) );
  NAND2_X1 U3178 ( .A1(n2441), .A2(n2440), .ZN(n2442) );
  AND2_X1 U3179 ( .A1(n2442), .A2(n2451), .ZN(n3001) );
  NAND2_X1 U3180 ( .A1(n2448), .A2(n3001), .ZN(n2443) );
  NAND2_X1 U3181 ( .A1(n2932), .A2(n3000), .ZN(n3795) );
  INV_X1 U3182 ( .A(n3795), .ZN(n2447) );
  NAND2_X1 U3183 ( .A1(n2944), .A2(n3953), .ZN(n3798) );
  NAND2_X1 U3184 ( .A1(n2432), .A2(REG1_REG_5__SCAN_IN), .ZN(n2456) );
  NAND2_X1 U3185 ( .A1(n3846), .A2(REG0_REG_5__SCAN_IN), .ZN(n2455) );
  INV_X1 U3186 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2450) );
  NAND2_X1 U3187 ( .A1(n2451), .A2(n2450), .ZN(n2452) );
  AND2_X1 U3188 ( .A1(n2458), .A2(n2452), .ZN(n3121) );
  NAND2_X1 U3189 ( .A1(n2617), .A2(n3121), .ZN(n2454) );
  NAND2_X1 U3190 ( .A1(n3845), .A2(REG2_REG_5__SCAN_IN), .ZN(n2453) );
  INV_X1 U3191 ( .A(n3119), .ZN(n2706) );
  NAND2_X1 U3192 ( .A1(n3046), .A2(n2706), .ZN(n3802) );
  INV_X1 U3193 ( .A(n3046), .ZN(n3952) );
  AND2_X1 U3194 ( .A1(n3119), .A2(n3952), .ZN(n3110) );
  INV_X1 U3195 ( .A(n3051), .ZN(n3021) );
  NAND2_X1 U3196 ( .A1(n3845), .A2(REG2_REG_6__SCAN_IN), .ZN(n2463) );
  NAND2_X1 U3197 ( .A1(n2432), .A2(REG1_REG_6__SCAN_IN), .ZN(n2462) );
  INV_X1 U3198 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2457) );
  NAND2_X1 U3199 ( .A1(n2458), .A2(n2457), .ZN(n2459) );
  AND2_X1 U3200 ( .A1(n2473), .A2(n2459), .ZN(n3091) );
  NAND2_X1 U3201 ( .A1(n2617), .A2(n3091), .ZN(n2461) );
  NAND2_X1 U3202 ( .A1(n3846), .A2(REG0_REG_6__SCAN_IN), .ZN(n2460) );
  NAND4_X1 U3203 ( .A1(n2463), .A2(n2462), .A3(n2461), .A4(n2460), .ZN(n3114)
         );
  NAND2_X1 U3204 ( .A1(n3021), .A2(n3114), .ZN(n3800) );
  NAND2_X1 U3205 ( .A1(n3045), .A2(n3800), .ZN(n2464) );
  INV_X1 U3206 ( .A(n3114), .ZN(n3133) );
  NAND2_X1 U3207 ( .A1(n3133), .A2(n3051), .ZN(n3804) );
  NAND2_X1 U3208 ( .A1(n3845), .A2(REG2_REG_7__SCAN_IN), .ZN(n2468) );
  NAND2_X1 U3209 ( .A1(n2656), .A2(REG1_REG_7__SCAN_IN), .ZN(n2467) );
  XNOR2_X1 U32100 ( .A(n2473), .B(REG3_REG_7__SCAN_IN), .ZN(n3104) );
  NAND2_X1 U32110 ( .A1(n2617), .A2(n3104), .ZN(n2466) );
  NAND2_X1 U32120 ( .A1(n3846), .A2(REG0_REG_7__SCAN_IN), .ZN(n2465) );
  NAND2_X1 U32130 ( .A1(n3185), .A2(n3137), .ZN(n3805) );
  INV_X1 U32140 ( .A(n3805), .ZN(n2469) );
  INV_X1 U32150 ( .A(n3137), .ZN(n2470) );
  NAND2_X1 U32160 ( .A1(n2470), .A2(n3951), .ZN(n3807) );
  NAND2_X1 U32170 ( .A1(n2656), .A2(REG1_REG_8__SCAN_IN), .ZN(n2478) );
  NAND2_X1 U32180 ( .A1(n3846), .A2(REG0_REG_8__SCAN_IN), .ZN(n2477) );
  INV_X1 U32190 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2472) );
  INV_X1 U32200 ( .A(REG3_REG_8__SCAN_IN), .ZN(n3183) );
  OAI21_X1 U32210 ( .B1(n2473), .B2(n2472), .A(n3183), .ZN(n2474) );
  AND2_X1 U32220 ( .A1(n2481), .A2(n2474), .ZN(n3188) );
  NAND2_X1 U32230 ( .A1(n2617), .A2(n3188), .ZN(n2476) );
  NAND2_X1 U32240 ( .A1(n3845), .A2(REG2_REG_8__SCAN_IN), .ZN(n2475) );
  INV_X1 U32250 ( .A(n3184), .ZN(n2713) );
  NAND2_X1 U32260 ( .A1(n3245), .A2(n2713), .ZN(n3810) );
  NAND2_X1 U32270 ( .A1(n3184), .A2(n3950), .ZN(n3806) );
  NAND2_X1 U32280 ( .A1(n3845), .A2(REG2_REG_9__SCAN_IN), .ZN(n2486) );
  NAND2_X1 U32290 ( .A1(n2432), .A2(REG1_REG_9__SCAN_IN), .ZN(n2485) );
  INV_X1 U32300 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2480) );
  NAND2_X1 U32310 ( .A1(n2481), .A2(n2480), .ZN(n2482) );
  AND2_X1 U32320 ( .A1(n2488), .A2(n2482), .ZN(n3246) );
  NAND2_X1 U32330 ( .A1(n2617), .A2(n3246), .ZN(n2484) );
  NAND2_X1 U32340 ( .A1(n3846), .A2(REG0_REG_9__SCAN_IN), .ZN(n2483) );
  NAND4_X1 U32350 ( .A1(n2486), .A2(n2485), .A3(n2484), .A4(n2483), .ZN(n3949)
         );
  AND2_X1 U32360 ( .A1(n3249), .A2(n3949), .ZN(n3814) );
  NAND2_X1 U32370 ( .A1(n3627), .A2(n3233), .ZN(n3811) );
  INV_X1 U32380 ( .A(n3264), .ZN(n3631) );
  NAND2_X1 U32390 ( .A1(n2432), .A2(REG1_REG_10__SCAN_IN), .ZN(n2493) );
  NAND2_X1 U32400 ( .A1(n3846), .A2(REG0_REG_10__SCAN_IN), .ZN(n2492) );
  NAND2_X1 U32410 ( .A1(n2488), .A2(n2487), .ZN(n2489) );
  AND2_X1 U32420 ( .A1(n2497), .A2(n2489), .ZN(n3628) );
  NAND2_X1 U32430 ( .A1(n2617), .A2(n3628), .ZN(n2491) );
  NAND2_X1 U32440 ( .A1(n3845), .A2(REG2_REG_10__SCAN_IN), .ZN(n2490) );
  NAND4_X1 U32450 ( .A1(n2493), .A2(n2492), .A3(n2491), .A4(n2490), .ZN(n3948)
         );
  NAND2_X1 U32460 ( .A1(n3631), .A2(n3948), .ZN(n3816) );
  NAND2_X1 U32470 ( .A1(n3216), .A2(n3816), .ZN(n2494) );
  NAND2_X1 U32480 ( .A1(n4297), .A2(n3264), .ZN(n3813) );
  INV_X1 U32490 ( .A(n4311), .ZN(n3272) );
  NAND2_X1 U32500 ( .A1(n2656), .A2(REG1_REG_11__SCAN_IN), .ZN(n2502) );
  NAND2_X1 U32510 ( .A1(n3846), .A2(REG0_REG_11__SCAN_IN), .ZN(n2501) );
  INV_X1 U32520 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2496) );
  NAND2_X1 U32530 ( .A1(n2497), .A2(n2496), .ZN(n2498) );
  AND2_X1 U32540 ( .A1(n2511), .A2(n2498), .ZN(n4315) );
  NAND2_X1 U32550 ( .A1(n2617), .A2(n4315), .ZN(n2500) );
  NAND2_X1 U32560 ( .A1(n3845), .A2(REG2_REG_11__SCAN_IN), .ZN(n2499) );
  INV_X1 U32570 ( .A(n3626), .ZN(n3947) );
  NAND2_X1 U32580 ( .A1(n3272), .A2(n3947), .ZN(n3817) );
  INV_X1 U32590 ( .A(n2723), .ZN(n4285) );
  NAND2_X1 U32600 ( .A1(n2656), .A2(REG1_REG_13__SCAN_IN), .ZN(n2510) );
  NAND2_X1 U32610 ( .A1(n3846), .A2(REG0_REG_13__SCAN_IN), .ZN(n2509) );
  INV_X1 U32620 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2504) );
  INV_X1 U32630 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2503) );
  OAI21_X1 U32640 ( .B1(n2511), .B2(n2504), .A(n2503), .ZN(n2506) );
  NAND2_X1 U32650 ( .A1(REG3_REG_12__SCAN_IN), .A2(REG3_REG_13__SCAN_IN), .ZN(
        n2505) );
  AND2_X1 U32660 ( .A1(n2506), .A2(n2519), .ZN(n4286) );
  NAND2_X1 U32670 ( .A1(n2617), .A2(n4286), .ZN(n2508) );
  NAND2_X1 U32680 ( .A1(n3845), .A2(REG2_REG_13__SCAN_IN), .ZN(n2507) );
  NAND4_X1 U32690 ( .A1(n2510), .A2(n2509), .A3(n2508), .A4(n2507), .ZN(n4249)
         );
  NAND2_X1 U32700 ( .A1(n4285), .A2(n4249), .ZN(n3891) );
  NAND2_X1 U32710 ( .A1(n3845), .A2(REG2_REG_12__SCAN_IN), .ZN(n2515) );
  NAND2_X1 U32720 ( .A1(n2432), .A2(REG1_REG_12__SCAN_IN), .ZN(n2514) );
  XNOR2_X1 U32730 ( .A(n2511), .B(REG3_REG_12__SCAN_IN), .ZN(n3425) );
  NAND2_X1 U32740 ( .A1(n2617), .A2(n3425), .ZN(n2513) );
  NAND2_X1 U32750 ( .A1(n3846), .A2(REG0_REG_12__SCAN_IN), .ZN(n2512) );
  NAND4_X1 U32760 ( .A1(n2515), .A2(n2514), .A3(n2513), .A4(n2512), .ZN(n4274)
         );
  NAND2_X1 U32770 ( .A1(n3421), .A2(n4274), .ZN(n4269) );
  NAND2_X1 U32780 ( .A1(n3626), .A2(n4311), .ZN(n3297) );
  INV_X1 U32790 ( .A(n4274), .ZN(n4299) );
  NAND2_X1 U32800 ( .A1(n4299), .A2(n3316), .ZN(n4268) );
  NAND2_X1 U32810 ( .A1(n3297), .A2(n4268), .ZN(n2517) );
  INV_X1 U32820 ( .A(n4249), .ZN(n3422) );
  NAND2_X1 U32830 ( .A1(n2723), .A2(n3422), .ZN(n3890) );
  INV_X1 U32840 ( .A(n3890), .ZN(n2516) );
  AOI21_X1 U32850 ( .B1(n2008), .B2(n2517), .A(n2516), .ZN(n3820) );
  INV_X1 U32860 ( .A(REG3_REG_14__SCAN_IN), .ZN(n3544) );
  NAND2_X1 U32870 ( .A1(n2519), .A2(n3544), .ZN(n2520) );
  NAND2_X1 U32880 ( .A1(n2526), .A2(n2520), .ZN(n4258) );
  OR2_X1 U32890 ( .A1(n2643), .A2(n4258), .ZN(n2524) );
  NAND2_X1 U32900 ( .A1(n2432), .A2(REG1_REG_14__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U32910 ( .A1(n3846), .A2(REG0_REG_14__SCAN_IN), .ZN(n2522) );
  NAND2_X1 U32920 ( .A1(n3845), .A2(REG2_REG_14__SCAN_IN), .ZN(n2521) );
  NAND2_X1 U32930 ( .A1(n4228), .A2(n4256), .ZN(n4232) );
  INV_X1 U32940 ( .A(n4228), .ZN(n4277) );
  INV_X1 U32950 ( .A(n4256), .ZN(n4252) );
  NAND2_X1 U32960 ( .A1(n4277), .A2(n4252), .ZN(n3823) );
  NAND2_X1 U32970 ( .A1(n4232), .A2(n3823), .ZN(n4244) );
  INV_X1 U32980 ( .A(n4244), .ZN(n4248) );
  INV_X1 U32990 ( .A(n4238), .ZN(n3774) );
  INV_X1 U33000 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4454) );
  NAND2_X1 U33010 ( .A1(n2526), .A2(n2525), .ZN(n2527) );
  NAND2_X1 U33020 ( .A1(n2533), .A2(n2527), .ZN(n3773) );
  OR2_X1 U33030 ( .A1(n3773), .A2(n2643), .ZN(n2529) );
  AOI22_X1 U33040 ( .A1(n3845), .A2(REG2_REG_15__SCAN_IN), .B1(n2432), .B2(
        REG1_REG_15__SCAN_IN), .ZN(n2528) );
  NAND2_X1 U33050 ( .A1(n3774), .A2(n4250), .ZN(n3822) );
  INV_X1 U33060 ( .A(n4250), .ZN(n3672) );
  NAND2_X1 U33070 ( .A1(n3672), .A2(n4238), .ZN(n3824) );
  NAND2_X1 U33080 ( .A1(n3822), .A2(n3824), .ZN(n3868) );
  INV_X1 U33090 ( .A(n4232), .ZN(n2530) );
  NOR2_X1 U33100 ( .A1(n3868), .A2(n2530), .ZN(n2531) );
  NAND2_X1 U33110 ( .A1(n4246), .A2(n2531), .ZN(n4230) );
  NAND2_X1 U33120 ( .A1(n4230), .A2(n3822), .ZN(n4214) );
  INV_X1 U33130 ( .A(n3671), .ZN(n4221) );
  NAND2_X1 U33140 ( .A1(n2533), .A2(n2532), .ZN(n2534) );
  AND2_X1 U33150 ( .A1(n2555), .A2(n2534), .ZN(n4220) );
  NAND2_X1 U33160 ( .A1(n4220), .A2(n2617), .ZN(n2537) );
  AOI22_X1 U33170 ( .A1(n3845), .A2(REG2_REG_16__SCAN_IN), .B1(n2656), .B2(
        REG1_REG_16__SCAN_IN), .ZN(n2536) );
  NAND2_X1 U33180 ( .A1(n3846), .A2(REG0_REG_16__SCAN_IN), .ZN(n2535) );
  NAND2_X1 U33190 ( .A1(n4221), .A2(n4229), .ZN(n3905) );
  NAND2_X1 U33200 ( .A1(n3671), .A2(n4203), .ZN(n3903) );
  NAND2_X1 U33210 ( .A1(n4214), .A2(n4211), .ZN(n2538) );
  NAND2_X1 U33220 ( .A1(n2547), .A2(n3639), .ZN(n2540) );
  AND2_X1 U33230 ( .A1(n2567), .A2(n2540), .ZN(n4163) );
  NAND2_X1 U33240 ( .A1(n4163), .A2(n2617), .ZN(n2545) );
  INV_X1 U33250 ( .A(REG0_REG_19__SCAN_IN), .ZN(n3581) );
  NAND2_X1 U33260 ( .A1(n2432), .A2(REG1_REG_19__SCAN_IN), .ZN(n2542) );
  NAND2_X1 U33270 ( .A1(n3845), .A2(REG2_REG_19__SCAN_IN), .ZN(n2541) );
  OAI211_X1 U33280 ( .C1(n2620), .C2(n3581), .A(n2542), .B(n2541), .ZN(n2543)
         );
  INV_X1 U33290 ( .A(n2543), .ZN(n2544) );
  NAND2_X1 U33300 ( .A1(n3946), .A2(n3640), .ZN(n2553) );
  INV_X1 U33310 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3751) );
  NAND2_X1 U33320 ( .A1(n2557), .A2(n3751), .ZN(n2546) );
  NAND2_X1 U33330 ( .A1(n2547), .A2(n2546), .ZN(n4193) );
  OR2_X1 U33340 ( .A1(n4193), .A2(n2643), .ZN(n2552) );
  INV_X1 U33350 ( .A(n2432), .ZN(n2646) );
  INV_X1 U33360 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4509) );
  NAND2_X1 U33370 ( .A1(n3845), .A2(REG2_REG_18__SCAN_IN), .ZN(n2549) );
  NAND2_X1 U33380 ( .A1(n3846), .A2(REG0_REG_18__SCAN_IN), .ZN(n2548) );
  OAI211_X1 U33390 ( .C1(n2646), .C2(n4509), .A(n2549), .B(n2548), .ZN(n2550)
         );
  INV_X1 U33400 ( .A(n2550), .ZN(n2551) );
  NAND2_X1 U33410 ( .A1(n4173), .A2(n4191), .ZN(n4168) );
  NAND2_X1 U33420 ( .A1(n2553), .A2(n4168), .ZN(n2562) );
  INV_X1 U33430 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2554) );
  NAND2_X1 U33440 ( .A1(n2555), .A2(n2554), .ZN(n2556) );
  NAND2_X1 U33450 ( .A1(n2557), .A2(n2556), .ZN(n4199) );
  OR2_X1 U33460 ( .A1(n4199), .A2(n2643), .ZN(n2560) );
  AOI22_X1 U33470 ( .A1(n2656), .A2(REG1_REG_17__SCAN_IN), .B1(n3846), .B2(
        REG0_REG_17__SCAN_IN), .ZN(n2559) );
  NAND2_X1 U33480 ( .A1(n3845), .A2(REG2_REG_17__SCAN_IN), .ZN(n2558) );
  AND2_X1 U33490 ( .A1(n4185), .A2(n3339), .ZN(n4166) );
  NAND2_X1 U33500 ( .A1(n4205), .A2(n4184), .ZN(n4167) );
  INV_X1 U33510 ( .A(n3339), .ZN(n4202) );
  NAND2_X1 U33520 ( .A1(n4217), .A2(n4202), .ZN(n4165) );
  AND2_X1 U3353 ( .A1(n4167), .A2(n4165), .ZN(n2563) );
  OR2_X1 U33540 ( .A1(n2563), .A2(n2562), .ZN(n2565) );
  NAND2_X1 U3355 ( .A1(n4187), .A2(n4172), .ZN(n2564) );
  NAND2_X1 U3356 ( .A1(n2565), .A2(n2564), .ZN(n4144) );
  NAND2_X1 U3357 ( .A1(n2567), .A2(n2083), .ZN(n2568) );
  NAND2_X1 U3358 ( .A1(n2583), .A2(n2568), .ZN(n4156) );
  INV_X1 U3359 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4157) );
  NAND2_X1 U3360 ( .A1(n3846), .A2(REG0_REG_20__SCAN_IN), .ZN(n2570) );
  NAND2_X1 U3361 ( .A1(n2432), .A2(REG1_REG_20__SCAN_IN), .ZN(n2569) );
  OAI211_X1 U3362 ( .C1(n2239), .C2(n4157), .A(n2570), .B(n2569), .ZN(n2571)
         );
  INV_X1 U3363 ( .A(n2571), .ZN(n2572) );
  NOR2_X1 U3364 ( .A1(n4129), .A2(n4147), .ZN(n2574) );
  NOR2_X1 U3365 ( .A1(n4144), .A2(n2574), .ZN(n3829) );
  NAND2_X1 U3366 ( .A1(n4129), .A2(n4147), .ZN(n3907) );
  NAND2_X1 U3367 ( .A1(n2575), .A2(n3907), .ZN(n4091) );
  INV_X1 U3368 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3649) );
  INV_X1 U3369 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3723) );
  OAI21_X1 U3370 ( .B1(n2583), .B2(n3649), .A(n3723), .ZN(n2577) );
  NAND2_X1 U3371 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2576) );
  AND2_X1 U3372 ( .A1(n2577), .A2(n2589), .ZN(n4118) );
  NAND2_X1 U3373 ( .A1(n4118), .A2(n2617), .ZN(n2582) );
  INV_X1 U3374 ( .A(REG1_REG_22__SCAN_IN), .ZN(n3593) );
  NAND2_X1 U3375 ( .A1(n3845), .A2(REG2_REG_22__SCAN_IN), .ZN(n2579) );
  NAND2_X1 U3376 ( .A1(n3846), .A2(REG0_REG_22__SCAN_IN), .ZN(n2578) );
  OAI211_X1 U3377 ( .C1(n2646), .C2(n3593), .A(n2579), .B(n2578), .ZN(n2580)
         );
  INV_X1 U3378 ( .A(n2580), .ZN(n2581) );
  OR2_X1 U3379 ( .A1(n4100), .A2(n4112), .ZN(n4095) );
  XNOR2_X1 U3380 ( .A(n2583), .B(REG3_REG_21__SCAN_IN), .ZN(n4126) );
  NAND2_X1 U3381 ( .A1(n4126), .A2(n2617), .ZN(n2588) );
  INV_X1 U3382 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4134) );
  NAND2_X1 U3383 ( .A1(n3846), .A2(REG0_REG_21__SCAN_IN), .ZN(n2585) );
  NAND2_X1 U3384 ( .A1(n2432), .A2(REG1_REG_21__SCAN_IN), .ZN(n2584) );
  OAI211_X1 U3385 ( .C1(n2239), .C2(n4134), .A(n2585), .B(n2584), .ZN(n2586)
         );
  INV_X1 U3386 ( .A(n2586), .ZN(n2587) );
  INV_X1 U3387 ( .A(n4128), .ZN(n3650) );
  OR2_X1 U3388 ( .A1(n4149), .A2(n3650), .ZN(n4093) );
  AND2_X1 U3389 ( .A1(n4095), .A2(n4093), .ZN(n3912) );
  NAND2_X1 U3390 ( .A1(n4091), .A2(n3912), .ZN(n2598) );
  NAND2_X1 U3391 ( .A1(n2589), .A2(n2084), .ZN(n2590) );
  NAND2_X1 U3392 ( .A1(n2600), .A2(n2590), .ZN(n3482) );
  INV_X1 U3393 ( .A(REG1_REG_23__SCAN_IN), .ZN(n3594) );
  NAND2_X1 U3394 ( .A1(n3845), .A2(REG2_REG_23__SCAN_IN), .ZN(n2592) );
  NAND2_X1 U3395 ( .A1(n3846), .A2(REG0_REG_23__SCAN_IN), .ZN(n2591) );
  OAI211_X1 U3396 ( .C1(n2646), .C2(n3594), .A(n2592), .B(n2591), .ZN(n2593)
         );
  INV_X1 U3397 ( .A(n2593), .ZN(n2594) );
  NAND2_X1 U3398 ( .A1(n2896), .A2(n3483), .ZN(n3864) );
  NAND2_X1 U3399 ( .A1(n4100), .A2(n4112), .ZN(n2596) );
  AND2_X1 U3400 ( .A1(n3864), .A2(n2596), .ZN(n3831) );
  AND2_X1 U3401 ( .A1(n4149), .A2(n3650), .ZN(n4092) );
  NAND2_X1 U3402 ( .A1(n4095), .A2(n4092), .ZN(n2597) );
  NAND2_X1 U3403 ( .A1(n2598), .A2(n3910), .ZN(n2599) );
  NAND2_X1 U3404 ( .A1(n4115), .A2(n4099), .ZN(n3865) );
  INV_X1 U3405 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3696) );
  NAND2_X1 U3406 ( .A1(n2600), .A2(n3696), .ZN(n2601) );
  NAND2_X1 U3407 ( .A1(n2608), .A2(n2601), .ZN(n3695) );
  INV_X1 U3408 ( .A(REG2_REG_24__SCAN_IN), .ZN(n3565) );
  NAND2_X1 U3409 ( .A1(n3846), .A2(REG0_REG_24__SCAN_IN), .ZN(n2603) );
  NAND2_X1 U3410 ( .A1(n2656), .A2(REG1_REG_24__SCAN_IN), .ZN(n2602) );
  OAI211_X1 U3411 ( .C1(n2239), .C2(n3565), .A(n2603), .B(n2602), .ZN(n2604)
         );
  INV_X1 U3412 ( .A(n2604), .ZN(n2605) );
  NOR2_X1 U3413 ( .A1(n4065), .A2(n4080), .ZN(n3861) );
  INV_X1 U3414 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3660) );
  NAND2_X1 U3415 ( .A1(n2608), .A2(n3660), .ZN(n2609) );
  NAND2_X1 U3416 ( .A1(n2615), .A2(n2609), .ZN(n3659) );
  INV_X1 U3417 ( .A(REG0_REG_25__SCAN_IN), .ZN(n3567) );
  NAND2_X1 U3418 ( .A1(n2432), .A2(REG1_REG_25__SCAN_IN), .ZN(n2611) );
  NAND2_X1 U3419 ( .A1(n3845), .A2(REG2_REG_25__SCAN_IN), .ZN(n2610) );
  OAI211_X1 U3420 ( .C1(n2620), .C2(n3567), .A(n2611), .B(n2610), .ZN(n2612)
         );
  INV_X1 U3421 ( .A(n2612), .ZN(n2613) );
  NAND2_X1 U3422 ( .A1(n4077), .A2(n3661), .ZN(n3870) );
  NAND2_X1 U3423 ( .A1(n4065), .A2(n4080), .ZN(n4060) );
  INV_X1 U3424 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3762) );
  NAND2_X1 U3425 ( .A1(n2615), .A2(n3762), .ZN(n2616) );
  INV_X1 U3426 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4410) );
  NAND2_X1 U3427 ( .A1(n2656), .A2(REG1_REG_26__SCAN_IN), .ZN(n2619) );
  NAND2_X1 U3428 ( .A1(n3845), .A2(REG2_REG_26__SCAN_IN), .ZN(n2618) );
  OAI211_X1 U3429 ( .C1(n2620), .C2(n4410), .A(n2619), .B(n2618), .ZN(n2621)
         );
  INV_X1 U3430 ( .A(n2621), .ZN(n2622) );
  OR2_X1 U3431 ( .A1(n3945), .A2(n4051), .ZN(n3869) );
  OR2_X1 U3432 ( .A1(n4077), .A2(n3661), .ZN(n4041) );
  NAND2_X1 U3433 ( .A1(n3945), .A2(n4051), .ZN(n3920) );
  NAND2_X1 U3434 ( .A1(n2623), .A2(n3920), .ZN(n4019) );
  INV_X1 U3435 ( .A(n2625), .ZN(n2624) );
  INV_X1 U3436 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3587) );
  NAND2_X1 U3437 ( .A1(n2625), .A2(n3587), .ZN(n2626) );
  NAND2_X1 U3438 ( .A1(n2634), .A2(n2626), .ZN(n4036) );
  INV_X1 U3439 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4035) );
  NAND2_X1 U3440 ( .A1(n2656), .A2(REG1_REG_27__SCAN_IN), .ZN(n2628) );
  NAND2_X1 U3441 ( .A1(n3846), .A2(REG0_REG_27__SCAN_IN), .ZN(n2627) );
  OAI211_X1 U3442 ( .C1(n4035), .C2(n2239), .A(n2628), .B(n2627), .ZN(n2629)
         );
  INV_X1 U3443 ( .A(n2629), .ZN(n2630) );
  NAND2_X1 U3444 ( .A1(n3763), .A2(n4032), .ZN(n3842) );
  INV_X1 U3445 ( .A(n4032), .ZN(n4022) );
  NAND2_X1 U3446 ( .A1(n4047), .A2(n4022), .ZN(n3838) );
  NAND2_X1 U3447 ( .A1(n3842), .A2(n3838), .ZN(n4029) );
  INV_X1 U3448 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2633) );
  NAND2_X1 U3449 ( .A1(n2634), .A2(n2633), .ZN(n2635) );
  NAND2_X1 U3450 ( .A1(n4012), .A2(n2635), .ZN(n3456) );
  INV_X1 U3451 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2638) );
  NAND2_X1 U3452 ( .A1(n3845), .A2(REG2_REG_28__SCAN_IN), .ZN(n2637) );
  NAND2_X1 U3453 ( .A1(n3846), .A2(REG0_REG_28__SCAN_IN), .ZN(n2636) );
  OAI211_X1 U3454 ( .C1(n2638), .C2(n2646), .A(n2637), .B(n2636), .ZN(n2639)
         );
  INV_X1 U3455 ( .A(n2639), .ZN(n2640) );
  NAND2_X1 U3456 ( .A1(n3944), .A2(n3435), .ZN(n3836) );
  NAND2_X1 U3457 ( .A1(n4025), .A2(n3446), .ZN(n3843) );
  NAND2_X1 U34580 ( .A1(n2642), .A2(n3843), .ZN(n2650) );
  NAND2_X1 U34590 ( .A1(n3845), .A2(REG2_REG_29__SCAN_IN), .ZN(n2645) );
  NAND2_X1 U3460 ( .A1(n3846), .A2(REG0_REG_29__SCAN_IN), .ZN(n2644) );
  OAI211_X1 U3461 ( .C1(n2646), .C2(n3570), .A(n2645), .B(n2644), .ZN(n2647)
         );
  INV_X1 U3462 ( .A(n2647), .ZN(n2648) );
  XNOR2_X1 U3463 ( .A(n3943), .B(n3835), .ZN(n3899) );
  XNOR2_X1 U3464 ( .A(n2650), .B(n3899), .ZN(n2667) );
  INV_X1 U3465 ( .A(n2865), .ZN(n4484) );
  NAND2_X1 U3466 ( .A1(n4484), .A2(n4482), .ZN(n2651) );
  NAND2_X1 U34670 ( .A1(n2652), .A2(IR_REG_31__SCAN_IN), .ZN(n2653) );
  MUX2_X1 U3468 ( .A(IR_REG_31__SCAN_IN), .B(n2653), .S(IR_REG_28__SCAN_IN), 
        .Z(n2654) );
  AND2_X1 U34690 ( .A1(n2655), .A2(n2654), .ZN(n4479) );
  NOR2_X2 U3470 ( .A1(n2660), .A2(n3935), .ZN(n4275) );
  NAND2_X1 U34710 ( .A1(n2656), .A2(REG1_REG_30__SCAN_IN), .ZN(n2659) );
  NAND2_X1 U3472 ( .A1(n3845), .A2(REG2_REG_30__SCAN_IN), .ZN(n2658) );
  NAND2_X1 U34730 ( .A1(n3846), .A2(REG0_REG_30__SCAN_IN), .ZN(n2657) );
  NAND3_X1 U3474 ( .A1(n2659), .A2(n2658), .A3(n2657), .ZN(n3942) );
  NOR2_X2 U34750 ( .A1(n2660), .A2(n4479), .ZN(n4276) );
  XNOR2_X1 U3476 ( .A(n2662), .B(n2661), .ZN(n3960) );
  INV_X1 U34770 ( .A(B_REG_SCAN_IN), .ZN(n2663) );
  OR2_X1 U3478 ( .A1(n3960), .A2(n2663), .ZN(n2664) );
  AND2_X1 U34790 ( .A1(n4276), .A2(n2664), .ZN(n3998) );
  INV_X1 U3480 ( .A(n2739), .ZN(n4483) );
  AOI22_X1 U34810 ( .A1(n3942), .A2(n3998), .B1(n4306), .B2(n3835), .ZN(n2665)
         );
  OAI21_X1 U3482 ( .B1(n4025), .B2(n4296), .A(n2665), .ZN(n2666) );
  AOI21_X1 U34830 ( .B1(n2667), .B2(n4281), .A(n2666), .ZN(n4011) );
  INV_X1 U3484 ( .A(n4481), .ZN(n2671) );
  NAND2_X1 U34850 ( .A1(n2671), .A2(B_REG_SCAN_IN), .ZN(n2674) );
  MUX2_X1 U3486 ( .A(n2674), .B(B_REG_SCAN_IN), .S(n2688), .Z(n2676) );
  NAND2_X1 U34870 ( .A1(n2013), .A2(IR_REG_31__SCAN_IN), .ZN(n2675) );
  NOR4_X1 U3488 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2685) );
  NOR4_X1 U34890 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_10__SCAN_IN), .ZN(n2684) );
  INV_X1 U3490 ( .A(D_REG_26__SCAN_IN), .ZN(n4624) );
  INV_X1 U34910 ( .A(D_REG_2__SCAN_IN), .ZN(n4629) );
  INV_X1 U3492 ( .A(D_REG_21__SCAN_IN), .ZN(n4626) );
  INV_X1 U34930 ( .A(D_REG_6__SCAN_IN), .ZN(n4627) );
  NAND4_X1 U3494 ( .A1(n4624), .A2(n4629), .A3(n4626), .A4(n4627), .ZN(n2682)
         );
  NOR4_X1 U34950 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_17__SCAN_IN), .A4(D_REG_18__SCAN_IN), .ZN(n2680) );
  NOR4_X1 U3496 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n2679) );
  NOR4_X1 U34970 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2678) );
  NOR4_X1 U3498 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2677) );
  NAND4_X1 U34990 ( .A1(n2680), .A2(n2679), .A3(n2678), .A4(n2677), .ZN(n2681)
         );
  NOR4_X1 U3500 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(n2682), 
        .A4(n2681), .ZN(n2683) );
  NAND3_X1 U35010 ( .A1(n2685), .A2(n2684), .A3(n2683), .ZN(n2686) );
  NAND2_X1 U3502 ( .A1(n2694), .A2(n2686), .ZN(n2879) );
  OAI21_X1 U35030 ( .B1(n2690), .B2(n3507), .A(n2689), .ZN(n2923) );
  NAND2_X1 U3504 ( .A1(n2923), .A2(STATE_REG_SCAN_IN), .ZN(n4631) );
  INV_X1 U35050 ( .A(n4631), .ZN(n2691) );
  NAND2_X1 U35060 ( .A1(n2865), .A2(n2739), .ZN(n2883) );
  NAND2_X1 U35070 ( .A1(n2883), .A2(n2882), .ZN(n2922) );
  INV_X1 U35080 ( .A(n2694), .ZN(n2767) );
  OAI22_X1 U35090 ( .A1(n2767), .A2(D_REG_1__SCAN_IN), .B1(n3415), .B2(n4481), 
        .ZN(n2878) );
  AND2_X1 U35100 ( .A1(n4484), .A2(n2739), .ZN(n4613) );
  NAND2_X1 U35110 ( .A1(n4658), .A2(n2693), .ZN(n2890) );
  INV_X1 U35120 ( .A(D_REG_0__SCAN_IN), .ZN(n3417) );
  NAND2_X1 U35130 ( .A1(n2694), .A2(n3417), .ZN(n2698) );
  INV_X1 U35140 ( .A(n3415), .ZN(n2695) );
  NAND2_X1 U35150 ( .A1(n2696), .A2(n2695), .ZN(n2697) );
  AND2_X1 U35160 ( .A1(n3466), .A2(n3956), .ZN(n2840) );
  NAND2_X1 U35170 ( .A1(n3877), .A2(n2840), .ZN(n3027) );
  NAND2_X1 U35180 ( .A1(n2892), .A2(n2868), .ZN(n3026) );
  NAND3_X1 U35190 ( .A1(n3027), .A2(n3026), .A3(n2699), .ZN(n3028) );
  INV_X1 U35200 ( .A(n3736), .ZN(n3034) );
  NAND2_X1 U35210 ( .A1(n2928), .A2(n3034), .ZN(n2700) );
  NAND2_X1 U35220 ( .A1(n3028), .A2(n2700), .ZN(n3069) );
  NAND2_X1 U35230 ( .A1(n3078), .A2(n3737), .ZN(n2701) );
  NAND2_X1 U35240 ( .A1(n3069), .A2(n2701), .ZN(n2703) );
  NAND2_X1 U35250 ( .A1(n2945), .A2(n3072), .ZN(n2702) );
  NAND2_X1 U35260 ( .A1(n3000), .A2(n3953), .ZN(n2704) );
  NAND2_X1 U35270 ( .A1(n3046), .A2(n3119), .ZN(n2705) );
  NAND2_X1 U35280 ( .A1(n3117), .A2(n2705), .ZN(n2708) );
  NAND2_X1 U35290 ( .A1(n2706), .A2(n3952), .ZN(n2707) );
  AND2_X1 U35300 ( .A1(n3051), .A2(n3114), .ZN(n2709) );
  INV_X1 U35310 ( .A(n3884), .ZN(n2710) );
  NAND2_X1 U35320 ( .A1(n3137), .A2(n3951), .ZN(n2711) );
  NAND2_X1 U35330 ( .A1(n3143), .A2(n2711), .ZN(n3155) );
  NAND2_X1 U35340 ( .A1(n3245), .A2(n3184), .ZN(n2712) );
  NAND2_X1 U35350 ( .A1(n3155), .A2(n2712), .ZN(n2715) );
  NAND2_X1 U35360 ( .A1(n2713), .A2(n3950), .ZN(n2714) );
  NAND2_X1 U35370 ( .A1(n2715), .A2(n2714), .ZN(n3201) );
  AND2_X1 U35380 ( .A1(n3233), .A2(n3949), .ZN(n2717) );
  NAND2_X1 U35390 ( .A1(n3627), .A2(n3249), .ZN(n2716) );
  NOR2_X1 U35400 ( .A1(n3264), .A2(n3948), .ZN(n2718) );
  AND2_X1 U35410 ( .A1(n3316), .A2(n4274), .ZN(n2719) );
  OR2_X1 U35420 ( .A1(n2723), .A2(n4249), .ZN(n2722) );
  NAND2_X1 U35430 ( .A1(n3626), .A2(n3272), .ZN(n3295) );
  OR2_X1 U35440 ( .A1(n2719), .A2(n3295), .ZN(n2721) );
  NAND2_X1 U35450 ( .A1(n4299), .A2(n3421), .ZN(n2720) );
  NAND2_X1 U35460 ( .A1(n4245), .A2(n4244), .ZN(n4243) );
  NAND2_X1 U35470 ( .A1(n4228), .A2(n4252), .ZN(n2725) );
  NAND2_X1 U35480 ( .A1(n4243), .A2(n2725), .ZN(n4227) );
  NAND2_X1 U35490 ( .A1(n4238), .A2(n4250), .ZN(n2726) );
  NAND2_X1 U35500 ( .A1(n4213), .A2(n2727), .ZN(n4212) );
  NAND2_X1 U35510 ( .A1(n4221), .A2(n4203), .ZN(n2728) );
  NAND2_X1 U35520 ( .A1(n4187), .A2(n3640), .ZN(n4140) );
  NAND2_X1 U35530 ( .A1(n4205), .A2(n4191), .ZN(n4138) );
  NAND2_X1 U35540 ( .A1(n4140), .A2(n4138), .ZN(n2729) );
  NAND2_X1 U35550 ( .A1(n4167), .A2(n4168), .ZN(n4183) );
  NAND2_X1 U35560 ( .A1(n3946), .A2(n4172), .ZN(n4139) );
  NAND2_X1 U35570 ( .A1(n4129), .A2(n4154), .ZN(n3866) );
  OAI211_X1 U35580 ( .C1(n2729), .C2(n4183), .A(n4139), .B(n3866), .ZN(n2730)
         );
  INV_X1 U35590 ( .A(n4129), .ZN(n4175) );
  NAND2_X1 U35600 ( .A1(n4175), .A2(n4147), .ZN(n3867) );
  NAND2_X1 U35610 ( .A1(n4149), .A2(n4128), .ZN(n2731) );
  INV_X1 U35620 ( .A(n4149), .ZN(n3724) );
  AOI22_X1 U35630 ( .A1(n4125), .A2(n2731), .B1(n3724), .B2(n3650), .ZN(n4108)
         );
  XNOR2_X1 U35640 ( .A(n4100), .B(n4112), .ZN(n4109) );
  NAND2_X1 U35650 ( .A1(n4108), .A2(n4109), .ZN(n4107) );
  NAND2_X1 U35660 ( .A1(n4107), .A2(n2732), .ZN(n4088) );
  NAND2_X1 U35670 ( .A1(n4115), .A2(n3483), .ZN(n2733) );
  INV_X1 U35680 ( .A(n4077), .ZN(n4045) );
  NOR2_X1 U35690 ( .A1(n4047), .A2(n4032), .ZN(n2737) );
  OAI22_X1 U35700 ( .A1(n4028), .A2(n2737), .B1(n3763), .B2(n4022), .ZN(n2747)
         );
  NAND2_X1 U35710 ( .A1(n3843), .A2(n3836), .ZN(n3860) );
  AOI22_X1 U35720 ( .A1(n2747), .A2(n3860), .B1(n3446), .B2(n3944), .ZN(n2738)
         );
  XNOR2_X1 U35730 ( .A(n2738), .B(n3899), .ZN(n4018) );
  XNOR2_X1 U35740 ( .A(n2981), .B(n4482), .ZN(n2740) );
  NAND2_X1 U35750 ( .A1(n2740), .A2(n2865), .ZN(n4303) );
  INV_X1 U35760 ( .A(n4658), .ZN(n4648) );
  NAND2_X1 U35770 ( .A1(n4684), .A2(n4665), .ZN(n4390) );
  NAND2_X1 U35780 ( .A1(n2742), .A2(n2741), .ZN(U3547) );
  INV_X1 U35790 ( .A(REG0_REG_29__SCAN_IN), .ZN(n3569) );
  NAND2_X1 U35800 ( .A1(n4675), .A2(n4665), .ZN(n4471) );
  NAND2_X1 U35810 ( .A1(n2746), .A2(n2745), .ZN(U3515) );
  XNOR2_X1 U3582 ( .A(n2747), .B(n3860), .ZN(n3461) );
  NAND2_X1 U3583 ( .A1(n3943), .A2(n4276), .ZN(n2750) );
  NAND2_X1 U3584 ( .A1(n4047), .A2(n4275), .ZN(n2749) );
  OAI211_X1 U3585 ( .C1(n3435), .C2(n4279), .A(n2750), .B(n2749), .ZN(n2751)
         );
  OAI21_X1 U3586 ( .B1(n3461), .B2(n4668), .A(n3457), .ZN(n2755) );
  OAI21_X1 U3587 ( .B1(n4034), .B2(n3435), .A(n2752), .ZN(n3454) );
  NAND2_X1 U3588 ( .A1(n2754), .A2(n2753), .ZN(U3514) );
  NAND2_X1 U3589 ( .A1(n4684), .A2(n4653), .ZN(n4395) );
  NAND2_X1 U3590 ( .A1(n2757), .A2(n2756), .ZN(U3546) );
  INV_X2 U3591 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X2 U3592 ( .A(n3955), .ZN(U4043) );
  MUX2_X1 U3593 ( .A(n2758), .B(n3063), .S(STATE_REG_SCAN_IN), .Z(n2759) );
  INV_X1 U3594 ( .A(n2759), .ZN(U3344) );
  INV_X1 U3595 ( .A(DATAI_21_), .ZN(n2761) );
  NAND2_X1 U3596 ( .A1(n3931), .A2(STATE_REG_SCAN_IN), .ZN(n2760) );
  OAI21_X1 U3597 ( .B1(STATE_REG_SCAN_IN), .B2(n2761), .A(n2760), .ZN(U3331)
         );
  INV_X1 U3598 ( .A(DATAI_26_), .ZN(n3489) );
  NAND2_X1 U3599 ( .A1(n3415), .A2(STATE_REG_SCAN_IN), .ZN(n2762) );
  OAI21_X1 U3600 ( .B1(STATE_REG_SCAN_IN), .B2(n3489), .A(n2762), .ZN(U3326)
         );
  INV_X1 U3601 ( .A(DATAI_31_), .ZN(n2766) );
  OR4_X1 U3602 ( .A1(n2764), .A2(IR_REG_30__SCAN_IN), .A3(n2763), .A4(U3149), 
        .ZN(n2765) );
  OAI21_X1 U3603 ( .B1(STATE_REG_SCAN_IN), .B2(n2766), .A(n2765), .ZN(U3321)
         );
  INV_X1 U3604 ( .A(D_REG_1__SCAN_IN), .ZN(n2769) );
  NOR3_X1 U3605 ( .A1(n4631), .A2(n3415), .A3(n4481), .ZN(n2768) );
  AOI21_X1 U3606 ( .B1(n4628), .B2(n2769), .A(n2768), .ZN(U3459) );
  INV_X1 U3607 ( .A(n3960), .ZN(n4480) );
  INV_X1 U3608 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2770) );
  AOI21_X1 U3609 ( .B1(n4480), .B2(n2770), .A(n3935), .ZN(n3963) );
  OAI21_X1 U3610 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4480), .A(n3963), .ZN(n2771)
         );
  MUX2_X1 U3611 ( .A(n2771), .B(n3963), .S(IR_REG_0__SCAN_IN), .Z(n2780) );
  OR2_X1 U3612 ( .A1(n2923), .A2(U3149), .ZN(n3940) );
  INV_X1 U3613 ( .A(n3940), .ZN(n2772) );
  OR2_X1 U3614 ( .A1(n2887), .A2(n2772), .ZN(n2776) );
  NAND2_X1 U3615 ( .A1(n2882), .A2(n2923), .ZN(n2773) );
  AND2_X1 U3616 ( .A1(n3850), .A2(n2773), .ZN(n2774) );
  INV_X1 U3617 ( .A(n2791), .ZN(n2779) );
  INV_X1 U3618 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2871) );
  NAND3_X1 U3619 ( .A1(n4584), .A2(IR_REG_0__SCAN_IN), .A3(n2871), .ZN(n2778)
         );
  INV_X1 U3620 ( .A(n2774), .ZN(n2775) );
  AOI22_X1 U3621 ( .A1(n4595), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n2777) );
  OAI211_X1 U3622 ( .C1(n2780), .C2(n2779), .A(n2778), .B(n2777), .ZN(U3240)
         );
  NOR2_X1 U3623 ( .A1(n4595), .A2(U4043), .ZN(U3148) );
  INV_X1 U3624 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n3526) );
  NAND2_X1 U3625 ( .A1(U4043), .A2(n3737), .ZN(n2781) );
  OAI21_X1 U3626 ( .B1(U4043), .B2(n3526), .A(n2781), .ZN(U3553) );
  INV_X1 U3627 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n3500) );
  NAND2_X1 U3628 ( .A1(U4043), .A2(n3114), .ZN(n2782) );
  OAI21_X1 U3629 ( .B1(U4043), .B2(n3500), .A(n2782), .ZN(U3556) );
  INV_X1 U3630 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n3525) );
  NAND2_X1 U3631 ( .A1(n4185), .A2(U4043), .ZN(n2783) );
  OAI21_X1 U3632 ( .B1(U4043), .B2(n3525), .A(n2783), .ZN(U3567) );
  AND2_X1 U3633 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n2796)
         );
  XNOR2_X1 U3634 ( .A(n2797), .B(n2796), .ZN(n2795) );
  INV_X1 U3635 ( .A(n4595), .ZN(n4563) );
  INV_X1 U3636 ( .A(ADDR_REG_1__SCAN_IN), .ZN(n2785) );
  INV_X1 U3637 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2784) );
  OAI22_X1 U3638 ( .A1(n4563), .A2(n2785), .B1(STATE_REG_SCAN_IN), .B2(n2784), 
        .ZN(n2786) );
  AOI21_X1 U3639 ( .B1(n4494), .B2(n4559), .A(n2786), .ZN(n2794) );
  AND2_X1 U3640 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3961)
         );
  NOR2_X1 U3641 ( .A1(n3960), .A2(n3935), .ZN(n2790) );
  NAND2_X1 U3642 ( .A1(n2792), .A2(n3961), .ZN(n2804) );
  OAI211_X1 U3643 ( .C1(n3961), .C2(n2792), .A(n4586), .B(n2804), .ZN(n2793)
         );
  OAI211_X1 U3644 ( .C1(n4590), .C2(n2795), .A(n2794), .B(n2793), .ZN(U3241)
         );
  NAND2_X1 U3645 ( .A1(n2797), .A2(n2796), .ZN(n2799) );
  NAND2_X1 U3646 ( .A1(n4494), .A2(REG1_REG_1__SCAN_IN), .ZN(n2798) );
  INV_X1 U3647 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3040) );
  XNOR2_X1 U3648 ( .A(n4493), .B(n3040), .ZN(n3964) );
  NAND2_X1 U3649 ( .A1(n3965), .A2(n3964), .ZN(n2801) );
  NAND2_X1 U3650 ( .A1(n4493), .A2(REG1_REG_2__SCAN_IN), .ZN(n2800) );
  NAND2_X2 U3651 ( .A1(n2801), .A2(n2800), .ZN(n2812) );
  XNOR2_X1 U3652 ( .A(n2811), .B(REG1_REG_3__SCAN_IN), .ZN(n2810) );
  INV_X1 U3653 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2802) );
  NAND2_X1 U3654 ( .A1(n4494), .A2(REG2_REG_1__SCAN_IN), .ZN(n2803) );
  NAND2_X1 U3655 ( .A1(n4493), .A2(REG2_REG_2__SCAN_IN), .ZN(n2805) );
  INV_X1 U3656 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3079) );
  XNOR2_X1 U3657 ( .A(n2817), .B(n3079), .ZN(n2808) );
  AOI22_X1 U3658 ( .A1(n4595), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n2806) );
  OAI21_X1 U3659 ( .B1(n4604), .B2(n2331), .A(n2806), .ZN(n2807) );
  AOI21_X1 U3660 ( .B1(n4586), .B2(n2808), .A(n2807), .ZN(n2809) );
  OAI21_X1 U3661 ( .B1(n2810), .B2(n4590), .A(n2809), .ZN(U3243) );
  NAND2_X1 U3662 ( .A1(n2811), .A2(REG1_REG_3__SCAN_IN), .ZN(n2814) );
  NAND2_X1 U3663 ( .A1(n2812), .A2(n4492), .ZN(n2813) );
  INV_X1 U3664 ( .A(n4529), .ZN(n2821) );
  INV_X1 U3665 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4679) );
  MUX2_X1 U3666 ( .A(REG1_REG_5__SCAN_IN), .B(n4679), .S(n2835), .Z(n2832) );
  NOR2_X2 U3667 ( .A1(n2833), .A2(n2832), .ZN(n2831) );
  INV_X1 U3668 ( .A(n2835), .ZN(n4491) );
  NOR2_X2 U3669 ( .A1(n2831), .A2(n2816), .ZN(n2850) );
  XNOR2_X1 U3670 ( .A(n2852), .B(REG1_REG_6__SCAN_IN), .ZN(n2827) );
  NAND2_X1 U3671 ( .A1(n2817), .A2(REG2_REG_3__SCAN_IN), .ZN(n2820) );
  NAND2_X1 U3672 ( .A1(n2818), .A2(n4492), .ZN(n2819) );
  NAND2_X1 U3673 ( .A1(n2820), .A2(n2819), .ZN(n2822) );
  XNOR2_X1 U3674 ( .A(n2822), .B(n2821), .ZN(n4527) );
  INV_X1 U3675 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3578) );
  MUX2_X1 U3676 ( .A(REG2_REG_5__SCAN_IN), .B(n3578), .S(n2835), .Z(n2829) );
  XOR2_X1 U3677 ( .A(n2855), .B(REG2_REG_6__SCAN_IN), .Z(n2825) );
  NAND2_X1 U3678 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3020) );
  NAND2_X1 U3679 ( .A1(n4595), .A2(ADDR_REG_6__SCAN_IN), .ZN(n2823) );
  OAI211_X1 U3680 ( .C1(n4604), .C2(n2062), .A(n3020), .B(n2823), .ZN(n2824)
         );
  AOI21_X1 U3681 ( .B1(n2825), .B2(n4586), .A(n2824), .ZN(n2826) );
  OAI21_X1 U3682 ( .B1(n2827), .B2(n4590), .A(n2826), .ZN(U3246) );
  AOI211_X1 U3683 ( .C1(n2830), .C2(n2829), .A(n4596), .B(n2828), .ZN(n2838)
         );
  AOI211_X1 U3684 ( .C1(n2833), .C2(n2832), .A(n4590), .B(n2831), .ZN(n2837)
         );
  NOR2_X1 U3685 ( .A1(STATE_REG_SCAN_IN), .A2(n2450), .ZN(n2962) );
  AOI21_X1 U3686 ( .B1(n4595), .B2(ADDR_REG_5__SCAN_IN), .A(n2962), .ZN(n2834)
         );
  OAI21_X1 U3687 ( .B1(n4604), .B2(n2835), .A(n2834), .ZN(n2836) );
  OR3_X1 U3688 ( .A1(n2838), .A2(n2837), .A3(n2836), .ZN(U3245) );
  INV_X1 U3689 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n3558) );
  NAND2_X1 U3690 ( .A1(n4100), .A2(U4043), .ZN(n2839) );
  OAI21_X1 U3691 ( .B1(U4043), .B2(n3558), .A(n2839), .ZN(U3572) );
  OR2_X1 U3692 ( .A1(n2840), .A2(n3877), .ZN(n2841) );
  NAND2_X1 U3693 ( .A1(n3027), .A2(n2841), .ZN(n2983) );
  NAND2_X1 U3694 ( .A1(n3956), .A2(n4275), .ZN(n2843) );
  NAND2_X1 U3695 ( .A1(n2892), .A2(n4306), .ZN(n2842) );
  OAI211_X1 U3696 ( .C1(n2928), .C2(n4298), .A(n2843), .B(n2842), .ZN(n2844)
         );
  INV_X1 U3697 ( .A(n2844), .ZN(n2847) );
  XNOR2_X1 U3698 ( .A(n3877), .B(n3784), .ZN(n2845) );
  NAND2_X1 U3699 ( .A1(n2845), .A2(n4281), .ZN(n2846) );
  OAI211_X1 U3700 ( .C1(n2983), .C2(n4303), .A(n2847), .B(n2846), .ZN(n2985)
         );
  OAI21_X1 U3701 ( .B1(n2898), .B2(n2864), .A(n3038), .ZN(n2989) );
  OAI22_X1 U3702 ( .A1(n2983), .A2(n4648), .B1(n2989), .B2(n4661), .ZN(n2848)
         );
  NOR2_X1 U3703 ( .A1(n2985), .A2(n2848), .ZN(n4647) );
  NAND2_X1 U3704 ( .A1(n4681), .A2(REG1_REG_1__SCAN_IN), .ZN(n2849) );
  OAI21_X1 U3705 ( .B1(n4647), .B2(n4681), .A(n2849), .ZN(U3519) );
  INV_X1 U3706 ( .A(n2850), .ZN(n2851) );
  AOI22_X2 U3707 ( .A1(n2852), .A2(REG1_REG_6__SCAN_IN), .B1(n4490), .B2(n2851), .ZN(n2970) );
  INV_X1 U3708 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4682) );
  XNOR2_X1 U3709 ( .A(n4489), .B(n4682), .ZN(n2853) );
  XNOR2_X1 U3710 ( .A(n2970), .B(n2853), .ZN(n2860) );
  INV_X1 U3711 ( .A(n4489), .ZN(n2971) );
  AND2_X1 U3712 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3105) );
  AOI21_X1 U3713 ( .B1(n4595), .B2(ADDR_REG_7__SCAN_IN), .A(n3105), .ZN(n2854)
         );
  OAI21_X1 U3714 ( .B1(n4604), .B2(n2971), .A(n2854), .ZN(n2859) );
  INV_X1 U3715 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3142) );
  MUX2_X1 U3716 ( .A(n3142), .B(REG2_REG_7__SCAN_IN), .S(n4489), .Z(n2856) );
  AOI211_X1 U3717 ( .C1(n2857), .C2(n2856), .A(n4596), .B(n2967), .ZN(n2858)
         );
  AOI211_X1 U3718 ( .C1(n2860), .C2(n4584), .A(n2859), .B(n2858), .ZN(n2861)
         );
  INV_X1 U3719 ( .A(n2861), .ZN(U3247) );
  INV_X1 U3720 ( .A(n2981), .ZN(n2863) );
  OAI22_X1 U3721 ( .A1(n2864), .A2(n3431), .B1(n3468), .B2(n3337), .ZN(n2866)
         );
  XNOR2_X1 U3722 ( .A(n2866), .B(n3433), .ZN(n2907) );
  BUF_X1 U3723 ( .A(n2956), .Z(n3263) );
  AOI22_X1 U3724 ( .A1(n2868), .A2(n2936), .B1(n2892), .B2(n3263), .ZN(n2908)
         );
  XNOR2_X1 U3725 ( .A(n2907), .B(n2908), .ZN(n2912) );
  NAND2_X1 U3726 ( .A1(n3956), .A2(n2956), .ZN(n2870) );
  NAND2_X1 U3727 ( .A1(n3466), .A2(n3393), .ZN(n2869) );
  INV_X1 U3728 ( .A(IR_REG_0__SCAN_IN), .ZN(n2872) );
  NOR2_X1 U3729 ( .A1(n2862), .A2(n2872), .ZN(n2873) );
  AOI21_X1 U3730 ( .B1(n3466), .B2(n3263), .A(n2873), .ZN(n2875) );
  NAND2_X1 U3731 ( .A1(n2936), .A2(n3956), .ZN(n2874) );
  NAND2_X1 U3732 ( .A1(n2875), .A2(n2874), .ZN(n3462) );
  NAND2_X1 U3733 ( .A1(n3463), .A2(n3462), .ZN(n2877) );
  NAND2_X1 U3734 ( .A1(n2308), .A2(n3396), .ZN(n2876) );
  NAND2_X1 U3735 ( .A1(n2877), .A2(n2876), .ZN(n2911) );
  XNOR2_X1 U3736 ( .A(n2912), .B(n2911), .ZN(n2895) );
  INV_X1 U3737 ( .A(n2878), .ZN(n2977) );
  NAND3_X1 U3738 ( .A1(n2977), .A2(n2880), .A3(n2879), .ZN(n2891) );
  INV_X1 U3739 ( .A(n2887), .ZN(n2881) );
  INV_X1 U3740 ( .A(n2889), .ZN(n2885) );
  AOI21_X1 U3741 ( .B1(n2883), .B2(n2901), .A(n2882), .ZN(n2884) );
  NAND2_X2 U3742 ( .A1(n2885), .A2(n2884), .ZN(n3782) );
  NOR2_X1 U3743 ( .A1(n2889), .A2(n2302), .ZN(n2886) );
  INV_X1 U3744 ( .A(n2928), .ZN(n3954) );
  AOI22_X1 U3745 ( .A1(n3749), .A2(n3956), .B1(n3750), .B2(n3954), .ZN(n2894)
         );
  INV_X1 U3746 ( .A(n2890), .ZN(n2888) );
  NAND2_X1 U3747 ( .A1(n2891), .A2(n2890), .ZN(n2924) );
  NAND2_X1 U3748 ( .A1(n2924), .A2(n2303), .ZN(n3735) );
  AOI22_X1 U3749 ( .A1(n3754), .A2(n2892), .B1(REG3_REG_1__SCAN_IN), .B2(n3735), .ZN(n2893) );
  OAI211_X1 U3750 ( .C1(n2895), .C2(n3782), .A(n2894), .B(n2893), .ZN(U3219)
         );
  INV_X1 U3751 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n3557) );
  NAND2_X1 U3752 ( .A1(n2896), .A2(U4043), .ZN(n2897) );
  OAI21_X1 U3753 ( .B1(U4043), .B2(n3557), .A(n2897), .ZN(U3573) );
  NAND2_X1 U3754 ( .A1(n2898), .A2(n3956), .ZN(n3786) );
  NAND2_X1 U3755 ( .A1(n3786), .A2(n3784), .ZN(n4619) );
  NAND2_X1 U3756 ( .A1(n4303), .A2(n4309), .ZN(n2900) );
  NOR2_X1 U3757 ( .A1(n3468), .A2(n4298), .ZN(n2899) );
  AOI21_X1 U3758 ( .B1(n4619), .B2(n2900), .A(n2899), .ZN(n4614) );
  AND2_X1 U3759 ( .A1(n3466), .A2(n2901), .ZN(n4617) );
  AOI21_X1 U3760 ( .B1(n4619), .B2(n4658), .A(n4617), .ZN(n2902) );
  AND2_X1 U3761 ( .A1(n4614), .A2(n2902), .ZN(n4645) );
  NAND2_X1 U3762 ( .A1(n4681), .A2(REG1_REG_0__SCAN_IN), .ZN(n2903) );
  OAI21_X1 U3763 ( .B1(n4681), .B2(n4645), .A(n2903), .ZN(U3518) );
  INV_X2 U3764 ( .A(n3392), .ZN(n3432) );
  INV_X1 U3765 ( .A(n2936), .ZN(n2959) );
  OAI22_X1 U3766 ( .A1(n3072), .A2(n3432), .B1(n2945), .B2(n2959), .ZN(n2938)
         );
  NAND2_X1 U3767 ( .A1(n3737), .A2(n3392), .ZN(n2905) );
  NAND2_X1 U3768 ( .A1(n3078), .A2(n3393), .ZN(n2904) );
  NAND2_X1 U3769 ( .A1(n2905), .A2(n2904), .ZN(n2906) );
  XOR2_X1 U3770 ( .A(n2938), .B(n2937), .Z(n2921) );
  INV_X1 U3771 ( .A(n2907), .ZN(n2909) );
  NOR2_X1 U3772 ( .A1(n2909), .A2(n2908), .ZN(n2910) );
  NAND2_X1 U3773 ( .A1(n3736), .A2(n3393), .ZN(n2913) );
  OAI21_X1 U3774 ( .B1(n2928), .B2(n3337), .A(n2913), .ZN(n2914) );
  XNOR2_X1 U3775 ( .A(n2914), .B(n3433), .ZN(n2917) );
  NAND2_X1 U3776 ( .A1(n3736), .A2(n3392), .ZN(n2915) );
  NOR2_X1 U3777 ( .A1(n2917), .A2(n2916), .ZN(n2918) );
  AOI21_X1 U3778 ( .B1(n2917), .B2(n2916), .A(n2918), .ZN(n3732) );
  NAND2_X1 U3779 ( .A1(n3729), .A2(n3732), .ZN(n3731) );
  INV_X1 U3780 ( .A(n2918), .ZN(n2919) );
  OAI21_X1 U3781 ( .B1(n2921), .B2(n2920), .A(n2941), .ZN(n2930) );
  INV_X1 U3782 ( .A(n3782), .ZN(n3733) );
  AOI22_X1 U3783 ( .A1(n3750), .A2(n3953), .B1(n3078), .B2(n3754), .ZN(n2927)
         );
  NAND4_X1 U3784 ( .A1(n2924), .A2(n2862), .A3(n2923), .A4(n2922), .ZN(n2925)
         );
  NAND2_X1 U3785 ( .A1(n2925), .A2(STATE_REG_SCAN_IN), .ZN(n3752) );
  MUX2_X1 U3786 ( .A(n3752), .B(STATE_REG_SCAN_IN), .S(REG3_REG_3__SCAN_IN), 
        .Z(n2926) );
  OAI211_X1 U3787 ( .C1(n2928), .C2(n3777), .A(n2927), .B(n2926), .ZN(n2929)
         );
  AOI21_X1 U3788 ( .B1(n2930), .B2(n3733), .A(n2929), .ZN(n2931) );
  INV_X1 U3789 ( .A(n2931), .ZN(U3215) );
  NAND2_X1 U3790 ( .A1(n3000), .A2(n3393), .ZN(n2934) );
  NAND2_X1 U3791 ( .A1(n3953), .A2(n3392), .ZN(n2933) );
  NAND2_X1 U3792 ( .A1(n2934), .A2(n2933), .ZN(n2935) );
  INV_X1 U3793 ( .A(n2937), .ZN(n2940) );
  INV_X1 U3794 ( .A(n2938), .ZN(n2939) );
  NAND2_X1 U3795 ( .A1(n2940), .A2(n2939), .ZN(n2943) );
  NAND2_X1 U3796 ( .A1(n2955), .A2(n3733), .ZN(n2950) );
  AOI21_X1 U3797 ( .B1(n2941), .B2(n2943), .A(n2942), .ZN(n2949) );
  NAND2_X1 U3798 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n4530) );
  OAI21_X1 U3799 ( .B1(n3775), .B2(n2944), .A(n4530), .ZN(n2947) );
  OAI22_X1 U3800 ( .A1(n3046), .A2(n3776), .B1(n3777), .B2(n2945), .ZN(n2946)
         );
  AOI211_X1 U3801 ( .C1(n3001), .C2(n3780), .A(n2947), .B(n2946), .ZN(n2948)
         );
  OAI21_X1 U3802 ( .B1(n2950), .B2(n2949), .A(n2948), .ZN(U3227) );
  INV_X1 U3803 ( .A(n2952), .ZN(n2953) );
  OR2_X1 U3804 ( .A1(n3119), .A2(n3431), .ZN(n2957) );
  XNOR2_X1 U3805 ( .A(n2958), .B(n3396), .ZN(n3008) );
  OR2_X1 U3806 ( .A1(n3119), .A2(n3432), .ZN(n2960) );
  OAI21_X1 U3807 ( .B1(n3046), .B2(n3436), .A(n2960), .ZN(n3009) );
  XNOR2_X1 U3808 ( .A(n3008), .B(n3009), .ZN(n3006) );
  XNOR2_X1 U3809 ( .A(n3007), .B(n3006), .ZN(n2965) );
  AOI22_X1 U3810 ( .A1(n3749), .A2(n3953), .B1(n3750), .B2(n3114), .ZN(n2964)
         );
  NOR2_X1 U3811 ( .A1(n3775), .A2(n3119), .ZN(n2961) );
  AOI211_X1 U3812 ( .C1(n3121), .C2(n3780), .A(n2962), .B(n2961), .ZN(n2963)
         );
  OAI211_X1 U3813 ( .C1(n2965), .C2(n3782), .A(n2964), .B(n2963), .ZN(U3224)
         );
  XNOR2_X1 U3814 ( .A(n3056), .B(REG2_REG_8__SCAN_IN), .ZN(n2976) );
  AND2_X1 U3815 ( .A1(U3149), .A2(REG3_REG_8__SCAN_IN), .ZN(n2969) );
  NOR2_X1 U3816 ( .A1(n4604), .A2(n3063), .ZN(n2968) );
  AOI211_X1 U3817 ( .C1(n4595), .C2(ADDR_REG_8__SCAN_IN), .A(n2969), .B(n2968), 
        .ZN(n2975) );
  INV_X1 U3818 ( .A(n3063), .ZN(n3055) );
  OAI211_X1 U3819 ( .C1(n2973), .C2(REG1_REG_8__SCAN_IN), .A(n3062), .B(n4584), 
        .ZN(n2974) );
  OAI211_X1 U3820 ( .C1(n2976), .C2(n4596), .A(n2975), .B(n2974), .ZN(U3248)
         );
  NAND3_X1 U3821 ( .A1(n2979), .A2(n2978), .A3(n2977), .ZN(n2980) );
  NAND2_X1 U3822 ( .A1(n4289), .A2(n2865), .ZN(n4192) );
  OR2_X1 U3823 ( .A1(n2981), .A2(n2865), .ZN(n3089) );
  INV_X1 U3824 ( .A(n3089), .ZN(n2982) );
  INV_X1 U3825 ( .A(n2983), .ZN(n2984) );
  AOI22_X1 U3826 ( .A1(n4620), .A2(n2984), .B1(REG3_REG_1__SCAN_IN), .B2(n4618), .ZN(n2988) );
  MUX2_X1 U3827 ( .A(REG2_REG_1__SCAN_IN), .B(n2985), .S(n4289), .Z(n2986) );
  INV_X1 U3828 ( .A(n2986), .ZN(n2987) );
  OAI211_X1 U3829 ( .C1(n4317), .C2(n2989), .A(n2988), .B(n2987), .ZN(U3289)
         );
  XNOR2_X1 U3830 ( .A(n3883), .B(n2991), .ZN(n2998) );
  NAND2_X1 U3831 ( .A1(n2992), .A2(n3883), .ZN(n2993) );
  NAND2_X1 U3832 ( .A1(n2994), .A2(n2993), .ZN(n3003) );
  AOI22_X1 U3833 ( .A1(n3952), .A2(n4276), .B1(n4275), .B2(n3737), .ZN(n2996)
         );
  NAND2_X1 U3834 ( .A1(n3000), .A2(n4306), .ZN(n2995) );
  OAI211_X1 U3835 ( .C1(n3003), .C2(n4303), .A(n2996), .B(n2995), .ZN(n2997)
         );
  AOI21_X1 U3836 ( .B1(n2998), .B2(n4281), .A(n2997), .ZN(n4655) );
  INV_X1 U3837 ( .A(n3076), .ZN(n2999) );
  AOI211_X1 U3838 ( .C1(n3000), .C2(n2999), .A(n4661), .B(n3120), .ZN(n4657)
         );
  AOI22_X1 U3839 ( .A1(n4657), .A2(n2865), .B1(n4618), .B2(n3001), .ZN(n3002)
         );
  AND2_X1 U3840 ( .A1(n4655), .A2(n3002), .ZN(n3005) );
  INV_X1 U3841 ( .A(n3003), .ZN(n4659) );
  AOI22_X1 U3842 ( .A1(n4659), .A2(n4620), .B1(REG2_REG_4__SCAN_IN), .B2(n4623), .ZN(n3004) );
  OAI21_X1 U3843 ( .B1(n3005), .B2(n4623), .A(n3004), .ZN(U3286) );
  NAND2_X1 U3844 ( .A1(n3007), .A2(n3006), .ZN(n3012) );
  INV_X1 U3845 ( .A(n3008), .ZN(n3010) );
  NAND2_X1 U3846 ( .A1(n3051), .A2(n3393), .ZN(n3014) );
  NAND2_X1 U3847 ( .A1(n3114), .A2(n3392), .ZN(n3013) );
  NAND2_X1 U3848 ( .A1(n3014), .A2(n3013), .ZN(n3015) );
  XNOR2_X1 U3849 ( .A(n3015), .B(n3396), .ZN(n3017) );
  AOI22_X1 U3850 ( .A1(n3399), .A2(n3114), .B1(n3051), .B2(n3392), .ZN(n3016)
         );
  NOR2_X1 U3851 ( .A1(n3017), .A2(n3016), .ZN(n3101) );
  INV_X1 U3852 ( .A(n3101), .ZN(n3018) );
  NAND2_X1 U3853 ( .A1(n3017), .A2(n3016), .ZN(n3100) );
  NAND2_X1 U3854 ( .A1(n3018), .A2(n3100), .ZN(n3019) );
  XNOR2_X1 U3855 ( .A(n2041), .B(n3019), .ZN(n3025) );
  OAI21_X1 U3856 ( .B1(n3775), .B2(n3021), .A(n3020), .ZN(n3023) );
  OAI22_X1 U3857 ( .A1(n3046), .A2(n3777), .B1(n3776), .B2(n3185), .ZN(n3022)
         );
  AOI211_X1 U3858 ( .C1(n3091), .C2(n3780), .A(n3023), .B(n3022), .ZN(n3024)
         );
  OAI21_X1 U3859 ( .B1(n3025), .B2(n3782), .A(n3024), .ZN(U3236) );
  NAND2_X1 U3860 ( .A1(n3027), .A2(n3026), .ZN(n3030) );
  INV_X1 U3861 ( .A(n3028), .ZN(n3029) );
  AOI21_X1 U3862 ( .B1(n3880), .B2(n3030), .A(n3029), .ZN(n4605) );
  OAI21_X1 U3863 ( .B1(n3880), .B2(n3032), .A(n3031), .ZN(n3037) );
  AOI22_X1 U3864 ( .A1(n2868), .A2(n4275), .B1(n4276), .B2(n3737), .ZN(n3033)
         );
  OAI21_X1 U3865 ( .B1(n3034), .B2(n4279), .A(n3033), .ZN(n3036) );
  NOR2_X1 U3866 ( .A1(n4605), .A2(n4303), .ZN(n3035) );
  AOI211_X1 U3867 ( .C1(n4281), .C2(n3037), .A(n3036), .B(n3035), .ZN(n4612)
         );
  OAI21_X1 U3868 ( .B1(n4605), .B2(n4648), .A(n4612), .ZN(n3085) );
  NAND2_X1 U3869 ( .A1(n3038), .A2(n3736), .ZN(n3039) );
  NAND2_X1 U3870 ( .A1(n3077), .A2(n3039), .ZN(n4606) );
  OAI22_X1 U3871 ( .A1(n4395), .A2(n4606), .B1(n4684), .B2(n3040), .ZN(n3041)
         );
  AOI21_X1 U3872 ( .B1(n3085), .B2(n4684), .A(n3041), .ZN(n3042) );
  INV_X1 U3873 ( .A(n3042), .ZN(U3520) );
  INV_X1 U3874 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n3527) );
  NAND2_X1 U3875 ( .A1(n4077), .A2(U4043), .ZN(n3043) );
  OAI21_X1 U3876 ( .B1(n3527), .B2(U4043), .A(n3043), .ZN(U3575) );
  NAND2_X1 U3877 ( .A1(n3804), .A2(n3800), .ZN(n3876) );
  XOR2_X1 U3878 ( .A(n3044), .B(n3876), .Z(n3095) );
  XNOR2_X1 U3879 ( .A(n3045), .B(n3876), .ZN(n3049) );
  OAI22_X1 U3880 ( .A1(n3046), .A2(n4296), .B1(n3185), .B2(n4298), .ZN(n3047)
         );
  AOI21_X1 U3881 ( .B1(n3051), .B2(n4306), .A(n3047), .ZN(n3048) );
  OAI21_X1 U3882 ( .B1(n3049), .B2(n4309), .A(n3048), .ZN(n3088) );
  AOI21_X1 U3883 ( .B1(n3095), .B2(n4665), .A(n3088), .ZN(n3131) );
  INV_X1 U3884 ( .A(n3138), .ZN(n3050) );
  AOI21_X1 U3885 ( .B1(n3051), .B2(n3118), .A(n3050), .ZN(n3129) );
  AOI22_X1 U3886 ( .A1(n3129), .A2(n4372), .B1(n4681), .B2(REG1_REG_6__SCAN_IN), .ZN(n3052) );
  OAI21_X1 U3887 ( .B1(n3131), .B2(n4681), .A(n3052), .ZN(U3524) );
  INV_X1 U3888 ( .A(n3053), .ZN(n3054) );
  INV_X1 U3889 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3057) );
  MUX2_X1 U3890 ( .A(n3057), .B(REG2_REG_9__SCAN_IN), .S(n4488), .Z(n3058) );
  AOI211_X1 U3891 ( .C1(n2053), .C2(n3058), .A(n4596), .B(n3162), .ZN(n3061)
         );
  INV_X1 U3892 ( .A(n4488), .ZN(n3165) );
  NAND2_X1 U3893 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n3247) );
  NAND2_X1 U3894 ( .A1(n4595), .A2(ADDR_REG_9__SCAN_IN), .ZN(n3059) );
  OAI211_X1 U3895 ( .C1(n4604), .C2(n3165), .A(n3247), .B(n3059), .ZN(n3060)
         );
  NOR2_X1 U3896 ( .A1(n3061), .A2(n3060), .ZN(n3068) );
  XOR2_X1 U3897 ( .A(REG1_REG_9__SCAN_IN), .B(n4488), .Z(n3065) );
  OAI211_X1 U3898 ( .C1(n3066), .C2(n3065), .A(n3166), .B(n4584), .ZN(n3067)
         );
  NAND2_X1 U3899 ( .A1(n3068), .A2(n3067), .ZN(U3249) );
  XNOR2_X1 U3900 ( .A(n3069), .B(n3882), .ZN(n4649) );
  INV_X1 U3901 ( .A(n4620), .ZN(n4294) );
  XNOR2_X1 U3902 ( .A(n3070), .B(n3882), .ZN(n3074) );
  AOI22_X1 U3903 ( .A1(n4275), .A2(n3954), .B1(n3953), .B2(n4276), .ZN(n3071)
         );
  OAI21_X1 U3904 ( .B1(n3072), .B2(n4279), .A(n3071), .ZN(n3073) );
  AOI21_X1 U3905 ( .B1(n3074), .B2(n4281), .A(n3073), .ZN(n3075) );
  OAI21_X1 U3906 ( .B1(n4649), .B2(n4303), .A(n3075), .ZN(n4650) );
  NAND2_X1 U3907 ( .A1(n4650), .A2(n4289), .ZN(n3082) );
  AOI21_X1 U3908 ( .B1(n3078), .B2(n3077), .A(n3076), .ZN(n4652) );
  OAI22_X1 U3909 ( .A1(n4289), .A2(n3079), .B1(REG3_REG_3__SCAN_IN), .B2(n4287), .ZN(n3080) );
  AOI21_X1 U3910 ( .B1(n4608), .B2(n4652), .A(n3080), .ZN(n3081) );
  OAI211_X1 U3911 ( .C1(n4649), .C2(n4294), .A(n3082), .B(n3081), .ZN(U3287)
         );
  INV_X1 U3912 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3083) );
  OAI22_X1 U3913 ( .A1(n4476), .A2(n4606), .B1(n4675), .B2(n3083), .ZN(n3084)
         );
  AOI21_X1 U3914 ( .B1(n3085), .B2(n4675), .A(n3084), .ZN(n3086) );
  INV_X1 U3915 ( .A(n3086), .ZN(U3471) );
  INV_X1 U3916 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n3499) );
  NAND2_X1 U3917 ( .A1(n4047), .A2(U4043), .ZN(n3087) );
  OAI21_X1 U3918 ( .B1(U4043), .B2(n3499), .A(n3087), .ZN(U3577) );
  INV_X1 U3919 ( .A(n3088), .ZN(n3097) );
  NAND2_X1 U3920 ( .A1(n4303), .A2(n3089), .ZN(n3090) );
  INV_X1 U3921 ( .A(n4242), .ZN(n4030) );
  INV_X1 U3922 ( .A(n3129), .ZN(n3093) );
  AOI22_X1 U3923 ( .A1(n4623), .A2(REG2_REG_6__SCAN_IN), .B1(n3091), .B2(n4618), .ZN(n3092) );
  OAI21_X1 U3924 ( .B1(n3093), .B2(n4317), .A(n3092), .ZN(n3094) );
  AOI21_X1 U3925 ( .B1(n3095), .B2(n4030), .A(n3094), .ZN(n3096) );
  OAI21_X1 U3926 ( .B1(n3097), .B2(n4623), .A(n3096), .ZN(U3284) );
  AOI22_X1 U3927 ( .A1(n3951), .A2(n3399), .B1(n3137), .B2(n3263), .ZN(n3171)
         );
  NAND2_X1 U3928 ( .A1(n3137), .A2(n3393), .ZN(n3098) );
  OAI21_X1 U3929 ( .B1(n3185), .B2(n3432), .A(n3098), .ZN(n3099) );
  XNOR2_X1 U3930 ( .A(n3099), .B(n3433), .ZN(n3173) );
  XOR2_X1 U3931 ( .A(n3171), .B(n3173), .Z(n3103) );
  AOI211_X1 U3932 ( .C1(n3103), .C2(n3102), .A(n3782), .B(n2044), .ZN(n3109)
         );
  INV_X1 U3933 ( .A(n3104), .ZN(n3141) );
  AOI22_X1 U3934 ( .A1(n3750), .A2(n3950), .B1(n3749), .B2(n3114), .ZN(n3107)
         );
  AOI21_X1 U3935 ( .B1(n3754), .B2(n3137), .A(n3105), .ZN(n3106) );
  OAI211_X1 U3936 ( .C1(n3752), .C2(n3141), .A(n3107), .B(n3106), .ZN(n3108)
         );
  OR2_X1 U3937 ( .A1(n3109), .A2(n3108), .ZN(U3210) );
  INV_X1 U3938 ( .A(n3110), .ZN(n3797) );
  AND2_X1 U3939 ( .A1(n3797), .A2(n3802), .ZN(n3881) );
  INV_X1 U3940 ( .A(n3881), .ZN(n3111) );
  XNOR2_X1 U3941 ( .A(n3112), .B(n3111), .ZN(n3113) );
  NAND2_X1 U3942 ( .A1(n3113), .A2(n4281), .ZN(n3116) );
  AOI22_X1 U3943 ( .A1(n3953), .A2(n4275), .B1(n4276), .B2(n3114), .ZN(n3115)
         );
  OAI211_X1 U3944 ( .C1(n4279), .C2(n3119), .A(n3116), .B(n3115), .ZN(n4663)
         );
  INV_X1 U3945 ( .A(n4663), .ZN(n3126) );
  XNOR2_X1 U3946 ( .A(n3117), .B(n3881), .ZN(n4666) );
  OAI21_X1 U3947 ( .B1(n3120), .B2(n3119), .A(n3118), .ZN(n4662) );
  NOR2_X1 U3948 ( .A1(n4662), .A2(n4317), .ZN(n3124) );
  INV_X1 U3949 ( .A(n3121), .ZN(n3122) );
  OAI22_X1 U3950 ( .A1(n4289), .A2(n3578), .B1(n3122), .B2(n4287), .ZN(n3123)
         );
  AOI211_X1 U3951 ( .C1(n4666), .C2(n4030), .A(n3124), .B(n3123), .ZN(n3125)
         );
  OAI21_X1 U3952 ( .B1(n3126), .B2(n4623), .A(n3125), .ZN(U3285) );
  INV_X1 U3953 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3127) );
  NOR2_X1 U3954 ( .A1(n4675), .A2(n3127), .ZN(n3128) );
  AOI21_X1 U3955 ( .B1(n3129), .B2(n4455), .A(n3128), .ZN(n3130) );
  OAI21_X1 U3956 ( .B1(n3131), .B2(n4673), .A(n3130), .ZN(U3479) );
  XOR2_X1 U3957 ( .A(n3132), .B(n3884), .Z(n3136) );
  OAI22_X1 U3958 ( .A1(n3133), .A2(n4296), .B1(n3245), .B2(n4298), .ZN(n3134)
         );
  AOI21_X1 U3959 ( .B1(n3137), .B2(n4306), .A(n3134), .ZN(n3135) );
  OAI21_X1 U3960 ( .B1(n3136), .B2(n4309), .A(n3135), .ZN(n4670) );
  INV_X1 U3961 ( .A(n4670), .ZN(n3150) );
  INV_X1 U3962 ( .A(n4192), .ZN(n3148) );
  NAND2_X1 U3963 ( .A1(n3138), .A2(n3137), .ZN(n3139) );
  NAND2_X1 U3964 ( .A1(n3139), .A2(n4653), .ZN(n3140) );
  NOR2_X1 U3965 ( .A1(n3156), .A2(n3140), .ZN(n4671) );
  OAI22_X1 U3966 ( .A1(n4289), .A2(n3142), .B1(n3141), .B2(n4287), .ZN(n3147)
         );
  INV_X1 U3967 ( .A(n3143), .ZN(n3145) );
  AND2_X1 U3968 ( .A1(n3144), .A2(n3884), .ZN(n4669) );
  NOR3_X1 U3969 ( .A1(n3145), .A2(n4669), .A3(n4242), .ZN(n3146) );
  AOI211_X1 U3970 ( .C1(n3148), .C2(n4671), .A(n3147), .B(n3146), .ZN(n3149)
         );
  OAI21_X1 U3971 ( .B1(n4623), .B2(n3150), .A(n3149), .ZN(U3283) );
  AND2_X1 U3972 ( .A1(n3810), .A2(n3806), .ZN(n3878) );
  XOR2_X1 U3973 ( .A(n3151), .B(n3878), .Z(n3154) );
  AOI22_X1 U3974 ( .A1(n3951), .A2(n4275), .B1(n4276), .B2(n3949), .ZN(n3152)
         );
  OAI21_X1 U3975 ( .B1(n3184), .B2(n4279), .A(n3152), .ZN(n3153) );
  AOI21_X1 U3976 ( .B1(n3154), .B2(n4281), .A(n3153), .ZN(n3191) );
  XOR2_X1 U3977 ( .A(n3155), .B(n3878), .Z(n3192) );
  INV_X1 U3978 ( .A(n3192), .ZN(n3160) );
  NOR2_X1 U3979 ( .A1(n3156), .A2(n3184), .ZN(n3157) );
  OR2_X1 U3980 ( .A1(n3207), .A2(n3157), .ZN(n3197) );
  AOI22_X1 U3981 ( .A1(n4623), .A2(REG2_REG_8__SCAN_IN), .B1(n3188), .B2(n4618), .ZN(n3158) );
  OAI21_X1 U3982 ( .B1(n3197), .B2(n4317), .A(n3158), .ZN(n3159) );
  AOI21_X1 U3983 ( .B1(n3160), .B2(n4030), .A(n3159), .ZN(n3161) );
  OAI21_X1 U3984 ( .B1(n4623), .B2(n3191), .A(n3161), .ZN(U3282) );
  XNOR2_X1 U3985 ( .A(n3279), .B(REG2_REG_10__SCAN_IN), .ZN(n3170) );
  NAND2_X1 U3986 ( .A1(U3149), .A2(REG3_REG_10__SCAN_IN), .ZN(n3629) );
  INV_X1 U3987 ( .A(n3629), .ZN(n3164) );
  INV_X1 U3988 ( .A(n4487), .ZN(n3287) );
  NOR2_X1 U3989 ( .A1(n4604), .A2(n3287), .ZN(n3163) );
  AOI211_X1 U3990 ( .C1(n4595), .C2(ADDR_REG_10__SCAN_IN), .A(n3164), .B(n3163), .ZN(n3169) );
  INV_X1 U3991 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3576) );
  XNOR2_X2 U3992 ( .A(n3286), .B(n3287), .ZN(n3167) );
  OAI211_X1 U3993 ( .C1(n3167), .C2(REG1_REG_10__SCAN_IN), .A(n3289), .B(n4584), .ZN(n3168) );
  OAI211_X1 U3994 ( .C1(n3170), .C2(n4596), .A(n3169), .B(n3168), .ZN(U3250)
         );
  INV_X1 U3995 ( .A(n3171), .ZN(n3172) );
  OR2_X1 U3996 ( .A1(n3184), .A2(n3431), .ZN(n3174) );
  OAI21_X1 U3997 ( .B1(n3245), .B2(n3337), .A(n3174), .ZN(n3175) );
  XNOR2_X1 U3998 ( .A(n3175), .B(n3433), .ZN(n3177) );
  OR2_X1 U3999 ( .A1(n3184), .A2(n3432), .ZN(n3176) );
  OAI21_X1 U4000 ( .B1(n3245), .B2(n3436), .A(n3176), .ZN(n3178) );
  NAND2_X1 U4001 ( .A1(n3177), .A2(n3178), .ZN(n3238) );
  NAND2_X1 U4002 ( .A1(n3242), .A2(n3238), .ZN(n3237) );
  INV_X1 U4003 ( .A(n3237), .ZN(n3182) );
  INV_X1 U4004 ( .A(n3177), .ZN(n3180) );
  INV_X1 U4005 ( .A(n3178), .ZN(n3179) );
  NAND2_X1 U4006 ( .A1(n3180), .A2(n3179), .ZN(n3239) );
  AOI21_X1 U4007 ( .B1(n3239), .B2(n3238), .A(n3242), .ZN(n3181) );
  AOI21_X1 U4008 ( .B1(n3182), .B2(n3239), .A(n3181), .ZN(n3190) );
  OAI22_X1 U4009 ( .A1(n3775), .A2(n3184), .B1(STATE_REG_SCAN_IN), .B2(n3183), 
        .ZN(n3187) );
  OAI22_X1 U4010 ( .A1(n3185), .A2(n3777), .B1(n3776), .B2(n3627), .ZN(n3186)
         );
  AOI211_X1 U4011 ( .C1(n3188), .C2(n3780), .A(n3187), .B(n3186), .ZN(n3189)
         );
  OAI21_X1 U4012 ( .B1(n3190), .B2(n3782), .A(n3189), .ZN(U3218) );
  OAI21_X1 U4013 ( .B1(n3192), .B2(n4668), .A(n3191), .ZN(n3199) );
  INV_X1 U4014 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3193) );
  OAI22_X1 U4015 ( .A1(n3197), .A2(n4395), .B1(n4684), .B2(n3193), .ZN(n3194)
         );
  AOI21_X1 U4016 ( .B1(n3199), .B2(n4684), .A(n3194), .ZN(n3195) );
  INV_X1 U4017 ( .A(n3195), .ZN(U3526) );
  INV_X1 U4018 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3196) );
  OAI22_X1 U4019 ( .A1(n3197), .A2(n4476), .B1(n4675), .B2(n3196), .ZN(n3198)
         );
  AOI21_X1 U4020 ( .B1(n3199), .B2(n4675), .A(n3198), .ZN(n3200) );
  INV_X1 U4021 ( .A(n3200), .ZN(U3483) );
  INV_X1 U4022 ( .A(n3814), .ZN(n3202) );
  NAND2_X1 U4023 ( .A1(n3202), .A2(n3811), .ZN(n3874) );
  XNOR2_X1 U4024 ( .A(n3201), .B(n3874), .ZN(n3232) );
  XNOR2_X1 U4025 ( .A(n3203), .B(n3874), .ZN(n3204) );
  NAND2_X1 U4026 ( .A1(n3204), .A2(n4281), .ZN(n3206) );
  AOI22_X1 U4027 ( .A1(n3950), .A2(n4275), .B1(n4276), .B2(n3948), .ZN(n3205)
         );
  OAI211_X1 U4028 ( .C1(n4279), .C2(n3249), .A(n3206), .B(n3205), .ZN(n3228)
         );
  INV_X1 U4029 ( .A(n3207), .ZN(n3209) );
  INV_X1 U4030 ( .A(n3222), .ZN(n3208) );
  AOI21_X1 U4031 ( .B1(n3233), .B2(n3209), .A(n3208), .ZN(n3229) );
  INV_X1 U4032 ( .A(n3229), .ZN(n3211) );
  AOI22_X1 U4033 ( .A1(n4623), .A2(REG2_REG_9__SCAN_IN), .B1(n3246), .B2(n4618), .ZN(n3210) );
  OAI21_X1 U4034 ( .B1(n3211), .B2(n4317), .A(n3210), .ZN(n3212) );
  AOI21_X1 U4035 ( .B1(n3228), .B2(n4289), .A(n3212), .ZN(n3213) );
  OAI21_X1 U4036 ( .B1(n4242), .B2(n3232), .A(n3213), .ZN(U3281) );
  NAND2_X1 U4037 ( .A1(n3228), .A2(n4684), .ZN(n3215) );
  AOI22_X1 U4038 ( .A1(n3229), .A2(n4372), .B1(REG1_REG_9__SCAN_IN), .B2(n4681), .ZN(n3214) );
  OAI211_X1 U4039 ( .C1(n3232), .C2(n4390), .A(n3215), .B(n3214), .ZN(U3527)
         );
  NAND2_X1 U4040 ( .A1(n3813), .A2(n3816), .ZN(n3875) );
  XNOR2_X1 U4041 ( .A(n3216), .B(n3875), .ZN(n3219) );
  OAI22_X1 U4042 ( .A1(n3627), .A2(n4296), .B1(n3626), .B2(n4298), .ZN(n3217)
         );
  AOI21_X1 U40430 ( .B1(n3264), .B2(n4306), .A(n3217), .ZN(n3218) );
  OAI21_X1 U4044 ( .B1(n3219), .B2(n4309), .A(n3218), .ZN(n3254) );
  INV_X1 U4045 ( .A(n3254), .ZN(n3227) );
  XNOR2_X1 U4046 ( .A(n3220), .B(n3875), .ZN(n3255) );
  INV_X1 U4047 ( .A(n4312), .ZN(n3221) );
  AOI21_X1 U4048 ( .B1(n3264), .B2(n3222), .A(n3221), .ZN(n3257) );
  INV_X1 U4049 ( .A(n3257), .ZN(n3224) );
  AOI22_X1 U4050 ( .A1(n4623), .A2(REG2_REG_10__SCAN_IN), .B1(n3628), .B2(
        n4618), .ZN(n3223) );
  OAI21_X1 U4051 ( .B1(n3224), .B2(n4317), .A(n3223), .ZN(n3225) );
  AOI21_X1 U4052 ( .B1(n3255), .B2(n4030), .A(n3225), .ZN(n3226) );
  OAI21_X1 U4053 ( .B1(n3227), .B2(n4623), .A(n3226), .ZN(U3280) );
  NAND2_X1 U4054 ( .A1(n3228), .A2(n4675), .ZN(n3231) );
  AOI22_X1 U4055 ( .A1(n3229), .A2(n4455), .B1(REG0_REG_9__SCAN_IN), .B2(n4673), .ZN(n3230) );
  OAI211_X1 U4056 ( .C1(n3232), .C2(n4471), .A(n3231), .B(n3230), .ZN(U3485)
         );
  OAI22_X1 U4057 ( .A1(n3249), .A2(n3432), .B1(n3627), .B2(n3436), .ZN(n3261)
         );
  NAND2_X1 U4058 ( .A1(n3233), .A2(n3393), .ZN(n3235) );
  NAND2_X1 U4059 ( .A1(n3949), .A2(n3263), .ZN(n3234) );
  NAND2_X1 U4060 ( .A1(n3235), .A2(n3234), .ZN(n3236) );
  XNOR2_X1 U4061 ( .A(n3236), .B(n3433), .ZN(n3260) );
  XOR2_X1 U4062 ( .A(n3261), .B(n3260), .Z(n3244) );
  NAND2_X1 U4063 ( .A1(n3237), .A2(n3239), .ZN(n3243) );
  AND2_X1 U4064 ( .A1(n3238), .A2(n3244), .ZN(n3241) );
  INV_X1 U4065 ( .A(n3244), .ZN(n3240) );
  OAI21_X1 U4066 ( .B1(n3244), .B2(n3243), .A(n3262), .ZN(n3252) );
  OAI22_X1 U4067 ( .A1(n3245), .A2(n3777), .B1(n3776), .B2(n4297), .ZN(n3251)
         );
  NAND2_X1 U4068 ( .A1(n3780), .A2(n3246), .ZN(n3248) );
  OAI211_X1 U4069 ( .C1(n3775), .C2(n3249), .A(n3248), .B(n3247), .ZN(n3250)
         );
  AOI211_X1 U4070 ( .C1(n3252), .C2(n3733), .A(n3251), .B(n3250), .ZN(n3253)
         );
  INV_X1 U4071 ( .A(n3253), .ZN(U3228) );
  AOI21_X1 U4072 ( .B1(n4665), .B2(n3255), .A(n3254), .ZN(n3259) );
  AOI22_X1 U4073 ( .A1(n3257), .A2(n4372), .B1(REG1_REG_10__SCAN_IN), .B2(
        n4681), .ZN(n3256) );
  OAI21_X1 U4074 ( .B1(n3259), .B2(n4681), .A(n3256), .ZN(U3528) );
  AOI22_X1 U4075 ( .A1(n3257), .A2(n4455), .B1(REG0_REG_10__SCAN_IN), .B2(
        n4673), .ZN(n3258) );
  OAI21_X1 U4076 ( .B1(n3259), .B2(n4673), .A(n3258), .ZN(U3487) );
  AOI22_X1 U4077 ( .A1(n3399), .A2(n3948), .B1(n3264), .B2(n3263), .ZN(n3267)
         );
  OAI22_X1 U4078 ( .A1(n3631), .A2(n3431), .B1(n4297), .B2(n3432), .ZN(n3265)
         );
  XNOR2_X1 U4079 ( .A(n3265), .B(n3433), .ZN(n3266) );
  XOR2_X1 U4080 ( .A(n3267), .B(n3266), .Z(n3625) );
  INV_X1 U4081 ( .A(n3266), .ZN(n3268) );
  OAI22_X1 U4082 ( .A1(n3272), .A2(n3431), .B1(n3626), .B2(n3432), .ZN(n3269)
         );
  XNOR2_X1 U4083 ( .A(n3269), .B(n3433), .ZN(n3311) );
  INV_X1 U4084 ( .A(n3307), .ZN(n3309) );
  XNOR2_X1 U4085 ( .A(n3311), .B(n3309), .ZN(n3270) );
  XNOR2_X1 U4086 ( .A(n3271), .B(n3270), .ZN(n3276) );
  NAND2_X1 U4087 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n3277) );
  OAI21_X1 U4088 ( .B1(n3775), .B2(n3272), .A(n3277), .ZN(n3274) );
  OAI22_X1 U4089 ( .A1(n4299), .A2(n3776), .B1(n3777), .B2(n4297), .ZN(n3273)
         );
  AOI211_X1 U4090 ( .C1(n4315), .C2(n3780), .A(n3274), .B(n3273), .ZN(n3275)
         );
  OAI21_X1 U4091 ( .B1(n3276), .B2(n3782), .A(n3275), .ZN(U3233) );
  INV_X1 U4092 ( .A(ADDR_REG_11__SCAN_IN), .ZN(n3278) );
  OAI21_X1 U4093 ( .B1(n4563), .B2(n3278), .A(n3277), .ZN(n3285) );
  AOI22_X1 U4094 ( .A1(n3279), .A2(REG2_REG_10__SCAN_IN), .B1(n4487), .B2(
        n2152), .ZN(n3283) );
  INV_X1 U4095 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3280) );
  MUX2_X1 U4096 ( .A(n3280), .B(REG2_REG_11__SCAN_IN), .S(n4486), .Z(n3282) );
  INV_X1 U4097 ( .A(n3974), .ZN(n3281) );
  AOI211_X1 U4098 ( .C1(n3283), .C2(n3282), .A(n4596), .B(n3281), .ZN(n3284)
         );
  AOI211_X1 U4099 ( .C1(n4559), .C2(n4486), .A(n3285), .B(n3284), .ZN(n3293)
         );
  INV_X1 U4100 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4393) );
  XNOR2_X1 U4101 ( .A(n4486), .B(n4393), .ZN(n3290) );
  OAI211_X1 U4102 ( .C1(n3291), .C2(n3290), .A(n3979), .B(n4584), .ZN(n3292)
         );
  NAND2_X1 U4103 ( .A1(n3293), .A2(n3292), .ZN(U3251) );
  OR2_X1 U4104 ( .A1(n3294), .A2(n4302), .ZN(n4300) );
  NAND2_X1 U4105 ( .A1(n4300), .A2(n3295), .ZN(n3296) );
  AND2_X1 U4106 ( .A1(n4268), .A2(n4269), .ZN(n3893) );
  XNOR2_X1 U4107 ( .A(n3296), .B(n3893), .ZN(n4472) );
  NAND2_X1 U4108 ( .A1(n3298), .A2(n3297), .ZN(n4271) );
  XOR2_X1 U4109 ( .A(n4271), .B(n3893), .Z(n3301) );
  OAI22_X1 U4110 ( .A1(n3422), .A2(n4298), .B1(n3626), .B2(n4296), .ZN(n3299)
         );
  AOI21_X1 U4111 ( .B1(n3316), .B2(n4306), .A(n3299), .ZN(n3300) );
  OAI21_X1 U4112 ( .B1(n3301), .B2(n4309), .A(n3300), .ZN(n4387) );
  NOR2_X1 U4113 ( .A1(n4314), .A2(n3421), .ZN(n4385) );
  INV_X1 U4114 ( .A(n3302), .ZN(n4384) );
  NOR3_X1 U4115 ( .A1(n4385), .A2(n4384), .A3(n4317), .ZN(n3305) );
  INV_X1 U4116 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3985) );
  INV_X1 U4117 ( .A(n3425), .ZN(n3303) );
  OAI22_X1 U4118 ( .A1(n4289), .A2(n3985), .B1(n3303), .B2(n4287), .ZN(n3304)
         );
  AOI211_X1 U4119 ( .C1(n4387), .C2(n4289), .A(n3305), .B(n3304), .ZN(n3306)
         );
  OAI21_X1 U4120 ( .B1(n4472), .B2(n4242), .A(n3306), .ZN(U3278) );
  NAND2_X1 U4121 ( .A1(n3308), .A2(n3307), .ZN(n3312) );
  INV_X1 U4122 ( .A(n3308), .ZN(n3310) );
  NAND2_X1 U4123 ( .A1(n3316), .A2(n3393), .ZN(n3314) );
  NAND2_X1 U4124 ( .A1(n4274), .A2(n3263), .ZN(n3313) );
  NAND2_X1 U4125 ( .A1(n3314), .A2(n3313), .ZN(n3315) );
  XNOR2_X1 U4126 ( .A(n3315), .B(n3396), .ZN(n3320) );
  INV_X1 U4127 ( .A(n3320), .ZN(n3318) );
  AOI22_X1 U4128 ( .A1(n3399), .A2(n4274), .B1(n3316), .B2(n3392), .ZN(n3319)
         );
  INV_X1 U4129 ( .A(n3319), .ZN(n3317) );
  NAND2_X1 U4130 ( .A1(n3318), .A2(n3317), .ZN(n3419) );
  OAI22_X1 U4131 ( .A1(n4285), .A2(n3431), .B1(n3422), .B2(n3432), .ZN(n3321)
         );
  XOR2_X1 U4132 ( .A(n3433), .B(n3321), .Z(n3713) );
  INV_X1 U4133 ( .A(n3713), .ZN(n3322) );
  OAI22_X1 U4134 ( .A1(n4285), .A2(n3337), .B1(n3422), .B2(n3436), .ZN(n3712)
         );
  NAND2_X1 U4135 ( .A1(n4256), .A2(n3393), .ZN(n3323) );
  OAI21_X1 U4136 ( .B1(n4228), .B2(n3337), .A(n3323), .ZN(n3324) );
  XNOR2_X1 U4137 ( .A(n3324), .B(n3433), .ZN(n3326) );
  NAND2_X1 U4138 ( .A1(n4256), .A2(n3392), .ZN(n3325) );
  OAI21_X1 U4139 ( .B1(n4228), .B2(n3436), .A(n3325), .ZN(n3327) );
  NAND2_X1 U4140 ( .A1(n3326), .A2(n3327), .ZN(n3470) );
  INV_X1 U4141 ( .A(n3326), .ZN(n3329) );
  INV_X1 U4142 ( .A(n3327), .ZN(n3328) );
  NAND2_X1 U4143 ( .A1(n3329), .A2(n3328), .ZN(n3469) );
  NAND2_X1 U4144 ( .A1(n4238), .A2(n3393), .ZN(n3332) );
  NAND2_X1 U4145 ( .A1(n4250), .A2(n3392), .ZN(n3331) );
  NAND2_X1 U4146 ( .A1(n3332), .A2(n3331), .ZN(n3333) );
  XNOR2_X1 U4147 ( .A(n3333), .B(n3433), .ZN(n3667) );
  NAND2_X1 U4148 ( .A1(n4221), .A2(n3392), .ZN(n3334) );
  OAI21_X1 U4149 ( .B1(n4229), .B2(n3436), .A(n3334), .ZN(n3681) );
  NAND2_X1 U4150 ( .A1(n4238), .A2(n3263), .ZN(n3336) );
  NAND2_X1 U4151 ( .A1(n3399), .A2(n4250), .ZN(n3335) );
  NAND2_X1 U4152 ( .A1(n3336), .A2(n3335), .ZN(n3771) );
  OR2_X1 U4153 ( .A1(n3681), .A2(n3771), .ZN(n3345) );
  OAI22_X1 U4154 ( .A1(n4217), .A2(n3337), .B1(n3431), .B2(n3339), .ZN(n3338)
         );
  XNOR2_X1 U4155 ( .A(n3338), .B(n3396), .ZN(n3683) );
  NOR2_X1 U4156 ( .A1(n3339), .A2(n3432), .ZN(n3340) );
  AOI21_X1 U4157 ( .B1(n4185), .B2(n3399), .A(n3340), .ZN(n3682) );
  NAND2_X1 U4158 ( .A1(n3683), .A2(n3682), .ZN(n3344) );
  OAI22_X1 U4159 ( .A1(n4229), .A2(n3432), .B1(n3671), .B2(n3431), .ZN(n3341)
         );
  XNOR2_X1 U4160 ( .A(n3341), .B(n3396), .ZN(n3669) );
  OAI21_X1 U4161 ( .B1(n3667), .B2(n3771), .A(n3681), .ZN(n3342) );
  NAND2_X1 U4162 ( .A1(n3669), .A2(n3342), .ZN(n3343) );
  OAI211_X1 U4163 ( .C1(n3667), .C2(n3345), .A(n3344), .B(n3343), .ZN(n3745)
         );
  INV_X1 U4164 ( .A(n3669), .ZN(n3680) );
  AND2_X1 U4165 ( .A1(n3667), .A2(n3771), .ZN(n3346) );
  AOI21_X1 U4166 ( .B1(n3680), .B2(n3681), .A(n3346), .ZN(n3743) );
  OAI22_X1 U4167 ( .A1(n4205), .A2(n3432), .B1(n3431), .B2(n4191), .ZN(n3347)
         );
  XNOR2_X1 U4168 ( .A(n3347), .B(n3433), .ZN(n3353) );
  OAI22_X1 U4169 ( .A1(n4205), .A2(n3436), .B1(n3432), .B2(n4191), .ZN(n3352)
         );
  NAND2_X1 U4170 ( .A1(n3353), .A2(n3352), .ZN(n3741) );
  INV_X1 U4171 ( .A(n3683), .ZN(n3349) );
  INV_X1 U4172 ( .A(n3682), .ZN(n3348) );
  NAND2_X1 U4173 ( .A1(n3349), .A2(n3348), .ZN(n3744) );
  OAI211_X1 U4174 ( .C1(n3745), .C2(n3743), .A(n3741), .B(n3744), .ZN(n3350)
         );
  INV_X1 U4175 ( .A(n3350), .ZN(n3351) );
  OR2_X1 U4176 ( .A1(n3353), .A2(n3352), .ZN(n3742) );
  OAI22_X1 U4177 ( .A1(n4187), .A2(n3436), .B1(n3432), .B2(n3640), .ZN(n3356)
         );
  OAI22_X1 U4178 ( .A1(n4187), .A2(n3432), .B1(n3431), .B2(n3640), .ZN(n3354)
         );
  XNOR2_X1 U4179 ( .A(n3354), .B(n3433), .ZN(n3355) );
  XOR2_X1 U4180 ( .A(n3356), .B(n3355), .Z(n3638) );
  NAND2_X1 U4181 ( .A1(n3360), .A2(n3359), .ZN(n3702) );
  NAND2_X1 U4182 ( .A1(n4129), .A2(n3392), .ZN(n3362) );
  NAND2_X1 U4183 ( .A1(n3393), .A2(n4154), .ZN(n3361) );
  NAND2_X1 U4184 ( .A1(n3362), .A2(n3361), .ZN(n3363) );
  XNOR2_X1 U4185 ( .A(n3363), .B(n3433), .ZN(n3366) );
  NAND2_X1 U4186 ( .A1(n4129), .A2(n3399), .ZN(n3365) );
  NAND2_X1 U4187 ( .A1(n3392), .A2(n4154), .ZN(n3364) );
  NAND2_X1 U4188 ( .A1(n3365), .A2(n3364), .ZN(n3367) );
  NAND2_X1 U4189 ( .A1(n3366), .A2(n3367), .ZN(n3703) );
  INV_X1 U4190 ( .A(n3366), .ZN(n3369) );
  INV_X1 U4191 ( .A(n3367), .ZN(n3368) );
  NAND2_X1 U4192 ( .A1(n3369), .A2(n3368), .ZN(n3705) );
  NAND2_X1 U4193 ( .A1(n4149), .A2(n3392), .ZN(n3371) );
  NAND2_X1 U4194 ( .A1(n3393), .A2(n4128), .ZN(n3370) );
  NAND2_X1 U4195 ( .A1(n3371), .A2(n3370), .ZN(n3372) );
  XNOR2_X1 U4196 ( .A(n3372), .B(n3433), .ZN(n3646) );
  NAND2_X1 U4197 ( .A1(n4149), .A2(n3399), .ZN(n3374) );
  NAND2_X1 U4198 ( .A1(n3392), .A2(n4128), .ZN(n3373) );
  NAND2_X1 U4199 ( .A1(n3374), .A2(n3373), .ZN(n3645) );
  NOR2_X1 U4200 ( .A1(n3646), .A2(n3645), .ZN(n3376) );
  NAND2_X1 U4201 ( .A1(n3646), .A2(n3645), .ZN(n3375) );
  OAI22_X1 U4202 ( .A1(n4131), .A2(n3432), .B1(n3431), .B2(n4112), .ZN(n3377)
         );
  XNOR2_X1 U4203 ( .A(n3377), .B(n3433), .ZN(n3380) );
  OAI22_X1 U4204 ( .A1(n4131), .A2(n3436), .B1(n3432), .B2(n4112), .ZN(n3379)
         );
  XNOR2_X1 U4205 ( .A(n3380), .B(n3379), .ZN(n3722) );
  OAI22_X1 U4206 ( .A1(n4115), .A2(n3432), .B1(n3483), .B2(n3431), .ZN(n3378)
         );
  XNOR2_X1 U4207 ( .A(n3378), .B(n3433), .ZN(n3384) );
  OAI22_X1 U4208 ( .A1(n4115), .A2(n3436), .B1(n3483), .B2(n3432), .ZN(n3383)
         );
  XNOR2_X1 U4209 ( .A(n3384), .B(n3383), .ZN(n3478) );
  NOR2_X1 U4210 ( .A1(n3380), .A2(n3379), .ZN(n3479) );
  NOR2_X1 U4211 ( .A1(n3478), .A2(n3479), .ZN(n3381) );
  NOR2_X1 U4212 ( .A1(n3432), .A2(n4080), .ZN(n3382) );
  AOI21_X1 U4213 ( .B1(n4065), .B2(n3399), .A(n3382), .ZN(n3388) );
  NAND2_X1 U4214 ( .A1(n3384), .A2(n3383), .ZN(n3387) );
  OAI22_X1 U4215 ( .A1(n4102), .A2(n3432), .B1(n4080), .B2(n3431), .ZN(n3386)
         );
  XNOR2_X1 U4216 ( .A(n3386), .B(n3433), .ZN(n3694) );
  NAND2_X1 U4217 ( .A1(n3692), .A2(n3694), .ZN(n3391) );
  NAND2_X1 U4218 ( .A1(n3480), .A2(n3387), .ZN(n3390) );
  INV_X1 U4219 ( .A(n3388), .ZN(n3389) );
  NAND2_X1 U4220 ( .A1(n3390), .A2(n3389), .ZN(n3690) );
  NAND2_X1 U4221 ( .A1(n3391), .A2(n3690), .ZN(n3658) );
  NAND2_X1 U4222 ( .A1(n4077), .A2(n3392), .ZN(n3395) );
  NAND2_X1 U4223 ( .A1(n3393), .A2(n4064), .ZN(n3394) );
  NAND2_X1 U4224 ( .A1(n3395), .A2(n3394), .ZN(n3397) );
  XNOR2_X1 U4225 ( .A(n3397), .B(n3396), .ZN(n3401) );
  AND2_X1 U4226 ( .A1(n3392), .A2(n4064), .ZN(n3398) );
  AOI21_X1 U4227 ( .B1(n4077), .B2(n3399), .A(n3398), .ZN(n3400) );
  NAND2_X1 U4228 ( .A1(n3401), .A2(n3400), .ZN(n3655) );
  NOR2_X1 U4229 ( .A1(n3401), .A2(n3400), .ZN(n3656) );
  OAI22_X1 U4230 ( .A1(n4067), .A2(n3432), .B1(n4051), .B2(n3431), .ZN(n3402)
         );
  XNOR2_X1 U4231 ( .A(n3402), .B(n3433), .ZN(n3403) );
  OAI22_X1 U4232 ( .A1(n4067), .A2(n3436), .B1(n4051), .B2(n3432), .ZN(n3404)
         );
  NAND2_X1 U4233 ( .A1(n3403), .A2(n3404), .ZN(n3759) );
  INV_X1 U4234 ( .A(n3403), .ZN(n3406) );
  INV_X1 U4235 ( .A(n3404), .ZN(n3405) );
  NAND2_X1 U4236 ( .A1(n3406), .A2(n3405), .ZN(n3760) );
  OAI22_X1 U4237 ( .A1(n3763), .A2(n3432), .B1(n3431), .B2(n4022), .ZN(n3407)
         );
  XNOR2_X1 U4238 ( .A(n3407), .B(n3433), .ZN(n3440) );
  OAI22_X1 U4239 ( .A1(n3763), .A2(n3436), .B1(n3432), .B2(n4022), .ZN(n3439)
         );
  XNOR2_X1 U4240 ( .A(n3440), .B(n3439), .ZN(n3430) );
  OAI22_X1 U4241 ( .A1(n4067), .A2(n3777), .B1(n3752), .B2(n4036), .ZN(n3408)
         );
  INV_X1 U4242 ( .A(n3408), .ZN(n3410) );
  AOI22_X1 U4243 ( .A1(n3754), .A2(n4032), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3409) );
  OAI211_X1 U4244 ( .C1(n4025), .C2(n3776), .A(n3410), .B(n3409), .ZN(n3411)
         );
  INV_X1 U4245 ( .A(n3411), .ZN(n3412) );
  OAI21_X1 U4246 ( .B1(n3413), .B2(n3782), .A(n3412), .ZN(U3211) );
  INV_X1 U4247 ( .A(DATAI_24_), .ZN(n3608) );
  NAND2_X1 U4248 ( .A1(n2688), .A2(STATE_REG_SCAN_IN), .ZN(n3414) );
  OAI21_X1 U4249 ( .B1(STATE_REG_SCAN_IN), .B2(n3608), .A(n3414), .ZN(U3328)
         );
  NOR3_X1 U4250 ( .A1(n2688), .A2(n4631), .A3(n3415), .ZN(n3416) );
  AOI21_X1 U4251 ( .B1(n4628), .B2(n3417), .A(n3416), .ZN(U3458) );
  NAND2_X1 U4252 ( .A1(n2050), .A2(n3419), .ZN(n3420) );
  XNOR2_X1 U4253 ( .A(n3418), .B(n3420), .ZN(n3427) );
  NAND2_X1 U4254 ( .A1(U3149), .A2(REG3_REG_12__SCAN_IN), .ZN(n3975) );
  OAI21_X1 U4255 ( .B1(n3775), .B2(n3421), .A(n3975), .ZN(n3424) );
  OAI22_X1 U4256 ( .A1(n3626), .A2(n3777), .B1(n3776), .B2(n3422), .ZN(n3423)
         );
  AOI211_X1 U4257 ( .C1(n3425), .C2(n3780), .A(n3424), .B(n3423), .ZN(n3426)
         );
  OAI21_X1 U4258 ( .B1(n3427), .B2(n3782), .A(n3426), .ZN(U3221) );
  INV_X1 U4259 ( .A(DATAI_30_), .ZN(n3541) );
  NAND2_X1 U4260 ( .A1(n3428), .A2(STATE_REG_SCAN_IN), .ZN(n3429) );
  OAI21_X1 U4261 ( .B1(STATE_REG_SCAN_IN), .B2(n3541), .A(n3429), .ZN(U3322)
         );
  OAI22_X1 U4262 ( .A1(n4025), .A2(n3432), .B1(n3431), .B2(n3435), .ZN(n3434)
         );
  XNOR2_X1 U4263 ( .A(n3434), .B(n3433), .ZN(n3438) );
  OAI22_X1 U4264 ( .A1(n4025), .A2(n3436), .B1(n3432), .B2(n3435), .ZN(n3437)
         );
  XNOR2_X1 U4265 ( .A(n3438), .B(n3437), .ZN(n3442) );
  NAND2_X1 U4266 ( .A1(n3442), .A2(n3733), .ZN(n3453) );
  AND2_X1 U4267 ( .A1(n3440), .A2(n3439), .ZN(n3443) );
  NOR3_X1 U4268 ( .A1(n3442), .A2(n3443), .A3(n3782), .ZN(n3441) );
  INV_X1 U4269 ( .A(n3442), .ZN(n3445) );
  INV_X1 U4270 ( .A(n3443), .ZN(n3444) );
  NOR3_X1 U4271 ( .A1(n3445), .A2(n3782), .A3(n3444), .ZN(n3450) );
  AOI22_X1 U4272 ( .A1(n3750), .A2(n3943), .B1(n4047), .B2(n3749), .ZN(n3448)
         );
  AOI22_X1 U4273 ( .A1(n3754), .A2(n3446), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3447) );
  OAI211_X1 U4274 ( .C1(n3752), .C2(n3456), .A(n3448), .B(n3447), .ZN(n3449)
         );
  NOR2_X1 U4275 ( .A1(n3450), .A2(n3449), .ZN(n3451) );
  OAI211_X1 U4276 ( .C1(n2309), .C2(n3453), .A(n3452), .B(n3451), .ZN(U3217)
         );
  INV_X1 U4277 ( .A(n3454), .ZN(n3460) );
  INV_X1 U4278 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3455) );
  OAI22_X1 U4279 ( .A1(n3456), .A2(n4287), .B1(n3455), .B2(n4289), .ZN(n3459)
         );
  NOR2_X1 U4280 ( .A1(n3457), .A2(n4623), .ZN(n3458) );
  XNOR2_X1 U4281 ( .A(n3463), .B(n3462), .ZN(n3957) );
  NAND2_X1 U4282 ( .A1(n3735), .A2(REG3_REG_0__SCAN_IN), .ZN(n3464) );
  OAI21_X1 U4283 ( .B1(n3782), .B2(n3957), .A(n3464), .ZN(n3465) );
  AOI21_X1 U4284 ( .B1(n3466), .B2(n3754), .A(n3465), .ZN(n3467) );
  OAI21_X1 U4285 ( .B1(n3468), .B2(n3776), .A(n3467), .ZN(U3229) );
  NAND2_X1 U4286 ( .A1(n3470), .A2(n3469), .ZN(n3471) );
  XNOR2_X1 U4287 ( .A(n3472), .B(n3471), .ZN(n3476) );
  AOI22_X1 U4288 ( .A1(n3750), .A2(n4250), .B1(n3749), .B2(n4249), .ZN(n3475)
         );
  NOR2_X1 U4289 ( .A1(n3544), .A2(STATE_REG_SCAN_IN), .ZN(n3988) );
  NOR2_X1 U4290 ( .A1(n3752), .A2(n4258), .ZN(n3473) );
  AOI211_X1 U4291 ( .C1(n4256), .C2(n3754), .A(n3988), .B(n3473), .ZN(n3474)
         );
  OAI211_X1 U4292 ( .C1(n3476), .C2(n3782), .A(n3475), .B(n3474), .ZN(U3212)
         );
  INV_X1 U4293 ( .A(n3477), .ZN(n3720) );
  OAI21_X1 U4294 ( .B1(n3720), .B2(n3479), .A(n3478), .ZN(n3481) );
  NAND3_X1 U4295 ( .A1(n3481), .A2(n3733), .A3(n3480), .ZN(n3487) );
  INV_X1 U4296 ( .A(n3482), .ZN(n4090) );
  OAI22_X1 U4297 ( .A1(n3775), .A2(n3483), .B1(STATE_REG_SCAN_IN), .B2(n2084), 
        .ZN(n3485) );
  OAI22_X1 U4298 ( .A1(n4102), .A2(n3776), .B1(n4131), .B2(n3777), .ZN(n3484)
         );
  AOI211_X1 U4299 ( .C1(n4090), .C2(n3780), .A(n3485), .B(n3484), .ZN(n3486)
         );
  NAND2_X1 U4300 ( .A1(n3487), .A2(n3486), .ZN(U3213) );
  AOI22_X1 U4301 ( .A1(n3489), .A2(keyinput45), .B1(n3608), .B2(keyinput46), 
        .ZN(n3488) );
  OAI221_X1 U4302 ( .B1(n3489), .B2(keyinput45), .C1(n3608), .C2(keyinput46), 
        .A(n3488), .ZN(n3497) );
  AOI22_X1 U4303 ( .A1(n4627), .A2(keyinput23), .B1(n4626), .B2(keyinput52), 
        .ZN(n3490) );
  OAI221_X1 U4304 ( .B1(n4627), .B2(keyinput23), .C1(n4626), .C2(keyinput52), 
        .A(n3490), .ZN(n3496) );
  INV_X1 U4305 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4495) );
  INV_X1 U4306 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3492) );
  AOI22_X1 U4307 ( .A1(n4495), .A2(keyinput28), .B1(keyinput56), .B2(n3492), 
        .ZN(n3491) );
  OAI221_X1 U4308 ( .B1(n4495), .B2(keyinput28), .C1(n3492), .C2(keyinput56), 
        .A(n3491), .ZN(n3495) );
  AOI22_X1 U4309 ( .A1(n4629), .A2(keyinput36), .B1(n4624), .B2(keyinput9), 
        .ZN(n3493) );
  OAI221_X1 U4310 ( .B1(n4629), .B2(keyinput36), .C1(n4624), .C2(keyinput9), 
        .A(n3493), .ZN(n3494) );
  NOR4_X1 U4311 ( .A1(n3497), .A2(n3496), .A3(n3495), .A4(n3494), .ZN(n3539)
         );
  INV_X1 U4312 ( .A(DATAI_11_), .ZN(n3609) );
  OAI22_X1 U4313 ( .A1(n3609), .A2(keyinput7), .B1(n3499), .B2(keyinput55), 
        .ZN(n3498) );
  AOI221_X1 U4314 ( .B1(n3609), .B2(keyinput7), .C1(keyinput55), .C2(n3499), 
        .A(n3498), .ZN(n3538) );
  XNOR2_X1 U4315 ( .A(n3500), .B(keyinput60), .ZN(n3511) );
  XNOR2_X1 U4316 ( .A(IR_REG_8__SCAN_IN), .B(keyinput53), .ZN(n3504) );
  XNOR2_X1 U4317 ( .A(IR_REG_7__SCAN_IN), .B(keyinput49), .ZN(n3503) );
  XNOR2_X1 U4318 ( .A(REG0_REG_10__SCAN_IN), .B(keyinput20), .ZN(n3502) );
  XNOR2_X1 U4319 ( .A(IR_REG_21__SCAN_IN), .B(keyinput48), .ZN(n3501) );
  NAND4_X1 U4320 ( .A1(n3504), .A2(n3503), .A3(n3502), .A4(n3501), .ZN(n3510)
         );
  INV_X1 U4321 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4208) );
  XNOR2_X1 U4322 ( .A(DATAI_7_), .B(keyinput22), .ZN(n3506) );
  NAND2_X1 U4323 ( .A1(n4208), .A2(keyinput0), .ZN(n3505) );
  OAI211_X1 U4324 ( .C1(n4208), .C2(keyinput0), .A(n3506), .B(n3505), .ZN(
        n3509) );
  XNOR2_X1 U4325 ( .A(n3507), .B(keyinput37), .ZN(n3508) );
  OR4_X1 U4326 ( .A1(n3511), .A2(n3510), .A3(n3509), .A4(n3508), .ZN(n3523) );
  INV_X1 U4327 ( .A(D_REG_23__SCAN_IN), .ZN(n4625) );
  XNOR2_X1 U4328 ( .A(n4625), .B(keyinput25), .ZN(n3522) );
  XNOR2_X1 U4329 ( .A(IR_REG_4__SCAN_IN), .B(keyinput15), .ZN(n3515) );
  XNOR2_X1 U4330 ( .A(REG3_REG_6__SCAN_IN), .B(keyinput63), .ZN(n3514) );
  XNOR2_X1 U4331 ( .A(DATAI_1_), .B(keyinput13), .ZN(n3513) );
  XNOR2_X1 U4332 ( .A(IR_REG_14__SCAN_IN), .B(keyinput32), .ZN(n3512) );
  NAND4_X1 U4333 ( .A1(n3515), .A2(n3514), .A3(n3513), .A4(n3512), .ZN(n3521)
         );
  XNOR2_X1 U4334 ( .A(IR_REG_9__SCAN_IN), .B(keyinput4), .ZN(n3519) );
  XNOR2_X1 U4335 ( .A(IR_REG_22__SCAN_IN), .B(keyinput16), .ZN(n3518) );
  XNOR2_X1 U4336 ( .A(IR_REG_20__SCAN_IN), .B(keyinput14), .ZN(n3517) );
  XNOR2_X1 U4337 ( .A(IR_REG_28__SCAN_IN), .B(keyinput33), .ZN(n3516) );
  NAND4_X1 U4338 ( .A1(n3519), .A2(n3518), .A3(n3517), .A4(n3516), .ZN(n3520)
         );
  NOR4_X1 U4339 ( .A1(n3523), .A2(n3522), .A3(n3521), .A4(n3520), .ZN(n3537)
         );
  AOI22_X1 U4340 ( .A1(n2450), .A2(keyinput24), .B1(keyinput38), .B2(n3525), 
        .ZN(n3524) );
  OAI221_X1 U4341 ( .B1(n2450), .B2(keyinput24), .C1(n3525), .C2(keyinput38), 
        .A(n3524), .ZN(n3535) );
  XOR2_X1 U4342 ( .A(keyinput3), .B(n3526), .Z(n3529) );
  XOR2_X1 U4343 ( .A(keyinput21), .B(n3527), .Z(n3528) );
  NAND2_X1 U4344 ( .A1(n3529), .A2(n3528), .ZN(n3534) );
  AOI22_X1 U4345 ( .A1(n2083), .A2(keyinput26), .B1(keyinput50), .B2(n3751), 
        .ZN(n3530) );
  OAI221_X1 U4346 ( .B1(n2083), .B2(keyinput26), .C1(n3751), .C2(keyinput50), 
        .A(n3530), .ZN(n3533) );
  AOI22_X1 U4347 ( .A1(n3587), .A2(keyinput1), .B1(keyinput17), .B2(n2084), 
        .ZN(n3531) );
  OAI221_X1 U4348 ( .B1(n3587), .B2(keyinput1), .C1(n2084), .C2(keyinput17), 
        .A(n3531), .ZN(n3532) );
  NOR4_X1 U4349 ( .A1(n3535), .A2(n3534), .A3(n3533), .A4(n3532), .ZN(n3536)
         );
  AND4_X1 U4350 ( .A1(n3539), .A2(n3538), .A3(n3537), .A4(n3536), .ZN(n3562)
         );
  INV_X1 U4351 ( .A(REG2_REG_23__SCAN_IN), .ZN(n3542) );
  AOI22_X1 U4352 ( .A1(n3542), .A2(keyinput31), .B1(keyinput40), .B2(n3541), 
        .ZN(n3540) );
  OAI221_X1 U4353 ( .B1(n3542), .B2(keyinput31), .C1(n3541), .C2(keyinput40), 
        .A(n3540), .ZN(n3553) );
  INV_X1 U4354 ( .A(DATAI_27_), .ZN(n3592) );
  AOI22_X1 U4355 ( .A1(n3592), .A2(keyinput29), .B1(n3544), .B2(keyinput19), 
        .ZN(n3543) );
  OAI221_X1 U4356 ( .B1(n3592), .B2(keyinput29), .C1(n3544), .C2(keyinput19), 
        .A(n3543), .ZN(n3552) );
  INV_X1 U4357 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3546) );
  AOI22_X1 U4358 ( .A1(n2785), .A2(keyinput54), .B1(n3546), .B2(keyinput62), 
        .ZN(n3545) );
  OAI221_X1 U4359 ( .B1(n2785), .B2(keyinput54), .C1(n3546), .C2(keyinput62), 
        .A(n3545), .ZN(n3551) );
  INV_X1 U4360 ( .A(ADDR_REG_8__SCAN_IN), .ZN(n3549) );
  INV_X1 U4361 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3548) );
  AOI22_X1 U4362 ( .A1(n3549), .A2(keyinput58), .B1(n3548), .B2(keyinput41), 
        .ZN(n3547) );
  OAI221_X1 U4363 ( .B1(n3549), .B2(keyinput58), .C1(n3548), .C2(keyinput41), 
        .A(n3547), .ZN(n3550) );
  NOR4_X1 U4364 ( .A1(n3553), .A2(n3552), .A3(n3551), .A4(n3550), .ZN(n3561)
         );
  INV_X1 U4365 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n3555) );
  INV_X1 U4366 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n4562) );
  OAI22_X1 U4367 ( .A1(n3555), .A2(keyinput11), .B1(n4562), .B2(keyinput51), 
        .ZN(n3554) );
  AOI221_X1 U4368 ( .B1(n3555), .B2(keyinput11), .C1(keyinput51), .C2(n4562), 
        .A(n3554), .ZN(n3560) );
  OAI22_X1 U4369 ( .A1(n3558), .A2(keyinput2), .B1(n3557), .B2(keyinput5), 
        .ZN(n3556) );
  AOI221_X1 U4370 ( .B1(n3558), .B2(keyinput2), .C1(keyinput5), .C2(n3557), 
        .A(n3556), .ZN(n3559) );
  AND4_X1 U4371 ( .A1(n3562), .A2(n3561), .A3(n3560), .A4(n3559), .ZN(n3622)
         );
  AOI22_X1 U4372 ( .A1(n3639), .A2(keyinput43), .B1(keyinput57), .B2(n3593), 
        .ZN(n3563) );
  OAI221_X1 U4373 ( .B1(n3639), .B2(keyinput43), .C1(n3593), .C2(keyinput57), 
        .A(n3563), .ZN(n3574) );
  AOI22_X1 U4374 ( .A1(n3594), .A2(keyinput44), .B1(keyinput30), .B2(n3565), 
        .ZN(n3564) );
  OAI221_X1 U4375 ( .B1(n3594), .B2(keyinput44), .C1(n3565), .C2(keyinput30), 
        .A(n3564), .ZN(n3573) );
  AOI22_X1 U4376 ( .A1(n3567), .A2(keyinput59), .B1(n4410), .B2(keyinput18), 
        .ZN(n3566) );
  OAI221_X1 U4377 ( .B1(n3567), .B2(keyinput59), .C1(n4410), .C2(keyinput18), 
        .A(n3566), .ZN(n3572) );
  AOI22_X1 U4378 ( .A1(n3570), .A2(keyinput35), .B1(keyinput47), .B2(n3569), 
        .ZN(n3568) );
  OAI221_X1 U4379 ( .B1(n3570), .B2(keyinput35), .C1(n3569), .C2(keyinput47), 
        .A(n3568), .ZN(n3571) );
  NOR4_X1 U4380 ( .A1(n3574), .A2(n3573), .A3(n3572), .A4(n3571), .ZN(n3621)
         );
  AOI22_X1 U4381 ( .A1(n3278), .A2(keyinput10), .B1(n3576), .B2(keyinput39), 
        .ZN(n3575) );
  OAI221_X1 U4382 ( .B1(n3278), .B2(keyinput10), .C1(n3576), .C2(keyinput39), 
        .A(n3575), .ZN(n3585) );
  INV_X1 U4383 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4544) );
  AOI22_X1 U4384 ( .A1(n4544), .A2(keyinput27), .B1(keyinput6), .B2(n3578), 
        .ZN(n3577) );
  OAI221_X1 U4385 ( .B1(n4544), .B2(keyinput27), .C1(n3578), .C2(keyinput6), 
        .A(n3577), .ZN(n3584) );
  INV_X1 U4386 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4388) );
  AOI22_X1 U4387 ( .A1(n2769), .A2(keyinput8), .B1(keyinput42), .B2(n4388), 
        .ZN(n3579) );
  OAI221_X1 U4388 ( .B1(n2769), .B2(keyinput8), .C1(n4388), .C2(keyinput42), 
        .A(n3579), .ZN(n3583) );
  INV_X1 U4389 ( .A(DATAI_13_), .ZN(n4641) );
  AOI22_X1 U4390 ( .A1(n4641), .A2(keyinput61), .B1(n3581), .B2(keyinput34), 
        .ZN(n3580) );
  OAI221_X1 U4391 ( .B1(n4641), .B2(keyinput61), .C1(n3581), .C2(keyinput34), 
        .A(n3580), .ZN(n3582) );
  NOR4_X1 U4392 ( .A1(n3585), .A2(n3584), .A3(n3583), .A4(n3582), .ZN(n3620)
         );
  NAND4_X1 U4393 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(n4626), .ZN(n3601) );
  INV_X1 U4394 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3586) );
  NAND4_X1 U4395 ( .A1(n3548), .A2(n3546), .A3(n3586), .A4(DATAI_7_), .ZN(
        n3591) );
  NOR4_X1 U4396 ( .A1(REG2_REG_19__SCAN_IN), .A2(REG3_REG_23__SCAN_IN), .A3(
        REG2_REG_18__SCAN_IN), .A4(n3587), .ZN(n3588) );
  NAND3_X1 U4397 ( .A1(n4208), .A2(D_REG_1__SCAN_IN), .A3(n3588), .ZN(n3590)
         );
  INV_X1 U4398 ( .A(DATAI_1_), .ZN(n3589) );
  OR4_X1 U4399 ( .A1(n3591), .A2(n3590), .A3(REG2_REG_5__SCAN_IN), .A4(n3589), 
        .ZN(n3600) );
  NAND4_X1 U4400 ( .A1(REG3_REG_20__SCAN_IN), .A2(REG3_REG_18__SCAN_IN), .A3(
        REG2_REG_23__SCAN_IN), .A4(DATAI_30_), .ZN(n3599) );
  NOR3_X1 U4401 ( .A1(REG3_REG_14__SCAN_IN), .A2(ADDR_REG_1__SCAN_IN), .A3(
        n3592), .ZN(n3597) );
  NOR4_X1 U4402 ( .A1(DATAI_13_), .A2(ADDR_REG_11__SCAN_IN), .A3(n4544), .A4(
        n4388), .ZN(n3596) );
  NOR4_X1 U4403 ( .A1(REG0_REG_19__SCAN_IN), .A2(n3594), .A3(n3639), .A4(n3593), .ZN(n3595) );
  NAND4_X1 U4404 ( .A1(ADDR_REG_8__SCAN_IN), .A2(n3597), .A3(n3596), .A4(n3595), .ZN(n3598) );
  NOR4_X1 U4405 ( .A1(n3601), .A2(n3600), .A3(n3599), .A4(n3598), .ZN(n3617)
         );
  NOR4_X1 U4406 ( .A1(D_REG_26__SCAN_IN), .A2(REG3_REG_6__SCAN_IN), .A3(
        REG1_REG_9__SCAN_IN), .A4(n2450), .ZN(n3607) );
  NAND4_X1 U4407 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .A3(
        IR_REG_20__SCAN_IN), .A4(IR_REG_23__SCAN_IN), .ZN(n3605) );
  NAND2_X1 U4408 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n3603)
         );
  OR4_X1 U4409 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_21__SCAN_IN), .A3(
        IR_REG_4__SCAN_IN), .A4(DATAO_REG_27__SCAN_IN), .ZN(n3602) );
  NOR4_X1 U4410 ( .A1(n3605), .A2(n3604), .A3(n3603), .A4(n3602), .ZN(n3606)
         );
  NAND2_X1 U4411 ( .A1(n3607), .A2(n3606), .ZN(n3615) );
  NAND4_X1 U4412 ( .A1(REG0_REG_29__SCAN_IN), .A2(DATAI_26_), .A3(
        DATAO_REG_6__SCAN_IN), .A4(n3608), .ZN(n3614) );
  NAND4_X1 U4413 ( .A1(DATAO_REG_3__SCAN_IN), .A2(ADDR_REG_3__SCAN_IN), .A3(
        ADDR_REG_15__SCAN_IN), .A4(n3609), .ZN(n3613) );
  NOR4_X1 U4414 ( .A1(REG1_REG_29__SCAN_IN), .A2(REG0_REG_25__SCAN_IN), .A3(
        REG2_REG_24__SCAN_IN), .A4(n4410), .ZN(n3611) );
  NOR3_X1 U4415 ( .A1(DATAO_REG_25__SCAN_IN), .A2(DATAO_REG_22__SCAN_IN), .A3(
        DATAO_REG_23__SCAN_IN), .ZN(n3610) );
  NAND3_X1 U4416 ( .A1(n3611), .A2(DATAO_REG_17__SCAN_IN), .A3(n3610), .ZN(
        n3612) );
  NOR4_X1 U4417 ( .A1(n3615), .A2(n3614), .A3(n3613), .A4(n3612), .ZN(n3616)
         );
  AOI21_X1 U4418 ( .B1(n3617), .B2(n3616), .A(keyinput12), .ZN(n3618) );
  MUX2_X1 U4419 ( .A(n3618), .B(keyinput12), .S(IR_REG_26__SCAN_IN), .Z(n3619)
         );
  NAND4_X1 U4420 ( .A1(n3622), .A2(n3621), .A3(n3620), .A4(n3619), .ZN(n3636)
         );
  AOI211_X1 U4421 ( .C1(n3625), .C2(n3624), .A(n3782), .B(n3623), .ZN(n3634)
         );
  OAI22_X1 U4422 ( .A1(n3627), .A2(n3777), .B1(n3776), .B2(n3626), .ZN(n3633)
         );
  NAND2_X1 U4423 ( .A1(n3780), .A2(n3628), .ZN(n3630) );
  OAI211_X1 U4424 ( .C1(n3775), .C2(n3631), .A(n3630), .B(n3629), .ZN(n3632)
         );
  NOR3_X1 U4425 ( .A1(n3634), .A2(n3633), .A3(n3632), .ZN(n3635) );
  XOR2_X1 U4426 ( .A(n3636), .B(n3635), .Z(U3214) );
  XOR2_X1 U4427 ( .A(n3638), .B(n3637), .Z(n3644) );
  AOI22_X1 U4428 ( .A1(n3749), .A2(n4173), .B1(n3750), .B2(n4129), .ZN(n3643)
         );
  NOR2_X1 U4429 ( .A1(n3639), .A2(STATE_REG_SCAN_IN), .ZN(n4520) );
  NOR2_X1 U4430 ( .A1(n3775), .A2(n3640), .ZN(n3641) );
  AOI211_X1 U4431 ( .C1(n4163), .C2(n3780), .A(n4520), .B(n3641), .ZN(n3642)
         );
  OAI211_X1 U4432 ( .C1(n3644), .C2(n3782), .A(n3643), .B(n3642), .ZN(U3216)
         );
  XNOR2_X1 U4433 ( .A(n3646), .B(n3645), .ZN(n3647) );
  XNOR2_X1 U4434 ( .A(n3648), .B(n3647), .ZN(n3654) );
  OAI22_X1 U4435 ( .A1(n3775), .A2(n3650), .B1(STATE_REG_SCAN_IN), .B2(n3649), 
        .ZN(n3652) );
  OAI22_X1 U4436 ( .A1(n4131), .A2(n3776), .B1(n4175), .B2(n3777), .ZN(n3651)
         );
  AOI211_X1 U4437 ( .C1(n4126), .C2(n3780), .A(n3652), .B(n3651), .ZN(n3653)
         );
  OAI21_X1 U4438 ( .B1(n3654), .B2(n3782), .A(n3653), .ZN(U3220) );
  NOR2_X1 U4439 ( .A1(n3656), .A2(n2117), .ZN(n3657) );
  XNOR2_X1 U4440 ( .A(n3658), .B(n3657), .ZN(n3665) );
  INV_X1 U4441 ( .A(n3659), .ZN(n4059) );
  OAI22_X1 U4442 ( .A1(n3775), .A2(n3661), .B1(STATE_REG_SCAN_IN), .B2(n3660), 
        .ZN(n3663) );
  OAI22_X1 U4443 ( .A1(n4067), .A2(n3776), .B1(n4102), .B2(n3777), .ZN(n3662)
         );
  AOI211_X1 U4444 ( .C1(n4059), .C2(n3780), .A(n3663), .B(n3662), .ZN(n3664)
         );
  OAI21_X1 U4445 ( .B1(n3665), .B2(n3782), .A(n3664), .ZN(U3222) );
  INV_X1 U4446 ( .A(n3771), .ZN(n3678) );
  INV_X1 U4447 ( .A(n3666), .ZN(n3668) );
  NAND2_X1 U4448 ( .A1(n3668), .A2(n3667), .ZN(n3768) );
  NOR2_X1 U4449 ( .A1(n3668), .A2(n3667), .ZN(n3770) );
  AOI21_X1 U4450 ( .B1(n3678), .B2(n3768), .A(n3770), .ZN(n3670) );
  XNOR2_X1 U4451 ( .A(n3669), .B(n3681), .ZN(n3677) );
  XNOR2_X1 U4452 ( .A(n3670), .B(n3677), .ZN(n3676) );
  NAND2_X1 U4453 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4564) );
  OAI21_X1 U4454 ( .B1(n3775), .B2(n3671), .A(n4564), .ZN(n3674) );
  OAI22_X1 U4455 ( .A1(n4217), .A2(n3776), .B1(n3777), .B2(n3672), .ZN(n3673)
         );
  AOI211_X1 U4456 ( .C1(n4220), .C2(n3780), .A(n3674), .B(n3673), .ZN(n3675)
         );
  OAI21_X1 U4457 ( .B1(n3676), .B2(n3782), .A(n3675), .ZN(U3223) );
  OAI211_X1 U4458 ( .C1(n3770), .C2(n3678), .A(n3677), .B(n3768), .ZN(n3679)
         );
  OAI21_X1 U4459 ( .B1(n3681), .B2(n3680), .A(n3679), .ZN(n3685) );
  XNOR2_X1 U4460 ( .A(n3683), .B(n3682), .ZN(n3684) );
  XNOR2_X1 U4461 ( .A(n3685), .B(n3684), .ZN(n3689) );
  AOI22_X1 U4462 ( .A1(n3750), .A2(n4173), .B1(n3749), .B2(n4203), .ZN(n3688)
         );
  AND2_X1 U4463 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4576) );
  NOR2_X1 U4464 ( .A1(n3752), .A2(n4199), .ZN(n3686) );
  AOI211_X1 U4465 ( .C1(n4202), .C2(n3754), .A(n4576), .B(n3686), .ZN(n3687)
         );
  OAI211_X1 U4466 ( .C1(n3689), .C2(n3782), .A(n3688), .B(n3687), .ZN(U3225)
         );
  NAND2_X1 U4467 ( .A1(n3691), .A2(n3692), .ZN(n3693) );
  XOR2_X1 U4468 ( .A(n3694), .B(n3693), .Z(n3700) );
  INV_X1 U4469 ( .A(n3695), .ZN(n4083) );
  OAI22_X1 U4470 ( .A1(n3775), .A2(n4080), .B1(STATE_REG_SCAN_IN), .B2(n3696), 
        .ZN(n3698) );
  OAI22_X1 U4471 ( .A1(n4045), .A2(n3776), .B1(n4115), .B2(n3777), .ZN(n3697)
         );
  AOI211_X1 U4472 ( .C1(n4083), .C2(n3780), .A(n3698), .B(n3697), .ZN(n3699)
         );
  OAI21_X1 U4473 ( .B1(n3700), .B2(n3782), .A(n3699), .ZN(U3226) );
  INV_X1 U4474 ( .A(n3701), .ZN(n3706) );
  AOI21_X1 U4475 ( .B1(n3705), .B2(n3703), .A(n3702), .ZN(n3704) );
  AOI21_X1 U4476 ( .B1(n3706), .B2(n3705), .A(n3704), .ZN(n3711) );
  INV_X1 U4477 ( .A(n4156), .ZN(n3709) );
  OAI22_X1 U4478 ( .A1(n3775), .A2(n4147), .B1(STATE_REG_SCAN_IN), .B2(n2083), 
        .ZN(n3708) );
  OAI22_X1 U4479 ( .A1(n3724), .A2(n3776), .B1(n3777), .B2(n4187), .ZN(n3707)
         );
  AOI211_X1 U4480 ( .C1(n3709), .C2(n3780), .A(n3708), .B(n3707), .ZN(n3710)
         );
  OAI21_X1 U4481 ( .B1(n3711), .B2(n3782), .A(n3710), .ZN(U3230) );
  XNOR2_X1 U4482 ( .A(n3713), .B(n3712), .ZN(n3714) );
  XNOR2_X1 U4483 ( .A(n3715), .B(n3714), .ZN(n3719) );
  AOI22_X1 U4484 ( .A1(n3749), .A2(n4274), .B1(n3750), .B2(n4277), .ZN(n3718)
         );
  AND2_X1 U4485 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n4541) );
  NOR2_X1 U4486 ( .A1(n3775), .A2(n4285), .ZN(n3716) );
  AOI211_X1 U4487 ( .C1(n4286), .C2(n3780), .A(n4541), .B(n3716), .ZN(n3717)
         );
  OAI211_X1 U4488 ( .C1(n3719), .C2(n3782), .A(n3718), .B(n3717), .ZN(U3231)
         );
  AOI21_X1 U4489 ( .B1(n3722), .B2(n3721), .A(n3720), .ZN(n3728) );
  OAI22_X1 U4490 ( .A1(n3775), .A2(n4112), .B1(STATE_REG_SCAN_IN), .B2(n3723), 
        .ZN(n3726) );
  OAI22_X1 U4491 ( .A1(n4115), .A2(n3776), .B1(n3724), .B2(n3777), .ZN(n3725)
         );
  AOI211_X1 U4492 ( .C1(n4118), .C2(n3780), .A(n3726), .B(n3725), .ZN(n3727)
         );
  OAI21_X1 U4493 ( .B1(n3728), .B2(n3782), .A(n3727), .ZN(U3232) );
  OAI21_X1 U4494 ( .B1(n3730), .B2(n3732), .A(n3731), .ZN(n3734) );
  NAND2_X1 U4495 ( .A1(n3734), .A2(n3733), .ZN(n3740) );
  AOI22_X1 U4496 ( .A1(n3754), .A2(n3736), .B1(REG3_REG_2__SCAN_IN), .B2(n3735), .ZN(n3739) );
  AOI22_X1 U4497 ( .A1(n3750), .A2(n3737), .B1(n3749), .B2(n2868), .ZN(n3738)
         );
  NAND3_X1 U4498 ( .A1(n3740), .A2(n3739), .A3(n3738), .ZN(U3234) );
  NAND2_X1 U4499 ( .A1(n3742), .A2(n3741), .ZN(n3748) );
  AND2_X1 U4500 ( .A1(n3666), .A2(n3743), .ZN(n3746) );
  OAI21_X1 U4501 ( .B1(n3746), .B2(n3745), .A(n3744), .ZN(n3747) );
  XOR2_X1 U4502 ( .A(n3748), .B(n3747), .Z(n3757) );
  AOI22_X1 U4503 ( .A1(n3750), .A2(n3946), .B1(n3749), .B2(n4185), .ZN(n3756)
         );
  NOR2_X1 U4504 ( .A1(n3751), .A2(STATE_REG_SCAN_IN), .ZN(n4594) );
  NOR2_X1 U4505 ( .A1(n3752), .A2(n4193), .ZN(n3753) );
  AOI211_X1 U4506 ( .C1(n4184), .C2(n3754), .A(n4594), .B(n3753), .ZN(n3755)
         );
  OAI211_X1 U4507 ( .C1(n3757), .C2(n3782), .A(n3756), .B(n3755), .ZN(U3235)
         );
  NAND2_X1 U4508 ( .A1(n3760), .A2(n3759), .ZN(n3761) );
  XNOR2_X1 U4509 ( .A(n3758), .B(n3761), .ZN(n3767) );
  OAI22_X1 U4510 ( .A1(n3775), .A2(n4051), .B1(STATE_REG_SCAN_IN), .B2(n3762), 
        .ZN(n3765) );
  OAI22_X1 U4511 ( .A1(n3763), .A2(n3776), .B1(n4045), .B2(n3777), .ZN(n3764)
         );
  AOI211_X1 U4512 ( .C1(n4052), .C2(n3780), .A(n3765), .B(n3764), .ZN(n3766)
         );
  OAI21_X1 U4513 ( .B1(n3767), .B2(n3782), .A(n3766), .ZN(U3237) );
  INV_X1 U4514 ( .A(n3768), .ZN(n3769) );
  NOR2_X1 U4515 ( .A1(n3770), .A2(n3769), .ZN(n3772) );
  XNOR2_X1 U4516 ( .A(n3772), .B(n3771), .ZN(n3783) );
  INV_X1 U4517 ( .A(n3773), .ZN(n4239) );
  NAND2_X1 U4518 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4560) );
  OAI21_X1 U4519 ( .B1(n3775), .B2(n3774), .A(n4560), .ZN(n3779) );
  OAI22_X1 U4520 ( .A1(n4228), .A2(n3777), .B1(n3776), .B2(n4229), .ZN(n3778)
         );
  AOI211_X1 U4521 ( .C1(n4239), .C2(n3780), .A(n3779), .B(n3778), .ZN(n3781)
         );
  OAI21_X1 U4522 ( .B1(n3783), .B2(n3782), .A(n3781), .ZN(U3238) );
  INV_X1 U4523 ( .A(n3784), .ZN(n3787) );
  OAI211_X1 U4524 ( .C1(n3787), .C2(n3931), .A(n3786), .B(n3785), .ZN(n3790)
         );
  NAND3_X1 U4525 ( .A1(n3790), .A2(n3789), .A3(n3788), .ZN(n3793) );
  NAND3_X1 U4526 ( .A1(n3793), .A2(n3792), .A3(n3791), .ZN(n3796) );
  NAND3_X1 U4527 ( .A1(n3796), .A2(n3795), .A3(n3794), .ZN(n3799) );
  NAND3_X1 U4528 ( .A1(n3799), .A2(n3798), .A3(n3797), .ZN(n3803) );
  INV_X1 U4529 ( .A(n3800), .ZN(n3801) );
  AOI21_X1 U4530 ( .B1(n3803), .B2(n3802), .A(n3801), .ZN(n3809) );
  NAND2_X1 U4531 ( .A1(n3805), .A2(n3804), .ZN(n3808) );
  OAI211_X1 U4532 ( .C1(n3809), .C2(n3808), .A(n3807), .B(n3806), .ZN(n3812)
         );
  AND3_X1 U4533 ( .A1(n3812), .A2(n3811), .A3(n3810), .ZN(n3815) );
  OAI21_X1 U4534 ( .B1(n3815), .B2(n3814), .A(n3813), .ZN(n3818) );
  NAND4_X1 U4535 ( .A1(n3818), .A2(n2008), .A3(n3817), .A4(n3816), .ZN(n3821)
         );
  NAND2_X1 U4536 ( .A1(n3824), .A2(n4232), .ZN(n3902) );
  INV_X1 U4537 ( .A(n3902), .ZN(n3819) );
  NAND3_X1 U4538 ( .A1(n3821), .A2(n3820), .A3(n3819), .ZN(n3827) );
  INV_X1 U4539 ( .A(n3822), .ZN(n3826) );
  INV_X1 U4540 ( .A(n3823), .ZN(n3825) );
  OAI21_X1 U4541 ( .B1(n3826), .B2(n3825), .A(n3824), .ZN(n3901) );
  NAND3_X1 U4542 ( .A1(n3827), .A2(n3903), .A3(n3901), .ZN(n3828) );
  AOI21_X1 U4543 ( .B1(n3828), .B2(n3905), .A(n3904), .ZN(n3830) );
  INV_X1 U4544 ( .A(n3829), .ZN(n3908) );
  INV_X1 U4545 ( .A(n4092), .ZN(n3863) );
  OAI211_X1 U4546 ( .C1(n3830), .C2(n3908), .A(n3907), .B(n3863), .ZN(n3833)
         );
  INV_X1 U4547 ( .A(n3831), .ZN(n3832) );
  AOI21_X1 U4548 ( .B1(n3833), .B2(n3912), .A(n3832), .ZN(n3834) );
  OR2_X1 U4549 ( .A1(n3861), .A2(n2257), .ZN(n3915) );
  OAI21_X1 U4550 ( .B1(n3834), .B2(n3915), .A(n3914), .ZN(n3841) );
  INV_X1 U4551 ( .A(n3835), .ZN(n3852) );
  INV_X1 U4552 ( .A(n3836), .ZN(n3837) );
  AOI21_X1 U4553 ( .B1(n3943), .B2(n3852), .A(n3837), .ZN(n3921) );
  INV_X1 U4554 ( .A(n3921), .ZN(n3840) );
  NAND2_X1 U4555 ( .A1(n3838), .A2(n3920), .ZN(n3839) );
  AOI211_X1 U4556 ( .C1(n3841), .C2(n3917), .A(n3840), .B(n3839), .ZN(n3859)
         );
  NAND2_X1 U4557 ( .A1(n3843), .A2(n3842), .ZN(n3919) );
  INV_X1 U4558 ( .A(n3942), .ZN(n3844) );
  AND2_X1 U4559 ( .A1(n3850), .A2(DATAI_30_), .ZN(n4005) );
  NAND2_X1 U4560 ( .A1(n3844), .A2(n4005), .ZN(n3851) );
  NAND2_X1 U4561 ( .A1(n2432), .A2(REG1_REG_31__SCAN_IN), .ZN(n3849) );
  NAND2_X1 U4562 ( .A1(n3845), .A2(REG2_REG_31__SCAN_IN), .ZN(n3848) );
  NAND2_X1 U4563 ( .A1(n3846), .A2(REG0_REG_31__SCAN_IN), .ZN(n3847) );
  NAND3_X1 U4564 ( .A1(n3849), .A2(n3848), .A3(n3847), .ZN(n3999) );
  NAND2_X1 U4565 ( .A1(n3850), .A2(DATAI_31_), .ZN(n4000) );
  NAND2_X1 U4566 ( .A1(n3999), .A2(n4000), .ZN(n3853) );
  AND2_X1 U4567 ( .A1(n3851), .A2(n3853), .ZN(n3871) );
  OAI21_X1 U4568 ( .B1(n3943), .B2(n3852), .A(n3871), .ZN(n3918) );
  AOI21_X1 U4569 ( .B1(n3921), .B2(n3919), .A(n3918), .ZN(n3923) );
  INV_X1 U4570 ( .A(n3923), .ZN(n3858) );
  INV_X1 U4571 ( .A(n3853), .ZN(n3857) );
  INV_X1 U4572 ( .A(n3999), .ZN(n3927) );
  INV_X1 U4573 ( .A(n4000), .ZN(n3854) );
  NAND2_X1 U4574 ( .A1(n3927), .A2(n3854), .ZN(n3856) );
  INV_X1 U4575 ( .A(n4005), .ZN(n3855) );
  NAND2_X1 U4576 ( .A1(n3942), .A2(n3855), .ZN(n3928) );
  AND2_X1 U4577 ( .A1(n3856), .A2(n3928), .ZN(n3872) );
  OAI22_X1 U4578 ( .A1(n3859), .A2(n3858), .B1(n3857), .B2(n3872), .ZN(n3933)
         );
  INV_X1 U4579 ( .A(n3860), .ZN(n3900) );
  INV_X1 U4580 ( .A(n4060), .ZN(n3862) );
  OR2_X1 U4581 ( .A1(n3862), .A2(n3861), .ZN(n4074) );
  INV_X1 U4582 ( .A(n4074), .ZN(n3897) );
  NAND2_X1 U4583 ( .A1(n3865), .A2(n3864), .ZN(n4098) );
  AND2_X1 U4584 ( .A1(n3867), .A2(n3866), .ZN(n4142) );
  INV_X1 U4585 ( .A(n4142), .ZN(n4145) );
  INV_X1 U4586 ( .A(n3868), .ZN(n4231) );
  NAND2_X1 U4587 ( .A1(n4140), .A2(n4139), .ZN(n4171) );
  AND2_X1 U4588 ( .A1(n4041), .A2(n3870), .ZN(n4063) );
  NAND4_X1 U4589 ( .A1(n4044), .A2(n4063), .A3(n3872), .A4(n3871), .ZN(n3873)
         );
  NOR2_X1 U4590 ( .A1(n3874), .A2(n3873), .ZN(n3889) );
  NOR2_X1 U4591 ( .A1(n3876), .A2(n3875), .ZN(n3888) );
  INV_X1 U4592 ( .A(n3877), .ZN(n3879) );
  NAND4_X1 U4593 ( .A1(n3881), .A2(n3880), .A3(n3879), .A4(n3878), .ZN(n3886)
         );
  NAND4_X1 U4594 ( .A1(n4302), .A2(n3884), .A3(n3883), .A4(n3882), .ZN(n3885)
         );
  NOR2_X1 U4595 ( .A1(n3886), .A2(n3885), .ZN(n3887) );
  NAND2_X1 U4596 ( .A1(n3891), .A2(n3890), .ZN(n4272) );
  NOR2_X1 U4597 ( .A1(n4183), .A2(n4272), .ZN(n3895) );
  INV_X1 U4598 ( .A(n4166), .ZN(n3892) );
  NAND2_X1 U4599 ( .A1(n3892), .A2(n4165), .ZN(n4201) );
  NOR2_X1 U4600 ( .A1(n4201), .A2(n4619), .ZN(n3894) );
  NAND3_X1 U4601 ( .A1(n3897), .A2(n4127), .A3(n3896), .ZN(n3898) );
  OAI21_X1 U4602 ( .B1(n4247), .B2(n3902), .A(n3901), .ZN(n3906) );
  AOI211_X1 U4603 ( .C1(n3906), .C2(n3905), .A(n2259), .B(n3904), .ZN(n3909)
         );
  OAI21_X1 U4604 ( .B1(n3909), .B2(n3908), .A(n3907), .ZN(n3913) );
  INV_X1 U4605 ( .A(n3910), .ZN(n3911) );
  AOI21_X1 U4606 ( .B1(n3913), .B2(n3912), .A(n3911), .ZN(n3916) );
  OAI21_X1 U4607 ( .B1(n3916), .B2(n3915), .A(n3914), .ZN(n3925) );
  NOR3_X1 U4608 ( .A1(n3919), .A2(n2254), .A3(n3918), .ZN(n3924) );
  NAND3_X1 U4609 ( .A1(n3921), .A2(n2632), .A3(n3920), .ZN(n3922) );
  AOI22_X1 U4610 ( .A1(n3925), .A2(n3924), .B1(n3923), .B2(n3922), .ZN(n3926)
         );
  AOI21_X1 U4611 ( .B1(n4005), .B2(n3927), .A(n3926), .ZN(n3930) );
  AOI21_X1 U4612 ( .B1(n3928), .B2(n3999), .A(n4000), .ZN(n3929) );
  OR2_X1 U4613 ( .A1(n3930), .A2(n3929), .ZN(n3932) );
  XNOR2_X1 U4614 ( .A(n3934), .B(n2865), .ZN(n3941) );
  NOR4_X1 U4615 ( .A1(n4631), .A2(n3936), .A3(n3960), .A4(n3935), .ZN(n3937)
         );
  NAND2_X1 U4616 ( .A1(n3937), .A2(n3263), .ZN(n3938) );
  OAI211_X1 U4617 ( .C1(n4482), .C2(n3940), .A(n3938), .B(B_REG_SCAN_IN), .ZN(
        n3939) );
  OAI21_X1 U4618 ( .B1(n3941), .B2(n3940), .A(n3939), .ZN(U3239) );
  MUX2_X1 U4619 ( .A(n3999), .B(DATAO_REG_31__SCAN_IN), .S(n3955), .Z(U3581)
         );
  MUX2_X1 U4620 ( .A(n3942), .B(DATAO_REG_30__SCAN_IN), .S(n3955), .Z(U3580)
         );
  MUX2_X1 U4621 ( .A(n3943), .B(DATAO_REG_29__SCAN_IN), .S(n3955), .Z(U3579)
         );
  MUX2_X1 U4622 ( .A(n3944), .B(DATAO_REG_28__SCAN_IN), .S(n3955), .Z(U3578)
         );
  MUX2_X1 U4623 ( .A(n3945), .B(DATAO_REG_26__SCAN_IN), .S(n3955), .Z(U3576)
         );
  MUX2_X1 U4624 ( .A(n4065), .B(DATAO_REG_24__SCAN_IN), .S(n3955), .Z(U3574)
         );
  MUX2_X1 U4625 ( .A(n4149), .B(DATAO_REG_21__SCAN_IN), .S(n3955), .Z(U3571)
         );
  MUX2_X1 U4626 ( .A(n4129), .B(DATAO_REG_20__SCAN_IN), .S(n3955), .Z(U3570)
         );
  MUX2_X1 U4627 ( .A(DATAO_REG_19__SCAN_IN), .B(n3946), .S(U4043), .Z(U3569)
         );
  MUX2_X1 U4628 ( .A(DATAO_REG_18__SCAN_IN), .B(n4173), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4629 ( .A(DATAO_REG_16__SCAN_IN), .B(n4203), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4630 ( .A(n4250), .B(DATAO_REG_15__SCAN_IN), .S(n3955), .Z(U3565)
         );
  MUX2_X1 U4631 ( .A(DATAO_REG_14__SCAN_IN), .B(n4277), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4632 ( .A(n4249), .B(DATAO_REG_13__SCAN_IN), .S(n3955), .Z(U3563)
         );
  MUX2_X1 U4633 ( .A(n4274), .B(DATAO_REG_12__SCAN_IN), .S(n3955), .Z(U3562)
         );
  MUX2_X1 U4634 ( .A(DATAO_REG_11__SCAN_IN), .B(n3947), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4635 ( .A(n3948), .B(DATAO_REG_10__SCAN_IN), .S(n3955), .Z(U3560)
         );
  MUX2_X1 U4636 ( .A(n3949), .B(DATAO_REG_9__SCAN_IN), .S(n3955), .Z(U3559) );
  MUX2_X1 U4637 ( .A(DATAO_REG_8__SCAN_IN), .B(n3950), .S(U4043), .Z(U3558) );
  MUX2_X1 U4638 ( .A(DATAO_REG_7__SCAN_IN), .B(n3951), .S(U4043), .Z(U3557) );
  MUX2_X1 U4639 ( .A(DATAO_REG_5__SCAN_IN), .B(n3952), .S(U4043), .Z(U3555) );
  MUX2_X1 U4640 ( .A(DATAO_REG_4__SCAN_IN), .B(n3953), .S(U4043), .Z(U3554) );
  MUX2_X1 U4641 ( .A(DATAO_REG_2__SCAN_IN), .B(n3954), .S(U4043), .Z(U3552) );
  MUX2_X1 U4642 ( .A(DATAO_REG_1__SCAN_IN), .B(n2868), .S(U4043), .Z(U3551) );
  MUX2_X1 U4643 ( .A(n3956), .B(DATAO_REG_0__SCAN_IN), .S(n3955), .Z(U3550) );
  INV_X1 U4644 ( .A(n3957), .ZN(n3958) );
  NAND2_X1 U4645 ( .A1(n3958), .A2(n3960), .ZN(n3959) );
  OAI211_X1 U4646 ( .C1(n3961), .C2(n3960), .A(n3959), .B(n4479), .ZN(n3962)
         );
  OAI211_X1 U4647 ( .C1(IR_REG_0__SCAN_IN), .C2(n3963), .A(n3962), .B(U4043), 
        .ZN(n4536) );
  AOI22_X1 U4648 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4595), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3972) );
  XOR2_X1 U4649 ( .A(n3964), .B(n3965), .Z(n3966) );
  AOI22_X1 U4650 ( .A1(n4493), .A2(n4559), .B1(n4584), .B2(n3966), .ZN(n3971)
         );
  OAI211_X1 U4651 ( .C1(n3969), .C2(n3968), .A(n4586), .B(n3967), .ZN(n3970)
         );
  NAND4_X1 U4652 ( .A1(n4536), .A2(n3972), .A3(n3971), .A4(n3970), .ZN(U3242)
         );
  XOR2_X1 U4653 ( .A(REG2_REG_12__SCAN_IN), .B(n3986), .Z(n3983) );
  INV_X1 U4654 ( .A(n3975), .ZN(n3977) );
  NOR2_X1 U4655 ( .A1(n4604), .A2(n2157), .ZN(n3976) );
  AOI211_X1 U4656 ( .C1(n4595), .C2(ADDR_REG_12__SCAN_IN), .A(n3977), .B(n3976), .ZN(n3982) );
  XNOR2_X1 U4657 ( .A(n3989), .B(n2157), .ZN(n3980) );
  OAI211_X1 U4658 ( .C1(n3980), .C2(REG1_REG_12__SCAN_IN), .A(n3991), .B(n4584), .ZN(n3981) );
  OAI211_X1 U4659 ( .C1(n3983), .C2(n4596), .A(n3982), .B(n3981), .ZN(U3252)
         );
  INV_X1 U4660 ( .A(n3992), .ZN(n4642) );
  NOR2_X1 U4661 ( .A1(n4544), .A2(n4642), .ZN(n4543) );
  OAI211_X1 U4662 ( .C1(n3987), .C2(REG2_REG_14__SCAN_IN), .A(n4499), .B(n4586), .ZN(n3997) );
  AOI21_X1 U4663 ( .B1(n4595), .B2(ADDR_REG_14__SCAN_IN), .A(n3988), .ZN(n3996) );
  NAND2_X1 U4664 ( .A1(n3989), .A2(n4485), .ZN(n3990) );
  INV_X1 U4665 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4382) );
  AOI22_X1 U4666 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4642), .B1(n3992), .B2(
        n4382), .ZN(n4539) );
  OAI211_X1 U4667 ( .C1(n3993), .C2(REG1_REG_14__SCAN_IN), .A(n4515), .B(n4584), .ZN(n3995) );
  NAND2_X1 U4668 ( .A1(n4559), .A2(n4512), .ZN(n3994) );
  NAND4_X1 U4669 ( .A1(n3997), .A2(n3996), .A3(n3995), .A4(n3994), .ZN(U3254)
         );
  NAND2_X1 U4670 ( .A1(n3999), .A2(n3998), .ZN(n4007) );
  OAI21_X1 U4671 ( .B1(n4000), .B2(n4279), .A(n4007), .ZN(n4396) );
  NAND2_X1 U4672 ( .A1(n4289), .A2(n4396), .ZN(n4002) );
  NAND2_X1 U4673 ( .A1(n4623), .A2(REG2_REG_31__SCAN_IN), .ZN(n4001) );
  OAI211_X1 U4674 ( .C1(n4399), .C2(n4317), .A(n4002), .B(n4001), .ZN(U3260)
         );
  INV_X1 U4675 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4010) );
  NAND2_X1 U4676 ( .A1(n4400), .A2(n4608), .ZN(n4009) );
  NAND2_X1 U4677 ( .A1(n4005), .A2(n4306), .ZN(n4006) );
  NAND2_X1 U4678 ( .A1(n4007), .A2(n4006), .ZN(n4401) );
  NAND2_X1 U4679 ( .A1(n4289), .A2(n4401), .ZN(n4008) );
  OAI211_X1 U4680 ( .C1(n4289), .C2(n4010), .A(n4009), .B(n4008), .ZN(U3261)
         );
  OAI21_X1 U4681 ( .B1(n4012), .B2(n4287), .A(n4011), .ZN(n4016) );
  INV_X1 U4682 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4013) );
  OAI22_X1 U4683 ( .A1(n4014), .A2(n4317), .B1(n4013), .B2(n4289), .ZN(n4015)
         );
  OAI21_X1 U4684 ( .B1(n4018), .B2(n4242), .A(n4017), .ZN(U3354) );
  NAND2_X1 U4685 ( .A1(n4019), .A2(n4029), .ZN(n4020) );
  NAND2_X1 U4686 ( .A1(n4021), .A2(n4020), .ZN(n4027) );
  OAI22_X1 U4687 ( .A1(n4067), .A2(n4296), .B1(n4022), .B2(n4279), .ZN(n4023)
         );
  INV_X1 U4688 ( .A(n4023), .ZN(n4024) );
  OAI21_X1 U4689 ( .B1(n4025), .B2(n4298), .A(n4024), .ZN(n4026) );
  AOI21_X1 U4690 ( .B1(n4027), .B2(n4281), .A(n4026), .ZN(n4328) );
  XOR2_X1 U4691 ( .A(n4029), .B(n4028), .Z(n4408) );
  INV_X1 U4692 ( .A(n4408), .ZN(n4031) );
  NAND2_X1 U4693 ( .A1(n4031), .A2(n4030), .ZN(n4039) );
  AND2_X1 U4694 ( .A1(n4050), .A2(n4032), .ZN(n4033) );
  NOR2_X1 U4695 ( .A1(n4034), .A2(n4033), .ZN(n4326) );
  OAI22_X1 U4696 ( .A1(n4036), .A2(n4287), .B1(n4035), .B2(n4289), .ZN(n4037)
         );
  AOI21_X1 U4697 ( .B1(n4326), .B2(n4608), .A(n4037), .ZN(n4038) );
  OAI211_X1 U4698 ( .C1(n4623), .C2(n4328), .A(n4039), .B(n4038), .ZN(U3263)
         );
  XNOR2_X1 U4699 ( .A(n4040), .B(n4044), .ZN(n4332) );
  INV_X1 U4700 ( .A(n4332), .ZN(n4056) );
  NAND2_X1 U4701 ( .A1(n4042), .A2(n4041), .ZN(n4043) );
  XOR2_X1 U4702 ( .A(n4044), .B(n4043), .Z(n4049) );
  OAI22_X1 U4703 ( .A1(n4045), .A2(n4296), .B1(n4051), .B2(n4279), .ZN(n4046)
         );
  AOI21_X1 U4704 ( .B1(n4276), .B2(n4047), .A(n4046), .ZN(n4048) );
  OAI21_X1 U4705 ( .B1(n4049), .B2(n4309), .A(n4048), .ZN(n4331) );
  OAI21_X1 U4706 ( .B1(n2021), .B2(n4051), .A(n4050), .ZN(n4412) );
  AOI22_X1 U4707 ( .A1(n4052), .A2(n4618), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4623), .ZN(n4053) );
  OAI21_X1 U4708 ( .B1(n4412), .B2(n4317), .A(n4053), .ZN(n4054) );
  AOI21_X1 U4709 ( .B1(n4331), .B2(n4289), .A(n4054), .ZN(n4055) );
  OAI21_X1 U4710 ( .B1(n4056), .B2(n4242), .A(n4055), .ZN(U3264) );
  XNOR2_X1 U4711 ( .A(n4057), .B(n4063), .ZN(n4417) );
  INV_X1 U4712 ( .A(n4082), .ZN(n4058) );
  AOI21_X1 U4713 ( .B1(n4064), .B2(n4058), .A(n2021), .ZN(n4415) );
  AOI22_X1 U4714 ( .A1(n4415), .A2(n4608), .B1(n4059), .B2(n4618), .ZN(n4072)
         );
  INV_X1 U4715 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4070) );
  NAND2_X1 U4716 ( .A1(n4061), .A2(n4060), .ZN(n4062) );
  XOR2_X1 U4717 ( .A(n4063), .B(n4062), .Z(n4069) );
  AOI22_X1 U4718 ( .A1(n4065), .A2(n4275), .B1(n4064), .B2(n4306), .ZN(n4066)
         );
  OAI21_X1 U4719 ( .B1(n4067), .B2(n4298), .A(n4066), .ZN(n4068) );
  AOI21_X1 U4720 ( .B1(n4069), .B2(n4281), .A(n4068), .ZN(n4335) );
  MUX2_X1 U4721 ( .A(n4070), .B(n4335), .S(n4289), .Z(n4071) );
  OAI211_X1 U4722 ( .C1(n4417), .C2(n4242), .A(n4072), .B(n4071), .ZN(U3265)
         );
  XNOR2_X1 U4723 ( .A(n4073), .B(n4074), .ZN(n4339) );
  INV_X1 U4724 ( .A(n4339), .ZN(n4087) );
  XNOR2_X1 U4725 ( .A(n4075), .B(n4074), .ZN(n4079) );
  OAI22_X1 U4726 ( .A1(n4115), .A2(n4296), .B1(n4080), .B2(n4279), .ZN(n4076)
         );
  AOI21_X1 U4727 ( .B1(n4077), .B2(n4276), .A(n4076), .ZN(n4078) );
  OAI21_X1 U4728 ( .B1(n4079), .B2(n4309), .A(n4078), .ZN(n4338) );
  NOR2_X1 U4729 ( .A1(n4089), .A2(n4080), .ZN(n4081) );
  OR2_X1 U4730 ( .A1(n4082), .A2(n4081), .ZN(n4421) );
  AOI22_X1 U4731 ( .A1(n4083), .A2(n4618), .B1(REG2_REG_24__SCAN_IN), .B2(
        n4623), .ZN(n4084) );
  OAI21_X1 U4732 ( .B1(n4421), .B2(n4317), .A(n4084), .ZN(n4085) );
  AOI21_X1 U4733 ( .B1(n4338), .B2(n4289), .A(n4085), .ZN(n4086) );
  OAI21_X1 U4734 ( .B1(n4087), .B2(n4242), .A(n4086), .ZN(U3266) );
  XNOR2_X1 U4735 ( .A(n4088), .B(n4098), .ZN(n4426) );
  AOI21_X1 U4736 ( .B1(n4099), .B2(n4346), .A(n4089), .ZN(n4424) );
  AOI22_X1 U4737 ( .A1(n4424), .A2(n4608), .B1(n4090), .B2(n4618), .ZN(n4106)
         );
  OR2_X1 U4738 ( .A1(n4091), .A2(n4092), .ZN(n4094) );
  NAND2_X1 U4739 ( .A1(n4094), .A2(n4093), .ZN(n4111) );
  INV_X1 U4740 ( .A(n4111), .ZN(n4096) );
  OAI21_X1 U4741 ( .B1(n4096), .B2(n4109), .A(n4095), .ZN(n4097) );
  XOR2_X1 U4742 ( .A(n4098), .B(n4097), .Z(n4104) );
  AOI22_X1 U4743 ( .A1(n4100), .A2(n4275), .B1(n4306), .B2(n4099), .ZN(n4101)
         );
  OAI21_X1 U4744 ( .B1(n4102), .B2(n4298), .A(n4101), .ZN(n4103) );
  MUX2_X1 U4745 ( .A(n3542), .B(n4342), .S(n4289), .Z(n4105) );
  OAI211_X1 U4746 ( .C1(n4426), .C2(n4242), .A(n4106), .B(n4105), .ZN(U3267)
         );
  OAI21_X1 U4747 ( .B1(n4108), .B2(n4109), .A(n4107), .ZN(n4430) );
  INV_X1 U4748 ( .A(n4109), .ZN(n4110) );
  XNOR2_X1 U4749 ( .A(n4111), .B(n4110), .ZN(n4117) );
  OR2_X1 U4750 ( .A1(n4279), .A2(n4112), .ZN(n4114) );
  NAND2_X1 U4751 ( .A1(n4149), .A2(n4275), .ZN(n4113) );
  OAI211_X1 U4752 ( .C1(n4115), .C2(n4298), .A(n4114), .B(n4113), .ZN(n4116)
         );
  AOI21_X1 U4753 ( .B1(n4117), .B2(n4281), .A(n4116), .ZN(n4348) );
  AOI22_X1 U4754 ( .A1(n4118), .A2(n4618), .B1(n4623), .B2(
        REG2_REG_22__SCAN_IN), .ZN(n4122) );
  NAND2_X1 U4755 ( .A1(n2225), .A2(n4120), .ZN(n4345) );
  NAND3_X1 U4756 ( .A1(n4346), .A2(n4608), .A3(n4345), .ZN(n4121) );
  OAI211_X1 U4757 ( .C1(n4348), .C2(n4623), .A(n4122), .B(n4121), .ZN(n4123)
         );
  INV_X1 U4758 ( .A(n4123), .ZN(n4124) );
  OAI21_X1 U4759 ( .B1(n4430), .B2(n4242), .A(n4124), .ZN(U3268) );
  XNOR2_X1 U4760 ( .A(n4125), .B(n4127), .ZN(n4435) );
  AOI21_X1 U4761 ( .B1(n4128), .B2(n4355), .A(n4119), .ZN(n4433) );
  AOI22_X1 U4762 ( .A1(n4433), .A2(n4608), .B1(n4126), .B2(n4618), .ZN(n4136)
         );
  XOR2_X1 U4763 ( .A(n4127), .B(n4091), .Z(n4133) );
  AOI22_X1 U4764 ( .A1(n4129), .A2(n4275), .B1(n4306), .B2(n4128), .ZN(n4130)
         );
  OAI21_X1 U4765 ( .B1(n4131), .B2(n4298), .A(n4130), .ZN(n4132) );
  AOI21_X1 U4766 ( .B1(n4133), .B2(n4281), .A(n4132), .ZN(n4351) );
  MUX2_X1 U4767 ( .A(n4351), .B(n4134), .S(n4623), .Z(n4135) );
  OAI211_X1 U4768 ( .C1(n4435), .C2(n4242), .A(n4136), .B(n4135), .ZN(U3269)
         );
  NAND2_X1 U4769 ( .A1(n4137), .A2(n4183), .ZN(n4180) );
  NAND2_X1 U4770 ( .A1(n4180), .A2(n4138), .ZN(n4161) );
  NAND2_X1 U4771 ( .A1(n4161), .A2(n4139), .ZN(n4141) );
  NAND2_X1 U4772 ( .A1(n4141), .A2(n4140), .ZN(n4143) );
  XNOR2_X1 U4773 ( .A(n4143), .B(n4142), .ZN(n4354) );
  INV_X1 U4774 ( .A(n4303), .ZN(n4153) );
  NOR2_X1 U4775 ( .A1(n2561), .A2(n4144), .ZN(n4146) );
  XNOR2_X1 U4776 ( .A(n4146), .B(n4145), .ZN(n4151) );
  OAI22_X1 U4777 ( .A1(n4187), .A2(n4296), .B1(n4147), .B2(n4279), .ZN(n4148)
         );
  AOI21_X1 U4778 ( .B1(n4149), .B2(n4276), .A(n4148), .ZN(n4150) );
  OAI21_X1 U4779 ( .B1(n4151), .B2(n4309), .A(n4150), .ZN(n4152) );
  AOI21_X1 U4780 ( .B1(n4354), .B2(n4153), .A(n4152), .ZN(n4358) );
  INV_X1 U4781 ( .A(n4162), .ZN(n4155) );
  NAND2_X1 U4782 ( .A1(n4155), .A2(n4154), .ZN(n4356) );
  AND3_X1 U4783 ( .A1(n4356), .A2(n4608), .A3(n4355), .ZN(n4159) );
  OAI22_X1 U4784 ( .A1(n4157), .A2(n4289), .B1(n4156), .B2(n4287), .ZN(n4158)
         );
  AOI211_X1 U4785 ( .C1(n4354), .C2(n4620), .A(n4159), .B(n4158), .ZN(n4160)
         );
  OAI21_X1 U4786 ( .B1(n4358), .B2(n4623), .A(n4160), .ZN(U3270) );
  XNOR2_X1 U4787 ( .A(n4161), .B(n4171), .ZN(n4441) );
  AOI21_X1 U4788 ( .B1(n4172), .B2(n2310), .A(n4162), .ZN(n4439) );
  AOI22_X1 U4789 ( .A1(n4439), .A2(n4608), .B1(n4163), .B2(n4618), .ZN(n4179)
         );
  OAI21_X1 U4790 ( .B1(n4164), .B2(n4166), .A(n4165), .ZN(n4182) );
  INV_X1 U4791 ( .A(n4167), .ZN(n4169) );
  OAI21_X1 U4792 ( .B1(n4182), .B2(n4169), .A(n4168), .ZN(n4170) );
  XOR2_X1 U4793 ( .A(n4171), .B(n4170), .Z(n4177) );
  AOI22_X1 U4794 ( .A1(n4173), .A2(n4275), .B1(n4172), .B2(n4306), .ZN(n4174)
         );
  OAI21_X1 U4795 ( .B1(n4175), .B2(n4298), .A(n4174), .ZN(n4176) );
  AOI21_X1 U4796 ( .B1(n4177), .B2(n4281), .A(n4176), .ZN(n4360) );
  MUX2_X1 U4797 ( .A(n4495), .B(n4360), .S(n4289), .Z(n4178) );
  OAI211_X1 U4798 ( .C1(n4441), .C2(n4242), .A(n4179), .B(n4178), .ZN(U3271)
         );
  OAI21_X1 U4799 ( .B1(n4137), .B2(n4183), .A(n4180), .ZN(n4181) );
  INV_X1 U4800 ( .A(n4181), .ZN(n4365) );
  XOR2_X1 U4801 ( .A(n4183), .B(n4182), .Z(n4189) );
  AOI22_X1 U4802 ( .A1(n4185), .A2(n4275), .B1(n4306), .B2(n4184), .ZN(n4186)
         );
  OAI21_X1 U4803 ( .B1(n4187), .B2(n4298), .A(n4186), .ZN(n4188) );
  AOI21_X1 U4804 ( .B1(n4189), .B2(n4281), .A(n4188), .ZN(n4364) );
  INV_X1 U4805 ( .A(n4364), .ZN(n4196) );
  OAI211_X1 U4806 ( .C1(n2233), .C2(n4191), .A(n4653), .B(n2310), .ZN(n4363)
         );
  NOR2_X1 U4807 ( .A1(n4363), .A2(n4192), .ZN(n4195) );
  OAI22_X1 U4808 ( .A1(n4289), .A2(n3492), .B1(n4193), .B2(n4287), .ZN(n4194)
         );
  AOI211_X1 U4809 ( .C1(n4196), .C2(n4289), .A(n4195), .B(n4194), .ZN(n4197)
         );
  OAI21_X1 U4810 ( .B1(n4365), .B2(n4242), .A(n4197), .ZN(U3272) );
  XNOR2_X1 U4811 ( .A(n4198), .B(n4201), .ZN(n4448) );
  AOI21_X1 U4812 ( .B1(n4202), .B2(n2019), .A(n2233), .ZN(n4446) );
  INV_X1 U4813 ( .A(n4199), .ZN(n4200) );
  AOI22_X1 U4814 ( .A1(n4446), .A2(n4608), .B1(n4200), .B2(n4618), .ZN(n4210)
         );
  XNOR2_X1 U4815 ( .A(n4164), .B(n4201), .ZN(n4207) );
  AOI22_X1 U4816 ( .A1(n4203), .A2(n4275), .B1(n4306), .B2(n4202), .ZN(n4204)
         );
  OAI21_X1 U4817 ( .B1(n4205), .B2(n4298), .A(n4204), .ZN(n4206) );
  AOI21_X1 U4818 ( .B1(n4207), .B2(n4281), .A(n4206), .ZN(n4443) );
  MUX2_X1 U4819 ( .A(n4208), .B(n4443), .S(n4289), .Z(n4209) );
  OAI211_X1 U4820 ( .C1(n4448), .C2(n4242), .A(n4210), .B(n4209), .ZN(U3273)
         );
  OAI21_X1 U4821 ( .B1(n4213), .B2(n2727), .A(n4212), .ZN(n4452) );
  XNOR2_X1 U4822 ( .A(n4214), .B(n2727), .ZN(n4219) );
  NAND2_X1 U4823 ( .A1(n4250), .A2(n4275), .ZN(n4216) );
  NAND2_X1 U4824 ( .A1(n4221), .A2(n4306), .ZN(n4215) );
  OAI211_X1 U4825 ( .C1(n4217), .C2(n4298), .A(n4216), .B(n4215), .ZN(n4218)
         );
  AOI21_X1 U4826 ( .B1(n4219), .B2(n4281), .A(n4218), .ZN(n4370) );
  AOI22_X1 U4827 ( .A1(n4623), .A2(REG2_REG_16__SCAN_IN), .B1(n4220), .B2(
        n4618), .ZN(n4224) );
  INV_X1 U4828 ( .A(n4237), .ZN(n4222) );
  NAND2_X1 U4829 ( .A1(n4222), .A2(n4221), .ZN(n4368) );
  NAND3_X1 U4830 ( .A1(n2019), .A2(n4608), .A3(n4368), .ZN(n4223) );
  OAI211_X1 U4831 ( .C1(n4370), .C2(n4623), .A(n4224), .B(n4223), .ZN(n4225)
         );
  INV_X1 U4832 ( .A(n4225), .ZN(n4226) );
  OAI21_X1 U4833 ( .B1(n4452), .B2(n4242), .A(n4226), .ZN(U3274) );
  XNOR2_X1 U4834 ( .A(n4227), .B(n4231), .ZN(n4459) );
  INV_X1 U4835 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4500) );
  OAI22_X1 U4836 ( .A1(n4229), .A2(n4298), .B1(n4228), .B2(n4296), .ZN(n4236)
         );
  INV_X1 U4837 ( .A(n4230), .ZN(n4234) );
  AOI21_X1 U4838 ( .B1(n4246), .B2(n4232), .A(n4231), .ZN(n4233) );
  NOR3_X1 U4839 ( .A1(n4234), .A2(n4233), .A3(n4309), .ZN(n4235) );
  AOI211_X1 U4840 ( .C1(n4306), .C2(n4238), .A(n4236), .B(n4235), .ZN(n4453)
         );
  MUX2_X1 U4841 ( .A(n4500), .B(n4453), .S(n4289), .Z(n4241) );
  AOI21_X1 U4842 ( .B1(n4238), .B2(n2043), .A(n4237), .ZN(n4456) );
  AOI22_X1 U4843 ( .A1(n4456), .A2(n4608), .B1(n4239), .B2(n4618), .ZN(n4240)
         );
  OAI211_X1 U4844 ( .C1(n4459), .C2(n4242), .A(n4241), .B(n4240), .ZN(U3275)
         );
  OAI21_X1 U4845 ( .B1(n4245), .B2(n4244), .A(n4243), .ZN(n4376) );
  INV_X1 U4846 ( .A(n4376), .ZN(n4264) );
  OAI21_X1 U4847 ( .B1(n4248), .B2(n4247), .A(n4246), .ZN(n4254) );
  AOI22_X1 U4848 ( .A1(n4250), .A2(n4276), .B1(n4275), .B2(n4249), .ZN(n4251)
         );
  OAI21_X1 U4849 ( .B1(n4252), .B2(n4279), .A(n4251), .ZN(n4253) );
  AOI21_X1 U4850 ( .B1(n4254), .B2(n4281), .A(n4253), .ZN(n4255) );
  OAI21_X1 U4851 ( .B1(n4264), .B2(n4303), .A(n4255), .ZN(n4375) );
  NAND2_X1 U4852 ( .A1(n4375), .A2(n4289), .ZN(n4263) );
  NAND2_X1 U4853 ( .A1(n4284), .A2(n4256), .ZN(n4257) );
  NAND2_X1 U4854 ( .A1(n2043), .A2(n4257), .ZN(n4463) );
  INV_X1 U4855 ( .A(n4463), .ZN(n4261) );
  INV_X1 U4856 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4259) );
  OAI22_X1 U4857 ( .A1(n4289), .A2(n4259), .B1(n4258), .B2(n4287), .ZN(n4260)
         );
  AOI21_X1 U4858 ( .B1(n4261), .B2(n4608), .A(n4260), .ZN(n4262) );
  OAI211_X1 U4859 ( .C1(n4264), .C2(n4294), .A(n4263), .B(n4262), .ZN(U3276)
         );
  NAND2_X1 U4860 ( .A1(n4266), .A2(n4265), .ZN(n4267) );
  XOR2_X1 U4861 ( .A(n4272), .B(n4267), .Z(n4379) );
  INV_X1 U4862 ( .A(n4268), .ZN(n4270) );
  OAI21_X1 U4863 ( .B1(n4271), .B2(n4270), .A(n4269), .ZN(n4273) );
  XNOR2_X1 U4864 ( .A(n4273), .B(n4272), .ZN(n4282) );
  AOI22_X1 U4865 ( .A1(n4277), .A2(n4276), .B1(n4275), .B2(n4274), .ZN(n4278)
         );
  OAI21_X1 U4866 ( .B1(n4285), .B2(n4279), .A(n4278), .ZN(n4280) );
  AOI21_X1 U4867 ( .B1(n4282), .B2(n4281), .A(n4280), .ZN(n4283) );
  OAI21_X1 U4868 ( .B1(n4379), .B2(n4303), .A(n4283), .ZN(n4380) );
  NAND2_X1 U4869 ( .A1(n4380), .A2(n4289), .ZN(n4293) );
  OAI21_X1 U4870 ( .B1(n4384), .B2(n4285), .A(n4284), .ZN(n4467) );
  INV_X1 U4871 ( .A(n4467), .ZN(n4291) );
  INV_X1 U4872 ( .A(n4286), .ZN(n4288) );
  OAI22_X1 U4873 ( .A1(n4289), .A2(n4544), .B1(n4288), .B2(n4287), .ZN(n4290)
         );
  AOI21_X1 U4874 ( .B1(n4291), .B2(n4608), .A(n4290), .ZN(n4292) );
  OAI211_X1 U4875 ( .C1(n4379), .C2(n4294), .A(n4293), .B(n4292), .ZN(U3277)
         );
  XOR2_X1 U4876 ( .A(n4295), .B(n4302), .Z(n4308) );
  OAI22_X1 U4877 ( .A1(n4299), .A2(n4298), .B1(n4297), .B2(n4296), .ZN(n4305)
         );
  INV_X1 U4878 ( .A(n4300), .ZN(n4301) );
  AOI21_X1 U4879 ( .B1(n4302), .B2(n3294), .A(n4301), .ZN(n4310) );
  NOR2_X1 U4880 ( .A1(n4310), .A2(n4303), .ZN(n4304) );
  AOI211_X1 U4881 ( .C1(n4306), .C2(n4311), .A(n4305), .B(n4304), .ZN(n4307)
         );
  OAI21_X1 U4882 ( .B1(n4309), .B2(n4308), .A(n4307), .ZN(n4391) );
  INV_X1 U4883 ( .A(n4391), .ZN(n4320) );
  INV_X1 U4884 ( .A(n4310), .ZN(n4392) );
  AND2_X1 U4885 ( .A1(n4312), .A2(n4311), .ZN(n4313) );
  OR2_X1 U4886 ( .A1(n4314), .A2(n4313), .ZN(n4477) );
  AOI22_X1 U4887 ( .A1(n4623), .A2(REG2_REG_11__SCAN_IN), .B1(n4315), .B2(
        n4618), .ZN(n4316) );
  OAI21_X1 U4888 ( .B1(n4477), .B2(n4317), .A(n4316), .ZN(n4318) );
  AOI21_X1 U4889 ( .B1(n4392), .B2(n4620), .A(n4318), .ZN(n4319) );
  OAI21_X1 U4890 ( .B1(n4320), .B2(n4623), .A(n4319), .ZN(U3279) );
  NAND2_X1 U4891 ( .A1(n4684), .A2(n4396), .ZN(n4322) );
  NAND2_X1 U4892 ( .A1(n4681), .A2(REG1_REG_31__SCAN_IN), .ZN(n4321) );
  OAI211_X1 U4893 ( .C1(n4399), .C2(n4395), .A(n4322), .B(n4321), .ZN(U3549)
         );
  INV_X1 U4894 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4325) );
  NAND2_X1 U4895 ( .A1(n4400), .A2(n4372), .ZN(n4324) );
  NAND2_X1 U4896 ( .A1(n4684), .A2(n4401), .ZN(n4323) );
  OAI211_X1 U4897 ( .C1(n4684), .C2(n4325), .A(n4324), .B(n4323), .ZN(U3548)
         );
  NAND2_X1 U4898 ( .A1(n4326), .A2(n4653), .ZN(n4327) );
  NAND2_X1 U4899 ( .A1(n4328), .A2(n4327), .ZN(n4405) );
  MUX2_X1 U4900 ( .A(REG1_REG_27__SCAN_IN), .B(n4405), .S(n4684), .Z(n4329) );
  INV_X1 U4901 ( .A(n4329), .ZN(n4330) );
  OAI21_X1 U4902 ( .B1(n4408), .B2(n4390), .A(n4330), .ZN(U3545) );
  INV_X1 U4903 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4333) );
  AOI21_X1 U4904 ( .B1(n4332), .B2(n4665), .A(n4331), .ZN(n4409) );
  MUX2_X1 U4905 ( .A(n4333), .B(n4409), .S(n4684), .Z(n4334) );
  OAI21_X1 U4906 ( .B1(n4395), .B2(n4412), .A(n4334), .ZN(U3544) );
  INV_X1 U4907 ( .A(n4335), .ZN(n4413) );
  MUX2_X1 U4908 ( .A(REG1_REG_25__SCAN_IN), .B(n4413), .S(n4684), .Z(n4336) );
  AOI21_X1 U4909 ( .B1(n4415), .B2(n4372), .A(n4336), .ZN(n4337) );
  OAI21_X1 U4910 ( .B1(n4417), .B2(n4390), .A(n4337), .ZN(U3543) );
  INV_X1 U4911 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4340) );
  AOI21_X1 U4912 ( .B1(n4339), .B2(n4665), .A(n4338), .ZN(n4418) );
  MUX2_X1 U4913 ( .A(n4340), .B(n4418), .S(n4684), .Z(n4341) );
  OAI21_X1 U4914 ( .B1(n4395), .B2(n4421), .A(n4341), .ZN(U3542) );
  INV_X1 U4915 ( .A(n4342), .ZN(n4422) );
  MUX2_X1 U4916 ( .A(REG1_REG_23__SCAN_IN), .B(n4422), .S(n4684), .Z(n4343) );
  AOI21_X1 U4917 ( .B1(n4424), .B2(n4372), .A(n4343), .ZN(n4344) );
  OAI21_X1 U4918 ( .B1(n4426), .B2(n4390), .A(n4344), .ZN(U3541) );
  NAND3_X1 U4919 ( .A1(n4346), .A2(n4653), .A3(n4345), .ZN(n4347) );
  NAND2_X1 U4920 ( .A1(n4348), .A2(n4347), .ZN(n4427) );
  MUX2_X1 U4921 ( .A(REG1_REG_22__SCAN_IN), .B(n4427), .S(n4684), .Z(n4349) );
  INV_X1 U4922 ( .A(n4349), .ZN(n4350) );
  OAI21_X1 U4923 ( .B1(n4430), .B2(n4390), .A(n4350), .ZN(U3540) );
  INV_X1 U4924 ( .A(n4351), .ZN(n4431) );
  MUX2_X1 U4925 ( .A(n4431), .B(REG1_REG_21__SCAN_IN), .S(n4681), .Z(n4352) );
  AOI21_X1 U4926 ( .B1(n4433), .B2(n4372), .A(n4352), .ZN(n4353) );
  OAI21_X1 U4927 ( .B1(n4435), .B2(n4390), .A(n4353), .ZN(U3539) );
  INV_X1 U4928 ( .A(n4354), .ZN(n4359) );
  NAND3_X1 U4929 ( .A1(n4356), .A2(n4653), .A3(n4355), .ZN(n4357) );
  OAI211_X1 U4930 ( .C1(n4359), .C2(n4648), .A(n4358), .B(n4357), .ZN(n4436)
         );
  MUX2_X1 U4931 ( .A(REG1_REG_20__SCAN_IN), .B(n4436), .S(n4684), .Z(U3538) );
  INV_X1 U4932 ( .A(n4360), .ZN(n4437) );
  MUX2_X1 U4933 ( .A(REG1_REG_19__SCAN_IN), .B(n4437), .S(n4684), .Z(n4361) );
  AOI21_X1 U4934 ( .B1(n4439), .B2(n4372), .A(n4361), .ZN(n4362) );
  OAI21_X1 U4935 ( .B1(n4390), .B2(n4441), .A(n4362), .ZN(U3537) );
  OAI211_X1 U4936 ( .C1(n4365), .C2(n4668), .A(n4364), .B(n4363), .ZN(n4442)
         );
  MUX2_X1 U4937 ( .A(REG1_REG_18__SCAN_IN), .B(n4442), .S(n4684), .Z(U3536) );
  INV_X1 U4938 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4510) );
  MUX2_X1 U4939 ( .A(n4510), .B(n4443), .S(n4684), .Z(n4367) );
  NAND2_X1 U4940 ( .A1(n4446), .A2(n4372), .ZN(n4366) );
  OAI211_X1 U4941 ( .C1(n4448), .C2(n4390), .A(n4367), .B(n4366), .ZN(U3535)
         );
  INV_X1 U4942 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4570) );
  NAND3_X1 U4943 ( .A1(n2019), .A2(n4653), .A3(n4368), .ZN(n4369) );
  AND2_X1 U4944 ( .A1(n4370), .A2(n4369), .ZN(n4449) );
  MUX2_X1 U4945 ( .A(n4570), .B(n4449), .S(n4684), .Z(n4371) );
  OAI21_X1 U4946 ( .B1(n4452), .B2(n4390), .A(n4371), .ZN(U3534) );
  INV_X1 U4947 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4516) );
  MUX2_X1 U4948 ( .A(n4516), .B(n4453), .S(n4684), .Z(n4374) );
  NAND2_X1 U4949 ( .A1(n4456), .A2(n4372), .ZN(n4373) );
  OAI211_X1 U4950 ( .C1(n4459), .C2(n4390), .A(n4374), .B(n4373), .ZN(U3533)
         );
  INV_X1 U4951 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4377) );
  AOI21_X1 U4952 ( .B1(n4658), .B2(n4376), .A(n4375), .ZN(n4460) );
  MUX2_X1 U4953 ( .A(n4377), .B(n4460), .S(n4684), .Z(n4378) );
  OAI21_X1 U4954 ( .B1(n4395), .B2(n4463), .A(n4378), .ZN(U3532) );
  INV_X1 U4955 ( .A(n4379), .ZN(n4381) );
  AOI21_X1 U4956 ( .B1(n4658), .B2(n4381), .A(n4380), .ZN(n4464) );
  MUX2_X1 U4957 ( .A(n4382), .B(n4464), .S(n4684), .Z(n4383) );
  OAI21_X1 U4958 ( .B1(n4395), .B2(n4467), .A(n4383), .ZN(U3531) );
  NOR3_X1 U4959 ( .A1(n4385), .A2(n4384), .A3(n4661), .ZN(n4386) );
  NOR2_X1 U4960 ( .A1(n4387), .A2(n4386), .ZN(n4468) );
  MUX2_X1 U4961 ( .A(n4388), .B(n4468), .S(n4684), .Z(n4389) );
  OAI21_X1 U4962 ( .B1(n4472), .B2(n4390), .A(n4389), .ZN(U3530) );
  AOI21_X1 U4963 ( .B1(n4658), .B2(n4392), .A(n4391), .ZN(n4473) );
  MUX2_X1 U4964 ( .A(n4393), .B(n4473), .S(n4684), .Z(n4394) );
  OAI21_X1 U4965 ( .B1(n4395), .B2(n4477), .A(n4394), .ZN(U3529) );
  NAND2_X1 U4966 ( .A1(n4675), .A2(n4396), .ZN(n4398) );
  NAND2_X1 U4967 ( .A1(n4673), .A2(REG0_REG_31__SCAN_IN), .ZN(n4397) );
  OAI211_X1 U4968 ( .C1(n4399), .C2(n4476), .A(n4398), .B(n4397), .ZN(U3517)
         );
  INV_X1 U4969 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4404) );
  NAND2_X1 U4970 ( .A1(n4400), .A2(n4455), .ZN(n4403) );
  NAND2_X1 U4971 ( .A1(n4675), .A2(n4401), .ZN(n4402) );
  OAI211_X1 U4972 ( .C1(n4675), .C2(n4404), .A(n4403), .B(n4402), .ZN(U3516)
         );
  MUX2_X1 U4973 ( .A(REG0_REG_27__SCAN_IN), .B(n4405), .S(n4675), .Z(n4406) );
  INV_X1 U4974 ( .A(n4406), .ZN(n4407) );
  OAI21_X1 U4975 ( .B1(n4408), .B2(n4471), .A(n4407), .ZN(U3513) );
  MUX2_X1 U4976 ( .A(n4410), .B(n4409), .S(n4675), .Z(n4411) );
  OAI21_X1 U4977 ( .B1(n4412), .B2(n4476), .A(n4411), .ZN(U3512) );
  MUX2_X1 U4978 ( .A(REG0_REG_25__SCAN_IN), .B(n4413), .S(n4675), .Z(n4414) );
  AOI21_X1 U4979 ( .B1(n4415), .B2(n4455), .A(n4414), .ZN(n4416) );
  OAI21_X1 U4980 ( .B1(n4417), .B2(n4471), .A(n4416), .ZN(U3511) );
  INV_X1 U4981 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4419) );
  MUX2_X1 U4982 ( .A(n4419), .B(n4418), .S(n4675), .Z(n4420) );
  OAI21_X1 U4983 ( .B1(n4421), .B2(n4476), .A(n4420), .ZN(U3510) );
  MUX2_X1 U4984 ( .A(REG0_REG_23__SCAN_IN), .B(n4422), .S(n4675), .Z(n4423) );
  AOI21_X1 U4985 ( .B1(n4424), .B2(n4455), .A(n4423), .ZN(n4425) );
  OAI21_X1 U4986 ( .B1(n4426), .B2(n4471), .A(n4425), .ZN(U3509) );
  MUX2_X1 U4987 ( .A(REG0_REG_22__SCAN_IN), .B(n4427), .S(n4675), .Z(n4428) );
  INV_X1 U4988 ( .A(n4428), .ZN(n4429) );
  OAI21_X1 U4989 ( .B1(n4430), .B2(n4471), .A(n4429), .ZN(U3508) );
  MUX2_X1 U4990 ( .A(n4431), .B(REG0_REG_21__SCAN_IN), .S(n4673), .Z(n4432) );
  AOI21_X1 U4991 ( .B1(n4433), .B2(n4455), .A(n4432), .ZN(n4434) );
  OAI21_X1 U4992 ( .B1(n4435), .B2(n4471), .A(n4434), .ZN(U3507) );
  MUX2_X1 U4993 ( .A(REG0_REG_20__SCAN_IN), .B(n4436), .S(n4675), .Z(U3506) );
  MUX2_X1 U4994 ( .A(REG0_REG_19__SCAN_IN), .B(n4437), .S(n4675), .Z(n4438) );
  AOI21_X1 U4995 ( .B1(n4439), .B2(n4455), .A(n4438), .ZN(n4440) );
  OAI21_X1 U4996 ( .B1(n4471), .B2(n4441), .A(n4440), .ZN(U3505) );
  MUX2_X1 U4997 ( .A(REG0_REG_18__SCAN_IN), .B(n4442), .S(n4675), .Z(U3503) );
  INV_X1 U4998 ( .A(n4443), .ZN(n4444) );
  MUX2_X1 U4999 ( .A(REG0_REG_17__SCAN_IN), .B(n4444), .S(n4675), .Z(n4445) );
  AOI21_X1 U5000 ( .B1(n4446), .B2(n4455), .A(n4445), .ZN(n4447) );
  OAI21_X1 U5001 ( .B1(n4448), .B2(n4471), .A(n4447), .ZN(U3501) );
  INV_X1 U5002 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4450) );
  MUX2_X1 U5003 ( .A(n4450), .B(n4449), .S(n4675), .Z(n4451) );
  OAI21_X1 U5004 ( .B1(n4452), .B2(n4471), .A(n4451), .ZN(U3499) );
  MUX2_X1 U5005 ( .A(n4454), .B(n4453), .S(n4675), .Z(n4458) );
  NAND2_X1 U5006 ( .A1(n4456), .A2(n4455), .ZN(n4457) );
  OAI211_X1 U5007 ( .C1(n4459), .C2(n4471), .A(n4458), .B(n4457), .ZN(U3497)
         );
  INV_X1 U5008 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4461) );
  MUX2_X1 U5009 ( .A(n4461), .B(n4460), .S(n4675), .Z(n4462) );
  OAI21_X1 U5010 ( .B1(n4463), .B2(n4476), .A(n4462), .ZN(U3495) );
  INV_X1 U5011 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4465) );
  MUX2_X1 U5012 ( .A(n4465), .B(n4464), .S(n4675), .Z(n4466) );
  OAI21_X1 U5013 ( .B1(n4467), .B2(n4476), .A(n4466), .ZN(U3493) );
  INV_X1 U5014 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4469) );
  MUX2_X1 U5015 ( .A(n4469), .B(n4468), .S(n4675), .Z(n4470) );
  OAI21_X1 U5016 ( .B1(n4472), .B2(n4471), .A(n4470), .ZN(U3491) );
  INV_X1 U5017 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4474) );
  MUX2_X1 U5018 ( .A(n4474), .B(n4473), .S(n4675), .Z(n4475) );
  OAI21_X1 U5019 ( .B1(n4477), .B2(n4476), .A(n4475), .ZN(U3489) );
  MUX2_X1 U5020 ( .A(n4478), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5021 ( .A(n4479), .B(DATAI_28_), .S(U3149), .Z(U3324) );
  MUX2_X1 U5022 ( .A(DATAI_27_), .B(n4480), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U5023 ( .A(n4481), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U5024 ( .A(n4482), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U5025 ( .A(DATAI_20_), .B(n4483), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5026 ( .A(n4484), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5027 ( .A(DATAI_14_), .B(n4512), .S(STATE_REG_SCAN_IN), .Z(U3338)
         );
  MUX2_X1 U5028 ( .A(n4485), .B(DATAI_12_), .S(U3149), .Z(U3340) );
  MUX2_X1 U5029 ( .A(n4486), .B(DATAI_11_), .S(U3149), .Z(U3341) );
  MUX2_X1 U5030 ( .A(n4487), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U5031 ( .A(n4488), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U5032 ( .A(n4489), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5033 ( .A(n4490), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5034 ( .A(n4491), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5035 ( .A(DATAI_4_), .B(n4529), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5036 ( .A(DATAI_3_), .B(n4492), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U5037 ( .A(DATAI_2_), .B(n4493), .S(STATE_REG_SCAN_IN), .Z(U3350) );
  MUX2_X1 U5038 ( .A(n4494), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U5039 ( .A(n4495), .B(REG2_REG_19__SCAN_IN), .S(n2865), .Z(n4508) );
  NAND2_X1 U5040 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4633), .ZN(n4506) );
  OAI21_X1 U5041 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4633), .A(n4506), .ZN(n4599) );
  INV_X1 U5042 ( .A(n4496), .ZN(n4497) );
  NAND2_X1 U5043 ( .A1(n4497), .A2(n4512), .ZN(n4498) );
  INV_X1 U5044 ( .A(n4558), .ZN(n4640) );
  AOI22_X1 U5045 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4640), .B1(n4558), .B2(
        n4500), .ZN(n4551) );
  AND2_X1 U5046 ( .A1(n4558), .A2(REG2_REG_15__SCAN_IN), .ZN(n4501) );
  INV_X1 U5047 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4567) );
  NAND2_X1 U5048 ( .A1(n4502), .A2(n4638), .ZN(n4503) );
  NOR2_X1 U5049 ( .A1(n4635), .A2(REG2_REG_17__SCAN_IN), .ZN(n4504) );
  AOI21_X1 U5050 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4635), .A(n4504), .ZN(n4579) );
  OR2_X1 U5051 ( .A1(n4635), .A2(REG2_REG_17__SCAN_IN), .ZN(n4505) );
  INV_X1 U5052 ( .A(n4506), .ZN(n4507) );
  AOI22_X1 U5053 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4603), .B1(n4633), .B2(
        n4509), .ZN(n4593) );
  AOI22_X1 U5054 ( .A1(n4635), .A2(REG1_REG_17__SCAN_IN), .B1(n4510), .B2(
        n4589), .ZN(n4582) );
  INV_X1 U5055 ( .A(n4511), .ZN(n4513) );
  AOI22_X1 U5056 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4640), .B1(n4558), .B2(
        n4516), .ZN(n4554) );
  NAND2_X1 U5057 ( .A1(n4517), .A2(n4638), .ZN(n4518) );
  XNOR2_X1 U5058 ( .A(n2865), .B(REG1_REG_19__SCAN_IN), .ZN(n4519) );
  AOI21_X1 U5059 ( .B1(n4595), .B2(ADDR_REG_19__SCAN_IN), .A(n4520), .ZN(n4521) );
  OAI21_X1 U5060 ( .B1(n4604), .B2(n2865), .A(n4521), .ZN(n4522) );
  INV_X1 U5061 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4524) );
  XNOR2_X1 U5062 ( .A(n4525), .B(n4524), .ZN(n4526) );
  NAND2_X1 U5063 ( .A1(n4584), .A2(n4526), .ZN(n4535) );
  XNOR2_X1 U5064 ( .A(n4527), .B(n2135), .ZN(n4528) );
  NAND2_X1 U5065 ( .A1(n4586), .A2(n4528), .ZN(n4534) );
  NAND2_X1 U5066 ( .A1(n4559), .A2(n4529), .ZN(n4533) );
  INV_X1 U5067 ( .A(n4530), .ZN(n4531) );
  AOI21_X1 U5068 ( .B1(n4595), .B2(ADDR_REG_4__SCAN_IN), .A(n4531), .ZN(n4532)
         );
  AND4_X1 U5069 ( .A1(n4535), .A2(n4534), .A3(n4533), .A4(n4532), .ZN(n4537)
         );
  NAND2_X1 U5070 ( .A1(n4537), .A2(n4536), .ZN(U3244) );
  AOI211_X1 U5071 ( .C1(n4540), .C2(n4539), .A(n4538), .B(n4590), .ZN(n4542)
         );
  AOI211_X1 U5072 ( .C1(n4595), .C2(ADDR_REG_13__SCAN_IN), .A(n4542), .B(n4541), .ZN(n4549) );
  AOI21_X1 U5073 ( .B1(n4544), .B2(n4642), .A(n4543), .ZN(n4547) );
  AOI21_X1 U5074 ( .B1(n4547), .B2(n4546), .A(n4596), .ZN(n4545) );
  OAI21_X1 U5075 ( .B1(n4547), .B2(n4546), .A(n4545), .ZN(n4548) );
  OAI211_X1 U5076 ( .C1(n4604), .C2(n4642), .A(n4549), .B(n4548), .ZN(U3253)
         );
  AOI211_X1 U5077 ( .C1(n4552), .C2(n4551), .A(n4550), .B(n4596), .ZN(n4557)
         );
  AOI211_X1 U5078 ( .C1(n4555), .C2(n4554), .A(n4553), .B(n4590), .ZN(n4556)
         );
  AOI211_X1 U5079 ( .C1(n4559), .C2(n4558), .A(n4557), .B(n4556), .ZN(n4561)
         );
  OAI211_X1 U5080 ( .C1(n4563), .C2(n4562), .A(n4561), .B(n4560), .ZN(U3255)
         );
  INV_X1 U5081 ( .A(n4564), .ZN(n4565) );
  AOI21_X1 U5082 ( .B1(n4595), .B2(ADDR_REG_16__SCAN_IN), .A(n4565), .ZN(n4575) );
  OAI21_X1 U5083 ( .B1(n4568), .B2(n4567), .A(n4566), .ZN(n4573) );
  OAI21_X1 U5084 ( .B1(n4571), .B2(n4570), .A(n4569), .ZN(n4572) );
  AOI22_X1 U5085 ( .A1(n4586), .A2(n4573), .B1(n4584), .B2(n4572), .ZN(n4574)
         );
  OAI211_X1 U5086 ( .C1(n4638), .C2(n4604), .A(n4575), .B(n4574), .ZN(U3256)
         );
  AOI21_X1 U5087 ( .B1(n4595), .B2(ADDR_REG_17__SCAN_IN), .A(n4576), .ZN(n4588) );
  OAI21_X1 U5088 ( .B1(n4579), .B2(n4578), .A(n4577), .ZN(n4585) );
  OAI21_X1 U5089 ( .B1(n4582), .B2(n4581), .A(n4580), .ZN(n4583) );
  AOI22_X1 U5090 ( .A1(n4586), .A2(n4585), .B1(n4584), .B2(n4583), .ZN(n4587)
         );
  OAI211_X1 U5091 ( .C1(n4589), .C2(n4604), .A(n4588), .B(n4587), .ZN(U3257)
         );
  INV_X1 U5092 ( .A(n4600), .ZN(n4601) );
  OAI211_X1 U5093 ( .C1(n4604), .C2(n4603), .A(n4602), .B(n4601), .ZN(U3258)
         );
  AOI22_X1 U5094 ( .A1(REG2_REG_2__SCAN_IN), .A2(n4623), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4618), .ZN(n4611) );
  INV_X1 U5095 ( .A(n4605), .ZN(n4609) );
  INV_X1 U5096 ( .A(n4606), .ZN(n4607) );
  AOI22_X1 U5097 ( .A1(n4609), .A2(n4620), .B1(n4608), .B2(n4607), .ZN(n4610)
         );
  OAI211_X1 U5098 ( .C1(n4623), .C2(n4612), .A(n4611), .B(n4610), .ZN(U3288)
         );
  INV_X1 U5099 ( .A(n4613), .ZN(n4616) );
  INV_X1 U5100 ( .A(n4614), .ZN(n4615) );
  AOI21_X1 U5101 ( .B1(n4617), .B2(n4616), .A(n4615), .ZN(n4622) );
  AOI22_X1 U5102 ( .A1(n4620), .A2(n4619), .B1(REG3_REG_0__SCAN_IN), .B2(n4618), .ZN(n4621) );
  OAI221_X1 U5103 ( .B1(n4623), .B2(n4622), .C1(n4289), .C2(n2770), .A(n4621), 
        .ZN(U3290) );
  AND2_X1 U5104 ( .A1(D_REG_31__SCAN_IN), .A2(n4628), .ZN(U3291) );
  AND2_X1 U5105 ( .A1(D_REG_30__SCAN_IN), .A2(n4628), .ZN(U3292) );
  AND2_X1 U5106 ( .A1(D_REG_29__SCAN_IN), .A2(n4628), .ZN(U3293) );
  AND2_X1 U5107 ( .A1(D_REG_28__SCAN_IN), .A2(n4628), .ZN(U3294) );
  AND2_X1 U5108 ( .A1(D_REG_27__SCAN_IN), .A2(n4628), .ZN(U3295) );
  INV_X1 U5109 ( .A(n4628), .ZN(n4630) );
  NOR2_X1 U5110 ( .A1(n4630), .A2(n4624), .ZN(U3296) );
  AND2_X1 U5111 ( .A1(D_REG_25__SCAN_IN), .A2(n4628), .ZN(U3297) );
  AND2_X1 U5112 ( .A1(D_REG_24__SCAN_IN), .A2(n4628), .ZN(U3298) );
  NOR2_X1 U5113 ( .A1(n4630), .A2(n4625), .ZN(U3299) );
  AND2_X1 U5114 ( .A1(D_REG_22__SCAN_IN), .A2(n4628), .ZN(U3300) );
  NOR2_X1 U5115 ( .A1(n4630), .A2(n4626), .ZN(U3301) );
  AND2_X1 U5116 ( .A1(D_REG_20__SCAN_IN), .A2(n4628), .ZN(U3302) );
  AND2_X1 U5117 ( .A1(D_REG_19__SCAN_IN), .A2(n4628), .ZN(U3303) );
  AND2_X1 U5118 ( .A1(D_REG_18__SCAN_IN), .A2(n4628), .ZN(U3304) );
  AND2_X1 U5119 ( .A1(D_REG_17__SCAN_IN), .A2(n4628), .ZN(U3305) );
  AND2_X1 U5120 ( .A1(D_REG_16__SCAN_IN), .A2(n4628), .ZN(U3306) );
  AND2_X1 U5121 ( .A1(D_REG_15__SCAN_IN), .A2(n4628), .ZN(U3307) );
  AND2_X1 U5122 ( .A1(D_REG_14__SCAN_IN), .A2(n4628), .ZN(U3308) );
  AND2_X1 U5123 ( .A1(D_REG_13__SCAN_IN), .A2(n4628), .ZN(U3309) );
  AND2_X1 U5124 ( .A1(D_REG_12__SCAN_IN), .A2(n4628), .ZN(U3310) );
  AND2_X1 U5125 ( .A1(D_REG_11__SCAN_IN), .A2(n4628), .ZN(U3311) );
  AND2_X1 U5126 ( .A1(D_REG_10__SCAN_IN), .A2(n4628), .ZN(U3312) );
  AND2_X1 U5127 ( .A1(D_REG_9__SCAN_IN), .A2(n4628), .ZN(U3313) );
  AND2_X1 U5128 ( .A1(D_REG_8__SCAN_IN), .A2(n4628), .ZN(U3314) );
  AND2_X1 U5129 ( .A1(D_REG_7__SCAN_IN), .A2(n4628), .ZN(U3315) );
  NOR2_X1 U5130 ( .A1(n4630), .A2(n4627), .ZN(U3316) );
  AND2_X1 U5131 ( .A1(D_REG_5__SCAN_IN), .A2(n4628), .ZN(U3317) );
  AND2_X1 U5132 ( .A1(D_REG_4__SCAN_IN), .A2(n4628), .ZN(U3318) );
  AND2_X1 U5133 ( .A1(D_REG_3__SCAN_IN), .A2(n4628), .ZN(U3319) );
  NOR2_X1 U5134 ( .A1(n4630), .A2(n4629), .ZN(U3320) );
  OAI21_X1 U5135 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4631), .ZN(
        n4632) );
  INV_X1 U5136 ( .A(n4632), .ZN(U3329) );
  OAI22_X1 U5137 ( .A1(U3149), .A2(n4633), .B1(DATAI_18_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4634) );
  INV_X1 U5138 ( .A(n4634), .ZN(U3334) );
  OAI22_X1 U5139 ( .A1(U3149), .A2(n4635), .B1(DATAI_17_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4636) );
  INV_X1 U5140 ( .A(n4636), .ZN(U3335) );
  AOI22_X1 U5141 ( .A1(STATE_REG_SCAN_IN), .A2(n4638), .B1(n4637), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5142 ( .A(DATAI_15_), .ZN(n4639) );
  AOI22_X1 U5143 ( .A1(STATE_REG_SCAN_IN), .A2(n4640), .B1(n4639), .B2(U3149), 
        .ZN(U3337) );
  AOI22_X1 U5144 ( .A1(STATE_REG_SCAN_IN), .A2(n4642), .B1(n4641), .B2(U3149), 
        .ZN(U3339) );
  OAI22_X1 U5145 ( .A1(U3149), .A2(IR_REG_0__SCAN_IN), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4643) );
  INV_X1 U5146 ( .A(n4643), .ZN(U3352) );
  INV_X1 U5147 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4644) );
  AOI22_X1 U5148 ( .A1(n4675), .A2(n4645), .B1(n4644), .B2(n4673), .ZN(U3467)
         );
  INV_X1 U5149 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4646) );
  AOI22_X1 U5150 ( .A1(n4675), .A2(n4647), .B1(n4646), .B2(n4673), .ZN(U3469)
         );
  NOR2_X1 U5151 ( .A1(n4649), .A2(n4648), .ZN(n4651) );
  AOI211_X1 U5152 ( .C1(n4653), .C2(n4652), .A(n4651), .B(n4650), .ZN(n4677)
         );
  INV_X1 U5153 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4654) );
  AOI22_X1 U5154 ( .A1(n4675), .A2(n4677), .B1(n4654), .B2(n4673), .ZN(U3473)
         );
  INV_X1 U5155 ( .A(n4655), .ZN(n4656) );
  AOI211_X1 U5156 ( .C1(n4659), .C2(n4658), .A(n4657), .B(n4656), .ZN(n4678)
         );
  INV_X1 U5157 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4660) );
  AOI22_X1 U5158 ( .A1(n4675), .A2(n4678), .B1(n4660), .B2(n4673), .ZN(U3475)
         );
  NOR2_X1 U5159 ( .A1(n4662), .A2(n4661), .ZN(n4664) );
  AOI211_X1 U5160 ( .C1(n4666), .C2(n4665), .A(n4664), .B(n4663), .ZN(n4680)
         );
  INV_X1 U5161 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4667) );
  AOI22_X1 U5162 ( .A1(n4675), .A2(n4680), .B1(n4667), .B2(n4673), .ZN(U3477)
         );
  NOR2_X1 U5163 ( .A1(n4669), .A2(n4668), .ZN(n4672) );
  AOI211_X1 U5164 ( .C1(n4672), .C2(n3143), .A(n4671), .B(n4670), .ZN(n4683)
         );
  INV_X1 U5165 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4674) );
  AOI22_X1 U5166 ( .A1(n4675), .A2(n4683), .B1(n4674), .B2(n4673), .ZN(U3481)
         );
  INV_X1 U5167 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4676) );
  AOI22_X1 U5168 ( .A1(n4684), .A2(n4677), .B1(n4676), .B2(n4681), .ZN(U3521)
         );
  AOI22_X1 U5169 ( .A1(n4684), .A2(n4678), .B1(n4524), .B2(n4681), .ZN(U3522)
         );
  AOI22_X1 U5170 ( .A1(n4684), .A2(n4680), .B1(n4679), .B2(n4681), .ZN(U3523)
         );
  AOI22_X1 U5171 ( .A1(n4684), .A2(n4683), .B1(n4682), .B2(n4681), .ZN(U3525)
         );
  CLKBUF_X1 U2252 ( .A(n2936), .Z(n3399) );
  CLKBUF_X1 U2427 ( .A(n2432), .Z(n2656) );
endmodule

